* SPICE3 file created from NOR2X1.ext - technology: sky130A

.subckt NOR2X1 Y A B VPB VNB
X0 a_198_181# a_164_908# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9366e+12p ps=1.294e+07u w=3e+06u l=150000u
X1 a_131_1005# a_164_908# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u M=2
X2 a_131_1005# a_343_383# a_198_181# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X3 a_198_181# a_343_383# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
.ends
