* SPICE3 file created from TIEHI.ext - technology: sky130A

.subckt TIEHI Y VDD GND
X0 VDD a_121_383 Y VDD pshort w=2 l=0.15 M=2
X1 a_121_383 a_121_383 GND GND nshort w=3 l=0.15
.ends
