// File: BUFX1.spi.BUFX1.pxi
// Created: Tue Oct 15 15:45:35 2024
// 
simulator lang=spectre
x_PM_BUFX1\%GND ( GND N_GND_c_10_p N_GND_c_32_p N_GND_c_46_p N_GND_c_4_p \
 N_GND_c_25_p N_GND_c_1_p N_GND_c_2_p N_GND_c_3_p N_GND_M0_noxref_s \
 N_GND_M1_noxref_s )  PM_BUFX1\%GND
x_PM_BUFX1\%VDD ( VDD N_VDD_c_81_p N_VDD_c_65_p N_VDD_c_73_p N_VDD_c_61_n \
 N_VDD_c_62_n N_VDD_c_63_n N_VDD_M2_noxref_s N_VDD_M3_noxref_d \
 N_VDD_M4_noxref_s N_VDD_M5_noxref_d )  PM_BUFX1\%VDD
x_PM_BUFX1\%noxref_3 ( N_noxref_3_c_108_n N_noxref_3_c_112_n \
 N_noxref_3_c_114_n N_noxref_3_c_184_p N_noxref_3_c_142_n N_noxref_3_c_144_n \
 N_noxref_3_c_117_n N_noxref_3_c_120_n N_noxref_3_M1_noxref_g \
 N_noxref_3_M4_noxref_g N_noxref_3_M5_noxref_g N_noxref_3_c_125_n \
 N_noxref_3_c_197_p N_noxref_3_c_198_p N_noxref_3_c_127_n N_noxref_3_c_155_n \
 N_noxref_3_c_156_n N_noxref_3_c_128_n N_noxref_3_c_190_p N_noxref_3_c_129_n \
 N_noxref_3_c_131_n N_noxref_3_c_132_n N_noxref_3_M0_noxref_d \
 N_noxref_3_M2_noxref_d )  PM_BUFX1\%noxref_3
x_PM_BUFX1\%A ( A A A A A A A N_A_c_210_n N_A_M0_noxref_g N_A_M2_noxref_g \
 N_A_M3_noxref_g N_A_c_215_n N_A_c_244_n N_A_c_245_n N_A_c_217_n N_A_c_233_n \
 N_A_c_234_n N_A_c_218_n N_A_c_252_n N_A_c_219_n N_A_c_221_n N_A_c_222_n )  \
 PM_BUFX1\%A
x_PM_BUFX1\%Y ( Y Y Y Y Y Y Y N_Y_c_259_n N_Y_c_282_n N_Y_c_269_n N_Y_c_271_n \
 N_Y_M1_noxref_d N_Y_M4_noxref_d )  PM_BUFX1\%Y
cc_1 ( N_GND_c_1_p N_VDD_c_61_n ) capacitor c=0.00989031f //x=4.07 //y=0 \
 //x2=4.07 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_62_n ) capacitor c=0.00989031f //x=0.63 //y=0 \
 //x2=0.74 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_63_n ) capacitor c=0.00962895f //x=2.22 //y=0 \
 //x2=2.22 //y2=7.4
cc_4 ( N_GND_c_4_p N_noxref_3_c_108_n ) capacitor c=2.8021e-19 //x=3.25 \
 //y=0.535 //x2=2.845 //y2=2.59
cc_5 ( N_GND_c_3_p N_noxref_3_c_108_n ) capacitor c=0.0424932f //x=2.22 //y=0 \
 //x2=2.845 //y2=2.59
cc_6 ( N_GND_M0_noxref_s N_noxref_3_c_108_n ) capacitor c=0.00261527f \
 //x=0.495 //y=0.37 //x2=2.845 //y2=2.59
cc_7 ( N_GND_M1_noxref_s N_noxref_3_c_108_n ) capacitor c=0.00380483f \
 //x=2.715 //y=0.37 //x2=2.845 //y2=2.59
cc_8 ( N_GND_c_3_p N_noxref_3_c_112_n ) capacitor c=9.11674e-19 //x=2.22 //y=0 \
 //x2=1.595 //y2=2.59
cc_9 ( N_GND_M0_noxref_s N_noxref_3_c_112_n ) capacitor c=0.00152335f \
 //x=0.495 //y=0.37 //x2=1.595 //y2=2.59
cc_10 ( N_GND_c_10_p N_noxref_3_c_114_n ) capacitor c=0.00180485f //x=4.07 \
 //y=0 //x2=1.395 //y2=2.08
cc_11 ( N_GND_c_3_p N_noxref_3_c_114_n ) capacitor c=0.0266238f //x=2.22 //y=0 \
 //x2=1.395 //y2=2.08
cc_12 ( N_GND_M0_noxref_s N_noxref_3_c_114_n ) capacitor c=0.00950196f \
 //x=0.495 //y=0.37 //x2=1.395 //y2=2.08
cc_13 ( N_GND_c_2_p N_noxref_3_c_117_n ) capacitor c=9.71e-19 //x=0.63 //y=0 \
 //x2=1.48 //y2=2.59
cc_14 ( N_GND_c_3_p N_noxref_3_c_117_n ) capacitor c=5.56859e-19 //x=2.22 \
 //y=0 //x2=1.48 //y2=2.59
cc_15 ( N_GND_M0_noxref_s N_noxref_3_c_117_n ) capacitor c=2.30929e-19 \
 //x=0.495 //y=0.37 //x2=1.48 //y2=2.59
cc_16 ( N_GND_c_10_p N_noxref_3_c_120_n ) capacitor c=0.00203213f //x=4.07 \
 //y=0 //x2=2.96 //y2=2.085
cc_17 ( N_GND_c_4_p N_noxref_3_c_120_n ) capacitor c=7.79915e-19 //x=3.25 \
 //y=0.535 //x2=2.96 //y2=2.085
cc_18 ( N_GND_c_1_p N_noxref_3_c_120_n ) capacitor c=0.00135052f //x=4.07 \
 //y=0 //x2=2.96 //y2=2.085
cc_19 ( N_GND_c_3_p N_noxref_3_c_120_n ) capacitor c=0.0264037f //x=2.22 //y=0 \
 //x2=2.96 //y2=2.085
cc_20 ( N_GND_M1_noxref_s N_noxref_3_c_120_n ) capacitor c=0.0105356f \
 //x=2.715 //y=0.37 //x2=2.96 //y2=2.085
cc_21 ( N_GND_c_4_p N_noxref_3_c_125_n ) capacitor c=0.0121126f //x=3.25 \
 //y=0.535 //x2=3.07 //y2=0.91
cc_22 ( N_GND_M1_noxref_s N_noxref_3_c_125_n ) capacitor c=0.0315727f \
 //x=2.715 //y=0.37 //x2=3.07 //y2=0.91
cc_23 ( N_GND_c_3_p N_noxref_3_c_127_n ) capacitor c=0.0038551f //x=2.22 //y=0 \
 //x2=3.07 //y2=1.92
cc_24 ( N_GND_M1_noxref_s N_noxref_3_c_128_n ) capacitor c=0.00483274f \
 //x=2.715 //y=0.37 //x2=3.445 //y2=0.755
cc_25 ( N_GND_c_25_p N_noxref_3_c_129_n ) capacitor c=0.0118602f //x=3.735 \
 //y=0.535 //x2=3.6 //y2=0.91
cc_26 ( N_GND_M1_noxref_s N_noxref_3_c_129_n ) capacitor c=0.0143355f \
 //x=2.715 //y=0.37 //x2=3.6 //y2=0.91
cc_27 ( N_GND_M1_noxref_s N_noxref_3_c_131_n ) capacitor c=0.0074042f \
 //x=2.715 //y=0.37 //x2=3.6 //y2=1.255
cc_28 ( N_GND_c_4_p N_noxref_3_c_132_n ) capacitor c=2.1838e-19 //x=3.25 \
 //y=0.535 //x2=2.96 //y2=2.085
cc_29 ( N_GND_c_3_p N_noxref_3_c_132_n ) capacitor c=0.0108179f //x=2.22 //y=0 \
 //x2=2.96 //y2=2.085
cc_30 ( N_GND_M1_noxref_s N_noxref_3_c_132_n ) capacitor c=0.00652238f \
 //x=2.715 //y=0.37 //x2=2.96 //y2=2.085
cc_31 ( N_GND_c_10_p N_noxref_3_M0_noxref_d ) capacitor c=0.00194883f //x=4.07 \
 //y=0 //x2=0.925 //y2=0.91
cc_32 ( N_GND_c_32_p N_noxref_3_M0_noxref_d ) capacitor c=0.0146043f //x=1.03 \
 //y=0.535 //x2=0.925 //y2=0.91
cc_33 ( N_GND_c_1_p N_noxref_3_M0_noxref_d ) capacitor c=2.29264e-19 //x=4.07 \
 //y=0 //x2=0.925 //y2=0.91
cc_34 ( N_GND_c_2_p N_noxref_3_M0_noxref_d ) capacitor c=0.0094373f //x=0.63 \
 //y=0 //x2=0.925 //y2=0.91
cc_35 ( N_GND_c_3_p N_noxref_3_M0_noxref_d ) capacitor c=0.00945919f //x=2.22 \
 //y=0 //x2=0.925 //y2=0.91
cc_36 ( N_GND_M0_noxref_s N_noxref_3_M0_noxref_d ) capacitor c=0.076995f \
 //x=0.495 //y=0.37 //x2=0.925 //y2=0.91
cc_37 ( N_GND_c_10_p N_A_c_210_n ) capacitor c=0.00203213f //x=4.07 //y=0 \
 //x2=0.74 //y2=2.085
cc_38 ( N_GND_c_32_p N_A_c_210_n ) capacitor c=8.01092e-19 //x=1.03 //y=0.535 \
 //x2=0.74 //y2=2.085
cc_39 ( N_GND_c_2_p N_A_c_210_n ) capacitor c=0.028767f //x=0.63 //y=0 \
 //x2=0.74 //y2=2.085
cc_40 ( N_GND_c_3_p N_A_c_210_n ) capacitor c=0.00133096f //x=2.22 //y=0 \
 //x2=0.74 //y2=2.085
cc_41 ( N_GND_M0_noxref_s N_A_c_210_n ) capacitor c=0.0107239f //x=0.495 \
 //y=0.37 //x2=0.74 //y2=2.085
cc_42 ( N_GND_c_32_p N_A_c_215_n ) capacitor c=0.0120496f //x=1.03 //y=0.535 \
 //x2=0.85 //y2=0.91
cc_43 ( N_GND_M0_noxref_s N_A_c_215_n ) capacitor c=0.0315727f //x=0.495 \
 //y=0.37 //x2=0.85 //y2=0.91
cc_44 ( N_GND_c_2_p N_A_c_217_n ) capacitor c=0.0124051f //x=0.63 //y=0 \
 //x2=0.85 //y2=1.92
cc_45 ( N_GND_M0_noxref_s N_A_c_218_n ) capacitor c=0.00483274f //x=0.495 \
 //y=0.37 //x2=1.225 //y2=0.755
cc_46 ( N_GND_c_46_p N_A_c_219_n ) capacitor c=0.0118602f //x=1.515 //y=0.535 \
 //x2=1.38 //y2=0.91
cc_47 ( N_GND_M0_noxref_s N_A_c_219_n ) capacitor c=0.0143355f //x=0.495 \
 //y=0.37 //x2=1.38 //y2=0.91
cc_48 ( N_GND_M0_noxref_s N_A_c_221_n ) capacitor c=0.0074042f //x=0.495 \
 //y=0.37 //x2=1.38 //y2=1.255
cc_49 ( N_GND_c_32_p N_A_c_222_n ) capacitor c=2.1838e-19 //x=1.03 //y=0.535 \
 //x2=0.74 //y2=2.085
cc_50 ( N_GND_c_2_p N_A_c_222_n ) capacitor c=0.0108179f //x=0.63 //y=0 \
 //x2=0.74 //y2=2.085
cc_51 ( N_GND_M0_noxref_s N_A_c_222_n ) capacitor c=0.00650244f //x=0.495 \
 //y=0.37 //x2=0.74 //y2=2.085
cc_52 ( N_GND_c_3_p Y ) capacitor c=9.57726e-19 //x=2.22 //y=0 //x2=3.7 \
 //y2=2.22
cc_53 ( N_GND_c_10_p N_Y_c_259_n ) capacitor c=0.0021242f //x=4.07 //y=0 \
 //x2=3.615 //y2=2.08
cc_54 ( N_GND_c_1_p N_Y_c_259_n ) capacitor c=0.029556f //x=4.07 //y=0 \
 //x2=3.615 //y2=2.08
cc_55 ( N_GND_M1_noxref_s N_Y_c_259_n ) capacitor c=0.00999304f //x=2.715 \
 //y=0.37 //x2=3.615 //y2=2.08
cc_56 ( N_GND_c_10_p N_Y_M1_noxref_d ) capacitor c=0.00194883f //x=4.07 //y=0 \
 //x2=3.145 //y2=0.91
cc_57 ( N_GND_c_4_p N_Y_M1_noxref_d ) capacitor c=0.0146043f //x=3.25 \
 //y=0.535 //x2=3.145 //y2=0.91
cc_58 ( N_GND_c_1_p N_Y_M1_noxref_d ) capacitor c=0.00973758f //x=4.07 //y=0 \
 //x2=3.145 //y2=0.91
cc_59 ( N_GND_c_3_p N_Y_M1_noxref_d ) capacitor c=0.00924905f //x=2.22 //y=0 \
 //x2=3.145 //y2=0.91
cc_60 ( N_GND_M1_noxref_s N_Y_M1_noxref_d ) capacitor c=0.076995f //x=2.715 \
 //y=0.37 //x2=3.145 //y2=0.91
cc_61 ( N_VDD_c_63_n N_noxref_3_c_108_n ) capacitor c=0.00382812f //x=2.22 \
 //y=7.4 //x2=2.845 //y2=2.59
cc_62 ( N_VDD_c_65_p N_noxref_3_c_142_n ) capacitor c=8.92854e-19 //x=1.47 \
 //y=7.4 //x2=1.395 //y2=4.58
cc_63 ( N_VDD_M3_noxref_d N_noxref_3_c_142_n ) capacitor c=0.00644908f \
 //x=1.41 //y=5.02 //x2=1.395 //y2=4.58
cc_64 ( N_VDD_c_62_n N_noxref_3_c_144_n ) capacitor c=0.0179238f //x=0.74 \
 //y=7.4 //x2=1.2 //y2=4.58
cc_65 ( N_VDD_c_62_n N_noxref_3_c_117_n ) capacitor c=4.80934e-19 //x=0.74 \
 //y=7.4 //x2=1.48 //y2=2.59
cc_66 ( N_VDD_c_63_n N_noxref_3_c_117_n ) capacitor c=0.0232484f //x=2.22 \
 //y=7.4 //x2=1.48 //y2=2.59
cc_67 ( N_VDD_c_61_n N_noxref_3_c_120_n ) capacitor c=0.00144809f //x=4.07 \
 //y=7.4 //x2=2.96 //y2=2.085
cc_68 ( N_VDD_c_63_n N_noxref_3_c_120_n ) capacitor c=0.0272885f //x=2.22 \
 //y=7.4 //x2=2.96 //y2=2.085
cc_69 ( N_VDD_M4_noxref_s N_noxref_3_c_120_n ) capacitor c=0.00938034f \
 //x=2.76 //y=5.02 //x2=2.96 //y2=2.085
cc_70 ( N_VDD_c_73_p N_noxref_3_M4_noxref_g ) capacitor c=0.00748034f //x=3.69 \
 //y=7.4 //x2=3.115 //y2=6.02
cc_71 ( N_VDD_c_63_n N_noxref_3_M4_noxref_g ) capacitor c=0.00653241f //x=2.22 \
 //y=7.4 //x2=3.115 //y2=6.02
cc_72 ( N_VDD_M4_noxref_s N_noxref_3_M4_noxref_g ) capacitor c=0.0528676f \
 //x=2.76 //y=5.02 //x2=3.115 //y2=6.02
cc_73 ( N_VDD_c_73_p N_noxref_3_M5_noxref_g ) capacitor c=0.00697478f //x=3.69 \
 //y=7.4 //x2=3.555 //y2=6.02
cc_74 ( N_VDD_M5_noxref_d N_noxref_3_M5_noxref_g ) capacitor c=0.0528676f \
 //x=3.63 //y=5.02 //x2=3.555 //y2=6.02
cc_75 ( N_VDD_c_61_n N_noxref_3_c_155_n ) capacitor c=0.0287802f //x=4.07 \
 //y=7.4 //x2=3.48 //y2=4.79
cc_76 ( N_VDD_c_63_n N_noxref_3_c_156_n ) capacitor c=0.011132f //x=2.22 \
 //y=7.4 //x2=3.19 //y2=4.79
cc_77 ( N_VDD_M4_noxref_s N_noxref_3_c_156_n ) capacitor c=0.00665831f \
 //x=2.76 //y=5.02 //x2=3.19 //y2=4.79
cc_78 ( N_VDD_c_81_p N_noxref_3_M2_noxref_d ) capacitor c=0.00722811f //x=4.07 \
 //y=7.4 //x2=0.97 //y2=5.02
cc_79 ( N_VDD_c_65_p N_noxref_3_M2_noxref_d ) capacitor c=0.0139004f //x=1.47 \
 //y=7.4 //x2=0.97 //y2=5.02
cc_80 ( N_VDD_c_61_n N_noxref_3_M2_noxref_d ) capacitor c=0.00135976f //x=4.07 \
 //y=7.4 //x2=0.97 //y2=5.02
cc_81 ( N_VDD_c_63_n N_noxref_3_M2_noxref_d ) capacitor c=0.0201812f //x=2.22 \
 //y=7.4 //x2=0.97 //y2=5.02
cc_82 ( N_VDD_M2_noxref_s N_noxref_3_M2_noxref_d ) capacitor c=0.0843065f \
 //x=0.54 //y=5.02 //x2=0.97 //y2=5.02
cc_83 ( N_VDD_M3_noxref_d N_noxref_3_M2_noxref_d ) capacitor c=0.0832641f \
 //x=1.41 //y=5.02 //x2=0.97 //y2=5.02
cc_84 ( N_VDD_c_62_n N_A_c_210_n ) capacitor c=0.0276175f //x=0.74 //y=7.4 \
 //x2=0.74 //y2=2.085
cc_85 ( N_VDD_c_63_n N_A_c_210_n ) capacitor c=0.00143749f //x=2.22 //y=7.4 \
 //x2=0.74 //y2=2.085
cc_86 ( N_VDD_M2_noxref_s N_A_c_210_n ) capacitor c=0.00938034f //x=0.54 \
 //y=5.02 //x2=0.74 //y2=2.085
cc_87 ( N_VDD_c_65_p N_A_M2_noxref_g ) capacitor c=0.00748034f //x=1.47 \
 //y=7.4 //x2=0.895 //y2=6.02
cc_88 ( N_VDD_c_62_n N_A_M2_noxref_g ) capacitor c=0.0241676f //x=0.74 //y=7.4 \
 //x2=0.895 //y2=6.02
cc_89 ( N_VDD_M2_noxref_s N_A_M2_noxref_g ) capacitor c=0.0528676f //x=0.54 \
 //y=5.02 //x2=0.895 //y2=6.02
cc_90 ( N_VDD_c_65_p N_A_M3_noxref_g ) capacitor c=0.00697478f //x=1.47 \
 //y=7.4 //x2=1.335 //y2=6.02
cc_91 ( N_VDD_M3_noxref_d N_A_M3_noxref_g ) capacitor c=0.0528676f //x=1.41 \
 //y=5.02 //x2=1.335 //y2=6.02
cc_92 ( N_VDD_c_63_n N_A_c_233_n ) capacitor c=0.0099588f //x=2.22 //y=7.4 \
 //x2=1.26 //y2=4.79
cc_93 ( N_VDD_c_62_n N_A_c_234_n ) capacitor c=0.011132f //x=0.74 //y=7.4 \
 //x2=0.97 //y2=4.79
cc_94 ( N_VDD_M2_noxref_s N_A_c_234_n ) capacitor c=0.00665831f //x=0.54 \
 //y=5.02 //x2=0.97 //y2=4.79
cc_95 ( N_VDD_c_61_n Y ) capacitor c=0.0232778f //x=4.07 //y=7.4 //x2=3.7 \
 //y2=2.22
cc_96 ( N_VDD_c_63_n Y ) capacitor c=4.80934e-19 //x=2.22 //y=7.4 //x2=3.7 \
 //y2=2.22
cc_97 ( N_VDD_c_73_p N_Y_c_269_n ) capacitor c=8.92854e-19 //x=3.69 //y=7.4 \
 //x2=3.615 //y2=4.58
cc_98 ( N_VDD_M5_noxref_d N_Y_c_269_n ) capacitor c=0.00644908f //x=3.63 \
 //y=5.02 //x2=3.615 //y2=4.58
cc_99 ( N_VDD_c_63_n N_Y_c_271_n ) capacitor c=0.017572f //x=2.22 //y=7.4 \
 //x2=3.42 //y2=4.58
cc_100 ( N_VDD_c_81_p N_Y_M4_noxref_d ) capacitor c=0.00722811f //x=4.07 \
 //y=7.4 //x2=3.19 //y2=5.02
cc_101 ( N_VDD_c_73_p N_Y_M4_noxref_d ) capacitor c=0.0139004f //x=3.69 \
 //y=7.4 //x2=3.19 //y2=5.02
cc_102 ( N_VDD_c_61_n N_Y_M4_noxref_d ) capacitor c=0.0219131f //x=4.07 \
 //y=7.4 //x2=3.19 //y2=5.02
cc_103 ( N_VDD_M4_noxref_s N_Y_M4_noxref_d ) capacitor c=0.0843065f //x=2.76 \
 //y=5.02 //x2=3.19 //y2=5.02
cc_104 ( N_VDD_M5_noxref_d N_Y_M4_noxref_d ) capacitor c=0.0832641f //x=3.63 \
 //y=5.02 //x2=3.19 //y2=5.02
cc_105 ( N_noxref_3_c_112_n N_A_c_210_n ) capacitor c=0.00730959f //x=1.595 \
 //y=2.59 //x2=0.74 //y2=2.085
cc_106 ( N_noxref_3_c_144_n N_A_c_210_n ) capacitor c=0.0250789f //x=1.2 \
 //y=4.58 //x2=0.74 //y2=2.085
cc_107 ( N_noxref_3_c_117_n N_A_c_210_n ) capacitor c=0.0712221f //x=1.48 \
 //y=2.59 //x2=0.74 //y2=2.085
cc_108 ( N_noxref_3_c_120_n N_A_c_210_n ) capacitor c=0.00109894f //x=2.96 \
 //y=2.085 //x2=0.74 //y2=2.085
cc_109 ( N_noxref_3_M0_noxref_d N_A_c_210_n ) capacitor c=0.0175773f //x=0.925 \
 //y=0.91 //x2=0.74 //y2=2.085
cc_110 ( N_noxref_3_M2_noxref_d N_A_M2_noxref_g ) capacitor c=0.0219309f \
 //x=0.97 //y=5.02 //x2=0.895 //y2=6.02
cc_111 ( N_noxref_3_M2_noxref_d N_A_M3_noxref_g ) capacitor c=0.021902f \
 //x=0.97 //y=5.02 //x2=1.335 //y2=6.02
cc_112 ( N_noxref_3_M0_noxref_d N_A_c_215_n ) capacitor c=0.00218556f \
 //x=0.925 //y=0.91 //x2=0.85 //y2=0.91
cc_113 ( N_noxref_3_M0_noxref_d N_A_c_244_n ) capacitor c=0.00347355f \
 //x=0.925 //y=0.91 //x2=0.85 //y2=1.255
cc_114 ( N_noxref_3_M0_noxref_d N_A_c_245_n ) capacitor c=0.00742431f \
 //x=0.925 //y=0.91 //x2=0.85 //y2=1.565
cc_115 ( N_noxref_3_M0_noxref_d N_A_c_217_n ) capacitor c=0.00957707f \
 //x=0.925 //y=0.91 //x2=0.85 //y2=1.92
cc_116 ( N_noxref_3_c_142_n N_A_c_233_n ) capacitor c=0.0107726f //x=1.395 \
 //y=4.58 //x2=1.26 //y2=4.79
cc_117 ( N_noxref_3_M2_noxref_d N_A_c_233_n ) capacitor c=0.0148755f //x=0.97 \
 //y=5.02 //x2=1.26 //y2=4.79
cc_118 ( N_noxref_3_c_144_n N_A_c_234_n ) capacitor c=0.00962086f //x=1.2 \
 //y=4.58 //x2=0.97 //y2=4.79
cc_119 ( N_noxref_3_M2_noxref_d N_A_c_234_n ) capacitor c=0.00307344f //x=0.97 \
 //y=5.02 //x2=0.97 //y2=4.79
cc_120 ( N_noxref_3_M0_noxref_d N_A_c_218_n ) capacitor c=0.00220879f \
 //x=0.925 //y=0.91 //x2=1.225 //y2=0.755
cc_121 ( N_noxref_3_c_114_n N_A_c_252_n ) capacitor c=0.0023507f //x=1.395 \
 //y=2.08 //x2=1.225 //y2=1.41
cc_122 ( N_noxref_3_M0_noxref_d N_A_c_252_n ) capacitor c=0.0138447f //x=0.925 \
 //y=0.91 //x2=1.225 //y2=1.41
cc_123 ( N_noxref_3_M0_noxref_d N_A_c_219_n ) capacitor c=0.00218624f \
 //x=0.925 //y=0.91 //x2=1.38 //y2=0.91
cc_124 ( N_noxref_3_M0_noxref_d N_A_c_221_n ) capacitor c=0.00601286f \
 //x=0.925 //y=0.91 //x2=1.38 //y2=1.255
cc_125 ( N_noxref_3_c_184_p N_A_c_222_n ) capacitor c=0.0167852f //x=1.195 \
 //y=2.08 //x2=0.74 //y2=2.085
cc_126 ( N_noxref_3_c_117_n N_A_c_222_n ) capacitor c=8.49451e-19 //x=1.48 \
 //y=2.59 //x2=0.74 //y2=2.085
cc_127 ( N_noxref_3_c_108_n Y ) capacitor c=0.00730959f //x=2.845 //y=2.59 \
 //x2=3.7 //y2=2.22
cc_128 ( N_noxref_3_c_117_n Y ) capacitor c=0.00108914f //x=1.48 //y=2.59 \
 //x2=3.7 //y2=2.22
cc_129 ( N_noxref_3_c_120_n Y ) capacitor c=0.0712221f //x=2.96 //y=2.085 \
 //x2=3.7 //y2=2.22
cc_130 ( N_noxref_3_c_132_n Y ) capacitor c=8.49451e-19 //x=2.96 //y=2.085 \
 //x2=3.7 //y2=2.22
cc_131 ( N_noxref_3_c_190_p N_Y_c_259_n ) capacitor c=0.0023507f //x=3.445 \
 //y=1.41 //x2=3.615 //y2=2.08
cc_132 ( N_noxref_3_c_132_n N_Y_c_282_n ) capacitor c=0.0167852f //x=2.96 \
 //y=2.085 //x2=3.415 //y2=2.08
cc_133 ( N_noxref_3_c_155_n N_Y_c_269_n ) capacitor c=0.0107726f //x=3.48 \
 //y=4.79 //x2=3.615 //y2=4.58
cc_134 ( N_noxref_3_c_120_n N_Y_c_271_n ) capacitor c=0.0253118f //x=2.96 \
 //y=2.085 //x2=3.42 //y2=4.58
cc_135 ( N_noxref_3_c_156_n N_Y_c_271_n ) capacitor c=0.00962086f //x=3.19 \
 //y=4.79 //x2=3.42 //y2=4.58
cc_136 ( N_noxref_3_c_120_n N_Y_M1_noxref_d ) capacitor c=0.0177062f //x=2.96 \
 //y=2.085 //x2=3.145 //y2=0.91
cc_137 ( N_noxref_3_c_125_n N_Y_M1_noxref_d ) capacitor c=0.00218556f //x=3.07 \
 //y=0.91 //x2=3.145 //y2=0.91
cc_138 ( N_noxref_3_c_197_p N_Y_M1_noxref_d ) capacitor c=0.00347355f //x=3.07 \
 //y=1.255 //x2=3.145 //y2=0.91
cc_139 ( N_noxref_3_c_198_p N_Y_M1_noxref_d ) capacitor c=0.00742431f //x=3.07 \
 //y=1.565 //x2=3.145 //y2=0.91
cc_140 ( N_noxref_3_c_127_n N_Y_M1_noxref_d ) capacitor c=0.00957707f //x=3.07 \
 //y=1.92 //x2=3.145 //y2=0.91
cc_141 ( N_noxref_3_c_128_n N_Y_M1_noxref_d ) capacitor c=0.00220879f \
 //x=3.445 //y=0.755 //x2=3.145 //y2=0.91
cc_142 ( N_noxref_3_c_190_p N_Y_M1_noxref_d ) capacitor c=0.0138447f //x=3.445 \
 //y=1.41 //x2=3.145 //y2=0.91
cc_143 ( N_noxref_3_c_129_n N_Y_M1_noxref_d ) capacitor c=0.00218624f //x=3.6 \
 //y=0.91 //x2=3.145 //y2=0.91
cc_144 ( N_noxref_3_c_131_n N_Y_M1_noxref_d ) capacitor c=0.00601286f //x=3.6 \
 //y=1.255 //x2=3.145 //y2=0.91
cc_145 ( N_noxref_3_M0_noxref_d N_Y_M1_noxref_d ) capacitor c=2.55525e-19 \
 //x=0.925 //y=0.91 //x2=3.145 //y2=0.91
cc_146 ( N_noxref_3_M4_noxref_g N_Y_M4_noxref_d ) capacitor c=0.0219309f \
 //x=3.115 //y=6.02 //x2=3.19 //y2=5.02
cc_147 ( N_noxref_3_M5_noxref_g N_Y_M4_noxref_d ) capacitor c=0.021902f \
 //x=3.555 //y=6.02 //x2=3.19 //y2=5.02
cc_148 ( N_noxref_3_c_155_n N_Y_M4_noxref_d ) capacitor c=0.0148755f //x=3.48 \
 //y=4.79 //x2=3.19 //y2=5.02
cc_149 ( N_noxref_3_c_156_n N_Y_M4_noxref_d ) capacitor c=0.00307344f //x=3.19 \
 //y=4.79 //x2=3.19 //y2=5.02
cc_150 ( N_noxref_3_M2_noxref_d N_Y_M4_noxref_d ) capacitor c=7.38512e-19 \
 //x=0.97 //y=5.02 //x2=3.19 //y2=5.02
