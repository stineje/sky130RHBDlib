* SPICE3 file created from TMRDFFSNRNQNX1.ext - technology: sky130A

.subckt TMRDFFSNRNQNX1 Q D CLK SN RN VDD GND
X0 VDD RN a_277_1004 VDD pshort w=2 l=0.15 M=2
X1 GND a_7973_1004 a_8749_75 GND nshort w=3 l=0.15
X2 a_6371_943 a_6049_1004 VDD VDD pshort w=2 l=0.15 M=2
X3 VDD a_7973_1004 a_7333_943 VDD pshort w=2 l=0.15 M=2
X4 VDD a_9897_1004 a_10219_943 VDD pshort w=2 l=0.15 M=2
X5 a_17533_1005 a_4125_1004 VDD VDD pshort w=2 l=0.15 M=2
X6 a_12143_943 CLK VDD VDD pshort w=2 l=0.15 M=2
X7 GND D a_91_75 GND nshort w=3 l=0.15
X8 a_15991_943 a_15669_1004 VDD VDD pshort w=2 l=0.15 M=2
X9 a_599_943 a_1561_943 VDD VDD pshort w=2 l=0.15 M=2
X10 VDD RN a_1561_943 VDD pshort w=2 l=0.15 M=2
X11 a_11916_182 RN a_11635_75 GND nshort w=3 l=0.15
X12 a_9897_1004 a_6371_943 VDD VDD pshort w=2 l=0.15 M=2
X13 a_4125_1004 a_599_943 VDD VDD pshort w=2 l=0.15 M=2
X14 a_9992_182 RN a_9711_75 GND nshort w=3 l=0.15
X15 VDD SN a_2201_1004 VDD pshort w=2 l=0.15 M=2
X16 a_4125_1004 a_4447_943 VDD VDD pshort w=2 l=0.15 M=2
X17 GND a_4125_1004 a_17428_73 GND nshort w=3 l=0.15
X18 VDD a_6371_943 a_6049_1004 VDD pshort w=2 l=0.15 M=2
X19 a_18197_1005 a_4125_1004 a_17533_1005 VDD pshort w=2 l=0.15 M=2
X20 a_1561_943 CLK VDD VDD pshort w=2 l=0.15 M=2
X21 GND a_11821_1004 a_13559_75 GND nshort w=3 l=0.15
X22 GND a_12143_943 a_15483_75 GND nshort w=3 l=0.15
X23 VDD a_599_943 a_277_1004 VDD pshort w=2 l=0.15 M=2
X24 a_13745_1004 SN VDD VDD pshort w=2 l=0.15 M=2
X25 a_17533_1005 a_9897_1004 VDD VDD pshort w=2 l=0.15 M=2
X26 a_12143_943 a_11821_1004 VDD VDD pshort w=2 l=0.15 M=2
X27 a_14802_182 CLK a_14521_75 GND nshort w=3 l=0.15
X28 VDD a_13745_1004 a_13105_943 VDD pshort w=2 l=0.15 M=2
X29 Q a_15669_1004 a_18094_73 GND nshort w=3 l=0.15
X30 a_10954_182 SN a_10673_75 GND nshort w=3 l=0.15
X31 a_15991_943 SN VDD VDD pshort w=2 l=0.15 M=2
X32 a_16726_182 SN a_16445_75 GND nshort w=3 l=0.15
X33 a_12878_182 CLK a_12597_75 GND nshort w=3 l=0.15
X34 a_15669_1004 a_12143_943 VDD VDD pshort w=2 l=0.15 M=2
X35 VDD a_1561_943 a_2201_1004 VDD pshort w=2 l=0.15 M=2
X36 a_4125_1004 RN VDD VDD pshort w=2 l=0.15 M=2
X37 VDD RN a_6049_1004 VDD pshort w=2 l=0.15 M=2
X38 a_7973_1004 a_7333_943 VDD VDD pshort w=2 l=0.15 M=2
X39 a_9897_1004 a_10219_943 VDD VDD pshort w=2 l=0.15 M=2
X40 GND a_15669_1004 a_16445_75 GND nshort w=3 l=0.15
X41 VDD a_13105_943 a_15991_943 VDD pshort w=2 l=0.15 M=2
X42 a_1561_943 a_2201_1004 VDD VDD pshort w=2 l=0.15 M=2
X43 a_2201_1004 a_1561_943 a_2296_182 GND nshort w=3 l=0.15
X44 a_372_182 RN a_91_75 GND nshort w=3 l=0.15
X45 a_18197_1005 a_15669_1004 a_17533_1005 VDD pshort w=2 l=0.15 M=2
X46 VDD a_4125_1004 a_4447_943 VDD pshort w=2 l=0.15 M=2
X47 a_6371_943 CLK VDD VDD pshort w=2 l=0.15 M=2
X48 a_4125_1004 a_4447_943 a_4220_182 GND nshort w=3 l=0.15
X49 VDD CLK a_7333_943 VDD pshort w=2 l=0.15 M=2
X50 a_6049_1004 D VDD VDD pshort w=2 l=0.15 M=2
X51 Q a_9897_1004 a_18197_1005 VDD pshort w=2 l=0.15 M=2
X52 a_13840_182 SN a_13559_75 GND nshort w=3 l=0.15
X53 a_277_1004 D VDD VDD pshort w=2 l=0.15 M=2
X54 a_15764_182 RN a_15483_75 GND nshort w=3 l=0.15
X55 VDD CLK a_13105_943 VDD pshort w=2 l=0.15 M=2
X56 a_10219_943 a_7333_943 VDD VDD pshort w=2 l=0.15 M=2
X57 VDD a_11821_1004 a_13745_1004 VDD pshort w=2 l=0.15 M=2
X58 VDD a_13105_943 a_12143_943 VDD pshort w=2 l=0.15 M=2
X59 a_15669_1004 RN VDD VDD pshort w=2 l=0.15 M=2
X60 VDD a_277_1004 a_599_943 VDD pshort w=2 l=0.15 M=2
X61 a_9897_1004 RN VDD VDD pshort w=2 l=0.15 M=2
X62 VDD RN a_11821_1004 VDD pshort w=2 l=0.15 M=2
X63 GND a_277_1004 a_2015_75 GND nshort w=3 l=0.15
X64 a_599_943 a_1561_943 a_1334_182 GND nshort w=3 l=0.15
X65 a_6371_943 a_7333_943 a_7106_182 GND nshort w=3 l=0.15
X66 a_13745_1004 a_13105_943 VDD VDD pshort w=2 l=0.15 M=2
X67 VDD SN a_4447_943 VDD pshort w=2 l=0.15 M=2
X68 a_1561_943 RN a_3258_182 GND nshort w=3 l=0.15
X69 a_18197_1005 a_15669_1004 Q VDD pshort w=2 l=0.15 M=2
X70 VDD a_15991_943 a_15669_1004 VDD pshort w=2 l=0.15 M=2
X71 a_6371_943 a_7333_943 VDD VDD pshort w=2 l=0.15 M=2
X72 VDD RN a_7333_943 VDD pshort w=2 l=0.15 M=2
X73 a_4447_943 a_1561_943 a_5182_182 GND nshort w=3 l=0.15
X74 VDD SN a_7973_1004 VDD pshort w=2 l=0.15 M=2
X75 a_11821_1004 a_12143_943 a_11916_182 GND nshort w=3 l=0.15
X76 Q a_9897_1004 a_17428_73 GND nshort w=3 l=0.15
X77 a_6049_1004 a_6371_943 a_6144_182 GND nshort w=3 l=0.15
X78 VDD CLK a_599_943 VDD pshort w=2 l=0.15 M=2
X79 a_9897_1004 a_10219_943 a_9992_182 GND nshort w=3 l=0.15
X80 VDD a_12143_943 a_11821_1004 VDD pshort w=2 l=0.15 M=2
X81 a_7973_1004 a_7333_943 a_8068_182 GND nshort w=3 l=0.15
X82 GND a_2201_1004 a_2977_75 GND nshort w=3 l=0.15
X83 VDD a_1561_943 a_4447_943 VDD pshort w=2 l=0.15 M=2
X84 GND a_277_1004 a_1053_75 GND nshort w=3 l=0.15
X85 VDD a_6049_1004 a_7973_1004 VDD pshort w=2 l=0.15 M=2
X86 VDD RN a_13105_943 VDD pshort w=2 l=0.15 M=2
X87 a_4220_182 RN a_3939_75 GND nshort w=3 l=0.15
X88 a_11821_1004 D VDD VDD pshort w=2 l=0.15 M=2
X89 a_10219_943 a_7333_943 a_10954_182 GND nshort w=3 l=0.15
X90 a_2296_182 SN a_2015_75 GND nshort w=3 l=0.15
X91 a_12143_943 a_13105_943 a_12878_182 GND nshort w=3 l=0.15
X92 a_13105_943 RN a_14802_182 GND nshort w=3 l=0.15
X93 GND a_599_943 a_3939_75 GND nshort w=3 l=0.15
X94 a_2201_1004 a_277_1004 VDD VDD pshort w=2 l=0.15 M=2
X95 a_7333_943 RN a_9030_182 GND nshort w=3 l=0.15
X96 a_5182_182 SN a_4901_75 GND nshort w=3 l=0.15
X97 a_15669_1004 a_15991_943 a_15764_182 GND nshort w=3 l=0.15
X98 a_7106_182 CLK a_6825_75 GND nshort w=3 l=0.15
X99 a_1334_182 CLK a_1053_75 GND nshort w=3 l=0.15
X100 a_3258_182 CLK a_2977_75 GND nshort w=3 l=0.15
X101 a_13745_1004 a_13105_943 a_13840_182 GND nshort w=3 l=0.15
X102 GND a_6049_1004 a_6825_75 GND nshort w=3 l=0.15
X103 VDD SN a_10219_943 VDD pshort w=2 l=0.15 M=2
X104 GND a_4125_1004 a_4901_75 GND nshort w=3 l=0.15
X105 GND a_15669_1004 a_18760_73 GND nshort w=3 l=0.15
X106 GND a_4125_1004 a_18094_73 GND nshort w=3 l=0.15
X107 a_6144_182 RN a_5863_75 GND nshort w=3 l=0.15
X108 GND D a_11635_75 GND nshort w=3 l=0.15
X109 a_15991_943 a_13105_943 a_16726_182 GND nshort w=3 l=0.15
X110 a_8068_182 SN a_7787_75 GND nshort w=3 l=0.15
X111 GND a_6049_1004 a_7787_75 GND nshort w=3 l=0.15
X112 GND a_6371_943 a_9711_75 GND nshort w=3 l=0.15
X113 Q a_9897_1004 a_18760_73 GND nshort w=3 l=0.15
X114 GND D a_5863_75 GND nshort w=3 l=0.15
X115 a_277_1004 a_599_943 a_372_182 GND nshort w=3 l=0.15
X116 a_9030_182 CLK a_8749_75 GND nshort w=3 l=0.15
X117 GND a_11821_1004 a_12597_75 GND nshort w=3 l=0.15
X118 GND a_13745_1004 a_14521_75 GND nshort w=3 l=0.15
X119 GND a_9897_1004 a_10673_75 GND nshort w=3 l=0.15
C0 a_15669_1004 VDD 2.64fF
C1 a_599_943 VDD 2.45fF
C2 D a_1561_943 4.46fF
C3 VDD a_4447_943 2.06fF
C4 a_12143_943 a_9897_1004 2.03fF
C5 RN SN 5.64fF
C6 VDD a_4125_1004 6.68fF
C7 a_7333_943 D 4.46fF
C8 RN a_4125_1004 2.01fF
C9 a_6371_943 VDD 2.46fF
C10 CLK D 11.68fF
C11 a_15991_943 VDD 2.06fF
C12 VDD a_11821_1004 2.38fF
C13 a_10219_943 VDD 2.05fF
C14 a_13745_1004 VDD 2.07fF
C15 VDD a_13105_943 2.67fF
C16 a_12143_943 SN 3.98fF
C17 a_9897_1004 CLK 3.04fF
C18 SN D 2.38fF
C19 a_599_943 a_1561_943 3.19fF
C20 D a_4125_1004 3.05fF
C21 RN VDD 2.54fF
C22 a_9897_1004 SN 2.92fF
C23 a_6049_1004 VDD 2.38fF
C24 a_9897_1004 a_4125_1004 5.26fF
C25 SN CLK 2.43fF
C26 a_12143_943 a_13105_943 3.19fF
C27 CLK a_4125_1004 11.67fF
C28 a_7333_943 a_6371_943 3.19fF
C29 a_12143_943 VDD 2.46fF
C30 SN a_599_943 2.03fF
C31 D VDD 3.62fF
C32 a_9897_1004 a_13105_943 4.45fF
C33 VDD a_1561_943 2.66fF
C34 SN a_4125_1004 2.63fF
C35 RN D 2.04fF
C36 a_7333_943 VDD 2.66fF
C37 a_9897_1004 VDD 4.10fF
C38 a_6371_943 SN 3.98fF
C39 VDD a_277_1004 2.25fF
C40 CLK VDD 5.05fF
C41 VDD a_7973_1004 2.07fF
C42 VDD a_2201_1004 2.07fF
C43 RN CLK 2.23fF
C44 SN GND 4.14fF
C45 RN GND 5.22fF
C46 VDD GND 45.75fF
.ends
