// File: dffsnx1_pcell.spi.pex
// Created: Tue Oct 15 15:56:17 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_DFFSNX1_PCELL\%noxref_1 ( 41 45 48 53 61 67 77 83 93 99 105 113 121 \
 136 140 143 146 149 151 153 154 155 156 157 158 )
c285 ( 158 0 ) capacitor c=0.0226075f //x=20.495 //y=0.875
c286 ( 157 0 ) capacitor c=0.0207407f //x=17.27 //y=0.865
c287 ( 156 0 ) capacitor c=0.0207407f //x=13.94 //y=0.865
c288 ( 155 0 ) capacitor c=0.0226205f //x=9.025 //y=0.875
c289 ( 154 0 ) capacitor c=0.0226323f //x=4.215 //y=0.875
c290 ( 153 0 ) capacitor c=0.0208404f //x=0.99 //y=0.865
c291 ( 152 0 ) capacitor c=0.00440144f //x=20.685 //y=0
c292 ( 151 0 ) capacitor c=0.105142f //x=19.61 //y=0
c293 ( 150 0 ) capacitor c=0.00440095f //x=17.46 //y=0
c294 ( 149 0 ) capacitor c=0.106174f //x=16.28 //y=0
c295 ( 148 0 ) capacitor c=0.00440095f //x=14.06 //y=0
c296 ( 146 0 ) capacitor c=0.108248f //x=12.95 //y=0
c297 ( 145 0 ) capacitor c=0.00440144f //x=9.25 //y=0
c298 ( 143 0 ) capacitor c=0.108235f //x=8.14 //y=0
c299 ( 142 0 ) capacitor c=0.00440144f //x=4.44 //y=0
c300 ( 140 0 ) capacitor c=0.105313f //x=3.33 //y=0
c301 ( 139 0 ) capacitor c=0.00440095f //x=1.18 //y=0
c302 ( 136 0 ) capacitor c=0.322261f //x=23.68 //y=0
c303 ( 121 0 ) capacitor c=0.0339325f //x=20.6 //y=0
c304 ( 113 0 ) capacitor c=0.0718026f //x=19.44 //y=0
c305 ( 105 0 ) capacitor c=0.0388888f //x=17.375 //y=0
c306 ( 99 0 ) capacitor c=0.0718026f //x=16.11 //y=0
c307 ( 93 0 ) capacitor c=0.0388888f //x=14.045 //y=0
c308 ( 83 0 ) capacitor c=0.133402f //x=12.78 //y=0
c309 ( 77 0 ) capacitor c=0.0339482f //x=9.13 //y=0
c310 ( 67 0 ) capacitor c=0.133515f //x=7.97 //y=0
c311 ( 61 0 ) capacitor c=0.0339482f //x=4.32 //y=0
c312 ( 53 0 ) capacitor c=0.0720582f //x=3.16 //y=0
c313 ( 48 0 ) capacitor c=0.179262f //x=0.74 //y=0
c314 ( 45 0 ) capacitor c=0.0426751f //x=1.095 //y=0
c315 ( 41 0 ) capacitor c=0.776195f //x=23.68 //y=0
r316 (  134 136 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=22.57 //y=0 //x2=23.68 //y2=0
r317 (  132 134 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.46 //y=0 //x2=22.57 //y2=0
r318 (  130 152 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.77 //y=0 //x2=20.685 //y2=0
r319 (  130 132 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=20.77 //y=0 //x2=21.46 //y2=0
r320 (  125 152 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.685 //y=0.17 //x2=20.685 //y2=0
r321 (  125 158 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=20.685 //y=0.17 //x2=20.685 //y2=0.965
r322 (  122 151 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.78 //y=0 //x2=19.61 //y2=0
r323 (  122 124 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.78 //y=0 //x2=20.35 //y2=0
r324 (  121 152 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.6 //y=0 //x2=20.685 //y2=0
r325 (  121 124 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=20.6 //y=0 //x2=20.35 //y2=0
r326 (  116 118 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.76 //y=0 //x2=18.87 //y2=0
r327 (  114 150 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.545 //y=0 //x2=17.46 //y2=0
r328 (  114 116 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=17.545 //y=0 //x2=17.76 //y2=0
r329 (  113 151 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.44 //y=0 //x2=19.61 //y2=0
r330 (  113 118 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.44 //y=0 //x2=18.87 //y2=0
r331 (  109 150 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.46 //y=0.17 //x2=17.46 //y2=0
r332 (  109 157 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=17.46 //y=0.17 //x2=17.46 //y2=0.955
r333 (  106 149 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.45 //y=0 //x2=16.28 //y2=0
r334 (  106 108 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=16.45 //y=0 //x2=16.65 //y2=0
r335 (  105 150 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.375 //y=0 //x2=17.46 //y2=0
r336 (  105 108 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=17.375 //y=0 //x2=16.65 //y2=0
r337 (  100 148 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.215 //y=0 //x2=14.13 //y2=0
r338 (  100 102 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=14.215 //y=0 //x2=15.17 //y2=0
r339 (  99 149 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.11 //y=0 //x2=16.28 //y2=0
r340 (  99 102 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=16.11 //y=0 //x2=15.17 //y2=0
r341 (  95 148 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.13 //y=0.17 //x2=14.13 //y2=0
r342 (  95 156 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=14.13 //y=0.17 //x2=14.13 //y2=0.955
r343 (  94 146 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=0 //x2=12.95 //y2=0
r344 (  93 148 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.045 //y=0 //x2=14.13 //y2=0
r345 (  93 94 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=14.045 //y=0 //x2=13.12 //y2=0
r346 (  88 90 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r347 (  86 88 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=10.36 //y=0 //x2=11.47 //y2=0
r348 (  84 145 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.3 //y=0 //x2=9.215 //y2=0
r349 (  84 86 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=9.3 //y=0 //x2=10.36 //y2=0
r350 (  83 146 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.95 //y2=0
r351 (  83 90 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.58 //y2=0
r352 (  79 145 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.215 //y=0.17 //x2=9.215 //y2=0
r353 (  79 155 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=9.215 //y=0.17 //x2=9.215 //y2=0.965
r354 (  78 143 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=0 //x2=8.14 //y2=0
r355 (  77 145 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.13 //y=0 //x2=9.215 //y2=0
r356 (  77 78 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=9.13 //y=0 //x2=8.31 //y2=0
r357 (  72 74 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r358 (  70 72 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=5.55 //y=0 //x2=6.66 //y2=0
r359 (  68 142 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.49 //y=0 //x2=4.405 //y2=0
r360 (  68 70 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=4.49 //y=0 //x2=5.55 //y2=0
r361 (  67 143 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=8.14 //y2=0
r362 (  67 74 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=7.77 //y2=0
r363 (  63 142 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.405 //y=0.17 //x2=4.405 //y2=0
r364 (  63 154 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=4.405 //y=0.17 //x2=4.405 //y2=0.965
r365 (  62 140 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=0 //x2=3.33 //y2=0
r366 (  61 142 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.32 //y=0 //x2=4.405 //y2=0
r367 (  61 62 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=4.32 //y=0 //x2=3.5 //y2=0
r368 (  56 58 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r369 (  54 139 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.18 //y2=0
r370 (  54 56 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.85 //y2=0
r371 (  53 140 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=3.33 //y2=0
r372 (  53 58 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r373 (  49 139 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r374 (  49 153 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.955
r375 (  45 139 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=1.18 //y2=0
r376 (  45 48 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=0.74 //y2=0
r377 (  41 136 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=0 //x2=23.68 //y2=0
r378 (  39 134 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=0 //x2=22.57 //y2=0
r379 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=0 //x2=23.68 //y2=0
r380 (  37 132 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.46 //y=0 //x2=21.46 //y2=0
r381 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.46 //y=0 //x2=22.57 //y2=0
r382 (  35 124 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=0 //x2=20.35 //y2=0
r383 (  35 37 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=0 //x2=21.46 //y2=0
r384 (  33 118 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=0 //x2=18.87 //y2=0
r385 (  33 35 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=0 //x2=20.35 //y2=0
r386 (  31 116 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=0 //x2=17.76 //y2=0
r387 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=0 //x2=18.87 //y2=0
r388 (  29 108 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=0 //x2=16.65 //y2=0
r389 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=0 //x2=17.76 //y2=0
r390 (  27 102 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r391 (  27 29 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.65 //y2=0
r392 (  25 148 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=0 //x2=14.06 //y2=0
r393 (  25 27 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=0 //x2=15.17 //y2=0
r394 (  23 90 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r395 (  23 25 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=0 //x2=14.06 //y2=0
r396 (  21 88 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r397 (  21 23 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=0 //x2=12.58 //y2=0
r398 (  19 86 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r399 (  19 21 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r400 (  17 145 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=0 //x2=9.25 //y2=0
r401 (  17 19 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=0 //x2=10.36 //y2=0
r402 (  15 74 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r403 (  15 17 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=9.25 //y2=0
r404 (  13 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r405 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r406 (  11 70 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r407 (  11 13 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r408 (  9 142 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r409 (  9 11 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.55 //y2=0
r410 (  7 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r411 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r412 (  5 56 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r413 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r414 (  2 48 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r415 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_DFFSNX1_PCELL\%noxref_1

subckt PM_DFFSNX1_PCELL\%noxref_2 ( 41 53 61 71 77 85 93 103 113 119 127 135 \
 145 155 161 169 179 189 193 203 213 235 245 253 266 270 273 279 285 289 294 \
 299 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 \
 318 319 )
c303 ( 319 0 ) capacitor c=0.0455453f //x=23.195 //y=5.02
c304 ( 318 0 ) capacitor c=0.0243052f //x=22.315 //y=5.02
c305 ( 317 0 ) capacitor c=0.0243052f //x=21.435 //y=5.02
c306 ( 316 0 ) capacitor c=0.0532751f //x=20.565 //y=5.02
c307 ( 315 0 ) capacitor c=0.0382117f //x=18.685 //y=5.02
c308 ( 314 0 ) capacitor c=0.024147f //x=17.805 //y=5.02
c309 ( 313 0 ) capacitor c=0.0493657f //x=16.935 //y=5.02
c310 ( 312 0 ) capacitor c=0.0381505f //x=15.355 //y=5.02
c311 ( 311 0 ) capacitor c=0.0240074f //x=14.475 //y=5.02
c312 ( 310 0 ) capacitor c=0.049209f //x=13.605 //y=5.02
c313 ( 309 0 ) capacitor c=0.0452179f //x=11.725 //y=5.02
c314 ( 308 0 ) capacitor c=0.024152f //x=10.845 //y=5.02
c315 ( 307 0 ) capacitor c=0.024152f //x=9.965 //y=5.02
c316 ( 306 0 ) capacitor c=0.053132f //x=9.095 //y=5.02
c317 ( 305 0 ) capacitor c=0.0452179f //x=6.915 //y=5.02
c318 ( 304 0 ) capacitor c=0.024152f //x=6.035 //y=5.02
c319 ( 303 0 ) capacitor c=0.02424f //x=5.155 //y=5.02
c320 ( 302 0 ) capacitor c=0.0532367f //x=4.285 //y=5.02
c321 ( 301 0 ) capacitor c=0.0381505f //x=2.405 //y=5.02
c322 ( 300 0 ) capacitor c=0.024246f //x=1.525 //y=5.02
c323 ( 299 0 ) capacitor c=0.053196f //x=0.655 //y=5.02
c324 ( 298 0 ) capacitor c=0.00591168f //x=23.34 //y=7.4
c325 ( 297 0 ) capacitor c=0.00591168f //x=22.46 //y=7.4
c326 ( 296 0 ) capacitor c=0.00591168f //x=21.58 //y=7.4
c327 ( 295 0 ) capacitor c=0.00591168f //x=20.7 //y=7.4
c328 ( 294 0 ) capacitor c=0.139422f //x=19.61 //y=7.4
c329 ( 293 0 ) capacitor c=0.00591168f //x=18.87 //y=7.4
c330 ( 291 0 ) capacitor c=0.00591168f //x=17.95 //y=7.4
c331 ( 290 0 ) capacitor c=0.00591168f //x=17.07 //y=7.4
c332 ( 289 0 ) capacitor c=0.116163f //x=16.28 //y=7.4
c333 ( 288 0 ) capacitor c=0.00591168f //x=15.5 //y=7.4
c334 ( 287 0 ) capacitor c=0.00591168f //x=14.62 //y=7.4
c335 ( 286 0 ) capacitor c=0.00591168f //x=13.74 //y=7.4
c336 ( 285 0 ) capacitor c=0.13452f //x=12.95 //y=7.4
c337 ( 284 0 ) capacitor c=0.00591168f //x=11.87 //y=7.4
c338 ( 283 0 ) capacitor c=0.00591168f //x=10.99 //y=7.4
c339 ( 282 0 ) capacitor c=0.00591168f //x=10.11 //y=7.4
c340 ( 281 0 ) capacitor c=0.00591168f //x=9.25 //y=7.4
c341 ( 279 0 ) capacitor c=0.155082f //x=8.14 //y=7.4
c342 ( 278 0 ) capacitor c=0.00591168f //x=7.06 //y=7.4
c343 ( 277 0 ) capacitor c=0.00591168f //x=6.18 //y=7.4
c344 ( 276 0 ) capacitor c=0.00591168f //x=5.3 //y=7.4
c345 ( 275 0 ) capacitor c=0.00591168f //x=4.44 //y=7.4
c346 ( 273 0 ) capacitor c=0.137403f //x=3.33 //y=7.4
c347 ( 272 0 ) capacitor c=0.00591168f //x=2.55 //y=7.4
c348 ( 271 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c349 ( 270 0 ) capacitor c=0.248311f //x=0.74 //y=7.4
c350 ( 266 0 ) capacitor c=0.272255f //x=23.68 //y=7.4
c351 ( 253 0 ) capacitor c=0.028513f //x=23.255 //y=7.4
c352 ( 245 0 ) capacitor c=0.0287069f //x=22.375 //y=7.4
c353 ( 235 0 ) capacitor c=0.0292055f //x=21.495 //y=7.4
c354 ( 225 0 ) capacitor c=0.0452081f //x=20.615 //y=7.4
c355 ( 221 0 ) capacitor c=0.0275781f //x=19.44 //y=7.4
c356 ( 213 0 ) capacitor c=0.0285035f //x=18.745 //y=7.4
c357 ( 203 0 ) capacitor c=0.0291038f //x=17.865 //y=7.4
c358 ( 193 0 ) capacitor c=0.0240981f //x=16.985 //y=7.4
c359 ( 189 0 ) capacitor c=0.0236224f //x=16.11 //y=7.4
c360 ( 179 0 ) capacitor c=0.0288598f //x=15.415 //y=7.4
c361 ( 169 0 ) capacitor c=0.0288369f //x=14.535 //y=7.4
c362 ( 161 0 ) capacitor c=0.0240981f //x=13.655 //y=7.4
c363 ( 155 0 ) capacitor c=0.0394667f //x=12.78 //y=7.4
c364 ( 145 0 ) capacitor c=0.0288488f //x=11.785 //y=7.4
c365 ( 135 0 ) capacitor c=0.0287514f //x=10.905 //y=7.4
c366 ( 127 0 ) capacitor c=0.0284966f //x=10.025 //y=7.4
c367 ( 119 0 ) capacitor c=0.0383672f //x=9.145 //y=7.4
c368 ( 113 0 ) capacitor c=0.0394667f //x=7.97 //y=7.4
c369 ( 103 0 ) capacitor c=0.0288488f //x=6.975 //y=7.4
c370 ( 93 0 ) capacitor c=0.0287505f //x=6.095 //y=7.4
c371 ( 85 0 ) capacitor c=0.028511f //x=5.215 //y=7.4
c372 ( 77 0 ) capacitor c=0.0383672f //x=4.335 //y=7.4
c373 ( 71 0 ) capacitor c=0.0236224f //x=3.16 //y=7.4
c374 ( 61 0 ) capacitor c=0.0288637f //x=2.465 //y=7.4
c375 ( 53 0 ) capacitor c=0.0286367f //x=1.585 //y=7.4
c376 ( 41 0 ) capacitor c=0.8559f //x=23.68 //y=7.4
r377 (  264 298 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.425 //y=7.4 //x2=23.34 //y2=7.4
r378 (  264 266 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=23.425 //y=7.4 //x2=23.68 //y2=7.4
r379 (  257 298 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.34 //y=7.23 //x2=23.34 //y2=7.4
r380 (  257 319 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=23.34 //y=7.23 //x2=23.34 //y2=6.745
r381 (  254 297 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.545 //y=7.4 //x2=22.46 //y2=7.4
r382 (  254 256 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=22.545 //y=7.4 //x2=22.57 //y2=7.4
r383 (  253 298 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.255 //y=7.4 //x2=23.34 //y2=7.4
r384 (  253 256 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=23.255 //y=7.4 //x2=22.57 //y2=7.4
r385 (  247 297 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.46 //y=7.23 //x2=22.46 //y2=7.4
r386 (  247 318 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.46 //y=7.23 //x2=22.46 //y2=6.745
r387 (  246 296 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.665 //y=7.4 //x2=21.58 //y2=7.4
r388 (  245 297 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.375 //y=7.4 //x2=22.46 //y2=7.4
r389 (  245 246 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.375 //y=7.4 //x2=21.665 //y2=7.4
r390 (  239 296 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.58 //y=7.23 //x2=21.58 //y2=7.4
r391 (  239 317 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.58 //y=7.23 //x2=21.58 //y2=6.745
r392 (  236 295 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.785 //y=7.4 //x2=20.7 //y2=7.4
r393 (  236 238 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=20.785 //y=7.4 //x2=21.46 //y2=7.4
r394 (  235 296 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.495 //y=7.4 //x2=21.58 //y2=7.4
r395 (  235 238 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=21.495 //y=7.4 //x2=21.46 //y2=7.4
r396 (  229 295 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.7 //y=7.23 //x2=20.7 //y2=7.4
r397 (  229 316 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=20.7 //y=7.23 //x2=20.7 //y2=6.405
r398 (  226 294 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.78 //y=7.4 //x2=19.61 //y2=7.4
r399 (  226 228 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.78 //y=7.4 //x2=20.35 //y2=7.4
r400 (  225 295 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.615 //y=7.4 //x2=20.7 //y2=7.4
r401 (  225 228 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.615 //y=7.4 //x2=20.35 //y2=7.4
r402 (  222 293 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.915 //y=7.4 //x2=18.83 //y2=7.4
r403 (  221 294 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.44 //y=7.4 //x2=19.61 //y2=7.4
r404 (  221 222 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=19.44 //y=7.4 //x2=18.915 //y2=7.4
r405 (  215 293 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.83 //y=7.23 //x2=18.83 //y2=7.4
r406 (  215 315 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=18.83 //y=7.23 //x2=18.83 //y2=6.745
r407 (  214 291 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.035 //y=7.4 //x2=17.95 //y2=7.4
r408 (  213 293 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.745 //y=7.4 //x2=18.83 //y2=7.4
r409 (  213 214 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=18.745 //y=7.4 //x2=18.035 //y2=7.4
r410 (  207 291 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.95 //y=7.23 //x2=17.95 //y2=7.4
r411 (  207 314 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.95 //y=7.23 //x2=17.95 //y2=6.745
r412 (  204 290 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.155 //y=7.4 //x2=17.07 //y2=7.4
r413 (  204 206 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=17.155 //y=7.4 //x2=17.76 //y2=7.4
r414 (  203 291 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.865 //y=7.4 //x2=17.95 //y2=7.4
r415 (  203 206 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=17.865 //y=7.4 //x2=17.76 //y2=7.4
r416 (  197 290 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.07 //y=7.23 //x2=17.07 //y2=7.4
r417 (  197 313 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=17.07 //y=7.23 //x2=17.07 //y2=6.405
r418 (  194 289 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.45 //y=7.4 //x2=16.28 //y2=7.4
r419 (  194 196 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=16.45 //y=7.4 //x2=16.65 //y2=7.4
r420 (  193 290 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.985 //y=7.4 //x2=17.07 //y2=7.4
r421 (  193 196 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=16.985 //y=7.4 //x2=16.65 //y2=7.4
r422 (  190 288 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.585 //y=7.4 //x2=15.5 //y2=7.4
r423 (  189 289 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.11 //y=7.4 //x2=16.28 //y2=7.4
r424 (  189 190 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=16.11 //y=7.4 //x2=15.585 //y2=7.4
r425 (  183 288 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.5 //y=7.23 //x2=15.5 //y2=7.4
r426 (  183 312 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.5 //y=7.23 //x2=15.5 //y2=6.745
r427 (  180 287 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.705 //y=7.4 //x2=14.62 //y2=7.4
r428 (  180 182 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=14.705 //y=7.4 //x2=15.17 //y2=7.4
r429 (  179 288 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.415 //y=7.4 //x2=15.5 //y2=7.4
r430 (  179 182 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=15.415 //y=7.4 //x2=15.17 //y2=7.4
r431 (  173 287 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.62 //y=7.23 //x2=14.62 //y2=7.4
r432 (  173 311 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.62 //y=7.23 //x2=14.62 //y2=6.745
r433 (  170 286 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.825 //y=7.4 //x2=13.74 //y2=7.4
r434 (  170 172 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=13.825 //y=7.4 //x2=14.06 //y2=7.4
r435 (  169 287 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.535 //y=7.4 //x2=14.62 //y2=7.4
r436 (  169 172 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=14.535 //y=7.4 //x2=14.06 //y2=7.4
r437 (  163 286 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.74 //y=7.23 //x2=13.74 //y2=7.4
r438 (  163 310 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=13.74 //y=7.23 //x2=13.74 //y2=6.405
r439 (  162 285 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=7.4 //x2=12.95 //y2=7.4
r440 (  161 286 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.655 //y=7.4 //x2=13.74 //y2=7.4
r441 (  161 162 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=13.655 //y=7.4 //x2=13.12 //y2=7.4
r442 (  156 284 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.955 //y=7.4 //x2=11.87 //y2=7.4
r443 (  156 158 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=11.955 //y=7.4 //x2=12.58 //y2=7.4
r444 (  155 285 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.95 //y2=7.4
r445 (  155 158 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.58 //y2=7.4
r446 (  149 284 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.87 //y=7.23 //x2=11.87 //y2=7.4
r447 (  149 309 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.87 //y=7.23 //x2=11.87 //y2=6.745
r448 (  146 283 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.075 //y=7.4 //x2=10.99 //y2=7.4
r449 (  146 148 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=11.075 //y=7.4 //x2=11.47 //y2=7.4
r450 (  145 284 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.785 //y=7.4 //x2=11.87 //y2=7.4
r451 (  145 148 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=11.785 //y=7.4 //x2=11.47 //y2=7.4
r452 (  139 283 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.99 //y=7.23 //x2=10.99 //y2=7.4
r453 (  139 308 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.99 //y=7.23 //x2=10.99 //y2=6.745
r454 (  136 282 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.195 //y=7.4 //x2=10.11 //y2=7.4
r455 (  136 138 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=10.195 //y=7.4 //x2=10.36 //y2=7.4
r456 (  135 283 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.905 //y=7.4 //x2=10.99 //y2=7.4
r457 (  135 138 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=10.905 //y=7.4 //x2=10.36 //y2=7.4
r458 (  129 282 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.11 //y=7.23 //x2=10.11 //y2=7.4
r459 (  129 307 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.11 //y=7.23 //x2=10.11 //y2=6.745
r460 (  128 281 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.315 //y=7.4 //x2=9.23 //y2=7.4
r461 (  127 282 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.025 //y=7.4 //x2=10.11 //y2=7.4
r462 (  127 128 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.025 //y=7.4 //x2=9.315 //y2=7.4
r463 (  121 281 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.23 //y=7.23 //x2=9.23 //y2=7.4
r464 (  121 306 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=9.23 //y=7.23 //x2=9.23 //y2=6.405
r465 (  120 279 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=7.4 //x2=8.14 //y2=7.4
r466 (  119 281 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.145 //y=7.4 //x2=9.23 //y2=7.4
r467 (  119 120 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=9.145 //y=7.4 //x2=8.31 //y2=7.4
r468 (  114 278 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.145 //y=7.4 //x2=7.06 //y2=7.4
r469 (  114 116 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=7.145 //y=7.4 //x2=7.77 //y2=7.4
r470 (  113 279 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=8.14 //y2=7.4
r471 (  113 116 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=7.77 //y2=7.4
r472 (  107 278 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.06 //y=7.23 //x2=7.06 //y2=7.4
r473 (  107 305 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.06 //y=7.23 //x2=7.06 //y2=6.745
r474 (  104 277 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.265 //y=7.4 //x2=6.18 //y2=7.4
r475 (  104 106 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=6.265 //y=7.4 //x2=6.66 //y2=7.4
r476 (  103 278 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.975 //y=7.4 //x2=7.06 //y2=7.4
r477 (  103 106 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=6.975 //y=7.4 //x2=6.66 //y2=7.4
r478 (  97 277 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.18 //y=7.23 //x2=6.18 //y2=7.4
r479 (  97 304 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.18 //y=7.23 //x2=6.18 //y2=6.745
r480 (  94 276 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.385 //y=7.4 //x2=5.3 //y2=7.4
r481 (  94 96 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=5.385 //y=7.4 //x2=5.55 //y2=7.4
r482 (  93 277 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.095 //y=7.4 //x2=6.18 //y2=7.4
r483 (  93 96 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=6.095 //y=7.4 //x2=5.55 //y2=7.4
r484 (  87 276 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.3 //y=7.23 //x2=5.3 //y2=7.4
r485 (  87 303 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=5.3 //y=7.23 //x2=5.3 //y2=6.745
r486 (  86 275 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.505 //y=7.4 //x2=4.42 //y2=7.4
r487 (  85 276 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.215 //y=7.4 //x2=5.3 //y2=7.4
r488 (  85 86 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.215 //y=7.4 //x2=4.505 //y2=7.4
r489 (  79 275 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.42 //y=7.23 //x2=4.42 //y2=7.4
r490 (  79 302 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.42 //y=7.23 //x2=4.42 //y2=6.405
r491 (  78 273 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r492 (  77 275 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.335 //y=7.4 //x2=4.42 //y2=7.4
r493 (  77 78 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=4.335 //y=7.4 //x2=3.5 //y2=7.4
r494 (  72 272 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.55 //y2=7.4
r495 (  72 74 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.96 //y2=7.4
r496 (  71 273 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r497 (  71 74 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r498 (  65 272 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r499 (  65 301 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.745
r500 (  62 271 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r501 (  62 64 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r502 (  61 272 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r503 (  61 64 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r504 (  55 271 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r505 (  55 300 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.745
r506 (  54 270 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r507 (  53 271 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r508 (  53 54 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r509 (  47 270 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r510 (  47 299 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.405
r511 (  41 266 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=7.4 //x2=23.68 //y2=7.4
r512 (  39 256 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=7.4 //x2=22.57 //y2=7.4
r513 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=7.4 //x2=23.68 //y2=7.4
r514 (  37 238 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.46 //y=7.4 //x2=21.46 //y2=7.4
r515 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.46 //y=7.4 //x2=22.57 //y2=7.4
r516 (  35 228 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=7.4 //x2=20.35 //y2=7.4
r517 (  35 37 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=7.4 //x2=21.46 //y2=7.4
r518 (  33 293 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=7.4 //x2=18.87 //y2=7.4
r519 (  33 35 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=7.4 //x2=20.35 //y2=7.4
r520 (  31 206 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=7.4 //x2=17.76 //y2=7.4
r521 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=7.4 //x2=18.87 //y2=7.4
r522 (  29 196 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=7.4 //x2=16.65 //y2=7.4
r523 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=7.4 //x2=17.76 //y2=7.4
r524 (  27 182 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r525 (  27 29 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.65 //y2=7.4
r526 (  25 172 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=7.4 //x2=14.06 //y2=7.4
r527 (  25 27 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=7.4 //x2=15.17 //y2=7.4
r528 (  23 158 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r529 (  23 25 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.4 //x2=14.06 //y2=7.4
r530 (  21 148 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r531 (  21 23 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=7.4 //x2=12.58 //y2=7.4
r532 (  19 138 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r533 (  19 21 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r534 (  17 281 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=7.4 //x2=9.25 //y2=7.4
r535 (  17 19 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=7.4 //x2=10.36 //y2=7.4
r536 (  15 116 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r537 (  15 17 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=9.25 //y2=7.4
r538 (  13 106 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r539 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r540 (  11 96 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r541 (  11 13 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r542 (  9 275 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r543 (  9 11 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.55 //y2=7.4
r544 (  7 74 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r545 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r546 (  5 64 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r547 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r548 (  2 270 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r549 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_DFFSNX1_PCELL\%noxref_2

subckt PM_DFFSNX1_PCELL\%noxref_3 ( 1 2 3 4 17 18 29 31 32 36 38 46 53 54 55 \
 56 57 58 59 60 61 62 63 64 66 72 73 74 75 79 80 81 82 83 85 91 92 93 94 114 \
 116 117 )
c240 ( 117 0 ) capacitor c=0.0220291f //x=1.965 //y=5.02
c241 ( 116 0 ) capacitor c=0.0217503f //x=1.085 //y=5.02
c242 ( 114 0 ) capacitor c=0.0084702f //x=1.96 //y=0.905
c243 ( 94 0 ) capacitor c=0.0556143f //x=9.525 //y=4.79
c244 ( 93 0 ) capacitor c=0.0293157f //x=9.815 //y=4.79
c245 ( 92 0 ) capacitor c=0.0347816f //x=9.48 //y=1.22
c246 ( 91 0 ) capacitor c=0.0187487f //x=9.48 //y=0.875
c247 ( 85 0 ) capacitor c=0.0137055f //x=9.325 //y=1.375
c248 ( 83 0 ) capacitor c=0.0149861f //x=9.325 //y=0.72
c249 ( 82 0 ) capacitor c=0.0965257f //x=8.95 //y=1.915
c250 ( 81 0 ) capacitor c=0.0229444f //x=8.95 //y=1.53
c251 ( 80 0 ) capacitor c=0.0234352f //x=8.95 //y=1.22
c252 ( 79 0 ) capacitor c=0.0198724f //x=8.95 //y=0.875
c253 ( 75 0 ) capacitor c=0.055995f //x=4.715 //y=4.79
c254 ( 74 0 ) capacitor c=0.0298189f //x=5.005 //y=4.79
c255 ( 73 0 ) capacitor c=0.0347816f //x=4.67 //y=1.22
c256 ( 72 0 ) capacitor c=0.0187487f //x=4.67 //y=0.875
c257 ( 66 0 ) capacitor c=0.0137055f //x=4.515 //y=1.375
c258 ( 64 0 ) capacitor c=0.0149861f //x=4.515 //y=0.72
c259 ( 63 0 ) capacitor c=0.0965245f //x=4.14 //y=1.915
c260 ( 62 0 ) capacitor c=0.0229444f //x=4.14 //y=1.53
c261 ( 61 0 ) capacitor c=0.0234352f //x=4.14 //y=1.22
c262 ( 60 0 ) capacitor c=0.0198724f //x=4.14 //y=0.875
c263 ( 59 0 ) capacitor c=0.110114f //x=9.89 //y=6.02
c264 ( 58 0 ) capacitor c=0.158956f //x=9.45 //y=6.02
c265 ( 57 0 ) capacitor c=0.110114f //x=5.08 //y=6.02
c266 ( 56 0 ) capacitor c=0.158956f //x=4.64 //y=6.02
c267 ( 53 0 ) capacitor c=0.0023043f //x=2.11 //y=5.2
c268 ( 46 0 ) capacitor c=0.10363f //x=9.25 //y=2.08
c269 ( 38 0 ) capacitor c=0.108245f //x=4.44 //y=2.08
c270 ( 36 0 ) capacitor c=0.114138f //x=2.59 //y=2.59
c271 ( 32 0 ) capacitor c=0.00550359f //x=2.235 //y=1.655
c272 ( 31 0 ) capacitor c=0.0140493f //x=2.505 //y=1.655
c273 ( 29 0 ) capacitor c=0.0140934f //x=2.505 //y=5.2
c274 ( 18 0 ) capacitor c=0.00387264f //x=1.315 //y=5.2
c275 ( 17 0 ) capacitor c=0.019002f //x=2.025 //y=5.2
c276 ( 4 0 ) capacitor c=0.012652f //x=4.705 //y=2.59
c277 ( 3 0 ) capacitor c=0.143287f //x=9.135 //y=2.59
c278 ( 2 0 ) capacitor c=0.0148669f //x=2.705 //y=2.59
c279 ( 1 0 ) capacitor c=0.0543359f //x=4.295 //y=2.59
r280 (  93 95 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.815 //y=4.79 //x2=9.89 //y2=4.865
r281 (  93 94 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=9.815 //y=4.79 //x2=9.525 //y2=4.79
r282 (  92 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.48 //y=1.22 //x2=9.44 //y2=1.375
r283 (  91 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.48 //y=0.875 //x2=9.44 //y2=0.72
r284 (  91 92 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.48 //y=0.875 //x2=9.48 //y2=1.22
r285 (  88 94 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.45 //y=4.865 //x2=9.525 //y2=4.79
r286 (  88 111 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=9.45 //y=4.865 //x2=9.25 //y2=4.7
r287 (  86 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.105 //y=1.375 //x2=8.99 //y2=1.375
r288 (  85 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.325 //y=1.375 //x2=9.44 //y2=1.375
r289 (  84 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.105 //y=0.72 //x2=8.99 //y2=0.72
r290 (  83 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.325 //y=0.72 //x2=9.44 //y2=0.72
r291 (  83 84 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=9.325 //y=0.72 //x2=9.105 //y2=0.72
r292 (  82 109 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.915 //x2=9.25 //y2=2.08
r293 (  81 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.53 //x2=8.99 //y2=1.375
r294 (  81 82 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.53 //x2=8.95 //y2=1.915
r295 (  80 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.22 //x2=8.99 //y2=1.375
r296 (  79 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=0.875 //x2=8.99 //y2=0.72
r297 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.95 //y=0.875 //x2=8.95 //y2=1.22
r298 (  74 76 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.005 //y=4.79 //x2=5.08 //y2=4.865
r299 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=5.005 //y=4.79 //x2=4.715 //y2=4.79
r300 (  73 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.67 //y=1.22 //x2=4.63 //y2=1.375
r301 (  72 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.67 //y=0.875 //x2=4.63 //y2=0.72
r302 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.67 //y=0.875 //x2=4.67 //y2=1.22
r303 (  69 75 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.64 //y=4.865 //x2=4.715 //y2=4.79
r304 (  69 103 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=4.64 //y=4.865 //x2=4.44 //y2=4.7
r305 (  67 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.295 //y=1.375 //x2=4.18 //y2=1.375
r306 (  66 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.515 //y=1.375 //x2=4.63 //y2=1.375
r307 (  65 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.295 //y=0.72 //x2=4.18 //y2=0.72
r308 (  64 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.515 //y=0.72 //x2=4.63 //y2=0.72
r309 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.515 //y=0.72 //x2=4.295 //y2=0.72
r310 (  63 101 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.915 //x2=4.44 //y2=2.08
r311 (  62 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.53 //x2=4.18 //y2=1.375
r312 (  62 63 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.53 //x2=4.14 //y2=1.915
r313 (  61 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.22 //x2=4.18 //y2=1.375
r314 (  60 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=0.875 //x2=4.18 //y2=0.72
r315 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.14 //y=0.875 //x2=4.14 //y2=1.22
r316 (  59 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.89 //y=6.02 //x2=9.89 //y2=4.865
r317 (  58 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.45 //y=6.02 //x2=9.45 //y2=4.865
r318 (  57 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.08 //y=6.02 //x2=5.08 //y2=4.865
r319 (  56 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.64 //y=6.02 //x2=4.64 //y2=4.865
r320 (  55 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.375 //x2=9.325 //y2=1.375
r321 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.375 //x2=9.105 //y2=1.375
r322 (  54 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.405 //y=1.375 //x2=4.515 //y2=1.375
r323 (  54 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.405 //y=1.375 //x2=4.295 //y2=1.375
r324 (  51 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=4.7 //x2=9.25 //y2=4.7
r325 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.59 //x2=9.25 //y2=4.7
r326 (  46 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=2.08 //x2=9.25 //y2=2.08
r327 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.08 //x2=9.25 //y2=2.59
r328 (  43 103 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=4.7 //x2=4.44 //y2=4.7
r329 (  41 43 ) resistor r=144.77 //w=0.187 //l=2.115 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.585 //x2=4.44 //y2=4.7
r330 (  38 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=2.08 //x2=4.44 //y2=2.08
r331 (  38 41 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.08 //x2=4.44 //y2=2.585
r332 (  34 36 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.115 //x2=2.59 //y2=2.59
r333 (  33 36 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=2.59
r334 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r335 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r336 (  30 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.195 //y=5.2 //x2=2.11 //y2=5.2
r337 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.59 //y2=5.115
r338 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.195 //y2=5.2
r339 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.235 //y2=1.655
r340 (  25 114 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r341 (  19 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.2
r342 (  19 117 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.725
r343 (  17 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=2.11 //y2=5.2
r344 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=1.315 //y2=5.2
r345 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.315 //y2=5.2
r346 (  11 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.23 //y2=5.725
r347 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.25 //y=2.59 //x2=9.25 //y2=2.59
r348 (  8 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=2.585 //x2=4.44 //y2=2.585
r349 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=2.59 //x2=2.59 //y2=2.59
r350 (  4 8 ) resistor r=0.164988 //w=0.206 //l=0.267488 //layer=m1 \
 //thickness=0.36 //x=4.705 //y=2.59 //x2=4.44 //y2=2.585
r351 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.135 //y=2.59 //x2=9.25 //y2=2.59
r352 (  3 4 ) resistor r=4.2271 //w=0.131 //l=4.43 //layer=m1 //thickness=0.36 \
 //x=9.135 //y=2.59 //x2=4.705 //y2=2.59
r353 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=2.59 //x2=2.59 //y2=2.59
r354 (  1 8 ) resistor r=0.0921728 //w=0.206 //l=0.147479 //layer=m1 \
 //thickness=0.36 //x=4.295 //y=2.59 //x2=4.44 //y2=2.585
r355 (  1 2 ) resistor r=1.51718 //w=0.131 //l=1.59 //layer=m1 \
 //thickness=0.36 //x=4.295 //y=2.59 //x2=2.705 //y2=2.59
ends PM_DFFSNX1_PCELL\%noxref_3

subckt PM_DFFSNX1_PCELL\%noxref_4 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 61 63 66 67 77 80 82 83 84 )
c160 ( 84 0 ) capacitor c=0.023087f //x=11.285 //y=5.02
c161 ( 83 0 ) capacitor c=0.023519f //x=10.405 //y=5.02
c162 ( 82 0 ) capacitor c=0.0224735f //x=9.525 //y=5.02
c163 ( 80 0 ) capacitor c=0.00872971f //x=11.535 //y=0.915
c164 ( 77 0 ) capacitor c=0.0588816f //x=14.06 //y=4.7
c165 ( 67 0 ) capacitor c=0.0318948f //x=14.395 //y=1.21
c166 ( 66 0 ) capacitor c=0.0187384f //x=14.395 //y=0.865
c167 ( 63 0 ) capacitor c=0.0141798f //x=14.24 //y=1.365
c168 ( 61 0 ) capacitor c=0.0149844f //x=14.24 //y=0.71
c169 ( 57 0 ) capacitor c=0.0813322f //x=13.865 //y=1.915
c170 ( 56 0 ) capacitor c=0.0229267f //x=13.865 //y=1.52
c171 ( 55 0 ) capacitor c=0.0234352f //x=13.865 //y=1.21
c172 ( 54 0 ) capacitor c=0.0199343f //x=13.865 //y=0.865
c173 ( 53 0 ) capacitor c=0.110275f //x=14.4 //y=6.02
c174 ( 52 0 ) capacitor c=0.154305f //x=13.96 //y=6.02
c175 ( 50 0 ) capacitor c=0.00106608f //x=11.43 //y=5.155
c176 ( 49 0 ) capacitor c=0.00207319f //x=10.55 //y=5.155
c177 ( 42 0 ) capacitor c=0.0900192f //x=14.06 //y=2.08
c178 ( 40 0 ) capacitor c=0.110109f //x=12.21 //y=2.59
c179 ( 36 0 ) capacitor c=0.00398962f //x=11.81 //y=1.665
c180 ( 35 0 ) capacitor c=0.0137288f //x=12.125 //y=1.665
c181 ( 29 0 ) capacitor c=0.0284988f //x=12.125 //y=5.155
c182 ( 21 0 ) capacitor c=0.0176454f //x=11.345 //y=5.155
c183 ( 14 0 ) capacitor c=0.00332903f //x=9.755 //y=5.155
c184 ( 13 0 ) capacitor c=0.0148427f //x=10.465 //y=5.155
c185 ( 2 0 ) capacitor c=0.00879187f //x=12.325 //y=2.59
c186 ( 1 0 ) capacitor c=0.0476269f //x=13.945 //y=2.59
r187 (  75 77 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=13.96 //y=4.7 //x2=14.06 //y2=4.7
r188 (  68 77 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=14.4 //y=4.865 //x2=14.06 //y2=4.7
r189 (  67 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.395 //y=1.21 //x2=14.355 //y2=1.365
r190 (  66 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.395 //y=0.865 //x2=14.355 //y2=0.71
r191 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.395 //y=0.865 //x2=14.395 //y2=1.21
r192 (  64 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.02 //y=1.365 //x2=13.905 //y2=1.365
r193 (  63 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.24 //y=1.365 //x2=14.355 //y2=1.365
r194 (  62 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.02 //y=0.71 //x2=13.905 //y2=0.71
r195 (  61 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.24 //y=0.71 //x2=14.355 //y2=0.71
r196 (  61 62 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=14.24 //y=0.71 //x2=14.02 //y2=0.71
r197 (  58 75 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=13.96 //y=4.865 //x2=13.96 //y2=4.7
r198 (  57 72 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.915 //x2=14.06 //y2=2.08
r199 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.52 //x2=13.905 //y2=1.365
r200 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.52 //x2=13.865 //y2=1.915
r201 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.21 //x2=13.905 //y2=1.365
r202 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=0.865 //x2=13.905 //y2=0.71
r203 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.865 //y=0.865 //x2=13.865 //y2=1.21
r204 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.4 //y=6.02 //x2=14.4 //y2=4.865
r205 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.96 //y=6.02 //x2=13.96 //y2=4.865
r206 (  51 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.13 //y=1.365 //x2=14.24 //y2=1.365
r207 (  51 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.13 //y=1.365 //x2=14.02 //y2=1.365
r208 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=4.7 //x2=14.06 //y2=4.7
r209 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.59 //x2=14.06 //y2=4.7
r210 (  42 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=2.08 //x2=14.06 //y2=2.08
r211 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.08 //x2=14.06 //y2=2.59
r212 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=12.21 //y=5.07 //x2=12.21 //y2=2.59
r213 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.75 //x2=12.21 //y2=2.59
r214 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.665 //x2=12.21 //y2=1.75
r215 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.665 //x2=11.81 //y2=1.665
r216 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.725 //y=1.58 //x2=11.81 //y2=1.665
r217 (  31 80 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=11.725 //y=1.58 //x2=11.725 //y2=1.01
r218 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.515 //y=5.155 //x2=11.43 //y2=5.155
r219 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.155 //x2=12.21 //y2=5.07
r220 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.155 //x2=11.515 //y2=5.155
r221 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.43 //y=5.24 //x2=11.43 //y2=5.155
r222 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.43 //y=5.24 //x2=11.43 //y2=5.725
r223 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.635 //y=5.155 //x2=10.55 //y2=5.155
r224 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.345 //y=5.155 //x2=11.43 //y2=5.155
r225 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.345 //y=5.155 //x2=10.635 //y2=5.155
r226 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.55 //y=5.24 //x2=10.55 //y2=5.155
r227 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.55 //y=5.24 //x2=10.55 //y2=5.725
r228 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.465 //y=5.155 //x2=10.55 //y2=5.155
r229 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.465 //y=5.155 //x2=9.755 //y2=5.155
r230 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.67 //y=5.24 //x2=9.755 //y2=5.155
r231 (  7 82 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.67 //y=5.24 //x2=9.67 //y2=5.725
r232 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=2.59 //x2=14.06 //y2=2.59
r233 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.21 //y=2.59 //x2=12.21 //y2=2.59
r234 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.325 //y=2.59 //x2=12.21 //y2=2.59
r235 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=2.59 //x2=14.06 //y2=2.59
r236 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=13.945 //y=2.59 //x2=12.325 //y2=2.59
ends PM_DFFSNX1_PCELL\%noxref_4

subckt PM_DFFSNX1_PCELL\%noxref_5 ( 1 2 8 15 17 23 24 25 26 27 28 29 30 31 33 \
 39 40 41 42 43 48 49 50 55 57 59 65 66 70 79 80 83 )
c198 ( 83 0 ) capacitor c=0.0331838f //x=14.83 //y=4.7
c199 ( 80 0 ) capacitor c=0.0279499f //x=14.8 //y=1.915
c200 ( 79 0 ) capacitor c=0.0425269f //x=14.8 //y=2.08
c201 ( 70 0 ) capacitor c=0.0334842f //x=5.55 //y=4.7
c202 ( 66 0 ) capacitor c=0.0429696f //x=15.365 //y=1.25
c203 ( 65 0 ) capacitor c=0.0192208f //x=15.365 //y=0.905
c204 ( 59 0 ) capacitor c=0.0148884f //x=15.21 //y=1.405
c205 ( 57 0 ) capacitor c=0.0157803f //x=15.21 //y=0.75
c206 ( 55 0 ) capacitor c=0.0299681f //x=15.205 //y=4.79
c207 ( 50 0 ) capacitor c=0.0205163f //x=14.835 //y=1.56
c208 ( 49 0 ) capacitor c=0.0168481f //x=14.835 //y=1.25
c209 ( 48 0 ) capacitor c=0.0174783f //x=14.835 //y=0.905
c210 ( 43 0 ) capacitor c=0.0245352f //x=5.885 //y=4.79
c211 ( 42 0 ) capacitor c=0.0826403f //x=5.64 //y=1.915
c212 ( 41 0 ) capacitor c=0.0170266f //x=5.64 //y=1.45
c213 ( 40 0 ) capacitor c=0.018609f //x=5.64 //y=1.22
c214 ( 39 0 ) capacitor c=0.0187309f //x=5.64 //y=0.91
c215 ( 33 0 ) capacitor c=0.014725f //x=5.485 //y=1.375
c216 ( 31 0 ) capacitor c=0.0146567f //x=5.485 //y=0.755
c217 ( 30 0 ) capacitor c=0.0335408f //x=5.115 //y=1.22
c218 ( 29 0 ) capacitor c=0.0173761f //x=5.115 //y=0.91
c219 ( 28 0 ) capacitor c=0.15358f //x=15.28 //y=6.02
c220 ( 27 0 ) capacitor c=0.110281f //x=14.84 //y=6.02
c221 ( 26 0 ) capacitor c=0.110114f //x=5.96 //y=6.02
c222 ( 25 0 ) capacitor c=0.11012f //x=5.52 //y=6.02
c223 ( 17 0 ) capacitor c=0.0726954f //x=14.8 //y=2.08
c224 ( 15 0 ) capacitor c=0.00369614f //x=14.8 //y=4.535
c225 ( 8 0 ) capacitor c=0.0979973f //x=5.55 //y=2.08
c226 ( 2 0 ) capacitor c=0.0154455f //x=5.665 //y=4.44
c227 ( 1 0 ) capacitor c=0.21665f //x=14.685 //y=4.44
r228 (  85 86 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=14.83 //y=4.79 //x2=14.83 //y2=4.865
r229 (  83 85 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=14.83 //y=4.7 //x2=14.83 //y2=4.79
r230 (  79 80 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=14.8 //y=2.08 //x2=14.8 //y2=1.915
r231 (  72 73 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=5.55 //y=4.79 //x2=5.55 //y2=4.865
r232 (  70 72 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=5.55 //y=4.7 //x2=5.55 //y2=4.79
r233 (  66 90 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.365 //y=1.25 //x2=15.325 //y2=1.405
r234 (  65 89 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.365 //y=0.905 //x2=15.325 //y2=0.75
r235 (  65 66 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.365 //y=0.905 //x2=15.365 //y2=1.25
r236 (  60 88 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.99 //y=1.405 //x2=14.875 //y2=1.405
r237 (  59 90 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.21 //y=1.405 //x2=15.325 //y2=1.405
r238 (  58 87 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.99 //y=0.75 //x2=14.875 //y2=0.75
r239 (  57 89 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.21 //y=0.75 //x2=15.325 //y2=0.75
r240 (  57 58 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.21 //y=0.75 //x2=14.99 //y2=0.75
r241 (  56 85 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=14.965 //y=4.79 //x2=14.83 //y2=4.79
r242 (  55 62 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.79 //x2=15.28 //y2=4.865
r243 (  55 56 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.79 //x2=14.965 //y2=4.79
r244 (  50 88 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.56 //x2=14.875 //y2=1.405
r245 (  50 80 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.56 //x2=14.835 //y2=1.915
r246 (  49 88 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.25 //x2=14.875 //y2=1.405
r247 (  48 87 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=0.905 //x2=14.875 //y2=0.75
r248 (  48 49 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.835 //y=0.905 //x2=14.835 //y2=1.25
r249 (  44 72 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=5.685 //y=4.79 //x2=5.55 //y2=4.79
r250 (  43 45 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.885 //y=4.79 //x2=5.96 //y2=4.865
r251 (  43 44 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=5.885 //y=4.79 //x2=5.685 //y2=4.79
r252 (  42 77 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.915 //x2=5.565 //y2=2.08
r253 (  41 75 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.45 //x2=5.6 //y2=1.375
r254 (  41 42 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.45 //x2=5.64 //y2=1.915
r255 (  40 75 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.22 //x2=5.6 //y2=1.375
r256 (  39 74 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.64 //y=0.91 //x2=5.6 //y2=0.755
r257 (  39 40 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=5.64 //y=0.91 //x2=5.64 //y2=1.22
r258 (  34 68 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.27 //y=1.375 //x2=5.155 //y2=1.375
r259 (  33 75 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.485 //y=1.375 //x2=5.6 //y2=1.375
r260 (  32 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.27 //y=0.755 //x2=5.155 //y2=0.755
r261 (  31 74 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.485 //y=0.755 //x2=5.6 //y2=0.755
r262 (  31 32 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=5.485 //y=0.755 //x2=5.27 //y2=0.755
r263 (  30 68 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.115 //y=1.22 //x2=5.155 //y2=1.375
r264 (  29 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.115 //y=0.91 //x2=5.155 //y2=0.755
r265 (  29 30 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=5.115 //y=0.91 //x2=5.115 //y2=1.22
r266 (  28 62 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.28 //y=6.02 //x2=15.28 //y2=4.865
r267 (  27 86 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.84 //y=6.02 //x2=14.84 //y2=4.865
r268 (  26 45 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.96 //y=6.02 //x2=5.96 //y2=4.865
r269 (  25 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.52 //y=6.02 //x2=5.52 //y2=4.865
r270 (  24 59 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.1 //y=1.405 //x2=15.21 //y2=1.405
r271 (  24 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.1 //y=1.405 //x2=14.99 //y2=1.405
r272 (  23 33 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=5.377 //y=1.375 //x2=5.485 //y2=1.375
r273 (  23 34 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=5.377 //y=1.375 //x2=5.27 //y2=1.375
r274 (  22 83 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.83 //y=4.7 //x2=14.83 //y2=4.7
r275 (  17 79 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.8 //y=2.08 //x2=14.8 //y2=2.08
r276 (  17 20 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=14.8 //y=2.08 //x2=14.8 //y2=4.44
r277 (  15 22 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=14.8 //y=4.535 //x2=14.815 //y2=4.7
r278 (  15 20 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=14.8 //y=4.535 //x2=14.8 //y2=4.44
r279 (  13 70 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=4.7 //x2=5.55 //y2=4.7
r280 (  11 13 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=5.55 //y=4.44 //x2=5.55 //y2=4.7
r281 (  8 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=2.08 //x2=5.55 //y2=2.08
r282 (  8 11 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li //thickness=0.1 \
 //x=5.55 //y=2.08 //x2=5.55 //y2=4.44
r283 (  6 20 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.8 //y=4.44 //x2=14.8 //y2=4.44
r284 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.55 //y=4.44 //x2=5.55 //y2=4.44
r285 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.665 //y=4.44 //x2=5.55 //y2=4.44
r286 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.685 //y=4.44 //x2=14.8 //y2=4.44
r287 (  1 2 ) resistor r=8.60687 //w=0.131 //l=9.02 //layer=m1 \
 //thickness=0.36 //x=14.685 //y=4.44 //x2=5.665 //y2=4.44
ends PM_DFFSNX1_PCELL\%noxref_5

subckt PM_DFFSNX1_PCELL\%noxref_6 ( 1 2 3 4 11 13 23 24 31 39 45 46 50 52 61 \
 62 64 65 67 68 69 70 71 72 73 74 75 80 82 84 90 91 92 93 94 95 99 101 104 105 \
 110 111 114 128 131 133 134 135 )
c285 ( 135 0 ) capacitor c=0.023087f //x=6.475 //y=5.02
c286 ( 134 0 ) capacitor c=0.023519f //x=5.595 //y=5.02
c287 ( 133 0 ) capacitor c=0.0224735f //x=4.715 //y=5.02
c288 ( 131 0 ) capacitor c=0.00853354f //x=6.725 //y=0.915
c289 ( 128 0 ) capacitor c=0.0597793f //x=17.39 //y=4.7
c290 ( 114 0 ) capacitor c=0.0331534f //x=1.88 //y=4.7
c291 ( 111 0 ) capacitor c=0.0279499f //x=1.85 //y=1.915
c292 ( 110 0 ) capacitor c=0.0437302f //x=1.85 //y=2.08
c293 ( 105 0 ) capacitor c=0.0318948f //x=17.725 //y=1.21
c294 ( 104 0 ) capacitor c=0.0187384f //x=17.725 //y=0.865
c295 ( 101 0 ) capacitor c=0.0141798f //x=17.57 //y=1.365
c296 ( 99 0 ) capacitor c=0.0149844f //x=17.57 //y=0.71
c297 ( 95 0 ) capacitor c=0.0813322f //x=17.195 //y=1.915
c298 ( 94 0 ) capacitor c=0.0229267f //x=17.195 //y=1.52
c299 ( 93 0 ) capacitor c=0.0234352f //x=17.195 //y=1.21
c300 ( 92 0 ) capacitor c=0.0199343f //x=17.195 //y=0.865
c301 ( 91 0 ) capacitor c=0.0429696f //x=2.415 //y=1.25
c302 ( 90 0 ) capacitor c=0.0192208f //x=2.415 //y=0.905
c303 ( 84 0 ) capacitor c=0.0158629f //x=2.26 //y=1.405
c304 ( 82 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c305 ( 80 0 ) capacitor c=0.0299681f //x=2.255 //y=4.79
c306 ( 75 0 ) capacitor c=0.0205163f //x=1.885 //y=1.56
c307 ( 74 0 ) capacitor c=0.0168481f //x=1.885 //y=1.25
c308 ( 73 0 ) capacitor c=0.0174783f //x=1.885 //y=0.905
c309 ( 72 0 ) capacitor c=0.110275f //x=17.73 //y=6.02
c310 ( 71 0 ) capacitor c=0.154305f //x=17.29 //y=6.02
c311 ( 70 0 ) capacitor c=0.15358f //x=2.33 //y=6.02
c312 ( 69 0 ) capacitor c=0.110281f //x=1.89 //y=6.02
c313 ( 65 0 ) capacitor c=0.0786338f //x=7.397 //y=3.905
c314 ( 64 0 ) capacitor c=0.0101843f //x=7.395 //y=4.07
c315 ( 62 0 ) capacitor c=0.00106608f //x=6.62 //y=5.155
c316 ( 61 0 ) capacitor c=0.00207162f //x=5.74 //y=5.155
c317 ( 52 0 ) capacitor c=0.0943029f //x=17.39 //y=2.08
c318 ( 50 0 ) capacitor c=0.0236247f //x=7.4 //y=5.07
c319 ( 46 0 ) capacitor c=0.00431225f //x=7 //y=1.665
c320 ( 45 0 ) capacitor c=0.0141453f //x=7.315 //y=1.665
c321 ( 39 0 ) capacitor c=0.0281378f //x=7.315 //y=5.155
c322 ( 31 0 ) capacitor c=0.0176454f //x=6.535 //y=5.155
c323 ( 24 0 ) capacitor c=0.00351598f //x=4.945 //y=5.155
c324 ( 23 0 ) capacitor c=0.0154196f //x=5.655 //y=5.155
c325 ( 13 0 ) capacitor c=0.0787953f //x=1.85 //y=2.08
c326 ( 11 0 ) capacitor c=0.00453889f //x=1.85 //y=4.535
c327 ( 4 0 ) capacitor c=0.00551102f //x=7.51 //y=4.07
c328 ( 3 0 ) capacitor c=0.180782f //x=17.275 //y=4.07
c329 ( 2 0 ) capacitor c=0.0180257f //x=1.965 //y=4.07
c330 ( 1 0 ) capacitor c=0.159166f //x=7.28 //y=4.07
r331 (  126 128 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=17.29 //y=4.7 //x2=17.39 //y2=4.7
r332 (  116 117 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.79 //x2=1.88 //y2=4.865
r333 (  114 116 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.7 //x2=1.88 //y2=4.79
r334 (  110 111 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r335 (  106 128 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=17.73 //y=4.865 //x2=17.39 //y2=4.7
r336 (  105 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.725 //y=1.21 //x2=17.685 //y2=1.365
r337 (  104 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.725 //y=0.865 //x2=17.685 //y2=0.71
r338 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.725 //y=0.865 //x2=17.725 //y2=1.21
r339 (  102 125 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.35 //y=1.365 //x2=17.235 //y2=1.365
r340 (  101 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.57 //y=1.365 //x2=17.685 //y2=1.365
r341 (  100 124 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.35 //y=0.71 //x2=17.235 //y2=0.71
r342 (  99 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.57 //y=0.71 //x2=17.685 //y2=0.71
r343 (  99 100 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.57 //y=0.71 //x2=17.35 //y2=0.71
r344 (  96 126 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.29 //y=4.865 //x2=17.29 //y2=4.7
r345 (  95 123 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.915 //x2=17.39 //y2=2.08
r346 (  94 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.52 //x2=17.235 //y2=1.365
r347 (  94 95 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.52 //x2=17.195 //y2=1.915
r348 (  93 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.21 //x2=17.235 //y2=1.365
r349 (  92 124 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=0.865 //x2=17.235 //y2=0.71
r350 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.195 //y=0.865 //x2=17.195 //y2=1.21
r351 (  91 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r352 (  90 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r353 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r354 (  85 119 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r355 (  84 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r356 (  83 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r357 (  82 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r358 (  82 83 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r359 (  81 116 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.015 //y=4.79 //x2=1.88 //y2=4.79
r360 (  80 87 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.33 //y2=4.865
r361 (  80 81 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.015 //y2=4.79
r362 (  75 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r363 (  75 111 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r364 (  74 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r365 (  73 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r366 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r367 (  72 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.73 //y=6.02 //x2=17.73 //y2=4.865
r368 (  71 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.29 //y=6.02 //x2=17.29 //y2=4.865
r369 (  70 87 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.02 //x2=2.33 //y2=4.865
r370 (  69 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.02 //x2=1.89 //y2=4.865
r371 (  68 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.46 //y=1.365 //x2=17.57 //y2=1.365
r372 (  68 102 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.46 //y=1.365 //x2=17.35 //y2=1.365
r373 (  67 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r374 (  67 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r375 (  64 66 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=7.397 //y=4.07 //x2=7.397 //y2=4.235
r376 (  64 65 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=7.397 //y=4.07 //x2=7.397 //y2=3.905
r377 (  60 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.88 //y=4.7 //x2=1.88 //y2=4.7
r378 (  57 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.39 //y=4.7 //x2=17.39 //y2=4.7
r379 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=17.39 //y=4.07 //x2=17.39 //y2=4.7
r380 (  52 123 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.39 //y=2.08 //x2=17.39 //y2=2.08
r381 (  52 55 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=17.39 //y=2.08 //x2=17.39 //y2=4.07
r382 (  50 66 ) resistor r=57.1551 //w=0.187 //l=0.835 //layer=li \
 //thickness=0.1 //x=7.4 //y=5.07 //x2=7.4 //y2=4.235
r383 (  47 65 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=7.4 //y=1.75 //x2=7.4 //y2=3.905
r384 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.665 //x2=7.4 //y2=1.75
r385 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.665 //x2=7 //y2=1.665
r386 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.915 //y=1.58 //x2=7 //y2=1.665
r387 (  41 131 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=6.915 //y=1.58 //x2=6.915 //y2=1.01
r388 (  40 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.705 //y=5.155 //x2=6.62 //y2=5.155
r389 (  39 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.155 //x2=7.4 //y2=5.07
r390 (  39 40 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.155 //x2=6.705 //y2=5.155
r391 (  33 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.62 //y=5.24 //x2=6.62 //y2=5.155
r392 (  33 135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.62 //y=5.24 //x2=6.62 //y2=5.725
r393 (  32 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.825 //y=5.155 //x2=5.74 //y2=5.155
r394 (  31 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.535 //y=5.155 //x2=6.62 //y2=5.155
r395 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.535 //y=5.155 //x2=5.825 //y2=5.155
r396 (  25 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.74 //y=5.24 //x2=5.74 //y2=5.155
r397 (  25 134 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=5.74 //y=5.24 //x2=5.74 //y2=5.725
r398 (  23 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.655 //y=5.155 //x2=5.74 //y2=5.155
r399 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.655 //y=5.155 //x2=4.945 //y2=5.155
r400 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.86 //y=5.24 //x2=4.945 //y2=5.155
r401 (  17 133 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.86 //y=5.24 //x2=4.86 //y2=5.725
r402 (  13 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r403 (  13 16 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.08 //x2=1.85 //y2=4.07
r404 (  11 60 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.865 //y2=4.7
r405 (  11 16 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.85 //y2=4.07
r406 (  10 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.39 //y=4.07 //x2=17.39 //y2=4.07
r407 (  8 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.395 //y=4.07 //x2=7.395 //y2=4.07
r408 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.85 //y=4.07 //x2=1.85 //y2=4.07
r409 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.51 //y=4.07 //x2=7.395 //y2=4.07
r410 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.275 //y=4.07 //x2=17.39 //y2=4.07
r411 (  3 4 ) resistor r=9.31775 //w=0.131 //l=9.765 //layer=m1 \
 //thickness=0.36 //x=17.275 //y=4.07 //x2=7.51 //y2=4.07
r412 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.965 //y=4.07 //x2=1.85 //y2=4.07
r413 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.28 //y=4.07 //x2=7.395 //y2=4.07
r414 (  1 2 ) resistor r=5.07156 //w=0.131 //l=5.315 //layer=m1 \
 //thickness=0.36 //x=7.28 //y=4.07 //x2=1.965 //y2=4.07
ends PM_DFFSNX1_PCELL\%noxref_6

subckt PM_DFFSNX1_PCELL\%noxref_7 ( 1 2 8 16 23 24 25 26 27 28 29 30 31 33 39 \
 40 41 42 43 48 49 50 52 58 59 60 61 62 70 81 )
c220 ( 81 0 ) capacitor c=0.0337728f //x=21.83 //y=4.7
c221 ( 70 0 ) capacitor c=0.0335551f //x=10.36 //y=4.7
c222 ( 62 0 ) capacitor c=0.025532f //x=22.165 //y=4.79
c223 ( 61 0 ) capacitor c=0.0831166f //x=21.92 //y=1.915
c224 ( 60 0 ) capacitor c=0.0170266f //x=21.92 //y=1.45
c225 ( 59 0 ) capacitor c=0.018609f //x=21.92 //y=1.22
c226 ( 58 0 ) capacitor c=0.0187309f //x=21.92 //y=0.91
c227 ( 52 0 ) capacitor c=0.014725f //x=21.765 //y=1.375
c228 ( 50 0 ) capacitor c=0.0146567f //x=21.765 //y=0.755
c229 ( 49 0 ) capacitor c=0.0335408f //x=21.395 //y=1.22
c230 ( 48 0 ) capacitor c=0.0173761f //x=21.395 //y=0.91
c231 ( 43 0 ) capacitor c=0.0245352f //x=10.695 //y=4.79
c232 ( 42 0 ) capacitor c=0.0826756f //x=10.45 //y=1.915
c233 ( 41 0 ) capacitor c=0.0170266f //x=10.45 //y=1.45
c234 ( 40 0 ) capacitor c=0.018609f //x=10.45 //y=1.22
c235 ( 39 0 ) capacitor c=0.0187309f //x=10.45 //y=0.91
c236 ( 33 0 ) capacitor c=0.014725f //x=10.295 //y=1.375
c237 ( 31 0 ) capacitor c=0.0146567f //x=10.295 //y=0.755
c238 ( 30 0 ) capacitor c=0.0335408f //x=9.925 //y=1.22
c239 ( 29 0 ) capacitor c=0.0173761f //x=9.925 //y=0.91
c240 ( 28 0 ) capacitor c=0.110114f //x=22.24 //y=6.02
c241 ( 27 0 ) capacitor c=0.11012f //x=21.8 //y=6.02
c242 ( 26 0 ) capacitor c=0.110114f //x=10.77 //y=6.02
c243 ( 25 0 ) capacitor c=0.11012f //x=10.33 //y=6.02
c244 ( 16 0 ) capacitor c=0.101396f //x=21.83 //y=2.08
c245 ( 8 0 ) capacitor c=0.094794f //x=10.36 //y=2.08
c246 ( 2 0 ) capacitor c=0.0160685f //x=10.475 //y=2.22
c247 ( 1 0 ) capacitor c=0.309704f //x=21.715 //y=2.22
r248 (  83 84 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=21.83 //y=4.79 //x2=21.83 //y2=4.865
r249 (  81 83 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=21.83 //y=4.7 //x2=21.83 //y2=4.79
r250 (  72 73 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=10.36 //y=4.79 //x2=10.36 //y2=4.865
r251 (  70 72 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=10.36 //y=4.7 //x2=10.36 //y2=4.79
r252 (  63 83 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=21.965 //y=4.79 //x2=21.83 //y2=4.79
r253 (  62 64 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=22.165 //y=4.79 //x2=22.24 //y2=4.865
r254 (  62 63 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=22.165 //y=4.79 //x2=21.965 //y2=4.79
r255 (  61 88 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.915 //x2=21.845 //y2=2.08
r256 (  60 86 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.45 //x2=21.88 //y2=1.375
r257 (  60 61 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.45 //x2=21.92 //y2=1.915
r258 (  59 86 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.22 //x2=21.88 //y2=1.375
r259 (  58 85 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.92 //y=0.91 //x2=21.88 //y2=0.755
r260 (  58 59 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.92 //y=0.91 //x2=21.92 //y2=1.22
r261 (  53 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.375 //x2=21.435 //y2=1.375
r262 (  52 86 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.765 //y=1.375 //x2=21.88 //y2=1.375
r263 (  51 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.755 //x2=21.435 //y2=0.755
r264 (  50 85 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.765 //y=0.755 //x2=21.88 //y2=0.755
r265 (  50 51 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=21.765 //y=0.755 //x2=21.55 //y2=0.755
r266 (  49 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.395 //y=1.22 //x2=21.435 //y2=1.375
r267 (  48 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.91 //x2=21.435 //y2=0.755
r268 (  48 49 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.91 //x2=21.395 //y2=1.22
r269 (  44 72 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=10.495 //y=4.79 //x2=10.36 //y2=4.79
r270 (  43 45 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.695 //y=4.79 //x2=10.77 //y2=4.865
r271 (  43 44 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=10.695 //y=4.79 //x2=10.495 //y2=4.79
r272 (  42 77 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.915 //x2=10.375 //y2=2.08
r273 (  41 75 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.45 //x2=10.41 //y2=1.375
r274 (  41 42 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.45 //x2=10.45 //y2=1.915
r275 (  40 75 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.22 //x2=10.41 //y2=1.375
r276 (  39 74 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.45 //y=0.91 //x2=10.41 //y2=0.755
r277 (  39 40 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=10.45 //y=0.91 //x2=10.45 //y2=1.22
r278 (  34 68 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.08 //y=1.375 //x2=9.965 //y2=1.375
r279 (  33 75 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.295 //y=1.375 //x2=10.41 //y2=1.375
r280 (  32 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.08 //y=0.755 //x2=9.965 //y2=0.755
r281 (  31 74 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.295 //y=0.755 //x2=10.41 //y2=0.755
r282 (  31 32 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=10.295 //y=0.755 //x2=10.08 //y2=0.755
r283 (  30 68 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.925 //y=1.22 //x2=9.965 //y2=1.375
r284 (  29 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.925 //y=0.91 //x2=9.965 //y2=0.755
r285 (  29 30 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=9.925 //y=0.91 //x2=9.925 //y2=1.22
r286 (  28 64 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.24 //y=6.02 //x2=22.24 //y2=4.865
r287 (  27 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.8 //y=6.02 //x2=21.8 //y2=4.865
r288 (  26 45 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.77 //y=6.02 //x2=10.77 //y2=4.865
r289 (  25 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.33 //y=6.02 //x2=10.33 //y2=4.865
r290 (  24 52 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=21.657 //y=1.375 //x2=21.765 //y2=1.375
r291 (  24 53 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=21.657 //y=1.375 //x2=21.55 //y2=1.375
r292 (  23 33 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=10.187 //y=1.375 //x2=10.295 //y2=1.375
r293 (  23 34 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=10.187 //y=1.375 //x2=10.08 //y2=1.375
r294 (  21 81 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.83 //y=4.7 //x2=21.83 //y2=4.7
r295 (  19 21 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.22 //x2=21.83 //y2=4.7
r296 (  16 88 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.83 //y=2.08 //x2=21.83 //y2=2.08
r297 (  16 19 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.08 //x2=21.83 //y2=2.22
r298 (  13 70 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=4.7 //x2=10.36 //y2=4.7
r299 (  11 13 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.22 //x2=10.36 //y2=4.7
r300 (  8 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=2.08 //x2=10.36 //y2=2.08
r301 (  8 11 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.08 //x2=10.36 //y2=2.22
r302 (  6 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.83 //y=2.22 //x2=21.83 //y2=2.22
r303 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=2.22 //x2=10.36 //y2=2.22
r304 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.475 //y=2.22 //x2=10.36 //y2=2.22
r305 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=2.22 //x2=21.83 //y2=2.22
r306 (  1 2 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=2.22 //x2=10.475 //y2=2.22
ends PM_DFFSNX1_PCELL\%noxref_7

subckt PM_DFFSNX1_PCELL\%noxref_8 ( 1 2 3 4 5 6 16 24 37 38 49 51 52 56 58 65 \
 66 67 68 69 70 71 72 73 74 78 79 80 85 87 90 91 95 96 97 102 104 107 108 112 \
 113 114 119 121 124 125 127 128 133 137 138 143 147 148 153 156 158 159 )
c326 ( 159 0 ) capacitor c=0.0220291f //x=14.915 //y=5.02
c327 ( 158 0 ) capacitor c=0.0217503f //x=14.035 //y=5.02
c328 ( 156 0 ) capacitor c=0.00866655f //x=14.91 //y=0.905
c329 ( 153 0 ) capacitor c=0.0617593f //x=22.94 //y=4.7
c330 ( 148 0 ) capacitor c=0.0273931f //x=22.94 //y=1.915
c331 ( 147 0 ) capacitor c=0.0471168f //x=22.94 //y=2.08
c332 ( 143 0 ) capacitor c=0.0587755f //x=11.47 //y=4.7
c333 ( 138 0 ) capacitor c=0.0273931f //x=11.47 //y=1.915
c334 ( 137 0 ) capacitor c=0.0462455f //x=11.47 //y=2.08
c335 ( 133 0 ) capacitor c=0.058931f //x=6.66 //y=4.7
c336 ( 128 0 ) capacitor c=0.0267105f //x=6.66 //y=1.915
c337 ( 127 0 ) capacitor c=0.0457054f //x=6.66 //y=2.08
c338 ( 125 0 ) capacitor c=0.0432517f //x=23.46 //y=1.26
c339 ( 124 0 ) capacitor c=0.0200379f //x=23.46 //y=0.915
c340 ( 121 0 ) capacitor c=0.0158629f //x=23.305 //y=1.415
c341 ( 119 0 ) capacitor c=0.0157803f //x=23.305 //y=0.76
c342 ( 114 0 ) capacitor c=0.0218028f //x=22.93 //y=1.57
c343 ( 113 0 ) capacitor c=0.0207459f //x=22.93 //y=1.26
c344 ( 112 0 ) capacitor c=0.0194308f //x=22.93 //y=0.915
c345 ( 108 0 ) capacitor c=0.0432517f //x=11.99 //y=1.26
c346 ( 107 0 ) capacitor c=0.0200379f //x=11.99 //y=0.915
c347 ( 104 0 ) capacitor c=0.0148873f //x=11.835 //y=1.415
c348 ( 102 0 ) capacitor c=0.0157803f //x=11.835 //y=0.76
c349 ( 97 0 ) capacitor c=0.0218028f //x=11.46 //y=1.57
c350 ( 96 0 ) capacitor c=0.0207459f //x=11.46 //y=1.26
c351 ( 95 0 ) capacitor c=0.0194308f //x=11.46 //y=0.915
c352 ( 91 0 ) capacitor c=0.0432517f //x=7.18 //y=1.26
c353 ( 90 0 ) capacitor c=0.0200379f //x=7.18 //y=0.915
c354 ( 87 0 ) capacitor c=0.0158629f //x=7.025 //y=1.415
c355 ( 85 0 ) capacitor c=0.0157803f //x=7.025 //y=0.76
c356 ( 80 0 ) capacitor c=0.0218028f //x=6.65 //y=1.57
c357 ( 79 0 ) capacitor c=0.0207459f //x=6.65 //y=1.26
c358 ( 78 0 ) capacitor c=0.0194308f //x=6.65 //y=0.915
c359 ( 74 0 ) capacitor c=0.158794f //x=23.12 //y=6.02
c360 ( 73 0 ) capacitor c=0.110114f //x=22.68 //y=6.02
c361 ( 72 0 ) capacitor c=0.158794f //x=11.65 //y=6.02
c362 ( 71 0 ) capacitor c=0.110114f //x=11.21 //y=6.02
c363 ( 70 0 ) capacitor c=0.158048f //x=6.84 //y=6.02
c364 ( 69 0 ) capacitor c=0.110114f //x=6.4 //y=6.02
c365 ( 65 0 ) capacitor c=0.0023043f //x=15.06 //y=5.2
c366 ( 58 0 ) capacitor c=0.0937219f //x=22.94 //y=2.08
c367 ( 56 0 ) capacitor c=0.111199f //x=15.54 //y=3.7
c368 ( 52 0 ) capacitor c=0.00404073f //x=15.185 //y=1.655
c369 ( 51 0 ) capacitor c=0.0122201f //x=15.455 //y=1.655
c370 ( 49 0 ) capacitor c=0.0140462f //x=15.455 //y=5.2
c371 ( 38 0 ) capacitor c=0.00251635f //x=14.265 //y=5.2
c372 ( 37 0 ) capacitor c=0.0143111f //x=14.975 //y=5.2
c373 ( 24 0 ) capacitor c=0.0857928f //x=11.47 //y=2.08
c374 ( 16 0 ) capacitor c=0.0865938f //x=6.66 //y=2.08
c375 ( 6 0 ) capacitor c=0.00472158f //x=15.655 //y=3.7
c376 ( 5 0 ) capacitor c=0.262578f //x=22.825 //y=3.7
c377 ( 4 0 ) capacitor c=0.00493991f //x=11.585 //y=3.7
c378 ( 3 0 ) capacitor c=0.0805272f //x=15.425 //y=3.7
c379 ( 2 0 ) capacitor c=0.0147097f //x=6.775 //y=3.7
c380 ( 1 0 ) capacitor c=0.105064f //x=11.355 //y=3.7
r381 (  147 148 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=22.94 //y=2.08 //x2=22.94 //y2=1.915
r382 (  137 138 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11.47 //y=2.08 //x2=11.47 //y2=1.915
r383 (  127 128 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.66 //y=2.08 //x2=6.66 //y2=1.915
r384 (  125 155 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.46 //y=1.26 //x2=23.42 //y2=1.415
r385 (  124 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.46 //y=0.915 //x2=23.42 //y2=0.76
r386 (  124 125 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.46 //y=0.915 //x2=23.46 //y2=1.26
r387 (  122 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.085 //y=1.415 //x2=22.97 //y2=1.415
r388 (  121 155 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.305 //y=1.415 //x2=23.42 //y2=1.415
r389 (  120 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.085 //y=0.76 //x2=22.97 //y2=0.76
r390 (  119 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.305 //y=0.76 //x2=23.42 //y2=0.76
r391 (  119 120 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=23.305 //y=0.76 //x2=23.085 //y2=0.76
r392 (  116 153 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=23.12 //y=4.865 //x2=22.94 //y2=4.7
r393 (  114 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.57 //x2=22.97 //y2=1.415
r394 (  114 148 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.57 //x2=22.93 //y2=1.915
r395 (  113 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.26 //x2=22.97 //y2=1.415
r396 (  112 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=0.915 //x2=22.97 //y2=0.76
r397 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.93 //y=0.915 //x2=22.93 //y2=1.26
r398 (  109 153 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=22.68 //y=4.865 //x2=22.94 //y2=4.7
r399 (  108 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.99 //y=1.26 //x2=11.95 //y2=1.415
r400 (  107 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.99 //y=0.915 //x2=11.95 //y2=0.76
r401 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.99 //y=0.915 //x2=11.99 //y2=1.26
r402 (  105 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.615 //y=1.415 //x2=11.5 //y2=1.415
r403 (  104 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.835 //y=1.415 //x2=11.95 //y2=1.415
r404 (  103 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.615 //y=0.76 //x2=11.5 //y2=0.76
r405 (  102 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.835 //y=0.76 //x2=11.95 //y2=0.76
r406 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=11.835 //y=0.76 //x2=11.615 //y2=0.76
r407 (  99 143 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=11.65 //y=4.865 //x2=11.47 //y2=4.7
r408 (  97 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.57 //x2=11.5 //y2=1.415
r409 (  97 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.57 //x2=11.46 //y2=1.915
r410 (  96 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.26 //x2=11.5 //y2=1.415
r411 (  95 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=0.915 //x2=11.5 //y2=0.76
r412 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.46 //y=0.915 //x2=11.46 //y2=1.26
r413 (  92 143 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=11.21 //y=4.865 //x2=11.47 //y2=4.7
r414 (  91 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.18 //y=1.26 //x2=7.14 //y2=1.415
r415 (  90 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.18 //y=0.915 //x2=7.14 //y2=0.76
r416 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.18 //y=0.915 //x2=7.18 //y2=1.26
r417 (  88 131 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.805 //y=1.415 //x2=6.69 //y2=1.415
r418 (  87 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.025 //y=1.415 //x2=7.14 //y2=1.415
r419 (  86 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.805 //y=0.76 //x2=6.69 //y2=0.76
r420 (  85 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.025 //y=0.76 //x2=7.14 //y2=0.76
r421 (  85 86 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.025 //y=0.76 //x2=6.805 //y2=0.76
r422 (  82 133 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=6.84 //y=4.865 //x2=6.66 //y2=4.7
r423 (  80 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.57 //x2=6.69 //y2=1.415
r424 (  80 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.57 //x2=6.65 //y2=1.915
r425 (  79 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.26 //x2=6.69 //y2=1.415
r426 (  78 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=0.915 //x2=6.69 //y2=0.76
r427 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.65 //y=0.915 //x2=6.65 //y2=1.26
r428 (  75 133 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=6.4 //y=4.865 //x2=6.66 //y2=4.7
r429 (  74 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.12 //y=6.02 //x2=23.12 //y2=4.865
r430 (  73 109 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.68 //y=6.02 //x2=22.68 //y2=4.865
r431 (  72 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.65 //y=6.02 //x2=11.65 //y2=4.865
r432 (  71 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.21 //y=6.02 //x2=11.21 //y2=4.865
r433 (  70 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.84 //y=6.02 //x2=6.84 //y2=4.865
r434 (  69 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.4 //y=6.02 //x2=6.4 //y2=4.865
r435 (  68 121 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.195 //y=1.415 //x2=23.305 //y2=1.415
r436 (  68 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.195 //y=1.415 //x2=23.085 //y2=1.415
r437 (  67 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.725 //y=1.415 //x2=11.835 //y2=1.415
r438 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.725 //y=1.415 //x2=11.615 //y2=1.415
r439 (  66 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.915 //y=1.415 //x2=7.025 //y2=1.415
r440 (  66 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.915 //y=1.415 //x2=6.805 //y2=1.415
r441 (  63 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.94 //y=4.7 //x2=22.94 //y2=4.7
r442 (  61 63 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=22.94 //y=3.7 //x2=22.94 //y2=4.7
r443 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.94 //y=2.08 //x2=22.94 //y2=2.08
r444 (  58 61 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=22.94 //y=2.08 //x2=22.94 //y2=3.7
r445 (  54 56 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=15.54 //y=5.115 //x2=15.54 //y2=3.7
r446 (  53 56 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=15.54 //y=1.74 //x2=15.54 //y2=3.7
r447 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.455 //y=1.655 //x2=15.54 //y2=1.74
r448 (  51 52 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=15.455 //y=1.655 //x2=15.185 //y2=1.655
r449 (  50 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.145 //y=5.2 //x2=15.06 //y2=5.2
r450 (  49 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.455 //y=5.2 //x2=15.54 //y2=5.115
r451 (  49 50 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=15.455 //y=5.2 //x2=15.145 //y2=5.2
r452 (  45 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.1 //y=1.57 //x2=15.185 //y2=1.655
r453 (  45 156 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=15.1 //y=1.57 //x2=15.1 //y2=1
r454 (  39 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.06 //y=5.285 //x2=15.06 //y2=5.2
r455 (  39 159 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=15.06 //y=5.285 //x2=15.06 //y2=5.725
r456 (  37 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.975 //y=5.2 //x2=15.06 //y2=5.2
r457 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=14.975 //y=5.2 //x2=14.265 //y2=5.2
r458 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.18 //y=5.285 //x2=14.265 //y2=5.2
r459 (  31 158 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=14.18 //y=5.285 //x2=14.18 //y2=5.725
r460 (  29 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=4.7 //x2=11.47 //y2=4.7
r461 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=11.47 //y=3.7 //x2=11.47 //y2=4.7
r462 (  24 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=2.08 //x2=11.47 //y2=2.08
r463 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=11.47 //y=2.08 //x2=11.47 //y2=3.7
r464 (  21 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=4.7 //x2=6.66 //y2=4.7
r465 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=6.66 //y=3.7 //x2=6.66 //y2=4.7
r466 (  16 127 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.08 //x2=6.66 //y2=2.08
r467 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.08 //x2=6.66 //y2=3.7
r468 (  14 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=22.94 //y=3.7 //x2=22.94 //y2=3.7
r469 (  12 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=3.7 //x2=15.54 //y2=3.7
r470 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.47 //y=3.7 //x2=11.47 //y2=3.7
r471 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=3.7 //x2=6.66 //y2=3.7
r472 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.655 //y=3.7 //x2=15.54 //y2=3.7
r473 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=22.825 //y=3.7 //x2=22.94 //y2=3.7
r474 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=22.825 //y=3.7 //x2=15.655 //y2=3.7
r475 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.585 //y=3.7 //x2=11.47 //y2=3.7
r476 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=3.7 //x2=15.54 //y2=3.7
r477 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=3.7 //x2=11.585 //y2=3.7
r478 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.775 //y=3.7 //x2=6.66 //y2=3.7
r479 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=3.7 //x2=11.47 //y2=3.7
r480 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=3.7 //x2=6.775 //y2=3.7
ends PM_DFFSNX1_PCELL\%noxref_8

subckt PM_DFFSNX1_PCELL\%noxref_9 ( 2 7 8 9 10 11 12 13 17 19 22 23 33 )
c57 ( 33 0 ) capacitor c=0.0667949f //x=1.11 //y=4.7
c58 ( 23 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c59 ( 22 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c60 ( 19 0 ) capacitor c=0.0141798f //x=1.29 //y=1.365
c61 ( 17 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c62 ( 13 0 ) capacitor c=0.0860049f //x=0.915 //y=1.915
c63 ( 12 0 ) capacitor c=0.0229722f //x=0.915 //y=1.52
c64 ( 11 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c65 ( 10 0 ) capacitor c=0.0199343f //x=0.915 //y=0.865
c66 ( 9 0 ) capacitor c=0.110275f //x=1.45 //y=6.02
c67 ( 8 0 ) capacitor c=0.154305f //x=1.01 //y=6.02
c68 ( 2 0 ) capacitor c=0.115639f //x=1.11 //y=2.08
r69 (  31 33 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.7 //x2=1.11 //y2=4.7
r70 (  24 33 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=1.45 //y=4.865 //x2=1.11 //y2=4.7
r71 (  23 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r72 (  22 34 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r73 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r74 (  20 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r75 (  19 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r76 (  18 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r77 (  17 34 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r78 (  17 18 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r79 (  14 31 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.865 //x2=1.01 //y2=4.7
r80 (  13 28 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r81 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r82 (  12 13 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r83 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r84 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r85 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r86 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.02 //x2=1.45 //y2=4.865
r87 (  8 14 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.02 //x2=1.01 //y2=4.865
r88 (  7 19 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r89 (  7 20 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r90 (  5 33 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r91 (  2 28 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r92 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=4.7
ends PM_DFFSNX1_PCELL\%noxref_9

subckt PM_DFFSNX1_PCELL\%noxref_10 ( 1 5 9 10 13 17 29 )
c48 ( 29 0 ) capacitor c=0.0632971f //x=0.56 //y=0.365
c49 ( 17 0 ) capacitor c=0.0072343f //x=2.635 //y=0.615
c50 ( 13 0 ) capacitor c=0.015427f //x=2.55 //y=0.53
c51 ( 10 0 ) capacitor c=0.00896024f //x=1.665 //y=1.495
c52 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c53 ( 5 0 ) capacitor c=0.0255599f //x=1.58 //y=1.58
c54 ( 1 0 ) capacitor c=0.0113547f //x=0.695 //y=1.495
r55 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r56 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r57 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r58 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=2.15 //y2=0.53
r59 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r60 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.15 //y2=0.53
r61 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r62 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r63 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r64 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r65 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r66 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r67 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r68 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r69 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r70 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_DFFSNX1_PCELL\%noxref_10

subckt PM_DFFSNX1_PCELL\%noxref_11 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0680128f //x=3.785 //y=0.375
c53 ( 17 0 ) capacitor c=0.018806f //x=5.775 //y=1.59
c54 ( 13 0 ) capacitor c=0.0155484f //x=5.775 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=4.89 //y=0.625
c56 ( 5 0 ) capacitor c=0.017077f //x=4.805 //y=1.59
c57 ( 1 0 ) capacitor c=0.00729042f //x=3.92 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.975 //y=1.59 //x2=4.89 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.975 //y=1.59 //x2=5.375 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.775 //y=1.59 //x2=5.86 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.775 //y=1.59 //x2=5.375 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.975 //y=0.54 //x2=4.89 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.975 //y=0.54 //x2=5.375 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.775 //y=0.54 //x2=5.86 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.775 //y=0.54 //x2=5.375 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.89 //y=1.505 //x2=4.89 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=4.89 //y=1.505 //x2=4.89 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=4.89 //y=0.625 //x2=4.89 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=4.89 //y=0.625 //x2=4.89 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.005 //y=1.59 //x2=3.92 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.005 //y=1.59 //x2=4.405 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.805 //y=1.59 //x2=4.89 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.805 //y=1.59 //x2=4.405 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.92 //y=1.505 //x2=3.92 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=3.92 //y=1.505 //x2=3.92 //y2=0.89
ends PM_DFFSNX1_PCELL\%noxref_11

subckt PM_DFFSNX1_PCELL\%noxref_12 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.041888f //x=6.295 //y=0.375
c54 ( 28 0 ) capacitor c=0.00460056f //x=5.19 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=6.43 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=7.4 //y=0.625
c57 ( 11 0 ) capacitor c=0.0145763f //x=7.315 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=6.43 //y=0.625
c59 ( 1 0 ) capacitor c=0.022894f //x=6.345 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.4 //y=0.625 //x2=7.4 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=7.4 //y=0.625 //x2=7.4 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.515 //y=0.54 //x2=6.43 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.515 //y=0.54 //x2=6.915 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.315 //y=0.54 //x2=7.4 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.315 //y=0.54 //x2=6.915 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.43 //y=1.08 //x2=6.43 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=6.43 //y=1.08 //x2=6.43 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.91 //x2=6.43 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.91 //x2=6.43 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.625 //x2=6.43 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.625 //x2=6.43 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.465 //y=0.995 //x2=5.38 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.345 //y=0.995 //x2=6.43 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=6.345 //y=0.995 //x2=5.465 //y2=0.995
ends PM_DFFSNX1_PCELL\%noxref_12

subckt PM_DFFSNX1_PCELL\%noxref_13 ( 1 5 9 13 17 35 )
c54 ( 35 0 ) capacitor c=0.0685332f //x=8.595 //y=0.375
c55 ( 17 0 ) capacitor c=0.0207646f //x=10.585 //y=1.59
c56 ( 13 0 ) capacitor c=0.0155144f //x=10.585 //y=0.54
c57 ( 9 0 ) capacitor c=0.00678203f //x=9.7 //y=0.625
c58 ( 5 0 ) capacitor c=0.0181938f //x=9.615 //y=1.59
c59 ( 1 0 ) capacitor c=0.00729042f //x=8.73 //y=1.505
r60 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.785 //y=1.59 //x2=9.7 //y2=1.63
r61 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.785 //y=1.59 //x2=10.185 //y2=1.59
r62 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.585 //y=1.59 //x2=10.67 //y2=1.59
r63 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.585 //y=1.59 //x2=10.185 //y2=1.59
r64 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.785 //y=0.54 //x2=9.7 //y2=0.5
r65 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.785 //y=0.54 //x2=10.185 //y2=0.54
r66 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.585 //y=0.54 //x2=10.67 //y2=0.54
r67 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.585 //y=0.54 //x2=10.185 //y2=0.54
r68 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.7 //y=1.505 //x2=9.7 //y2=1.63
r69 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.7 //y=1.505 //x2=9.7 //y2=0.89
r70 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.7 //y=0.625 //x2=9.7 //y2=0.5
r71 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=9.7 //y=0.625 //x2=9.7 //y2=0.89
r72 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.815 //y=1.59 //x2=8.73 //y2=1.63
r73 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.815 //y=1.59 //x2=9.215 //y2=1.59
r74 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.615 //y=1.59 //x2=9.7 //y2=1.63
r75 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.615 //y=1.59 //x2=9.215 //y2=1.59
r76 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.73 //y=1.505 //x2=8.73 //y2=1.63
r77 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.73 //y=1.505 //x2=8.73 //y2=0.89
ends PM_DFFSNX1_PCELL\%noxref_13

subckt PM_DFFSNX1_PCELL\%noxref_14 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0414744f //x=11.105 //y=0.375
c54 ( 28 0 ) capacitor c=0.00461914f //x=10 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=11.24 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=12.21 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144274f //x=12.125 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=11.24 //y=0.625
c59 ( 1 0 ) capacitor c=0.0220663f //x=11.155 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=12.21 //y=0.625 //x2=12.21 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=12.21 //y=0.625 //x2=12.21 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.325 //y=0.54 //x2=11.24 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.325 //y=0.54 //x2=11.725 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.125 //y=0.54 //x2=12.21 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.125 //y=0.54 //x2=11.725 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.24 //y=1.08 //x2=11.24 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=11.24 //y=1.08 //x2=11.24 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.91 //x2=11.24 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.91 //x2=11.24 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.625 //x2=11.24 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.625 //x2=11.24 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.275 //y=0.995 //x2=10.19 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.155 //y=0.995 //x2=11.24 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=11.155 //y=0.995 //x2=10.275 //y2=0.995
ends PM_DFFSNX1_PCELL\%noxref_14

subckt PM_DFFSNX1_PCELL\%noxref_15 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632682f //x=13.51 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=15.585 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=15.5 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=14.615 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=14.615 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=14.53 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=13.645 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=15.585 //y=0.615 //x2=15.585 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.585 //y=0.615 //x2=15.585 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.7 //y=0.53 //x2=14.615 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.7 //y=0.53 //x2=15.1 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.5 //y=0.53 //x2=15.585 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.5 //y=0.53 //x2=15.1 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.615 //y=1.495 //x2=14.615 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=14.615 //y=1.495 //x2=14.615 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=14.615 //y=0.615 //x2=14.615 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=14.615 //y=0.615 //x2=14.615 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.73 //y=1.58 //x2=13.645 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.73 //y=1.58 //x2=14.13 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.53 //y=1.58 //x2=14.615 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.53 //y=1.58 //x2=14.13 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=13.645 //y=1.495 //x2=13.645 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.645 //y=1.495 //x2=13.645 //y2=0.88
ends PM_DFFSNX1_PCELL\%noxref_15

subckt PM_DFFSNX1_PCELL\%noxref_16 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 \
 34 )
c72 ( 34 0 ) capacitor c=0.0332623f //x=18.16 //y=4.7
c73 ( 31 0 ) capacitor c=0.0279499f //x=18.13 //y=1.915
c74 ( 30 0 ) capacitor c=0.0425269f //x=18.13 //y=2.08
c75 ( 28 0 ) capacitor c=0.0429696f //x=18.695 //y=1.25
c76 ( 27 0 ) capacitor c=0.0192208f //x=18.695 //y=0.905
c77 ( 21 0 ) capacitor c=0.0148884f //x=18.54 //y=1.405
c78 ( 19 0 ) capacitor c=0.0157803f //x=18.54 //y=0.75
c79 ( 17 0 ) capacitor c=0.0306375f //x=18.535 //y=4.79
c80 ( 12 0 ) capacitor c=0.0205163f //x=18.165 //y=1.56
c81 ( 11 0 ) capacitor c=0.0168481f //x=18.165 //y=1.25
c82 ( 10 0 ) capacitor c=0.0174783f //x=18.165 //y=0.905
c83 ( 9 0 ) capacitor c=0.15358f //x=18.61 //y=6.02
c84 ( 8 0 ) capacitor c=0.110281f //x=18.17 //y=6.02
c85 ( 3 0 ) capacitor c=0.0772741f //x=18.13 //y=2.08
c86 ( 1 0 ) capacitor c=0.00453889f //x=18.13 //y=4.535
r87 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=18.16 //y=4.79 //x2=18.16 //y2=4.865
r88 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=18.16 //y=4.7 //x2=18.16 //y2=4.79
r89 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=18.13 //y=2.08 //x2=18.13 //y2=1.915
r90 (  28 41 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.695 //y=1.25 //x2=18.655 //y2=1.405
r91 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.695 //y=0.905 //x2=18.655 //y2=0.75
r92 (  27 28 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.695 //y=0.905 //x2=18.695 //y2=1.25
r93 (  22 39 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.32 //y=1.405 //x2=18.205 //y2=1.405
r94 (  21 41 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.54 //y=1.405 //x2=18.655 //y2=1.405
r95 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.32 //y=0.75 //x2=18.205 //y2=0.75
r96 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.54 //y=0.75 //x2=18.655 //y2=0.75
r97 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.54 //y=0.75 //x2=18.32 //y2=0.75
r98 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=18.295 //y=4.79 //x2=18.16 //y2=4.79
r99 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.79 //x2=18.61 //y2=4.865
r100 (  17 18 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.79 //x2=18.295 //y2=4.79
r101 (  12 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.56 //x2=18.205 //y2=1.405
r102 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.56 //x2=18.165 //y2=1.915
r103 (  11 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.25 //x2=18.205 //y2=1.405
r104 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=0.905 //x2=18.205 //y2=0.75
r105 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.165 //y=0.905 //x2=18.165 //y2=1.25
r106 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.61 //y=6.02 //x2=18.61 //y2=4.865
r107 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.17 //y=6.02 //x2=18.17 //y2=4.865
r108 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.43 //y=1.405 //x2=18.54 //y2=1.405
r109 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.43 //y=1.405 //x2=18.32 //y2=1.405
r110 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.16 //y=4.7 //x2=18.16 //y2=4.7
r111 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.13 //y=2.08 //x2=18.13 //y2=2.08
r112 (  1 6 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.535 //x2=18.145 //y2=4.7
r113 (  1 3 ) resistor r=168.043 //w=0.187 //l=2.455 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.535 //x2=18.13 //y2=2.08
ends PM_DFFSNX1_PCELL\%noxref_16

subckt PM_DFFSNX1_PCELL\%noxref_17 ( 7 8 19 21 22 24 25 26 28 29 )
c74 ( 29 0 ) capacitor c=0.0220291f //x=18.245 //y=5.02
c75 ( 28 0 ) capacitor c=0.0217503f //x=17.365 //y=5.02
c76 ( 26 0 ) capacitor c=0.0084702f //x=18.24 //y=0.905
c77 ( 25 0 ) capacitor c=0.0024826f //x=18.39 //y=5.2
c78 ( 24 0 ) capacitor c=0.115479f //x=18.87 //y=5.115
c79 ( 22 0 ) capacitor c=0.00404073f //x=18.515 //y=1.655
c80 ( 21 0 ) capacitor c=0.0122201f //x=18.785 //y=1.655
c81 ( 19 0 ) capacitor c=0.0143719f //x=18.785 //y=5.2
c82 ( 8 0 ) capacitor c=0.00272496f //x=17.595 //y=5.2
c83 ( 7 0 ) capacitor c=0.0155386f //x=18.305 //y=5.2
r84 (  23 24 ) resistor r=231.016 //w=0.187 //l=3.375 //layer=li \
 //thickness=0.1 //x=18.87 //y=1.74 //x2=18.87 //y2=5.115
r85 (  21 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.785 //y=1.655 //x2=18.87 //y2=1.74
r86 (  21 22 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=18.785 //y=1.655 //x2=18.515 //y2=1.655
r87 (  20 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=18.475 //y=5.2 //x2=18.39 //y2=5.2
r88 (  19 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.785 //y=5.2 //x2=18.87 //y2=5.115
r89 (  19 20 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=18.785 //y=5.2 //x2=18.475 //y2=5.2
r90 (  15 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.43 //y=1.57 //x2=18.515 //y2=1.655
r91 (  15 26 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=18.43 //y=1.57 //x2=18.43 //y2=1
r92 (  9 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=18.39 //y=5.285 //x2=18.39 //y2=5.2
r93 (  9 29 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li //thickness=0.1 \
 //x=18.39 //y=5.285 //x2=18.39 //y2=5.725
r94 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=18.305 //y=5.2 //x2=18.39 //y2=5.2
r95 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=18.305 //y=5.2 //x2=17.595 //y2=5.2
r96 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.51 //y=5.285 //x2=17.595 //y2=5.2
r97 (  1 28 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li //thickness=0.1 \
 //x=17.51 //y=5.285 //x2=17.51 //y2=5.725
ends PM_DFFSNX1_PCELL\%noxref_17

subckt PM_DFFSNX1_PCELL\%noxref_18 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632684f //x=16.84 //y=0.365
c53 ( 17 0 ) capacitor c=0.0072343f //x=18.915 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=18.83 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=17.945 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=17.945 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=17.86 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=16.975 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=18.915 //y=0.615 //x2=18.915 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.915 //y=0.615 //x2=18.915 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.03 //y=0.53 //x2=17.945 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.03 //y=0.53 //x2=18.43 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.83 //y=0.53 //x2=18.915 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.83 //y=0.53 //x2=18.43 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=17.945 //y=1.495 //x2=17.945 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=17.945 //y=1.495 //x2=17.945 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=17.945 //y=0.615 //x2=17.945 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=17.945 //y=0.615 //x2=17.945 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.06 //y=1.58 //x2=16.975 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.06 //y=1.58 //x2=17.46 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.86 //y=1.58 //x2=17.945 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.86 //y=1.58 //x2=17.46 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=16.975 //y=1.495 //x2=16.975 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=16.975 //y=1.495 //x2=16.975 //y2=0.88
ends PM_DFFSNX1_PCELL\%noxref_18

subckt PM_DFFSNX1_PCELL\%noxref_19 ( 2 7 8 9 10 11 12 13 14 16 22 23 24 25 )
c61 ( 25 0 ) capacitor c=0.0562318f //x=20.995 //y=4.79
c62 ( 24 0 ) capacitor c=0.0305765f //x=21.285 //y=4.79
c63 ( 23 0 ) capacitor c=0.0347816f //x=20.95 //y=1.22
c64 ( 22 0 ) capacitor c=0.0187487f //x=20.95 //y=0.875
c65 ( 16 0 ) capacitor c=0.0137055f //x=20.795 //y=1.375
c66 ( 14 0 ) capacitor c=0.0149861f //x=20.795 //y=0.72
c67 ( 13 0 ) capacitor c=0.096037f //x=20.42 //y=1.915
c68 ( 12 0 ) capacitor c=0.0228993f //x=20.42 //y=1.53
c69 ( 11 0 ) capacitor c=0.0234352f //x=20.42 //y=1.22
c70 ( 10 0 ) capacitor c=0.0198724f //x=20.42 //y=0.875
c71 ( 9 0 ) capacitor c=0.110114f //x=21.36 //y=6.02
c72 ( 8 0 ) capacitor c=0.158956f //x=20.92 //y=6.02
c73 ( 2 0 ) capacitor c=0.10896f //x=20.72 //y=2.08
r74 (  24 26 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.285 //y=4.79 //x2=21.36 //y2=4.865
r75 (  24 25 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=21.285 //y=4.79 //x2=20.995 //y2=4.79
r76 (  23 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.95 //y=1.22 //x2=20.91 //y2=1.375
r77 (  22 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.95 //y=0.875 //x2=20.91 //y2=0.72
r78 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.95 //y=0.875 //x2=20.95 //y2=1.22
r79 (  19 25 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.92 //y=4.865 //x2=20.995 //y2=4.79
r80 (  19 34 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=20.92 //y=4.865 //x2=20.72 //y2=4.7
r81 (  17 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.575 //y=1.375 //x2=20.46 //y2=1.375
r82 (  16 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.795 //y=1.375 //x2=20.91 //y2=1.375
r83 (  15 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.575 //y=0.72 //x2=20.46 //y2=0.72
r84 (  14 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.795 //y=0.72 //x2=20.91 //y2=0.72
r85 (  14 15 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.795 //y=0.72 //x2=20.575 //y2=0.72
r86 (  13 32 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.915 //x2=20.72 //y2=2.08
r87 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.53 //x2=20.46 //y2=1.375
r88 (  12 13 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.53 //x2=20.42 //y2=1.915
r89 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.22 //x2=20.46 //y2=1.375
r90 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=0.875 //x2=20.46 //y2=0.72
r91 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.42 //y=0.875 //x2=20.42 //y2=1.22
r92 (  9 26 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.36 //y=6.02 //x2=21.36 //y2=4.865
r93 (  8 19 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.92 //y=6.02 //x2=20.92 //y2=4.865
r94 (  7 16 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.685 //y=1.375 //x2=20.795 //y2=1.375
r95 (  7 17 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.685 //y=1.375 //x2=20.575 //y2=1.375
r96 (  5 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.72 //y=4.7 //x2=20.72 //y2=4.7
r97 (  2 32 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.72 //y=2.08 //x2=20.72 //y2=2.08
r98 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=20.72 //y=2.08 //x2=20.72 //y2=4.7
ends PM_DFFSNX1_PCELL\%noxref_19

subckt PM_DFFSNX1_PCELL\%noxref_20 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0686352f //x=20.065 //y=0.375
c51 ( 17 0 ) capacitor c=0.0182323f //x=22.055 //y=1.59
c52 ( 13 0 ) capacitor c=0.0155478f //x=22.055 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=21.17 //y=0.625
c54 ( 5 0 ) capacitor c=0.0164013f //x=21.085 //y=1.59
c55 ( 1 0 ) capacitor c=0.00696517f //x=20.2 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.255 //y=1.59 //x2=21.17 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.255 //y=1.59 //x2=21.655 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.055 //y=1.59 //x2=22.14 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.055 //y=1.59 //x2=21.655 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.255 //y=0.54 //x2=21.17 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.255 //y=0.54 //x2=21.655 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.055 //y=0.54 //x2=22.14 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.055 //y=0.54 //x2=21.655 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=21.17 //y=1.505 //x2=21.17 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=21.17 //y=1.505 //x2=21.17 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=21.17 //y=0.625 //x2=21.17 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=21.17 //y=0.625 //x2=21.17 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.285 //y=1.59 //x2=20.2 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.285 //y=1.59 //x2=20.685 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.085 //y=1.59 //x2=21.17 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.085 //y=1.59 //x2=20.685 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.2 //y=1.505 //x2=20.2 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=20.2 //y=1.505 //x2=20.2 //y2=0.89
ends PM_DFFSNX1_PCELL\%noxref_20

subckt PM_DFFSNX1_PCELL\%noxref_21 ( 7 8 15 23 29 30 32 33 34 35 37 38 39 )
c77 ( 39 0 ) capacitor c=0.023087f //x=22.755 //y=5.02
c78 ( 38 0 ) capacitor c=0.023519f //x=21.875 //y=5.02
c79 ( 37 0 ) capacitor c=0.0224735f //x=20.995 //y=5.02
c80 ( 35 0 ) capacitor c=0.00853354f //x=23.005 //y=0.915
c81 ( 34 0 ) capacitor c=0.00125237f //x=22.9 //y=5.155
c82 ( 33 0 ) capacitor c=0.00243871f //x=22.02 //y=5.155
c83 ( 32 0 ) capacitor c=0.134057f //x=23.68 //y=5.07
c84 ( 30 0 ) capacitor c=0.00777616f //x=23.28 //y=1.665
c85 ( 29 0 ) capacitor c=0.0191287f //x=23.595 //y=1.665
c86 ( 23 0 ) capacitor c=0.0349602f //x=23.595 //y=5.155
c87 ( 15 0 ) capacitor c=0.0191592f //x=22.815 //y=5.155
c88 ( 8 0 ) capacitor c=0.00369455f //x=21.225 //y=5.155
c89 ( 7 0 ) capacitor c=0.0161734f //x=21.935 //y=5.155
r90 (  31 32 ) resistor r=227.251 //w=0.187 //l=3.32 //layer=li \
 //thickness=0.1 //x=23.68 //y=1.75 //x2=23.68 //y2=5.07
r91 (  29 31 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.595 //y=1.665 //x2=23.68 //y2=1.75
r92 (  29 30 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=23.595 //y=1.665 //x2=23.28 //y2=1.665
r93 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.195 //y=1.58 //x2=23.28 //y2=1.665
r94 (  25 35 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=23.195 //y=1.58 //x2=23.195 //y2=1.01
r95 (  24 34 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.985 //y=5.155 //x2=22.9 //y2=5.155
r96 (  23 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.595 //y=5.155 //x2=23.68 //y2=5.07
r97 (  23 24 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li //thickness=0.1 \
 //x=23.595 //y=5.155 //x2=22.985 //y2=5.155
r98 (  17 34 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.9 //y=5.24 //x2=22.9 //y2=5.155
r99 (  17 39 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.9 //y=5.24 //x2=22.9 //y2=5.725
r100 (  16 33 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.105 //y=5.155 //x2=22.02 //y2=5.155
r101 (  15 34 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.815 //y=5.155 //x2=22.9 //y2=5.155
r102 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.815 //y=5.155 //x2=22.105 //y2=5.155
r103 (  9 33 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.02 //y=5.24 //x2=22.02 //y2=5.155
r104 (  9 38 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.02 //y=5.24 //x2=22.02 //y2=5.725
r105 (  7 33 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=21.935 //y=5.155 //x2=22.02 //y2=5.155
r106 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=21.935 //y=5.155 //x2=21.225 //y2=5.155
r107 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.14 //y=5.24 //x2=21.225 //y2=5.155
r108 (  1 37 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.14 //y=5.24 //x2=21.14 //y2=5.725
ends PM_DFFSNX1_PCELL\%noxref_21

subckt PM_DFFSNX1_PCELL\%noxref_22 ( 1 3 11 15 25 28 29 )
c50 ( 29 0 ) capacitor c=0.0429573f //x=22.575 //y=0.375
c51 ( 28 0 ) capacitor c=0.00457437f //x=21.47 //y=0.91
c52 ( 25 0 ) capacitor c=0.00156479f //x=22.71 //y=0.995
c53 ( 15 0 ) capacitor c=0.00737666f //x=23.68 //y=0.625
c54 ( 11 0 ) capacitor c=0.0150034f //x=23.595 //y=0.54
c55 ( 3 0 ) capacitor c=0.00718386f //x=22.71 //y=0.625
c56 ( 1 0 ) capacitor c=0.0246097f //x=22.625 //y=0.995
r57 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.68 //y=0.625 //x2=23.68 //y2=0.5
r58 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=23.68 //y=0.625 //x2=23.68 //y2=0.89
r59 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.795 //y=0.54 //x2=22.71 //y2=0.5
r60 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.795 //y=0.54 //x2=23.195 //y2=0.54
r61 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.595 //y=0.54 //x2=23.68 //y2=0.5
r62 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.595 //y=0.54 //x2=23.195 //y2=0.54
r63 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.71 //y=1.08 //x2=22.71 //y2=0.995
r64 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=22.71 //y=1.08 //x2=22.71 //y2=1.23
r65 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.91 //x2=22.71 //y2=0.995
r66 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.91 //x2=22.71 //y2=0.89
r67 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.625 //x2=22.71 //y2=0.5
r68 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.625 //x2=22.71 //y2=0.89
r69 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.745 //y=0.995 //x2=21.66 //y2=0.995
r70 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.625 //y=0.995 //x2=22.71 //y2=0.995
r71 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=22.625 //y=0.995 //x2=21.745 //y2=0.995
ends PM_DFFSNX1_PCELL\%noxref_22

