* SPICE3 file created from FA.ext - technology: sky130A

.subckt FA SUM COUT A B CIN VDD GND
M1000 a_5767_1050.t4 A.t0 VDD.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_3461_1051.t3 CIN.t0 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_6401_209.t1 a_5767_1050.t5 VDD.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_6858_209.t2 a_6401_209.t3 a_6791_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD.t31 CIN.t1 a_4657_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_575_1051.t2 A.t3 VDD.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 GND a_3027_990.t3 a_3442_101.t0 nshort w=-1.605u l=1.765u
+  ad=10.9968p pd=79.06u as=0p ps=0u
M1007 a_836_209.t3 a_185_209.t3 a_1241_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t7 B.t0 a_807_990.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_6791_1051.t1 a_5291_209.t3 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 COUT a_6858_209.t4 GND.t7 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1011 VDD.t3 a_836_209.t7 a_2795_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VDD.t15 a_836_209.t8 a_2405_209.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_807_990.t1 B.t1 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t9 a_4657_1050.t5 a_5291_209.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_185_209.t2 A.t4 VDD.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_3027_990.t2 CIN.t2 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 SUM.t2 a_3027_990.t4 a_2795_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_3461_1051.t0 a_2405_209.t3 SUM.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 COUT.t2 a_6858_209.t5 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VDD.t14 a_836_209.t9 a_4657_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t6 B.t4 a_5767_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 SUM a_2405_209.t4 a_3442_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.14u as=0p ps=0u
M1023 a_2795_1051.t2 a_836_209.t10 VDD.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VDD.t13 CIN.t4 a_3461_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_575_1051.t0 a_807_990.t3 a_836_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_4657_1050.t1 CIN.t5 VDD.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1241_1051.t1 B.t5 VDD.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 VDD.t2 a_5291_209.t5 a_6791_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 GND CIN.t6 a_4552_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1030 VDD.t16 a_5767_1050.t7 a_6401_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_6791_1051.t3 a_6401_209.t5 a_6858_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 GND a_836_209.t13 a_2776_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_2405_209.t1 a_836_209.t11 VDD.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_4657_1050.t3 a_836_209.t12 VDD.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_836_209.t5 a_807_990.t4 a_575_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_5291_209.t1 a_4657_1050.t6 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1241_1051.t2 a_185_209.t5 a_836_209.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 GND a_807_990.t5 a_1222_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1039 SUM CIN.t8 a_2776_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1040 GND B.t7 a_5662_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1041 VDD.t22 A.t6 a_575_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VDD.t20 A.t7 a_185_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 SUM.t3 a_2405_209.t5 a_3461_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_5767_1050.t1 B.t6 VDD.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 GND A.t2 a_556_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1046 VDD.t26 CIN.t7 a_3027_990.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 VDD.t25 A.t8 a_5767_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_2795_1051.t0 a_3027_990.t5 SUM.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 VDD.t1 B.t8 a_1241_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 VDD.t19 a_6858_209.t6 COUT.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 A B 0.85fF
C1 VDD SUM 0.53fF
C2 A SUM 0.26fF
C3 VDD CIN 0.88fF
C4 A CIN 0.54fF
C5 B SUM 0.24fF
C6 B CIN 1.51fF
C7 SUM CIN 0.62fF
C8 COUT VDD 0.76fF
C9 VDD A 0.58fF
C10 VDD B 1.29fF
R0 A.n5 A.t7 512.525
R1 A.n0 A.t3 480.392
R2 A.n1 A.t8 472.359
R3 A.n0 A.t6 403.272
R4 A.n1 A.t0 384.527
R5 A.n5 A.t4 371.139
R6 A.n6 A.t1 290.093
R7 A.n2 A.n1 213.314
R8 A.n3 A.t2 183.422
R9 A.n3 A.n2 171.69
R10 A.n4 A.n3 156.359
R11 A.n2 A.t5 141.114
R12 A.n6 A.n5 93.541
R13 A.n7 A.n4 77.859
R14 A.n7 A.n6 76
R15 A.n4 A.n0 45.7
R16 A.n7 A 0.046
R17 VDD.n434 VDD.n432 144.705
R18 VDD.n493 VDD.n491 144.705
R19 VDD.n551 VDD.n549 144.705
R20 VDD.n618 VDD.n616 144.705
R21 VDD.n643 VDD.n641 144.705
R22 VDD.n386 VDD.n384 144.705
R23 VDD.n701 VDD.n699 144.705
R24 VDD.n340 VDD.n338 144.705
R25 VDD.n279 VDD.n277 144.705
R26 VDD.n233 VDD.n231 144.705
R27 VDD.n172 VDD.n170 144.705
R28 VDD.n126 VDD.n124 144.705
R29 VDD.n68 VDD.n66 144.705
R30 VDD.n26 VDD.n25 77.792
R31 VDD.n35 VDD.n34 77.792
R32 VDD.n131 VDD.n130 77.792
R33 VDD.n141 VDD.n140 77.792
R34 VDD.n238 VDD.n237 77.792
R35 VDD.n247 VDD.n246 77.792
R36 VDD.n345 VDD.n344 77.792
R37 VDD.n355 VDD.n354 77.792
R38 VDD.n633 VDD.n632 77.792
R39 VDD.n622 VDD.n621 77.792
R40 VDD.n587 VDD.n586 77.792
R41 VDD.n577 VDD.n576 77.792
R42 VDD.n424 VDD.n423 77.792
R43 VDD.n413 VDD.n412 77.792
R44 VDD.n29 VDD.n23 76.145
R45 VDD.n29 VDD.n28 76
R46 VDD.n33 VDD.n32 76
R47 VDD.n39 VDD.n38 76
R48 VDD.n43 VDD.n42 76
R49 VDD.n70 VDD.n69 76
R50 VDD.n74 VDD.n73 76
R51 VDD.n78 VDD.n77 76
R52 VDD.n82 VDD.n81 76
R53 VDD.n87 VDD.n86 76
R54 VDD.n94 VDD.n93 76
R55 VDD.n98 VDD.n97 76
R56 VDD.n102 VDD.n101 76
R57 VDD.n128 VDD.n127 76
R58 VDD.n134 VDD.n133 76
R59 VDD.n138 VDD.n137 76
R60 VDD.n144 VDD.n143 76
R61 VDD.n148 VDD.n147 76
R62 VDD.n174 VDD.n173 76
R63 VDD.n179 VDD.n178 76
R64 VDD.n184 VDD.n183 76
R65 VDD.n190 VDD.n189 76
R66 VDD.n195 VDD.n194 76
R67 VDD.n200 VDD.n199 76
R68 VDD.n205 VDD.n204 76
R69 VDD.n209 VDD.n208 76
R70 VDD.n235 VDD.n234 76
R71 VDD.n241 VDD.n240 76
R72 VDD.n245 VDD.n244 76
R73 VDD.n251 VDD.n250 76
R74 VDD.n255 VDD.n254 76
R75 VDD.n281 VDD.n280 76
R76 VDD.n286 VDD.n285 76
R77 VDD.n291 VDD.n290 76
R78 VDD.n297 VDD.n296 76
R79 VDD.n302 VDD.n301 76
R80 VDD.n307 VDD.n306 76
R81 VDD.n312 VDD.n311 76
R82 VDD.n316 VDD.n315 76
R83 VDD.n342 VDD.n341 76
R84 VDD.n348 VDD.n347 76
R85 VDD.n352 VDD.n351 76
R86 VDD.n358 VDD.n357 76
R87 VDD.n362 VDD.n361 76
R88 VDD.n388 VDD.n387 76
R89 VDD.n752 VDD.n751 76
R90 VDD.n748 VDD.n747 76
R91 VDD.n744 VDD.n743 76
R92 VDD.n740 VDD.n739 76
R93 VDD.n735 VDD.n734 76
R94 VDD.n728 VDD.n727 76
R95 VDD.n724 VDD.n723 76
R96 VDD.n698 VDD.n697 76
R97 VDD.n694 VDD.n693 76
R98 VDD.n690 VDD.n689 76
R99 VDD.n686 VDD.n685 76
R100 VDD.n682 VDD.n681 76
R101 VDD.n677 VDD.n676 76
R102 VDD.n670 VDD.n669 76
R103 VDD.n666 VDD.n665 76
R104 VDD.n640 VDD.n639 76
R105 VDD.n636 VDD.n635 76
R106 VDD.n630 VDD.n629 76
R107 VDD.n626 VDD.n625 76
R108 VDD.n620 VDD.n619 76
R109 VDD.n594 VDD.n593 76
R110 VDD.n590 VDD.n589 76
R111 VDD.n584 VDD.n583 76
R112 VDD.n580 VDD.n579 76
R113 VDD.n574 VDD.n573 76
R114 VDD.n548 VDD.n547 76
R115 VDD.n544 VDD.n543 76
R116 VDD.n540 VDD.n539 76
R117 VDD.n536 VDD.n535 76
R118 VDD.n532 VDD.n531 76
R119 VDD.n527 VDD.n526 76
R120 VDD.n520 VDD.n519 76
R121 VDD.n516 VDD.n515 76
R122 VDD.n490 VDD.n489 76
R123 VDD.n486 VDD.n485 76
R124 VDD.n482 VDD.n481 76
R125 VDD.n478 VDD.n477 76
R126 VDD.n474 VDD.n473 76
R127 VDD.n469 VDD.n468 76
R128 VDD.n462 VDD.n461 76
R129 VDD.n458 VDD.n457 76
R130 VDD.n431 VDD.n430 76
R131 VDD.n427 VDD.n426 76
R132 VDD.n421 VDD.n420 76
R133 VDD.n417 VDD.n416 76
R134 VDD.n411 VDD.n410 76
R135 VDD.n464 VDD.n463 65.585
R136 VDD.n522 VDD.n521 65.585
R137 VDD.n672 VDD.n671 65.585
R138 VDD.n730 VDD.n729 65.585
R139 VDD.n415 VDD.t21 55.106
R140 VDD.n422 VDD.t20 55.106
R141 VDD.n575 VDD.t18 55.106
R142 VDD.n585 VDD.t7 55.106
R143 VDD.n624 VDD.t29 55.106
R144 VDD.n631 VDD.t15 55.106
R145 VDD.n353 VDD.t5 55.106
R146 VDD.n343 VDD.t26 55.106
R147 VDD.n308 VDD.t10 55.106
R148 VDD.n249 VDD.t4 55.106
R149 VDD.n236 VDD.t9 55.106
R150 VDD.n201 VDD.t11 55.106
R151 VDD.n139 VDD.t30 55.106
R152 VDD.n129 VDD.t16 55.106
R153 VDD.n37 VDD.t12 55.106
R154 VDD.n24 VDD.t19 55.106
R155 VDD.n282 VDD.t14 55.106
R156 VDD.n177 VDD.t25 55.106
R157 VDD.n89 VDD.n88 41.183
R158 VDD.n293 VDD.n292 40.824
R159 VDD.n188 VDD.n187 40.824
R160 VDD.n498 VDD.n497 36.774
R161 VDD.n556 VDD.n555 36.774
R162 VDD.n599 VDD.n598 36.774
R163 VDD.n648 VDD.n647 36.774
R164 VDD.n706 VDD.n705 36.774
R165 VDD.n367 VDD.n366 36.774
R166 VDD.n321 VDD.n320 36.774
R167 VDD.n260 VDD.n259 36.774
R168 VDD.n214 VDD.n213 36.774
R169 VDD.n153 VDD.n152 36.774
R170 VDD.n107 VDD.n106 36.774
R171 VDD.n48 VDD.n47 36.774
R172 VDD.n450 VDD.n449 36.774
R173 VDD.n181 VDD.n180 36.608
R174 VDD.n288 VDD.n287 36.608
R175 VDD.n91 VDD.n90 32.032
R176 VDD.n197 VDD.n196 32.032
R177 VDD.n304 VDD.n303 32.032
R178 VDD.n732 VDD.n731 32.032
R179 VDD.n674 VDD.n673 32.032
R180 VDD.n524 VDD.n523 32.032
R181 VDD.n466 VDD.n465 32.032
R182 VDD.n410 VDD.n407 21.841
R183 VDD.n23 VDD.n20 21.841
R184 VDD.n463 VDD.t24 14.282
R185 VDD.n463 VDD.t22 14.282
R186 VDD.n521 VDD.t17 14.282
R187 VDD.n521 VDD.t1 14.282
R188 VDD.n671 VDD.t27 14.282
R189 VDD.n671 VDD.t3 14.282
R190 VDD.n729 VDD.t0 14.282
R191 VDD.n729 VDD.t13 14.282
R192 VDD.n292 VDD.t28 14.282
R193 VDD.n292 VDD.t31 14.282
R194 VDD.n187 VDD.t23 14.282
R195 VDD.n187 VDD.t6 14.282
R196 VDD.n88 VDD.t8 14.282
R197 VDD.n88 VDD.t2 14.282
R198 VDD.n407 VDD.n390 14.167
R199 VDD.n390 VDD.n389 14.167
R200 VDD.n513 VDD.n495 14.167
R201 VDD.n495 VDD.n494 14.167
R202 VDD.n571 VDD.n553 14.167
R203 VDD.n553 VDD.n552 14.167
R204 VDD.n614 VDD.n596 14.167
R205 VDD.n596 VDD.n595 14.167
R206 VDD.n663 VDD.n645 14.167
R207 VDD.n645 VDD.n644 14.167
R208 VDD.n721 VDD.n703 14.167
R209 VDD.n703 VDD.n702 14.167
R210 VDD.n382 VDD.n364 14.167
R211 VDD.n364 VDD.n363 14.167
R212 VDD.n336 VDD.n318 14.167
R213 VDD.n318 VDD.n317 14.167
R214 VDD.n275 VDD.n257 14.167
R215 VDD.n257 VDD.n256 14.167
R216 VDD.n229 VDD.n211 14.167
R217 VDD.n211 VDD.n210 14.167
R218 VDD.n168 VDD.n150 14.167
R219 VDD.n150 VDD.n149 14.167
R220 VDD.n122 VDD.n104 14.167
R221 VDD.n104 VDD.n103 14.167
R222 VDD.n64 VDD.n45 14.167
R223 VDD.n45 VDD.n44 14.167
R224 VDD.n455 VDD.n436 14.167
R225 VDD.n436 VDD.n435 14.167
R226 VDD.n20 VDD.n19 14.167
R227 VDD.n19 VDD.n17 14.167
R228 VDD.n69 VDD.n65 14.167
R229 VDD.n127 VDD.n123 14.167
R230 VDD.n173 VDD.n169 14.167
R231 VDD.n234 VDD.n230 14.167
R232 VDD.n280 VDD.n276 14.167
R233 VDD.n341 VDD.n337 14.167
R234 VDD.n387 VDD.n383 14.167
R235 VDD.n723 VDD.n722 14.167
R236 VDD.n665 VDD.n664 14.167
R237 VDD.n619 VDD.n615 14.167
R238 VDD.n573 VDD.n572 14.167
R239 VDD.n515 VDD.n514 14.167
R240 VDD.n457 VDD.n456 14.167
R241 VDD.n23 VDD.n22 13.653
R242 VDD.n22 VDD.n21 13.653
R243 VDD.n28 VDD.n27 13.653
R244 VDD.n27 VDD.n26 13.653
R245 VDD.n32 VDD.n31 13.653
R246 VDD.n31 VDD.n30 13.653
R247 VDD.n38 VDD.n36 13.653
R248 VDD.n36 VDD.n35 13.653
R249 VDD.n42 VDD.n41 13.653
R250 VDD.n41 VDD.n40 13.653
R251 VDD.n69 VDD.n68 13.653
R252 VDD.n68 VDD.n67 13.653
R253 VDD.n73 VDD.n72 13.653
R254 VDD.n72 VDD.n71 13.653
R255 VDD.n77 VDD.n76 13.653
R256 VDD.n76 VDD.n75 13.653
R257 VDD.n81 VDD.n80 13.653
R258 VDD.n80 VDD.n79 13.653
R259 VDD.n86 VDD.n85 13.653
R260 VDD.n85 VDD.n84 13.653
R261 VDD.n93 VDD.n92 13.653
R262 VDD.n92 VDD.n91 13.653
R263 VDD.n97 VDD.n96 13.653
R264 VDD.n96 VDD.n95 13.653
R265 VDD.n101 VDD.n100 13.653
R266 VDD.n100 VDD.n99 13.653
R267 VDD.n127 VDD.n126 13.653
R268 VDD.n126 VDD.n125 13.653
R269 VDD.n133 VDD.n132 13.653
R270 VDD.n132 VDD.n131 13.653
R271 VDD.n137 VDD.n136 13.653
R272 VDD.n136 VDD.n135 13.653
R273 VDD.n143 VDD.n142 13.653
R274 VDD.n142 VDD.n141 13.653
R275 VDD.n147 VDD.n146 13.653
R276 VDD.n146 VDD.n145 13.653
R277 VDD.n173 VDD.n172 13.653
R278 VDD.n172 VDD.n171 13.653
R279 VDD.n178 VDD.n176 13.653
R280 VDD.n176 VDD.n175 13.653
R281 VDD.n183 VDD.n182 13.653
R282 VDD.n182 VDD.n181 13.653
R283 VDD.n189 VDD.n186 13.653
R284 VDD.n186 VDD.n185 13.653
R285 VDD.n194 VDD.n193 13.653
R286 VDD.n193 VDD.n192 13.653
R287 VDD.n199 VDD.n198 13.653
R288 VDD.n198 VDD.n197 13.653
R289 VDD.n204 VDD.n203 13.653
R290 VDD.n203 VDD.n202 13.653
R291 VDD.n208 VDD.n207 13.653
R292 VDD.n207 VDD.n206 13.653
R293 VDD.n234 VDD.n233 13.653
R294 VDD.n233 VDD.n232 13.653
R295 VDD.n240 VDD.n239 13.653
R296 VDD.n239 VDD.n238 13.653
R297 VDD.n244 VDD.n243 13.653
R298 VDD.n243 VDD.n242 13.653
R299 VDD.n250 VDD.n248 13.653
R300 VDD.n248 VDD.n247 13.653
R301 VDD.n254 VDD.n253 13.653
R302 VDD.n253 VDD.n252 13.653
R303 VDD.n280 VDD.n279 13.653
R304 VDD.n279 VDD.n278 13.653
R305 VDD.n285 VDD.n284 13.653
R306 VDD.n284 VDD.n283 13.653
R307 VDD.n290 VDD.n289 13.653
R308 VDD.n289 VDD.n288 13.653
R309 VDD.n296 VDD.n295 13.653
R310 VDD.n295 VDD.n294 13.653
R311 VDD.n301 VDD.n300 13.653
R312 VDD.n300 VDD.n299 13.653
R313 VDD.n306 VDD.n305 13.653
R314 VDD.n305 VDD.n304 13.653
R315 VDD.n311 VDD.n310 13.653
R316 VDD.n310 VDD.n309 13.653
R317 VDD.n315 VDD.n314 13.653
R318 VDD.n314 VDD.n313 13.653
R319 VDD.n341 VDD.n340 13.653
R320 VDD.n340 VDD.n339 13.653
R321 VDD.n347 VDD.n346 13.653
R322 VDD.n346 VDD.n345 13.653
R323 VDD.n351 VDD.n350 13.653
R324 VDD.n350 VDD.n349 13.653
R325 VDD.n357 VDD.n356 13.653
R326 VDD.n356 VDD.n355 13.653
R327 VDD.n361 VDD.n360 13.653
R328 VDD.n360 VDD.n359 13.653
R329 VDD.n387 VDD.n386 13.653
R330 VDD.n386 VDD.n385 13.653
R331 VDD.n751 VDD.n750 13.653
R332 VDD.n750 VDD.n749 13.653
R333 VDD.n747 VDD.n746 13.653
R334 VDD.n746 VDD.n745 13.653
R335 VDD.n743 VDD.n742 13.653
R336 VDD.n742 VDD.n741 13.653
R337 VDD.n739 VDD.n738 13.653
R338 VDD.n738 VDD.n737 13.653
R339 VDD.n734 VDD.n733 13.653
R340 VDD.n733 VDD.n732 13.653
R341 VDD.n727 VDD.n726 13.653
R342 VDD.n726 VDD.n725 13.653
R343 VDD.n723 VDD.n701 13.653
R344 VDD.n701 VDD.n700 13.653
R345 VDD.n697 VDD.n696 13.653
R346 VDD.n696 VDD.n695 13.653
R347 VDD.n693 VDD.n692 13.653
R348 VDD.n692 VDD.n691 13.653
R349 VDD.n689 VDD.n688 13.653
R350 VDD.n688 VDD.n687 13.653
R351 VDD.n685 VDD.n684 13.653
R352 VDD.n684 VDD.n683 13.653
R353 VDD.n681 VDD.n680 13.653
R354 VDD.n680 VDD.n679 13.653
R355 VDD.n676 VDD.n675 13.653
R356 VDD.n675 VDD.n674 13.653
R357 VDD.n669 VDD.n668 13.653
R358 VDD.n668 VDD.n667 13.653
R359 VDD.n665 VDD.n643 13.653
R360 VDD.n643 VDD.n642 13.653
R361 VDD.n639 VDD.n638 13.653
R362 VDD.n638 VDD.n637 13.653
R363 VDD.n635 VDD.n634 13.653
R364 VDD.n634 VDD.n633 13.653
R365 VDD.n629 VDD.n628 13.653
R366 VDD.n628 VDD.n627 13.653
R367 VDD.n625 VDD.n623 13.653
R368 VDD.n623 VDD.n622 13.653
R369 VDD.n619 VDD.n618 13.653
R370 VDD.n618 VDD.n617 13.653
R371 VDD.n593 VDD.n592 13.653
R372 VDD.n592 VDD.n591 13.653
R373 VDD.n589 VDD.n588 13.653
R374 VDD.n588 VDD.n587 13.653
R375 VDD.n583 VDD.n582 13.653
R376 VDD.n582 VDD.n581 13.653
R377 VDD.n579 VDD.n578 13.653
R378 VDD.n578 VDD.n577 13.653
R379 VDD.n573 VDD.n551 13.653
R380 VDD.n551 VDD.n550 13.653
R381 VDD.n547 VDD.n546 13.653
R382 VDD.n546 VDD.n545 13.653
R383 VDD.n543 VDD.n542 13.653
R384 VDD.n542 VDD.n541 13.653
R385 VDD.n539 VDD.n538 13.653
R386 VDD.n538 VDD.n537 13.653
R387 VDD.n535 VDD.n534 13.653
R388 VDD.n534 VDD.n533 13.653
R389 VDD.n531 VDD.n530 13.653
R390 VDD.n530 VDD.n529 13.653
R391 VDD.n526 VDD.n525 13.653
R392 VDD.n525 VDD.n524 13.653
R393 VDD.n519 VDD.n518 13.653
R394 VDD.n518 VDD.n517 13.653
R395 VDD.n515 VDD.n493 13.653
R396 VDD.n493 VDD.n492 13.653
R397 VDD.n489 VDD.n488 13.653
R398 VDD.n488 VDD.n487 13.653
R399 VDD.n485 VDD.n484 13.653
R400 VDD.n484 VDD.n483 13.653
R401 VDD.n481 VDD.n480 13.653
R402 VDD.n480 VDD.n479 13.653
R403 VDD.n477 VDD.n476 13.653
R404 VDD.n476 VDD.n475 13.653
R405 VDD.n473 VDD.n472 13.653
R406 VDD.n472 VDD.n471 13.653
R407 VDD.n468 VDD.n467 13.653
R408 VDD.n467 VDD.n466 13.653
R409 VDD.n461 VDD.n460 13.653
R410 VDD.n460 VDD.n459 13.653
R411 VDD.n457 VDD.n434 13.653
R412 VDD.n434 VDD.n433 13.653
R413 VDD.n430 VDD.n429 13.653
R414 VDD.n429 VDD.n428 13.653
R415 VDD.n426 VDD.n425 13.653
R416 VDD.n425 VDD.n424 13.653
R417 VDD.n420 VDD.n419 13.653
R418 VDD.n419 VDD.n418 13.653
R419 VDD.n416 VDD.n414 13.653
R420 VDD.n414 VDD.n413 13.653
R421 VDD.n410 VDD.n409 13.653
R422 VDD.n409 VDD.n408 13.653
R423 VDD.n4 VDD.n2 12.915
R424 VDD.n4 VDD.n3 12.66
R425 VDD.n12 VDD.n11 12.343
R426 VDD.n12 VDD.n9 12.343
R427 VDD.n7 VDD.n6 12.343
R428 VDD.n189 VDD.n188 8.658
R429 VDD.n296 VDD.n293 8.658
R430 VDD.n514 VDD.n513 7.674
R431 VDD.n572 VDD.n571 7.674
R432 VDD.n615 VDD.n614 7.674
R433 VDD.n664 VDD.n663 7.674
R434 VDD.n722 VDD.n721 7.674
R435 VDD.n383 VDD.n382 7.674
R436 VDD.n337 VDD.n336 7.674
R437 VDD.n276 VDD.n275 7.674
R438 VDD.n230 VDD.n229 7.674
R439 VDD.n169 VDD.n168 7.674
R440 VDD.n123 VDD.n122 7.674
R441 VDD.n65 VDD.n64 7.674
R442 VDD.n456 VDD.n455 7.674
R443 VDD.n59 VDD.n58 7.5
R444 VDD.n53 VDD.n52 7.5
R445 VDD.n55 VDD.n54 7.5
R446 VDD.n50 VDD.n49 7.5
R447 VDD.n64 VDD.n63 7.5
R448 VDD.n117 VDD.n116 7.5
R449 VDD.n111 VDD.n110 7.5
R450 VDD.n113 VDD.n112 7.5
R451 VDD.n119 VDD.n109 7.5
R452 VDD.n119 VDD.n107 7.5
R453 VDD.n122 VDD.n121 7.5
R454 VDD.n163 VDD.n162 7.5
R455 VDD.n157 VDD.n156 7.5
R456 VDD.n159 VDD.n158 7.5
R457 VDD.n165 VDD.n155 7.5
R458 VDD.n165 VDD.n153 7.5
R459 VDD.n168 VDD.n167 7.5
R460 VDD.n224 VDD.n223 7.5
R461 VDD.n218 VDD.n217 7.5
R462 VDD.n220 VDD.n219 7.5
R463 VDD.n226 VDD.n216 7.5
R464 VDD.n226 VDD.n214 7.5
R465 VDD.n229 VDD.n228 7.5
R466 VDD.n270 VDD.n269 7.5
R467 VDD.n264 VDD.n263 7.5
R468 VDD.n266 VDD.n265 7.5
R469 VDD.n272 VDD.n262 7.5
R470 VDD.n272 VDD.n260 7.5
R471 VDD.n275 VDD.n274 7.5
R472 VDD.n331 VDD.n330 7.5
R473 VDD.n325 VDD.n324 7.5
R474 VDD.n327 VDD.n326 7.5
R475 VDD.n333 VDD.n323 7.5
R476 VDD.n333 VDD.n321 7.5
R477 VDD.n336 VDD.n335 7.5
R478 VDD.n377 VDD.n376 7.5
R479 VDD.n371 VDD.n370 7.5
R480 VDD.n373 VDD.n372 7.5
R481 VDD.n379 VDD.n369 7.5
R482 VDD.n379 VDD.n367 7.5
R483 VDD.n382 VDD.n381 7.5
R484 VDD.n716 VDD.n715 7.5
R485 VDD.n710 VDD.n709 7.5
R486 VDD.n712 VDD.n711 7.5
R487 VDD.n718 VDD.n708 7.5
R488 VDD.n718 VDD.n706 7.5
R489 VDD.n721 VDD.n720 7.5
R490 VDD.n658 VDD.n657 7.5
R491 VDD.n652 VDD.n651 7.5
R492 VDD.n654 VDD.n653 7.5
R493 VDD.n660 VDD.n650 7.5
R494 VDD.n660 VDD.n648 7.5
R495 VDD.n663 VDD.n662 7.5
R496 VDD.n609 VDD.n608 7.5
R497 VDD.n603 VDD.n602 7.5
R498 VDD.n605 VDD.n604 7.5
R499 VDD.n611 VDD.n601 7.5
R500 VDD.n611 VDD.n599 7.5
R501 VDD.n614 VDD.n613 7.5
R502 VDD.n566 VDD.n565 7.5
R503 VDD.n560 VDD.n559 7.5
R504 VDD.n562 VDD.n561 7.5
R505 VDD.n568 VDD.n558 7.5
R506 VDD.n568 VDD.n556 7.5
R507 VDD.n571 VDD.n570 7.5
R508 VDD.n508 VDD.n507 7.5
R509 VDD.n502 VDD.n501 7.5
R510 VDD.n504 VDD.n503 7.5
R511 VDD.n510 VDD.n500 7.5
R512 VDD.n510 VDD.n498 7.5
R513 VDD.n513 VDD.n512 7.5
R514 VDD.n440 VDD.n439 7.5
R515 VDD.n443 VDD.n442 7.5
R516 VDD.n445 VDD.n444 7.5
R517 VDD.n448 VDD.n447 7.5
R518 VDD.n455 VDD.n454 7.5
R519 VDD.n402 VDD.n401 7.5
R520 VDD.n396 VDD.n395 7.5
R521 VDD.n398 VDD.n397 7.5
R522 VDD.n404 VDD.n394 7.5
R523 VDD.n404 VDD.n392 7.5
R524 VDD.n407 VDD.n406 7.5
R525 VDD.n20 VDD.n16 7.5
R526 VDD.n2 VDD.n1 7.5
R527 VDD.n6 VDD.n5 7.5
R528 VDD.n11 VDD.n10 7.5
R529 VDD.n19 VDD.n18 7.5
R530 VDD.n14 VDD.n0 7.5
R531 VDD.n51 VDD.n48 6.772
R532 VDD.n62 VDD.n46 6.772
R533 VDD.n60 VDD.n57 6.772
R534 VDD.n56 VDD.n53 6.772
R535 VDD.n120 VDD.n105 6.772
R536 VDD.n118 VDD.n115 6.772
R537 VDD.n114 VDD.n111 6.772
R538 VDD.n166 VDD.n151 6.772
R539 VDD.n164 VDD.n161 6.772
R540 VDD.n160 VDD.n157 6.772
R541 VDD.n227 VDD.n212 6.772
R542 VDD.n225 VDD.n222 6.772
R543 VDD.n221 VDD.n218 6.772
R544 VDD.n273 VDD.n258 6.772
R545 VDD.n271 VDD.n268 6.772
R546 VDD.n267 VDD.n264 6.772
R547 VDD.n334 VDD.n319 6.772
R548 VDD.n332 VDD.n329 6.772
R549 VDD.n328 VDD.n325 6.772
R550 VDD.n380 VDD.n365 6.772
R551 VDD.n378 VDD.n375 6.772
R552 VDD.n374 VDD.n371 6.772
R553 VDD.n719 VDD.n704 6.772
R554 VDD.n717 VDD.n714 6.772
R555 VDD.n713 VDD.n710 6.772
R556 VDD.n661 VDD.n646 6.772
R557 VDD.n659 VDD.n656 6.772
R558 VDD.n655 VDD.n652 6.772
R559 VDD.n612 VDD.n597 6.772
R560 VDD.n610 VDD.n607 6.772
R561 VDD.n606 VDD.n603 6.772
R562 VDD.n569 VDD.n554 6.772
R563 VDD.n567 VDD.n564 6.772
R564 VDD.n563 VDD.n560 6.772
R565 VDD.n511 VDD.n496 6.772
R566 VDD.n509 VDD.n506 6.772
R567 VDD.n505 VDD.n502 6.772
R568 VDD.n405 VDD.n391 6.772
R569 VDD.n403 VDD.n400 6.772
R570 VDD.n399 VDD.n396 6.772
R571 VDD.n51 VDD.n50 6.772
R572 VDD.n56 VDD.n55 6.772
R573 VDD.n60 VDD.n59 6.772
R574 VDD.n63 VDD.n62 6.772
R575 VDD.n114 VDD.n113 6.772
R576 VDD.n118 VDD.n117 6.772
R577 VDD.n121 VDD.n120 6.772
R578 VDD.n160 VDD.n159 6.772
R579 VDD.n164 VDD.n163 6.772
R580 VDD.n167 VDD.n166 6.772
R581 VDD.n221 VDD.n220 6.772
R582 VDD.n225 VDD.n224 6.772
R583 VDD.n228 VDD.n227 6.772
R584 VDD.n267 VDD.n266 6.772
R585 VDD.n271 VDD.n270 6.772
R586 VDD.n274 VDD.n273 6.772
R587 VDD.n328 VDD.n327 6.772
R588 VDD.n332 VDD.n331 6.772
R589 VDD.n335 VDD.n334 6.772
R590 VDD.n374 VDD.n373 6.772
R591 VDD.n378 VDD.n377 6.772
R592 VDD.n381 VDD.n380 6.772
R593 VDD.n713 VDD.n712 6.772
R594 VDD.n717 VDD.n716 6.772
R595 VDD.n720 VDD.n719 6.772
R596 VDD.n655 VDD.n654 6.772
R597 VDD.n659 VDD.n658 6.772
R598 VDD.n662 VDD.n661 6.772
R599 VDD.n606 VDD.n605 6.772
R600 VDD.n610 VDD.n609 6.772
R601 VDD.n613 VDD.n612 6.772
R602 VDD.n563 VDD.n562 6.772
R603 VDD.n567 VDD.n566 6.772
R604 VDD.n570 VDD.n569 6.772
R605 VDD.n505 VDD.n504 6.772
R606 VDD.n509 VDD.n508 6.772
R607 VDD.n512 VDD.n511 6.772
R608 VDD.n399 VDD.n398 6.772
R609 VDD.n403 VDD.n402 6.772
R610 VDD.n406 VDD.n405 6.772
R611 VDD.n454 VDD.n453 6.772
R612 VDD.n441 VDD.n438 6.772
R613 VDD.n446 VDD.n443 6.772
R614 VDD.n451 VDD.n448 6.772
R615 VDD.n451 VDD.n450 6.772
R616 VDD.n446 VDD.n445 6.772
R617 VDD.n441 VDD.n440 6.772
R618 VDD.n453 VDD.n437 6.772
R619 VDD.n16 VDD.n15 6.458
R620 VDD.n109 VDD.n108 6.202
R621 VDD.n155 VDD.n154 6.202
R622 VDD.n216 VDD.n215 6.202
R623 VDD.n262 VDD.n261 6.202
R624 VDD.n323 VDD.n322 6.202
R625 VDD.n369 VDD.n368 6.202
R626 VDD.n708 VDD.n707 6.202
R627 VDD.n650 VDD.n649 6.202
R628 VDD.n601 VDD.n600 6.202
R629 VDD.n558 VDD.n557 6.202
R630 VDD.n500 VDD.n499 6.202
R631 VDD.n394 VDD.n393 6.202
R632 VDD.n93 VDD.n89 5.903
R633 VDD.n734 VDD.n730 5.903
R634 VDD.n676 VDD.n672 5.903
R635 VDD.n526 VDD.n522 5.903
R636 VDD.n468 VDD.n464 5.903
R637 VDD.n84 VDD.n83 4.576
R638 VDD.n192 VDD.n191 4.576
R639 VDD.n299 VDD.n298 4.576
R640 VDD.n737 VDD.n736 4.576
R641 VDD.n679 VDD.n678 4.576
R642 VDD.n529 VDD.n528 4.576
R643 VDD.n471 VDD.n470 4.576
R644 VDD.n204 VDD.n201 2.754
R645 VDD.n311 VDD.n308 2.754
R646 VDD.n178 VDD.n177 2.361
R647 VDD.n285 VDD.n282 2.361
R648 VDD.n28 VDD.n24 1.967
R649 VDD.n38 VDD.n37 1.967
R650 VDD.n133 VDD.n129 1.967
R651 VDD.n143 VDD.n139 1.967
R652 VDD.n240 VDD.n236 1.967
R653 VDD.n250 VDD.n249 1.967
R654 VDD.n347 VDD.n343 1.967
R655 VDD.n357 VDD.n353 1.967
R656 VDD.n635 VDD.n631 1.967
R657 VDD.n625 VDD.n624 1.967
R658 VDD.n589 VDD.n585 1.967
R659 VDD.n579 VDD.n575 1.967
R660 VDD.n426 VDD.n422 1.967
R661 VDD.n416 VDD.n415 1.967
R662 VDD.n14 VDD.n7 1.329
R663 VDD.n14 VDD.n8 1.329
R664 VDD.n14 VDD.n12 1.329
R665 VDD.n14 VDD.n13 1.329
R666 VDD.n15 VDD.n14 0.696
R667 VDD.n14 VDD.n4 0.696
R668 VDD.n61 VDD.n60 0.365
R669 VDD.n61 VDD.n56 0.365
R670 VDD.n61 VDD.n51 0.365
R671 VDD.n62 VDD.n61 0.365
R672 VDD.n119 VDD.n118 0.365
R673 VDD.n119 VDD.n114 0.365
R674 VDD.n120 VDD.n119 0.365
R675 VDD.n165 VDD.n164 0.365
R676 VDD.n165 VDD.n160 0.365
R677 VDD.n166 VDD.n165 0.365
R678 VDD.n226 VDD.n225 0.365
R679 VDD.n226 VDD.n221 0.365
R680 VDD.n227 VDD.n226 0.365
R681 VDD.n272 VDD.n271 0.365
R682 VDD.n272 VDD.n267 0.365
R683 VDD.n273 VDD.n272 0.365
R684 VDD.n333 VDD.n332 0.365
R685 VDD.n333 VDD.n328 0.365
R686 VDD.n334 VDD.n333 0.365
R687 VDD.n379 VDD.n378 0.365
R688 VDD.n379 VDD.n374 0.365
R689 VDD.n380 VDD.n379 0.365
R690 VDD.n718 VDD.n717 0.365
R691 VDD.n718 VDD.n713 0.365
R692 VDD.n719 VDD.n718 0.365
R693 VDD.n660 VDD.n659 0.365
R694 VDD.n660 VDD.n655 0.365
R695 VDD.n661 VDD.n660 0.365
R696 VDD.n611 VDD.n610 0.365
R697 VDD.n611 VDD.n606 0.365
R698 VDD.n612 VDD.n611 0.365
R699 VDD.n568 VDD.n567 0.365
R700 VDD.n568 VDD.n563 0.365
R701 VDD.n569 VDD.n568 0.365
R702 VDD.n510 VDD.n509 0.365
R703 VDD.n510 VDD.n505 0.365
R704 VDD.n511 VDD.n510 0.365
R705 VDD.n404 VDD.n403 0.365
R706 VDD.n404 VDD.n399 0.365
R707 VDD.n405 VDD.n404 0.365
R708 VDD.n452 VDD.n451 0.365
R709 VDD.n452 VDD.n446 0.365
R710 VDD.n452 VDD.n441 0.365
R711 VDD.n453 VDD.n452 0.365
R712 VDD.n70 VDD.n43 0.29
R713 VDD.n128 VDD.n102 0.29
R714 VDD.n174 VDD.n148 0.29
R715 VDD.n235 VDD.n209 0.29
R716 VDD.n281 VDD.n255 0.29
R717 VDD.n342 VDD.n316 0.29
R718 VDD.n388 VDD.n362 0.29
R719 VDD.n724 VDD.n698 0.29
R720 VDD.n666 VDD.n640 0.29
R721 VDD.n620 VDD.n594 0.29
R722 VDD.n574 VDD.n548 0.29
R723 VDD.n516 VDD.n490 0.29
R724 VDD.n458 VDD.n431 0.29
R725 VDD.n411 VDD 0.207
R726 VDD.n87 VDD.n82 0.181
R727 VDD.n195 VDD.n190 0.181
R728 VDD.n302 VDD.n297 0.181
R729 VDD.n744 VDD.n740 0.181
R730 VDD.n686 VDD.n682 0.181
R731 VDD.n536 VDD.n532 0.181
R732 VDD.n478 VDD.n474 0.181
R733 VDD.n33 VDD.n29 0.157
R734 VDD.n39 VDD.n33 0.157
R735 VDD.n138 VDD.n134 0.157
R736 VDD.n144 VDD.n138 0.157
R737 VDD.n245 VDD.n241 0.157
R738 VDD.n251 VDD.n245 0.157
R739 VDD.n352 VDD.n348 0.157
R740 VDD.n358 VDD.n352 0.157
R741 VDD.n636 VDD.n630 0.157
R742 VDD.n630 VDD.n626 0.157
R743 VDD.n590 VDD.n584 0.157
R744 VDD.n584 VDD.n580 0.157
R745 VDD.n427 VDD.n421 0.157
R746 VDD.n421 VDD.n417 0.157
R747 VDD.n43 VDD.n39 0.145
R748 VDD.n74 VDD.n70 0.145
R749 VDD.n78 VDD.n74 0.145
R750 VDD.n82 VDD.n78 0.145
R751 VDD.n94 VDD.n87 0.145
R752 VDD.n98 VDD.n94 0.145
R753 VDD.n102 VDD.n98 0.145
R754 VDD.n134 VDD.n128 0.145
R755 VDD.n148 VDD.n144 0.145
R756 VDD.n179 VDD.n174 0.145
R757 VDD.n184 VDD.n179 0.145
R758 VDD.n190 VDD.n184 0.145
R759 VDD.n200 VDD.n195 0.145
R760 VDD.n205 VDD.n200 0.145
R761 VDD.n209 VDD.n205 0.145
R762 VDD.n241 VDD.n235 0.145
R763 VDD.n255 VDD.n251 0.145
R764 VDD.n286 VDD.n281 0.145
R765 VDD.n291 VDD.n286 0.145
R766 VDD.n297 VDD.n291 0.145
R767 VDD.n307 VDD.n302 0.145
R768 VDD.n312 VDD.n307 0.145
R769 VDD.n316 VDD.n312 0.145
R770 VDD.n348 VDD.n342 0.145
R771 VDD.n362 VDD.n358 0.145
R772 VDD.n752 VDD.n748 0.145
R773 VDD.n748 VDD.n744 0.145
R774 VDD.n740 VDD.n735 0.145
R775 VDD.n735 VDD.n728 0.145
R776 VDD.n728 VDD.n724 0.145
R777 VDD.n698 VDD.n694 0.145
R778 VDD.n694 VDD.n690 0.145
R779 VDD.n690 VDD.n686 0.145
R780 VDD.n682 VDD.n677 0.145
R781 VDD.n677 VDD.n670 0.145
R782 VDD.n670 VDD.n666 0.145
R783 VDD.n640 VDD.n636 0.145
R784 VDD.n626 VDD.n620 0.145
R785 VDD.n594 VDD.n590 0.145
R786 VDD.n580 VDD.n574 0.145
R787 VDD.n548 VDD.n544 0.145
R788 VDD.n544 VDD.n540 0.145
R789 VDD.n540 VDD.n536 0.145
R790 VDD.n532 VDD.n527 0.145
R791 VDD.n527 VDD.n520 0.145
R792 VDD.n520 VDD.n516 0.145
R793 VDD.n490 VDD.n486 0.145
R794 VDD.n486 VDD.n482 0.145
R795 VDD.n482 VDD.n478 0.145
R796 VDD.n474 VDD.n469 0.145
R797 VDD.n469 VDD.n462 0.145
R798 VDD.n462 VDD.n458 0.145
R799 VDD.n431 VDD.n427 0.145
R800 VDD.n417 VDD.n411 0.145
R801 VDD VDD.n388 0.078
R802 VDD VDD.n752 0.066
R803 a_5767_1050.n0 a_5767_1050.t7 512.525
R804 a_5767_1050.n0 a_5767_1050.t5 371.139
R805 a_5767_1050.n1 a_5767_1050.t6 210.434
R806 a_5767_1050.n6 a_5767_1050.n5 184.039
R807 a_5767_1050.n8 a_5767_1050.n6 179.052
R808 a_5767_1050.n1 a_5767_1050.n0 173.2
R809 a_5767_1050.n6 a_5767_1050.n1 153.043
R810 a_5767_1050.n8 a_5767_1050.n7 76.002
R811 a_5767_1050.n5 a_5767_1050.n4 30
R812 a_5767_1050.n3 a_5767_1050.n2 24.383
R813 a_5767_1050.n5 a_5767_1050.n3 23.684
R814 a_5767_1050.n7 a_5767_1050.t0 14.282
R815 a_5767_1050.n7 a_5767_1050.t1 14.282
R816 a_5767_1050.n9 a_5767_1050.t3 14.282
R817 a_5767_1050.t4 a_5767_1050.n9 14.282
R818 a_5767_1050.n9 a_5767_1050.n8 12.848
R819 CIN.n2 CIN.t2 512.525
R820 CIN.n0 CIN.t1 480.392
R821 CIN.n5 CIN.t0 480.392
R822 CIN.n0 CIN.t5 403.272
R823 CIN.n5 CIN.t4 403.272
R824 CIN.n3 CIN.t8 372.349
R825 CIN.n2 CIN.t7 371.139
R826 CIN.n1 CIN.t6 336.586
R827 CIN.n3 CIN.t3 157.328
R828 CIN.n4 CIN.n3 132.764
R829 CIN.n6 CIN.n5 124.375
R830 CIN.n4 CIN.n2 93.541
R831 CIN.n6 CIN.n4 76
R832 CIN.n7 CIN.n1 76
R833 CIN.n1 CIN.n0 45.341
R834 CIN CIN.n6 1.269
R835 CIN.n7 CIN 0.046
R836 a_3461_1051.t2 a_3461_1051.n0 101.66
R837 a_3461_1051.n0 a_3461_1051.t0 101.659
R838 a_3461_1051.n0 a_3461_1051.t1 14.294
R839 a_3461_1051.n0 a_3461_1051.t3 14.282
R840 a_6401_209.n0 a_6401_209.t5 470.752
R841 a_6401_209.n0 a_6401_209.t3 384.527
R842 a_6401_209.n1 a_6401_209.t4 214.619
R843 a_6401_209.n7 a_6401_209.n6 184.006
R844 a_6401_209.n6 a_6401_209.n5 179.015
R845 a_6401_209.n6 a_6401_209.n1 153.859
R846 a_6401_209.n1 a_6401_209.n0 136.726
R847 a_6401_209.n5 a_6401_209.n4 30
R848 a_6401_209.n3 a_6401_209.n2 24.383
R849 a_6401_209.n5 a_6401_209.n3 23.684
R850 a_6401_209.n7 a_6401_209.t0 14.282
R851 a_6401_209.t1 a_6401_209.n7 14.282
R852 a_6791_1051.t0 a_6791_1051.n0 101.66
R853 a_6791_1051.n0 a_6791_1051.t3 101.659
R854 a_6791_1051.n0 a_6791_1051.t2 14.294
R855 a_6791_1051.n0 a_6791_1051.t1 14.282
R856 a_6858_209.n0 a_6858_209.t6 512.525
R857 a_6858_209.n0 a_6858_209.t5 371.139
R858 a_6858_209.n1 a_6858_209.t4 210.434
R859 a_6858_209.n11 a_6858_209.n10 191.888
R860 a_6858_209.n1 a_6858_209.n0 173.2
R861 a_6858_209.n10 a_6858_209.n1 153.043
R862 a_6858_209.n10 a_6858_209.n9 135.634
R863 a_6858_209.n9 a_6858_209.n8 118.016
R864 a_6858_209.n4 a_6858_209.n2 80.526
R865 a_6858_209.n9 a_6858_209.n4 48.405
R866 a_6858_209.n8 a_6858_209.n7 30
R867 a_6858_209.n4 a_6858_209.n3 30
R868 a_6858_209.n6 a_6858_209.n5 24.383
R869 a_6858_209.n8 a_6858_209.n6 23.684
R870 a_6858_209.n11 a_6858_209.t1 14.282
R871 a_6858_209.t2 a_6858_209.n11 14.282
R872 GND.n32 GND.n30 219.745
R873 GND.n276 GND.n275 219.745
R874 GND.n309 GND.n307 219.745
R875 GND.n339 GND.n337 219.745
R876 GND.n369 GND.n367 219.745
R877 GND.n402 GND.n400 219.745
R878 GND.n432 GND.n430 219.745
R879 GND.n237 GND.n235 219.745
R880 GND.n205 GND.n203 219.745
R881 GND.n172 GND.n170 219.745
R882 GND.n139 GND.n137 219.745
R883 GND.n109 GND.n107 219.745
R884 GND.n76 GND.n75 219.745
R885 GND.n32 GND.n31 85.529
R886 GND.n276 GND.n274 85.529
R887 GND.n309 GND.n308 85.529
R888 GND.n339 GND.n338 85.529
R889 GND.n369 GND.n368 85.529
R890 GND.n402 GND.n401 85.529
R891 GND.n432 GND.n431 85.529
R892 GND.n237 GND.n236 85.529
R893 GND.n205 GND.n204 85.529
R894 GND.n172 GND.n171 85.529
R895 GND.n139 GND.n138 85.529
R896 GND.n109 GND.n108 85.529
R897 GND.n76 GND.n74 85.529
R898 GND.n127 GND.n126 84.842
R899 GND.n440 GND.n439 84.842
R900 GND.n410 GND.n409 84.842
R901 GND.n317 GND.n316 84.842
R902 GND.n9 GND.n1 76.145
R903 GND.n244 GND.n243 76
R904 GND.n9 GND.n8 76
R905 GND.n17 GND.n16 76
R906 GND.n26 GND.n25 76
R907 GND.n29 GND.n28 76
R908 GND.n36 GND.n35 76
R909 GND.n43 GND.n42 76
R910 GND.n49 GND.n48 76
R911 GND.n52 GND.n51 76
R912 GND.n58 GND.n57 76
R913 GND.n63 GND.n62 76
R914 GND.n70 GND.n69 76
R915 GND.n73 GND.n72 76
R916 GND.n80 GND.n79 76
R917 GND.n88 GND.n87 76
R918 GND.n96 GND.n95 76
R919 GND.n103 GND.n102 76
R920 GND.n106 GND.n105 76
R921 GND.n113 GND.n112 76
R922 GND.n116 GND.n115 76
R923 GND.n119 GND.n118 76
R924 GND.n122 GND.n121 76
R925 GND.n125 GND.n124 76
R926 GND.n130 GND.n129 76
R927 GND.n133 GND.n132 76
R928 GND.n136 GND.n135 76
R929 GND.n143 GND.n142 76
R930 GND.n151 GND.n150 76
R931 GND.n159 GND.n158 76
R932 GND.n166 GND.n165 76
R933 GND.n169 GND.n168 76
R934 GND.n176 GND.n175 76
R935 GND.n179 GND.n178 76
R936 GND.n182 GND.n181 76
R937 GND.n185 GND.n184 76
R938 GND.n188 GND.n187 76
R939 GND.n196 GND.n195 76
R940 GND.n199 GND.n198 76
R941 GND.n202 GND.n201 76
R942 GND.n209 GND.n208 76
R943 GND.n216 GND.n215 76
R944 GND.n224 GND.n223 76
R945 GND.n231 GND.n230 76
R946 GND.n234 GND.n233 76
R947 GND.n241 GND.n240 76
R948 GND.n455 GND.n454 76
R949 GND.n452 GND.n451 76
R950 GND.n449 GND.n448 76
R951 GND.n446 GND.n445 76
R952 GND.n443 GND.n442 76
R953 GND.n438 GND.n437 76
R954 GND.n435 GND.n434 76
R955 GND.n428 GND.n427 76
R956 GND.n425 GND.n424 76
R957 GND.n422 GND.n421 76
R958 GND.n419 GND.n418 76
R959 GND.n416 GND.n415 76
R960 GND.n413 GND.n412 76
R961 GND.n408 GND.n407 76
R962 GND.n405 GND.n404 76
R963 GND.n398 GND.n397 76
R964 GND.n395 GND.n394 76
R965 GND.n387 GND.n386 76
R966 GND.n379 GND.n378 76
R967 GND.n372 GND.n371 76
R968 GND.n365 GND.n364 76
R969 GND.n362 GND.n361 76
R970 GND.n355 GND.n354 76
R971 GND.n349 GND.n348 76
R972 GND.n342 GND.n341 76
R973 GND.n335 GND.n334 76
R974 GND.n332 GND.n331 76
R975 GND.n329 GND.n328 76
R976 GND.n326 GND.n325 76
R977 GND.n323 GND.n322 76
R978 GND.n320 GND.n319 76
R979 GND.n315 GND.n314 76
R980 GND.n312 GND.n311 76
R981 GND.n305 GND.n304 76
R982 GND.n302 GND.n301 76
R983 GND.n299 GND.n298 76
R984 GND.n296 GND.n295 76
R985 GND.n293 GND.n292 76
R986 GND.n290 GND.n289 76
R987 GND.n282 GND.n281 76
R988 GND.n279 GND.n278 76
R989 GND.n272 GND.n271 76
R990 GND.n269 GND.n268 76
R991 GND.n261 GND.n260 76
R992 GND.n253 GND.n252 76
R993 GND.n193 GND.n192 63.835
R994 GND.n287 GND.n286 63.835
R995 GND.n211 GND.t6 39.413
R996 GND.n22 GND.t7 39.412
R997 GND.n249 GND.t11 39.412
R998 GND.n5 GND.n4 35.01
R999 GND.n84 GND.n83 35.01
R1000 GND.n147 GND.n146 35.01
R1001 GND.n391 GND.n390 35.01
R1002 GND.n265 GND.n264 35.01
R1003 GND.n82 GND.n81 29.127
R1004 GND.n145 GND.n144 29.127
R1005 GND.n389 GND.n388 29.127
R1006 GND.n192 GND.n191 28.421
R1007 GND.n286 GND.n285 28.421
R1008 GND.n192 GND.n190 25.263
R1009 GND.n286 GND.n284 25.263
R1010 GND.n190 GND.n189 24.383
R1011 GND.n284 GND.n283 24.383
R1012 GND.n91 GND.t10 20.794
R1013 GND.n154 GND.t0 20.794
R1014 GND.n382 GND.t14 20.794
R1015 GND.n6 GND.n5 19.735
R1016 GND.n14 GND.n13 19.735
R1017 GND.n24 GND.n23 19.735
R1018 GND.n60 GND.n59 19.735
R1019 GND.n55 GND.n54 19.735
R1020 GND.n47 GND.n46 19.735
R1021 GND.n40 GND.n39 19.735
R1022 GND.n68 GND.n67 19.735
R1023 GND.n85 GND.n84 19.735
R1024 GND.n93 GND.n92 19.735
R1025 GND.n101 GND.n100 19.735
R1026 GND.n148 GND.n147 19.735
R1027 GND.n156 GND.n155 19.735
R1028 GND.n164 GND.n163 19.735
R1029 GND.n213 GND.n212 19.735
R1030 GND.n222 GND.n221 19.735
R1031 GND.n229 GND.n228 19.735
R1032 GND.n392 GND.n391 19.735
R1033 GND.n384 GND.n383 19.735
R1034 GND.n377 GND.n376 19.735
R1035 GND.n359 GND.n358 19.735
R1036 GND.n353 GND.n352 19.735
R1037 GND.n347 GND.n346 19.735
R1038 GND.n266 GND.n265 19.735
R1039 GND.n258 GND.n257 19.735
R1040 GND.n251 GND.n250 19.735
R1041 GND.n46 GND.t8 19.724
R1042 GND.n59 GND.t4 19.724
R1043 GND.n5 GND.n3 19.017
R1044 GND.n84 GND.n82 19.017
R1045 GND.n147 GND.n145 19.017
R1046 GND.n391 GND.n389 19.017
R1047 GND.n265 GND.n263 19.017
R1048 GND.n351 GND.t1 18.552
R1049 GND.n227 GND.n226 18.345
R1050 GND.n22 GND.n21 17.185
R1051 GND.n249 GND.n248 17.185
R1052 GND.n211 GND.n210 17.185
R1053 GND.n35 GND.n33 14.167
R1054 GND.n79 GND.n77 14.167
R1055 GND.n112 GND.n110 14.167
R1056 GND.n142 GND.n140 14.167
R1057 GND.n175 GND.n173 14.167
R1058 GND.n208 GND.n206 14.167
R1059 GND.n240 GND.n238 14.167
R1060 GND.n434 GND.n433 14.167
R1061 GND.n404 GND.n403 14.167
R1062 GND.n371 GND.n370 14.167
R1063 GND.n341 GND.n340 14.167
R1064 GND.n311 GND.n310 14.167
R1065 GND.n278 GND.n277 14.167
R1066 GND.n252 GND.n245 13.653
R1067 GND.n260 GND.n259 13.653
R1068 GND.n268 GND.n267 13.653
R1069 GND.n271 GND.n270 13.653
R1070 GND.n278 GND.n273 13.653
R1071 GND.n281 GND.n280 13.653
R1072 GND.n289 GND.n288 13.653
R1073 GND.n292 GND.n291 13.653
R1074 GND.n295 GND.n294 13.653
R1075 GND.n298 GND.n297 13.653
R1076 GND.n301 GND.n300 13.653
R1077 GND.n304 GND.n303 13.653
R1078 GND.n311 GND.n306 13.653
R1079 GND.n314 GND.n313 13.653
R1080 GND.n319 GND.n318 13.653
R1081 GND.n322 GND.n321 13.653
R1082 GND.n325 GND.n324 13.653
R1083 GND.n328 GND.n327 13.653
R1084 GND.n331 GND.n330 13.653
R1085 GND.n334 GND.n333 13.653
R1086 GND.n341 GND.n336 13.653
R1087 GND.n348 GND.n343 13.653
R1088 GND.n354 GND.n350 13.653
R1089 GND.n361 GND.n360 13.653
R1090 GND.n364 GND.n363 13.653
R1091 GND.n371 GND.n366 13.653
R1092 GND.n378 GND.n373 13.653
R1093 GND.n386 GND.n385 13.653
R1094 GND.n394 GND.n393 13.653
R1095 GND.n397 GND.n396 13.653
R1096 GND.n404 GND.n399 13.653
R1097 GND.n407 GND.n406 13.653
R1098 GND.n412 GND.n411 13.653
R1099 GND.n415 GND.n414 13.653
R1100 GND.n418 GND.n417 13.653
R1101 GND.n421 GND.n420 13.653
R1102 GND.n424 GND.n423 13.653
R1103 GND.n427 GND.n426 13.653
R1104 GND.n434 GND.n429 13.653
R1105 GND.n437 GND.n436 13.653
R1106 GND.n442 GND.n441 13.653
R1107 GND.n445 GND.n444 13.653
R1108 GND.n448 GND.n447 13.653
R1109 GND.n451 GND.n450 13.653
R1110 GND.n454 GND.n453 13.653
R1111 GND.n240 GND.n239 13.653
R1112 GND.n233 GND.n232 13.653
R1113 GND.n230 GND.n225 13.653
R1114 GND.n223 GND.n217 13.653
R1115 GND.n215 GND.n214 13.653
R1116 GND.n208 GND.n207 13.653
R1117 GND.n201 GND.n200 13.653
R1118 GND.n198 GND.n197 13.653
R1119 GND.n195 GND.n194 13.653
R1120 GND.n187 GND.n186 13.653
R1121 GND.n184 GND.n183 13.653
R1122 GND.n181 GND.n180 13.653
R1123 GND.n178 GND.n177 13.653
R1124 GND.n175 GND.n174 13.653
R1125 GND.n168 GND.n167 13.653
R1126 GND.n165 GND.n160 13.653
R1127 GND.n158 GND.n157 13.653
R1128 GND.n150 GND.n149 13.653
R1129 GND.n142 GND.n141 13.653
R1130 GND.n135 GND.n134 13.653
R1131 GND.n132 GND.n131 13.653
R1132 GND.n129 GND.n128 13.653
R1133 GND.n124 GND.n123 13.653
R1134 GND.n121 GND.n120 13.653
R1135 GND.n118 GND.n117 13.653
R1136 GND.n115 GND.n114 13.653
R1137 GND.n112 GND.n111 13.653
R1138 GND.n105 GND.n104 13.653
R1139 GND.n102 GND.n97 13.653
R1140 GND.n95 GND.n94 13.653
R1141 GND.n87 GND.n86 13.653
R1142 GND.n79 GND.n78 13.653
R1143 GND.n72 GND.n71 13.653
R1144 GND.n69 GND.n64 13.653
R1145 GND.n62 GND.n61 13.653
R1146 GND.n57 GND.n56 13.653
R1147 GND.n51 GND.n50 13.653
R1148 GND.n48 GND.n44 13.653
R1149 GND.n42 GND.n41 13.653
R1150 GND.n35 GND.n34 13.653
R1151 GND.n28 GND.n27 13.653
R1152 GND.n25 GND.n18 13.653
R1153 GND.n16 GND.n15 13.653
R1154 GND.n8 GND.n7 13.653
R1155 GND.n346 GND.n345 13.608
R1156 GND.n67 GND.n66 12.837
R1157 GND.n100 GND.n99 12.837
R1158 GND.n163 GND.n162 12.837
R1159 GND.n376 GND.n375 12.837
R1160 GND.n39 GND.n38 11.605
R1161 GND.n358 GND.n357 10.853
R1162 GND.n357 GND.n356 10.417
R1163 GND.n38 GND.n37 9.809
R1164 GND.n57 GND.n55 8.854
R1165 GND.n345 GND.n344 7.858
R1166 GND.n66 GND.n65 7.566
R1167 GND.n99 GND.n98 7.566
R1168 GND.n162 GND.n161 7.566
R1169 GND.n375 GND.n374 7.566
R1170 GND.n3 GND.n2 7.5
R1171 GND.n12 GND.n11 7.5
R1172 GND.n220 GND.n219 7.5
R1173 GND.n263 GND.n262 7.5
R1174 GND.n256 GND.n255 7.5
R1175 GND.n33 GND.n32 7.312
R1176 GND.n277 GND.n276 7.312
R1177 GND.n310 GND.n309 7.312
R1178 GND.n340 GND.n339 7.312
R1179 GND.n370 GND.n369 7.312
R1180 GND.n403 GND.n402 7.312
R1181 GND.n433 GND.n432 7.312
R1182 GND.n238 GND.n237 7.312
R1183 GND.n206 GND.n205 7.312
R1184 GND.n173 GND.n172 7.312
R1185 GND.n140 GND.n139 7.312
R1186 GND.n110 GND.n109 7.312
R1187 GND.n77 GND.n76 7.312
R1188 GND.t8 GND.n45 7.04
R1189 GND.n228 GND.n227 6.358
R1190 GND.n212 GND.n211 6.139
R1191 GND.n23 GND.n22 6.139
R1192 GND.n250 GND.n249 6.139
R1193 GND.n54 GND.n53 5.774
R1194 GND.n20 GND.n19 4.551
R1195 GND.n90 GND.n89 4.551
R1196 GND.n153 GND.n152 4.551
R1197 GND.n381 GND.n380 4.551
R1198 GND.n247 GND.n246 4.551
R1199 GND.n8 GND.n6 3.935
R1200 GND.n48 GND.n47 3.935
R1201 GND.n62 GND.n60 3.935
R1202 GND.n87 GND.n85 3.935
R1203 GND.n129 GND.n127 3.935
R1204 GND.n150 GND.n148 3.935
R1205 GND.n195 GND.n193 3.935
R1206 GND.n230 GND.n229 3.935
R1207 GND.n442 GND.n440 3.935
R1208 GND.n412 GND.n410 3.935
R1209 GND.n394 GND.n392 3.935
R1210 GND.n348 GND.n347 3.935
R1211 GND.n319 GND.n317 3.935
R1212 GND.n289 GND.n287 3.935
R1213 GND.n268 GND.n266 3.935
R1214 GND.n25 GND.n24 3.541
R1215 GND.n102 GND.n101 3.541
R1216 GND.n165 GND.n164 3.541
R1217 GND.n215 GND.n213 3.541
R1218 GND.n378 GND.n377 3.541
R1219 GND.n361 GND.n359 3.541
R1220 GND.n252 GND.n251 3.541
R1221 GND.t7 GND.n20 2.238
R1222 GND.t10 GND.n90 2.238
R1223 GND.t0 GND.n153 2.238
R1224 GND.t14 GND.n381 2.238
R1225 GND.t11 GND.n247 2.238
R1226 GND.n11 GND.n10 1.935
R1227 GND.n219 GND.n218 1.935
R1228 GND.n255 GND.n254 1.935
R1229 GND.n42 GND.n40 0.983
R1230 GND.n69 GND.n68 0.983
R1231 GND.n1 GND.n0 0.596
R1232 GND.n243 GND.n242 0.596
R1233 GND.n13 GND.n12 0.358
R1234 GND.n92 GND.n91 0.358
R1235 GND.n155 GND.n154 0.358
R1236 GND.n221 GND.n220 0.358
R1237 GND.n383 GND.n382 0.358
R1238 GND.n352 GND.n351 0.358
R1239 GND.n257 GND.n256 0.358
R1240 GND.n36 GND.n29 0.29
R1241 GND.n80 GND.n73 0.29
R1242 GND.n113 GND.n106 0.29
R1243 GND.n143 GND.n136 0.29
R1244 GND.n176 GND.n169 0.29
R1245 GND.n209 GND.n202 0.29
R1246 GND.n241 GND.n234 0.29
R1247 GND.n435 GND.n428 0.29
R1248 GND.n405 GND.n398 0.29
R1249 GND.n372 GND.n365 0.29
R1250 GND.n342 GND.n335 0.29
R1251 GND.n312 GND.n305 0.29
R1252 GND.n279 GND.n272 0.29
R1253 GND.n244 GND 0.207
R1254 GND.n16 GND.n14 0.196
R1255 GND.n95 GND.n93 0.196
R1256 GND.n158 GND.n156 0.196
R1257 GND.n223 GND.n222 0.196
R1258 GND.n386 GND.n384 0.196
R1259 GND.n354 GND.n353 0.196
R1260 GND.n260 GND.n258 0.196
R1261 GND.n58 GND.n52 0.181
R1262 GND.n125 GND.n122 0.181
R1263 GND.n188 GND.n185 0.181
R1264 GND.n449 GND.n446 0.181
R1265 GND.n419 GND.n416 0.181
R1266 GND.n326 GND.n323 0.181
R1267 GND.n296 GND.n293 0.181
R1268 GND.n17 GND.n9 0.157
R1269 GND.n26 GND.n17 0.157
R1270 GND.n96 GND.n88 0.157
R1271 GND.n103 GND.n96 0.157
R1272 GND.n159 GND.n151 0.157
R1273 GND.n166 GND.n159 0.157
R1274 GND.n224 GND.n216 0.157
R1275 GND.n231 GND.n224 0.157
R1276 GND.n395 GND.n387 0.157
R1277 GND.n387 GND.n379 0.157
R1278 GND.n362 GND.n355 0.157
R1279 GND.n355 GND.n349 0.157
R1280 GND.n269 GND.n261 0.157
R1281 GND.n261 GND.n253 0.157
R1282 GND.n29 GND.n26 0.145
R1283 GND.n43 GND.n36 0.145
R1284 GND.n49 GND.n43 0.145
R1285 GND.n52 GND.n49 0.145
R1286 GND.n63 GND.n58 0.145
R1287 GND.n70 GND.n63 0.145
R1288 GND.n73 GND.n70 0.145
R1289 GND.n88 GND.n80 0.145
R1290 GND.n106 GND.n103 0.145
R1291 GND.n116 GND.n113 0.145
R1292 GND.n119 GND.n116 0.145
R1293 GND.n122 GND.n119 0.145
R1294 GND.n130 GND.n125 0.145
R1295 GND.n133 GND.n130 0.145
R1296 GND.n136 GND.n133 0.145
R1297 GND.n151 GND.n143 0.145
R1298 GND.n169 GND.n166 0.145
R1299 GND.n179 GND.n176 0.145
R1300 GND.n182 GND.n179 0.145
R1301 GND.n185 GND.n182 0.145
R1302 GND.n196 GND.n188 0.145
R1303 GND.n199 GND.n196 0.145
R1304 GND.n202 GND.n199 0.145
R1305 GND.n216 GND.n209 0.145
R1306 GND.n234 GND.n231 0.145
R1307 GND.n455 GND.n452 0.145
R1308 GND.n452 GND.n449 0.145
R1309 GND.n446 GND.n443 0.145
R1310 GND.n443 GND.n438 0.145
R1311 GND.n438 GND.n435 0.145
R1312 GND.n428 GND.n425 0.145
R1313 GND.n425 GND.n422 0.145
R1314 GND.n422 GND.n419 0.145
R1315 GND.n416 GND.n413 0.145
R1316 GND.n413 GND.n408 0.145
R1317 GND.n408 GND.n405 0.145
R1318 GND.n398 GND.n395 0.145
R1319 GND.n379 GND.n372 0.145
R1320 GND.n365 GND.n362 0.145
R1321 GND.n349 GND.n342 0.145
R1322 GND.n335 GND.n332 0.145
R1323 GND.n332 GND.n329 0.145
R1324 GND.n329 GND.n326 0.145
R1325 GND.n323 GND.n320 0.145
R1326 GND.n320 GND.n315 0.145
R1327 GND.n315 GND.n312 0.145
R1328 GND.n305 GND.n302 0.145
R1329 GND.n302 GND.n299 0.145
R1330 GND.n299 GND.n296 0.145
R1331 GND.n293 GND.n290 0.145
R1332 GND.n290 GND.n282 0.145
R1333 GND.n282 GND.n279 0.145
R1334 GND.n272 GND.n269 0.145
R1335 GND.n253 GND.n244 0.145
R1336 GND GND.n241 0.078
R1337 GND GND.n455 0.066
R1338 a_185_209.n0 a_185_209.t3 477.179
R1339 a_185_209.n0 a_185_209.t5 406.485
R1340 a_185_209.n1 a_185_209.t4 269.148
R1341 a_185_209.n3 a_185_209.n2 200.754
R1342 a_185_209.n4 a_185_209.n3 184.006
R1343 a_185_209.n3 a_185_209.n1 156.579
R1344 a_185_209.n1 a_185_209.n0 125.359
R1345 a_185_209.n4 a_185_209.t1 14.282
R1346 a_185_209.t2 a_185_209.n4 14.282
R1347 a_556_101.t0 a_556_101.n1 34.62
R1348 a_556_101.t0 a_556_101.n0 8.137
R1349 a_556_101.t0 a_556_101.n2 4.69
R1350 a_4657_1050.n1 a_4657_1050.t5 512.525
R1351 a_4657_1050.n1 a_4657_1050.t6 371.139
R1352 a_4657_1050.n2 a_4657_1050.t7 210.434
R1353 a_4657_1050.n4 a_4657_1050.n3 205.778
R1354 a_4657_1050.n5 a_4657_1050.n4 179.052
R1355 a_4657_1050.n2 a_4657_1050.n1 173.2
R1356 a_4657_1050.n4 a_4657_1050.n2 153.043
R1357 a_4657_1050.n6 a_4657_1050.n5 76.001
R1358 a_4657_1050.n0 a_4657_1050.t0 14.282
R1359 a_4657_1050.n0 a_4657_1050.t3 14.282
R1360 a_4657_1050.t2 a_4657_1050.n6 14.282
R1361 a_4657_1050.n6 a_4657_1050.t1 14.282
R1362 a_4657_1050.n5 a_4657_1050.n0 12.85
R1363 a_836_209.n1 a_836_209.t8 512.525
R1364 a_836_209.n2 a_836_209.t10 480.392
R1365 a_836_209.n5 a_836_209.t9 472.359
R1366 a_836_209.n2 a_836_209.t7 403.272
R1367 a_836_209.n5 a_836_209.t12 384.527
R1368 a_836_209.n1 a_836_209.t11 371.139
R1369 a_836_209.n3 a_836_209.t13 336.586
R1370 a_836_209.n18 a_836_209.n16 217.115
R1371 a_836_209.n6 a_836_209.n5 216.272
R1372 a_836_209.n14 a_836_209.n13 210.593
R1373 a_836_209.n14 a_836_209.n9 165.336
R1374 a_836_209.n16 a_836_209.n0 165.336
R1375 a_836_209.n7 a_836_209.n6 160.932
R1376 a_836_209.n4 a_836_209.n3 153.859
R1377 a_836_209.n6 a_836_209.t6 141.114
R1378 a_836_209.n7 a_836_209.t14 136.929
R1379 a_836_209.n8 a_836_209.n7 106.211
R1380 a_836_209.n4 a_836_209.n1 93.541
R1381 a_836_209.n15 a_836_209.n8 78.675
R1382 a_836_209.n16 a_836_209.n15 78.403
R1383 a_836_209.n15 a_836_209.n14 76
R1384 a_836_209.n8 a_836_209.n4 53.105
R1385 a_836_209.n3 a_836_209.n2 45.7
R1386 a_836_209.n13 a_836_209.n12 30
R1387 a_836_209.n11 a_836_209.n10 24.383
R1388 a_836_209.n13 a_836_209.n11 23.684
R1389 a_836_209.n18 a_836_209.n17 15.218
R1390 a_836_209.n9 a_836_209.t4 14.282
R1391 a_836_209.n9 a_836_209.t3 14.282
R1392 a_836_209.n0 a_836_209.t0 14.282
R1393 a_836_209.n0 a_836_209.t5 14.282
R1394 a_836_209.n19 a_836_209.n18 12.014
R1395 a_4552_101.n12 a_4552_101.n11 26.811
R1396 a_4552_101.n6 a_4552_101.n5 24.977
R1397 a_4552_101.n2 a_4552_101.n1 24.877
R1398 a_4552_101.t0 a_4552_101.n2 12.677
R1399 a_4552_101.t0 a_4552_101.n3 11.595
R1400 a_4552_101.t1 a_4552_101.n8 8.137
R1401 a_4552_101.t0 a_4552_101.n4 7.273
R1402 a_4552_101.t0 a_4552_101.n0 6.109
R1403 a_4552_101.t1 a_4552_101.n7 4.864
R1404 a_4552_101.t0 a_4552_101.n12 2.074
R1405 a_4552_101.n7 a_4552_101.n6 1.13
R1406 a_4552_101.n12 a_4552_101.t1 0.937
R1407 a_4552_101.t1 a_4552_101.n10 0.804
R1408 a_4552_101.n10 a_4552_101.n9 0.136
R1409 a_575_1051.n0 a_575_1051.t0 101.66
R1410 a_575_1051.n0 a_575_1051.t1 101.66
R1411 a_575_1051.n0 a_575_1051.t3 14.294
R1412 a_575_1051.t2 a_575_1051.n0 14.282
R1413 a_1241_1051.t2 a_1241_1051.n0 101.663
R1414 a_1241_1051.n0 a_1241_1051.t0 101.661
R1415 a_1241_1051.n0 a_1241_1051.t3 14.294
R1416 a_1241_1051.n0 a_1241_1051.t1 14.282
R1417 B.n2 B.t1 512.525
R1418 B.n6 B.t5 480.392
R1419 B.n0 B.t4 480.392
R1420 B.n6 B.t8 403.272
R1421 B.n0 B.t6 403.272
R1422 B.n4 B.t3 372.349
R1423 B.n2 B.t0 371.139
R1424 B.n1 B.t7 363.924
R1425 B.n4 B.t2 157.328
R1426 B.n5 B.n4 132.764
R1427 B.n7 B.n6 121.7
R1428 B.n3 B.n1 112.241
R1429 B.n7 B.n5 78.675
R1430 B.n3 B.n2 63.745
R1431 B.n5 B.n3 27.338
R1432 B.n1 B.n0 15.545
R1433 B.n7 B 0.046
R1434 a_807_990.n0 a_807_990.t4 477.179
R1435 a_807_990.n0 a_807_990.t3 406.485
R1436 a_807_990.n4 a_807_990.t5 384.505
R1437 a_807_990.n5 a_807_990.n0 228.016
R1438 a_807_990.n4 a_807_990.n3 167.985
R1439 a_807_990.n6 a_807_990.n5 130.9
R1440 a_807_990.n5 a_807_990.n4 79.658
R1441 a_807_990.n3 a_807_990.n2 22.578
R1442 a_807_990.t2 a_807_990.n6 14.282
R1443 a_807_990.n6 a_807_990.t1 14.282
R1444 a_807_990.n3 a_807_990.n1 8.58
R1445 a_5291_209.n0 a_5291_209.t3 486.819
R1446 a_5291_209.n0 a_5291_209.t5 384.527
R1447 a_5291_209.n1 a_5291_209.t4 223.948
R1448 a_5291_209.n4 a_5291_209.n3 210.559
R1449 a_5291_209.n3 a_5291_209.n2 174.201
R1450 a_5291_209.n1 a_5291_209.n0 159.653
R1451 a_5291_209.n3 a_5291_209.n1 157.396
R1452 a_5291_209.t2 a_5291_209.n4 14.282
R1453 a_5291_209.n4 a_5291_209.t1 14.282
R1454 a_2795_1051.n0 a_2795_1051.t0 101.66
R1455 a_2795_1051.n0 a_2795_1051.t3 101.66
R1456 a_2795_1051.n0 a_2795_1051.t1 14.294
R1457 a_2795_1051.t2 a_2795_1051.n0 14.282
R1458 a_2405_209.n0 a_2405_209.t5 477.179
R1459 a_2405_209.n0 a_2405_209.t3 406.485
R1460 a_2405_209.n1 a_2405_209.t4 269.148
R1461 a_2405_209.n3 a_2405_209.n2 200.754
R1462 a_2405_209.n4 a_2405_209.n3 184.006
R1463 a_2405_209.n3 a_2405_209.n1 156.579
R1464 a_2405_209.n1 a_2405_209.n0 125.359
R1465 a_2405_209.t2 a_2405_209.n4 14.282
R1466 a_2405_209.n4 a_2405_209.t1 14.282
R1467 a_1222_101.t0 a_1222_101.n1 34.62
R1468 a_1222_101.t0 a_1222_101.n0 8.137
R1469 a_1222_101.t0 a_1222_101.n2 4.69
R1470 a_3027_990.n0 a_3027_990.t4 477.179
R1471 a_3027_990.n0 a_3027_990.t5 406.485
R1472 a_3027_990.n4 a_3027_990.t3 384.505
R1473 a_3027_990.n5 a_3027_990.n0 228.016
R1474 a_3027_990.n4 a_3027_990.n3 167.985
R1475 a_3027_990.n6 a_3027_990.n5 130.9
R1476 a_3027_990.n5 a_3027_990.n4 79.658
R1477 a_3027_990.n3 a_3027_990.n2 22.578
R1478 a_3027_990.n6 a_3027_990.t1 14.282
R1479 a_3027_990.t2 a_3027_990.n6 14.282
R1480 a_3027_990.n3 a_3027_990.n1 8.58
R1481 a_3442_101.n5 a_3442_101.n4 24.877
R1482 a_3442_101.t0 a_3442_101.n5 12.677
R1483 a_3442_101.t0 a_3442_101.n3 11.595
R1484 a_3442_101.t0 a_3442_101.n6 8.137
R1485 a_3442_101.n2 a_3442_101.n0 4.031
R1486 a_3442_101.n2 a_3442_101.n1 3.644
R1487 a_3442_101.t0 a_3442_101.n2 1.093
R1488 a_5662_101.t0 a_5662_101.n1 34.62
R1489 a_5662_101.t0 a_5662_101.n0 8.137
R1490 a_5662_101.t0 a_5662_101.n2 4.69
R1491 COUT.n2 COUT.n1 200.754
R1492 COUT.n2 COUT.n0 184.007
R1493 COUT.n3 COUT.n2 76
R1494 COUT.n0 COUT.t1 14.282
R1495 COUT.n0 COUT.t2 14.282
R1496 COUT.n3 COUT 0.046
R1497 SUM.n2 SUM.n1 232.332
R1498 SUM.n8 SUM.n7 210.593
R1499 SUM.n2 SUM.n0 165.336
R1500 SUM.n8 SUM.n3 165.336
R1501 SUM SUM.n8 78.357
R1502 SUM.n9 SUM.n2 76
R1503 SUM.n7 SUM.n6 30
R1504 SUM.n5 SUM.n4 24.383
R1505 SUM.n7 SUM.n5 23.684
R1506 SUM.n0 SUM.t4 14.282
R1507 SUM.n0 SUM.t3 14.282
R1508 SUM.n3 SUM.t1 14.282
R1509 SUM.n3 SUM.t2 14.282
R1510 SUM.n9 SUM 0.046
R1511 a_2776_101.t0 a_2776_101.n1 34.62
R1512 a_2776_101.t0 a_2776_101.n0 8.137
R1513 a_2776_101.t0 a_2776_101.n2 4.69
C11 VDD GND 29.86fF
C12 a_2776_101.n0 GND 0.06fF
C13 a_2776_101.n1 GND 0.15fF
C14 a_2776_101.n2 GND 0.05fF
C15 SUM.n0 GND 1.21fF
C16 SUM.n1 GND 0.72fF
C17 SUM.n2 GND 0.86fF
C18 SUM.n3 GND 1.21fF
C19 SUM.n4 GND 0.07fF
C20 SUM.n5 GND 0.10fF
C21 SUM.n6 GND 0.06fF
C22 SUM.n7 GND 0.54fF
C23 SUM.n8 GND 0.82fF
C24 SUM.n9 GND 0.05fF
C25 a_5662_101.n0 GND 0.06fF
C26 a_5662_101.n1 GND 0.14fF
C27 a_5662_101.n2 GND 0.05fF
C28 a_3442_101.n0 GND 0.09fF
C29 a_3442_101.n1 GND 0.03fF
C30 a_3442_101.n2 GND 0.01fF
C31 a_3442_101.n3 GND 0.07fF
C32 a_3442_101.n4 GND 0.12fF
C33 a_3442_101.n5 GND 0.07fF
C34 a_3442_101.n6 GND 0.06fF
C35 a_3027_990.n0 GND 1.33fF
C36 a_3027_990.n1 GND 0.08fF
C37 a_3027_990.n2 GND 0.10fF
C38 a_3027_990.n3 GND 0.42fF
C39 a_3027_990.n4 GND 1.60fF
C40 a_3027_990.n5 GND 1.61fF
C41 a_3027_990.n6 GND 1.26fF
C42 a_1222_101.n0 GND 0.06fF
C43 a_1222_101.n1 GND 0.14fF
C44 a_1222_101.n2 GND 0.05fF
C45 a_2405_209.n0 GND 0.63fF
C46 a_2405_209.n1 GND 1.45fF
C47 a_2405_209.n2 GND 0.55fF
C48 a_2405_209.n3 GND 1.56fF
C49 a_2405_209.n4 GND 1.17fF
C50 a_2795_1051.n0 GND 0.52fF
C51 a_5291_209.n0 GND 0.46fF
C52 a_5291_209.t4 GND 0.52fF
C53 a_5291_209.n1 GND 1.11fF
C54 a_5291_209.n2 GND 0.35fF
C55 a_5291_209.n3 GND 1.20fF
C56 a_5291_209.n4 GND 0.86fF
C57 a_807_990.n0 GND 1.24fF
C58 a_807_990.n1 GND 0.07fF
C59 a_807_990.n2 GND 0.09fF
C60 a_807_990.n3 GND 0.39fF
C61 a_807_990.n4 GND 1.48fF
C62 a_807_990.n5 GND 1.50fF
C63 a_807_990.n6 GND 1.17fF
C64 a_1241_1051.n0 GND 0.52fF
C65 a_575_1051.n0 GND 0.52fF
C66 a_4552_101.n0 GND 0.03fF
C67 a_4552_101.n1 GND 0.12fF
C68 a_4552_101.n2 GND 0.07fF
C69 a_4552_101.n3 GND 0.07fF
C70 a_4552_101.n4 GND 0.00fF
C71 a_4552_101.n5 GND 0.05fF
C72 a_4552_101.n6 GND 0.06fF
C73 a_4552_101.n7 GND 0.02fF
C74 a_4552_101.n8 GND 0.06fF
C75 a_4552_101.n9 GND 0.09fF
C76 a_4552_101.n10 GND 0.21fF
C77 a_4552_101.t1 GND 0.28fF
C78 a_4552_101.n11 GND 0.11fF
C79 a_4552_101.n12 GND 0.00fF
C80 a_836_209.n0 GND 1.06fF
C81 a_836_209.n1 GND 0.44fF
C82 a_836_209.n2 GND 0.50fF
C83 a_836_209.n3 GND 1.02fF
C84 a_836_209.n4 GND 0.67fF
C85 a_836_209.n5 GND 0.73fF
C86 a_836_209.t6 GND 0.69fF
C87 a_836_209.n6 GND 2.20fF
C88 a_836_209.t14 GND 0.69fF
C89 a_836_209.n7 GND 2.01fF
C90 a_836_209.n8 GND 0.31fF
C91 a_836_209.n9 GND 1.06fF
C92 a_836_209.n10 GND 0.06fF
C93 a_836_209.n11 GND 0.09fF
C94 a_836_209.n12 GND 0.05fF
C95 a_836_209.n13 GND 0.48fF
C96 a_836_209.n14 GND 0.70fF
C97 a_836_209.n15 GND 1.90fF
C98 a_836_209.n16 GND 0.73fF
C99 a_836_209.n17 GND 0.13fF
C100 a_836_209.n18 GND 0.46fF
C101 a_836_209.n19 GND 0.07fF
C102 a_4657_1050.n0 GND 0.45fF
C103 a_4657_1050.n1 GND 0.32fF
C104 a_4657_1050.t7 GND 0.43fF
C105 a_4657_1050.n2 GND 0.49fF
C106 a_4657_1050.n3 GND 0.31fF
C107 a_4657_1050.n4 GND 0.51fF
C108 a_4657_1050.n5 GND 0.29fF
C109 a_4657_1050.n6 GND 0.53fF
C110 a_556_101.n0 GND 0.06fF
C111 a_556_101.n1 GND 0.14fF
C112 a_556_101.n2 GND 0.05fF
C113 a_185_209.n0 GND 0.55fF
C114 a_185_209.t4 GND 0.69fF
C115 a_185_209.n1 GND 1.27fF
C116 a_185_209.n2 GND 0.48fF
C117 a_185_209.n3 GND 1.36fF
C118 a_185_209.n4 GND 1.02fF
C119 a_6858_209.n0 GND 0.31fF
C120 a_6858_209.n1 GND 0.48fF
C121 a_6858_209.n2 GND 0.05fF
C122 a_6858_209.n3 GND 0.03fF
C123 a_6858_209.n4 GND 0.11fF
C124 a_6858_209.n5 GND 0.03fF
C125 a_6858_209.n6 GND 0.05fF
C126 a_6858_209.n7 GND 0.03fF
C127 a_6858_209.n8 GND 0.15fF
C128 a_6858_209.n9 GND 0.30fF
C129 a_6858_209.n10 GND 0.44fF
C130 a_6858_209.n11 GND 0.58fF
C131 a_6791_1051.n0 GND 0.55fF
C132 a_6401_209.n0 GND 0.38fF
C133 a_6401_209.t4 GND 0.52fF
C134 a_6401_209.n1 GND 0.63fF
C135 a_6401_209.n2 GND 0.04fF
C136 a_6401_209.n3 GND 0.06fF
C137 a_6401_209.n4 GND 0.04fF
C138 a_6401_209.n5 GND 0.26fF
C139 a_6401_209.n6 GND 0.70fF
C140 a_6401_209.n7 GND 0.78fF
C141 a_3461_1051.n0 GND 0.52fF
C142 a_5767_1050.n0 GND 0.33fF
C143 a_5767_1050.t6 GND 0.45fF
C144 a_5767_1050.n1 GND 0.51fF
C145 a_5767_1050.n2 GND 0.04fF
C146 a_5767_1050.n3 GND 0.05fF
C147 a_5767_1050.n4 GND 0.03fF
C148 a_5767_1050.n5 GND 0.24fF
C149 a_5767_1050.n6 GND 0.51fF
C150 a_5767_1050.n7 GND 0.56fF
C151 a_5767_1050.n8 GND 0.30fF
C152 a_5767_1050.n9 GND 0.47fF
C153 VDD.n0 GND 0.12fF
C154 VDD.n1 GND 0.02fF
C155 VDD.n2 GND 0.02fF
C156 VDD.n3 GND 0.04fF
C157 VDD.n4 GND 0.01fF
C158 VDD.n5 GND 0.02fF
C159 VDD.n6 GND 0.02fF
C160 VDD.n9 GND 0.02fF
C161 VDD.n10 GND 0.02fF
C162 VDD.n11 GND 0.02fF
C163 VDD.n14 GND 0.45fF
C164 VDD.n16 GND 0.03fF
C165 VDD.n17 GND 0.02fF
C166 VDD.n18 GND 0.02fF
C167 VDD.n19 GND 0.02fF
C168 VDD.n20 GND 0.03fF
C169 VDD.n21 GND 0.27fF
C170 VDD.n22 GND 0.02fF
C171 VDD.n23 GND 0.03fF
C172 VDD.n24 GND 0.06fF
C173 VDD.n25 GND 0.15fF
C174 VDD.n26 GND 0.20fF
C175 VDD.n27 GND 0.01fF
C176 VDD.n28 GND 0.01fF
C177 VDD.n29 GND 0.07fF
C178 VDD.n30 GND 0.16fF
C179 VDD.n31 GND 0.01fF
C180 VDD.n32 GND 0.02fF
C181 VDD.n33 GND 0.02fF
C182 VDD.n34 GND 0.15fF
C183 VDD.n35 GND 0.20fF
C184 VDD.n36 GND 0.01fF
C185 VDD.n37 GND 0.06fF
C186 VDD.n38 GND 0.01fF
C187 VDD.n39 GND 0.02fF
C188 VDD.n40 GND 0.27fF
C189 VDD.n41 GND 0.01fF
C190 VDD.n42 GND 0.02fF
C191 VDD.n43 GND 0.03fF
C192 VDD.n44 GND 0.02fF
C193 VDD.n45 GND 0.02fF
C194 VDD.n46 GND 0.02fF
C195 VDD.n47 GND 0.18fF
C196 VDD.n48 GND 0.04fF
C197 VDD.n49 GND 0.04fF
C198 VDD.n50 GND 0.02fF
C199 VDD.n52 GND 0.02fF
C200 VDD.n53 GND 0.02fF
C201 VDD.n54 GND 0.02fF
C202 VDD.n55 GND 0.02fF
C203 VDD.n57 GND 0.02fF
C204 VDD.n58 GND 0.02fF
C205 VDD.n59 GND 0.02fF
C206 VDD.n61 GND 0.27fF
C207 VDD.n63 GND 0.02fF
C208 VDD.n64 GND 0.02fF
C209 VDD.n65 GND 0.03fF
C210 VDD.n66 GND 0.02fF
C211 VDD.n67 GND 0.27fF
C212 VDD.n68 GND 0.01fF
C213 VDD.n69 GND 0.02fF
C214 VDD.n70 GND 0.03fF
C215 VDD.n71 GND 0.27fF
C216 VDD.n72 GND 0.01fF
C217 VDD.n73 GND 0.02fF
C218 VDD.n74 GND 0.02fF
C219 VDD.n75 GND 0.27fF
C220 VDD.n76 GND 0.01fF
C221 VDD.n77 GND 0.02fF
C222 VDD.n78 GND 0.02fF
C223 VDD.n79 GND 0.30fF
C224 VDD.n80 GND 0.01fF
C225 VDD.n81 GND 0.03fF
C226 VDD.n82 GND 0.03fF
C227 VDD.n83 GND 0.17fF
C228 VDD.n84 GND 0.14fF
C229 VDD.n85 GND 0.01fF
C230 VDD.n86 GND 0.02fF
C231 VDD.n87 GND 0.03fF
C232 VDD.n88 GND 0.10fF
C233 VDD.n89 GND 0.02fF
C234 VDD.n90 GND 0.13fF
C235 VDD.n91 GND 0.16fF
C236 VDD.n92 GND 0.01fF
C237 VDD.n93 GND 0.02fF
C238 VDD.n94 GND 0.02fF
C239 VDD.n95 GND 0.24fF
C240 VDD.n96 GND 0.01fF
C241 VDD.n97 GND 0.02fF
C242 VDD.n98 GND 0.02fF
C243 VDD.n99 GND 0.27fF
C244 VDD.n100 GND 0.01fF
C245 VDD.n101 GND 0.02fF
C246 VDD.n102 GND 0.03fF
C247 VDD.n103 GND 0.02fF
C248 VDD.n104 GND 0.02fF
C249 VDD.n105 GND 0.02fF
C250 VDD.n106 GND 0.18fF
C251 VDD.n107 GND 0.04fF
C252 VDD.n108 GND 0.03fF
C253 VDD.n109 GND 0.02fF
C254 VDD.n110 GND 0.02fF
C255 VDD.n111 GND 0.02fF
C256 VDD.n112 GND 0.02fF
C257 VDD.n113 GND 0.02fF
C258 VDD.n115 GND 0.02fF
C259 VDD.n116 GND 0.02fF
C260 VDD.n117 GND 0.02fF
C261 VDD.n119 GND 0.27fF
C262 VDD.n121 GND 0.02fF
C263 VDD.n122 GND 0.02fF
C264 VDD.n123 GND 0.03fF
C265 VDD.n124 GND 0.02fF
C266 VDD.n125 GND 0.27fF
C267 VDD.n126 GND 0.01fF
C268 VDD.n127 GND 0.02fF
C269 VDD.n128 GND 0.03fF
C270 VDD.n129 GND 0.06fF
C271 VDD.n130 GND 0.15fF
C272 VDD.n131 GND 0.20fF
C273 VDD.n132 GND 0.01fF
C274 VDD.n133 GND 0.01fF
C275 VDD.n134 GND 0.02fF
C276 VDD.n135 GND 0.16fF
C277 VDD.n136 GND 0.01fF
C278 VDD.n137 GND 0.02fF
C279 VDD.n138 GND 0.02fF
C280 VDD.n139 GND 0.06fF
C281 VDD.n140 GND 0.15fF
C282 VDD.n141 GND 0.20fF
C283 VDD.n142 GND 0.01fF
C284 VDD.n143 GND 0.01fF
C285 VDD.n144 GND 0.02fF
C286 VDD.n145 GND 0.27fF
C287 VDD.n146 GND 0.01fF
C288 VDD.n147 GND 0.02fF
C289 VDD.n148 GND 0.03fF
C290 VDD.n149 GND 0.02fF
C291 VDD.n150 GND 0.02fF
C292 VDD.n151 GND 0.02fF
C293 VDD.n152 GND 0.18fF
C294 VDD.n153 GND 0.04fF
C295 VDD.n154 GND 0.03fF
C296 VDD.n155 GND 0.02fF
C297 VDD.n156 GND 0.02fF
C298 VDD.n157 GND 0.02fF
C299 VDD.n158 GND 0.02fF
C300 VDD.n159 GND 0.02fF
C301 VDD.n161 GND 0.02fF
C302 VDD.n162 GND 0.02fF
C303 VDD.n163 GND 0.02fF
C304 VDD.n165 GND 0.27fF
C305 VDD.n167 GND 0.02fF
C306 VDD.n168 GND 0.02fF
C307 VDD.n169 GND 0.03fF
C308 VDD.n170 GND 0.02fF
C309 VDD.n171 GND 0.27fF
C310 VDD.n172 GND 0.01fF
C311 VDD.n173 GND 0.02fF
C312 VDD.n174 GND 0.03fF
C313 VDD.n175 GND 0.24fF
C314 VDD.n176 GND 0.01fF
C315 VDD.n177 GND 0.05fF
C316 VDD.n178 GND 0.01fF
C317 VDD.n179 GND 0.02fF
C318 VDD.n180 GND 0.13fF
C319 VDD.n181 GND 0.16fF
C320 VDD.n182 GND 0.01fF
C321 VDD.n183 GND 0.02fF
C322 VDD.n184 GND 0.02fF
C323 VDD.n185 GND 0.30fF
C324 VDD.n186 GND 0.01fF
C325 VDD.n187 GND 0.10fF
C326 VDD.n188 GND 0.02fF
C327 VDD.n189 GND 0.02fF
C328 VDD.n190 GND 0.03fF
C329 VDD.n191 GND 0.17fF
C330 VDD.n192 GND 0.14fF
C331 VDD.n193 GND 0.01fF
C332 VDD.n194 GND 0.02fF
C333 VDD.n195 GND 0.03fF
C334 VDD.n196 GND 0.13fF
C335 VDD.n197 GND 0.16fF
C336 VDD.n198 GND 0.01fF
C337 VDD.n199 GND 0.02fF
C338 VDD.n200 GND 0.02fF
C339 VDD.n201 GND 0.06fF
C340 VDD.n202 GND 0.24fF
C341 VDD.n203 GND 0.01fF
C342 VDD.n204 GND 0.01fF
C343 VDD.n205 GND 0.02fF
C344 VDD.n206 GND 0.27fF
C345 VDD.n207 GND 0.01fF
C346 VDD.n208 GND 0.02fF
C347 VDD.n209 GND 0.03fF
C348 VDD.n210 GND 0.02fF
C349 VDD.n211 GND 0.02fF
C350 VDD.n212 GND 0.02fF
C351 VDD.n213 GND 0.18fF
C352 VDD.n214 GND 0.04fF
C353 VDD.n215 GND 0.03fF
C354 VDD.n216 GND 0.02fF
C355 VDD.n217 GND 0.02fF
C356 VDD.n218 GND 0.02fF
C357 VDD.n219 GND 0.02fF
C358 VDD.n220 GND 0.02fF
C359 VDD.n222 GND 0.02fF
C360 VDD.n223 GND 0.02fF
C361 VDD.n224 GND 0.02fF
C362 VDD.n226 GND 0.27fF
C363 VDD.n228 GND 0.02fF
C364 VDD.n229 GND 0.02fF
C365 VDD.n230 GND 0.03fF
C366 VDD.n231 GND 0.02fF
C367 VDD.n232 GND 0.27fF
C368 VDD.n233 GND 0.01fF
C369 VDD.n234 GND 0.02fF
C370 VDD.n235 GND 0.03fF
C371 VDD.n236 GND 0.06fF
C372 VDD.n237 GND 0.15fF
C373 VDD.n238 GND 0.20fF
C374 VDD.n239 GND 0.01fF
C375 VDD.n240 GND 0.01fF
C376 VDD.n241 GND 0.02fF
C377 VDD.n242 GND 0.16fF
C378 VDD.n243 GND 0.01fF
C379 VDD.n244 GND 0.02fF
C380 VDD.n245 GND 0.02fF
C381 VDD.n246 GND 0.15fF
C382 VDD.n247 GND 0.20fF
C383 VDD.n248 GND 0.01fF
C384 VDD.n249 GND 0.06fF
C385 VDD.n250 GND 0.01fF
C386 VDD.n251 GND 0.02fF
C387 VDD.n252 GND 0.27fF
C388 VDD.n253 GND 0.01fF
C389 VDD.n254 GND 0.02fF
C390 VDD.n255 GND 0.03fF
C391 VDD.n256 GND 0.02fF
C392 VDD.n257 GND 0.02fF
C393 VDD.n258 GND 0.02fF
C394 VDD.n259 GND 0.18fF
C395 VDD.n260 GND 0.04fF
C396 VDD.n261 GND 0.03fF
C397 VDD.n262 GND 0.02fF
C398 VDD.n263 GND 0.02fF
C399 VDD.n264 GND 0.02fF
C400 VDD.n265 GND 0.02fF
C401 VDD.n266 GND 0.02fF
C402 VDD.n268 GND 0.02fF
C403 VDD.n269 GND 0.02fF
C404 VDD.n270 GND 0.02fF
C405 VDD.n272 GND 0.27fF
C406 VDD.n274 GND 0.02fF
C407 VDD.n275 GND 0.02fF
C408 VDD.n276 GND 0.03fF
C409 VDD.n277 GND 0.02fF
C410 VDD.n278 GND 0.27fF
C411 VDD.n279 GND 0.01fF
C412 VDD.n280 GND 0.02fF
C413 VDD.n281 GND 0.03fF
C414 VDD.n282 GND 0.05fF
C415 VDD.n283 GND 0.24fF
C416 VDD.n284 GND 0.01fF
C417 VDD.n285 GND 0.01fF
C418 VDD.n286 GND 0.02fF
C419 VDD.n287 GND 0.13fF
C420 VDD.n288 GND 0.16fF
C421 VDD.n289 GND 0.01fF
C422 VDD.n290 GND 0.02fF
C423 VDD.n291 GND 0.02fF
C424 VDD.n292 GND 0.10fF
C425 VDD.n293 GND 0.02fF
C426 VDD.n294 GND 0.30fF
C427 VDD.n295 GND 0.01fF
C428 VDD.n296 GND 0.02fF
C429 VDD.n297 GND 0.03fF
C430 VDD.n298 GND 0.17fF
C431 VDD.n299 GND 0.14fF
C432 VDD.n300 GND 0.01fF
C433 VDD.n301 GND 0.02fF
C434 VDD.n302 GND 0.03fF
C435 VDD.n303 GND 0.13fF
C436 VDD.n304 GND 0.16fF
C437 VDD.n305 GND 0.01fF
C438 VDD.n306 GND 0.02fF
C439 VDD.n307 GND 0.02fF
C440 VDD.n308 GND 0.06fF
C441 VDD.n309 GND 0.24fF
C442 VDD.n310 GND 0.01fF
C443 VDD.n311 GND 0.01fF
C444 VDD.n312 GND 0.02fF
C445 VDD.n313 GND 0.27fF
C446 VDD.n314 GND 0.01fF
C447 VDD.n315 GND 0.02fF
C448 VDD.n316 GND 0.03fF
C449 VDD.n317 GND 0.02fF
C450 VDD.n318 GND 0.02fF
C451 VDD.n319 GND 0.02fF
C452 VDD.n320 GND 0.18fF
C453 VDD.n321 GND 0.04fF
C454 VDD.n322 GND 0.03fF
C455 VDD.n323 GND 0.02fF
C456 VDD.n324 GND 0.02fF
C457 VDD.n325 GND 0.02fF
C458 VDD.n326 GND 0.02fF
C459 VDD.n327 GND 0.02fF
C460 VDD.n329 GND 0.02fF
C461 VDD.n330 GND 0.02fF
C462 VDD.n331 GND 0.02fF
C463 VDD.n333 GND 0.27fF
C464 VDD.n335 GND 0.02fF
C465 VDD.n336 GND 0.02fF
C466 VDD.n337 GND 0.03fF
C467 VDD.n338 GND 0.02fF
C468 VDD.n339 GND 0.27fF
C469 VDD.n340 GND 0.01fF
C470 VDD.n341 GND 0.02fF
C471 VDD.n342 GND 0.03fF
C472 VDD.n343 GND 0.06fF
C473 VDD.n344 GND 0.15fF
C474 VDD.n345 GND 0.20fF
C475 VDD.n346 GND 0.01fF
C476 VDD.n347 GND 0.01fF
C477 VDD.n348 GND 0.02fF
C478 VDD.n349 GND 0.16fF
C479 VDD.n350 GND 0.01fF
C480 VDD.n351 GND 0.02fF
C481 VDD.n352 GND 0.02fF
C482 VDD.n353 GND 0.06fF
C483 VDD.n354 GND 0.15fF
C484 VDD.n355 GND 0.20fF
C485 VDD.n356 GND 0.01fF
C486 VDD.n357 GND 0.01fF
C487 VDD.n358 GND 0.02fF
C488 VDD.n359 GND 0.27fF
C489 VDD.n360 GND 0.01fF
C490 VDD.n361 GND 0.02fF
C491 VDD.n362 GND 0.03fF
C492 VDD.n363 GND 0.02fF
C493 VDD.n364 GND 0.02fF
C494 VDD.n365 GND 0.02fF
C495 VDD.n366 GND 0.18fF
C496 VDD.n367 GND 0.04fF
C497 VDD.n368 GND 0.03fF
C498 VDD.n369 GND 0.02fF
C499 VDD.n370 GND 0.02fF
C500 VDD.n371 GND 0.02fF
C501 VDD.n372 GND 0.02fF
C502 VDD.n373 GND 0.02fF
C503 VDD.n375 GND 0.02fF
C504 VDD.n376 GND 0.02fF
C505 VDD.n377 GND 0.02fF
C506 VDD.n379 GND 0.27fF
C507 VDD.n381 GND 0.02fF
C508 VDD.n382 GND 0.02fF
C509 VDD.n383 GND 0.03fF
C510 VDD.n384 GND 0.02fF
C511 VDD.n385 GND 0.27fF
C512 VDD.n386 GND 0.01fF
C513 VDD.n387 GND 0.02fF
C514 VDD.n388 GND 0.03fF
C515 VDD.n389 GND 0.02fF
C516 VDD.n390 GND 0.02fF
C517 VDD.n391 GND 0.02fF
C518 VDD.n392 GND 0.12fF
C519 VDD.n393 GND 0.03fF
C520 VDD.n394 GND 0.02fF
C521 VDD.n395 GND 0.02fF
C522 VDD.n396 GND 0.02fF
C523 VDD.n397 GND 0.02fF
C524 VDD.n398 GND 0.02fF
C525 VDD.n400 GND 0.02fF
C526 VDD.n401 GND 0.02fF
C527 VDD.n402 GND 0.02fF
C528 VDD.n404 GND 0.45fF
C529 VDD.n406 GND 0.03fF
C530 VDD.n407 GND 0.03fF
C531 VDD.n408 GND 0.27fF
C532 VDD.n409 GND 0.02fF
C533 VDD.n410 GND 0.03fF
C534 VDD.n411 GND 0.03fF
C535 VDD.n412 GND 0.15fF
C536 VDD.n413 GND 0.20fF
C537 VDD.n414 GND 0.01fF
C538 VDD.n415 GND 0.06fF
C539 VDD.n416 GND 0.01fF
C540 VDD.n417 GND 0.02fF
C541 VDD.n418 GND 0.16fF
C542 VDD.n419 GND 0.01fF
C543 VDD.n420 GND 0.02fF
C544 VDD.n421 GND 0.02fF
C545 VDD.n422 GND 0.06fF
C546 VDD.n423 GND 0.15fF
C547 VDD.n424 GND 0.20fF
C548 VDD.n425 GND 0.01fF
C549 VDD.n426 GND 0.01fF
C550 VDD.n427 GND 0.02fF
C551 VDD.n428 GND 0.27fF
C552 VDD.n429 GND 0.01fF
C553 VDD.n430 GND 0.02fF
C554 VDD.n431 GND 0.03fF
C555 VDD.n432 GND 0.02fF
C556 VDD.n433 GND 0.27fF
C557 VDD.n434 GND 0.01fF
C558 VDD.n435 GND 0.02fF
C559 VDD.n436 GND 0.02fF
C560 VDD.n437 GND 0.02fF
C561 VDD.n438 GND 0.02fF
C562 VDD.n439 GND 0.02fF
C563 VDD.n440 GND 0.02fF
C564 VDD.n442 GND 0.02fF
C565 VDD.n443 GND 0.02fF
C566 VDD.n444 GND 0.02fF
C567 VDD.n445 GND 0.02fF
C568 VDD.n447 GND 0.04fF
C569 VDD.n448 GND 0.02fF
C570 VDD.n449 GND 0.18fF
C571 VDD.n450 GND 0.04fF
C572 VDD.n452 GND 0.27fF
C573 VDD.n454 GND 0.02fF
C574 VDD.n455 GND 0.02fF
C575 VDD.n456 GND 0.03fF
C576 VDD.n457 GND 0.02fF
C577 VDD.n458 GND 0.03fF
C578 VDD.n459 GND 0.24fF
C579 VDD.n460 GND 0.01fF
C580 VDD.n461 GND 0.02fF
C581 VDD.n462 GND 0.02fF
C582 VDD.n463 GND 0.10fF
C583 VDD.n464 GND 0.03fF
C584 VDD.n465 GND 0.13fF
C585 VDD.n466 GND 0.16fF
C586 VDD.n467 GND 0.01fF
C587 VDD.n468 GND 0.02fF
C588 VDD.n469 GND 0.02fF
C589 VDD.n470 GND 0.17fF
C590 VDD.n471 GND 0.14fF
C591 VDD.n472 GND 0.01fF
C592 VDD.n473 GND 0.02fF
C593 VDD.n474 GND 0.03fF
C594 VDD.n475 GND 0.30fF
C595 VDD.n476 GND 0.01fF
C596 VDD.n477 GND 0.03fF
C597 VDD.n478 GND 0.03fF
C598 VDD.n479 GND 0.27fF
C599 VDD.n480 GND 0.01fF
C600 VDD.n481 GND 0.02fF
C601 VDD.n482 GND 0.02fF
C602 VDD.n483 GND 0.27fF
C603 VDD.n484 GND 0.01fF
C604 VDD.n485 GND 0.02fF
C605 VDD.n486 GND 0.02fF
C606 VDD.n487 GND 0.27fF
C607 VDD.n488 GND 0.01fF
C608 VDD.n489 GND 0.02fF
C609 VDD.n490 GND 0.03fF
C610 VDD.n491 GND 0.02fF
C611 VDD.n492 GND 0.27fF
C612 VDD.n493 GND 0.01fF
C613 VDD.n494 GND 0.02fF
C614 VDD.n495 GND 0.02fF
C615 VDD.n496 GND 0.02fF
C616 VDD.n497 GND 0.21fF
C617 VDD.n498 GND 0.04fF
C618 VDD.n499 GND 0.03fF
C619 VDD.n500 GND 0.02fF
C620 VDD.n501 GND 0.02fF
C621 VDD.n502 GND 0.02fF
C622 VDD.n503 GND 0.02fF
C623 VDD.n504 GND 0.02fF
C624 VDD.n506 GND 0.02fF
C625 VDD.n507 GND 0.02fF
C626 VDD.n508 GND 0.02fF
C627 VDD.n510 GND 0.27fF
C628 VDD.n512 GND 0.02fF
C629 VDD.n513 GND 0.02fF
C630 VDD.n514 GND 0.03fF
C631 VDD.n515 GND 0.02fF
C632 VDD.n516 GND 0.03fF
C633 VDD.n517 GND 0.24fF
C634 VDD.n518 GND 0.01fF
C635 VDD.n519 GND 0.02fF
C636 VDD.n520 GND 0.02fF
C637 VDD.n521 GND 0.10fF
C638 VDD.n522 GND 0.03fF
C639 VDD.n523 GND 0.13fF
C640 VDD.n524 GND 0.16fF
C641 VDD.n525 GND 0.01fF
C642 VDD.n526 GND 0.02fF
C643 VDD.n527 GND 0.02fF
C644 VDD.n528 GND 0.17fF
C645 VDD.n529 GND 0.14fF
C646 VDD.n530 GND 0.01fF
C647 VDD.n531 GND 0.02fF
C648 VDD.n532 GND 0.03fF
C649 VDD.n533 GND 0.30fF
C650 VDD.n534 GND 0.01fF
C651 VDD.n535 GND 0.03fF
C652 VDD.n536 GND 0.03fF
C653 VDD.n537 GND 0.27fF
C654 VDD.n538 GND 0.01fF
C655 VDD.n539 GND 0.02fF
C656 VDD.n540 GND 0.02fF
C657 VDD.n541 GND 0.27fF
C658 VDD.n542 GND 0.01fF
C659 VDD.n543 GND 0.02fF
C660 VDD.n544 GND 0.02fF
C661 VDD.n545 GND 0.27fF
C662 VDD.n546 GND 0.01fF
C663 VDD.n547 GND 0.02fF
C664 VDD.n548 GND 0.03fF
C665 VDD.n549 GND 0.02fF
C666 VDD.n550 GND 0.27fF
C667 VDD.n551 GND 0.01fF
C668 VDD.n552 GND 0.02fF
C669 VDD.n553 GND 0.02fF
C670 VDD.n554 GND 0.02fF
C671 VDD.n555 GND 0.18fF
C672 VDD.n556 GND 0.04fF
C673 VDD.n557 GND 0.03fF
C674 VDD.n558 GND 0.02fF
C675 VDD.n559 GND 0.02fF
C676 VDD.n560 GND 0.02fF
C677 VDD.n561 GND 0.02fF
C678 VDD.n562 GND 0.02fF
C679 VDD.n564 GND 0.02fF
C680 VDD.n565 GND 0.02fF
C681 VDD.n566 GND 0.02fF
C682 VDD.n568 GND 0.27fF
C683 VDD.n570 GND 0.02fF
C684 VDD.n571 GND 0.02fF
C685 VDD.n572 GND 0.03fF
C686 VDD.n573 GND 0.02fF
C687 VDD.n574 GND 0.03fF
C688 VDD.n575 GND 0.06fF
C689 VDD.n576 GND 0.15fF
C690 VDD.n577 GND 0.20fF
C691 VDD.n578 GND 0.01fF
C692 VDD.n579 GND 0.01fF
C693 VDD.n580 GND 0.02fF
C694 VDD.n581 GND 0.16fF
C695 VDD.n582 GND 0.01fF
C696 VDD.n583 GND 0.02fF
C697 VDD.n584 GND 0.02fF
C698 VDD.n585 GND 0.06fF
C699 VDD.n586 GND 0.15fF
C700 VDD.n587 GND 0.20fF
C701 VDD.n588 GND 0.01fF
C702 VDD.n589 GND 0.01fF
C703 VDD.n590 GND 0.02fF
C704 VDD.n591 GND 0.27fF
C705 VDD.n592 GND 0.01fF
C706 VDD.n593 GND 0.02fF
C707 VDD.n594 GND 0.03fF
C708 VDD.n595 GND 0.02fF
C709 VDD.n596 GND 0.02fF
C710 VDD.n597 GND 0.02fF
C711 VDD.n598 GND 0.14fF
C712 VDD.n599 GND 0.04fF
C713 VDD.n600 GND 0.03fF
C714 VDD.n601 GND 0.02fF
C715 VDD.n602 GND 0.02fF
C716 VDD.n603 GND 0.02fF
C717 VDD.n604 GND 0.02fF
C718 VDD.n605 GND 0.02fF
C719 VDD.n607 GND 0.02fF
C720 VDD.n608 GND 0.02fF
C721 VDD.n609 GND 0.02fF
C722 VDD.n611 GND 0.27fF
C723 VDD.n613 GND 0.02fF
C724 VDD.n614 GND 0.02fF
C725 VDD.n615 GND 0.03fF
C726 VDD.n616 GND 0.02fF
C727 VDD.n617 GND 0.27fF
C728 VDD.n618 GND 0.01fF
C729 VDD.n619 GND 0.02fF
C730 VDD.n620 GND 0.03fF
C731 VDD.n621 GND 0.15fF
C732 VDD.n622 GND 0.20fF
C733 VDD.n623 GND 0.01fF
C734 VDD.n624 GND 0.06fF
C735 VDD.n625 GND 0.01fF
C736 VDD.n626 GND 0.02fF
C737 VDD.n627 GND 0.16fF
C738 VDD.n628 GND 0.01fF
C739 VDD.n629 GND 0.02fF
C740 VDD.n630 GND 0.02fF
C741 VDD.n631 GND 0.06fF
C742 VDD.n632 GND 0.15fF
C743 VDD.n633 GND 0.20fF
C744 VDD.n634 GND 0.01fF
C745 VDD.n635 GND 0.01fF
C746 VDD.n636 GND 0.02fF
C747 VDD.n637 GND 0.27fF
C748 VDD.n638 GND 0.01fF
C749 VDD.n639 GND 0.02fF
C750 VDD.n640 GND 0.03fF
C751 VDD.n641 GND 0.02fF
C752 VDD.n642 GND 0.27fF
C753 VDD.n643 GND 0.01fF
C754 VDD.n644 GND 0.02fF
C755 VDD.n645 GND 0.02fF
C756 VDD.n646 GND 0.02fF
C757 VDD.n647 GND 0.18fF
C758 VDD.n648 GND 0.04fF
C759 VDD.n649 GND 0.03fF
C760 VDD.n650 GND 0.02fF
C761 VDD.n651 GND 0.02fF
C762 VDD.n652 GND 0.02fF
C763 VDD.n653 GND 0.02fF
C764 VDD.n654 GND 0.02fF
C765 VDD.n656 GND 0.02fF
C766 VDD.n657 GND 0.02fF
C767 VDD.n658 GND 0.02fF
C768 VDD.n660 GND 0.27fF
C769 VDD.n662 GND 0.02fF
C770 VDD.n663 GND 0.02fF
C771 VDD.n664 GND 0.03fF
C772 VDD.n665 GND 0.02fF
C773 VDD.n666 GND 0.03fF
C774 VDD.n667 GND 0.24fF
C775 VDD.n668 GND 0.01fF
C776 VDD.n669 GND 0.02fF
C777 VDD.n670 GND 0.02fF
C778 VDD.n671 GND 0.10fF
C779 VDD.n672 GND 0.03fF
C780 VDD.n673 GND 0.13fF
C781 VDD.n674 GND 0.16fF
C782 VDD.n675 GND 0.01fF
C783 VDD.n676 GND 0.02fF
C784 VDD.n677 GND 0.02fF
C785 VDD.n678 GND 0.17fF
C786 VDD.n679 GND 0.14fF
C787 VDD.n680 GND 0.01fF
C788 VDD.n681 GND 0.02fF
C789 VDD.n682 GND 0.03fF
C790 VDD.n683 GND 0.30fF
C791 VDD.n684 GND 0.01fF
C792 VDD.n685 GND 0.03fF
C793 VDD.n686 GND 0.03fF
C794 VDD.n687 GND 0.27fF
C795 VDD.n688 GND 0.01fF
C796 VDD.n689 GND 0.02fF
C797 VDD.n690 GND 0.02fF
C798 VDD.n691 GND 0.27fF
C799 VDD.n692 GND 0.01fF
C800 VDD.n693 GND 0.02fF
C801 VDD.n694 GND 0.02fF
C802 VDD.n695 GND 0.27fF
C803 VDD.n696 GND 0.01fF
C804 VDD.n697 GND 0.02fF
C805 VDD.n698 GND 0.03fF
C806 VDD.n699 GND 0.02fF
C807 VDD.n700 GND 0.27fF
C808 VDD.n701 GND 0.01fF
C809 VDD.n702 GND 0.02fF
C810 VDD.n703 GND 0.02fF
C811 VDD.n704 GND 0.02fF
C812 VDD.n705 GND 0.21fF
C813 VDD.n706 GND 0.04fF
C814 VDD.n707 GND 0.03fF
C815 VDD.n708 GND 0.02fF
C816 VDD.n709 GND 0.02fF
C817 VDD.n710 GND 0.02fF
C818 VDD.n711 GND 0.02fF
C819 VDD.n712 GND 0.02fF
C820 VDD.n714 GND 0.02fF
C821 VDD.n715 GND 0.02fF
C822 VDD.n716 GND 0.02fF
C823 VDD.n718 GND 0.27fF
C824 VDD.n720 GND 0.02fF
C825 VDD.n721 GND 0.02fF
C826 VDD.n722 GND 0.03fF
C827 VDD.n723 GND 0.02fF
C828 VDD.n724 GND 0.03fF
C829 VDD.n725 GND 0.24fF
C830 VDD.n726 GND 0.01fF
C831 VDD.n727 GND 0.02fF
C832 VDD.n728 GND 0.02fF
C833 VDD.n729 GND 0.10fF
C834 VDD.n730 GND 0.03fF
C835 VDD.n731 GND 0.13fF
C836 VDD.n732 GND 0.16fF
C837 VDD.n733 GND 0.01fF
C838 VDD.n734 GND 0.02fF
C839 VDD.n735 GND 0.02fF
C840 VDD.n736 GND 0.17fF
C841 VDD.n737 GND 0.14fF
C842 VDD.n738 GND 0.01fF
C843 VDD.n739 GND 0.02fF
C844 VDD.n740 GND 0.03fF
C845 VDD.n741 GND 0.30fF
C846 VDD.n742 GND 0.01fF
C847 VDD.n743 GND 0.03fF
C848 VDD.n744 GND 0.03fF
C849 VDD.n745 GND 0.27fF
C850 VDD.n746 GND 0.01fF
C851 VDD.n747 GND 0.02fF
C852 VDD.n748 GND 0.02fF
C853 VDD.n749 GND 0.27fF
C854 VDD.n750 GND 0.01fF
C855 VDD.n751 GND 0.02fF
C856 VDD.n752 GND 0.02fF
.ends
