// File: DFFSNRNX1.spi.DFFSNRNX1.pxi
// Created: Tue Oct 15 15:47:46 2024
// 
simulator lang=spectre
x_PM_DFFSNRNX1\%GND ( GND N_GND_c_8_p N_GND_c_118_p N_GND_c_1_p N_GND_c_9_p \
 N_GND_c_10_p N_GND_c_14_p N_GND_c_15_p N_GND_c_38_p N_GND_c_45_p N_GND_c_52_p \
 N_GND_c_65_p N_GND_c_72_p N_GND_c_84_p N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p \
 N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p N_GND_M0_noxref_d N_GND_M3_noxref_d \
 N_GND_M6_noxref_d N_GND_M9_noxref_d N_GND_M12_noxref_d N_GND_M15_noxref_d )  \
 PM_DFFSNRNX1\%GND
x_PM_DFFSNRNX1\%VDD ( VDD N_VDD_c_316_p N_VDD_c_309_n N_VDD_c_317_p \
 N_VDD_c_318_p N_VDD_c_324_p N_VDD_c_328_p N_VDD_c_462_p N_VDD_c_337_p \
 N_VDD_c_407_p N_VDD_c_425_p N_VDD_c_429_p N_VDD_c_465_p N_VDD_c_341_p \
 N_VDD_c_366_p N_VDD_c_372_p N_VDD_c_376_p N_VDD_c_468_p N_VDD_c_382_p \
 N_VDD_c_411_p N_VDD_c_493_p N_VDD_c_478_p N_VDD_c_479_p N_VDD_c_439_p \
 N_VDD_c_497_p N_VDD_c_510_p N_VDD_c_514_p N_VDD_c_556_p N_VDD_c_519_p \
 N_VDD_c_548_p N_VDD_c_588_p N_VDD_c_310_n N_VDD_c_311_n N_VDD_c_312_n \
 N_VDD_c_313_n N_VDD_c_314_n N_VDD_c_315_n N_VDD_M18_noxref_s \
 N_VDD_M19_noxref_d N_VDD_M21_noxref_d N_VDD_M23_noxref_d N_VDD_M24_noxref_s \
 N_VDD_M25_noxref_d N_VDD_M27_noxref_d N_VDD_M29_noxref_d N_VDD_M30_noxref_s \
 N_VDD_M31_noxref_d N_VDD_M33_noxref_d N_VDD_M35_noxref_d N_VDD_M36_noxref_s \
 N_VDD_M37_noxref_d N_VDD_M39_noxref_d N_VDD_M41_noxref_d N_VDD_M42_noxref_s \
 N_VDD_M43_noxref_d N_VDD_M45_noxref_d N_VDD_M47_noxref_d N_VDD_M48_noxref_s \
 N_VDD_M49_noxref_d N_VDD_M51_noxref_d N_VDD_M53_noxref_d )  PM_DFFSNRNX1\%VDD
x_PM_DFFSNRNX1\%noxref_3 ( N_noxref_3_c_651_n N_noxref_3_c_655_n \
 N_noxref_3_c_656_n N_noxref_3_c_660_n N_noxref_3_c_685_n N_noxref_3_c_689_n \
 N_noxref_3_c_691_n N_noxref_3_c_695_n N_noxref_3_c_661_n N_noxref_3_c_770_p \
 N_noxref_3_c_699_n N_noxref_3_c_662_n N_noxref_3_c_663_n N_noxref_3_c_817_p \
 N_noxref_3_c_781_p N_noxref_3_M3_noxref_g N_noxref_3_M6_noxref_g \
 N_noxref_3_M24_noxref_g N_noxref_3_M25_noxref_g N_noxref_3_M30_noxref_g \
 N_noxref_3_M31_noxref_g N_noxref_3_c_664_n N_noxref_3_c_666_n \
 N_noxref_3_c_667_n N_noxref_3_c_668_n N_noxref_3_c_669_n N_noxref_3_c_670_n \
 N_noxref_3_c_671_n N_noxref_3_c_673_n N_noxref_3_c_747_p N_noxref_3_c_714_n \
 N_noxref_3_c_674_n N_noxref_3_c_676_n N_noxref_3_c_677_n N_noxref_3_c_678_n \
 N_noxref_3_c_679_n N_noxref_3_c_680_n N_noxref_3_c_681_n N_noxref_3_c_683_n \
 N_noxref_3_c_736_p N_noxref_3_c_716_n N_noxref_3_M2_noxref_d \
 N_noxref_3_M18_noxref_d N_noxref_3_M20_noxref_d N_noxref_3_M22_noxref_d )  \
 PM_DFFSNRNX1\%noxref_3
x_PM_DFFSNRNX1\%noxref_4 ( N_noxref_4_c_902_n N_noxref_4_c_955_n \
 N_noxref_4_c_916_n N_noxref_4_c_920_n N_noxref_4_c_922_n N_noxref_4_c_926_n \
 N_noxref_4_c_903_n N_noxref_4_c_1000_p N_noxref_4_c_930_n N_noxref_4_c_904_n \
 N_noxref_4_c_1010_p N_noxref_4_c_1018_p N_noxref_4_M9_noxref_g \
 N_noxref_4_M36_noxref_g N_noxref_4_M37_noxref_g N_noxref_4_c_905_n \
 N_noxref_4_c_907_n N_noxref_4_c_908_n N_noxref_4_c_909_n N_noxref_4_c_910_n \
 N_noxref_4_c_911_n N_noxref_4_c_912_n N_noxref_4_c_914_n N_noxref_4_c_968_p \
 N_noxref_4_c_938_n N_noxref_4_M8_noxref_d N_noxref_4_M30_noxref_d \
 N_noxref_4_M32_noxref_d N_noxref_4_M34_noxref_d )  PM_DFFSNRNX1\%noxref_4
x_PM_DFFSNRNX1\%CLK ( N_CLK_c_1062_n N_CLK_c_1079_n CLK CLK CLK CLK CLK \
 N_CLK_c_1063_n N_CLK_c_1064_n N_CLK_M4_noxref_g N_CLK_M10_noxref_g \
 N_CLK_M26_noxref_g N_CLK_M27_noxref_g N_CLK_M38_noxref_g N_CLK_M39_noxref_g \
 N_CLK_c_1091_n N_CLK_c_1094_n N_CLK_c_1218_p N_CLK_c_1225_p N_CLK_c_1096_n \
 N_CLK_c_1097_n N_CLK_c_1098_n N_CLK_c_1099_n N_CLK_c_1143_p N_CLK_c_1118_n \
 N_CLK_c_1121_n N_CLK_c_1241_p N_CLK_c_1248_p N_CLK_c_1123_n N_CLK_c_1124_n \
 N_CLK_c_1125_n N_CLK_c_1126_n N_CLK_c_1151_p N_CLK_c_1102_n N_CLK_c_1128_n )  \
 PM_DFFSNRNX1\%CLK
x_PM_DFFSNRNX1\%noxref_6 ( N_noxref_6_c_1253_n N_noxref_6_c_1254_n \
 N_noxref_6_c_1255_n N_noxref_6_c_1325_n N_noxref_6_c_1256_n \
 N_noxref_6_c_1272_n N_noxref_6_c_1276_n N_noxref_6_c_1278_n \
 N_noxref_6_c_1282_n N_noxref_6_c_1257_n N_noxref_6_c_1335_n \
 N_noxref_6_c_1286_n N_noxref_6_c_1258_n N_noxref_6_c_1375_n \
 N_noxref_6_c_1457_p N_noxref_6_M2_noxref_g N_noxref_6_M12_noxref_g \
 N_noxref_6_M22_noxref_g N_noxref_6_M23_noxref_g N_noxref_6_M42_noxref_g \
 N_noxref_6_M43_noxref_g N_noxref_6_c_1342_n N_noxref_6_c_1343_n \
 N_noxref_6_c_1344_n N_noxref_6_c_1345_n N_noxref_6_c_1346_n \
 N_noxref_6_c_1348_n N_noxref_6_c_1349_n N_noxref_6_c_1259_n \
 N_noxref_6_c_1261_n N_noxref_6_c_1262_n N_noxref_6_c_1263_n \
 N_noxref_6_c_1264_n N_noxref_6_c_1265_n N_noxref_6_c_1266_n \
 N_noxref_6_c_1268_n N_noxref_6_c_1402_p N_noxref_6_c_1298_n \
 N_noxref_6_c_1351_n N_noxref_6_c_1352_n N_noxref_6_c_1354_n \
 N_noxref_6_M5_noxref_d N_noxref_6_M24_noxref_d N_noxref_6_M26_noxref_d \
 N_noxref_6_M28_noxref_d )  PM_DFFSNRNX1\%noxref_6
x_PM_DFFSNRNX1\%RN ( N_RN_c_1514_n N_RN_c_1515_n N_RN_c_1536_n N_RN_c_1542_n \
 RN RN RN RN RN RN RN RN RN RN RN RN RN N_RN_c_1516_n N_RN_c_1517_n \
 N_RN_c_1518_n N_RN_M1_noxref_g N_RN_M11_noxref_g N_RN_M13_noxref_g \
 N_RN_M20_noxref_g N_RN_M21_noxref_g N_RN_M40_noxref_g N_RN_M41_noxref_g \
 N_RN_M44_noxref_g N_RN_M45_noxref_g N_RN_c_1755_p N_RN_c_1757_p N_RN_c_1781_p \
 N_RN_c_1788_p N_RN_c_1644_n N_RN_c_1645_n N_RN_c_1646_n N_RN_c_1647_n \
 N_RN_c_1578_n N_RN_c_1603_n N_RN_c_1604_n N_RN_c_1605_n N_RN_c_1724_p \
 N_RN_c_1706_p N_RN_c_1726_p N_RN_c_1707_p N_RN_c_1651_n N_RN_c_1654_n \
 N_RN_c_1811_p N_RN_c_1818_p N_RN_c_1656_n N_RN_c_1657_n N_RN_c_1658_n \
 N_RN_c_1659_n N_RN_c_1674_p N_RN_c_1579_n N_RN_c_1606_n N_RN_c_1608_n \
 N_RN_c_1609_n N_RN_c_1663_n )  PM_DFFSNRNX1\%RN
x_PM_DFFSNRNX1\%QN ( N_QN_c_1823_n N_QN_c_1892_p QN QN QN QN QN QN QN QN \
 N_QN_c_1838_n N_QN_c_1842_n N_QN_c_1844_n N_QN_c_1848_n N_QN_c_1824_n \
 N_QN_c_1894_p N_QN_c_1825_n N_QN_c_1887_n N_QN_c_1936_p N_QN_M15_noxref_g \
 N_QN_M48_noxref_g N_QN_M49_noxref_g N_QN_c_1826_n N_QN_c_1828_n N_QN_c_1829_n \
 N_QN_c_1830_n N_QN_c_1831_n N_QN_c_1832_n N_QN_c_1833_n N_QN_c_1835_n \
 N_QN_c_1901_p N_QN_c_1859_n N_QN_M14_noxref_d N_QN_M42_noxref_d \
 N_QN_M44_noxref_d N_QN_M46_noxref_d )  PM_DFFSNRNX1\%QN
x_PM_DFFSNRNX1\%SN ( N_SN_c_1980_n N_SN_c_1990_n SN SN SN SN SN SN \
 N_SN_c_1991_n N_SN_c_1992_n N_SN_M7_noxref_g N_SN_M16_noxref_g \
 N_SN_M32_noxref_g N_SN_M33_noxref_g N_SN_M50_noxref_g N_SN_M51_noxref_g \
 N_SN_c_2014_n N_SN_c_2017_n N_SN_c_2157_p N_SN_c_2165_p N_SN_c_2019_n \
 N_SN_c_2020_n N_SN_c_2021_n N_SN_c_2022_n N_SN_c_2039_n N_SN_c_2075_n \
 N_SN_c_2078_n N_SN_c_2197_p N_SN_c_2204_p N_SN_c_2080_n N_SN_c_2081_n \
 N_SN_c_2082_n N_SN_c_2083_n N_SN_c_2093_p N_SN_c_2024_n N_SN_c_2085_n )  \
 PM_DFFSNRNX1\%SN
x_PM_DFFSNRNX1\%noxref_10 ( N_noxref_10_c_2214_n N_noxref_10_c_2308_n \
 N_noxref_10_c_2215_n N_noxref_10_c_2278_n N_noxref_10_c_2216_n \
 N_noxref_10_c_2223_n N_noxref_10_c_2209_n N_noxref_10_c_2317_n \
 N_noxref_10_c_2210_n N_noxref_10_c_2225_n N_noxref_10_c_2229_n \
 N_noxref_10_c_2231_n N_noxref_10_c_2235_n N_noxref_10_c_2211_n \
 N_noxref_10_c_2450_n N_noxref_10_c_2239_n N_noxref_10_c_2212_n \
 N_noxref_10_c_2241_n N_noxref_10_c_2326_n N_noxref_10_c_2413_n \
 N_noxref_10_M5_noxref_g N_noxref_10_M8_noxref_g N_noxref_10_M17_noxref_g \
 N_noxref_10_M28_noxref_g N_noxref_10_M29_noxref_g N_noxref_10_M34_noxref_g \
 N_noxref_10_M35_noxref_g N_noxref_10_M52_noxref_g N_noxref_10_M53_noxref_g \
 N_noxref_10_c_2330_n N_noxref_10_c_2331_n N_noxref_10_c_2332_n \
 N_noxref_10_c_2370_n N_noxref_10_c_2371_n N_noxref_10_c_2373_n \
 N_noxref_10_c_2374_n N_noxref_10_c_2291_n N_noxref_10_c_2292_n \
 N_noxref_10_c_2293_n N_noxref_10_c_2294_n N_noxref_10_c_2295_n \
 N_noxref_10_c_2297_n N_noxref_10_c_2298_n N_noxref_10_c_2465_n \
 N_noxref_10_c_2466_n N_noxref_10_c_2467_n N_noxref_10_c_2506_p \
 N_noxref_10_c_2497_p N_noxref_10_c_2508_p N_noxref_10_c_2498_p \
 N_noxref_10_c_2275_n N_noxref_10_c_2335_n N_noxref_10_c_2336_n \
 N_noxref_10_c_2300_n N_noxref_10_c_2301_n N_noxref_10_c_2303_n \
 N_noxref_10_c_2475_n N_noxref_10_c_2477_n N_noxref_10_c_2478_n \
 N_noxref_10_M11_noxref_d N_noxref_10_M36_noxref_d N_noxref_10_M38_noxref_d \
 N_noxref_10_M40_noxref_d )  PM_DFFSNRNX1\%noxref_10
x_PM_DFFSNRNX1\%Q ( N_Q_c_2549_n N_Q_c_2588_n Q Q Q Q Q Q Q Q Q Q Q Q Q \
 N_Q_c_2550_n N_Q_c_2556_n N_Q_c_2560_n N_Q_c_2562_n N_Q_c_2566_n N_Q_c_2551_n \
 N_Q_c_2701_p N_Q_c_2649_n N_Q_c_2671_n N_Q_M14_noxref_g N_Q_M46_noxref_g \
 N_Q_M47_noxref_g N_Q_c_2598_n N_Q_c_2599_n N_Q_c_2600_n N_Q_c_2627_n \
 N_Q_c_2628_n N_Q_c_2630_n N_Q_c_2631_n N_Q_c_2601_n N_Q_c_2603_n N_Q_c_2604_n \
 N_Q_M17_noxref_d N_Q_M48_noxref_d N_Q_M50_noxref_d N_Q_M52_noxref_d )  \
 PM_DFFSNRNX1\%Q
x_PM_DFFSNRNX1\%D ( D D D D D D N_D_c_2706_n N_D_M0_noxref_g N_D_M18_noxref_g \
 N_D_M19_noxref_g N_D_c_2707_n N_D_c_2709_n N_D_c_2710_n N_D_c_2711_n \
 N_D_c_2712_n N_D_c_2713_n N_D_c_2714_n N_D_c_2716_n N_D_c_2729_n N_D_c_2724_n \
 )  PM_DFFSNRNX1\%D
x_PM_DFFSNRNX1\%noxref_13 ( N_noxref_13_c_2790_n N_noxref_13_c_2762_n \
 N_noxref_13_c_2766_n N_noxref_13_c_2769_n N_noxref_13_c_2781_n \
 N_noxref_13_M0_noxref_s )  PM_DFFSNRNX1\%noxref_13
x_PM_DFFSNRNX1\%noxref_14 ( N_noxref_14_c_2808_n N_noxref_14_c_2811_n \
 N_noxref_14_c_2814_n N_noxref_14_c_2817_n N_noxref_14_c_2825_n \
 N_noxref_14_M1_noxref_d N_noxref_14_M2_noxref_s )  PM_DFFSNRNX1\%noxref_14
x_PM_DFFSNRNX1\%noxref_15 ( N_noxref_15_c_2877_n N_noxref_15_c_2861_n \
 N_noxref_15_c_2865_n N_noxref_15_c_2868_n N_noxref_15_c_2888_n \
 N_noxref_15_M3_noxref_s )  PM_DFFSNRNX1\%noxref_15
x_PM_DFFSNRNX1\%noxref_16 ( N_noxref_16_c_2913_n N_noxref_16_c_2916_n \
 N_noxref_16_c_2919_n N_noxref_16_c_2922_n N_noxref_16_c_2945_n \
 N_noxref_16_M4_noxref_d N_noxref_16_M5_noxref_s )  PM_DFFSNRNX1\%noxref_16
x_PM_DFFSNRNX1\%noxref_17 ( N_noxref_17_c_2983_n N_noxref_17_c_2967_n \
 N_noxref_17_c_2971_n N_noxref_17_c_2974_n N_noxref_17_c_2997_n \
 N_noxref_17_M6_noxref_s )  PM_DFFSNRNX1\%noxref_17
x_PM_DFFSNRNX1\%noxref_18 ( N_noxref_18_c_3021_n N_noxref_18_c_3024_n \
 N_noxref_18_c_3027_n N_noxref_18_c_3030_n N_noxref_18_c_3038_n \
 N_noxref_18_M7_noxref_d N_noxref_18_M8_noxref_s )  PM_DFFSNRNX1\%noxref_18
x_PM_DFFSNRNX1\%noxref_19 ( N_noxref_19_c_3091_n N_noxref_19_c_3075_n \
 N_noxref_19_c_3079_n N_noxref_19_c_3082_n N_noxref_19_c_3105_n \
 N_noxref_19_M9_noxref_s )  PM_DFFSNRNX1\%noxref_19
x_PM_DFFSNRNX1\%noxref_20 ( N_noxref_20_c_3125_n N_noxref_20_c_3128_n \
 N_noxref_20_c_3131_n N_noxref_20_c_3134_n N_noxref_20_c_3156_n \
 N_noxref_20_M10_noxref_d N_noxref_20_M11_noxref_s )  PM_DFFSNRNX1\%noxref_20
x_PM_DFFSNRNX1\%noxref_21 ( N_noxref_21_c_3195_n N_noxref_21_c_3179_n \
 N_noxref_21_c_3183_n N_noxref_21_c_3186_n N_noxref_21_c_3207_n \
 N_noxref_21_M12_noxref_s )  PM_DFFSNRNX1\%noxref_21
x_PM_DFFSNRNX1\%noxref_22 ( N_noxref_22_c_3229_n N_noxref_22_c_3232_n \
 N_noxref_22_c_3235_n N_noxref_22_c_3238_n N_noxref_22_c_3258_n \
 N_noxref_22_M13_noxref_d N_noxref_22_M14_noxref_s )  PM_DFFSNRNX1\%noxref_22
x_PM_DFFSNRNX1\%noxref_23 ( N_noxref_23_c_3297_n N_noxref_23_c_3283_n \
 N_noxref_23_c_3287_n N_noxref_23_c_3290_n N_noxref_23_c_3313_n \
 N_noxref_23_M15_noxref_s )  PM_DFFSNRNX1\%noxref_23
x_PM_DFFSNRNX1\%noxref_24 ( N_noxref_24_c_3333_n N_noxref_24_c_3335_n \
 N_noxref_24_c_3338_n N_noxref_24_c_3340_n N_noxref_24_c_3361_n \
 N_noxref_24_M16_noxref_d N_noxref_24_M17_noxref_s )  PM_DFFSNRNX1\%noxref_24
cc_1 ( N_GND_c_1_p N_VDD_c_309_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_310_n ) capacitor c=0.00989031f //x=28.12 //y=0 \
 //x2=28.12 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_311_n ) capacitor c=0.00891658f //x=4.81 //y=0 \
 //x2=4.81 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_312_n ) capacitor c=0.00474978f //x=9.62 //y=0 \
 //x2=9.62 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_313_n ) capacitor c=0.0057235f //x=14.43 //y=0 \
 //x2=14.43 //y2=7.4
cc_6 ( N_GND_c_6_p N_VDD_c_314_n ) capacitor c=0.0057235f //x=19.24 //y=0 \
 //x2=19.24 //y2=7.4
cc_7 ( N_GND_c_7_p N_VDD_c_315_n ) capacitor c=0.0057235f //x=24.05 //y=0 \
 //x2=24.05 //y2=7.4
cc_8 ( N_GND_c_8_p N_noxref_3_c_651_n ) capacitor c=0.0137933f //x=28.12 //y=0 \
 //x2=5.805 //y2=2.965
cc_9 ( N_GND_c_9_p N_noxref_3_c_651_n ) capacitor c=0.0019736f //x=4.64 //y=0 \
 //x2=5.805 //y2=2.965
cc_10 ( N_GND_c_10_p N_noxref_3_c_651_n ) capacitor c=0.00184044f //x=5.8 \
 //y=0 //x2=5.805 //y2=2.965
cc_11 ( N_GND_c_3_p N_noxref_3_c_651_n ) capacitor c=0.014386f //x=4.81 //y=0 \
 //x2=5.805 //y2=2.965
cc_12 ( N_GND_c_8_p N_noxref_3_c_655_n ) capacitor c=0.00197533f //x=28.12 \
 //y=0 //x2=4.185 //y2=2.965
cc_13 ( N_GND_c_8_p N_noxref_3_c_656_n ) capacitor c=0.0371387f //x=28.12 \
 //y=0 //x2=10.615 //y2=2.965
cc_14 ( N_GND_c_14_p N_noxref_3_c_656_n ) capacitor c=0.00285709f //x=9.45 \
 //y=0 //x2=10.615 //y2=2.965
cc_15 ( N_GND_c_15_p N_noxref_3_c_656_n ) capacitor c=0.00184044f //x=10.61 \
 //y=0 //x2=10.615 //y2=2.965
cc_16 ( N_GND_c_4_p N_noxref_3_c_656_n ) capacitor c=0.014386f //x=9.62 //y=0 \
 //x2=10.615 //y2=2.965
cc_17 ( N_GND_c_8_p N_noxref_3_c_660_n ) capacitor c=0.00182434f //x=28.12 \
 //y=0 //x2=6.035 //y2=2.965
cc_18 ( N_GND_c_3_p N_noxref_3_c_661_n ) capacitor c=0.0459494f //x=4.81 //y=0 \
 //x2=3.985 //y2=1.665
cc_19 ( N_GND_c_3_p N_noxref_3_c_662_n ) capacitor c=0.0179249f //x=4.81 //y=0 \
 //x2=5.92 //y2=2.08
cc_20 ( N_GND_c_4_p N_noxref_3_c_663_n ) capacitor c=0.0176137f //x=9.62 //y=0 \
 //x2=10.73 //y2=2.08
cc_21 ( N_GND_c_10_p N_noxref_3_c_664_n ) capacitor c=0.00132755f //x=5.8 \
 //y=0 //x2=5.62 //y2=0.875
cc_22 ( N_GND_M3_noxref_d N_noxref_3_c_664_n ) capacitor c=0.00211996f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=0.875
cc_23 ( N_GND_M3_noxref_d N_noxref_3_c_666_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=1.22
cc_24 ( N_GND_c_3_p N_noxref_3_c_667_n ) capacitor c=0.00204716f //x=4.81 \
 //y=0 //x2=5.62 //y2=1.53
cc_25 ( N_GND_c_3_p N_noxref_3_c_668_n ) capacitor c=0.0126573f //x=4.81 //y=0 \
 //x2=5.62 //y2=1.915
cc_26 ( N_GND_M3_noxref_d N_noxref_3_c_669_n ) capacitor c=0.0131341f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=0.72
cc_27 ( N_GND_M3_noxref_d N_noxref_3_c_670_n ) capacitor c=0.00193146f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=1.375
cc_28 ( N_GND_c_14_p N_noxref_3_c_671_n ) capacitor c=0.00129018f //x=9.45 \
 //y=0 //x2=6.15 //y2=0.875
cc_29 ( N_GND_M3_noxref_d N_noxref_3_c_671_n ) capacitor c=0.00257848f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=0.875
cc_30 ( N_GND_M3_noxref_d N_noxref_3_c_673_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=1.22
cc_31 ( N_GND_c_15_p N_noxref_3_c_674_n ) capacitor c=0.00132755f //x=10.61 \
 //y=0 //x2=10.43 //y2=0.875
cc_32 ( N_GND_M6_noxref_d N_noxref_3_c_674_n ) capacitor c=0.00211996f \
 //x=10.505 //y=0.875 //x2=10.43 //y2=0.875
cc_33 ( N_GND_M6_noxref_d N_noxref_3_c_676_n ) capacitor c=0.00255985f \
 //x=10.505 //y=0.875 //x2=10.43 //y2=1.22
cc_34 ( N_GND_c_4_p N_noxref_3_c_677_n ) capacitor c=0.00204716f //x=9.62 \
 //y=0 //x2=10.43 //y2=1.53
cc_35 ( N_GND_c_4_p N_noxref_3_c_678_n ) capacitor c=0.0126573f //x=9.62 //y=0 \
 //x2=10.43 //y2=1.915
cc_36 ( N_GND_M6_noxref_d N_noxref_3_c_679_n ) capacitor c=0.0131341f \
 //x=10.505 //y=0.875 //x2=10.805 //y2=0.72
cc_37 ( N_GND_M6_noxref_d N_noxref_3_c_680_n ) capacitor c=0.00193146f \
 //x=10.505 //y=0.875 //x2=10.805 //y2=1.375
cc_38 ( N_GND_c_38_p N_noxref_3_c_681_n ) capacitor c=0.00129018f //x=14.26 \
 //y=0 //x2=10.96 //y2=0.875
cc_39 ( N_GND_M6_noxref_d N_noxref_3_c_681_n ) capacitor c=0.00257848f \
 //x=10.505 //y=0.875 //x2=10.96 //y2=0.875
cc_40 ( N_GND_M6_noxref_d N_noxref_3_c_683_n ) capacitor c=0.00255985f \
 //x=10.505 //y=0.875 //x2=10.96 //y2=1.22
cc_41 ( N_GND_c_3_p N_noxref_3_M2_noxref_d ) capacitor c=0.00591582f //x=4.81 \
 //y=0 //x2=3.395 //y2=0.915
cc_42 ( N_GND_c_5_p N_noxref_4_c_902_n ) capacitor c=0.00750857f //x=14.43 \
 //y=0 //x2=15.425 //y2=2.96
cc_43 ( N_GND_c_5_p N_noxref_4_c_903_n ) capacitor c=0.0432345f //x=14.43 \
 //y=0 //x2=13.605 //y2=1.665
cc_44 ( N_GND_c_5_p N_noxref_4_c_904_n ) capacitor c=0.0153336f //x=14.43 \
 //y=0 //x2=15.54 //y2=2.08
cc_45 ( N_GND_c_45_p N_noxref_4_c_905_n ) capacitor c=0.00132755f //x=15.42 \
 //y=0 //x2=15.24 //y2=0.875
cc_46 ( N_GND_M9_noxref_d N_noxref_4_c_905_n ) capacitor c=0.00211996f \
 //x=15.315 //y=0.875 //x2=15.24 //y2=0.875
cc_47 ( N_GND_M9_noxref_d N_noxref_4_c_907_n ) capacitor c=0.00255985f \
 //x=15.315 //y=0.875 //x2=15.24 //y2=1.22
cc_48 ( N_GND_c_5_p N_noxref_4_c_908_n ) capacitor c=0.00204716f //x=14.43 \
 //y=0 //x2=15.24 //y2=1.53
cc_49 ( N_GND_c_5_p N_noxref_4_c_909_n ) capacitor c=0.0126573f //x=14.43 \
 //y=0 //x2=15.24 //y2=1.915
cc_50 ( N_GND_M9_noxref_d N_noxref_4_c_910_n ) capacitor c=0.0131341f \
 //x=15.315 //y=0.875 //x2=15.615 //y2=0.72
cc_51 ( N_GND_M9_noxref_d N_noxref_4_c_911_n ) capacitor c=0.00193146f \
 //x=15.315 //y=0.875 //x2=15.615 //y2=1.375
cc_52 ( N_GND_c_52_p N_noxref_4_c_912_n ) capacitor c=0.00129018f //x=19.07 \
 //y=0 //x2=15.77 //y2=0.875
cc_53 ( N_GND_M9_noxref_d N_noxref_4_c_912_n ) capacitor c=0.00257848f \
 //x=15.315 //y=0.875 //x2=15.77 //y2=0.875
cc_54 ( N_GND_M9_noxref_d N_noxref_4_c_914_n ) capacitor c=0.00255985f \
 //x=15.315 //y=0.875 //x2=15.77 //y2=1.22
cc_55 ( N_GND_c_5_p N_noxref_4_M8_noxref_d ) capacitor c=0.00591582f //x=14.43 \
 //y=0 //x2=13.015 //y2=0.915
cc_56 ( N_GND_c_8_p N_CLK_c_1062_n ) capacitor c=0.0284311f //x=28.12 //y=0 \
 //x2=16.535 //y2=3.33
cc_57 ( N_GND_c_3_p N_CLK_c_1063_n ) capacitor c=7.64246e-19 //x=4.81 //y=0 \
 //x2=7.03 //y2=2.08
cc_58 ( N_GND_c_5_p N_CLK_c_1064_n ) capacitor c=6.4925e-19 //x=14.43 //y=0 \
 //x2=16.65 //y2=2.08
cc_59 ( N_GND_c_8_p N_noxref_6_c_1253_n ) capacitor c=0.00825249f //x=28.12 \
 //y=0 //x2=8.765 //y2=3.7
cc_60 ( N_GND_c_8_p N_noxref_6_c_1254_n ) capacitor c=0.00154647f //x=28.12 \
 //y=0 //x2=3.445 //y2=3.7
cc_61 ( N_GND_c_6_p N_noxref_6_c_1255_n ) capacitor c=0.0034979f //x=19.24 \
 //y=0 //x2=20.235 //y2=3.7
cc_62 ( N_GND_c_3_p N_noxref_6_c_1256_n ) capacitor c=9.53263e-19 //x=4.81 \
 //y=0 //x2=3.33 //y2=2.08
cc_63 ( N_GND_c_4_p N_noxref_6_c_1257_n ) capacitor c=0.0455868f //x=9.62 \
 //y=0 //x2=8.795 //y2=1.665
cc_64 ( N_GND_c_6_p N_noxref_6_c_1258_n ) capacitor c=0.0153336f //x=19.24 \
 //y=0 //x2=20.35 //y2=2.08
cc_65 ( N_GND_c_65_p N_noxref_6_c_1259_n ) capacitor c=0.00132755f //x=20.23 \
 //y=0 //x2=20.05 //y2=0.875
cc_66 ( N_GND_M12_noxref_d N_noxref_6_c_1259_n ) capacitor c=0.00211996f \
 //x=20.125 //y=0.875 //x2=20.05 //y2=0.875
cc_67 ( N_GND_M12_noxref_d N_noxref_6_c_1261_n ) capacitor c=0.00255985f \
 //x=20.125 //y=0.875 //x2=20.05 //y2=1.22
cc_68 ( N_GND_c_6_p N_noxref_6_c_1262_n ) capacitor c=0.00204716f //x=19.24 \
 //y=0 //x2=20.05 //y2=1.53
cc_69 ( N_GND_c_6_p N_noxref_6_c_1263_n ) capacitor c=0.0126573f //x=19.24 \
 //y=0 //x2=20.05 //y2=1.915
cc_70 ( N_GND_M12_noxref_d N_noxref_6_c_1264_n ) capacitor c=0.0131341f \
 //x=20.125 //y=0.875 //x2=20.425 //y2=0.72
cc_71 ( N_GND_M12_noxref_d N_noxref_6_c_1265_n ) capacitor c=0.00193146f \
 //x=20.125 //y=0.875 //x2=20.425 //y2=1.375
cc_72 ( N_GND_c_72_p N_noxref_6_c_1266_n ) capacitor c=0.00129018f //x=23.88 \
 //y=0 //x2=20.58 //y2=0.875
cc_73 ( N_GND_M12_noxref_d N_noxref_6_c_1266_n ) capacitor c=0.00257848f \
 //x=20.125 //y=0.875 //x2=20.58 //y2=0.875
cc_74 ( N_GND_M12_noxref_d N_noxref_6_c_1268_n ) capacitor c=0.00255985f \
 //x=20.125 //y=0.875 //x2=20.58 //y2=1.22
cc_75 ( N_GND_c_4_p N_noxref_6_M5_noxref_d ) capacitor c=0.00591582f //x=9.62 \
 //y=0 //x2=8.205 //y2=0.915
cc_76 ( N_GND_c_8_p N_RN_c_1514_n ) capacitor c=0.00571459f //x=28.12 //y=0 \
 //x2=17.645 //y2=4.44
cc_77 ( N_GND_c_8_p N_RN_c_1515_n ) capacitor c=0.00132659f //x=28.12 //y=0 \
 //x2=2.335 //y2=4.44
cc_78 ( N_GND_c_1_p N_RN_c_1516_n ) capacitor c=7.64246e-19 //x=0.74 //y=0 \
 //x2=2.22 //y2=2.08
cc_79 ( N_GND_c_6_p N_RN_c_1517_n ) capacitor c=7.09207e-19 //x=19.24 //y=0 \
 //x2=17.76 //y2=2.08
cc_80 ( N_GND_c_6_p N_RN_c_1518_n ) capacitor c=6.4925e-19 //x=19.24 //y=0 \
 //x2=21.46 //y2=2.08
cc_81 ( N_GND_c_7_p N_QN_c_1823_n ) capacitor c=0.00505527f //x=24.05 //y=0 \
 //x2=25.045 //y2=3.33
cc_82 ( N_GND_c_7_p N_QN_c_1824_n ) capacitor c=0.0432429f //x=24.05 //y=0 \
 //x2=23.225 //y2=1.665
cc_83 ( N_GND_c_7_p N_QN_c_1825_n ) capacitor c=0.0152529f //x=24.05 //y=0 \
 //x2=25.16 //y2=2.08
cc_84 ( N_GND_c_84_p N_QN_c_1826_n ) capacitor c=0.00132755f //x=25.04 //y=0 \
 //x2=24.86 //y2=0.875
cc_85 ( N_GND_M15_noxref_d N_QN_c_1826_n ) capacitor c=0.00211996f //x=24.935 \
 //y=0.875 //x2=24.86 //y2=0.875
cc_86 ( N_GND_M15_noxref_d N_QN_c_1828_n ) capacitor c=0.00255985f //x=24.935 \
 //y=0.875 //x2=24.86 //y2=1.22
cc_87 ( N_GND_c_7_p N_QN_c_1829_n ) capacitor c=0.00204716f //x=24.05 //y=0 \
 //x2=24.86 //y2=1.53
cc_88 ( N_GND_c_7_p N_QN_c_1830_n ) capacitor c=0.0126573f //x=24.05 //y=0 \
 //x2=24.86 //y2=1.915
cc_89 ( N_GND_M15_noxref_d N_QN_c_1831_n ) capacitor c=0.0131341f //x=24.935 \
 //y=0.875 //x2=25.235 //y2=0.72
cc_90 ( N_GND_M15_noxref_d N_QN_c_1832_n ) capacitor c=0.00193146f //x=24.935 \
 //y=0.875 //x2=25.235 //y2=1.375
cc_91 ( N_GND_c_2_p N_QN_c_1833_n ) capacitor c=0.00129018f //x=28.12 //y=0 \
 //x2=25.39 //y2=0.875
cc_92 ( N_GND_M15_noxref_d N_QN_c_1833_n ) capacitor c=0.00257848f //x=24.935 \
 //y=0.875 //x2=25.39 //y2=0.875
cc_93 ( N_GND_M15_noxref_d N_QN_c_1835_n ) capacitor c=0.00255985f //x=24.935 \
 //y=0.875 //x2=25.39 //y2=1.22
cc_94 ( N_GND_c_7_p N_QN_M14_noxref_d ) capacitor c=0.00591582f //x=24.05 \
 //y=0 //x2=22.635 //y2=0.915
cc_95 ( N_GND_c_8_p N_SN_c_1980_n ) capacitor c=0.120604f //x=28.12 //y=0 \
 //x2=26.155 //y2=2.59
cc_96 ( N_GND_c_38_p N_SN_c_1980_n ) capacitor c=0.00342161f //x=14.26 //y=0 \
 //x2=26.155 //y2=2.59
cc_97 ( N_GND_c_45_p N_SN_c_1980_n ) capacitor c=0.00221947f //x=15.42 //y=0 \
 //x2=26.155 //y2=2.59
cc_98 ( N_GND_c_52_p N_SN_c_1980_n ) capacitor c=0.00344363f //x=19.07 //y=0 \
 //x2=26.155 //y2=2.59
cc_99 ( N_GND_c_65_p N_SN_c_1980_n ) capacitor c=0.00221947f //x=20.23 //y=0 \
 //x2=26.155 //y2=2.59
cc_100 ( N_GND_c_72_p N_SN_c_1980_n ) capacitor c=0.00344363f //x=23.88 //y=0 \
 //x2=26.155 //y2=2.59
cc_101 ( N_GND_c_84_p N_SN_c_1980_n ) capacitor c=0.00221947f //x=25.04 //y=0 \
 //x2=26.155 //y2=2.59
cc_102 ( N_GND_c_5_p N_SN_c_1980_n ) capacitor c=0.0338055f //x=14.43 //y=0 \
 //x2=26.155 //y2=2.59
cc_103 ( N_GND_c_6_p N_SN_c_1980_n ) capacitor c=0.0377057f //x=19.24 //y=0 \
 //x2=26.155 //y2=2.59
cc_104 ( N_GND_c_7_p N_SN_c_1980_n ) capacitor c=0.0360747f //x=24.05 //y=0 \
 //x2=26.155 //y2=2.59
cc_105 ( N_GND_c_8_p N_SN_c_1990_n ) capacitor c=0.00219703f //x=28.12 //y=0 \
 //x2=11.955 //y2=2.59
cc_106 ( N_GND_c_4_p N_SN_c_1991_n ) capacitor c=9.22578e-19 //x=9.62 //y=0 \
 //x2=11.84 //y2=2.08
cc_107 ( N_GND_c_7_p N_SN_c_1992_n ) capacitor c=6.9062e-19 //x=24.05 //y=0 \
 //x2=26.27 //y2=2.08
cc_108 ( N_GND_c_4_p N_noxref_10_c_2209_n ) capacitor c=9.53263e-19 //x=9.62 \
 //y=0 //x2=8.14 //y2=2.08
cc_109 ( N_GND_c_5_p N_noxref_10_c_2210_n ) capacitor c=7.95208e-19 //x=14.43 \
 //y=0 //x2=12.95 //y2=2.08
cc_110 ( N_GND_c_6_p N_noxref_10_c_2211_n ) capacitor c=0.0433371f //x=19.24 \
 //y=0 //x2=18.415 //y2=1.665
cc_111 ( N_GND_c_2_p N_noxref_10_c_2212_n ) capacitor c=0.00128267f //x=28.12 \
 //y=0 //x2=27.38 //y2=2.08
cc_112 ( N_GND_c_6_p N_noxref_10_M11_noxref_d ) capacitor c=0.00591582f \
 //x=19.24 //y=0 //x2=17.825 //y2=0.915
cc_113 ( N_GND_c_8_p N_Q_c_2549_n ) capacitor c=0.0135088f //x=28.12 //y=0 \
 //x2=28.005 //y2=3.7
cc_114 ( N_GND_c_7_p N_Q_c_2550_n ) capacitor c=7.09207e-19 //x=24.05 //y=0 \
 //x2=22.57 //y2=2.08
cc_115 ( N_GND_c_2_p N_Q_c_2551_n ) capacitor c=0.0461865f //x=28.12 //y=0 \
 //x2=28.035 //y2=1.665
cc_116 ( N_GND_c_2_p N_Q_M17_noxref_d ) capacitor c=0.00593061f //x=28.12 \
 //y=0 //x2=27.445 //y2=0.915
cc_117 ( N_GND_c_1_p N_D_c_2706_n ) capacitor c=0.0180363f //x=0.74 //y=0 \
 //x2=1.11 //y2=2.08
cc_118 ( N_GND_c_118_p N_D_c_2707_n ) capacitor c=0.00132755f //x=0.99 //y=0 \
 //x2=0.81 //y2=0.875
cc_119 ( N_GND_M0_noxref_d N_D_c_2707_n ) capacitor c=0.00211996f //x=0.885 \
 //y=0.875 //x2=0.81 //y2=0.875
cc_120 ( N_GND_M0_noxref_d N_D_c_2709_n ) capacitor c=0.00255985f //x=0.885 \
 //y=0.875 //x2=0.81 //y2=1.22
cc_121 ( N_GND_c_1_p N_D_c_2710_n ) capacitor c=0.00295461f //x=0.74 //y=0 \
 //x2=0.81 //y2=1.53
cc_122 ( N_GND_c_1_p N_D_c_2711_n ) capacitor c=0.0134214f //x=0.74 //y=0 \
 //x2=0.81 //y2=1.915
cc_123 ( N_GND_M0_noxref_d N_D_c_2712_n ) capacitor c=0.0131341f //x=0.885 \
 //y=0.875 //x2=1.185 //y2=0.72
cc_124 ( N_GND_M0_noxref_d N_D_c_2713_n ) capacitor c=0.00193146f //x=0.885 \
 //y=0.875 //x2=1.185 //y2=1.375
cc_125 ( N_GND_c_9_p N_D_c_2714_n ) capacitor c=0.00129018f //x=4.64 //y=0 \
 //x2=1.34 //y2=0.875
cc_126 ( N_GND_M0_noxref_d N_D_c_2714_n ) capacitor c=0.00257848f //x=0.885 \
 //y=0.875 //x2=1.34 //y2=0.875
cc_127 ( N_GND_M0_noxref_d N_D_c_2716_n ) capacitor c=0.00255985f //x=0.885 \
 //y=0.875 //x2=1.34 //y2=1.22
cc_128 ( N_GND_c_8_p N_noxref_13_c_2762_n ) capacitor c=0.00710541f //x=28.12 \
 //y=0 //x2=1.475 //y2=1.59
cc_129 ( N_GND_c_118_p N_noxref_13_c_2762_n ) capacitor c=0.00110021f //x=0.99 \
 //y=0 //x2=1.475 //y2=1.59
cc_130 ( N_GND_c_9_p N_noxref_13_c_2762_n ) capacitor c=0.00179185f //x=4.64 \
 //y=0 //x2=1.475 //y2=1.59
cc_131 ( N_GND_M0_noxref_d N_noxref_13_c_2762_n ) capacitor c=0.00900091f \
 //x=0.885 //y=0.875 //x2=1.475 //y2=1.59
cc_132 ( N_GND_c_8_p N_noxref_13_c_2766_n ) capacitor c=0.00709506f //x=28.12 \
 //y=0 //x2=1.56 //y2=0.625
cc_133 ( N_GND_c_9_p N_noxref_13_c_2766_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=1.56 //y2=0.625
cc_134 ( N_GND_M0_noxref_d N_noxref_13_c_2766_n ) capacitor c=0.033954f \
 //x=0.885 //y=0.875 //x2=1.56 //y2=0.625
cc_135 ( N_GND_c_8_p N_noxref_13_c_2769_n ) capacitor c=0.0169144f //x=28.12 \
 //y=0 //x2=2.445 //y2=0.54
cc_136 ( N_GND_c_9_p N_noxref_13_c_2769_n ) capacitor c=0.0356078f //x=4.64 \
 //y=0 //x2=2.445 //y2=0.54
cc_137 ( N_GND_c_2_p N_noxref_13_c_2769_n ) capacitor c=0.00265129f //x=28.12 \
 //y=0 //x2=2.445 //y2=0.54
cc_138 ( N_GND_c_8_p N_noxref_13_M0_noxref_s ) capacitor c=0.0126182f \
 //x=28.12 //y=0 //x2=0.455 //y2=0.375
cc_139 ( N_GND_c_118_p N_noxref_13_M0_noxref_s ) capacitor c=0.0140218f \
 //x=0.99 //y=0 //x2=0.455 //y2=0.375
cc_140 ( N_GND_c_1_p N_noxref_13_M0_noxref_s ) capacitor c=0.0712607f //x=0.74 \
 //y=0 //x2=0.455 //y2=0.375
cc_141 ( N_GND_c_9_p N_noxref_13_M0_noxref_s ) capacitor c=0.0131422f //x=4.64 \
 //y=0 //x2=0.455 //y2=0.375
cc_142 ( N_GND_c_3_p N_noxref_13_M0_noxref_s ) capacitor c=3.31601e-19 \
 //x=4.81 //y=0 //x2=0.455 //y2=0.375
cc_143 ( N_GND_M0_noxref_d N_noxref_13_M0_noxref_s ) capacitor c=0.033718f \
 //x=0.885 //y=0.875 //x2=0.455 //y2=0.375
cc_144 ( N_GND_c_8_p N_noxref_14_c_2808_n ) capacitor c=0.00667057f //x=28.12 \
 //y=0 //x2=3.015 //y2=0.995
cc_145 ( N_GND_c_9_p N_noxref_14_c_2808_n ) capacitor c=0.00829979f //x=4.64 \
 //y=0 //x2=3.015 //y2=0.995
cc_146 ( N_GND_c_2_p N_noxref_14_c_2808_n ) capacitor c=3.54249e-19 //x=28.12 \
 //y=0 //x2=3.015 //y2=0.995
cc_147 ( N_GND_c_8_p N_noxref_14_c_2811_n ) capacitor c=0.00583375f //x=28.12 \
 //y=0 //x2=3.1 //y2=0.625
cc_148 ( N_GND_c_9_p N_noxref_14_c_2811_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=3.1 //y2=0.625
cc_149 ( N_GND_M0_noxref_d N_noxref_14_c_2811_n ) capacitor c=6.21394e-19 \
 //x=0.885 //y=0.875 //x2=3.1 //y2=0.625
cc_150 ( N_GND_c_8_p N_noxref_14_c_2814_n ) capacitor c=0.0121495f //x=28.12 \
 //y=0 //x2=3.985 //y2=0.54
cc_151 ( N_GND_c_9_p N_noxref_14_c_2814_n ) capacitor c=0.0362581f //x=4.64 \
 //y=0 //x2=3.985 //y2=0.54
cc_152 ( N_GND_c_2_p N_noxref_14_c_2814_n ) capacitor c=0.00283214f //x=28.12 \
 //y=0 //x2=3.985 //y2=0.54
cc_153 ( N_GND_c_8_p N_noxref_14_c_2817_n ) capacitor c=0.00276729f //x=28.12 \
 //y=0 //x2=4.07 //y2=0.625
cc_154 ( N_GND_c_9_p N_noxref_14_c_2817_n ) capacitor c=0.0141921f //x=4.64 \
 //y=0 //x2=4.07 //y2=0.625
cc_155 ( N_GND_c_3_p N_noxref_14_c_2817_n ) capacitor c=0.0404137f //x=4.81 \
 //y=0 //x2=4.07 //y2=0.625
cc_156 ( N_GND_M0_noxref_d N_noxref_14_M1_noxref_d ) capacitor c=0.00162435f \
 //x=0.885 //y=0.875 //x2=1.86 //y2=0.91
cc_157 ( N_GND_c_1_p N_noxref_14_M2_noxref_s ) capacitor c=8.16352e-19 \
 //x=0.74 //y=0 //x2=2.965 //y2=0.375
cc_158 ( N_GND_c_3_p N_noxref_14_M2_noxref_s ) capacitor c=0.00183204f \
 //x=4.81 //y=0 //x2=2.965 //y2=0.375
cc_159 ( N_GND_c_8_p N_noxref_15_c_2861_n ) capacitor c=0.00540769f //x=28.12 \
 //y=0 //x2=6.285 //y2=1.59
cc_160 ( N_GND_c_10_p N_noxref_15_c_2861_n ) capacitor c=0.00111539f //x=5.8 \
 //y=0 //x2=6.285 //y2=1.59
cc_161 ( N_GND_c_14_p N_noxref_15_c_2861_n ) capacitor c=0.00180703f //x=9.45 \
 //y=0 //x2=6.285 //y2=1.59
cc_162 ( N_GND_M3_noxref_d N_noxref_15_c_2861_n ) capacitor c=0.00879948f \
 //x=5.695 //y=0.875 //x2=6.285 //y2=1.59
cc_163 ( N_GND_c_8_p N_noxref_15_c_2865_n ) capacitor c=0.00277721f //x=28.12 \
 //y=0 //x2=6.37 //y2=0.625
cc_164 ( N_GND_c_14_p N_noxref_15_c_2865_n ) capacitor c=0.0142595f //x=9.45 \
 //y=0 //x2=6.37 //y2=0.625
cc_165 ( N_GND_M3_noxref_d N_noxref_15_c_2865_n ) capacitor c=0.033954f \
 //x=5.695 //y=0.875 //x2=6.37 //y2=0.625
cc_166 ( N_GND_c_8_p N_noxref_15_c_2868_n ) capacitor c=0.0113743f //x=28.12 \
 //y=0 //x2=7.255 //y2=0.54
cc_167 ( N_GND_c_14_p N_noxref_15_c_2868_n ) capacitor c=0.0361685f //x=9.45 \
 //y=0 //x2=7.255 //y2=0.54
cc_168 ( N_GND_c_2_p N_noxref_15_c_2868_n ) capacitor c=0.00265129f //x=28.12 \
 //y=0 //x2=7.255 //y2=0.54
cc_169 ( N_GND_c_8_p N_noxref_15_M3_noxref_s ) capacitor c=0.00554931f \
 //x=28.12 //y=0 //x2=5.265 //y2=0.375
cc_170 ( N_GND_c_10_p N_noxref_15_M3_noxref_s ) capacitor c=0.0142595f //x=5.8 \
 //y=0 //x2=5.265 //y2=0.375
cc_171 ( N_GND_c_14_p N_noxref_15_M3_noxref_s ) capacitor c=0.0138379f \
 //x=9.45 //y=0 //x2=5.265 //y2=0.375
cc_172 ( N_GND_c_3_p N_noxref_15_M3_noxref_s ) capacitor c=0.0696963f //x=4.81 \
 //y=0 //x2=5.265 //y2=0.375
cc_173 ( N_GND_c_4_p N_noxref_15_M3_noxref_s ) capacitor c=3.31601e-19 \
 //x=9.62 //y=0 //x2=5.265 //y2=0.375
cc_174 ( N_GND_M3_noxref_d N_noxref_15_M3_noxref_s ) capacitor c=0.033718f \
 //x=5.695 //y=0.875 //x2=5.265 //y2=0.375
cc_175 ( N_GND_c_8_p N_noxref_16_c_2913_n ) capacitor c=0.00375578f //x=28.12 \
 //y=0 //x2=7.825 //y2=0.995
cc_176 ( N_GND_c_14_p N_noxref_16_c_2913_n ) capacitor c=0.00944923f //x=9.45 \
 //y=0 //x2=7.825 //y2=0.995
cc_177 ( N_GND_c_2_p N_noxref_16_c_2913_n ) capacitor c=3.54249e-19 //x=28.12 \
 //y=0 //x2=7.825 //y2=0.995
cc_178 ( N_GND_c_8_p N_noxref_16_c_2916_n ) capacitor c=0.00277721f //x=28.12 \
 //y=0 //x2=7.91 //y2=0.625
cc_179 ( N_GND_c_14_p N_noxref_16_c_2916_n ) capacitor c=0.0142595f //x=9.45 \
 //y=0 //x2=7.91 //y2=0.625
cc_180 ( N_GND_M3_noxref_d N_noxref_16_c_2916_n ) capacitor c=6.21394e-19 \
 //x=5.695 //y=0.875 //x2=7.91 //y2=0.625
cc_181 ( N_GND_c_8_p N_noxref_16_c_2919_n ) capacitor c=0.0114539f //x=28.12 \
 //y=0 //x2=8.795 //y2=0.54
cc_182 ( N_GND_c_14_p N_noxref_16_c_2919_n ) capacitor c=0.0365594f //x=9.45 \
 //y=0 //x2=8.795 //y2=0.54
cc_183 ( N_GND_c_2_p N_noxref_16_c_2919_n ) capacitor c=0.00283214f //x=28.12 \
 //y=0 //x2=8.795 //y2=0.54
cc_184 ( N_GND_c_8_p N_noxref_16_c_2922_n ) capacitor c=0.00277585f //x=28.12 \
 //y=0 //x2=8.88 //y2=0.625
cc_185 ( N_GND_c_14_p N_noxref_16_c_2922_n ) capacitor c=0.014198f //x=9.45 \
 //y=0 //x2=8.88 //y2=0.625
cc_186 ( N_GND_c_4_p N_noxref_16_c_2922_n ) capacitor c=0.0404137f //x=9.62 \
 //y=0 //x2=8.88 //y2=0.625
cc_187 ( N_GND_M3_noxref_d N_noxref_16_M4_noxref_d ) capacitor c=0.00162435f \
 //x=5.695 //y=0.875 //x2=6.67 //y2=0.91
cc_188 ( N_GND_c_3_p N_noxref_16_M5_noxref_s ) capacitor c=8.16352e-19 \
 //x=4.81 //y=0 //x2=7.775 //y2=0.375
cc_189 ( N_GND_c_4_p N_noxref_16_M5_noxref_s ) capacitor c=0.00183204f \
 //x=9.62 //y=0 //x2=7.775 //y2=0.375
cc_190 ( N_GND_c_8_p N_noxref_17_c_2967_n ) capacitor c=0.00543225f //x=28.12 \
 //y=0 //x2=11.095 //y2=1.59
cc_191 ( N_GND_c_15_p N_noxref_17_c_2967_n ) capacitor c=0.00111539f //x=10.61 \
 //y=0 //x2=11.095 //y2=1.59
cc_192 ( N_GND_c_38_p N_noxref_17_c_2967_n ) capacitor c=0.0018074f //x=14.26 \
 //y=0 //x2=11.095 //y2=1.59
cc_193 ( N_GND_M6_noxref_d N_noxref_17_c_2967_n ) capacitor c=0.00879948f \
 //x=10.505 //y=0.875 //x2=11.095 //y2=1.59
cc_194 ( N_GND_c_8_p N_noxref_17_c_2971_n ) capacitor c=0.00287639f //x=28.12 \
 //y=0 //x2=11.18 //y2=0.625
cc_195 ( N_GND_c_38_p N_noxref_17_c_2971_n ) capacitor c=0.014327f //x=14.26 \
 //y=0 //x2=11.18 //y2=0.625
cc_196 ( N_GND_M6_noxref_d N_noxref_17_c_2971_n ) capacitor c=0.033954f \
 //x=10.505 //y=0.875 //x2=11.18 //y2=0.625
cc_197 ( N_GND_c_8_p N_noxref_17_c_2974_n ) capacitor c=0.0113713f //x=28.12 \
 //y=0 //x2=12.065 //y2=0.54
cc_198 ( N_GND_c_38_p N_noxref_17_c_2974_n ) capacitor c=0.0361671f //x=14.26 \
 //y=0 //x2=12.065 //y2=0.54
cc_199 ( N_GND_c_2_p N_noxref_17_c_2974_n ) capacitor c=0.00265129f //x=28.12 \
 //y=0 //x2=12.065 //y2=0.54
cc_200 ( N_GND_c_8_p N_noxref_17_M6_noxref_s ) capacitor c=0.00543443f \
 //x=28.12 //y=0 //x2=10.075 //y2=0.375
cc_201 ( N_GND_c_15_p N_noxref_17_M6_noxref_s ) capacitor c=0.0142595f \
 //x=10.61 //y=0 //x2=10.075 //y2=0.375
cc_202 ( N_GND_c_38_p N_noxref_17_M6_noxref_s ) capacitor c=0.0137569f \
 //x=14.26 //y=0 //x2=10.075 //y2=0.375
cc_203 ( N_GND_c_4_p N_noxref_17_M6_noxref_s ) capacitor c=0.0696963f //x=9.62 \
 //y=0 //x2=10.075 //y2=0.375
cc_204 ( N_GND_c_5_p N_noxref_17_M6_noxref_s ) capacitor c=3.31601e-19 \
 //x=14.43 //y=0 //x2=10.075 //y2=0.375
cc_205 ( N_GND_M6_noxref_d N_noxref_17_M6_noxref_s ) capacitor c=0.033718f \
 //x=10.505 //y=0.875 //x2=10.075 //y2=0.375
cc_206 ( N_GND_c_8_p N_noxref_18_c_3021_n ) capacitor c=0.00364762f //x=28.12 \
 //y=0 //x2=12.635 //y2=0.995
cc_207 ( N_GND_c_38_p N_noxref_18_c_3021_n ) capacitor c=0.00940048f //x=14.26 \
 //y=0 //x2=12.635 //y2=0.995
cc_208 ( N_GND_c_2_p N_noxref_18_c_3021_n ) capacitor c=3.54249e-19 //x=28.12 \
 //y=0 //x2=12.635 //y2=0.995
cc_209 ( N_GND_c_8_p N_noxref_18_c_3024_n ) capacitor c=0.00266608f //x=28.12 \
 //y=0 //x2=12.72 //y2=0.625
cc_210 ( N_GND_c_38_p N_noxref_18_c_3024_n ) capacitor c=0.0141814f //x=14.26 \
 //y=0 //x2=12.72 //y2=0.625
cc_211 ( N_GND_M6_noxref_d N_noxref_18_c_3024_n ) capacitor c=6.21394e-19 \
 //x=10.505 //y=0.875 //x2=12.72 //y2=0.625
cc_212 ( N_GND_c_8_p N_noxref_18_c_3027_n ) capacitor c=0.0110123f //x=28.12 \
 //y=0 //x2=13.605 //y2=0.54
cc_213 ( N_GND_c_38_p N_noxref_18_c_3027_n ) capacitor c=0.0364696f //x=14.26 \
 //y=0 //x2=13.605 //y2=0.54
cc_214 ( N_GND_c_2_p N_noxref_18_c_3027_n ) capacitor c=0.00283214f //x=28.12 \
 //y=0 //x2=13.605 //y2=0.54
cc_215 ( N_GND_c_8_p N_noxref_18_c_3030_n ) capacitor c=0.00266421f //x=28.12 \
 //y=0 //x2=13.69 //y2=0.625
cc_216 ( N_GND_c_38_p N_noxref_18_c_3030_n ) capacitor c=0.0141195f //x=14.26 \
 //y=0 //x2=13.69 //y2=0.625
cc_217 ( N_GND_c_5_p N_noxref_18_c_3030_n ) capacitor c=0.0404137f //x=14.43 \
 //y=0 //x2=13.69 //y2=0.625
cc_218 ( N_GND_M6_noxref_d N_noxref_18_M7_noxref_d ) capacitor c=0.00162435f \
 //x=10.505 //y=0.875 //x2=11.48 //y2=0.91
cc_219 ( N_GND_c_4_p N_noxref_18_M8_noxref_s ) capacitor c=8.16352e-19 \
 //x=9.62 //y=0 //x2=12.585 //y2=0.375
cc_220 ( N_GND_c_5_p N_noxref_18_M8_noxref_s ) capacitor c=0.00183204f \
 //x=14.43 //y=0 //x2=12.585 //y2=0.375
cc_221 ( N_GND_c_8_p N_noxref_19_c_3075_n ) capacitor c=0.00529827f //x=28.12 \
 //y=0 //x2=15.905 //y2=1.59
cc_222 ( N_GND_c_45_p N_noxref_19_c_3075_n ) capacitor c=0.00111496f //x=15.42 \
 //y=0 //x2=15.905 //y2=1.59
cc_223 ( N_GND_c_52_p N_noxref_19_c_3075_n ) capacitor c=0.0018066f //x=19.07 \
 //y=0 //x2=15.905 //y2=1.59
cc_224 ( N_GND_M9_noxref_d N_noxref_19_c_3075_n ) capacitor c=0.00869643f \
 //x=15.315 //y=0.875 //x2=15.905 //y2=1.59
cc_225 ( N_GND_c_8_p N_noxref_19_c_3079_n ) capacitor c=0.00266608f //x=28.12 \
 //y=0 //x2=15.99 //y2=0.625
cc_226 ( N_GND_c_52_p N_noxref_19_c_3079_n ) capacitor c=0.0141814f //x=19.07 \
 //y=0 //x2=15.99 //y2=0.625
cc_227 ( N_GND_M9_noxref_d N_noxref_19_c_3079_n ) capacitor c=0.033954f \
 //x=15.315 //y=0.875 //x2=15.99 //y2=0.625
cc_228 ( N_GND_c_8_p N_noxref_19_c_3082_n ) capacitor c=0.0109327f //x=28.12 \
 //y=0 //x2=16.875 //y2=0.54
cc_229 ( N_GND_c_52_p N_noxref_19_c_3082_n ) capacitor c=0.0361235f //x=19.07 \
 //y=0 //x2=16.875 //y2=0.54
cc_230 ( N_GND_c_2_p N_noxref_19_c_3082_n ) capacitor c=0.00265129f //x=28.12 \
 //y=0 //x2=16.875 //y2=0.54
cc_231 ( N_GND_c_8_p N_noxref_19_M9_noxref_s ) capacitor c=0.00532331f \
 //x=28.12 //y=0 //x2=14.885 //y2=0.375
cc_232 ( N_GND_c_45_p N_noxref_19_M9_noxref_s ) capacitor c=0.0141814f \
 //x=15.42 //y=0 //x2=14.885 //y2=0.375
cc_233 ( N_GND_c_52_p N_noxref_19_M9_noxref_s ) capacitor c=0.0132355f \
 //x=19.07 //y=0 //x2=14.885 //y2=0.375
cc_234 ( N_GND_c_5_p N_noxref_19_M9_noxref_s ) capacitor c=0.0696963f \
 //x=14.43 //y=0 //x2=14.885 //y2=0.375
cc_235 ( N_GND_c_6_p N_noxref_19_M9_noxref_s ) capacitor c=3.31601e-19 \
 //x=19.24 //y=0 //x2=14.885 //y2=0.375
cc_236 ( N_GND_M9_noxref_d N_noxref_19_M9_noxref_s ) capacitor c=0.033718f \
 //x=15.315 //y=0.875 //x2=14.885 //y2=0.375
cc_237 ( N_GND_c_8_p N_noxref_20_c_3125_n ) capacitor c=0.00364762f //x=28.12 \
 //y=0 //x2=17.445 //y2=0.995
cc_238 ( N_GND_c_52_p N_noxref_20_c_3125_n ) capacitor c=0.00940048f //x=19.07 \
 //y=0 //x2=17.445 //y2=0.995
cc_239 ( N_GND_c_2_p N_noxref_20_c_3125_n ) capacitor c=3.54249e-19 //x=28.12 \
 //y=0 //x2=17.445 //y2=0.995
cc_240 ( N_GND_c_8_p N_noxref_20_c_3128_n ) capacitor c=0.00266608f //x=28.12 \
 //y=0 //x2=17.53 //y2=0.625
cc_241 ( N_GND_c_52_p N_noxref_20_c_3128_n ) capacitor c=0.0141814f //x=19.07 \
 //y=0 //x2=17.53 //y2=0.625
cc_242 ( N_GND_M9_noxref_d N_noxref_20_c_3128_n ) capacitor c=6.21394e-19 \
 //x=15.315 //y=0.875 //x2=17.53 //y2=0.625
cc_243 ( N_GND_c_8_p N_noxref_20_c_3131_n ) capacitor c=0.0110123f //x=28.12 \
 //y=0 //x2=18.415 //y2=0.54
cc_244 ( N_GND_c_52_p N_noxref_20_c_3131_n ) capacitor c=0.0365163f //x=19.07 \
 //y=0 //x2=18.415 //y2=0.54
cc_245 ( N_GND_c_2_p N_noxref_20_c_3131_n ) capacitor c=0.00283214f //x=28.12 \
 //y=0 //x2=18.415 //y2=0.54
cc_246 ( N_GND_c_8_p N_noxref_20_c_3134_n ) capacitor c=0.00266421f //x=28.12 \
 //y=0 //x2=18.5 //y2=0.625
cc_247 ( N_GND_c_52_p N_noxref_20_c_3134_n ) capacitor c=0.0141195f //x=19.07 \
 //y=0 //x2=18.5 //y2=0.625
cc_248 ( N_GND_c_6_p N_noxref_20_c_3134_n ) capacitor c=0.0404137f //x=19.24 \
 //y=0 //x2=18.5 //y2=0.625
cc_249 ( N_GND_M9_noxref_d N_noxref_20_M10_noxref_d ) capacitor c=0.00162435f \
 //x=15.315 //y=0.875 //x2=16.29 //y2=0.91
cc_250 ( N_GND_c_5_p N_noxref_20_M11_noxref_s ) capacitor c=8.16352e-19 \
 //x=14.43 //y=0 //x2=17.395 //y2=0.375
cc_251 ( N_GND_c_6_p N_noxref_20_M11_noxref_s ) capacitor c=0.00183204f \
 //x=19.24 //y=0 //x2=17.395 //y2=0.375
cc_252 ( N_GND_c_8_p N_noxref_21_c_3179_n ) capacitor c=0.00529827f //x=28.12 \
 //y=0 //x2=20.715 //y2=1.59
cc_253 ( N_GND_c_65_p N_noxref_21_c_3179_n ) capacitor c=0.00111496f //x=20.23 \
 //y=0 //x2=20.715 //y2=1.59
cc_254 ( N_GND_c_72_p N_noxref_21_c_3179_n ) capacitor c=0.0018066f //x=23.88 \
 //y=0 //x2=20.715 //y2=1.59
cc_255 ( N_GND_M12_noxref_d N_noxref_21_c_3179_n ) capacitor c=0.00869643f \
 //x=20.125 //y=0.875 //x2=20.715 //y2=1.59
cc_256 ( N_GND_c_8_p N_noxref_21_c_3183_n ) capacitor c=0.00266608f //x=28.12 \
 //y=0 //x2=20.8 //y2=0.625
cc_257 ( N_GND_c_72_p N_noxref_21_c_3183_n ) capacitor c=0.0141814f //x=23.88 \
 //y=0 //x2=20.8 //y2=0.625
cc_258 ( N_GND_M12_noxref_d N_noxref_21_c_3183_n ) capacitor c=0.033954f \
 //x=20.125 //y=0.875 //x2=20.8 //y2=0.625
cc_259 ( N_GND_c_8_p N_noxref_21_c_3186_n ) capacitor c=0.0109327f //x=28.12 \
 //y=0 //x2=21.685 //y2=0.54
cc_260 ( N_GND_c_72_p N_noxref_21_c_3186_n ) capacitor c=0.0361235f //x=23.88 \
 //y=0 //x2=21.685 //y2=0.54
cc_261 ( N_GND_c_2_p N_noxref_21_c_3186_n ) capacitor c=0.00265129f //x=28.12 \
 //y=0 //x2=21.685 //y2=0.54
cc_262 ( N_GND_c_8_p N_noxref_21_M12_noxref_s ) capacitor c=0.00532331f \
 //x=28.12 //y=0 //x2=19.695 //y2=0.375
cc_263 ( N_GND_c_65_p N_noxref_21_M12_noxref_s ) capacitor c=0.0141814f \
 //x=20.23 //y=0 //x2=19.695 //y2=0.375
cc_264 ( N_GND_c_72_p N_noxref_21_M12_noxref_s ) capacitor c=0.0132355f \
 //x=23.88 //y=0 //x2=19.695 //y2=0.375
cc_265 ( N_GND_c_6_p N_noxref_21_M12_noxref_s ) capacitor c=0.0696963f \
 //x=19.24 //y=0 //x2=19.695 //y2=0.375
cc_266 ( N_GND_c_7_p N_noxref_21_M12_noxref_s ) capacitor c=3.31601e-19 \
 //x=24.05 //y=0 //x2=19.695 //y2=0.375
cc_267 ( N_GND_M12_noxref_d N_noxref_21_M12_noxref_s ) capacitor c=0.033718f \
 //x=20.125 //y=0.875 //x2=19.695 //y2=0.375
cc_268 ( N_GND_c_8_p N_noxref_22_c_3229_n ) capacitor c=0.00364762f //x=28.12 \
 //y=0 //x2=22.255 //y2=0.995
cc_269 ( N_GND_c_72_p N_noxref_22_c_3229_n ) capacitor c=0.00940048f //x=23.88 \
 //y=0 //x2=22.255 //y2=0.995
cc_270 ( N_GND_c_2_p N_noxref_22_c_3229_n ) capacitor c=3.54249e-19 //x=28.12 \
 //y=0 //x2=22.255 //y2=0.995
cc_271 ( N_GND_c_8_p N_noxref_22_c_3232_n ) capacitor c=0.00266608f //x=28.12 \
 //y=0 //x2=22.34 //y2=0.625
cc_272 ( N_GND_c_72_p N_noxref_22_c_3232_n ) capacitor c=0.0141814f //x=23.88 \
 //y=0 //x2=22.34 //y2=0.625
cc_273 ( N_GND_M12_noxref_d N_noxref_22_c_3232_n ) capacitor c=6.21394e-19 \
 //x=20.125 //y=0.875 //x2=22.34 //y2=0.625
cc_274 ( N_GND_c_8_p N_noxref_22_c_3235_n ) capacitor c=0.0110123f //x=28.12 \
 //y=0 //x2=23.225 //y2=0.54
cc_275 ( N_GND_c_72_p N_noxref_22_c_3235_n ) capacitor c=0.0364696f //x=23.88 \
 //y=0 //x2=23.225 //y2=0.54
cc_276 ( N_GND_c_2_p N_noxref_22_c_3235_n ) capacitor c=0.00283214f //x=28.12 \
 //y=0 //x2=23.225 //y2=0.54
cc_277 ( N_GND_c_8_p N_noxref_22_c_3238_n ) capacitor c=0.00266421f //x=28.12 \
 //y=0 //x2=23.31 //y2=0.625
cc_278 ( N_GND_c_72_p N_noxref_22_c_3238_n ) capacitor c=0.0141195f //x=23.88 \
 //y=0 //x2=23.31 //y2=0.625
cc_279 ( N_GND_c_7_p N_noxref_22_c_3238_n ) capacitor c=0.0404137f //x=24.05 \
 //y=0 //x2=23.31 //y2=0.625
cc_280 ( N_GND_M12_noxref_d N_noxref_22_M13_noxref_d ) capacitor c=0.00162435f \
 //x=20.125 //y=0.875 //x2=21.1 //y2=0.91
cc_281 ( N_GND_c_6_p N_noxref_22_M14_noxref_s ) capacitor c=8.16352e-19 \
 //x=19.24 //y=0 //x2=22.205 //y2=0.375
cc_282 ( N_GND_c_7_p N_noxref_22_M14_noxref_s ) capacitor c=0.00183204f \
 //x=24.05 //y=0 //x2=22.205 //y2=0.375
cc_283 ( N_GND_c_8_p N_noxref_23_c_3283_n ) capacitor c=0.00529827f //x=28.12 \
 //y=0 //x2=25.525 //y2=1.59
cc_284 ( N_GND_c_84_p N_noxref_23_c_3283_n ) capacitor c=0.00111496f //x=25.04 \
 //y=0 //x2=25.525 //y2=1.59
cc_285 ( N_GND_c_2_p N_noxref_23_c_3283_n ) capacitor c=0.0018066f //x=28.12 \
 //y=0 //x2=25.525 //y2=1.59
cc_286 ( N_GND_M15_noxref_d N_noxref_23_c_3283_n ) capacitor c=0.00869643f \
 //x=24.935 //y=0.875 //x2=25.525 //y2=1.59
cc_287 ( N_GND_c_8_p N_noxref_23_c_3287_n ) capacitor c=0.00266608f //x=28.12 \
 //y=0 //x2=25.61 //y2=0.625
cc_288 ( N_GND_c_2_p N_noxref_23_c_3287_n ) capacitor c=0.0141814f //x=28.12 \
 //y=0 //x2=25.61 //y2=0.625
cc_289 ( N_GND_M15_noxref_d N_noxref_23_c_3287_n ) capacitor c=0.033954f \
 //x=24.935 //y=0.875 //x2=25.61 //y2=0.625
cc_290 ( N_GND_c_8_p N_noxref_23_c_3290_n ) capacitor c=0.0110426f //x=28.12 \
 //y=0 //x2=26.495 //y2=0.54
cc_291 ( N_GND_c_2_p N_noxref_23_c_3290_n ) capacitor c=0.0385273f //x=28.12 \
 //y=0 //x2=26.495 //y2=0.54
cc_292 ( N_GND_c_8_p N_noxref_23_M15_noxref_s ) capacitor c=0.00563707f \
 //x=28.12 //y=0 //x2=24.505 //y2=0.375
cc_293 ( N_GND_c_84_p N_noxref_23_M15_noxref_s ) capacitor c=0.0141814f \
 //x=25.04 //y=0 //x2=24.505 //y2=0.375
cc_294 ( N_GND_c_2_p N_noxref_23_M15_noxref_s ) capacitor c=0.0129524f \
 //x=28.12 //y=0 //x2=24.505 //y2=0.375
cc_295 ( N_GND_c_7_p N_noxref_23_M15_noxref_s ) capacitor c=0.0696963f \
 //x=24.05 //y=0 //x2=24.505 //y2=0.375
cc_296 ( N_GND_M15_noxref_d N_noxref_23_M15_noxref_s ) capacitor c=0.033718f \
 //x=24.935 //y=0.875 //x2=24.505 //y2=0.375
cc_297 ( N_GND_c_8_p N_noxref_24_c_3333_n ) capacitor c=0.00394306f //x=28.12 \
 //y=0 //x2=27.065 //y2=0.995
cc_298 ( N_GND_c_2_p N_noxref_24_c_3333_n ) capacitor c=0.00865404f //x=28.12 \
 //y=0 //x2=27.065 //y2=0.995
cc_299 ( N_GND_c_8_p N_noxref_24_c_3335_n ) capacitor c=0.00296961f //x=28.12 \
 //y=0 //x2=27.15 //y2=0.625
cc_300 ( N_GND_c_2_p N_noxref_24_c_3335_n ) capacitor c=0.0140218f //x=28.12 \
 //y=0 //x2=27.15 //y2=0.625
cc_301 ( N_GND_M15_noxref_d N_noxref_24_c_3335_n ) capacitor c=6.21394e-19 \
 //x=24.935 //y=0.875 //x2=27.15 //y2=0.625
cc_302 ( N_GND_c_8_p N_noxref_24_c_3338_n ) capacitor c=0.0122137f //x=28.12 \
 //y=0 //x2=28.035 //y2=0.54
cc_303 ( N_GND_c_2_p N_noxref_24_c_3338_n ) capacitor c=0.0388692f //x=28.12 \
 //y=0 //x2=28.035 //y2=0.54
cc_304 ( N_GND_c_8_p N_noxref_24_c_3340_n ) capacitor c=0.00296179f //x=28.12 \
 //y=0 //x2=28.12 //y2=0.625
cc_305 ( N_GND_c_2_p N_noxref_24_c_3340_n ) capacitor c=0.0549101f //x=28.12 \
 //y=0 //x2=28.12 //y2=0.625
cc_306 ( N_GND_M15_noxref_d N_noxref_24_M16_noxref_d ) capacitor c=0.00162435f \
 //x=24.935 //y=0.875 //x2=25.91 //y2=0.91
cc_307 ( N_GND_c_2_p N_noxref_24_M17_noxref_s ) capacitor c=0.00183576f \
 //x=28.12 //y=0 //x2=27.015 //y2=0.375
cc_308 ( N_GND_c_7_p N_noxref_24_M17_noxref_s ) capacitor c=8.16352e-19 \
 //x=24.05 //y=0 //x2=27.015 //y2=0.375
cc_309 ( N_VDD_c_316_p N_noxref_3_c_685_n ) capacitor c=0.00557756f //x=28.12 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_310 ( N_VDD_c_317_p N_noxref_3_c_685_n ) capacitor c=4.18223e-19 //x=1.885 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_311 ( N_VDD_c_318_p N_noxref_3_c_685_n ) capacitor c=4.31906e-19 //x=2.765 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_312 ( N_VDD_M19_noxref_d N_noxref_3_c_685_n ) capacitor c=0.0119114f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_313 ( N_VDD_c_309_n N_noxref_3_c_689_n ) capacitor c=0.00880189f //x=0.74 \
 //y=7.4 //x2=1.615 //y2=5.155
cc_314 ( N_VDD_M18_noxref_s N_noxref_3_c_689_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_315 ( N_VDD_c_316_p N_noxref_3_c_691_n ) capacitor c=0.0044221f //x=28.12 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_316 ( N_VDD_c_318_p N_noxref_3_c_691_n ) capacitor c=4.31931e-19 //x=2.765 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_317 ( N_VDD_c_324_p N_noxref_3_c_691_n ) capacitor c=4.31931e-19 //x=3.645 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_318 ( N_VDD_M21_noxref_d N_noxref_3_c_691_n ) capacitor c=0.0112985f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_319 ( N_VDD_c_316_p N_noxref_3_c_695_n ) capacitor c=0.00434174f //x=28.12 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_320 ( N_VDD_c_324_p N_noxref_3_c_695_n ) capacitor c=7.46626e-19 //x=3.645 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_321 ( N_VDD_c_328_p N_noxref_3_c_695_n ) capacitor c=0.00198565f //x=4.64 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_322 ( N_VDD_M23_noxref_d N_noxref_3_c_695_n ) capacitor c=0.0112985f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_323 ( N_VDD_c_311_n N_noxref_3_c_699_n ) capacitor c=0.043403f //x=4.81 \
 //y=7.4 //x2=4.07 //y2=2.965
cc_324 ( N_VDD_c_316_p N_noxref_3_c_662_n ) capacitor c=9.10347e-19 //x=28.12 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_325 ( N_VDD_c_311_n N_noxref_3_c_662_n ) capacitor c=0.0140736f //x=4.81 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_326 ( N_VDD_M24_noxref_s N_noxref_3_c_662_n ) capacitor c=0.0120327f \
 //x=5.765 //y=5.02 //x2=5.92 //y2=2.08
cc_327 ( N_VDD_c_316_p N_noxref_3_c_663_n ) capacitor c=9.10347e-19 //x=28.12 \
 //y=7.4 //x2=10.73 //y2=2.08
cc_328 ( N_VDD_c_312_n N_noxref_3_c_663_n ) capacitor c=0.0134015f //x=9.62 \
 //y=7.4 //x2=10.73 //y2=2.08
cc_329 ( N_VDD_M30_noxref_s N_noxref_3_c_663_n ) capacitor c=0.0125322f \
 //x=10.575 //y=5.02 //x2=10.73 //y2=2.08
cc_330 ( N_VDD_c_337_p N_noxref_3_M24_noxref_g ) capacitor c=0.00749687f \
 //x=6.695 //y=7.4 //x2=6.12 //y2=6.02
cc_331 ( N_VDD_M24_noxref_s N_noxref_3_M24_noxref_g ) capacitor c=0.0477201f \
 //x=5.765 //y=5.02 //x2=6.12 //y2=6.02
cc_332 ( N_VDD_c_337_p N_noxref_3_M25_noxref_g ) capacitor c=0.00675175f \
 //x=6.695 //y=7.4 //x2=6.56 //y2=6.02
cc_333 ( N_VDD_M25_noxref_d N_noxref_3_M25_noxref_g ) capacitor c=0.015318f \
 //x=6.635 //y=5.02 //x2=6.56 //y2=6.02
cc_334 ( N_VDD_c_341_p N_noxref_3_M30_noxref_g ) capacitor c=0.00749687f \
 //x=11.505 //y=7.4 //x2=10.93 //y2=6.02
cc_335 ( N_VDD_M30_noxref_s N_noxref_3_M30_noxref_g ) capacitor c=0.0477201f \
 //x=10.575 //y=5.02 //x2=10.93 //y2=6.02
cc_336 ( N_VDD_c_341_p N_noxref_3_M31_noxref_g ) capacitor c=0.00675175f \
 //x=11.505 //y=7.4 //x2=11.37 //y2=6.02
cc_337 ( N_VDD_M31_noxref_d N_noxref_3_M31_noxref_g ) capacitor c=0.015318f \
 //x=11.445 //y=5.02 //x2=11.37 //y2=6.02
cc_338 ( N_VDD_c_311_n N_noxref_3_c_714_n ) capacitor c=0.00757682f //x=4.81 \
 //y=7.4 //x2=6.195 //y2=4.79
cc_339 ( N_VDD_M24_noxref_s N_noxref_3_c_714_n ) capacitor c=0.00444914f \
 //x=5.765 //y=5.02 //x2=6.195 //y2=4.79
cc_340 ( N_VDD_c_312_n N_noxref_3_c_716_n ) capacitor c=0.0076931f //x=9.62 \
 //y=7.4 //x2=11.005 //y2=4.79
cc_341 ( N_VDD_M30_noxref_s N_noxref_3_c_716_n ) capacitor c=0.00444914f \
 //x=10.575 //y=5.02 //x2=11.005 //y2=4.79
cc_342 ( N_VDD_c_316_p N_noxref_3_M18_noxref_d ) capacitor c=0.00706456f \
 //x=28.12 //y=7.4 //x2=1.385 //y2=5.02
cc_343 ( N_VDD_c_317_p N_noxref_3_M18_noxref_d ) capacitor c=0.0138437f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_344 ( N_VDD_M19_noxref_d N_noxref_3_M18_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_345 ( N_VDD_c_316_p N_noxref_3_M20_noxref_d ) capacitor c=0.00275186f \
 //x=28.12 //y=7.4 //x2=2.265 //y2=5.02
cc_346 ( N_VDD_c_318_p N_noxref_3_M20_noxref_d ) capacitor c=0.0140346f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_347 ( N_VDD_c_311_n N_noxref_3_M20_noxref_d ) capacitor c=4.9285e-19 \
 //x=4.81 //y=7.4 //x2=2.265 //y2=5.02
cc_348 ( N_VDD_M18_noxref_s N_noxref_3_M20_noxref_d ) capacitor c=0.00130656f \
 //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_349 ( N_VDD_M19_noxref_d N_noxref_3_M20_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_350 ( N_VDD_M21_noxref_d N_noxref_3_M20_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_351 ( N_VDD_c_316_p N_noxref_3_M22_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=3.145 //y2=5.02
cc_352 ( N_VDD_c_324_p N_noxref_3_M22_noxref_d ) capacitor c=0.0137384f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_353 ( N_VDD_c_311_n N_noxref_3_M22_noxref_d ) capacitor c=0.00939849f \
 //x=4.81 //y=7.4 //x2=3.145 //y2=5.02
cc_354 ( N_VDD_M21_noxref_d N_noxref_3_M22_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_355 ( N_VDD_M23_noxref_d N_noxref_3_M22_noxref_d ) capacitor c=0.0664752f \
 //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_356 ( N_VDD_M24_noxref_s N_noxref_3_M22_noxref_d ) capacitor c=3.57641e-19 \
 //x=5.765 //y=5.02 //x2=3.145 //y2=5.02
cc_357 ( N_VDD_c_316_p N_noxref_4_c_916_n ) capacitor c=0.00444892f //x=28.12 \
 //y=7.4 //x2=11.945 //y2=5.155
cc_358 ( N_VDD_c_341_p N_noxref_4_c_916_n ) capacitor c=4.31931e-19 //x=11.505 \
 //y=7.4 //x2=11.945 //y2=5.155
cc_359 ( N_VDD_c_366_p N_noxref_4_c_916_n ) capacitor c=4.31931e-19 //x=12.385 \
 //y=7.4 //x2=11.945 //y2=5.155
cc_360 ( N_VDD_M31_noxref_d N_noxref_4_c_916_n ) capacitor c=0.0112985f \
 //x=11.445 //y=5.02 //x2=11.945 //y2=5.155
cc_361 ( N_VDD_c_312_n N_noxref_4_c_920_n ) capacitor c=0.00863585f //x=9.62 \
 //y=7.4 //x2=11.235 //y2=5.155
cc_362 ( N_VDD_M30_noxref_s N_noxref_4_c_920_n ) capacitor c=0.0831083f \
 //x=10.575 //y=5.02 //x2=11.235 //y2=5.155
cc_363 ( N_VDD_c_316_p N_noxref_4_c_922_n ) capacitor c=0.0044221f //x=28.12 \
 //y=7.4 //x2=12.825 //y2=5.155
cc_364 ( N_VDD_c_366_p N_noxref_4_c_922_n ) capacitor c=4.31931e-19 //x=12.385 \
 //y=7.4 //x2=12.825 //y2=5.155
cc_365 ( N_VDD_c_372_p N_noxref_4_c_922_n ) capacitor c=4.31931e-19 //x=13.265 \
 //y=7.4 //x2=12.825 //y2=5.155
cc_366 ( N_VDD_M33_noxref_d N_noxref_4_c_922_n ) capacitor c=0.0112985f \
 //x=12.325 //y=5.02 //x2=12.825 //y2=5.155
cc_367 ( N_VDD_c_316_p N_noxref_4_c_926_n ) capacitor c=0.00434174f //x=28.12 \
 //y=7.4 //x2=13.605 //y2=5.155
cc_368 ( N_VDD_c_372_p N_noxref_4_c_926_n ) capacitor c=7.46626e-19 //x=13.265 \
 //y=7.4 //x2=13.605 //y2=5.155
cc_369 ( N_VDD_c_376_p N_noxref_4_c_926_n ) capacitor c=0.00198565f //x=14.26 \
 //y=7.4 //x2=13.605 //y2=5.155
cc_370 ( N_VDD_M35_noxref_d N_noxref_4_c_926_n ) capacitor c=0.0112985f \
 //x=13.205 //y=5.02 //x2=13.605 //y2=5.155
cc_371 ( N_VDD_c_313_n N_noxref_4_c_930_n ) capacitor c=0.0427356f //x=14.43 \
 //y=7.4 //x2=13.69 //y2=2.96
cc_372 ( N_VDD_c_316_p N_noxref_4_c_904_n ) capacitor c=9.10347e-19 //x=28.12 \
 //y=7.4 //x2=15.54 //y2=2.08
cc_373 ( N_VDD_c_313_n N_noxref_4_c_904_n ) capacitor c=0.0133888f //x=14.43 \
 //y=7.4 //x2=15.54 //y2=2.08
cc_374 ( N_VDD_M36_noxref_s N_noxref_4_c_904_n ) capacitor c=0.0125322f \
 //x=15.385 //y=5.02 //x2=15.54 //y2=2.08
cc_375 ( N_VDD_c_382_p N_noxref_4_M36_noxref_g ) capacitor c=0.00749687f \
 //x=16.315 //y=7.4 //x2=15.74 //y2=6.02
cc_376 ( N_VDD_M36_noxref_s N_noxref_4_M36_noxref_g ) capacitor c=0.0477201f \
 //x=15.385 //y=5.02 //x2=15.74 //y2=6.02
cc_377 ( N_VDD_c_382_p N_noxref_4_M37_noxref_g ) capacitor c=0.00675175f \
 //x=16.315 //y=7.4 //x2=16.18 //y2=6.02
cc_378 ( N_VDD_M37_noxref_d N_noxref_4_M37_noxref_g ) capacitor c=0.015318f \
 //x=16.255 //y=5.02 //x2=16.18 //y2=6.02
cc_379 ( N_VDD_c_313_n N_noxref_4_c_938_n ) capacitor c=0.00757682f //x=14.43 \
 //y=7.4 //x2=15.815 //y2=4.79
cc_380 ( N_VDD_M36_noxref_s N_noxref_4_c_938_n ) capacitor c=0.00444914f \
 //x=15.385 //y=5.02 //x2=15.815 //y2=4.79
cc_381 ( N_VDD_c_316_p N_noxref_4_M30_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=11.005 //y2=5.02
cc_382 ( N_VDD_c_341_p N_noxref_4_M30_noxref_d ) capacitor c=0.014035f \
 //x=11.505 //y=7.4 //x2=11.005 //y2=5.02
cc_383 ( N_VDD_M31_noxref_d N_noxref_4_M30_noxref_d ) capacitor c=0.0664752f \
 //x=11.445 //y=5.02 //x2=11.005 //y2=5.02
cc_384 ( N_VDD_c_316_p N_noxref_4_M32_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=11.885 //y2=5.02
cc_385 ( N_VDD_c_366_p N_noxref_4_M32_noxref_d ) capacitor c=0.014035f \
 //x=12.385 //y=7.4 //x2=11.885 //y2=5.02
cc_386 ( N_VDD_c_313_n N_noxref_4_M32_noxref_d ) capacitor c=4.9285e-19 \
 //x=14.43 //y=7.4 //x2=11.885 //y2=5.02
cc_387 ( N_VDD_M30_noxref_s N_noxref_4_M32_noxref_d ) capacitor c=0.00130656f \
 //x=10.575 //y=5.02 //x2=11.885 //y2=5.02
cc_388 ( N_VDD_M31_noxref_d N_noxref_4_M32_noxref_d ) capacitor c=0.0664752f \
 //x=11.445 //y=5.02 //x2=11.885 //y2=5.02
cc_389 ( N_VDD_M33_noxref_d N_noxref_4_M32_noxref_d ) capacitor c=0.0664752f \
 //x=12.325 //y=5.02 //x2=11.885 //y2=5.02
cc_390 ( N_VDD_c_316_p N_noxref_4_M34_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=12.765 //y2=5.02
cc_391 ( N_VDD_c_372_p N_noxref_4_M34_noxref_d ) capacitor c=0.014035f \
 //x=13.265 //y=7.4 //x2=12.765 //y2=5.02
cc_392 ( N_VDD_c_313_n N_noxref_4_M34_noxref_d ) capacitor c=0.00939849f \
 //x=14.43 //y=7.4 //x2=12.765 //y2=5.02
cc_393 ( N_VDD_M33_noxref_d N_noxref_4_M34_noxref_d ) capacitor c=0.0664752f \
 //x=12.325 //y=5.02 //x2=12.765 //y2=5.02
cc_394 ( N_VDD_M35_noxref_d N_noxref_4_M34_noxref_d ) capacitor c=0.0664752f \
 //x=13.205 //y=5.02 //x2=12.765 //y2=5.02
cc_395 ( N_VDD_M36_noxref_s N_noxref_4_M34_noxref_d ) capacitor c=3.57641e-19 \
 //x=15.385 //y=5.02 //x2=12.765 //y2=5.02
cc_396 ( N_VDD_c_316_p N_CLK_c_1063_n ) capacitor c=2.03486e-19 //x=28.12 \
 //y=7.4 //x2=7.03 //y2=2.08
cc_397 ( N_VDD_c_311_n N_CLK_c_1063_n ) capacitor c=6.95672e-19 //x=4.81 \
 //y=7.4 //x2=7.03 //y2=2.08
cc_398 ( N_VDD_c_316_p N_CLK_c_1064_n ) capacitor c=2.03486e-19 //x=28.12 \
 //y=7.4 //x2=16.65 //y2=2.08
cc_399 ( N_VDD_c_313_n N_CLK_c_1064_n ) capacitor c=6.29521e-19 //x=14.43 \
 //y=7.4 //x2=16.65 //y2=2.08
cc_400 ( N_VDD_c_407_p N_CLK_M26_noxref_g ) capacitor c=0.00676195f //x=7.575 \
 //y=7.4 //x2=7 //y2=6.02
cc_401 ( N_VDD_M25_noxref_d N_CLK_M26_noxref_g ) capacitor c=0.015318f \
 //x=6.635 //y=5.02 //x2=7 //y2=6.02
cc_402 ( N_VDD_c_407_p N_CLK_M27_noxref_g ) capacitor c=0.00675175f //x=7.575 \
 //y=7.4 //x2=7.44 //y2=6.02
cc_403 ( N_VDD_M27_noxref_d N_CLK_M27_noxref_g ) capacitor c=0.015318f \
 //x=7.515 //y=5.02 //x2=7.44 //y2=6.02
cc_404 ( N_VDD_c_411_p N_CLK_M38_noxref_g ) capacitor c=0.00676195f //x=17.195 \
 //y=7.4 //x2=16.62 //y2=6.02
cc_405 ( N_VDD_M37_noxref_d N_CLK_M38_noxref_g ) capacitor c=0.015318f \
 //x=16.255 //y=5.02 //x2=16.62 //y2=6.02
cc_406 ( N_VDD_c_411_p N_CLK_M39_noxref_g ) capacitor c=0.00675175f //x=17.195 \
 //y=7.4 //x2=17.06 //y2=6.02
cc_407 ( N_VDD_M39_noxref_d N_CLK_M39_noxref_g ) capacitor c=0.015318f \
 //x=17.135 //y=5.02 //x2=17.06 //y2=6.02
cc_408 ( N_VDD_c_311_n N_noxref_6_c_1253_n ) capacitor c=0.00686843f //x=4.81 \
 //y=7.4 //x2=8.765 //y2=3.7
cc_409 ( N_VDD_c_311_n N_noxref_6_c_1256_n ) capacitor c=7.23426e-19 //x=4.81 \
 //y=7.4 //x2=3.33 //y2=2.08
cc_410 ( N_VDD_c_316_p N_noxref_6_c_1272_n ) capacitor c=0.00444892f //x=28.12 \
 //y=7.4 //x2=7.135 //y2=5.155
cc_411 ( N_VDD_c_337_p N_noxref_6_c_1272_n ) capacitor c=4.31931e-19 //x=6.695 \
 //y=7.4 //x2=7.135 //y2=5.155
cc_412 ( N_VDD_c_407_p N_noxref_6_c_1272_n ) capacitor c=4.31931e-19 //x=7.575 \
 //y=7.4 //x2=7.135 //y2=5.155
cc_413 ( N_VDD_M25_noxref_d N_noxref_6_c_1272_n ) capacitor c=0.0112985f \
 //x=6.635 //y=5.02 //x2=7.135 //y2=5.155
cc_414 ( N_VDD_c_311_n N_noxref_6_c_1276_n ) capacitor c=0.00863585f //x=4.81 \
 //y=7.4 //x2=6.425 //y2=5.155
cc_415 ( N_VDD_M24_noxref_s N_noxref_6_c_1276_n ) capacitor c=0.0831083f \
 //x=5.765 //y=5.02 //x2=6.425 //y2=5.155
cc_416 ( N_VDD_c_316_p N_noxref_6_c_1278_n ) capacitor c=0.0044221f //x=28.12 \
 //y=7.4 //x2=8.015 //y2=5.155
cc_417 ( N_VDD_c_407_p N_noxref_6_c_1278_n ) capacitor c=4.31931e-19 //x=7.575 \
 //y=7.4 //x2=8.015 //y2=5.155
cc_418 ( N_VDD_c_425_p N_noxref_6_c_1278_n ) capacitor c=4.31931e-19 //x=8.455 \
 //y=7.4 //x2=8.015 //y2=5.155
cc_419 ( N_VDD_M27_noxref_d N_noxref_6_c_1278_n ) capacitor c=0.0112985f \
 //x=7.515 //y=5.02 //x2=8.015 //y2=5.155
cc_420 ( N_VDD_c_316_p N_noxref_6_c_1282_n ) capacitor c=0.00434174f //x=28.12 \
 //y=7.4 //x2=8.795 //y2=5.155
cc_421 ( N_VDD_c_425_p N_noxref_6_c_1282_n ) capacitor c=7.46626e-19 //x=8.455 \
 //y=7.4 //x2=8.795 //y2=5.155
cc_422 ( N_VDD_c_429_p N_noxref_6_c_1282_n ) capacitor c=0.00198565f //x=9.45 \
 //y=7.4 //x2=8.795 //y2=5.155
cc_423 ( N_VDD_M29_noxref_d N_noxref_6_c_1282_n ) capacitor c=0.0112985f \
 //x=8.395 //y=5.02 //x2=8.795 //y2=5.155
cc_424 ( N_VDD_c_312_n N_noxref_6_c_1286_n ) capacitor c=0.0427358f //x=9.62 \
 //y=7.4 //x2=8.88 //y2=3.7
cc_425 ( N_VDD_c_316_p N_noxref_6_c_1258_n ) capacitor c=9.10347e-19 //x=28.12 \
 //y=7.4 //x2=20.35 //y2=2.08
cc_426 ( N_VDD_c_314_n N_noxref_6_c_1258_n ) capacitor c=0.013309f //x=19.24 \
 //y=7.4 //x2=20.35 //y2=2.08
cc_427 ( N_VDD_M42_noxref_s N_noxref_6_c_1258_n ) capacitor c=0.0120327f \
 //x=20.195 //y=5.02 //x2=20.35 //y2=2.08
cc_428 ( N_VDD_c_324_p N_noxref_6_M22_noxref_g ) capacitor c=0.00675175f \
 //x=3.645 //y=7.4 //x2=3.07 //y2=6.02
cc_429 ( N_VDD_M21_noxref_d N_noxref_6_M22_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=3.07 //y2=6.02
cc_430 ( N_VDD_c_324_p N_noxref_6_M23_noxref_g ) capacitor c=0.00675379f \
 //x=3.645 //y=7.4 //x2=3.51 //y2=6.02
cc_431 ( N_VDD_M23_noxref_d N_noxref_6_M23_noxref_g ) capacitor c=0.0394719f \
 //x=3.585 //y=5.02 //x2=3.51 //y2=6.02
cc_432 ( N_VDD_c_439_p N_noxref_6_M42_noxref_g ) capacitor c=0.00749687f \
 //x=21.125 //y=7.4 //x2=20.55 //y2=6.02
cc_433 ( N_VDD_M42_noxref_s N_noxref_6_M42_noxref_g ) capacitor c=0.0477201f \
 //x=20.195 //y=5.02 //x2=20.55 //y2=6.02
cc_434 ( N_VDD_c_439_p N_noxref_6_M43_noxref_g ) capacitor c=0.00675175f \
 //x=21.125 //y=7.4 //x2=20.99 //y2=6.02
cc_435 ( N_VDD_M43_noxref_d N_noxref_6_M43_noxref_g ) capacitor c=0.015318f \
 //x=21.065 //y=5.02 //x2=20.99 //y2=6.02
cc_436 ( N_VDD_c_314_n N_noxref_6_c_1298_n ) capacitor c=0.00757682f //x=19.24 \
 //y=7.4 //x2=20.625 //y2=4.79
cc_437 ( N_VDD_M42_noxref_s N_noxref_6_c_1298_n ) capacitor c=0.00444914f \
 //x=20.195 //y=5.02 //x2=20.625 //y2=4.79
cc_438 ( N_VDD_c_316_p N_noxref_6_M24_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=6.195 //y2=5.02
cc_439 ( N_VDD_c_337_p N_noxref_6_M24_noxref_d ) capacitor c=0.014035f \
 //x=6.695 //y=7.4 //x2=6.195 //y2=5.02
cc_440 ( N_VDD_M25_noxref_d N_noxref_6_M24_noxref_d ) capacitor c=0.0664752f \
 //x=6.635 //y=5.02 //x2=6.195 //y2=5.02
cc_441 ( N_VDD_c_316_p N_noxref_6_M26_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=7.075 //y2=5.02
cc_442 ( N_VDD_c_407_p N_noxref_6_M26_noxref_d ) capacitor c=0.014035f \
 //x=7.575 //y=7.4 //x2=7.075 //y2=5.02
cc_443 ( N_VDD_c_312_n N_noxref_6_M26_noxref_d ) capacitor c=4.9285e-19 \
 //x=9.62 //y=7.4 //x2=7.075 //y2=5.02
cc_444 ( N_VDD_M24_noxref_s N_noxref_6_M26_noxref_d ) capacitor c=0.00130656f \
 //x=5.765 //y=5.02 //x2=7.075 //y2=5.02
cc_445 ( N_VDD_M25_noxref_d N_noxref_6_M26_noxref_d ) capacitor c=0.0664752f \
 //x=6.635 //y=5.02 //x2=7.075 //y2=5.02
cc_446 ( N_VDD_M27_noxref_d N_noxref_6_M26_noxref_d ) capacitor c=0.0664752f \
 //x=7.515 //y=5.02 //x2=7.075 //y2=5.02
cc_447 ( N_VDD_c_316_p N_noxref_6_M28_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=7.955 //y2=5.02
cc_448 ( N_VDD_c_425_p N_noxref_6_M28_noxref_d ) capacitor c=0.014035f \
 //x=8.455 //y=7.4 //x2=7.955 //y2=5.02
cc_449 ( N_VDD_c_312_n N_noxref_6_M28_noxref_d ) capacitor c=0.00939849f \
 //x=9.62 //y=7.4 //x2=7.955 //y2=5.02
cc_450 ( N_VDD_M27_noxref_d N_noxref_6_M28_noxref_d ) capacitor c=0.0664752f \
 //x=7.515 //y=5.02 //x2=7.955 //y2=5.02
cc_451 ( N_VDD_M29_noxref_d N_noxref_6_M28_noxref_d ) capacitor c=0.0664752f \
 //x=8.395 //y=5.02 //x2=7.955 //y2=5.02
cc_452 ( N_VDD_M30_noxref_s N_noxref_6_M28_noxref_d ) capacitor c=3.57641e-19 \
 //x=10.575 //y=5.02 //x2=7.955 //y2=5.02
cc_453 ( N_VDD_c_316_p N_RN_c_1514_n ) capacitor c=0.115493f //x=28.12 //y=7.4 \
 //x2=17.645 //y2=4.44
cc_454 ( N_VDD_c_328_p N_RN_c_1514_n ) capacitor c=0.00258496f //x=4.64 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_455 ( N_VDD_c_462_p N_RN_c_1514_n ) capacitor c=0.00328994f //x=5.815 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_456 ( N_VDD_c_337_p N_RN_c_1514_n ) capacitor c=0.00135925f //x=6.695 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_457 ( N_VDD_c_429_p N_RN_c_1514_n ) capacitor c=0.00258496f //x=9.45 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_458 ( N_VDD_c_465_p N_RN_c_1514_n ) capacitor c=0.00328994f //x=10.625 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_459 ( N_VDD_c_341_p N_RN_c_1514_n ) capacitor c=0.00135925f //x=11.505 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_460 ( N_VDD_c_376_p N_RN_c_1514_n ) capacitor c=0.00258496f //x=14.26 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_461 ( N_VDD_c_468_p N_RN_c_1514_n ) capacitor c=0.00328994f //x=15.435 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_462 ( N_VDD_c_382_p N_RN_c_1514_n ) capacitor c=0.00135925f //x=16.315 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_463 ( N_VDD_c_311_n N_RN_c_1514_n ) capacitor c=0.0375613f //x=4.81 //y=7.4 \
 //x2=17.645 //y2=4.44
cc_464 ( N_VDD_c_312_n N_RN_c_1514_n ) capacitor c=0.0389825f //x=9.62 //y=7.4 \
 //x2=17.645 //y2=4.44
cc_465 ( N_VDD_c_313_n N_RN_c_1514_n ) capacitor c=0.0389825f //x=14.43 \
 //y=7.4 //x2=17.645 //y2=4.44
cc_466 ( N_VDD_M24_noxref_s N_RN_c_1514_n ) capacitor c=0.00179496f //x=5.765 \
 //y=5.02 //x2=17.645 //y2=4.44
cc_467 ( N_VDD_M30_noxref_s N_RN_c_1514_n ) capacitor c=0.00179496f //x=10.575 \
 //y=5.02 //x2=17.645 //y2=4.44
cc_468 ( N_VDD_M36_noxref_s N_RN_c_1514_n ) capacitor c=0.00179496f //x=15.385 \
 //y=5.02 //x2=17.645 //y2=4.44
cc_469 ( N_VDD_c_316_p N_RN_c_1515_n ) capacitor c=0.00146066f //x=28.12 \
 //y=7.4 //x2=2.335 //y2=4.44
cc_470 ( N_VDD_c_316_p N_RN_c_1536_n ) capacitor c=0.0282652f //x=28.12 \
 //y=7.4 //x2=21.345 //y2=4.44
cc_471 ( N_VDD_c_478_p N_RN_c_1536_n ) capacitor c=0.00258496f //x=19.07 \
 //y=7.4 //x2=21.345 //y2=4.44
cc_472 ( N_VDD_c_479_p N_RN_c_1536_n ) capacitor c=0.00328994f //x=20.245 \
 //y=7.4 //x2=21.345 //y2=4.44
cc_473 ( N_VDD_c_439_p N_RN_c_1536_n ) capacitor c=0.00135925f //x=21.125 \
 //y=7.4 //x2=21.345 //y2=4.44
cc_474 ( N_VDD_c_314_n N_RN_c_1536_n ) capacitor c=0.0389825f //x=19.24 \
 //y=7.4 //x2=21.345 //y2=4.44
cc_475 ( N_VDD_M42_noxref_s N_RN_c_1536_n ) capacitor c=0.00179496f //x=20.195 \
 //y=5.02 //x2=21.345 //y2=4.44
cc_476 ( N_VDD_c_316_p N_RN_c_1542_n ) capacitor c=0.00110755f //x=28.12 \
 //y=7.4 //x2=17.875 //y2=4.44
cc_477 ( N_VDD_c_316_p N_RN_c_1516_n ) capacitor c=2.03287e-19 //x=28.12 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_478 ( N_VDD_c_309_n N_RN_c_1516_n ) capacitor c=8.7832e-19 //x=0.74 //y=7.4 \
 //x2=2.22 //y2=2.08
cc_479 ( N_VDD_c_314_n N_RN_c_1517_n ) capacitor c=6.89593e-19 //x=19.24 \
 //y=7.4 //x2=17.76 //y2=2.08
cc_480 ( N_VDD_c_316_p N_RN_c_1518_n ) capacitor c=2.03287e-19 //x=28.12 \
 //y=7.4 //x2=21.46 //y2=2.08
cc_481 ( N_VDD_c_314_n N_RN_c_1518_n ) capacitor c=6.41871e-19 //x=19.24 \
 //y=7.4 //x2=21.46 //y2=2.08
cc_482 ( N_VDD_c_318_p N_RN_M20_noxref_g ) capacitor c=0.00676195f //x=2.765 \
 //y=7.4 //x2=2.19 //y2=6.02
cc_483 ( N_VDD_M19_noxref_d N_RN_M20_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=2.19 //y2=6.02
cc_484 ( N_VDD_c_318_p N_RN_M21_noxref_g ) capacitor c=0.00675175f //x=2.765 \
 //y=7.4 //x2=2.63 //y2=6.02
cc_485 ( N_VDD_M21_noxref_d N_RN_M21_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=2.63 //y2=6.02
cc_486 ( N_VDD_c_493_p N_RN_M40_noxref_g ) capacitor c=0.00675175f //x=18.075 \
 //y=7.4 //x2=17.5 //y2=6.02
cc_487 ( N_VDD_M39_noxref_d N_RN_M40_noxref_g ) capacitor c=0.015318f \
 //x=17.135 //y=5.02 //x2=17.5 //y2=6.02
cc_488 ( N_VDD_c_493_p N_RN_M41_noxref_g ) capacitor c=0.00675379f //x=18.075 \
 //y=7.4 //x2=17.94 //y2=6.02
cc_489 ( N_VDD_M41_noxref_d N_RN_M41_noxref_g ) capacitor c=0.0394719f \
 //x=18.015 //y=5.02 //x2=17.94 //y2=6.02
cc_490 ( N_VDD_c_497_p N_RN_M44_noxref_g ) capacitor c=0.00676195f //x=22.005 \
 //y=7.4 //x2=21.43 //y2=6.02
cc_491 ( N_VDD_M43_noxref_d N_RN_M44_noxref_g ) capacitor c=0.015318f \
 //x=21.065 //y=5.02 //x2=21.43 //y2=6.02
cc_492 ( N_VDD_c_497_p N_RN_M45_noxref_g ) capacitor c=0.00675175f //x=22.005 \
 //y=7.4 //x2=21.87 //y2=6.02
cc_493 ( N_VDD_M45_noxref_d N_RN_M45_noxref_g ) capacitor c=0.015318f \
 //x=21.945 //y=5.02 //x2=21.87 //y2=6.02
cc_494 ( N_VDD_c_315_n QN ) capacitor c=0.045031f //x=24.05 //y=7.4 //x2=23.31 \
 //y2=2.22
cc_495 ( N_VDD_c_316_p N_QN_c_1838_n ) capacitor c=0.00444751f //x=28.12 \
 //y=7.4 //x2=21.565 //y2=5.155
cc_496 ( N_VDD_c_439_p N_QN_c_1838_n ) capacitor c=4.31931e-19 //x=21.125 \
 //y=7.4 //x2=21.565 //y2=5.155
cc_497 ( N_VDD_c_497_p N_QN_c_1838_n ) capacitor c=4.31906e-19 //x=22.005 \
 //y=7.4 //x2=21.565 //y2=5.155
cc_498 ( N_VDD_M43_noxref_d N_QN_c_1838_n ) capacitor c=0.0112985f //x=21.065 \
 //y=5.02 //x2=21.565 //y2=5.155
cc_499 ( N_VDD_c_314_n N_QN_c_1842_n ) capacitor c=0.00863585f //x=19.24 \
 //y=7.4 //x2=20.855 //y2=5.155
cc_500 ( N_VDD_M42_noxref_s N_QN_c_1842_n ) capacitor c=0.0831083f //x=20.195 \
 //y=5.02 //x2=20.855 //y2=5.155
cc_501 ( N_VDD_c_316_p N_QN_c_1844_n ) capacitor c=0.00448996f //x=28.12 \
 //y=7.4 //x2=22.445 //y2=5.155
cc_502 ( N_VDD_c_497_p N_QN_c_1844_n ) capacitor c=4.32228e-19 //x=22.005 \
 //y=7.4 //x2=22.445 //y2=5.155
cc_503 ( N_VDD_c_510_p N_QN_c_1844_n ) capacitor c=4.32228e-19 //x=22.885 \
 //y=7.4 //x2=22.445 //y2=5.155
cc_504 ( N_VDD_M45_noxref_d N_QN_c_1844_n ) capacitor c=0.0115147f //x=21.945 \
 //y=5.02 //x2=22.445 //y2=5.155
cc_505 ( N_VDD_c_316_p N_QN_c_1848_n ) capacitor c=0.00442621f //x=28.12 \
 //y=7.4 //x2=23.225 //y2=5.155
cc_506 ( N_VDD_c_510_p N_QN_c_1848_n ) capacitor c=7.47666e-19 //x=22.885 \
 //y=7.4 //x2=23.225 //y2=5.155
cc_507 ( N_VDD_c_514_p N_QN_c_1848_n ) capacitor c=0.00198981f //x=23.88 \
 //y=7.4 //x2=23.225 //y2=5.155
cc_508 ( N_VDD_M47_noxref_d N_QN_c_1848_n ) capacitor c=0.0115147f //x=22.825 \
 //y=5.02 //x2=23.225 //y2=5.155
cc_509 ( N_VDD_c_316_p N_QN_c_1825_n ) capacitor c=9.23542e-19 //x=28.12 \
 //y=7.4 //x2=25.16 //y2=2.08
cc_510 ( N_VDD_c_315_n N_QN_c_1825_n ) capacitor c=0.0160291f //x=24.05 \
 //y=7.4 //x2=25.16 //y2=2.08
cc_511 ( N_VDD_M48_noxref_s N_QN_c_1825_n ) capacitor c=0.0123142f //x=25.005 \
 //y=5.02 //x2=25.16 //y2=2.08
cc_512 ( N_VDD_c_519_p N_QN_M48_noxref_g ) capacitor c=0.00749687f //x=25.935 \
 //y=7.4 //x2=25.36 //y2=6.02
cc_513 ( N_VDD_M48_noxref_s N_QN_M48_noxref_g ) capacitor c=0.0477201f \
 //x=25.005 //y=5.02 //x2=25.36 //y2=6.02
cc_514 ( N_VDD_c_519_p N_QN_M49_noxref_g ) capacitor c=0.00675175f //x=25.935 \
 //y=7.4 //x2=25.8 //y2=6.02
cc_515 ( N_VDD_M49_noxref_d N_QN_M49_noxref_g ) capacitor c=0.015318f \
 //x=25.875 //y=5.02 //x2=25.8 //y2=6.02
cc_516 ( N_VDD_c_315_n N_QN_c_1859_n ) capacitor c=0.00757682f //x=24.05 \
 //y=7.4 //x2=25.435 //y2=4.79
cc_517 ( N_VDD_M48_noxref_s N_QN_c_1859_n ) capacitor c=0.00445134f //x=25.005 \
 //y=5.02 //x2=25.435 //y2=4.79
cc_518 ( N_VDD_c_316_p N_QN_M42_noxref_d ) capacitor c=0.00275235f //x=28.12 \
 //y=7.4 //x2=20.625 //y2=5.02
cc_519 ( N_VDD_c_439_p N_QN_M42_noxref_d ) capacitor c=0.014035f //x=21.125 \
 //y=7.4 //x2=20.625 //y2=5.02
cc_520 ( N_VDD_M43_noxref_d N_QN_M42_noxref_d ) capacitor c=0.0664752f \
 //x=21.065 //y=5.02 //x2=20.625 //y2=5.02
cc_521 ( N_VDD_c_316_p N_QN_M44_noxref_d ) capacitor c=0.00282723f //x=28.12 \
 //y=7.4 //x2=21.505 //y2=5.02
cc_522 ( N_VDD_c_497_p N_QN_M44_noxref_d ) capacitor c=0.0140856f //x=22.005 \
 //y=7.4 //x2=21.505 //y2=5.02
cc_523 ( N_VDD_c_315_n N_QN_M44_noxref_d ) capacitor c=4.9285e-19 //x=24.05 \
 //y=7.4 //x2=21.505 //y2=5.02
cc_524 ( N_VDD_M42_noxref_s N_QN_M44_noxref_d ) capacitor c=0.00130656f \
 //x=20.195 //y=5.02 //x2=21.505 //y2=5.02
cc_525 ( N_VDD_M43_noxref_d N_QN_M44_noxref_d ) capacitor c=0.0664752f \
 //x=21.065 //y=5.02 //x2=21.505 //y2=5.02
cc_526 ( N_VDD_M45_noxref_d N_QN_M44_noxref_d ) capacitor c=0.0664752f \
 //x=21.945 //y=5.02 //x2=21.505 //y2=5.02
cc_527 ( N_VDD_c_316_p N_QN_M46_noxref_d ) capacitor c=0.00285091f //x=28.12 \
 //y=7.4 //x2=22.385 //y2=5.02
cc_528 ( N_VDD_c_510_p N_QN_M46_noxref_d ) capacitor c=0.0138051f //x=22.885 \
 //y=7.4 //x2=22.385 //y2=5.02
cc_529 ( N_VDD_c_315_n N_QN_M46_noxref_d ) capacitor c=0.00939849f //x=24.05 \
 //y=7.4 //x2=22.385 //y2=5.02
cc_530 ( N_VDD_M45_noxref_d N_QN_M46_noxref_d ) capacitor c=0.0664752f \
 //x=21.945 //y=5.02 //x2=22.385 //y2=5.02
cc_531 ( N_VDD_M47_noxref_d N_QN_M46_noxref_d ) capacitor c=0.0664752f \
 //x=22.825 //y=5.02 //x2=22.385 //y2=5.02
cc_532 ( N_VDD_M48_noxref_s N_QN_M46_noxref_d ) capacitor c=3.57641e-19 \
 //x=25.005 //y=5.02 //x2=22.385 //y2=5.02
cc_533 ( N_VDD_c_316_p N_SN_c_1991_n ) capacitor c=2.03486e-19 //x=28.12 \
 //y=7.4 //x2=11.84 //y2=2.08
cc_534 ( N_VDD_c_312_n N_SN_c_1991_n ) capacitor c=6.19572e-19 //x=9.62 \
 //y=7.4 //x2=11.84 //y2=2.08
cc_535 ( N_VDD_c_316_p N_SN_c_1992_n ) capacitor c=2.05828e-19 //x=28.12 \
 //y=7.4 //x2=26.27 //y2=2.08
cc_536 ( N_VDD_c_315_n N_SN_c_1992_n ) capacitor c=7.34568e-19 //x=24.05 \
 //y=7.4 //x2=26.27 //y2=2.08
cc_537 ( N_VDD_c_366_p N_SN_M32_noxref_g ) capacitor c=0.00676195f //x=12.385 \
 //y=7.4 //x2=11.81 //y2=6.02
cc_538 ( N_VDD_M31_noxref_d N_SN_M32_noxref_g ) capacitor c=0.015318f \
 //x=11.445 //y=5.02 //x2=11.81 //y2=6.02
cc_539 ( N_VDD_c_366_p N_SN_M33_noxref_g ) capacitor c=0.00675175f //x=12.385 \
 //y=7.4 //x2=12.25 //y2=6.02
cc_540 ( N_VDD_M33_noxref_d N_SN_M33_noxref_g ) capacitor c=0.015318f \
 //x=12.325 //y=5.02 //x2=12.25 //y2=6.02
cc_541 ( N_VDD_c_548_p N_SN_M50_noxref_g ) capacitor c=0.00676195f //x=26.815 \
 //y=7.4 //x2=26.24 //y2=6.02
cc_542 ( N_VDD_M49_noxref_d N_SN_M50_noxref_g ) capacitor c=0.015318f \
 //x=25.875 //y=5.02 //x2=26.24 //y2=6.02
cc_543 ( N_VDD_c_548_p N_SN_M51_noxref_g ) capacitor c=0.00675175f //x=26.815 \
 //y=7.4 //x2=26.68 //y2=6.02
cc_544 ( N_VDD_M51_noxref_d N_SN_M51_noxref_g ) capacitor c=0.015318f \
 //x=26.755 //y=5.02 //x2=26.68 //y2=6.02
cc_545 ( N_VDD_c_312_n N_noxref_10_c_2214_n ) capacitor c=0.0140578f //x=9.62 \
 //y=7.4 //x2=12.835 //y2=4.07
cc_546 ( N_VDD_c_313_n N_noxref_10_c_2215_n ) capacitor c=0.0140578f //x=14.43 \
 //y=7.4 //x2=18.385 //y2=4.07
cc_547 ( N_VDD_c_316_p N_noxref_10_c_2216_n ) capacitor c=0.0524622f //x=28.12 \
 //y=7.4 //x2=27.265 //y2=4.07
cc_548 ( N_VDD_c_514_p N_noxref_10_c_2216_n ) capacitor c=0.00214241f \
 //x=23.88 //y=7.4 //x2=27.265 //y2=4.07
cc_549 ( N_VDD_c_556_p N_noxref_10_c_2216_n ) capacitor c=0.0027159f \
 //x=25.055 //y=7.4 //x2=27.265 //y2=4.07
cc_550 ( N_VDD_c_519_p N_noxref_10_c_2216_n ) capacitor c=0.00113459f \
 //x=25.935 //y=7.4 //x2=27.265 //y2=4.07
cc_551 ( N_VDD_c_314_n N_noxref_10_c_2216_n ) capacitor c=0.0140578f //x=19.24 \
 //y=7.4 //x2=27.265 //y2=4.07
cc_552 ( N_VDD_c_315_n N_noxref_10_c_2216_n ) capacitor c=0.0269494f //x=24.05 \
 //y=7.4 //x2=27.265 //y2=4.07
cc_553 ( N_VDD_M48_noxref_s N_noxref_10_c_2216_n ) capacitor c=0.00122826f \
 //x=25.005 //y=5.02 //x2=27.265 //y2=4.07
cc_554 ( N_VDD_c_314_n N_noxref_10_c_2223_n ) capacitor c=0.00104972f \
 //x=19.24 //y=7.4 //x2=18.615 //y2=4.07
cc_555 ( N_VDD_c_313_n N_noxref_10_c_2210_n ) capacitor c=5.93913e-19 \
 //x=14.43 //y=7.4 //x2=12.95 //y2=2.08
cc_556 ( N_VDD_c_316_p N_noxref_10_c_2225_n ) capacitor c=0.00444892f \
 //x=28.12 //y=7.4 //x2=16.755 //y2=5.155
cc_557 ( N_VDD_c_382_p N_noxref_10_c_2225_n ) capacitor c=4.31931e-19 \
 //x=16.315 //y=7.4 //x2=16.755 //y2=5.155
cc_558 ( N_VDD_c_411_p N_noxref_10_c_2225_n ) capacitor c=4.31931e-19 \
 //x=17.195 //y=7.4 //x2=16.755 //y2=5.155
cc_559 ( N_VDD_M37_noxref_d N_noxref_10_c_2225_n ) capacitor c=0.0112985f \
 //x=16.255 //y=5.02 //x2=16.755 //y2=5.155
cc_560 ( N_VDD_c_313_n N_noxref_10_c_2229_n ) capacitor c=0.00863585f \
 //x=14.43 //y=7.4 //x2=16.045 //y2=5.155
cc_561 ( N_VDD_M36_noxref_s N_noxref_10_c_2229_n ) capacitor c=0.0831083f \
 //x=15.385 //y=5.02 //x2=16.045 //y2=5.155
cc_562 ( N_VDD_c_316_p N_noxref_10_c_2231_n ) capacitor c=0.0044221f //x=28.12 \
 //y=7.4 //x2=17.635 //y2=5.155
cc_563 ( N_VDD_c_411_p N_noxref_10_c_2231_n ) capacitor c=4.31931e-19 \
 //x=17.195 //y=7.4 //x2=17.635 //y2=5.155
cc_564 ( N_VDD_c_493_p N_noxref_10_c_2231_n ) capacitor c=4.31931e-19 \
 //x=18.075 //y=7.4 //x2=17.635 //y2=5.155
cc_565 ( N_VDD_M39_noxref_d N_noxref_10_c_2231_n ) capacitor c=0.0112985f \
 //x=17.135 //y=5.02 //x2=17.635 //y2=5.155
cc_566 ( N_VDD_c_316_p N_noxref_10_c_2235_n ) capacitor c=0.00434116f \
 //x=28.12 //y=7.4 //x2=18.415 //y2=5.155
cc_567 ( N_VDD_c_493_p N_noxref_10_c_2235_n ) capacitor c=7.46549e-19 \
 //x=18.075 //y=7.4 //x2=18.415 //y2=5.155
cc_568 ( N_VDD_c_478_p N_noxref_10_c_2235_n ) capacitor c=0.00198565f \
 //x=19.07 //y=7.4 //x2=18.415 //y2=5.155
cc_569 ( N_VDD_M41_noxref_d N_noxref_10_c_2235_n ) capacitor c=0.0112985f \
 //x=18.015 //y=5.02 //x2=18.415 //y2=5.155
cc_570 ( N_VDD_c_314_n N_noxref_10_c_2239_n ) capacitor c=0.042763f //x=19.24 \
 //y=7.4 //x2=18.5 //y2=4.07
cc_571 ( N_VDD_c_310_n N_noxref_10_c_2212_n ) capacitor c=9.3395e-19 //x=28.12 \
 //y=7.4 //x2=27.38 //y2=2.08
cc_572 ( N_VDD_c_312_n N_noxref_10_c_2241_n ) capacitor c=5.93454e-19 //x=9.62 \
 //y=7.4 //x2=8.135 //y2=4.07
cc_573 ( N_VDD_c_425_p N_noxref_10_M28_noxref_g ) capacitor c=0.00675175f \
 //x=8.455 //y=7.4 //x2=7.88 //y2=6.02
cc_574 ( N_VDD_M27_noxref_d N_noxref_10_M28_noxref_g ) capacitor c=0.015318f \
 //x=7.515 //y=5.02 //x2=7.88 //y2=6.02
cc_575 ( N_VDD_c_425_p N_noxref_10_M29_noxref_g ) capacitor c=0.00675379f \
 //x=8.455 //y=7.4 //x2=8.32 //y2=6.02
cc_576 ( N_VDD_M29_noxref_d N_noxref_10_M29_noxref_g ) capacitor c=0.0394719f \
 //x=8.395 //y=5.02 //x2=8.32 //y2=6.02
cc_577 ( N_VDD_c_372_p N_noxref_10_M34_noxref_g ) capacitor c=0.00675175f \
 //x=13.265 //y=7.4 //x2=12.69 //y2=6.02
cc_578 ( N_VDD_M33_noxref_d N_noxref_10_M34_noxref_g ) capacitor c=0.015318f \
 //x=12.325 //y=5.02 //x2=12.69 //y2=6.02
cc_579 ( N_VDD_c_372_p N_noxref_10_M35_noxref_g ) capacitor c=0.00675379f \
 //x=13.265 //y=7.4 //x2=13.13 //y2=6.02
cc_580 ( N_VDD_M35_noxref_d N_noxref_10_M35_noxref_g ) capacitor c=0.0394719f \
 //x=13.205 //y=5.02 //x2=13.13 //y2=6.02
cc_581 ( N_VDD_c_588_p N_noxref_10_M52_noxref_g ) capacitor c=0.00675175f \
 //x=27.695 //y=7.4 //x2=27.12 //y2=6.02
cc_582 ( N_VDD_M51_noxref_d N_noxref_10_M52_noxref_g ) capacitor c=0.015318f \
 //x=26.755 //y=5.02 //x2=27.12 //y2=6.02
cc_583 ( N_VDD_c_588_p N_noxref_10_M53_noxref_g ) capacitor c=0.00675379f \
 //x=27.695 //y=7.4 //x2=27.56 //y2=6.02
cc_584 ( N_VDD_M53_noxref_d N_noxref_10_M53_noxref_g ) capacitor c=0.0394719f \
 //x=27.635 //y=5.02 //x2=27.56 //y2=6.02
cc_585 ( N_VDD_c_316_p N_noxref_10_M36_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=15.815 //y2=5.02
cc_586 ( N_VDD_c_382_p N_noxref_10_M36_noxref_d ) capacitor c=0.014035f \
 //x=16.315 //y=7.4 //x2=15.815 //y2=5.02
cc_587 ( N_VDD_M37_noxref_d N_noxref_10_M36_noxref_d ) capacitor c=0.0664752f \
 //x=16.255 //y=5.02 //x2=15.815 //y2=5.02
cc_588 ( N_VDD_c_316_p N_noxref_10_M38_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=16.695 //y2=5.02
cc_589 ( N_VDD_c_411_p N_noxref_10_M38_noxref_d ) capacitor c=0.014035f \
 //x=17.195 //y=7.4 //x2=16.695 //y2=5.02
cc_590 ( N_VDD_c_314_n N_noxref_10_M38_noxref_d ) capacitor c=4.9285e-19 \
 //x=19.24 //y=7.4 //x2=16.695 //y2=5.02
cc_591 ( N_VDD_M36_noxref_s N_noxref_10_M38_noxref_d ) capacitor c=0.00130656f \
 //x=15.385 //y=5.02 //x2=16.695 //y2=5.02
cc_592 ( N_VDD_M37_noxref_d N_noxref_10_M38_noxref_d ) capacitor c=0.0664752f \
 //x=16.255 //y=5.02 //x2=16.695 //y2=5.02
cc_593 ( N_VDD_M39_noxref_d N_noxref_10_M38_noxref_d ) capacitor c=0.0664752f \
 //x=17.135 //y=5.02 //x2=16.695 //y2=5.02
cc_594 ( N_VDD_c_316_p N_noxref_10_M40_noxref_d ) capacitor c=0.00274449f \
 //x=28.12 //y=7.4 //x2=17.575 //y2=5.02
cc_595 ( N_VDD_c_493_p N_noxref_10_M40_noxref_d ) capacitor c=0.0140295f \
 //x=18.075 //y=7.4 //x2=17.575 //y2=5.02
cc_596 ( N_VDD_c_314_n N_noxref_10_M40_noxref_d ) capacitor c=0.00939849f \
 //x=19.24 //y=7.4 //x2=17.575 //y2=5.02
cc_597 ( N_VDD_M39_noxref_d N_noxref_10_M40_noxref_d ) capacitor c=0.0664752f \
 //x=17.135 //y=5.02 //x2=17.575 //y2=5.02
cc_598 ( N_VDD_M41_noxref_d N_noxref_10_M40_noxref_d ) capacitor c=0.0664752f \
 //x=18.015 //y=5.02 //x2=17.575 //y2=5.02
cc_599 ( N_VDD_M42_noxref_s N_noxref_10_M40_noxref_d ) capacitor c=3.57641e-19 \
 //x=20.195 //y=5.02 //x2=17.575 //y2=5.02
cc_600 ( N_VDD_c_316_p N_Q_c_2549_n ) capacitor c=0.0226671f //x=28.12 //y=7.4 \
 //x2=28.005 //y2=3.7
cc_601 ( N_VDD_c_310_n Q ) capacitor c=0.0459745f //x=28.12 //y=7.4 //x2=28.12 \
 //y2=2.22
cc_602 ( N_VDD_c_315_n N_Q_c_2550_n ) capacitor c=0.00114628f //x=24.05 \
 //y=7.4 //x2=22.57 //y2=2.08
cc_603 ( N_VDD_c_316_p N_Q_c_2556_n ) capacitor c=0.004515f //x=28.12 //y=7.4 \
 //x2=26.375 //y2=5.155
cc_604 ( N_VDD_c_519_p N_Q_c_2556_n ) capacitor c=4.32228e-19 //x=25.935 \
 //y=7.4 //x2=26.375 //y2=5.155
cc_605 ( N_VDD_c_548_p N_Q_c_2556_n ) capacitor c=4.32228e-19 //x=26.815 \
 //y=7.4 //x2=26.375 //y2=5.155
cc_606 ( N_VDD_M49_noxref_d N_Q_c_2556_n ) capacitor c=0.0115147f //x=25.875 \
 //y=5.02 //x2=26.375 //y2=5.155
cc_607 ( N_VDD_c_315_n N_Q_c_2560_n ) capacitor c=0.00863585f //x=24.05 \
 //y=7.4 //x2=25.665 //y2=5.155
cc_608 ( N_VDD_M48_noxref_s N_Q_c_2560_n ) capacitor c=0.0831083f //x=25.005 \
 //y=5.02 //x2=25.665 //y2=5.155
cc_609 ( N_VDD_c_316_p N_Q_c_2562_n ) capacitor c=0.00448996f //x=28.12 \
 //y=7.4 //x2=27.255 //y2=5.155
cc_610 ( N_VDD_c_548_p N_Q_c_2562_n ) capacitor c=4.32228e-19 //x=26.815 \
 //y=7.4 //x2=27.255 //y2=5.155
cc_611 ( N_VDD_c_588_p N_Q_c_2562_n ) capacitor c=4.32228e-19 //x=27.695 \
 //y=7.4 //x2=27.255 //y2=5.155
cc_612 ( N_VDD_M51_noxref_d N_Q_c_2562_n ) capacitor c=0.0115147f //x=26.755 \
 //y=5.02 //x2=27.255 //y2=5.155
cc_613 ( N_VDD_c_316_p N_Q_c_2566_n ) capacitor c=0.00448978f //x=28.12 \
 //y=7.4 //x2=28.035 //y2=5.155
cc_614 ( N_VDD_c_588_p N_Q_c_2566_n ) capacitor c=7.40594e-19 //x=27.695 \
 //y=7.4 //x2=28.035 //y2=5.155
cc_615 ( N_VDD_c_310_n N_Q_c_2566_n ) capacitor c=0.00179956f //x=28.12 \
 //y=7.4 //x2=28.035 //y2=5.155
cc_616 ( N_VDD_M53_noxref_d N_Q_c_2566_n ) capacitor c=0.0116565f //x=27.635 \
 //y=5.02 //x2=28.035 //y2=5.155
cc_617 ( N_VDD_c_510_p N_Q_M46_noxref_g ) capacitor c=0.00675175f //x=22.885 \
 //y=7.4 //x2=22.31 //y2=6.02
cc_618 ( N_VDD_M45_noxref_d N_Q_M46_noxref_g ) capacitor c=0.015318f \
 //x=21.945 //y=5.02 //x2=22.31 //y2=6.02
cc_619 ( N_VDD_c_510_p N_Q_M47_noxref_g ) capacitor c=0.00675379f //x=22.885 \
 //y=7.4 //x2=22.75 //y2=6.02
cc_620 ( N_VDD_M47_noxref_d N_Q_M47_noxref_g ) capacitor c=0.0394719f \
 //x=22.825 //y=5.02 //x2=22.75 //y2=6.02
cc_621 ( N_VDD_c_316_p N_Q_M48_noxref_d ) capacitor c=0.00285091f //x=28.12 \
 //y=7.4 //x2=25.435 //y2=5.02
cc_622 ( N_VDD_c_519_p N_Q_M48_noxref_d ) capacitor c=0.0141016f //x=25.935 \
 //y=7.4 //x2=25.435 //y2=5.02
cc_623 ( N_VDD_M49_noxref_d N_Q_M48_noxref_d ) capacitor c=0.0664752f \
 //x=25.875 //y=5.02 //x2=25.435 //y2=5.02
cc_624 ( N_VDD_c_316_p N_Q_M50_noxref_d ) capacitor c=0.00285091f //x=28.12 \
 //y=7.4 //x2=26.315 //y2=5.02
cc_625 ( N_VDD_c_548_p N_Q_M50_noxref_d ) capacitor c=0.0141016f //x=26.815 \
 //y=7.4 //x2=26.315 //y2=5.02
cc_626 ( N_VDD_c_310_n N_Q_M50_noxref_d ) capacitor c=4.9285e-19 //x=28.12 \
 //y=7.4 //x2=26.315 //y2=5.02
cc_627 ( N_VDD_M48_noxref_s N_Q_M50_noxref_d ) capacitor c=0.00130656f \
 //x=25.005 //y=5.02 //x2=26.315 //y2=5.02
cc_628 ( N_VDD_M49_noxref_d N_Q_M50_noxref_d ) capacitor c=0.0664752f \
 //x=25.875 //y=5.02 //x2=26.315 //y2=5.02
cc_629 ( N_VDD_M51_noxref_d N_Q_M50_noxref_d ) capacitor c=0.0664752f \
 //x=26.755 //y=5.02 //x2=26.315 //y2=5.02
cc_630 ( N_VDD_c_316_p N_Q_M52_noxref_d ) capacitor c=0.00284366f //x=28.12 \
 //y=7.4 //x2=27.195 //y2=5.02
cc_631 ( N_VDD_c_588_p N_Q_M52_noxref_d ) capacitor c=0.0138002f //x=27.695 \
 //y=7.4 //x2=27.195 //y2=5.02
cc_632 ( N_VDD_c_310_n N_Q_M52_noxref_d ) capacitor c=0.00963505f //x=28.12 \
 //y=7.4 //x2=27.195 //y2=5.02
cc_633 ( N_VDD_M51_noxref_d N_Q_M52_noxref_d ) capacitor c=0.0664752f \
 //x=26.755 //y=5.02 //x2=27.195 //y2=5.02
cc_634 ( N_VDD_M53_noxref_d N_Q_M52_noxref_d ) capacitor c=0.0664752f \
 //x=27.635 //y=5.02 //x2=27.195 //y2=5.02
cc_635 ( N_VDD_c_316_p N_D_c_2706_n ) capacitor c=0.00112336f //x=28.12 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_636 ( N_VDD_c_309_n N_D_c_2706_n ) capacitor c=0.0165592f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_637 ( N_VDD_M18_noxref_s N_D_c_2706_n ) capacitor c=0.0130213f //x=0.955 \
 //y=5.02 //x2=1.11 //y2=2.08
cc_638 ( N_VDD_c_317_p N_D_M18_noxref_g ) capacitor c=0.00749687f //x=1.885 \
 //y=7.4 //x2=1.31 //y2=6.02
cc_639 ( N_VDD_M18_noxref_s N_D_M18_noxref_g ) capacitor c=0.0477201f \
 //x=0.955 //y=5.02 //x2=1.31 //y2=6.02
cc_640 ( N_VDD_c_317_p N_D_M19_noxref_g ) capacitor c=0.00675175f //x=1.885 \
 //y=7.4 //x2=1.75 //y2=6.02
cc_641 ( N_VDD_M19_noxref_d N_D_M19_noxref_g ) capacitor c=0.015318f //x=1.825 \
 //y=5.02 //x2=1.75 //y2=6.02
cc_642 ( N_VDD_c_309_n N_D_c_2724_n ) capacitor c=0.00757682f //x=0.74 //y=7.4 \
 //x2=1.385 //y2=4.79
cc_643 ( N_VDD_M18_noxref_s N_D_c_2724_n ) capacitor c=0.00442959f //x=0.955 \
 //y=5.02 //x2=1.385 //y2=4.79
cc_644 ( N_noxref_3_c_656_n N_noxref_4_c_955_n ) capacitor c=0.00556843f \
 //x=10.615 //y=2.965 //x2=13.805 //y2=2.96
cc_645 ( N_noxref_3_M31_noxref_g N_noxref_4_c_916_n ) capacitor c=0.0168349f \
 //x=11.37 //y=6.02 //x2=11.945 //y2=5.155
cc_646 ( N_noxref_3_M30_noxref_g N_noxref_4_c_920_n ) capacitor c=0.0213876f \
 //x=10.93 //y=6.02 //x2=11.235 //y2=5.155
cc_647 ( N_noxref_3_c_736_p N_noxref_4_c_920_n ) capacitor c=0.00428486f \
 //x=11.295 //y=4.79 //x2=11.235 //y2=5.155
cc_648 ( N_noxref_3_M31_noxref_g N_noxref_4_M30_noxref_d ) capacitor \
 c=0.0180032f //x=11.37 //y=6.02 //x2=11.005 //y2=5.02
cc_649 ( N_noxref_3_c_656_n N_CLK_c_1062_n ) capacitor c=0.33849f //x=10.615 \
 //y=2.965 //x2=16.535 //y2=3.33
cc_650 ( N_noxref_3_c_663_n N_CLK_c_1062_n ) capacitor c=0.0216421f //x=10.73 \
 //y=2.08 //x2=16.535 //y2=3.33
cc_651 ( N_noxref_3_c_656_n N_CLK_c_1079_n ) capacitor c=0.0294585f //x=10.615 \
 //y=2.965 //x2=7.145 //y2=3.33
cc_652 ( N_noxref_3_c_662_n N_CLK_c_1079_n ) capacitor c=0.00526349f //x=5.92 \
 //y=2.08 //x2=7.145 //y2=3.33
cc_653 ( N_noxref_3_c_656_n N_CLK_c_1063_n ) capacitor c=0.0253594f //x=10.615 \
 //y=2.965 //x2=7.03 //y2=2.08
cc_654 ( N_noxref_3_c_660_n N_CLK_c_1063_n ) capacitor c=9.95819e-19 //x=6.035 \
 //y=2.965 //x2=7.03 //y2=2.08
cc_655 ( N_noxref_3_c_699_n N_CLK_c_1063_n ) capacitor c=5.06912e-19 //x=4.07 \
 //y=2.965 //x2=7.03 //y2=2.08
cc_656 ( N_noxref_3_c_662_n N_CLK_c_1063_n ) capacitor c=0.0487554f //x=5.92 \
 //y=2.08 //x2=7.03 //y2=2.08
cc_657 ( N_noxref_3_c_668_n N_CLK_c_1063_n ) capacitor c=0.00238338f //x=5.62 \
 //y=1.915 //x2=7.03 //y2=2.08
cc_658 ( N_noxref_3_c_747_p N_CLK_c_1063_n ) capacitor c=0.00147352f //x=6.485 \
 //y=4.79 //x2=7.03 //y2=2.08
cc_659 ( N_noxref_3_c_714_n N_CLK_c_1063_n ) capacitor c=0.00142741f //x=6.195 \
 //y=4.79 //x2=7.03 //y2=2.08
cc_660 ( N_noxref_3_M24_noxref_g N_CLK_M26_noxref_g ) capacitor c=0.0105869f \
 //x=6.12 //y=6.02 //x2=7 //y2=6.02
cc_661 ( N_noxref_3_M25_noxref_g N_CLK_M26_noxref_g ) capacitor c=0.10632f \
 //x=6.56 //y=6.02 //x2=7 //y2=6.02
cc_662 ( N_noxref_3_M25_noxref_g N_CLK_M27_noxref_g ) capacitor c=0.0101598f \
 //x=6.56 //y=6.02 //x2=7.44 //y2=6.02
cc_663 ( N_noxref_3_c_664_n N_CLK_c_1091_n ) capacitor c=5.72482e-19 //x=5.62 \
 //y=0.875 //x2=6.595 //y2=0.91
cc_664 ( N_noxref_3_c_666_n N_CLK_c_1091_n ) capacitor c=0.00149976f //x=5.62 \
 //y=1.22 //x2=6.595 //y2=0.91
cc_665 ( N_noxref_3_c_671_n N_CLK_c_1091_n ) capacitor c=0.0160123f //x=6.15 \
 //y=0.875 //x2=6.595 //y2=0.91
cc_666 ( N_noxref_3_c_667_n N_CLK_c_1094_n ) capacitor c=0.00111227f //x=5.62 \
 //y=1.53 //x2=6.595 //y2=1.22
cc_667 ( N_noxref_3_c_673_n N_CLK_c_1094_n ) capacitor c=0.0124075f //x=6.15 \
 //y=1.22 //x2=6.595 //y2=1.22
cc_668 ( N_noxref_3_c_671_n N_CLK_c_1096_n ) capacitor c=0.00103227f //x=6.15 \
 //y=0.875 //x2=7.12 //y2=0.91
cc_669 ( N_noxref_3_c_673_n N_CLK_c_1097_n ) capacitor c=0.0010154f //x=6.15 \
 //y=1.22 //x2=7.12 //y2=1.22
cc_670 ( N_noxref_3_c_673_n N_CLK_c_1098_n ) capacitor c=9.23422e-19 //x=6.15 \
 //y=1.22 //x2=7.12 //y2=1.45
cc_671 ( N_noxref_3_c_656_n N_CLK_c_1099_n ) capacitor c=0.00231387f \
 //x=10.615 //y=2.965 //x2=7.12 //y2=1.915
cc_672 ( N_noxref_3_c_662_n N_CLK_c_1099_n ) capacitor c=0.00231304f //x=5.92 \
 //y=2.08 //x2=7.12 //y2=1.915
cc_673 ( N_noxref_3_c_668_n N_CLK_c_1099_n ) capacitor c=0.00964411f //x=5.62 \
 //y=1.915 //x2=7.12 //y2=1.915
cc_674 ( N_noxref_3_c_662_n N_CLK_c_1102_n ) capacitor c=0.00183762f //x=5.92 \
 //y=2.08 //x2=7.03 //y2=4.7
cc_675 ( N_noxref_3_c_747_p N_CLK_c_1102_n ) capacitor c=0.0168581f //x=6.485 \
 //y=4.79 //x2=7.03 //y2=4.7
cc_676 ( N_noxref_3_c_714_n N_CLK_c_1102_n ) capacitor c=0.00484466f //x=6.195 \
 //y=4.79 //x2=7.03 //y2=4.7
cc_677 ( N_noxref_3_c_651_n N_noxref_6_c_1253_n ) capacitor c=0.0743044f \
 //x=5.805 //y=2.965 //x2=8.765 //y2=3.7
cc_678 ( N_noxref_3_c_655_n N_noxref_6_c_1253_n ) capacitor c=0.0136944f \
 //x=4.185 //y=2.965 //x2=8.765 //y2=3.7
cc_679 ( N_noxref_3_c_656_n N_noxref_6_c_1253_n ) capacitor c=0.053052f \
 //x=10.615 //y=2.965 //x2=8.765 //y2=3.7
cc_680 ( N_noxref_3_c_660_n N_noxref_6_c_1253_n ) capacitor c=0.0123989f \
 //x=6.035 //y=2.965 //x2=8.765 //y2=3.7
cc_681 ( N_noxref_3_c_770_p N_noxref_6_c_1253_n ) capacitor c=0.0042996f \
 //x=3.67 //y=1.665 //x2=8.765 //y2=3.7
cc_682 ( N_noxref_3_c_699_n N_noxref_6_c_1253_n ) capacitor c=0.0237485f \
 //x=4.07 //y=2.965 //x2=8.765 //y2=3.7
cc_683 ( N_noxref_3_c_662_n N_noxref_6_c_1253_n ) capacitor c=0.024705f \
 //x=5.92 //y=2.08 //x2=8.765 //y2=3.7
cc_684 ( N_noxref_3_c_699_n N_noxref_6_c_1254_n ) capacitor c=0.00179385f \
 //x=4.07 //y=2.965 //x2=3.445 //y2=3.7
cc_685 ( N_noxref_3_c_656_n N_noxref_6_c_1255_n ) capacitor c=0.0117239f \
 //x=10.615 //y=2.965 //x2=20.235 //y2=3.7
cc_686 ( N_noxref_3_c_663_n N_noxref_6_c_1255_n ) capacitor c=0.0197627f \
 //x=10.73 //y=2.08 //x2=20.235 //y2=3.7
cc_687 ( N_noxref_3_c_656_n N_noxref_6_c_1325_n ) capacitor c=4.83387e-19 \
 //x=10.615 //y=2.965 //x2=8.995 //y2=3.7
cc_688 ( N_noxref_3_c_663_n N_noxref_6_c_1325_n ) capacitor c=7.01366e-19 \
 //x=10.73 //y=2.08 //x2=8.995 //y2=3.7
cc_689 ( N_noxref_3_c_655_n N_noxref_6_c_1256_n ) capacitor c=0.00687545f \
 //x=4.185 //y=2.965 //x2=3.33 //y2=2.08
cc_690 ( N_noxref_3_c_699_n N_noxref_6_c_1256_n ) capacitor c=0.0857427f \
 //x=4.07 //y=2.965 //x2=3.33 //y2=2.08
cc_691 ( N_noxref_3_c_662_n N_noxref_6_c_1256_n ) capacitor c=0.00105582f \
 //x=5.92 //y=2.08 //x2=3.33 //y2=2.08
cc_692 ( N_noxref_3_c_781_p N_noxref_6_c_1256_n ) capacitor c=0.016476f \
 //x=3.29 //y=5.155 //x2=3.33 //y2=2.08
cc_693 ( N_noxref_3_M25_noxref_g N_noxref_6_c_1272_n ) capacitor c=0.0168349f \
 //x=6.56 //y=6.02 //x2=7.135 //y2=5.155
cc_694 ( N_noxref_3_c_695_n N_noxref_6_c_1276_n ) capacitor c=3.10026e-19 \
 //x=3.985 //y=5.155 //x2=6.425 //y2=5.155
cc_695 ( N_noxref_3_M24_noxref_g N_noxref_6_c_1276_n ) capacitor c=0.0213876f \
 //x=6.12 //y=6.02 //x2=6.425 //y2=5.155
cc_696 ( N_noxref_3_c_747_p N_noxref_6_c_1276_n ) capacitor c=0.00428486f \
 //x=6.485 //y=4.79 //x2=6.425 //y2=5.155
cc_697 ( N_noxref_3_c_656_n N_noxref_6_c_1335_n ) capacitor c=0.00835258f \
 //x=10.615 //y=2.965 //x2=8.48 //y2=1.665
cc_698 ( N_noxref_3_c_656_n N_noxref_6_c_1286_n ) capacitor c=0.024355f \
 //x=10.615 //y=2.965 //x2=8.88 //y2=3.7
cc_699 ( N_noxref_3_c_663_n N_noxref_6_c_1286_n ) capacitor c=0.0109419f \
 //x=10.73 //y=2.08 //x2=8.88 //y2=3.7
cc_700 ( N_noxref_3_c_691_n N_noxref_6_M22_noxref_g ) capacitor c=0.01736f \
 //x=3.205 //y=5.155 //x2=3.07 //y2=6.02
cc_701 ( N_noxref_3_M22_noxref_d N_noxref_6_M22_noxref_g ) capacitor \
 c=0.0180032f //x=3.145 //y=5.02 //x2=3.07 //y2=6.02
cc_702 ( N_noxref_3_c_695_n N_noxref_6_M23_noxref_g ) capacitor c=0.0194981f \
 //x=3.985 //y=5.155 //x2=3.51 //y2=6.02
cc_703 ( N_noxref_3_M22_noxref_d N_noxref_6_M23_noxref_g ) capacitor \
 c=0.0194246f //x=3.145 //y=5.02 //x2=3.51 //y2=6.02
cc_704 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1342_n ) capacitor c=0.00217566f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=0.915
cc_705 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1343_n ) capacitor c=0.0034598f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=1.26
cc_706 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1344_n ) capacitor c=0.00544291f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=1.57
cc_707 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1345_n ) capacitor c=0.00241102f \
 //x=3.395 //y=0.915 //x2=3.695 //y2=0.76
cc_708 ( N_noxref_3_c_661_n N_noxref_6_c_1346_n ) capacitor c=0.00359704f \
 //x=3.985 //y=1.665 //x2=3.695 //y2=1.415
cc_709 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1346_n ) capacitor c=0.0140297f \
 //x=3.395 //y=0.915 //x2=3.695 //y2=1.415
cc_710 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1348_n ) capacitor c=0.00219619f \
 //x=3.395 //y=0.915 //x2=3.85 //y2=0.915
cc_711 ( N_noxref_3_c_661_n N_noxref_6_c_1349_n ) capacitor c=0.00457401f \
 //x=3.985 //y=1.665 //x2=3.85 //y2=1.26
cc_712 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1349_n ) capacitor c=0.00603828f \
 //x=3.395 //y=0.915 //x2=3.85 //y2=1.26
cc_713 ( N_noxref_3_c_699_n N_noxref_6_c_1351_n ) capacitor c=0.00877984f \
 //x=4.07 //y=2.965 //x2=3.33 //y2=2.08
cc_714 ( N_noxref_3_c_699_n N_noxref_6_c_1352_n ) capacitor c=0.00283672f \
 //x=4.07 //y=2.965 //x2=3.33 //y2=1.915
cc_715 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1352_n ) capacitor c=0.00661782f \
 //x=3.395 //y=0.915 //x2=3.33 //y2=1.915
cc_716 ( N_noxref_3_c_695_n N_noxref_6_c_1354_n ) capacitor c=0.00201851f \
 //x=3.985 //y=5.155 //x2=3.33 //y2=4.7
cc_717 ( N_noxref_3_c_699_n N_noxref_6_c_1354_n ) capacitor c=0.013693f \
 //x=4.07 //y=2.965 //x2=3.33 //y2=4.7
cc_718 ( N_noxref_3_c_781_p N_noxref_6_c_1354_n ) capacitor c=0.00475601f \
 //x=3.29 //y=5.155 //x2=3.33 //y2=4.7
cc_719 ( N_noxref_3_M25_noxref_g N_noxref_6_M24_noxref_d ) capacitor \
 c=0.0180032f //x=6.56 //y=6.02 //x2=6.195 //y2=5.02
cc_720 ( N_noxref_3_c_651_n N_RN_c_1514_n ) capacitor c=0.00385587f //x=5.805 \
 //y=2.965 //x2=17.645 //y2=4.44
cc_721 ( N_noxref_3_c_655_n N_RN_c_1514_n ) capacitor c=3.67454e-19 //x=4.185 \
 //y=2.965 //x2=17.645 //y2=4.44
cc_722 ( N_noxref_3_c_656_n N_RN_c_1514_n ) capacitor c=0.00397392f //x=10.615 \
 //y=2.965 //x2=17.645 //y2=4.44
cc_723 ( N_noxref_3_c_660_n N_RN_c_1514_n ) capacitor c=2.47225e-19 //x=6.035 \
 //y=2.965 //x2=17.645 //y2=4.44
cc_724 ( N_noxref_3_c_695_n N_RN_c_1514_n ) capacitor c=0.0183122f //x=3.985 \
 //y=5.155 //x2=17.645 //y2=4.44
cc_725 ( N_noxref_3_c_699_n N_RN_c_1514_n ) capacitor c=0.023368f //x=4.07 \
 //y=2.965 //x2=17.645 //y2=4.44
cc_726 ( N_noxref_3_c_662_n N_RN_c_1514_n ) capacitor c=0.0232115f //x=5.92 \
 //y=2.08 //x2=17.645 //y2=4.44
cc_727 ( N_noxref_3_c_663_n N_RN_c_1514_n ) capacitor c=0.0208709f //x=10.73 \
 //y=2.08 //x2=17.645 //y2=4.44
cc_728 ( N_noxref_3_c_817_p N_RN_c_1514_n ) capacitor c=0.0306894f //x=2.41 \
 //y=5.155 //x2=17.645 //y2=4.44
cc_729 ( N_noxref_3_c_714_n N_RN_c_1514_n ) capacitor c=0.0169569f //x=6.195 \
 //y=4.79 //x2=17.645 //y2=4.44
cc_730 ( N_noxref_3_c_716_n N_RN_c_1514_n ) capacitor c=0.0166984f //x=11.005 \
 //y=4.79 //x2=17.645 //y2=4.44
cc_731 ( N_noxref_3_c_685_n N_RN_c_1515_n ) capacitor c=0.00325717f //x=2.325 \
 //y=5.155 //x2=2.335 //y2=4.44
cc_732 ( N_noxref_3_c_685_n N_RN_c_1516_n ) capacitor c=0.0143918f //x=2.325 \
 //y=5.155 //x2=2.22 //y2=2.08
cc_733 ( N_noxref_3_c_699_n N_RN_c_1516_n ) capacitor c=0.0032755f //x=4.07 \
 //y=2.965 //x2=2.22 //y2=2.08
cc_734 ( N_noxref_3_c_685_n N_RN_M20_noxref_g ) capacitor c=0.016514f \
 //x=2.325 //y=5.155 //x2=2.19 //y2=6.02
cc_735 ( N_noxref_3_M20_noxref_d N_RN_M20_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.19 //y2=6.02
cc_736 ( N_noxref_3_c_691_n N_RN_M21_noxref_g ) capacitor c=0.01736f //x=3.205 \
 //y=5.155 //x2=2.63 //y2=6.02
cc_737 ( N_noxref_3_M20_noxref_d N_RN_M21_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.63 //y2=6.02
cc_738 ( N_noxref_3_c_817_p N_RN_c_1578_n ) capacitor c=0.00426767f //x=2.41 \
 //y=5.155 //x2=2.555 //y2=4.79
cc_739 ( N_noxref_3_c_685_n N_RN_c_1579_n ) capacitor c=0.00322046f //x=2.325 \
 //y=5.155 //x2=2.22 //y2=4.7
cc_740 ( N_noxref_3_c_663_n N_SN_c_1990_n ) capacitor c=0.00526349f //x=10.73 \
 //y=2.08 //x2=11.955 //y2=2.59
cc_741 ( N_noxref_3_c_656_n N_SN_c_1991_n ) capacitor c=0.00316035f //x=10.615 \
 //y=2.965 //x2=11.84 //y2=2.08
cc_742 ( N_noxref_3_c_663_n N_SN_c_1991_n ) capacitor c=0.0456411f //x=10.73 \
 //y=2.08 //x2=11.84 //y2=2.08
cc_743 ( N_noxref_3_c_678_n N_SN_c_1991_n ) capacitor c=0.00238338f //x=10.43 \
 //y=1.915 //x2=11.84 //y2=2.08
cc_744 ( N_noxref_3_c_736_p N_SN_c_1991_n ) capacitor c=0.00147352f //x=11.295 \
 //y=4.79 //x2=11.84 //y2=2.08
cc_745 ( N_noxref_3_c_716_n N_SN_c_1991_n ) capacitor c=0.00142741f //x=11.005 \
 //y=4.79 //x2=11.84 //y2=2.08
cc_746 ( N_noxref_3_M30_noxref_g N_SN_M32_noxref_g ) capacitor c=0.0105869f \
 //x=10.93 //y=6.02 //x2=11.81 //y2=6.02
cc_747 ( N_noxref_3_M31_noxref_g N_SN_M32_noxref_g ) capacitor c=0.10632f \
 //x=11.37 //y=6.02 //x2=11.81 //y2=6.02
cc_748 ( N_noxref_3_M31_noxref_g N_SN_M33_noxref_g ) capacitor c=0.0101598f \
 //x=11.37 //y=6.02 //x2=12.25 //y2=6.02
cc_749 ( N_noxref_3_c_674_n N_SN_c_2014_n ) capacitor c=5.72482e-19 //x=10.43 \
 //y=0.875 //x2=11.405 //y2=0.91
cc_750 ( N_noxref_3_c_676_n N_SN_c_2014_n ) capacitor c=0.00149976f //x=10.43 \
 //y=1.22 //x2=11.405 //y2=0.91
cc_751 ( N_noxref_3_c_681_n N_SN_c_2014_n ) capacitor c=0.0160123f //x=10.96 \
 //y=0.875 //x2=11.405 //y2=0.91
cc_752 ( N_noxref_3_c_677_n N_SN_c_2017_n ) capacitor c=0.00111227f //x=10.43 \
 //y=1.53 //x2=11.405 //y2=1.22
cc_753 ( N_noxref_3_c_683_n N_SN_c_2017_n ) capacitor c=0.0124075f //x=10.96 \
 //y=1.22 //x2=11.405 //y2=1.22
cc_754 ( N_noxref_3_c_681_n N_SN_c_2019_n ) capacitor c=0.00103227f //x=10.96 \
 //y=0.875 //x2=11.93 //y2=0.91
cc_755 ( N_noxref_3_c_683_n N_SN_c_2020_n ) capacitor c=0.0010154f //x=10.96 \
 //y=1.22 //x2=11.93 //y2=1.22
cc_756 ( N_noxref_3_c_683_n N_SN_c_2021_n ) capacitor c=9.23422e-19 //x=10.96 \
 //y=1.22 //x2=11.93 //y2=1.45
cc_757 ( N_noxref_3_c_663_n N_SN_c_2022_n ) capacitor c=0.00231304f //x=10.73 \
 //y=2.08 //x2=11.93 //y2=1.915
cc_758 ( N_noxref_3_c_678_n N_SN_c_2022_n ) capacitor c=0.00964411f //x=10.43 \
 //y=1.915 //x2=11.93 //y2=1.915
cc_759 ( N_noxref_3_c_663_n N_SN_c_2024_n ) capacitor c=0.00183762f //x=10.73 \
 //y=2.08 //x2=11.84 //y2=4.7
cc_760 ( N_noxref_3_c_736_p N_SN_c_2024_n ) capacitor c=0.0168581f //x=11.295 \
 //y=4.79 //x2=11.84 //y2=4.7
cc_761 ( N_noxref_3_c_716_n N_SN_c_2024_n ) capacitor c=0.00484466f //x=11.005 \
 //y=4.79 //x2=11.84 //y2=4.7
cc_762 ( N_noxref_3_c_663_n N_noxref_10_c_2214_n ) capacitor c=0.0194977f \
 //x=10.73 //y=2.08 //x2=12.835 //y2=4.07
cc_763 ( N_noxref_3_c_656_n N_noxref_10_c_2209_n ) capacitor c=0.0224183f \
 //x=10.615 //y=2.965 //x2=8.14 //y2=2.08
cc_764 ( N_noxref_3_c_662_n N_noxref_10_c_2209_n ) capacitor c=0.0010353f \
 //x=5.92 //y=2.08 //x2=8.14 //y2=2.08
cc_765 ( N_noxref_3_c_663_n N_noxref_10_c_2209_n ) capacitor c=6.87018e-19 \
 //x=10.73 //y=2.08 //x2=8.14 //y2=2.08
cc_766 ( N_noxref_3_c_663_n N_noxref_10_c_2210_n ) capacitor c=0.00128592f \
 //x=10.73 //y=2.08 //x2=12.95 //y2=2.08
cc_767 ( N_noxref_3_c_662_n N_noxref_10_c_2241_n ) capacitor c=3.2187e-19 \
 //x=5.92 //y=2.08 //x2=8.135 //y2=4.07
cc_768 ( N_noxref_3_c_656_n N_noxref_10_c_2275_n ) capacitor c=0.0018253f \
 //x=10.615 //y=2.965 //x2=8.14 //y2=2.08
cc_769 ( N_noxref_3_c_689_n N_D_M18_noxref_g ) capacitor c=0.0213876f \
 //x=1.615 //y=5.155 //x2=1.31 //y2=6.02
cc_770 ( N_noxref_3_c_685_n N_D_M19_noxref_g ) capacitor c=0.0204065f \
 //x=2.325 //y=5.155 //x2=1.75 //y2=6.02
cc_771 ( N_noxref_3_M18_noxref_d N_D_M19_noxref_g ) capacitor c=0.0180032f \
 //x=1.385 //y=5.02 //x2=1.75 //y2=6.02
cc_772 ( N_noxref_3_c_689_n N_D_c_2729_n ) capacitor c=0.00437952f //x=1.615 \
 //y=5.155 //x2=1.675 //y2=4.79
cc_773 ( N_noxref_3_M2_noxref_d N_noxref_13_M0_noxref_s ) capacitor \
 c=0.00309936f //x=3.395 //y=0.915 //x2=0.455 //y2=0.375
cc_774 ( N_noxref_3_c_661_n N_noxref_14_c_2814_n ) capacitor c=0.00467111f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_775 ( N_noxref_3_M2_noxref_d N_noxref_14_c_2814_n ) capacitor c=0.0118029f \
 //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_776 ( N_noxref_3_c_770_p N_noxref_14_c_2825_n ) capacitor c=0.0200405f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_777 ( N_noxref_3_M2_noxref_d N_noxref_14_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_778 ( N_noxref_3_c_661_n N_noxref_14_M2_noxref_s ) capacitor c=0.0205066f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_779 ( N_noxref_3_M2_noxref_d N_noxref_14_M2_noxref_s ) capacitor \
 c=0.0426368f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
cc_780 ( N_noxref_3_c_651_n N_noxref_15_c_2877_n ) capacitor c=0.00323545f \
 //x=5.805 //y=2.965 //x2=5.4 //y2=1.505
cc_781 ( N_noxref_3_c_661_n N_noxref_15_c_2877_n ) capacitor c=3.84569e-19 \
 //x=3.985 //y=1.665 //x2=5.4 //y2=1.505
cc_782 ( N_noxref_3_c_668_n N_noxref_15_c_2877_n ) capacitor c=0.0034165f \
 //x=5.62 //y=1.915 //x2=5.4 //y2=1.505
cc_783 ( N_noxref_3_c_651_n N_noxref_15_c_2861_n ) capacitor c=0.00724023f \
 //x=5.805 //y=2.965 //x2=6.285 //y2=1.59
cc_784 ( N_noxref_3_c_656_n N_noxref_15_c_2861_n ) capacitor c=0.00395948f \
 //x=10.615 //y=2.965 //x2=6.285 //y2=1.59
cc_785 ( N_noxref_3_c_660_n N_noxref_15_c_2861_n ) capacitor c=0.00158887f \
 //x=6.035 //y=2.965 //x2=6.285 //y2=1.59
cc_786 ( N_noxref_3_c_662_n N_noxref_15_c_2861_n ) capacitor c=0.0119604f \
 //x=5.92 //y=2.08 //x2=6.285 //y2=1.59
cc_787 ( N_noxref_3_c_667_n N_noxref_15_c_2861_n ) capacitor c=0.00703864f \
 //x=5.62 //y=1.53 //x2=6.285 //y2=1.59
cc_788 ( N_noxref_3_c_668_n N_noxref_15_c_2861_n ) capacitor c=0.0224281f \
 //x=5.62 //y=1.915 //x2=6.285 //y2=1.59
cc_789 ( N_noxref_3_c_670_n N_noxref_15_c_2861_n ) capacitor c=0.00708583f \
 //x=5.995 //y=1.375 //x2=6.285 //y2=1.59
cc_790 ( N_noxref_3_c_673_n N_noxref_15_c_2861_n ) capacitor c=0.00698822f \
 //x=6.15 //y=1.22 //x2=6.285 //y2=1.59
cc_791 ( N_noxref_3_c_656_n N_noxref_15_c_2888_n ) capacitor c=0.0109188f \
 //x=10.615 //y=2.965 //x2=7.255 //y2=1.59
cc_792 ( N_noxref_3_c_656_n N_noxref_15_M3_noxref_s ) capacitor c=0.00625215f \
 //x=10.615 //y=2.965 //x2=5.265 //y2=0.375
cc_793 ( N_noxref_3_c_664_n N_noxref_15_M3_noxref_s ) capacitor c=0.0327271f \
 //x=5.62 //y=0.875 //x2=5.265 //y2=0.375
cc_794 ( N_noxref_3_c_667_n N_noxref_15_M3_noxref_s ) capacitor c=7.99997e-19 \
 //x=5.62 //y=1.53 //x2=5.265 //y2=0.375
cc_795 ( N_noxref_3_c_668_n N_noxref_15_M3_noxref_s ) capacitor c=0.00122123f \
 //x=5.62 //y=1.915 //x2=5.265 //y2=0.375
cc_796 ( N_noxref_3_c_671_n N_noxref_15_M3_noxref_s ) capacitor c=0.0121427f \
 //x=6.15 //y=0.875 //x2=5.265 //y2=0.375
cc_797 ( N_noxref_3_M2_noxref_d N_noxref_15_M3_noxref_s ) capacitor \
 c=2.55333e-19 //x=3.395 //y=0.915 //x2=5.265 //y2=0.375
cc_798 ( N_noxref_3_c_656_n N_noxref_16_c_2913_n ) capacitor c=0.00382437f \
 //x=10.615 //y=2.965 //x2=7.825 //y2=0.995
cc_799 ( N_noxref_3_c_656_n N_noxref_16_c_2919_n ) capacitor c=6.56577e-19 \
 //x=10.615 //y=2.965 //x2=8.795 //y2=0.54
cc_800 ( N_noxref_3_c_656_n N_noxref_16_M5_noxref_s ) capacitor c=0.00323545f \
 //x=10.615 //y=2.965 //x2=7.775 //y2=0.375
cc_801 ( N_noxref_3_c_656_n N_noxref_17_c_2983_n ) capacitor c=0.00323545f \
 //x=10.615 //y=2.965 //x2=10.21 //y2=1.505
cc_802 ( N_noxref_3_c_678_n N_noxref_17_c_2983_n ) capacitor c=0.0034165f \
 //x=10.43 //y=1.915 //x2=10.21 //y2=1.505
cc_803 ( N_noxref_3_c_656_n N_noxref_17_c_2967_n ) capacitor c=0.00929348f \
 //x=10.615 //y=2.965 //x2=11.095 //y2=1.59
cc_804 ( N_noxref_3_c_663_n N_noxref_17_c_2967_n ) capacitor c=0.0119604f \
 //x=10.73 //y=2.08 //x2=11.095 //y2=1.59
cc_805 ( N_noxref_3_c_677_n N_noxref_17_c_2967_n ) capacitor c=0.00703864f \
 //x=10.43 //y=1.53 //x2=11.095 //y2=1.59
cc_806 ( N_noxref_3_c_678_n N_noxref_17_c_2967_n ) capacitor c=0.0224281f \
 //x=10.43 //y=1.915 //x2=11.095 //y2=1.59
cc_807 ( N_noxref_3_c_680_n N_noxref_17_c_2967_n ) capacitor c=0.00708583f \
 //x=10.805 //y=1.375 //x2=11.095 //y2=1.59
cc_808 ( N_noxref_3_c_683_n N_noxref_17_c_2967_n ) capacitor c=0.00698822f \
 //x=10.96 //y=1.22 //x2=11.095 //y2=1.59
cc_809 ( N_noxref_3_c_674_n N_noxref_17_M6_noxref_s ) capacitor c=0.0327271f \
 //x=10.43 //y=0.875 //x2=10.075 //y2=0.375
cc_810 ( N_noxref_3_c_677_n N_noxref_17_M6_noxref_s ) capacitor c=7.99997e-19 \
 //x=10.43 //y=1.53 //x2=10.075 //y2=0.375
cc_811 ( N_noxref_3_c_678_n N_noxref_17_M6_noxref_s ) capacitor c=0.00122123f \
 //x=10.43 //y=1.915 //x2=10.075 //y2=0.375
cc_812 ( N_noxref_3_c_681_n N_noxref_17_M6_noxref_s ) capacitor c=0.0121427f \
 //x=10.96 //y=0.875 //x2=10.075 //y2=0.375
cc_813 ( N_noxref_4_c_902_n N_CLK_c_1062_n ) capacitor c=0.174212f //x=15.425 \
 //y=2.96 //x2=16.535 //y2=3.33
cc_814 ( N_noxref_4_c_955_n N_CLK_c_1062_n ) capacitor c=0.0294052f //x=13.805 \
 //y=2.96 //x2=16.535 //y2=3.33
cc_815 ( N_noxref_4_c_930_n N_CLK_c_1062_n ) capacitor c=0.0205776f //x=13.69 \
 //y=2.96 //x2=16.535 //y2=3.33
cc_816 ( N_noxref_4_c_904_n N_CLK_c_1062_n ) capacitor c=0.0229269f //x=15.54 \
 //y=2.08 //x2=16.535 //y2=3.33
cc_817 ( N_noxref_4_c_902_n N_CLK_c_1064_n ) capacitor c=0.00520283f \
 //x=15.425 //y=2.96 //x2=16.65 //y2=2.08
cc_818 ( N_noxref_4_c_930_n N_CLK_c_1064_n ) capacitor c=5.24823e-19 //x=13.69 \
 //y=2.96 //x2=16.65 //y2=2.08
cc_819 ( N_noxref_4_c_904_n N_CLK_c_1064_n ) capacitor c=0.0442053f //x=15.54 \
 //y=2.08 //x2=16.65 //y2=2.08
cc_820 ( N_noxref_4_c_909_n N_CLK_c_1064_n ) capacitor c=0.00238338f //x=15.24 \
 //y=1.915 //x2=16.65 //y2=2.08
cc_821 ( N_noxref_4_c_968_p N_CLK_c_1064_n ) capacitor c=0.00147352f \
 //x=16.105 //y=4.79 //x2=16.65 //y2=2.08
cc_822 ( N_noxref_4_c_938_n N_CLK_c_1064_n ) capacitor c=0.00142741f \
 //x=15.815 //y=4.79 //x2=16.65 //y2=2.08
cc_823 ( N_noxref_4_M36_noxref_g N_CLK_M38_noxref_g ) capacitor c=0.0105869f \
 //x=15.74 //y=6.02 //x2=16.62 //y2=6.02
cc_824 ( N_noxref_4_M37_noxref_g N_CLK_M38_noxref_g ) capacitor c=0.10632f \
 //x=16.18 //y=6.02 //x2=16.62 //y2=6.02
cc_825 ( N_noxref_4_M37_noxref_g N_CLK_M39_noxref_g ) capacitor c=0.0101598f \
 //x=16.18 //y=6.02 //x2=17.06 //y2=6.02
cc_826 ( N_noxref_4_c_905_n N_CLK_c_1118_n ) capacitor c=5.72482e-19 //x=15.24 \
 //y=0.875 //x2=16.215 //y2=0.91
cc_827 ( N_noxref_4_c_907_n N_CLK_c_1118_n ) capacitor c=0.00149976f //x=15.24 \
 //y=1.22 //x2=16.215 //y2=0.91
cc_828 ( N_noxref_4_c_912_n N_CLK_c_1118_n ) capacitor c=0.0160123f //x=15.77 \
 //y=0.875 //x2=16.215 //y2=0.91
cc_829 ( N_noxref_4_c_908_n N_CLK_c_1121_n ) capacitor c=0.00111227f //x=15.24 \
 //y=1.53 //x2=16.215 //y2=1.22
cc_830 ( N_noxref_4_c_914_n N_CLK_c_1121_n ) capacitor c=0.0124075f //x=15.77 \
 //y=1.22 //x2=16.215 //y2=1.22
cc_831 ( N_noxref_4_c_912_n N_CLK_c_1123_n ) capacitor c=0.00103227f //x=15.77 \
 //y=0.875 //x2=16.74 //y2=0.91
cc_832 ( N_noxref_4_c_914_n N_CLK_c_1124_n ) capacitor c=0.0010154f //x=15.77 \
 //y=1.22 //x2=16.74 //y2=1.22
cc_833 ( N_noxref_4_c_914_n N_CLK_c_1125_n ) capacitor c=9.23422e-19 //x=15.77 \
 //y=1.22 //x2=16.74 //y2=1.45
cc_834 ( N_noxref_4_c_904_n N_CLK_c_1126_n ) capacitor c=0.00231304f //x=15.54 \
 //y=2.08 //x2=16.74 //y2=1.915
cc_835 ( N_noxref_4_c_909_n N_CLK_c_1126_n ) capacitor c=0.00964411f //x=15.24 \
 //y=1.915 //x2=16.74 //y2=1.915
cc_836 ( N_noxref_4_c_904_n N_CLK_c_1128_n ) capacitor c=0.00183762f //x=15.54 \
 //y=2.08 //x2=16.65 //y2=4.7
cc_837 ( N_noxref_4_c_968_p N_CLK_c_1128_n ) capacitor c=0.0168581f //x=16.105 \
 //y=4.79 //x2=16.65 //y2=4.7
cc_838 ( N_noxref_4_c_938_n N_CLK_c_1128_n ) capacitor c=0.00484466f \
 //x=15.815 //y=4.79 //x2=16.65 //y2=4.7
cc_839 ( N_noxref_4_c_902_n N_noxref_6_c_1255_n ) capacitor c=0.0116525f \
 //x=15.425 //y=2.96 //x2=20.235 //y2=3.7
cc_840 ( N_noxref_4_c_955_n N_noxref_6_c_1255_n ) capacitor c=7.98461e-19 \
 //x=13.805 //y=2.96 //x2=20.235 //y2=3.7
cc_841 ( N_noxref_4_c_930_n N_noxref_6_c_1255_n ) capacitor c=0.0187698f \
 //x=13.69 //y=2.96 //x2=20.235 //y2=3.7
cc_842 ( N_noxref_4_c_904_n N_noxref_6_c_1255_n ) capacitor c=0.0197889f \
 //x=15.54 //y=2.08 //x2=20.235 //y2=3.7
cc_843 ( N_noxref_4_c_920_n N_noxref_6_c_1282_n ) capacitor c=3.10026e-19 \
 //x=11.235 //y=5.155 //x2=8.795 //y2=5.155
cc_844 ( N_noxref_4_c_916_n N_RN_c_1514_n ) capacitor c=0.032141f //x=11.945 \
 //y=5.155 //x2=17.645 //y2=4.44
cc_845 ( N_noxref_4_c_920_n N_RN_c_1514_n ) capacitor c=0.0230136f //x=11.235 \
 //y=5.155 //x2=17.645 //y2=4.44
cc_846 ( N_noxref_4_c_926_n N_RN_c_1514_n ) capacitor c=0.0183122f //x=13.605 \
 //y=5.155 //x2=17.645 //y2=4.44
cc_847 ( N_noxref_4_c_930_n N_RN_c_1514_n ) capacitor c=0.0210274f //x=13.69 \
 //y=2.96 //x2=17.645 //y2=4.44
cc_848 ( N_noxref_4_c_904_n N_RN_c_1514_n ) capacitor c=0.0208709f //x=15.54 \
 //y=2.08 //x2=17.645 //y2=4.44
cc_849 ( N_noxref_4_c_938_n N_RN_c_1514_n ) capacitor c=0.0166984f //x=15.815 \
 //y=4.79 //x2=17.645 //y2=4.44
cc_850 ( N_noxref_4_c_904_n N_RN_c_1517_n ) capacitor c=0.00132243f //x=15.54 \
 //y=2.08 //x2=17.76 //y2=2.08
cc_851 ( N_noxref_4_c_902_n N_SN_c_1980_n ) capacitor c=0.172536f //x=15.425 \
 //y=2.96 //x2=26.155 //y2=2.59
cc_852 ( N_noxref_4_c_955_n N_SN_c_1980_n ) capacitor c=0.0292376f //x=13.805 \
 //y=2.96 //x2=26.155 //y2=2.59
cc_853 ( N_noxref_4_c_1000_p N_SN_c_1980_n ) capacitor c=0.0115788f //x=13.29 \
 //y=1.665 //x2=26.155 //y2=2.59
cc_854 ( N_noxref_4_c_930_n N_SN_c_1980_n ) capacitor c=0.0228083f //x=13.69 \
 //y=2.96 //x2=26.155 //y2=2.59
cc_855 ( N_noxref_4_c_904_n N_SN_c_1980_n ) capacitor c=0.024186f //x=15.54 \
 //y=2.08 //x2=26.155 //y2=2.59
cc_856 ( N_noxref_4_c_909_n N_SN_c_1980_n ) capacitor c=0.00712164f //x=15.24 \
 //y=1.915 //x2=26.155 //y2=2.59
cc_857 ( N_noxref_4_c_916_n N_SN_c_1991_n ) capacitor c=0.0144268f //x=11.945 \
 //y=5.155 //x2=11.84 //y2=2.08
cc_858 ( N_noxref_4_c_930_n N_SN_c_1991_n ) capacitor c=0.00265678f //x=13.69 \
 //y=2.96 //x2=11.84 //y2=2.08
cc_859 ( N_noxref_4_c_916_n N_SN_M32_noxref_g ) capacitor c=0.0165266f \
 //x=11.945 //y=5.155 //x2=11.81 //y2=6.02
cc_860 ( N_noxref_4_M32_noxref_d N_SN_M32_noxref_g ) capacitor c=0.0180032f \
 //x=11.885 //y=5.02 //x2=11.81 //y2=6.02
cc_861 ( N_noxref_4_c_922_n N_SN_M33_noxref_g ) capacitor c=0.01736f \
 //x=12.825 //y=5.155 //x2=12.25 //y2=6.02
cc_862 ( N_noxref_4_M32_noxref_d N_SN_M33_noxref_g ) capacitor c=0.0180032f \
 //x=11.885 //y=5.02 //x2=12.25 //y2=6.02
cc_863 ( N_noxref_4_c_1010_p N_SN_c_2039_n ) capacitor c=0.00426767f //x=12.03 \
 //y=5.155 //x2=12.175 //y2=4.79
cc_864 ( N_noxref_4_c_916_n N_SN_c_2024_n ) capacitor c=0.00322054f //x=11.945 \
 //y=5.155 //x2=11.84 //y2=4.7
cc_865 ( N_noxref_4_c_930_n N_noxref_10_c_2215_n ) capacitor c=0.0181982f \
 //x=13.69 //y=2.96 //x2=18.385 //y2=4.07
cc_866 ( N_noxref_4_c_904_n N_noxref_10_c_2215_n ) capacitor c=0.019517f \
 //x=15.54 //y=2.08 //x2=18.385 //y2=4.07
cc_867 ( N_noxref_4_c_930_n N_noxref_10_c_2278_n ) capacitor c=0.00179385f \
 //x=13.69 //y=2.96 //x2=13.065 //y2=4.07
cc_868 ( N_noxref_4_c_955_n N_noxref_10_c_2210_n ) capacitor c=0.00458487f \
 //x=13.805 //y=2.96 //x2=12.95 //y2=2.08
cc_869 ( N_noxref_4_c_930_n N_noxref_10_c_2210_n ) capacitor c=0.0790607f \
 //x=13.69 //y=2.96 //x2=12.95 //y2=2.08
cc_870 ( N_noxref_4_c_904_n N_noxref_10_c_2210_n ) capacitor c=8.48165e-19 \
 //x=15.54 //y=2.08 //x2=12.95 //y2=2.08
cc_871 ( N_noxref_4_c_1018_p N_noxref_10_c_2210_n ) capacitor c=0.0171303f \
 //x=12.91 //y=5.155 //x2=12.95 //y2=2.08
cc_872 ( N_noxref_4_M37_noxref_g N_noxref_10_c_2225_n ) capacitor c=0.0168349f \
 //x=16.18 //y=6.02 //x2=16.755 //y2=5.155
cc_873 ( N_noxref_4_c_926_n N_noxref_10_c_2229_n ) capacitor c=3.10026e-19 \
 //x=13.605 //y=5.155 //x2=16.045 //y2=5.155
cc_874 ( N_noxref_4_M36_noxref_g N_noxref_10_c_2229_n ) capacitor c=0.0213876f \
 //x=15.74 //y=6.02 //x2=16.045 //y2=5.155
cc_875 ( N_noxref_4_c_968_p N_noxref_10_c_2229_n ) capacitor c=0.00428486f \
 //x=16.105 //y=4.79 //x2=16.045 //y2=5.155
cc_876 ( N_noxref_4_c_922_n N_noxref_10_M34_noxref_g ) capacitor c=0.01736f \
 //x=12.825 //y=5.155 //x2=12.69 //y2=6.02
cc_877 ( N_noxref_4_M34_noxref_d N_noxref_10_M34_noxref_g ) capacitor \
 c=0.0180032f //x=12.765 //y=5.02 //x2=12.69 //y2=6.02
cc_878 ( N_noxref_4_c_926_n N_noxref_10_M35_noxref_g ) capacitor c=0.0194981f \
 //x=13.605 //y=5.155 //x2=13.13 //y2=6.02
cc_879 ( N_noxref_4_M34_noxref_d N_noxref_10_M35_noxref_g ) capacitor \
 c=0.0194246f //x=12.765 //y=5.02 //x2=13.13 //y2=6.02
cc_880 ( N_noxref_4_M8_noxref_d N_noxref_10_c_2291_n ) capacitor c=0.00217566f \
 //x=13.015 //y=0.915 //x2=12.94 //y2=0.915
cc_881 ( N_noxref_4_M8_noxref_d N_noxref_10_c_2292_n ) capacitor c=0.0034598f \
 //x=13.015 //y=0.915 //x2=12.94 //y2=1.26
cc_882 ( N_noxref_4_M8_noxref_d N_noxref_10_c_2293_n ) capacitor c=0.00544291f \
 //x=13.015 //y=0.915 //x2=12.94 //y2=1.57
cc_883 ( N_noxref_4_M8_noxref_d N_noxref_10_c_2294_n ) capacitor c=0.00241102f \
 //x=13.015 //y=0.915 //x2=13.315 //y2=0.76
cc_884 ( N_noxref_4_c_903_n N_noxref_10_c_2295_n ) capacitor c=0.00359704f \
 //x=13.605 //y=1.665 //x2=13.315 //y2=1.415
cc_885 ( N_noxref_4_M8_noxref_d N_noxref_10_c_2295_n ) capacitor c=0.0140297f \
 //x=13.015 //y=0.915 //x2=13.315 //y2=1.415
cc_886 ( N_noxref_4_M8_noxref_d N_noxref_10_c_2297_n ) capacitor c=0.00219619f \
 //x=13.015 //y=0.915 //x2=13.47 //y2=0.915
cc_887 ( N_noxref_4_c_903_n N_noxref_10_c_2298_n ) capacitor c=0.00457401f \
 //x=13.605 //y=1.665 //x2=13.47 //y2=1.26
cc_888 ( N_noxref_4_M8_noxref_d N_noxref_10_c_2298_n ) capacitor c=0.00603828f \
 //x=13.015 //y=0.915 //x2=13.47 //y2=1.26
cc_889 ( N_noxref_4_c_930_n N_noxref_10_c_2300_n ) capacitor c=0.00877984f \
 //x=13.69 //y=2.96 //x2=12.95 //y2=2.08
cc_890 ( N_noxref_4_c_930_n N_noxref_10_c_2301_n ) capacitor c=0.00283672f \
 //x=13.69 //y=2.96 //x2=12.95 //y2=1.915
cc_891 ( N_noxref_4_M8_noxref_d N_noxref_10_c_2301_n ) capacitor c=0.00661782f \
 //x=13.015 //y=0.915 //x2=12.95 //y2=1.915
cc_892 ( N_noxref_4_c_926_n N_noxref_10_c_2303_n ) capacitor c=0.00201851f \
 //x=13.605 //y=5.155 //x2=12.95 //y2=4.7
cc_893 ( N_noxref_4_c_930_n N_noxref_10_c_2303_n ) capacitor c=0.013844f \
 //x=13.69 //y=2.96 //x2=12.95 //y2=4.7
cc_894 ( N_noxref_4_c_1018_p N_noxref_10_c_2303_n ) capacitor c=0.00475601f \
 //x=12.91 //y=5.155 //x2=12.95 //y2=4.7
cc_895 ( N_noxref_4_M37_noxref_g N_noxref_10_M36_noxref_d ) capacitor \
 c=0.0180032f //x=16.18 //y=6.02 //x2=15.815 //y2=5.02
cc_896 ( N_noxref_4_M8_noxref_d N_noxref_17_M6_noxref_s ) capacitor \
 c=0.00309936f //x=13.015 //y=0.915 //x2=10.075 //y2=0.375
cc_897 ( N_noxref_4_c_903_n N_noxref_18_c_3027_n ) capacitor c=0.00461497f \
 //x=13.605 //y=1.665 //x2=13.605 //y2=0.54
cc_898 ( N_noxref_4_M8_noxref_d N_noxref_18_c_3027_n ) capacitor c=0.0116817f \
 //x=13.015 //y=0.915 //x2=13.605 //y2=0.54
cc_899 ( N_noxref_4_c_1000_p N_noxref_18_c_3038_n ) capacitor c=0.0200405f \
 //x=13.29 //y=1.665 //x2=12.72 //y2=0.995
cc_900 ( N_noxref_4_M8_noxref_d N_noxref_18_M7_noxref_d ) capacitor \
 c=5.27807e-19 //x=13.015 //y=0.915 //x2=11.48 //y2=0.91
cc_901 ( N_noxref_4_c_903_n N_noxref_18_M8_noxref_s ) capacitor c=0.0201579f \
 //x=13.605 //y=1.665 //x2=12.585 //y2=0.375
cc_902 ( N_noxref_4_M8_noxref_d N_noxref_18_M8_noxref_s ) capacitor \
 c=0.0426368f //x=13.015 //y=0.915 //x2=12.585 //y2=0.375
cc_903 ( N_noxref_4_c_903_n N_noxref_19_c_3091_n ) capacitor c=3.84569e-19 \
 //x=13.605 //y=1.665 //x2=15.02 //y2=1.505
cc_904 ( N_noxref_4_c_909_n N_noxref_19_c_3091_n ) capacitor c=0.0034165f \
 //x=15.24 //y=1.915 //x2=15.02 //y2=1.505
cc_905 ( N_noxref_4_c_904_n N_noxref_19_c_3075_n ) capacitor c=0.0117982f \
 //x=15.54 //y=2.08 //x2=15.905 //y2=1.59
cc_906 ( N_noxref_4_c_908_n N_noxref_19_c_3075_n ) capacitor c=0.00703864f \
 //x=15.24 //y=1.53 //x2=15.905 //y2=1.59
cc_907 ( N_noxref_4_c_909_n N_noxref_19_c_3075_n ) capacitor c=0.0215834f \
 //x=15.24 //y=1.915 //x2=15.905 //y2=1.59
cc_908 ( N_noxref_4_c_911_n N_noxref_19_c_3075_n ) capacitor c=0.00708583f \
 //x=15.615 //y=1.375 //x2=15.905 //y2=1.59
cc_909 ( N_noxref_4_c_914_n N_noxref_19_c_3075_n ) capacitor c=0.00698822f \
 //x=15.77 //y=1.22 //x2=15.905 //y2=1.59
cc_910 ( N_noxref_4_c_905_n N_noxref_19_M9_noxref_s ) capacitor c=0.0327271f \
 //x=15.24 //y=0.875 //x2=14.885 //y2=0.375
cc_911 ( N_noxref_4_c_908_n N_noxref_19_M9_noxref_s ) capacitor c=7.99997e-19 \
 //x=15.24 //y=1.53 //x2=14.885 //y2=0.375
cc_912 ( N_noxref_4_c_909_n N_noxref_19_M9_noxref_s ) capacitor c=0.00122123f \
 //x=15.24 //y=1.915 //x2=14.885 //y2=0.375
cc_913 ( N_noxref_4_c_912_n N_noxref_19_M9_noxref_s ) capacitor c=0.0121427f \
 //x=15.77 //y=0.875 //x2=14.885 //y2=0.375
cc_914 ( N_noxref_4_M8_noxref_d N_noxref_19_M9_noxref_s ) capacitor \
 c=2.55333e-19 //x=13.015 //y=0.915 //x2=14.885 //y2=0.375
cc_915 ( N_CLK_c_1062_n N_noxref_6_c_1253_n ) capacitor c=0.14131f //x=16.535 \
 //y=3.33 //x2=8.765 //y2=3.7
cc_916 ( N_CLK_c_1079_n N_noxref_6_c_1253_n ) capacitor c=0.029189f //x=7.145 \
 //y=3.33 //x2=8.765 //y2=3.7
cc_917 ( N_CLK_c_1063_n N_noxref_6_c_1253_n ) capacitor c=0.0231796f //x=7.03 \
 //y=2.08 //x2=8.765 //y2=3.7
cc_918 ( N_CLK_c_1062_n N_noxref_6_c_1255_n ) capacitor c=0.697076f //x=16.535 \
 //y=3.33 //x2=20.235 //y2=3.7
cc_919 ( N_CLK_c_1064_n N_noxref_6_c_1255_n ) capacitor c=0.0208745f //x=16.65 \
 //y=2.08 //x2=20.235 //y2=3.7
cc_920 ( N_CLK_c_1062_n N_noxref_6_c_1325_n ) capacitor c=0.0268461f \
 //x=16.535 //y=3.33 //x2=8.995 //y2=3.7
cc_921 ( N_CLK_c_1063_n N_noxref_6_c_1272_n ) capacitor c=0.0144268f //x=7.03 \
 //y=2.08 //x2=7.135 //y2=5.155
cc_922 ( N_CLK_M26_noxref_g N_noxref_6_c_1272_n ) capacitor c=0.0165266f //x=7 \
 //y=6.02 //x2=7.135 //y2=5.155
cc_923 ( N_CLK_c_1102_n N_noxref_6_c_1272_n ) capacitor c=0.00322054f //x=7.03 \
 //y=4.7 //x2=7.135 //y2=5.155
cc_924 ( N_CLK_M27_noxref_g N_noxref_6_c_1278_n ) capacitor c=0.01736f \
 //x=7.44 //y=6.02 //x2=8.015 //y2=5.155
cc_925 ( N_CLK_c_1062_n N_noxref_6_c_1286_n ) capacitor c=0.0205384f \
 //x=16.535 //y=3.33 //x2=8.88 //y2=3.7
cc_926 ( N_CLK_c_1063_n N_noxref_6_c_1286_n ) capacitor c=0.00286753f //x=7.03 \
 //y=2.08 //x2=8.88 //y2=3.7
cc_927 ( N_CLK_c_1143_p N_noxref_6_c_1375_n ) capacitor c=0.00426767f \
 //x=7.365 //y=4.79 //x2=7.22 //y2=5.155
cc_928 ( N_CLK_M26_noxref_g N_noxref_6_M26_noxref_d ) capacitor c=0.0180032f \
 //x=7 //y=6.02 //x2=7.075 //y2=5.02
cc_929 ( N_CLK_M27_noxref_g N_noxref_6_M26_noxref_d ) capacitor c=0.0180032f \
 //x=7.44 //y=6.02 //x2=7.075 //y2=5.02
cc_930 ( N_CLK_c_1062_n N_RN_c_1514_n ) capacitor c=0.00660904f //x=16.535 \
 //y=3.33 //x2=17.645 //y2=4.44
cc_931 ( N_CLK_c_1079_n N_RN_c_1514_n ) capacitor c=7.33995e-19 //x=7.145 \
 //y=3.33 //x2=17.645 //y2=4.44
cc_932 ( N_CLK_c_1063_n N_RN_c_1514_n ) capacitor c=0.0233868f //x=7.03 \
 //y=2.08 //x2=17.645 //y2=4.44
cc_933 ( N_CLK_c_1064_n N_RN_c_1514_n ) capacitor c=0.0210462f //x=16.65 \
 //y=2.08 //x2=17.645 //y2=4.44
cc_934 ( N_CLK_c_1143_p N_RN_c_1514_n ) capacitor c=0.0085986f //x=7.365 \
 //y=4.79 //x2=17.645 //y2=4.44
cc_935 ( N_CLK_c_1151_p N_RN_c_1514_n ) capacitor c=0.0085986f //x=16.985 \
 //y=4.79 //x2=17.645 //y2=4.44
cc_936 ( N_CLK_c_1102_n N_RN_c_1514_n ) capacitor c=0.00293313f //x=7.03 \
 //y=4.7 //x2=17.645 //y2=4.44
cc_937 ( N_CLK_c_1128_n N_RN_c_1514_n ) capacitor c=0.00293313f //x=16.65 \
 //y=4.7 //x2=17.645 //y2=4.44
cc_938 ( N_CLK_c_1064_n N_RN_c_1542_n ) capacitor c=0.00153281f //x=16.65 \
 //y=2.08 //x2=17.875 //y2=4.44
cc_939 ( N_CLK_c_1062_n N_RN_c_1517_n ) capacitor c=0.00526349f //x=16.535 \
 //y=3.33 //x2=17.76 //y2=2.08
cc_940 ( N_CLK_c_1064_n N_RN_c_1517_n ) capacitor c=0.0464118f //x=16.65 \
 //y=2.08 //x2=17.76 //y2=2.08
cc_941 ( N_CLK_c_1126_n N_RN_c_1517_n ) capacitor c=0.0023343f //x=16.74 \
 //y=1.915 //x2=17.76 //y2=2.08
cc_942 ( N_CLK_c_1128_n N_RN_c_1517_n ) capacitor c=0.00141297f //x=16.65 \
 //y=4.7 //x2=17.76 //y2=2.08
cc_943 ( N_CLK_M38_noxref_g N_RN_M40_noxref_g ) capacitor c=0.0101598f \
 //x=16.62 //y=6.02 //x2=17.5 //y2=6.02
cc_944 ( N_CLK_M39_noxref_g N_RN_M40_noxref_g ) capacitor c=0.0602553f \
 //x=17.06 //y=6.02 //x2=17.5 //y2=6.02
cc_945 ( N_CLK_M39_noxref_g N_RN_M41_noxref_g ) capacitor c=0.0101598f \
 //x=17.06 //y=6.02 //x2=17.94 //y2=6.02
cc_946 ( N_CLK_c_1123_n N_RN_c_1603_n ) capacitor c=0.00456962f //x=16.74 \
 //y=0.91 //x2=17.75 //y2=0.915
cc_947 ( N_CLK_c_1124_n N_RN_c_1604_n ) capacitor c=0.00438372f //x=16.74 \
 //y=1.22 //x2=17.75 //y2=1.26
cc_948 ( N_CLK_c_1125_n N_RN_c_1605_n ) capacitor c=0.00438372f //x=16.74 \
 //y=1.45 //x2=17.75 //y2=1.57
cc_949 ( N_CLK_c_1064_n N_RN_c_1606_n ) capacitor c=0.00228632f //x=16.65 \
 //y=2.08 //x2=17.76 //y2=2.08
cc_950 ( N_CLK_c_1126_n N_RN_c_1606_n ) capacitor c=0.00933826f //x=16.74 \
 //y=1.915 //x2=17.76 //y2=2.08
cc_951 ( N_CLK_c_1126_n N_RN_c_1608_n ) capacitor c=0.00438372f //x=16.74 \
 //y=1.915 //x2=17.76 //y2=1.915
cc_952 ( N_CLK_c_1064_n N_RN_c_1609_n ) capacitor c=0.00219458f //x=16.65 \
 //y=2.08 //x2=17.76 //y2=4.7
cc_953 ( N_CLK_c_1151_p N_RN_c_1609_n ) capacitor c=0.0611812f //x=16.985 \
 //y=4.79 //x2=17.76 //y2=4.7
cc_954 ( N_CLK_c_1128_n N_RN_c_1609_n ) capacitor c=0.00487508f //x=16.65 \
 //y=4.7 //x2=17.76 //y2=4.7
cc_955 ( N_CLK_c_1062_n N_SN_c_1980_n ) capacitor c=0.128638f //x=16.535 \
 //y=3.33 //x2=26.155 //y2=2.59
cc_956 ( N_CLK_c_1064_n N_SN_c_1980_n ) capacitor c=0.0251844f //x=16.65 \
 //y=2.08 //x2=26.155 //y2=2.59
cc_957 ( N_CLK_c_1126_n N_SN_c_1980_n ) capacitor c=0.00263139f //x=16.74 \
 //y=1.915 //x2=26.155 //y2=2.59
cc_958 ( N_CLK_c_1062_n N_SN_c_1990_n ) capacitor c=0.0133087f //x=16.535 \
 //y=3.33 //x2=11.955 //y2=2.59
cc_959 ( N_CLK_c_1062_n N_SN_c_1991_n ) capacitor c=0.0217085f //x=16.535 \
 //y=3.33 //x2=11.84 //y2=2.08
cc_960 ( N_CLK_c_1062_n N_noxref_10_c_2214_n ) capacitor c=0.0347141f \
 //x=16.535 //y=3.33 //x2=12.835 //y2=4.07
cc_961 ( N_CLK_c_1062_n N_noxref_10_c_2308_n ) capacitor c=7.00757e-19 \
 //x=16.535 //y=3.33 //x2=8.25 //y2=4.07
cc_962 ( N_CLK_c_1063_n N_noxref_10_c_2308_n ) capacitor c=0.00528706f \
 //x=7.03 //y=2.08 //x2=8.25 //y2=4.07
cc_963 ( N_CLK_c_1062_n N_noxref_10_c_2215_n ) capacitor c=0.0257572f \
 //x=16.535 //y=3.33 //x2=18.385 //y2=4.07
cc_964 ( N_CLK_c_1064_n N_noxref_10_c_2215_n ) capacitor c=0.0190126f \
 //x=16.65 //y=2.08 //x2=18.385 //y2=4.07
cc_965 ( N_CLK_c_1062_n N_noxref_10_c_2278_n ) capacitor c=4.7279e-19 \
 //x=16.535 //y=3.33 //x2=13.065 //y2=4.07
cc_966 ( N_CLK_c_1062_n N_noxref_10_c_2209_n ) capacitor c=0.0179796f \
 //x=16.535 //y=3.33 //x2=8.14 //y2=2.08
cc_967 ( N_CLK_c_1079_n N_noxref_10_c_2209_n ) capacitor c=0.00128547f \
 //x=7.145 //y=3.33 //x2=8.14 //y2=2.08
cc_968 ( N_CLK_c_1063_n N_noxref_10_c_2209_n ) capacitor c=0.0322045f //x=7.03 \
 //y=2.08 //x2=8.14 //y2=2.08
cc_969 ( N_CLK_c_1099_n N_noxref_10_c_2209_n ) capacitor c=0.0023343f //x=7.12 \
 //y=1.915 //x2=8.14 //y2=2.08
cc_970 ( N_CLK_c_1063_n N_noxref_10_c_2317_n ) capacitor c=0.00867715f \
 //x=7.03 //y=2.08 //x2=8.14 //y2=4.7
cc_971 ( N_CLK_c_1102_n N_noxref_10_c_2317_n ) capacitor c=0.00142741f \
 //x=7.03 //y=4.7 //x2=8.14 //y2=4.7
cc_972 ( N_CLK_c_1062_n N_noxref_10_c_2210_n ) capacitor c=0.0203592f \
 //x=16.535 //y=3.33 //x2=12.95 //y2=2.08
cc_973 ( N_CLK_c_1064_n N_noxref_10_c_2225_n ) capacitor c=0.0144268f \
 //x=16.65 //y=2.08 //x2=16.755 //y2=5.155
cc_974 ( N_CLK_M38_noxref_g N_noxref_10_c_2225_n ) capacitor c=0.0165266f \
 //x=16.62 //y=6.02 //x2=16.755 //y2=5.155
cc_975 ( N_CLK_c_1128_n N_noxref_10_c_2225_n ) capacitor c=0.00322054f \
 //x=16.65 //y=4.7 //x2=16.755 //y2=5.155
cc_976 ( N_CLK_M39_noxref_g N_noxref_10_c_2231_n ) capacitor c=0.01736f \
 //x=17.06 //y=6.02 //x2=17.635 //y2=5.155
cc_977 ( N_CLK_c_1064_n N_noxref_10_c_2239_n ) capacitor c=0.00315138f \
 //x=16.65 //y=2.08 //x2=18.5 //y2=4.07
cc_978 ( N_CLK_c_1063_n N_noxref_10_c_2241_n ) capacitor c=0.00609925f \
 //x=7.03 //y=2.08 //x2=8.135 //y2=4.07
cc_979 ( N_CLK_c_1151_p N_noxref_10_c_2326_n ) capacitor c=0.00426767f \
 //x=16.985 //y=4.79 //x2=16.84 //y2=5.155
cc_980 ( N_CLK_M26_noxref_g N_noxref_10_M28_noxref_g ) capacitor c=0.0101598f \
 //x=7 //y=6.02 //x2=7.88 //y2=6.02
cc_981 ( N_CLK_M27_noxref_g N_noxref_10_M28_noxref_g ) capacitor c=0.0602553f \
 //x=7.44 //y=6.02 //x2=7.88 //y2=6.02
cc_982 ( N_CLK_M27_noxref_g N_noxref_10_M29_noxref_g ) capacitor c=0.0101598f \
 //x=7.44 //y=6.02 //x2=8.32 //y2=6.02
cc_983 ( N_CLK_c_1096_n N_noxref_10_c_2330_n ) capacitor c=0.00456962f \
 //x=7.12 //y=0.91 //x2=8.13 //y2=0.915
cc_984 ( N_CLK_c_1097_n N_noxref_10_c_2331_n ) capacitor c=0.00438372f \
 //x=7.12 //y=1.22 //x2=8.13 //y2=1.26
cc_985 ( N_CLK_c_1098_n N_noxref_10_c_2332_n ) capacitor c=0.00438372f \
 //x=7.12 //y=1.45 //x2=8.13 //y2=1.57
cc_986 ( N_CLK_c_1063_n N_noxref_10_c_2275_n ) capacitor c=0.00228632f \
 //x=7.03 //y=2.08 //x2=8.14 //y2=2.08
cc_987 ( N_CLK_c_1099_n N_noxref_10_c_2275_n ) capacitor c=0.00933826f \
 //x=7.12 //y=1.915 //x2=8.14 //y2=2.08
cc_988 ( N_CLK_c_1099_n N_noxref_10_c_2335_n ) capacitor c=0.00438372f \
 //x=7.12 //y=1.915 //x2=8.14 //y2=1.915
cc_989 ( N_CLK_c_1063_n N_noxref_10_c_2336_n ) capacitor c=0.00219458f \
 //x=7.03 //y=2.08 //x2=8.14 //y2=4.7
cc_990 ( N_CLK_c_1143_p N_noxref_10_c_2336_n ) capacitor c=0.0611812f \
 //x=7.365 //y=4.79 //x2=8.14 //y2=4.7
cc_991 ( N_CLK_c_1102_n N_noxref_10_c_2336_n ) capacitor c=0.00487508f \
 //x=7.03 //y=4.7 //x2=8.14 //y2=4.7
cc_992 ( N_CLK_M38_noxref_g N_noxref_10_M38_noxref_d ) capacitor c=0.0180032f \
 //x=16.62 //y=6.02 //x2=16.695 //y2=5.02
cc_993 ( N_CLK_M39_noxref_g N_noxref_10_M38_noxref_d ) capacitor c=0.0180032f \
 //x=17.06 //y=6.02 //x2=16.695 //y2=5.02
cc_994 ( N_CLK_c_1091_n N_noxref_15_c_2868_n ) capacitor c=0.0167228f \
 //x=6.595 //y=0.91 //x2=7.255 //y2=0.54
cc_995 ( N_CLK_c_1096_n N_noxref_15_c_2868_n ) capacitor c=0.00534519f \
 //x=7.12 //y=0.91 //x2=7.255 //y2=0.54
cc_996 ( N_CLK_c_1063_n N_noxref_15_c_2888_n ) capacitor c=0.0124901f //x=7.03 \
 //y=2.08 //x2=7.255 //y2=1.59
cc_997 ( N_CLK_c_1094_n N_noxref_15_c_2888_n ) capacitor c=0.0153476f \
 //x=6.595 //y=1.22 //x2=7.255 //y2=1.59
cc_998 ( N_CLK_c_1099_n N_noxref_15_c_2888_n ) capacitor c=0.0223834f //x=7.12 \
 //y=1.915 //x2=7.255 //y2=1.59
cc_999 ( N_CLK_c_1091_n N_noxref_15_M3_noxref_s ) capacitor c=0.00798959f \
 //x=6.595 //y=0.91 //x2=5.265 //y2=0.375
cc_1000 ( N_CLK_c_1098_n N_noxref_15_M3_noxref_s ) capacitor c=0.00212176f \
 //x=7.12 //y=1.45 //x2=5.265 //y2=0.375
cc_1001 ( N_CLK_c_1099_n N_noxref_15_M3_noxref_s ) capacitor c=0.00298115f \
 //x=7.12 //y=1.915 //x2=5.265 //y2=0.375
cc_1002 ( N_CLK_c_1218_p N_noxref_16_c_2913_n ) capacitor c=2.14837e-19 \
 //x=6.965 //y=0.755 //x2=7.825 //y2=0.995
cc_1003 ( N_CLK_c_1096_n N_noxref_16_c_2913_n ) capacitor c=0.00123426f \
 //x=7.12 //y=0.91 //x2=7.825 //y2=0.995
cc_1004 ( N_CLK_c_1097_n N_noxref_16_c_2913_n ) capacitor c=0.0129288f \
 //x=7.12 //y=1.22 //x2=7.825 //y2=0.995
cc_1005 ( N_CLK_c_1098_n N_noxref_16_c_2913_n ) capacitor c=0.00142359f \
 //x=7.12 //y=1.45 //x2=7.825 //y2=0.995
cc_1006 ( N_CLK_c_1091_n N_noxref_16_M4_noxref_d ) capacitor c=0.00223875f \
 //x=6.595 //y=0.91 //x2=6.67 //y2=0.91
cc_1007 ( N_CLK_c_1094_n N_noxref_16_M4_noxref_d ) capacitor c=0.00262485f \
 //x=6.595 //y=1.22 //x2=6.67 //y2=0.91
cc_1008 ( N_CLK_c_1218_p N_noxref_16_M4_noxref_d ) capacitor c=0.00220746f \
 //x=6.965 //y=0.755 //x2=6.67 //y2=0.91
cc_1009 ( N_CLK_c_1225_p N_noxref_16_M4_noxref_d ) capacitor c=0.00194798f \
 //x=6.965 //y=1.375 //x2=6.67 //y2=0.91
cc_1010 ( N_CLK_c_1096_n N_noxref_16_M4_noxref_d ) capacitor c=0.00198465f \
 //x=7.12 //y=0.91 //x2=6.67 //y2=0.91
cc_1011 ( N_CLK_c_1097_n N_noxref_16_M4_noxref_d ) capacitor c=0.00128384f \
 //x=7.12 //y=1.22 //x2=6.67 //y2=0.91
cc_1012 ( N_CLK_c_1096_n N_noxref_16_M5_noxref_s ) capacitor c=7.21316e-19 \
 //x=7.12 //y=0.91 //x2=7.775 //y2=0.375
cc_1013 ( N_CLK_c_1097_n N_noxref_16_M5_noxref_s ) capacitor c=0.00348171f \
 //x=7.12 //y=1.22 //x2=7.775 //y2=0.375
cc_1014 ( N_CLK_c_1062_n N_noxref_17_c_2967_n ) capacitor c=0.00263604f \
 //x=16.535 //y=3.33 //x2=11.095 //y2=1.59
cc_1015 ( N_CLK_c_1062_n N_noxref_17_c_2997_n ) capacitor c=0.00504206f \
 //x=16.535 //y=3.33 //x2=12.065 //y2=1.59
cc_1016 ( N_CLK_c_1062_n N_noxref_17_M6_noxref_s ) capacitor c=0.00243521f \
 //x=16.535 //y=3.33 //x2=10.075 //y2=0.375
cc_1017 ( N_CLK_c_1118_n N_noxref_19_c_3082_n ) capacitor c=0.0167228f \
 //x=16.215 //y=0.91 //x2=16.875 //y2=0.54
cc_1018 ( N_CLK_c_1123_n N_noxref_19_c_3082_n ) capacitor c=0.00534519f \
 //x=16.74 //y=0.91 //x2=16.875 //y2=0.54
cc_1019 ( N_CLK_c_1064_n N_noxref_19_c_3105_n ) capacitor c=0.012061f \
 //x=16.65 //y=2.08 //x2=16.875 //y2=1.59
cc_1020 ( N_CLK_c_1121_n N_noxref_19_c_3105_n ) capacitor c=0.0153476f \
 //x=16.215 //y=1.22 //x2=16.875 //y2=1.59
cc_1021 ( N_CLK_c_1126_n N_noxref_19_c_3105_n ) capacitor c=0.0219329f \
 //x=16.74 //y=1.915 //x2=16.875 //y2=1.59
cc_1022 ( N_CLK_c_1118_n N_noxref_19_M9_noxref_s ) capacitor c=0.00798959f \
 //x=16.215 //y=0.91 //x2=14.885 //y2=0.375
cc_1023 ( N_CLK_c_1125_n N_noxref_19_M9_noxref_s ) capacitor c=0.00212176f \
 //x=16.74 //y=1.45 //x2=14.885 //y2=0.375
cc_1024 ( N_CLK_c_1126_n N_noxref_19_M9_noxref_s ) capacitor c=0.00298115f \
 //x=16.74 //y=1.915 //x2=14.885 //y2=0.375
cc_1025 ( N_CLK_c_1241_p N_noxref_20_c_3125_n ) capacitor c=2.14837e-19 \
 //x=16.585 //y=0.755 //x2=17.445 //y2=0.995
cc_1026 ( N_CLK_c_1123_n N_noxref_20_c_3125_n ) capacitor c=0.00123426f \
 //x=16.74 //y=0.91 //x2=17.445 //y2=0.995
cc_1027 ( N_CLK_c_1124_n N_noxref_20_c_3125_n ) capacitor c=0.0129288f \
 //x=16.74 //y=1.22 //x2=17.445 //y2=0.995
cc_1028 ( N_CLK_c_1125_n N_noxref_20_c_3125_n ) capacitor c=0.00142359f \
 //x=16.74 //y=1.45 //x2=17.445 //y2=0.995
cc_1029 ( N_CLK_c_1118_n N_noxref_20_M10_noxref_d ) capacitor c=0.00223875f \
 //x=16.215 //y=0.91 //x2=16.29 //y2=0.91
cc_1030 ( N_CLK_c_1121_n N_noxref_20_M10_noxref_d ) capacitor c=0.00262485f \
 //x=16.215 //y=1.22 //x2=16.29 //y2=0.91
cc_1031 ( N_CLK_c_1241_p N_noxref_20_M10_noxref_d ) capacitor c=0.00220746f \
 //x=16.585 //y=0.755 //x2=16.29 //y2=0.91
cc_1032 ( N_CLK_c_1248_p N_noxref_20_M10_noxref_d ) capacitor c=0.00194798f \
 //x=16.585 //y=1.375 //x2=16.29 //y2=0.91
cc_1033 ( N_CLK_c_1123_n N_noxref_20_M10_noxref_d ) capacitor c=0.00198465f \
 //x=16.74 //y=0.91 //x2=16.29 //y2=0.91
cc_1034 ( N_CLK_c_1124_n N_noxref_20_M10_noxref_d ) capacitor c=0.00128384f \
 //x=16.74 //y=1.22 //x2=16.29 //y2=0.91
cc_1035 ( N_CLK_c_1123_n N_noxref_20_M11_noxref_s ) capacitor c=7.21316e-19 \
 //x=16.74 //y=0.91 //x2=17.395 //y2=0.375
cc_1036 ( N_CLK_c_1124_n N_noxref_20_M11_noxref_s ) capacitor c=0.00348171f \
 //x=16.74 //y=1.22 //x2=17.395 //y2=0.375
cc_1037 ( N_noxref_6_c_1253_n N_RN_c_1514_n ) capacitor c=0.199363f //x=8.765 \
 //y=3.7 //x2=17.645 //y2=4.44
cc_1038 ( N_noxref_6_c_1254_n N_RN_c_1514_n ) capacitor c=0.0134983f //x=3.445 \
 //y=3.7 //x2=17.645 //y2=4.44
cc_1039 ( N_noxref_6_c_1255_n N_RN_c_1514_n ) capacitor c=0.0638008f \
 //x=20.235 //y=3.7 //x2=17.645 //y2=4.44
cc_1040 ( N_noxref_6_c_1325_n N_RN_c_1514_n ) capacitor c=4.78746e-19 \
 //x=8.995 //y=3.7 //x2=17.645 //y2=4.44
cc_1041 ( N_noxref_6_c_1256_n N_RN_c_1514_n ) capacitor c=0.0226638f //x=3.33 \
 //y=2.08 //x2=17.645 //y2=4.44
cc_1042 ( N_noxref_6_c_1272_n N_RN_c_1514_n ) capacitor c=0.032089f //x=7.135 \
 //y=5.155 //x2=17.645 //y2=4.44
cc_1043 ( N_noxref_6_c_1276_n N_RN_c_1514_n ) capacitor c=0.0230136f //x=6.425 \
 //y=5.155 //x2=17.645 //y2=4.44
cc_1044 ( N_noxref_6_c_1282_n N_RN_c_1514_n ) capacitor c=0.0183122f //x=8.795 \
 //y=5.155 //x2=17.645 //y2=4.44
cc_1045 ( N_noxref_6_c_1286_n N_RN_c_1514_n ) capacitor c=0.0210274f //x=8.88 \
 //y=3.7 //x2=17.645 //y2=4.44
cc_1046 ( N_noxref_6_c_1354_n N_RN_c_1514_n ) capacitor c=0.00988777f //x=3.33 \
 //y=4.7 //x2=17.645 //y2=4.44
cc_1047 ( N_noxref_6_c_1256_n N_RN_c_1515_n ) capacitor c=0.00153281f //x=3.33 \
 //y=2.08 //x2=2.335 //y2=4.44
cc_1048 ( N_noxref_6_c_1255_n N_RN_c_1536_n ) capacitor c=0.0157795f \
 //x=20.235 //y=3.7 //x2=21.345 //y2=4.44
cc_1049 ( N_noxref_6_c_1258_n N_RN_c_1536_n ) capacitor c=0.0218124f //x=20.35 \
 //y=2.08 //x2=21.345 //y2=4.44
cc_1050 ( N_noxref_6_c_1298_n N_RN_c_1536_n ) capacitor c=0.0168397f \
 //x=20.625 //y=4.79 //x2=21.345 //y2=4.44
cc_1051 ( N_noxref_6_c_1255_n N_RN_c_1542_n ) capacitor c=4.66937e-19 \
 //x=20.235 //y=3.7 //x2=17.875 //y2=4.44
cc_1052 ( N_noxref_6_c_1254_n N_RN_c_1516_n ) capacitor c=0.00526349f \
 //x=3.445 //y=3.7 //x2=2.22 //y2=2.08
cc_1053 ( N_noxref_6_c_1256_n N_RN_c_1516_n ) capacitor c=0.0535967f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_1054 ( N_noxref_6_c_1351_n N_RN_c_1516_n ) capacitor c=0.00228632f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_1055 ( N_noxref_6_c_1354_n N_RN_c_1516_n ) capacitor c=0.00218014f //x=3.33 \
 //y=4.7 //x2=2.22 //y2=2.08
cc_1056 ( N_noxref_6_c_1255_n N_RN_c_1517_n ) capacitor c=0.0218601f \
 //x=20.235 //y=3.7 //x2=17.76 //y2=2.08
cc_1057 ( N_noxref_6_c_1258_n N_RN_c_1517_n ) capacitor c=8.87185e-19 \
 //x=20.35 //y=2.08 //x2=17.76 //y2=2.08
cc_1058 ( N_noxref_6_c_1255_n N_RN_c_1518_n ) capacitor c=0.0027353f \
 //x=20.235 //y=3.7 //x2=21.46 //y2=2.08
cc_1059 ( N_noxref_6_c_1258_n N_RN_c_1518_n ) capacitor c=0.049364f //x=20.35 \
 //y=2.08 //x2=21.46 //y2=2.08
cc_1060 ( N_noxref_6_c_1263_n N_RN_c_1518_n ) capacitor c=0.00238338f \
 //x=20.05 //y=1.915 //x2=21.46 //y2=2.08
cc_1061 ( N_noxref_6_c_1402_p N_RN_c_1518_n ) capacitor c=0.00147352f \
 //x=20.915 //y=4.79 //x2=21.46 //y2=2.08
cc_1062 ( N_noxref_6_c_1298_n N_RN_c_1518_n ) capacitor c=0.00141297f \
 //x=20.625 //y=4.79 //x2=21.46 //y2=2.08
cc_1063 ( N_noxref_6_M22_noxref_g N_RN_M20_noxref_g ) capacitor c=0.0101598f \
 //x=3.07 //y=6.02 //x2=2.19 //y2=6.02
cc_1064 ( N_noxref_6_M22_noxref_g N_RN_M21_noxref_g ) capacitor c=0.0602553f \
 //x=3.07 //y=6.02 //x2=2.63 //y2=6.02
cc_1065 ( N_noxref_6_M23_noxref_g N_RN_M21_noxref_g ) capacitor c=0.0101598f \
 //x=3.51 //y=6.02 //x2=2.63 //y2=6.02
cc_1066 ( N_noxref_6_M42_noxref_g N_RN_M44_noxref_g ) capacitor c=0.0105869f \
 //x=20.55 //y=6.02 //x2=21.43 //y2=6.02
cc_1067 ( N_noxref_6_M43_noxref_g N_RN_M44_noxref_g ) capacitor c=0.10632f \
 //x=20.99 //y=6.02 //x2=21.43 //y2=6.02
cc_1068 ( N_noxref_6_M43_noxref_g N_RN_M45_noxref_g ) capacitor c=0.0101598f \
 //x=20.99 //y=6.02 //x2=21.87 //y2=6.02
cc_1069 ( N_noxref_6_c_1342_n N_RN_c_1644_n ) capacitor c=0.00456962f //x=3.32 \
 //y=0.915 //x2=2.31 //y2=0.91
cc_1070 ( N_noxref_6_c_1343_n N_RN_c_1645_n ) capacitor c=0.00438372f //x=3.32 \
 //y=1.26 //x2=2.31 //y2=1.22
cc_1071 ( N_noxref_6_c_1344_n N_RN_c_1646_n ) capacitor c=0.00438372f //x=3.32 \
 //y=1.57 //x2=2.31 //y2=1.45
cc_1072 ( N_noxref_6_c_1256_n N_RN_c_1647_n ) capacitor c=0.0023343f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_1073 ( N_noxref_6_c_1351_n N_RN_c_1647_n ) capacitor c=0.00933826f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_1074 ( N_noxref_6_c_1352_n N_RN_c_1647_n ) capacitor c=0.00438372f //x=3.33 \
 //y=1.915 //x2=2.31 //y2=1.915
cc_1075 ( N_noxref_6_c_1354_n N_RN_c_1578_n ) capacitor c=0.0611812f //x=3.33 \
 //y=4.7 //x2=2.555 //y2=4.79
cc_1076 ( N_noxref_6_c_1259_n N_RN_c_1651_n ) capacitor c=5.72482e-19 \
 //x=20.05 //y=0.875 //x2=21.025 //y2=0.91
cc_1077 ( N_noxref_6_c_1261_n N_RN_c_1651_n ) capacitor c=0.00149976f \
 //x=20.05 //y=1.22 //x2=21.025 //y2=0.91
cc_1078 ( N_noxref_6_c_1266_n N_RN_c_1651_n ) capacitor c=0.0160123f //x=20.58 \
 //y=0.875 //x2=21.025 //y2=0.91
cc_1079 ( N_noxref_6_c_1262_n N_RN_c_1654_n ) capacitor c=0.00111227f \
 //x=20.05 //y=1.53 //x2=21.025 //y2=1.22
cc_1080 ( N_noxref_6_c_1268_n N_RN_c_1654_n ) capacitor c=0.0124075f //x=20.58 \
 //y=1.22 //x2=21.025 //y2=1.22
cc_1081 ( N_noxref_6_c_1266_n N_RN_c_1656_n ) capacitor c=0.00103227f \
 //x=20.58 //y=0.875 //x2=21.55 //y2=0.91
cc_1082 ( N_noxref_6_c_1268_n N_RN_c_1657_n ) capacitor c=0.0010154f //x=20.58 \
 //y=1.22 //x2=21.55 //y2=1.22
cc_1083 ( N_noxref_6_c_1268_n N_RN_c_1658_n ) capacitor c=9.23422e-19 \
 //x=20.58 //y=1.22 //x2=21.55 //y2=1.45
cc_1084 ( N_noxref_6_c_1258_n N_RN_c_1659_n ) capacitor c=0.00231304f \
 //x=20.35 //y=2.08 //x2=21.55 //y2=1.915
cc_1085 ( N_noxref_6_c_1263_n N_RN_c_1659_n ) capacitor c=0.00964411f \
 //x=20.05 //y=1.915 //x2=21.55 //y2=1.915
cc_1086 ( N_noxref_6_c_1256_n N_RN_c_1579_n ) capacitor c=0.00142741f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=4.7
cc_1087 ( N_noxref_6_c_1354_n N_RN_c_1579_n ) capacitor c=0.00487508f //x=3.33 \
 //y=4.7 //x2=2.22 //y2=4.7
cc_1088 ( N_noxref_6_c_1258_n N_RN_c_1663_n ) capacitor c=0.00183762f \
 //x=20.35 //y=2.08 //x2=21.46 //y2=4.7
cc_1089 ( N_noxref_6_c_1402_p N_RN_c_1663_n ) capacitor c=0.0168581f \
 //x=20.915 //y=4.79 //x2=21.46 //y2=4.7
cc_1090 ( N_noxref_6_c_1298_n N_RN_c_1663_n ) capacitor c=0.00484466f \
 //x=20.625 //y=4.79 //x2=21.46 //y2=4.7
cc_1091 ( N_noxref_6_M43_noxref_g N_QN_c_1838_n ) capacitor c=0.0168349f \
 //x=20.99 //y=6.02 //x2=21.565 //y2=5.155
cc_1092 ( N_noxref_6_M42_noxref_g N_QN_c_1842_n ) capacitor c=0.0213876f \
 //x=20.55 //y=6.02 //x2=20.855 //y2=5.155
cc_1093 ( N_noxref_6_c_1402_p N_QN_c_1842_n ) capacitor c=0.00428486f \
 //x=20.915 //y=4.79 //x2=20.855 //y2=5.155
cc_1094 ( N_noxref_6_M43_noxref_g N_QN_M42_noxref_d ) capacitor c=0.0180032f \
 //x=20.99 //y=6.02 //x2=20.625 //y2=5.02
cc_1095 ( N_noxref_6_c_1255_n N_SN_c_1980_n ) capacitor c=0.122715f //x=20.235 \
 //y=3.7 //x2=26.155 //y2=2.59
cc_1096 ( N_noxref_6_c_1258_n N_SN_c_1980_n ) capacitor c=0.0263038f //x=20.35 \
 //y=2.08 //x2=26.155 //y2=2.59
cc_1097 ( N_noxref_6_c_1263_n N_SN_c_1980_n ) capacitor c=0.00537379f \
 //x=20.05 //y=1.915 //x2=26.155 //y2=2.59
cc_1098 ( N_noxref_6_c_1255_n N_SN_c_1990_n ) capacitor c=7.19251e-19 \
 //x=20.235 //y=3.7 //x2=11.955 //y2=2.59
cc_1099 ( N_noxref_6_c_1255_n N_SN_c_1991_n ) capacitor c=0.0190398f \
 //x=20.235 //y=3.7 //x2=11.84 //y2=2.08
cc_1100 ( N_noxref_6_c_1286_n N_SN_c_1991_n ) capacitor c=5.91559e-19 //x=8.88 \
 //y=3.7 //x2=11.84 //y2=2.08
cc_1101 ( N_noxref_6_c_1253_n N_noxref_10_c_2214_n ) capacitor c=0.0450244f \
 //x=8.765 //y=3.7 //x2=12.835 //y2=4.07
cc_1102 ( N_noxref_6_c_1255_n N_noxref_10_c_2214_n ) capacitor c=0.339801f \
 //x=20.235 //y=3.7 //x2=12.835 //y2=4.07
cc_1103 ( N_noxref_6_c_1325_n N_noxref_10_c_2214_n ) capacitor c=0.026809f \
 //x=8.995 //y=3.7 //x2=12.835 //y2=4.07
cc_1104 ( N_noxref_6_c_1286_n N_noxref_10_c_2214_n ) capacitor c=0.0200135f \
 //x=8.88 //y=3.7 //x2=12.835 //y2=4.07
cc_1105 ( N_noxref_6_c_1253_n N_noxref_10_c_2308_n ) capacitor c=0.0295035f \
 //x=8.765 //y=3.7 //x2=8.25 //y2=4.07
cc_1106 ( N_noxref_6_c_1286_n N_noxref_10_c_2308_n ) capacitor c=0.00178442f \
 //x=8.88 //y=3.7 //x2=8.25 //y2=4.07
cc_1107 ( N_noxref_6_c_1255_n N_noxref_10_c_2215_n ) capacitor c=0.468089f \
 //x=20.235 //y=3.7 //x2=18.385 //y2=4.07
cc_1108 ( N_noxref_6_c_1255_n N_noxref_10_c_2278_n ) capacitor c=0.0268959f \
 //x=20.235 //y=3.7 //x2=13.065 //y2=4.07
cc_1109 ( N_noxref_6_c_1255_n N_noxref_10_c_2216_n ) capacitor c=0.176507f \
 //x=20.235 //y=3.7 //x2=27.265 //y2=4.07
cc_1110 ( N_noxref_6_c_1258_n N_noxref_10_c_2216_n ) capacitor c=0.0213324f \
 //x=20.35 //y=2.08 //x2=27.265 //y2=4.07
cc_1111 ( N_noxref_6_c_1255_n N_noxref_10_c_2223_n ) capacitor c=0.0268461f \
 //x=20.235 //y=3.7 //x2=18.615 //y2=4.07
cc_1112 ( N_noxref_6_c_1258_n N_noxref_10_c_2223_n ) capacitor c=3.50683e-19 \
 //x=20.35 //y=2.08 //x2=18.615 //y2=4.07
cc_1113 ( N_noxref_6_c_1253_n N_noxref_10_c_2209_n ) capacitor c=0.0177645f \
 //x=8.765 //y=3.7 //x2=8.14 //y2=2.08
cc_1114 ( N_noxref_6_c_1325_n N_noxref_10_c_2209_n ) capacitor c=0.00179385f \
 //x=8.995 //y=3.7 //x2=8.14 //y2=2.08
cc_1115 ( N_noxref_6_c_1286_n N_noxref_10_c_2209_n ) capacitor c=0.0794709f \
 //x=8.88 //y=3.7 //x2=8.14 //y2=2.08
cc_1116 ( N_noxref_6_c_1457_p N_noxref_10_c_2317_n ) capacitor c=0.0166016f \
 //x=8.1 //y=5.155 //x2=8.14 //y2=4.7
cc_1117 ( N_noxref_6_c_1255_n N_noxref_10_c_2210_n ) capacitor c=0.019837f \
 //x=20.235 //y=3.7 //x2=12.95 //y2=2.08
cc_1118 ( N_noxref_6_c_1255_n N_noxref_10_c_2239_n ) capacitor c=0.0251381f \
 //x=20.235 //y=3.7 //x2=18.5 //y2=4.07
cc_1119 ( N_noxref_6_c_1258_n N_noxref_10_c_2239_n ) capacitor c=0.0142589f \
 //x=20.35 //y=2.08 //x2=18.5 //y2=4.07
cc_1120 ( N_noxref_6_c_1253_n N_noxref_10_c_2241_n ) capacitor c=0.00221254f \
 //x=8.765 //y=3.7 //x2=8.135 //y2=4.07
cc_1121 ( N_noxref_6_c_1286_n N_noxref_10_c_2241_n ) capacitor c=3.94811e-19 \
 //x=8.88 //y=3.7 //x2=8.135 //y2=4.07
cc_1122 ( N_noxref_6_c_1457_p N_noxref_10_c_2241_n ) capacitor c=2.67208e-19 \
 //x=8.1 //y=5.155 //x2=8.135 //y2=4.07
cc_1123 ( N_noxref_6_c_1278_n N_noxref_10_M28_noxref_g ) capacitor c=0.01736f \
 //x=8.015 //y=5.155 //x2=7.88 //y2=6.02
cc_1124 ( N_noxref_6_M28_noxref_d N_noxref_10_M28_noxref_g ) capacitor \
 c=0.0180032f //x=7.955 //y=5.02 //x2=7.88 //y2=6.02
cc_1125 ( N_noxref_6_c_1282_n N_noxref_10_M29_noxref_g ) capacitor \
 c=0.0194981f //x=8.795 //y=5.155 //x2=8.32 //y2=6.02
cc_1126 ( N_noxref_6_M28_noxref_d N_noxref_10_M29_noxref_g ) capacitor \
 c=0.0194246f //x=7.955 //y=5.02 //x2=8.32 //y2=6.02
cc_1127 ( N_noxref_6_M5_noxref_d N_noxref_10_c_2330_n ) capacitor \
 c=0.00217566f //x=8.205 //y=0.915 //x2=8.13 //y2=0.915
cc_1128 ( N_noxref_6_M5_noxref_d N_noxref_10_c_2331_n ) capacitor c=0.0034598f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=1.26
cc_1129 ( N_noxref_6_M5_noxref_d N_noxref_10_c_2332_n ) capacitor \
 c=0.00544291f //x=8.205 //y=0.915 //x2=8.13 //y2=1.57
cc_1130 ( N_noxref_6_M5_noxref_d N_noxref_10_c_2370_n ) capacitor \
 c=0.00241102f //x=8.205 //y=0.915 //x2=8.505 //y2=0.76
cc_1131 ( N_noxref_6_c_1257_n N_noxref_10_c_2371_n ) capacitor c=0.00359704f \
 //x=8.795 //y=1.665 //x2=8.505 //y2=1.415
cc_1132 ( N_noxref_6_M5_noxref_d N_noxref_10_c_2371_n ) capacitor c=0.0140297f \
 //x=8.205 //y=0.915 //x2=8.505 //y2=1.415
cc_1133 ( N_noxref_6_M5_noxref_d N_noxref_10_c_2373_n ) capacitor \
 c=0.00219619f //x=8.205 //y=0.915 //x2=8.66 //y2=0.915
cc_1134 ( N_noxref_6_c_1257_n N_noxref_10_c_2374_n ) capacitor c=0.00457401f \
 //x=8.795 //y=1.665 //x2=8.66 //y2=1.26
cc_1135 ( N_noxref_6_M5_noxref_d N_noxref_10_c_2374_n ) capacitor \
 c=0.00603828f //x=8.205 //y=0.915 //x2=8.66 //y2=1.26
cc_1136 ( N_noxref_6_c_1286_n N_noxref_10_c_2275_n ) capacitor c=0.00877984f \
 //x=8.88 //y=3.7 //x2=8.14 //y2=2.08
cc_1137 ( N_noxref_6_c_1286_n N_noxref_10_c_2335_n ) capacitor c=0.00283672f \
 //x=8.88 //y=3.7 //x2=8.14 //y2=1.915
cc_1138 ( N_noxref_6_M5_noxref_d N_noxref_10_c_2335_n ) capacitor \
 c=0.00661782f //x=8.205 //y=0.915 //x2=8.14 //y2=1.915
cc_1139 ( N_noxref_6_c_1282_n N_noxref_10_c_2336_n ) capacitor c=0.00201851f \
 //x=8.795 //y=5.155 //x2=8.14 //y2=4.7
cc_1140 ( N_noxref_6_c_1286_n N_noxref_10_c_2336_n ) capacitor c=0.013844f \
 //x=8.88 //y=3.7 //x2=8.14 //y2=4.7
cc_1141 ( N_noxref_6_c_1457_p N_noxref_10_c_2336_n ) capacitor c=0.0046827f \
 //x=8.1 //y=5.155 //x2=8.14 //y2=4.7
cc_1142 ( N_noxref_6_c_1255_n N_Q_c_2588_n ) capacitor c=0.00740361f \
 //x=20.235 //y=3.7 //x2=22.685 //y2=3.7
cc_1143 ( N_noxref_6_c_1258_n N_Q_c_2550_n ) capacitor c=0.00135527f //x=20.35 \
 //y=2.08 //x2=22.57 //y2=2.08
cc_1144 ( N_noxref_6_c_1256_n N_D_c_2706_n ) capacitor c=0.00181863f //x=3.33 \
 //y=2.08 //x2=1.11 //y2=2.08
cc_1145 ( N_noxref_6_c_1256_n N_noxref_14_c_2814_n ) capacitor c=0.00209081f \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_1146 ( N_noxref_6_c_1342_n N_noxref_14_c_2814_n ) capacitor c=0.0194423f \
 //x=3.32 //y=0.915 //x2=3.985 //y2=0.54
cc_1147 ( N_noxref_6_c_1348_n N_noxref_14_c_2814_n ) capacitor c=0.00656458f \
 //x=3.85 //y=0.915 //x2=3.985 //y2=0.54
cc_1148 ( N_noxref_6_c_1351_n N_noxref_14_c_2814_n ) capacitor c=2.20712e-19 \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_1149 ( N_noxref_6_c_1343_n N_noxref_14_c_2825_n ) capacitor c=0.00538829f \
 //x=3.32 //y=1.26 //x2=3.1 //y2=0.995
cc_1150 ( N_noxref_6_c_1342_n N_noxref_14_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=0.915 //x2=2.965 //y2=0.375
cc_1151 ( N_noxref_6_c_1344_n N_noxref_14_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=1.57 //x2=2.965 //y2=0.375
cc_1152 ( N_noxref_6_c_1348_n N_noxref_14_M2_noxref_s ) capacitor c=0.0143002f \
 //x=3.85 //y=0.915 //x2=2.965 //y2=0.375
cc_1153 ( N_noxref_6_c_1349_n N_noxref_14_M2_noxref_s ) capacitor \
 c=0.00290153f //x=3.85 //y=1.26 //x2=2.965 //y2=0.375
cc_1154 ( N_noxref_6_M5_noxref_d N_noxref_15_M3_noxref_s ) capacitor \
 c=0.00309936f //x=8.205 //y=0.915 //x2=5.265 //y2=0.375
cc_1155 ( N_noxref_6_c_1257_n N_noxref_16_c_2919_n ) capacitor c=0.00464321f \
 //x=8.795 //y=1.665 //x2=8.795 //y2=0.54
cc_1156 ( N_noxref_6_M5_noxref_d N_noxref_16_c_2919_n ) capacitor c=0.0117414f \
 //x=8.205 //y=0.915 //x2=8.795 //y2=0.54
cc_1157 ( N_noxref_6_c_1335_n N_noxref_16_c_2945_n ) capacitor c=0.0200405f \
 //x=8.48 //y=1.665 //x2=7.91 //y2=0.995
cc_1158 ( N_noxref_6_M5_noxref_d N_noxref_16_M4_noxref_d ) capacitor \
 c=5.27807e-19 //x=8.205 //y=0.915 //x2=6.67 //y2=0.91
cc_1159 ( N_noxref_6_c_1257_n N_noxref_16_M5_noxref_s ) capacitor c=0.0205309f \
 //x=8.795 //y=1.665 //x2=7.775 //y2=0.375
cc_1160 ( N_noxref_6_M5_noxref_d N_noxref_16_M5_noxref_s ) capacitor \
 c=0.0426368f //x=8.205 //y=0.915 //x2=7.775 //y2=0.375
cc_1161 ( N_noxref_6_c_1257_n N_noxref_17_c_2983_n ) capacitor c=3.84569e-19 \
 //x=8.795 //y=1.665 //x2=10.21 //y2=1.505
cc_1162 ( N_noxref_6_M5_noxref_d N_noxref_17_M6_noxref_s ) capacitor \
 c=2.55333e-19 //x=8.205 //y=0.915 //x2=10.075 //y2=0.375
cc_1163 ( N_noxref_6_c_1263_n N_noxref_21_c_3195_n ) capacitor c=0.0034165f \
 //x=20.05 //y=1.915 //x2=19.83 //y2=1.505
cc_1164 ( N_noxref_6_c_1258_n N_noxref_21_c_3179_n ) capacitor c=0.0122624f \
 //x=20.35 //y=2.08 //x2=20.715 //y2=1.59
cc_1165 ( N_noxref_6_c_1262_n N_noxref_21_c_3179_n ) capacitor c=0.00703864f \
 //x=20.05 //y=1.53 //x2=20.715 //y2=1.59
cc_1166 ( N_noxref_6_c_1263_n N_noxref_21_c_3179_n ) capacitor c=0.0215834f \
 //x=20.05 //y=1.915 //x2=20.715 //y2=1.59
cc_1167 ( N_noxref_6_c_1265_n N_noxref_21_c_3179_n ) capacitor c=0.00708583f \
 //x=20.425 //y=1.375 //x2=20.715 //y2=1.59
cc_1168 ( N_noxref_6_c_1268_n N_noxref_21_c_3179_n ) capacitor c=0.00698822f \
 //x=20.58 //y=1.22 //x2=20.715 //y2=1.59
cc_1169 ( N_noxref_6_c_1259_n N_noxref_21_M12_noxref_s ) capacitor \
 c=0.0327271f //x=20.05 //y=0.875 //x2=19.695 //y2=0.375
cc_1170 ( N_noxref_6_c_1262_n N_noxref_21_M12_noxref_s ) capacitor \
 c=7.99997e-19 //x=20.05 //y=1.53 //x2=19.695 //y2=0.375
cc_1171 ( N_noxref_6_c_1263_n N_noxref_21_M12_noxref_s ) capacitor \
 c=0.00122123f //x=20.05 //y=1.915 //x2=19.695 //y2=0.375
cc_1172 ( N_noxref_6_c_1266_n N_noxref_21_M12_noxref_s ) capacitor \
 c=0.0121427f //x=20.58 //y=0.875 //x2=19.695 //y2=0.375
cc_1173 ( N_RN_c_1518_n QN ) capacitor c=0.00326636f //x=21.46 //y=2.08 \
 //x2=23.31 //y2=2.22
cc_1174 ( N_RN_c_1536_n N_QN_c_1838_n ) capacitor c=0.00241768f //x=21.345 \
 //y=4.44 //x2=21.565 //y2=5.155
cc_1175 ( N_RN_c_1518_n N_QN_c_1838_n ) capacitor c=0.014564f //x=21.46 \
 //y=2.08 //x2=21.565 //y2=5.155
cc_1176 ( N_RN_M44_noxref_g N_QN_c_1838_n ) capacitor c=0.016514f //x=21.43 \
 //y=6.02 //x2=21.565 //y2=5.155
cc_1177 ( N_RN_c_1663_n N_QN_c_1838_n ) capacitor c=0.00322046f //x=21.46 \
 //y=4.7 //x2=21.565 //y2=5.155
cc_1178 ( N_RN_c_1536_n N_QN_c_1842_n ) capacitor c=0.0219114f //x=21.345 \
 //y=4.44 //x2=20.855 //y2=5.155
cc_1179 ( N_RN_M45_noxref_g N_QN_c_1844_n ) capacitor c=0.0184045f //x=21.87 \
 //y=6.02 //x2=22.445 //y2=5.155
cc_1180 ( N_RN_c_1536_n N_QN_c_1887_n ) capacitor c=0.00101864f //x=21.345 \
 //y=4.44 //x2=21.65 //y2=5.155
cc_1181 ( N_RN_c_1674_p N_QN_c_1887_n ) capacitor c=0.00427771f //x=21.795 \
 //y=4.79 //x2=21.65 //y2=5.155
cc_1182 ( N_RN_M44_noxref_g N_QN_M44_noxref_d ) capacitor c=0.0180032f \
 //x=21.43 //y=6.02 //x2=21.505 //y2=5.02
cc_1183 ( N_RN_M45_noxref_g N_QN_M44_noxref_d ) capacitor c=0.0180032f \
 //x=21.87 //y=6.02 //x2=21.505 //y2=5.02
cc_1184 ( N_RN_c_1536_n N_SN_c_1980_n ) capacitor c=0.00602392f //x=21.345 \
 //y=4.44 //x2=26.155 //y2=2.59
cc_1185 ( N_RN_c_1517_n N_SN_c_1980_n ) capacitor c=0.0253613f //x=17.76 \
 //y=2.08 //x2=26.155 //y2=2.59
cc_1186 ( N_RN_c_1518_n N_SN_c_1980_n ) capacitor c=0.0273718f //x=21.46 \
 //y=2.08 //x2=26.155 //y2=2.59
cc_1187 ( N_RN_c_1659_n N_SN_c_1980_n ) capacitor c=0.00233308f //x=21.55 \
 //y=1.915 //x2=26.155 //y2=2.59
cc_1188 ( N_RN_c_1606_n N_SN_c_1980_n ) capacitor c=0.00232725f //x=17.76 \
 //y=2.08 //x2=26.155 //y2=2.59
cc_1189 ( N_RN_c_1514_n N_SN_c_1991_n ) capacitor c=0.0210462f //x=17.645 \
 //y=4.44 //x2=11.84 //y2=2.08
cc_1190 ( N_RN_c_1514_n N_SN_c_2039_n ) capacitor c=0.0085986f //x=17.645 \
 //y=4.44 //x2=12.175 //y2=4.79
cc_1191 ( N_RN_c_1514_n N_SN_c_2024_n ) capacitor c=0.00293313f //x=17.645 \
 //y=4.44 //x2=11.84 //y2=4.7
cc_1192 ( N_RN_c_1514_n N_noxref_10_c_2214_n ) capacitor c=0.398867f \
 //x=17.645 //y=4.44 //x2=12.835 //y2=4.07
cc_1193 ( N_RN_c_1514_n N_noxref_10_c_2308_n ) capacitor c=0.0291412f \
 //x=17.645 //y=4.44 //x2=8.25 //y2=4.07
cc_1194 ( N_RN_c_1514_n N_noxref_10_c_2215_n ) capacitor c=0.398418f \
 //x=17.645 //y=4.44 //x2=18.385 //y2=4.07
cc_1195 ( N_RN_c_1536_n N_noxref_10_c_2215_n ) capacitor c=0.0442407f \
 //x=21.345 //y=4.44 //x2=18.385 //y2=4.07
cc_1196 ( N_RN_c_1542_n N_noxref_10_c_2215_n ) capacitor c=0.0268623f \
 //x=17.875 //y=4.44 //x2=18.385 //y2=4.07
cc_1197 ( N_RN_c_1517_n N_noxref_10_c_2215_n ) capacitor c=0.0198123f \
 //x=17.76 //y=2.08 //x2=18.385 //y2=4.07
cc_1198 ( N_RN_c_1514_n N_noxref_10_c_2278_n ) capacitor c=0.0265199f \
 //x=17.645 //y=4.44 //x2=13.065 //y2=4.07
cc_1199 ( N_RN_c_1536_n N_noxref_10_c_2216_n ) capacitor c=0.268165f \
 //x=21.345 //y=4.44 //x2=27.265 //y2=4.07
cc_1200 ( N_RN_c_1518_n N_noxref_10_c_2216_n ) capacitor c=0.0256971f \
 //x=21.46 //y=2.08 //x2=27.265 //y2=4.07
cc_1201 ( N_RN_c_1674_p N_noxref_10_c_2216_n ) capacitor c=0.00483006f \
 //x=21.795 //y=4.79 //x2=27.265 //y2=4.07
cc_1202 ( N_RN_c_1536_n N_noxref_10_c_2223_n ) capacitor c=0.0265915f \
 //x=21.345 //y=4.44 //x2=18.615 //y2=4.07
cc_1203 ( N_RN_c_1517_n N_noxref_10_c_2223_n ) capacitor c=0.00179385f \
 //x=17.76 //y=2.08 //x2=18.615 //y2=4.07
cc_1204 ( N_RN_c_1514_n N_noxref_10_c_2317_n ) capacitor c=0.0197679f \
 //x=17.645 //y=4.44 //x2=8.14 //y2=4.7
cc_1205 ( N_RN_c_1514_n N_noxref_10_c_2210_n ) capacitor c=0.0218403f \
 //x=17.645 //y=4.44 //x2=12.95 //y2=2.08
cc_1206 ( N_RN_c_1514_n N_noxref_10_c_2225_n ) capacitor c=0.0311077f \
 //x=17.645 //y=4.44 //x2=16.755 //y2=5.155
cc_1207 ( N_RN_c_1514_n N_noxref_10_c_2229_n ) capacitor c=0.0230136f \
 //x=17.645 //y=4.44 //x2=16.045 //y2=5.155
cc_1208 ( N_RN_M40_noxref_g N_noxref_10_c_2231_n ) capacitor c=0.01736f \
 //x=17.5 //y=6.02 //x2=17.635 //y2=5.155
cc_1209 ( N_RN_c_1536_n N_noxref_10_c_2235_n ) capacitor c=0.0173131f \
 //x=21.345 //y=4.44 //x2=18.415 //y2=5.155
cc_1210 ( N_RN_c_1542_n N_noxref_10_c_2235_n ) capacitor c=0.00124956f \
 //x=17.875 //y=4.44 //x2=18.415 //y2=5.155
cc_1211 ( N_RN_M41_noxref_g N_noxref_10_c_2235_n ) capacitor c=0.0194918f \
 //x=17.94 //y=6.02 //x2=18.415 //y2=5.155
cc_1212 ( N_RN_c_1609_n N_noxref_10_c_2235_n ) capacitor c=0.00201851f \
 //x=17.76 //y=4.7 //x2=18.415 //y2=5.155
cc_1213 ( N_RN_c_1706_p N_noxref_10_c_2211_n ) capacitor c=0.00359704f \
 //x=18.125 //y=1.415 //x2=18.415 //y2=1.665
cc_1214 ( N_RN_c_1707_p N_noxref_10_c_2211_n ) capacitor c=0.00457401f \
 //x=18.28 //y=1.26 //x2=18.415 //y2=1.665
cc_1215 ( N_RN_c_1536_n N_noxref_10_c_2239_n ) capacitor c=0.022862f \
 //x=21.345 //y=4.44 //x2=18.5 //y2=4.07
cc_1216 ( N_RN_c_1542_n N_noxref_10_c_2239_n ) capacitor c=0.00118555f \
 //x=17.875 //y=4.44 //x2=18.5 //y2=4.07
cc_1217 ( N_RN_c_1517_n N_noxref_10_c_2239_n ) capacitor c=0.081883f //x=17.76 \
 //y=2.08 //x2=18.5 //y2=4.07
cc_1218 ( N_RN_c_1518_n N_noxref_10_c_2239_n ) capacitor c=7.03136e-19 \
 //x=21.46 //y=2.08 //x2=18.5 //y2=4.07
cc_1219 ( N_RN_c_1606_n N_noxref_10_c_2239_n ) capacitor c=0.00877984f \
 //x=17.76 //y=2.08 //x2=18.5 //y2=4.07
cc_1220 ( N_RN_c_1608_n N_noxref_10_c_2239_n ) capacitor c=0.00283672f \
 //x=17.76 //y=1.915 //x2=18.5 //y2=4.07
cc_1221 ( N_RN_c_1609_n N_noxref_10_c_2239_n ) capacitor c=0.013693f //x=17.76 \
 //y=4.7 //x2=18.5 //y2=4.07
cc_1222 ( N_RN_c_1514_n N_noxref_10_c_2241_n ) capacitor c=0.00215288f \
 //x=17.645 //y=4.44 //x2=8.135 //y2=4.07
cc_1223 ( N_RN_c_1542_n N_noxref_10_c_2413_n ) capacitor c=0.00125695f \
 //x=17.875 //y=4.44 //x2=17.72 //y2=5.155
cc_1224 ( N_RN_c_1517_n N_noxref_10_c_2413_n ) capacitor c=0.0165698f \
 //x=17.76 //y=2.08 //x2=17.72 //y2=5.155
cc_1225 ( N_RN_c_1609_n N_noxref_10_c_2413_n ) capacitor c=0.00475592f \
 //x=17.76 //y=4.7 //x2=17.72 //y2=5.155
cc_1226 ( N_RN_c_1514_n N_noxref_10_c_2336_n ) capacitor c=0.011194f \
 //x=17.645 //y=4.44 //x2=8.14 //y2=4.7
cc_1227 ( N_RN_c_1514_n N_noxref_10_c_2303_n ) capacitor c=0.0111881f \
 //x=17.645 //y=4.44 //x2=12.95 //y2=4.7
cc_1228 ( N_RN_c_1603_n N_noxref_10_M11_noxref_d ) capacitor c=0.00217566f \
 //x=17.75 //y=0.915 //x2=17.825 //y2=0.915
cc_1229 ( N_RN_c_1604_n N_noxref_10_M11_noxref_d ) capacitor c=0.0034598f \
 //x=17.75 //y=1.26 //x2=17.825 //y2=0.915
cc_1230 ( N_RN_c_1605_n N_noxref_10_M11_noxref_d ) capacitor c=0.00544291f \
 //x=17.75 //y=1.57 //x2=17.825 //y2=0.915
cc_1231 ( N_RN_c_1724_p N_noxref_10_M11_noxref_d ) capacitor c=0.00241102f \
 //x=18.125 //y=0.76 //x2=17.825 //y2=0.915
cc_1232 ( N_RN_c_1706_p N_noxref_10_M11_noxref_d ) capacitor c=0.0140297f \
 //x=18.125 //y=1.415 //x2=17.825 //y2=0.915
cc_1233 ( N_RN_c_1726_p N_noxref_10_M11_noxref_d ) capacitor c=0.00219619f \
 //x=18.28 //y=0.915 //x2=17.825 //y2=0.915
cc_1234 ( N_RN_c_1707_p N_noxref_10_M11_noxref_d ) capacitor c=0.00603828f \
 //x=18.28 //y=1.26 //x2=17.825 //y2=0.915
cc_1235 ( N_RN_c_1608_n N_noxref_10_M11_noxref_d ) capacitor c=0.00661782f \
 //x=17.76 //y=1.915 //x2=17.825 //y2=0.915
cc_1236 ( N_RN_M40_noxref_g N_noxref_10_M40_noxref_d ) capacitor c=0.0180032f \
 //x=17.5 //y=6.02 //x2=17.575 //y2=5.02
cc_1237 ( N_RN_M41_noxref_g N_noxref_10_M40_noxref_d ) capacitor c=0.0194246f \
 //x=17.94 //y=6.02 //x2=17.575 //y2=5.02
cc_1238 ( N_RN_c_1518_n N_Q_c_2588_n ) capacitor c=0.0027353f //x=21.46 \
 //y=2.08 //x2=22.685 //y2=3.7
cc_1239 ( N_RN_c_1536_n N_Q_c_2550_n ) capacitor c=0.00551083f //x=21.345 \
 //y=4.44 //x2=22.57 //y2=2.08
cc_1240 ( N_RN_c_1518_n N_Q_c_2550_n ) capacitor c=0.0502572f //x=21.46 \
 //y=2.08 //x2=22.57 //y2=2.08
cc_1241 ( N_RN_c_1659_n N_Q_c_2550_n ) capacitor c=0.0023343f //x=21.55 \
 //y=1.915 //x2=22.57 //y2=2.08
cc_1242 ( N_RN_c_1663_n N_Q_c_2550_n ) capacitor c=0.00142741f //x=21.46 \
 //y=4.7 //x2=22.57 //y2=2.08
cc_1243 ( N_RN_M44_noxref_g N_Q_M46_noxref_g ) capacitor c=0.0101598f \
 //x=21.43 //y=6.02 //x2=22.31 //y2=6.02
cc_1244 ( N_RN_M45_noxref_g N_Q_M46_noxref_g ) capacitor c=0.0602553f \
 //x=21.87 //y=6.02 //x2=22.31 //y2=6.02
cc_1245 ( N_RN_M45_noxref_g N_Q_M47_noxref_g ) capacitor c=0.0101598f \
 //x=21.87 //y=6.02 //x2=22.75 //y2=6.02
cc_1246 ( N_RN_c_1656_n N_Q_c_2598_n ) capacitor c=0.00456962f //x=21.55 \
 //y=0.91 //x2=22.56 //y2=0.915
cc_1247 ( N_RN_c_1657_n N_Q_c_2599_n ) capacitor c=0.00438372f //x=21.55 \
 //y=1.22 //x2=22.56 //y2=1.26
cc_1248 ( N_RN_c_1658_n N_Q_c_2600_n ) capacitor c=0.00438372f //x=21.55 \
 //y=1.45 //x2=22.56 //y2=1.57
cc_1249 ( N_RN_c_1518_n N_Q_c_2601_n ) capacitor c=0.00228632f //x=21.46 \
 //y=2.08 //x2=22.57 //y2=2.08
cc_1250 ( N_RN_c_1659_n N_Q_c_2601_n ) capacitor c=0.00933826f //x=21.55 \
 //y=1.915 //x2=22.57 //y2=2.08
cc_1251 ( N_RN_c_1659_n N_Q_c_2603_n ) capacitor c=0.00438372f //x=21.55 \
 //y=1.915 //x2=22.57 //y2=1.915
cc_1252 ( N_RN_c_1518_n N_Q_c_2604_n ) capacitor c=0.00218014f //x=21.46 \
 //y=2.08 //x2=22.57 //y2=4.7
cc_1253 ( N_RN_c_1674_p N_Q_c_2604_n ) capacitor c=0.0611812f //x=21.795 \
 //y=4.79 //x2=22.57 //y2=4.7
cc_1254 ( N_RN_c_1663_n N_Q_c_2604_n ) capacitor c=0.00487508f //x=21.46 \
 //y=4.7 //x2=22.57 //y2=4.7
cc_1255 ( N_RN_c_1515_n N_D_c_2706_n ) capacitor c=0.00551083f //x=2.335 \
 //y=4.44 //x2=1.11 //y2=2.08
cc_1256 ( N_RN_c_1516_n N_D_c_2706_n ) capacitor c=0.0563464f //x=2.22 \
 //y=2.08 //x2=1.11 //y2=2.08
cc_1257 ( N_RN_c_1647_n N_D_c_2706_n ) capacitor c=0.00231304f //x=2.31 \
 //y=1.915 //x2=1.11 //y2=2.08
cc_1258 ( N_RN_c_1579_n N_D_c_2706_n ) capacitor c=0.00183762f //x=2.22 \
 //y=4.7 //x2=1.11 //y2=2.08
cc_1259 ( N_RN_M20_noxref_g N_D_M18_noxref_g ) capacitor c=0.0105869f //x=2.19 \
 //y=6.02 //x2=1.31 //y2=6.02
cc_1260 ( N_RN_M20_noxref_g N_D_M19_noxref_g ) capacitor c=0.10632f //x=2.19 \
 //y=6.02 //x2=1.75 //y2=6.02
cc_1261 ( N_RN_M21_noxref_g N_D_M19_noxref_g ) capacitor c=0.0101598f //x=2.63 \
 //y=6.02 //x2=1.75 //y2=6.02
cc_1262 ( N_RN_c_1755_p N_D_c_2707_n ) capacitor c=5.72482e-19 //x=1.785 \
 //y=0.91 //x2=0.81 //y2=0.875
cc_1263 ( N_RN_c_1755_p N_D_c_2709_n ) capacitor c=0.00149976f //x=1.785 \
 //y=0.91 //x2=0.81 //y2=1.22
cc_1264 ( N_RN_c_1757_p N_D_c_2710_n ) capacitor c=0.00111227f //x=1.785 \
 //y=1.22 //x2=0.81 //y2=1.53
cc_1265 ( N_RN_c_1516_n N_D_c_2711_n ) capacitor c=0.00238338f //x=2.22 \
 //y=2.08 //x2=0.81 //y2=1.915
cc_1266 ( N_RN_c_1647_n N_D_c_2711_n ) capacitor c=0.00964411f //x=2.31 \
 //y=1.915 //x2=0.81 //y2=1.915
cc_1267 ( N_RN_c_1755_p N_D_c_2714_n ) capacitor c=0.0160123f //x=1.785 \
 //y=0.91 //x2=1.34 //y2=0.875
cc_1268 ( N_RN_c_1644_n N_D_c_2714_n ) capacitor c=0.00103227f //x=2.31 \
 //y=0.91 //x2=1.34 //y2=0.875
cc_1269 ( N_RN_c_1757_p N_D_c_2716_n ) capacitor c=0.0124075f //x=1.785 \
 //y=1.22 //x2=1.34 //y2=1.22
cc_1270 ( N_RN_c_1645_n N_D_c_2716_n ) capacitor c=0.0010154f //x=2.31 \
 //y=1.22 //x2=1.34 //y2=1.22
cc_1271 ( N_RN_c_1646_n N_D_c_2716_n ) capacitor c=9.23422e-19 //x=2.31 \
 //y=1.45 //x2=1.34 //y2=1.22
cc_1272 ( N_RN_c_1516_n N_D_c_2729_n ) capacitor c=0.00147352f //x=2.22 \
 //y=2.08 //x2=1.675 //y2=4.79
cc_1273 ( N_RN_c_1579_n N_D_c_2729_n ) capacitor c=0.0168581f //x=2.22 //y=4.7 \
 //x2=1.675 //y2=4.79
cc_1274 ( N_RN_c_1516_n N_D_c_2724_n ) capacitor c=0.00141297f //x=2.22 \
 //y=2.08 //x2=1.385 //y2=4.79
cc_1275 ( N_RN_c_1579_n N_D_c_2724_n ) capacitor c=0.00484466f //x=2.22 \
 //y=4.7 //x2=1.385 //y2=4.79
cc_1276 ( N_RN_c_1755_p N_noxref_13_c_2769_n ) capacitor c=0.0167228f \
 //x=1.785 //y=0.91 //x2=2.445 //y2=0.54
cc_1277 ( N_RN_c_1644_n N_noxref_13_c_2769_n ) capacitor c=0.00534519f \
 //x=2.31 //y=0.91 //x2=2.445 //y2=0.54
cc_1278 ( N_RN_c_1514_n N_noxref_13_c_2781_n ) capacitor c=0.00136783f \
 //x=17.645 //y=4.44 //x2=2.445 //y2=1.59
cc_1279 ( N_RN_c_1515_n N_noxref_13_c_2781_n ) capacitor c=0.00102601f \
 //x=2.335 //y=4.44 //x2=2.445 //y2=1.59
cc_1280 ( N_RN_c_1516_n N_noxref_13_c_2781_n ) capacitor c=0.012374f //x=2.22 \
 //y=2.08 //x2=2.445 //y2=1.59
cc_1281 ( N_RN_c_1757_p N_noxref_13_c_2781_n ) capacitor c=0.0153476f \
 //x=1.785 //y=1.22 //x2=2.445 //y2=1.59
cc_1282 ( N_RN_c_1647_n N_noxref_13_c_2781_n ) capacitor c=0.0231679f //x=2.31 \
 //y=1.915 //x2=2.445 //y2=1.59
cc_1283 ( N_RN_c_1514_n N_noxref_13_M0_noxref_s ) capacitor c=9.40017e-19 \
 //x=17.645 //y=4.44 //x2=0.455 //y2=0.375
cc_1284 ( N_RN_c_1755_p N_noxref_13_M0_noxref_s ) capacitor c=0.00798959f \
 //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_1285 ( N_RN_c_1646_n N_noxref_13_M0_noxref_s ) capacitor c=0.00212176f \
 //x=2.31 //y=1.45 //x2=0.455 //y2=0.375
cc_1286 ( N_RN_c_1647_n N_noxref_13_M0_noxref_s ) capacitor c=0.00298115f \
 //x=2.31 //y=1.915 //x2=0.455 //y2=0.375
cc_1287 ( N_RN_c_1514_n N_noxref_14_c_2808_n ) capacitor c=0.00133627f \
 //x=17.645 //y=4.44 //x2=3.015 //y2=0.995
cc_1288 ( N_RN_c_1781_p N_noxref_14_c_2808_n ) capacitor c=2.14837e-19 \
 //x=2.155 //y=0.755 //x2=3.015 //y2=0.995
cc_1289 ( N_RN_c_1644_n N_noxref_14_c_2808_n ) capacitor c=0.00123426f \
 //x=2.31 //y=0.91 //x2=3.015 //y2=0.995
cc_1290 ( N_RN_c_1645_n N_noxref_14_c_2808_n ) capacitor c=0.0129288f //x=2.31 \
 //y=1.22 //x2=3.015 //y2=0.995
cc_1291 ( N_RN_c_1646_n N_noxref_14_c_2808_n ) capacitor c=0.00142359f \
 //x=2.31 //y=1.45 //x2=3.015 //y2=0.995
cc_1292 ( N_RN_c_1755_p N_noxref_14_M1_noxref_d ) capacitor c=0.00223875f \
 //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_1293 ( N_RN_c_1757_p N_noxref_14_M1_noxref_d ) capacitor c=0.00262485f \
 //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_1294 ( N_RN_c_1781_p N_noxref_14_M1_noxref_d ) capacitor c=0.00220746f \
 //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_1295 ( N_RN_c_1788_p N_noxref_14_M1_noxref_d ) capacitor c=0.00194798f \
 //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_1296 ( N_RN_c_1644_n N_noxref_14_M1_noxref_d ) capacitor c=0.00198465f \
 //x=2.31 //y=0.91 //x2=1.86 //y2=0.91
cc_1297 ( N_RN_c_1645_n N_noxref_14_M1_noxref_d ) capacitor c=0.00128384f \
 //x=2.31 //y=1.22 //x2=1.86 //y2=0.91
cc_1298 ( N_RN_c_1514_n N_noxref_14_M2_noxref_s ) capacitor c=9.61379e-19 \
 //x=17.645 //y=4.44 //x2=2.965 //y2=0.375
cc_1299 ( N_RN_c_1644_n N_noxref_14_M2_noxref_s ) capacitor c=7.21316e-19 \
 //x=2.31 //y=0.91 //x2=2.965 //y2=0.375
cc_1300 ( N_RN_c_1645_n N_noxref_14_M2_noxref_s ) capacitor c=0.00348171f \
 //x=2.31 //y=1.22 //x2=2.965 //y2=0.375
cc_1301 ( N_RN_c_1517_n N_noxref_20_c_3131_n ) capacitor c=0.0020642f \
 //x=17.76 //y=2.08 //x2=18.415 //y2=0.54
cc_1302 ( N_RN_c_1603_n N_noxref_20_c_3131_n ) capacitor c=0.0194423f \
 //x=17.75 //y=0.915 //x2=18.415 //y2=0.54
cc_1303 ( N_RN_c_1726_p N_noxref_20_c_3131_n ) capacitor c=0.00656458f \
 //x=18.28 //y=0.915 //x2=18.415 //y2=0.54
cc_1304 ( N_RN_c_1606_n N_noxref_20_c_3131_n ) capacitor c=2.20712e-19 \
 //x=17.76 //y=2.08 //x2=18.415 //y2=0.54
cc_1305 ( N_RN_c_1604_n N_noxref_20_c_3156_n ) capacitor c=0.00538829f \
 //x=17.75 //y=1.26 //x2=17.53 //y2=0.995
cc_1306 ( N_RN_c_1603_n N_noxref_20_M11_noxref_s ) capacitor c=0.00538829f \
 //x=17.75 //y=0.915 //x2=17.395 //y2=0.375
cc_1307 ( N_RN_c_1605_n N_noxref_20_M11_noxref_s ) capacitor c=0.00538829f \
 //x=17.75 //y=1.57 //x2=17.395 //y2=0.375
cc_1308 ( N_RN_c_1726_p N_noxref_20_M11_noxref_s ) capacitor c=0.0143002f \
 //x=18.28 //y=0.915 //x2=17.395 //y2=0.375
cc_1309 ( N_RN_c_1707_p N_noxref_20_M11_noxref_s ) capacitor c=0.00290153f \
 //x=18.28 //y=1.26 //x2=17.395 //y2=0.375
cc_1310 ( N_RN_c_1651_n N_noxref_21_c_3186_n ) capacitor c=0.0167228f \
 //x=21.025 //y=0.91 //x2=21.685 //y2=0.54
cc_1311 ( N_RN_c_1656_n N_noxref_21_c_3186_n ) capacitor c=0.00534519f \
 //x=21.55 //y=0.91 //x2=21.685 //y2=0.54
cc_1312 ( N_RN_c_1518_n N_noxref_21_c_3207_n ) capacitor c=0.012334f //x=21.46 \
 //y=2.08 //x2=21.685 //y2=1.59
cc_1313 ( N_RN_c_1654_n N_noxref_21_c_3207_n ) capacitor c=0.0153476f \
 //x=21.025 //y=1.22 //x2=21.685 //y2=1.59
cc_1314 ( N_RN_c_1659_n N_noxref_21_c_3207_n ) capacitor c=0.0219329f \
 //x=21.55 //y=1.915 //x2=21.685 //y2=1.59
cc_1315 ( N_RN_c_1651_n N_noxref_21_M12_noxref_s ) capacitor c=0.00798959f \
 //x=21.025 //y=0.91 //x2=19.695 //y2=0.375
cc_1316 ( N_RN_c_1658_n N_noxref_21_M12_noxref_s ) capacitor c=0.00212176f \
 //x=21.55 //y=1.45 //x2=19.695 //y2=0.375
cc_1317 ( N_RN_c_1659_n N_noxref_21_M12_noxref_s ) capacitor c=0.00298115f \
 //x=21.55 //y=1.915 //x2=19.695 //y2=0.375
cc_1318 ( N_RN_c_1811_p N_noxref_22_c_3229_n ) capacitor c=2.14837e-19 \
 //x=21.395 //y=0.755 //x2=22.255 //y2=0.995
cc_1319 ( N_RN_c_1656_n N_noxref_22_c_3229_n ) capacitor c=0.00123426f \
 //x=21.55 //y=0.91 //x2=22.255 //y2=0.995
cc_1320 ( N_RN_c_1657_n N_noxref_22_c_3229_n ) capacitor c=0.0129288f \
 //x=21.55 //y=1.22 //x2=22.255 //y2=0.995
cc_1321 ( N_RN_c_1658_n N_noxref_22_c_3229_n ) capacitor c=0.00142359f \
 //x=21.55 //y=1.45 //x2=22.255 //y2=0.995
cc_1322 ( N_RN_c_1651_n N_noxref_22_M13_noxref_d ) capacitor c=0.00223875f \
 //x=21.025 //y=0.91 //x2=21.1 //y2=0.91
cc_1323 ( N_RN_c_1654_n N_noxref_22_M13_noxref_d ) capacitor c=0.00262485f \
 //x=21.025 //y=1.22 //x2=21.1 //y2=0.91
cc_1324 ( N_RN_c_1811_p N_noxref_22_M13_noxref_d ) capacitor c=0.00220746f \
 //x=21.395 //y=0.755 //x2=21.1 //y2=0.91
cc_1325 ( N_RN_c_1818_p N_noxref_22_M13_noxref_d ) capacitor c=0.00194798f \
 //x=21.395 //y=1.375 //x2=21.1 //y2=0.91
cc_1326 ( N_RN_c_1656_n N_noxref_22_M13_noxref_d ) capacitor c=0.00198465f \
 //x=21.55 //y=0.91 //x2=21.1 //y2=0.91
cc_1327 ( N_RN_c_1657_n N_noxref_22_M13_noxref_d ) capacitor c=0.00128384f \
 //x=21.55 //y=1.22 //x2=21.1 //y2=0.91
cc_1328 ( N_RN_c_1656_n N_noxref_22_M14_noxref_s ) capacitor c=7.21316e-19 \
 //x=21.55 //y=0.91 //x2=22.205 //y2=0.375
cc_1329 ( N_RN_c_1657_n N_noxref_22_M14_noxref_s ) capacitor c=0.00348171f \
 //x=21.55 //y=1.22 //x2=22.205 //y2=0.375
cc_1330 ( N_QN_c_1823_n N_SN_c_1980_n ) capacitor c=0.0844361f //x=25.045 \
 //y=3.33 //x2=26.155 //y2=2.59
cc_1331 ( N_QN_c_1892_p N_SN_c_1980_n ) capacitor c=0.0133526f //x=23.425 \
 //y=3.33 //x2=26.155 //y2=2.59
cc_1332 ( QN N_SN_c_1980_n ) capacitor c=0.0236318f //x=23.31 //y=2.22 \
 //x2=26.155 //y2=2.59
cc_1333 ( N_QN_c_1894_p N_SN_c_1980_n ) capacitor c=0.0115788f //x=22.91 \
 //y=1.665 //x2=26.155 //y2=2.59
cc_1334 ( N_QN_c_1825_n N_SN_c_1980_n ) capacitor c=0.0262948f //x=25.16 \
 //y=2.08 //x2=26.155 //y2=2.59
cc_1335 ( N_QN_c_1830_n N_SN_c_1980_n ) capacitor c=0.00565297f //x=24.86 \
 //y=1.915 //x2=26.155 //y2=2.59
cc_1336 ( N_QN_c_1823_n N_SN_c_1992_n ) capacitor c=0.00520283f //x=25.045 \
 //y=3.33 //x2=26.27 //y2=2.08
cc_1337 ( QN N_SN_c_1992_n ) capacitor c=5.77178e-19 //x=23.31 //y=2.22 \
 //x2=26.27 //y2=2.08
cc_1338 ( N_QN_c_1825_n N_SN_c_1992_n ) capacitor c=0.0489575f //x=25.16 \
 //y=2.08 //x2=26.27 //y2=2.08
cc_1339 ( N_QN_c_1830_n N_SN_c_1992_n ) capacitor c=0.00238338f //x=24.86 \
 //y=1.915 //x2=26.27 //y2=2.08
cc_1340 ( N_QN_c_1901_p N_SN_c_1992_n ) capacitor c=0.00147352f //x=25.725 \
 //y=4.79 //x2=26.27 //y2=2.08
cc_1341 ( N_QN_c_1859_n N_SN_c_1992_n ) capacitor c=0.00142741f //x=25.435 \
 //y=4.79 //x2=26.27 //y2=2.08
cc_1342 ( N_QN_M48_noxref_g N_SN_M50_noxref_g ) capacitor c=0.0105869f \
 //x=25.36 //y=6.02 //x2=26.24 //y2=6.02
cc_1343 ( N_QN_M49_noxref_g N_SN_M50_noxref_g ) capacitor c=0.10632f //x=25.8 \
 //y=6.02 //x2=26.24 //y2=6.02
cc_1344 ( N_QN_M49_noxref_g N_SN_M51_noxref_g ) capacitor c=0.0101598f \
 //x=25.8 //y=6.02 //x2=26.68 //y2=6.02
cc_1345 ( N_QN_c_1826_n N_SN_c_2075_n ) capacitor c=5.72482e-19 //x=24.86 \
 //y=0.875 //x2=25.835 //y2=0.91
cc_1346 ( N_QN_c_1828_n N_SN_c_2075_n ) capacitor c=0.00149976f //x=24.86 \
 //y=1.22 //x2=25.835 //y2=0.91
cc_1347 ( N_QN_c_1833_n N_SN_c_2075_n ) capacitor c=0.0160123f //x=25.39 \
 //y=0.875 //x2=25.835 //y2=0.91
cc_1348 ( N_QN_c_1829_n N_SN_c_2078_n ) capacitor c=0.00111227f //x=24.86 \
 //y=1.53 //x2=25.835 //y2=1.22
cc_1349 ( N_QN_c_1835_n N_SN_c_2078_n ) capacitor c=0.0124075f //x=25.39 \
 //y=1.22 //x2=25.835 //y2=1.22
cc_1350 ( N_QN_c_1833_n N_SN_c_2080_n ) capacitor c=0.00103227f //x=25.39 \
 //y=0.875 //x2=26.36 //y2=0.91
cc_1351 ( N_QN_c_1835_n N_SN_c_2081_n ) capacitor c=0.0010154f //x=25.39 \
 //y=1.22 //x2=26.36 //y2=1.22
cc_1352 ( N_QN_c_1835_n N_SN_c_2082_n ) capacitor c=9.23422e-19 //x=25.39 \
 //y=1.22 //x2=26.36 //y2=1.45
cc_1353 ( N_QN_c_1825_n N_SN_c_2083_n ) capacitor c=0.00231304f //x=25.16 \
 //y=2.08 //x2=26.36 //y2=1.915
cc_1354 ( N_QN_c_1830_n N_SN_c_2083_n ) capacitor c=0.00964411f //x=24.86 \
 //y=1.915 //x2=26.36 //y2=1.915
cc_1355 ( N_QN_c_1825_n N_SN_c_2085_n ) capacitor c=0.00183762f //x=25.16 \
 //y=2.08 //x2=26.27 //y2=4.7
cc_1356 ( N_QN_c_1901_p N_SN_c_2085_n ) capacitor c=0.0168581f //x=25.725 \
 //y=4.79 //x2=26.27 //y2=4.7
cc_1357 ( N_QN_c_1859_n N_SN_c_2085_n ) capacitor c=0.00484466f //x=25.435 \
 //y=4.79 //x2=26.27 //y2=4.7
cc_1358 ( N_QN_c_1823_n N_noxref_10_c_2216_n ) capacitor c=0.0106705f \
 //x=25.045 //y=3.33 //x2=27.265 //y2=4.07
cc_1359 ( N_QN_c_1892_p N_noxref_10_c_2216_n ) capacitor c=7.97799e-19 \
 //x=23.425 //y=3.33 //x2=27.265 //y2=4.07
cc_1360 ( QN N_noxref_10_c_2216_n ) capacitor c=0.0232919f //x=23.31 //y=2.22 \
 //x2=27.265 //y2=4.07
cc_1361 ( N_QN_c_1848_n N_noxref_10_c_2216_n ) capacitor c=0.0138556f \
 //x=23.225 //y=5.155 //x2=27.265 //y2=4.07
cc_1362 ( N_QN_c_1825_n N_noxref_10_c_2216_n ) capacitor c=0.0234593f \
 //x=25.16 //y=2.08 //x2=27.265 //y2=4.07
cc_1363 ( N_QN_c_1887_n N_noxref_10_c_2216_n ) capacitor c=0.0229907f \
 //x=21.65 //y=5.155 //x2=27.265 //y2=4.07
cc_1364 ( N_QN_c_1859_n N_noxref_10_c_2216_n ) capacitor c=0.0131995f \
 //x=25.435 //y=4.79 //x2=27.265 //y2=4.07
cc_1365 ( N_QN_c_1842_n N_noxref_10_c_2235_n ) capacitor c=3.10026e-19 \
 //x=20.855 //y=5.155 //x2=18.415 //y2=5.155
cc_1366 ( N_QN_c_1825_n N_noxref_10_c_2212_n ) capacitor c=0.00153442f \
 //x=25.16 //y=2.08 //x2=27.38 //y2=2.08
cc_1367 ( N_QN_c_1823_n N_Q_c_2549_n ) capacitor c=0.176086f //x=25.045 \
 //y=3.33 //x2=28.005 //y2=3.7
cc_1368 ( N_QN_c_1892_p N_Q_c_2549_n ) capacitor c=0.029467f //x=23.425 \
 //y=3.33 //x2=28.005 //y2=3.7
cc_1369 ( QN N_Q_c_2549_n ) capacitor c=0.0206044f //x=23.31 //y=2.22 \
 //x2=28.005 //y2=3.7
cc_1370 ( N_QN_c_1825_n N_Q_c_2549_n ) capacitor c=0.0215974f //x=25.16 \
 //y=2.08 //x2=28.005 //y2=3.7
cc_1371 ( QN N_Q_c_2588_n ) capacitor c=0.00131333f //x=23.31 //y=2.22 \
 //x2=22.685 //y2=3.7
cc_1372 ( N_QN_c_1892_p N_Q_c_2550_n ) capacitor c=0.00720056f //x=23.425 \
 //y=3.33 //x2=22.57 //y2=2.08
cc_1373 ( QN N_Q_c_2550_n ) capacitor c=0.082926f //x=23.31 //y=2.22 \
 //x2=22.57 //y2=2.08
cc_1374 ( N_QN_c_1825_n N_Q_c_2550_n ) capacitor c=9.66956e-19 //x=25.16 \
 //y=2.08 //x2=22.57 //y2=2.08
cc_1375 ( N_QN_c_1936_p N_Q_c_2550_n ) capacitor c=0.0168082f //x=22.53 \
 //y=5.155 //x2=22.57 //y2=2.08
cc_1376 ( N_QN_M49_noxref_g N_Q_c_2556_n ) capacitor c=0.0178794f //x=25.8 \
 //y=6.02 //x2=26.375 //y2=5.155
cc_1377 ( N_QN_c_1848_n N_Q_c_2560_n ) capacitor c=3.10026e-19 //x=23.225 \
 //y=5.155 //x2=25.665 //y2=5.155
cc_1378 ( N_QN_M48_noxref_g N_Q_c_2560_n ) capacitor c=0.0213876f //x=25.36 \
 //y=6.02 //x2=25.665 //y2=5.155
cc_1379 ( N_QN_c_1901_p N_Q_c_2560_n ) capacitor c=0.00429591f //x=25.725 \
 //y=4.79 //x2=25.665 //y2=5.155
cc_1380 ( N_QN_c_1844_n N_Q_M46_noxref_g ) capacitor c=0.0184045f //x=22.445 \
 //y=5.155 //x2=22.31 //y2=6.02
cc_1381 ( N_QN_M46_noxref_d N_Q_M46_noxref_g ) capacitor c=0.0180032f \
 //x=22.385 //y=5.02 //x2=22.31 //y2=6.02
cc_1382 ( N_QN_c_1848_n N_Q_M47_noxref_g ) capacitor c=0.0205426f //x=23.225 \
 //y=5.155 //x2=22.75 //y2=6.02
cc_1383 ( N_QN_M46_noxref_d N_Q_M47_noxref_g ) capacitor c=0.0194246f \
 //x=22.385 //y=5.02 //x2=22.75 //y2=6.02
cc_1384 ( N_QN_M14_noxref_d N_Q_c_2598_n ) capacitor c=0.00217566f //x=22.635 \
 //y=0.915 //x2=22.56 //y2=0.915
cc_1385 ( N_QN_M14_noxref_d N_Q_c_2599_n ) capacitor c=0.0034598f //x=22.635 \
 //y=0.915 //x2=22.56 //y2=1.26
cc_1386 ( N_QN_M14_noxref_d N_Q_c_2600_n ) capacitor c=0.00544291f //x=22.635 \
 //y=0.915 //x2=22.56 //y2=1.57
cc_1387 ( N_QN_M14_noxref_d N_Q_c_2627_n ) capacitor c=0.00241102f //x=22.635 \
 //y=0.915 //x2=22.935 //y2=0.76
cc_1388 ( N_QN_c_1824_n N_Q_c_2628_n ) capacitor c=0.00359704f //x=23.225 \
 //y=1.665 //x2=22.935 //y2=1.415
cc_1389 ( N_QN_M14_noxref_d N_Q_c_2628_n ) capacitor c=0.0140297f //x=22.635 \
 //y=0.915 //x2=22.935 //y2=1.415
cc_1390 ( N_QN_M14_noxref_d N_Q_c_2630_n ) capacitor c=0.00219619f //x=22.635 \
 //y=0.915 //x2=23.09 //y2=0.915
cc_1391 ( N_QN_c_1824_n N_Q_c_2631_n ) capacitor c=0.00457401f //x=23.225 \
 //y=1.665 //x2=23.09 //y2=1.26
cc_1392 ( N_QN_M14_noxref_d N_Q_c_2631_n ) capacitor c=0.00603828f //x=22.635 \
 //y=0.915 //x2=23.09 //y2=1.26
cc_1393 ( QN N_Q_c_2601_n ) capacitor c=0.00877984f //x=23.31 //y=2.22 \
 //x2=22.57 //y2=2.08
cc_1394 ( QN N_Q_c_2603_n ) capacitor c=0.00283672f //x=23.31 //y=2.22 \
 //x2=22.57 //y2=1.915
cc_1395 ( N_QN_M14_noxref_d N_Q_c_2603_n ) capacitor c=0.00661782f //x=22.635 \
 //y=0.915 //x2=22.57 //y2=1.915
cc_1396 ( QN N_Q_c_2604_n ) capacitor c=0.013693f //x=23.31 //y=2.22 \
 //x2=22.57 //y2=4.7
cc_1397 ( N_QN_c_1848_n N_Q_c_2604_n ) capacitor c=0.00201851f //x=23.225 \
 //y=5.155 //x2=22.57 //y2=4.7
cc_1398 ( N_QN_c_1936_p N_Q_c_2604_n ) capacitor c=0.00475729f //x=22.53 \
 //y=5.155 //x2=22.57 //y2=4.7
cc_1399 ( N_QN_M49_noxref_g N_Q_M48_noxref_d ) capacitor c=0.0180032f //x=25.8 \
 //y=6.02 //x2=25.435 //y2=5.02
cc_1400 ( N_QN_M14_noxref_d N_noxref_21_M12_noxref_s ) capacitor c=0.00309936f \
 //x=22.635 //y=0.915 //x2=19.695 //y2=0.375
cc_1401 ( N_QN_c_1824_n N_noxref_22_c_3235_n ) capacitor c=0.00461497f \
 //x=23.225 //y=1.665 //x2=23.225 //y2=0.54
cc_1402 ( N_QN_M14_noxref_d N_noxref_22_c_3235_n ) capacitor c=0.0116817f \
 //x=22.635 //y=0.915 //x2=23.225 //y2=0.54
cc_1403 ( N_QN_c_1894_p N_noxref_22_c_3258_n ) capacitor c=0.0200405f \
 //x=22.91 //y=1.665 //x2=22.34 //y2=0.995
cc_1404 ( N_QN_M14_noxref_d N_noxref_22_M13_noxref_d ) capacitor c=5.27807e-19 \
 //x=22.635 //y=0.915 //x2=21.1 //y2=0.91
cc_1405 ( N_QN_c_1824_n N_noxref_22_M14_noxref_s ) capacitor c=0.0201579f \
 //x=23.225 //y=1.665 //x2=22.205 //y2=0.375
cc_1406 ( N_QN_M14_noxref_d N_noxref_22_M14_noxref_s ) capacitor c=0.0426368f \
 //x=22.635 //y=0.915 //x2=22.205 //y2=0.375
cc_1407 ( N_QN_c_1824_n N_noxref_23_c_3297_n ) capacitor c=3.84569e-19 \
 //x=23.225 //y=1.665 //x2=24.64 //y2=1.505
cc_1408 ( N_QN_c_1830_n N_noxref_23_c_3297_n ) capacitor c=0.0034165f \
 //x=24.86 //y=1.915 //x2=24.64 //y2=1.505
cc_1409 ( N_QN_c_1825_n N_noxref_23_c_3283_n ) capacitor c=0.0122624f \
 //x=25.16 //y=2.08 //x2=25.525 //y2=1.59
cc_1410 ( N_QN_c_1829_n N_noxref_23_c_3283_n ) capacitor c=0.00703864f \
 //x=24.86 //y=1.53 //x2=25.525 //y2=1.59
cc_1411 ( N_QN_c_1830_n N_noxref_23_c_3283_n ) capacitor c=0.0215834f \
 //x=24.86 //y=1.915 //x2=25.525 //y2=1.59
cc_1412 ( N_QN_c_1832_n N_noxref_23_c_3283_n ) capacitor c=0.00708583f \
 //x=25.235 //y=1.375 //x2=25.525 //y2=1.59
cc_1413 ( N_QN_c_1835_n N_noxref_23_c_3283_n ) capacitor c=0.00698822f \
 //x=25.39 //y=1.22 //x2=25.525 //y2=1.59
cc_1414 ( N_QN_c_1826_n N_noxref_23_M15_noxref_s ) capacitor c=0.0327271f \
 //x=24.86 //y=0.875 //x2=24.505 //y2=0.375
cc_1415 ( N_QN_c_1829_n N_noxref_23_M15_noxref_s ) capacitor c=7.99997e-19 \
 //x=24.86 //y=1.53 //x2=24.505 //y2=0.375
cc_1416 ( N_QN_c_1830_n N_noxref_23_M15_noxref_s ) capacitor c=0.00122123f \
 //x=24.86 //y=1.915 //x2=24.505 //y2=0.375
cc_1417 ( N_QN_c_1833_n N_noxref_23_M15_noxref_s ) capacitor c=0.0121427f \
 //x=25.39 //y=0.875 //x2=24.505 //y2=0.375
cc_1418 ( N_QN_M14_noxref_d N_noxref_23_M15_noxref_s ) capacitor c=2.55333e-19 \
 //x=22.635 //y=0.915 //x2=24.505 //y2=0.375
cc_1419 ( N_SN_c_1991_n N_noxref_10_c_2214_n ) capacitor c=0.0190126f \
 //x=11.84 //y=2.08 //x2=12.835 //y2=4.07
cc_1420 ( N_SN_c_1980_n N_noxref_10_c_2215_n ) capacitor c=0.00948333f \
 //x=26.155 //y=2.59 //x2=18.385 //y2=4.07
cc_1421 ( N_SN_c_1991_n N_noxref_10_c_2278_n ) capacitor c=0.00128547f \
 //x=11.84 //y=2.08 //x2=13.065 //y2=4.07
cc_1422 ( N_SN_c_1980_n N_noxref_10_c_2216_n ) capacitor c=0.0565371f \
 //x=26.155 //y=2.59 //x2=27.265 //y2=4.07
cc_1423 ( N_SN_c_1992_n N_noxref_10_c_2216_n ) capacitor c=0.0242403f \
 //x=26.27 //y=2.08 //x2=27.265 //y2=4.07
cc_1424 ( N_SN_c_2093_p N_noxref_10_c_2216_n ) capacitor c=0.0067704f \
 //x=26.605 //y=4.79 //x2=27.265 //y2=4.07
cc_1425 ( N_SN_c_2085_n N_noxref_10_c_2216_n ) capacitor c=0.00230259f \
 //x=26.27 //y=4.7 //x2=27.265 //y2=4.07
cc_1426 ( N_SN_c_1980_n N_noxref_10_c_2223_n ) capacitor c=3.16222e-19 \
 //x=26.155 //y=2.59 //x2=18.615 //y2=4.07
cc_1427 ( N_SN_c_1980_n N_noxref_10_c_2210_n ) capacitor c=0.0238423f \
 //x=26.155 //y=2.59 //x2=12.95 //y2=2.08
cc_1428 ( N_SN_c_1990_n N_noxref_10_c_2210_n ) capacitor c=0.00128547f \
 //x=11.955 //y=2.59 //x2=12.95 //y2=2.08
cc_1429 ( N_SN_c_1991_n N_noxref_10_c_2210_n ) capacitor c=0.0452955f \
 //x=11.84 //y=2.08 //x2=12.95 //y2=2.08
cc_1430 ( N_SN_c_2022_n N_noxref_10_c_2210_n ) capacitor c=0.0023343f \
 //x=11.93 //y=1.915 //x2=12.95 //y2=2.08
cc_1431 ( N_SN_c_2024_n N_noxref_10_c_2210_n ) capacitor c=0.00142741f \
 //x=11.84 //y=4.7 //x2=12.95 //y2=2.08
cc_1432 ( N_SN_c_1980_n N_noxref_10_c_2450_n ) capacitor c=0.0115788f \
 //x=26.155 //y=2.59 //x2=18.1 //y2=1.665
cc_1433 ( N_SN_c_1980_n N_noxref_10_c_2239_n ) capacitor c=0.024834f \
 //x=26.155 //y=2.59 //x2=18.5 //y2=4.07
cc_1434 ( N_SN_c_1980_n N_noxref_10_c_2212_n ) capacitor c=0.00526349f \
 //x=26.155 //y=2.59 //x2=27.38 //y2=2.08
cc_1435 ( N_SN_c_1992_n N_noxref_10_c_2212_n ) capacitor c=0.0511494f \
 //x=26.27 //y=2.08 //x2=27.38 //y2=2.08
cc_1436 ( N_SN_c_2083_n N_noxref_10_c_2212_n ) capacitor c=0.0023343f \
 //x=26.36 //y=1.915 //x2=27.38 //y2=2.08
cc_1437 ( N_SN_c_2085_n N_noxref_10_c_2212_n ) capacitor c=0.00142741f \
 //x=26.27 //y=4.7 //x2=27.38 //y2=2.08
cc_1438 ( N_SN_M32_noxref_g N_noxref_10_M34_noxref_g ) capacitor c=0.0101598f \
 //x=11.81 //y=6.02 //x2=12.69 //y2=6.02
cc_1439 ( N_SN_M33_noxref_g N_noxref_10_M34_noxref_g ) capacitor c=0.0602553f \
 //x=12.25 //y=6.02 //x2=12.69 //y2=6.02
cc_1440 ( N_SN_M33_noxref_g N_noxref_10_M35_noxref_g ) capacitor c=0.0101598f \
 //x=12.25 //y=6.02 //x2=13.13 //y2=6.02
cc_1441 ( N_SN_M50_noxref_g N_noxref_10_M52_noxref_g ) capacitor c=0.0101598f \
 //x=26.24 //y=6.02 //x2=27.12 //y2=6.02
cc_1442 ( N_SN_M51_noxref_g N_noxref_10_M52_noxref_g ) capacitor c=0.0602553f \
 //x=26.68 //y=6.02 //x2=27.12 //y2=6.02
cc_1443 ( N_SN_M51_noxref_g N_noxref_10_M53_noxref_g ) capacitor c=0.0101598f \
 //x=26.68 //y=6.02 //x2=27.56 //y2=6.02
cc_1444 ( N_SN_c_2019_n N_noxref_10_c_2291_n ) capacitor c=0.00456962f \
 //x=11.93 //y=0.91 //x2=12.94 //y2=0.915
cc_1445 ( N_SN_c_2020_n N_noxref_10_c_2292_n ) capacitor c=0.00438372f \
 //x=11.93 //y=1.22 //x2=12.94 //y2=1.26
cc_1446 ( N_SN_c_2021_n N_noxref_10_c_2293_n ) capacitor c=0.00438372f \
 //x=11.93 //y=1.45 //x2=12.94 //y2=1.57
cc_1447 ( N_SN_c_2080_n N_noxref_10_c_2465_n ) capacitor c=0.00456962f \
 //x=26.36 //y=0.91 //x2=27.37 //y2=0.915
cc_1448 ( N_SN_c_2081_n N_noxref_10_c_2466_n ) capacitor c=0.00438372f \
 //x=26.36 //y=1.22 //x2=27.37 //y2=1.26
cc_1449 ( N_SN_c_2082_n N_noxref_10_c_2467_n ) capacitor c=0.00438372f \
 //x=26.36 //y=1.45 //x2=27.37 //y2=1.57
cc_1450 ( N_SN_c_1980_n N_noxref_10_c_2300_n ) capacitor c=0.00232725f \
 //x=26.155 //y=2.59 //x2=12.95 //y2=2.08
cc_1451 ( N_SN_c_1991_n N_noxref_10_c_2300_n ) capacitor c=0.00228632f \
 //x=11.84 //y=2.08 //x2=12.95 //y2=2.08
cc_1452 ( N_SN_c_2022_n N_noxref_10_c_2300_n ) capacitor c=0.00933826f \
 //x=11.93 //y=1.915 //x2=12.95 //y2=2.08
cc_1453 ( N_SN_c_2022_n N_noxref_10_c_2301_n ) capacitor c=0.00438372f \
 //x=11.93 //y=1.915 //x2=12.95 //y2=1.915
cc_1454 ( N_SN_c_1991_n N_noxref_10_c_2303_n ) capacitor c=0.00219458f \
 //x=11.84 //y=2.08 //x2=12.95 //y2=4.7
cc_1455 ( N_SN_c_2039_n N_noxref_10_c_2303_n ) capacitor c=0.0611812f \
 //x=12.175 //y=4.79 //x2=12.95 //y2=4.7
cc_1456 ( N_SN_c_2024_n N_noxref_10_c_2303_n ) capacitor c=0.00487508f \
 //x=11.84 //y=4.7 //x2=12.95 //y2=4.7
cc_1457 ( N_SN_c_1992_n N_noxref_10_c_2475_n ) capacitor c=0.00228632f \
 //x=26.27 //y=2.08 //x2=27.38 //y2=2.08
cc_1458 ( N_SN_c_2083_n N_noxref_10_c_2475_n ) capacitor c=0.00933826f \
 //x=26.36 //y=1.915 //x2=27.38 //y2=2.08
cc_1459 ( N_SN_c_2083_n N_noxref_10_c_2477_n ) capacitor c=0.00438372f \
 //x=26.36 //y=1.915 //x2=27.38 //y2=1.915
cc_1460 ( N_SN_c_1992_n N_noxref_10_c_2478_n ) capacitor c=0.00219458f \
 //x=26.27 //y=2.08 //x2=27.38 //y2=4.7
cc_1461 ( N_SN_c_2093_p N_noxref_10_c_2478_n ) capacitor c=0.0611812f \
 //x=26.605 //y=4.79 //x2=27.38 //y2=4.7
cc_1462 ( N_SN_c_2085_n N_noxref_10_c_2478_n ) capacitor c=0.00487508f \
 //x=26.27 //y=4.7 //x2=27.38 //y2=4.7
cc_1463 ( N_SN_c_1980_n N_Q_c_2549_n ) capacitor c=0.0534079f //x=26.155 \
 //y=2.59 //x2=28.005 //y2=3.7
cc_1464 ( N_SN_c_1992_n N_Q_c_2549_n ) capacitor c=0.0229885f //x=26.27 \
 //y=2.08 //x2=28.005 //y2=3.7
cc_1465 ( N_SN_c_1980_n N_Q_c_2588_n ) capacitor c=0.00777466f //x=26.155 \
 //y=2.59 //x2=22.685 //y2=3.7
cc_1466 ( N_SN_c_1992_n Q ) capacitor c=0.00376573f //x=26.27 //y=2.08 \
 //x2=28.12 //y2=2.22
cc_1467 ( N_SN_c_1980_n N_Q_c_2550_n ) capacitor c=0.025454f //x=26.155 \
 //y=2.59 //x2=22.57 //y2=2.08
cc_1468 ( N_SN_c_1992_n N_Q_c_2556_n ) capacitor c=0.0148665f //x=26.27 \
 //y=2.08 //x2=26.375 //y2=5.155
cc_1469 ( N_SN_M50_noxref_g N_Q_c_2556_n ) capacitor c=0.0166659f //x=26.24 \
 //y=6.02 //x2=26.375 //y2=5.155
cc_1470 ( N_SN_c_2085_n N_Q_c_2556_n ) capacitor c=0.00322396f //x=26.27 \
 //y=4.7 //x2=26.375 //y2=5.155
cc_1471 ( N_SN_M51_noxref_g N_Q_c_2562_n ) capacitor c=0.0184045f //x=26.68 \
 //y=6.02 //x2=27.255 //y2=5.155
cc_1472 ( N_SN_c_2093_p N_Q_c_2649_n ) capacitor c=0.00427862f //x=26.605 \
 //y=4.79 //x2=26.46 //y2=5.155
cc_1473 ( N_SN_c_1980_n N_Q_c_2601_n ) capacitor c=0.00232725f //x=26.155 \
 //y=2.59 //x2=22.57 //y2=2.08
cc_1474 ( N_SN_M50_noxref_g N_Q_M50_noxref_d ) capacitor c=0.0180032f \
 //x=26.24 //y=6.02 //x2=26.315 //y2=5.02
cc_1475 ( N_SN_M51_noxref_g N_Q_M50_noxref_d ) capacitor c=0.0180032f \
 //x=26.68 //y=6.02 //x2=26.315 //y2=5.02
cc_1476 ( N_SN_c_2014_n N_noxref_17_c_2974_n ) capacitor c=0.0167228f \
 //x=11.405 //y=0.91 //x2=12.065 //y2=0.54
cc_1477 ( N_SN_c_2019_n N_noxref_17_c_2974_n ) capacitor c=0.00534519f \
 //x=11.93 //y=0.91 //x2=12.065 //y2=0.54
cc_1478 ( N_SN_c_1980_n N_noxref_17_c_2997_n ) capacitor c=0.0029635f \
 //x=26.155 //y=2.59 //x2=12.065 //y2=1.59
cc_1479 ( N_SN_c_1990_n N_noxref_17_c_2997_n ) capacitor c=0.00236045f \
 //x=11.955 //y=2.59 //x2=12.065 //y2=1.59
cc_1480 ( N_SN_c_1991_n N_noxref_17_c_2997_n ) capacitor c=0.0120444f \
 //x=11.84 //y=2.08 //x2=12.065 //y2=1.59
cc_1481 ( N_SN_c_2017_n N_noxref_17_c_2997_n ) capacitor c=0.0153476f \
 //x=11.405 //y=1.22 //x2=12.065 //y2=1.59
cc_1482 ( N_SN_c_2022_n N_noxref_17_c_2997_n ) capacitor c=0.0219169f \
 //x=11.93 //y=1.915 //x2=12.065 //y2=1.59
cc_1483 ( N_SN_c_1980_n N_noxref_17_M6_noxref_s ) capacitor c=0.0041843f \
 //x=26.155 //y=2.59 //x2=10.075 //y2=0.375
cc_1484 ( N_SN_c_2014_n N_noxref_17_M6_noxref_s ) capacitor c=0.00798959f \
 //x=11.405 //y=0.91 //x2=10.075 //y2=0.375
cc_1485 ( N_SN_c_2021_n N_noxref_17_M6_noxref_s ) capacitor c=0.00212176f \
 //x=11.93 //y=1.45 //x2=10.075 //y2=0.375
cc_1486 ( N_SN_c_2022_n N_noxref_17_M6_noxref_s ) capacitor c=0.00298115f \
 //x=11.93 //y=1.915 //x2=10.075 //y2=0.375
cc_1487 ( N_SN_c_1980_n N_noxref_18_c_3021_n ) capacitor c=0.00494691f \
 //x=26.155 //y=2.59 //x2=12.635 //y2=0.995
cc_1488 ( N_SN_c_2157_p N_noxref_18_c_3021_n ) capacitor c=2.14837e-19 \
 //x=11.775 //y=0.755 //x2=12.635 //y2=0.995
cc_1489 ( N_SN_c_2019_n N_noxref_18_c_3021_n ) capacitor c=0.00123426f \
 //x=11.93 //y=0.91 //x2=12.635 //y2=0.995
cc_1490 ( N_SN_c_2020_n N_noxref_18_c_3021_n ) capacitor c=0.0129288f \
 //x=11.93 //y=1.22 //x2=12.635 //y2=0.995
cc_1491 ( N_SN_c_2021_n N_noxref_18_c_3021_n ) capacitor c=0.00142359f \
 //x=11.93 //y=1.45 //x2=12.635 //y2=0.995
cc_1492 ( N_SN_c_1980_n N_noxref_18_c_3027_n ) capacitor c=8.29806e-19 \
 //x=26.155 //y=2.59 //x2=13.605 //y2=0.54
cc_1493 ( N_SN_c_2014_n N_noxref_18_M7_noxref_d ) capacitor c=0.00223875f \
 //x=11.405 //y=0.91 //x2=11.48 //y2=0.91
cc_1494 ( N_SN_c_2017_n N_noxref_18_M7_noxref_d ) capacitor c=0.00262485f \
 //x=11.405 //y=1.22 //x2=11.48 //y2=0.91
cc_1495 ( N_SN_c_2157_p N_noxref_18_M7_noxref_d ) capacitor c=0.00220746f \
 //x=11.775 //y=0.755 //x2=11.48 //y2=0.91
cc_1496 ( N_SN_c_2165_p N_noxref_18_M7_noxref_d ) capacitor c=0.00194798f \
 //x=11.775 //y=1.375 //x2=11.48 //y2=0.91
cc_1497 ( N_SN_c_2019_n N_noxref_18_M7_noxref_d ) capacitor c=0.00198465f \
 //x=11.93 //y=0.91 //x2=11.48 //y2=0.91
cc_1498 ( N_SN_c_2020_n N_noxref_18_M7_noxref_d ) capacitor c=0.00128384f \
 //x=11.93 //y=1.22 //x2=11.48 //y2=0.91
cc_1499 ( N_SN_c_1980_n N_noxref_18_M8_noxref_s ) capacitor c=0.00448771f \
 //x=26.155 //y=2.59 //x2=12.585 //y2=0.375
cc_1500 ( N_SN_c_2019_n N_noxref_18_M8_noxref_s ) capacitor c=7.21316e-19 \
 //x=11.93 //y=0.91 //x2=12.585 //y2=0.375
cc_1501 ( N_SN_c_2020_n N_noxref_18_M8_noxref_s ) capacitor c=0.00348171f \
 //x=11.93 //y=1.22 //x2=12.585 //y2=0.375
cc_1502 ( N_SN_c_1980_n N_noxref_19_c_3091_n ) capacitor c=0.00448771f \
 //x=26.155 //y=2.59 //x2=15.02 //y2=1.505
cc_1503 ( N_SN_c_1980_n N_noxref_19_c_3075_n ) capacitor c=0.0163649f \
 //x=26.155 //y=2.59 //x2=15.905 //y2=1.59
cc_1504 ( N_SN_c_1980_n N_noxref_19_c_3105_n ) capacitor c=0.0144126f \
 //x=26.155 //y=2.59 //x2=16.875 //y2=1.59
cc_1505 ( N_SN_c_1980_n N_noxref_19_M9_noxref_s ) capacitor c=0.00867201f \
 //x=26.155 //y=2.59 //x2=14.885 //y2=0.375
cc_1506 ( N_SN_c_1980_n N_noxref_20_c_3125_n ) capacitor c=0.00494691f \
 //x=26.155 //y=2.59 //x2=17.445 //y2=0.995
cc_1507 ( N_SN_c_1980_n N_noxref_20_c_3131_n ) capacitor c=8.29806e-19 \
 //x=26.155 //y=2.59 //x2=18.415 //y2=0.54
cc_1508 ( N_SN_c_1980_n N_noxref_20_M11_noxref_s ) capacitor c=0.00448771f \
 //x=26.155 //y=2.59 //x2=17.395 //y2=0.375
cc_1509 ( N_SN_c_1980_n N_noxref_21_c_3195_n ) capacitor c=0.00448771f \
 //x=26.155 //y=2.59 //x2=19.83 //y2=1.505
cc_1510 ( N_SN_c_1980_n N_noxref_21_c_3179_n ) capacitor c=0.0163649f \
 //x=26.155 //y=2.59 //x2=20.715 //y2=1.59
cc_1511 ( N_SN_c_1980_n N_noxref_21_c_3207_n ) capacitor c=0.0144126f \
 //x=26.155 //y=2.59 //x2=21.685 //y2=1.59
cc_1512 ( N_SN_c_1980_n N_noxref_21_M12_noxref_s ) capacitor c=0.00867201f \
 //x=26.155 //y=2.59 //x2=19.695 //y2=0.375
cc_1513 ( N_SN_c_1980_n N_noxref_22_c_3229_n ) capacitor c=0.00494691f \
 //x=26.155 //y=2.59 //x2=22.255 //y2=0.995
cc_1514 ( N_SN_c_1980_n N_noxref_22_c_3235_n ) capacitor c=8.29806e-19 \
 //x=26.155 //y=2.59 //x2=23.225 //y2=0.54
cc_1515 ( N_SN_c_1980_n N_noxref_22_M14_noxref_s ) capacitor c=0.00448771f \
 //x=26.155 //y=2.59 //x2=22.205 //y2=0.375
cc_1516 ( N_SN_c_1980_n N_noxref_23_c_3297_n ) capacitor c=0.00448771f \
 //x=26.155 //y=2.59 //x2=24.64 //y2=1.505
cc_1517 ( N_SN_c_1980_n N_noxref_23_c_3283_n ) capacitor c=0.0163649f \
 //x=26.155 //y=2.59 //x2=25.525 //y2=1.59
cc_1518 ( N_SN_c_2075_n N_noxref_23_c_3290_n ) capacitor c=0.0167228f \
 //x=25.835 //y=0.91 //x2=26.495 //y2=0.54
cc_1519 ( N_SN_c_2080_n N_noxref_23_c_3290_n ) capacitor c=0.00534519f \
 //x=26.36 //y=0.91 //x2=26.495 //y2=0.54
cc_1520 ( N_SN_c_1980_n N_noxref_23_c_3313_n ) capacitor c=0.0125159f \
 //x=26.155 //y=2.59 //x2=26.495 //y2=1.59
cc_1521 ( N_SN_c_1992_n N_noxref_23_c_3313_n ) capacitor c=0.0123163f \
 //x=26.27 //y=2.08 //x2=26.495 //y2=1.59
cc_1522 ( N_SN_c_2078_n N_noxref_23_c_3313_n ) capacitor c=0.0153476f \
 //x=25.835 //y=1.22 //x2=26.495 //y2=1.59
cc_1523 ( N_SN_c_2083_n N_noxref_23_c_3313_n ) capacitor c=0.0221623f \
 //x=26.36 //y=1.915 //x2=26.495 //y2=1.59
cc_1524 ( N_SN_c_1980_n N_noxref_23_M15_noxref_s ) capacitor c=0.00448771f \
 //x=26.155 //y=2.59 //x2=24.505 //y2=0.375
cc_1525 ( N_SN_c_2075_n N_noxref_23_M15_noxref_s ) capacitor c=0.00798959f \
 //x=25.835 //y=0.91 //x2=24.505 //y2=0.375
cc_1526 ( N_SN_c_2082_n N_noxref_23_M15_noxref_s ) capacitor c=0.00212176f \
 //x=26.36 //y=1.45 //x2=24.505 //y2=0.375
cc_1527 ( N_SN_c_2083_n N_noxref_23_M15_noxref_s ) capacitor c=0.00298115f \
 //x=26.36 //y=1.915 //x2=24.505 //y2=0.375
cc_1528 ( N_SN_c_2197_p N_noxref_24_c_3333_n ) capacitor c=2.14837e-19 \
 //x=26.205 //y=0.755 //x2=27.065 //y2=0.995
cc_1529 ( N_SN_c_2080_n N_noxref_24_c_3333_n ) capacitor c=0.00123426f \
 //x=26.36 //y=0.91 //x2=27.065 //y2=0.995
cc_1530 ( N_SN_c_2081_n N_noxref_24_c_3333_n ) capacitor c=0.0129288f \
 //x=26.36 //y=1.22 //x2=27.065 //y2=0.995
cc_1531 ( N_SN_c_2082_n N_noxref_24_c_3333_n ) capacitor c=0.00142359f \
 //x=26.36 //y=1.45 //x2=27.065 //y2=0.995
cc_1532 ( N_SN_c_2075_n N_noxref_24_M16_noxref_d ) capacitor c=0.00223875f \
 //x=25.835 //y=0.91 //x2=25.91 //y2=0.91
cc_1533 ( N_SN_c_2078_n N_noxref_24_M16_noxref_d ) capacitor c=0.00262485f \
 //x=25.835 //y=1.22 //x2=25.91 //y2=0.91
cc_1534 ( N_SN_c_2197_p N_noxref_24_M16_noxref_d ) capacitor c=0.00220746f \
 //x=26.205 //y=0.755 //x2=25.91 //y2=0.91
cc_1535 ( N_SN_c_2204_p N_noxref_24_M16_noxref_d ) capacitor c=0.00194798f \
 //x=26.205 //y=1.375 //x2=25.91 //y2=0.91
cc_1536 ( N_SN_c_2080_n N_noxref_24_M16_noxref_d ) capacitor c=0.00198465f \
 //x=26.36 //y=0.91 //x2=25.91 //y2=0.91
cc_1537 ( N_SN_c_2081_n N_noxref_24_M16_noxref_d ) capacitor c=0.00128384f \
 //x=26.36 //y=1.22 //x2=25.91 //y2=0.91
cc_1538 ( N_SN_c_2080_n N_noxref_24_M17_noxref_s ) capacitor c=7.21316e-19 \
 //x=26.36 //y=0.91 //x2=27.015 //y2=0.375
cc_1539 ( N_SN_c_2081_n N_noxref_24_M17_noxref_s ) capacitor c=0.00348171f \
 //x=26.36 //y=1.22 //x2=27.015 //y2=0.375
cc_1540 ( N_noxref_10_c_2216_n N_Q_c_2549_n ) capacitor c=0.433554f //x=27.265 \
 //y=4.07 //x2=28.005 //y2=3.7
cc_1541 ( N_noxref_10_c_2212_n N_Q_c_2549_n ) capacitor c=0.027223f //x=27.38 \
 //y=2.08 //x2=28.005 //y2=3.7
cc_1542 ( N_noxref_10_c_2478_n N_Q_c_2549_n ) capacitor c=0.0018324f //x=27.38 \
 //y=4.7 //x2=28.005 //y2=3.7
cc_1543 ( N_noxref_10_c_2216_n N_Q_c_2588_n ) capacitor c=0.0292842f \
 //x=27.265 //y=4.07 //x2=22.685 //y2=3.7
cc_1544 ( N_noxref_10_c_2216_n Q ) capacitor c=0.00642908f //x=27.265 //y=4.07 \
 //x2=28.12 //y2=2.22
cc_1545 ( N_noxref_10_c_2212_n Q ) capacitor c=0.0880964f //x=27.38 //y=2.08 \
 //x2=28.12 //y2=2.22
cc_1546 ( N_noxref_10_c_2475_n Q ) capacitor c=0.00877984f //x=27.38 //y=2.08 \
 //x2=28.12 //y2=2.22
cc_1547 ( N_noxref_10_c_2477_n Q ) capacitor c=0.00283672f //x=27.38 //y=1.915 \
 //x2=28.12 //y2=2.22
cc_1548 ( N_noxref_10_c_2478_n Q ) capacitor c=0.013844f //x=27.38 //y=4.7 \
 //x2=28.12 //y2=2.22
cc_1549 ( N_noxref_10_c_2216_n N_Q_c_2550_n ) capacitor c=0.0237491f \
 //x=27.265 //y=4.07 //x2=22.57 //y2=2.08
cc_1550 ( N_noxref_10_c_2216_n N_Q_c_2556_n ) capacitor c=0.0236892f \
 //x=27.265 //y=4.07 //x2=26.375 //y2=5.155
cc_1551 ( N_noxref_10_c_2216_n N_Q_c_2560_n ) capacitor c=0.0173f //x=27.265 \
 //y=4.07 //x2=25.665 //y2=5.155
cc_1552 ( N_noxref_10_M52_noxref_g N_Q_c_2562_n ) capacitor c=0.0184045f \
 //x=27.12 //y=6.02 //x2=27.255 //y2=5.155
cc_1553 ( N_noxref_10_c_2216_n N_Q_c_2566_n ) capacitor c=0.00181724f \
 //x=27.265 //y=4.07 //x2=28.035 //y2=5.155
cc_1554 ( N_noxref_10_M53_noxref_g N_Q_c_2566_n ) capacitor c=0.0211056f \
 //x=27.56 //y=6.02 //x2=28.035 //y2=5.155
cc_1555 ( N_noxref_10_c_2478_n N_Q_c_2566_n ) capacitor c=0.00201851f \
 //x=27.38 //y=4.7 //x2=28.035 //y2=5.155
cc_1556 ( N_noxref_10_c_2497_p N_Q_c_2551_n ) capacitor c=0.00359704f \
 //x=27.745 //y=1.415 //x2=28.035 //y2=1.665
cc_1557 ( N_noxref_10_c_2498_p N_Q_c_2551_n ) capacitor c=0.00457401f //x=27.9 \
 //y=1.26 //x2=28.035 //y2=1.665
cc_1558 ( N_noxref_10_c_2216_n N_Q_c_2671_n ) capacitor c=7.87932e-19 \
 //x=27.265 //y=4.07 //x2=27.34 //y2=5.155
cc_1559 ( N_noxref_10_c_2212_n N_Q_c_2671_n ) capacitor c=0.0169174f //x=27.38 \
 //y=2.08 //x2=27.34 //y2=5.155
cc_1560 ( N_noxref_10_c_2478_n N_Q_c_2671_n ) capacitor c=0.0047572f //x=27.38 \
 //y=4.7 //x2=27.34 //y2=5.155
cc_1561 ( N_noxref_10_c_2216_n N_Q_c_2604_n ) capacitor c=0.00775263f \
 //x=27.265 //y=4.07 //x2=22.57 //y2=4.7
cc_1562 ( N_noxref_10_c_2465_n N_Q_M17_noxref_d ) capacitor c=0.00217566f \
 //x=27.37 //y=0.915 //x2=27.445 //y2=0.915
cc_1563 ( N_noxref_10_c_2466_n N_Q_M17_noxref_d ) capacitor c=0.0034598f \
 //x=27.37 //y=1.26 //x2=27.445 //y2=0.915
cc_1564 ( N_noxref_10_c_2467_n N_Q_M17_noxref_d ) capacitor c=0.00544291f \
 //x=27.37 //y=1.57 //x2=27.445 //y2=0.915
cc_1565 ( N_noxref_10_c_2506_p N_Q_M17_noxref_d ) capacitor c=0.00241102f \
 //x=27.745 //y=0.76 //x2=27.445 //y2=0.915
cc_1566 ( N_noxref_10_c_2497_p N_Q_M17_noxref_d ) capacitor c=0.0140297f \
 //x=27.745 //y=1.415 //x2=27.445 //y2=0.915
cc_1567 ( N_noxref_10_c_2508_p N_Q_M17_noxref_d ) capacitor c=0.00219619f \
 //x=27.9 //y=0.915 //x2=27.445 //y2=0.915
cc_1568 ( N_noxref_10_c_2498_p N_Q_M17_noxref_d ) capacitor c=0.00603828f \
 //x=27.9 //y=1.26 //x2=27.445 //y2=0.915
cc_1569 ( N_noxref_10_c_2477_n N_Q_M17_noxref_d ) capacitor c=0.00661782f \
 //x=27.38 //y=1.915 //x2=27.445 //y2=0.915
cc_1570 ( N_noxref_10_M52_noxref_g N_Q_M52_noxref_d ) capacitor c=0.0180032f \
 //x=27.12 //y=6.02 //x2=27.195 //y2=5.02
cc_1571 ( N_noxref_10_M53_noxref_g N_Q_M52_noxref_d ) capacitor c=0.0194246f \
 //x=27.56 //y=6.02 //x2=27.195 //y2=5.02
cc_1572 ( N_noxref_10_c_2209_n N_noxref_16_c_2919_n ) capacitor c=0.00207747f \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_1573 ( N_noxref_10_c_2330_n N_noxref_16_c_2919_n ) capacitor c=0.0194423f \
 //x=8.13 //y=0.915 //x2=8.795 //y2=0.54
cc_1574 ( N_noxref_10_c_2373_n N_noxref_16_c_2919_n ) capacitor c=0.00656458f \
 //x=8.66 //y=0.915 //x2=8.795 //y2=0.54
cc_1575 ( N_noxref_10_c_2275_n N_noxref_16_c_2919_n ) capacitor c=2.20712e-19 \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_1576 ( N_noxref_10_c_2331_n N_noxref_16_c_2945_n ) capacitor c=0.00538829f \
 //x=8.13 //y=1.26 //x2=7.91 //y2=0.995
cc_1577 ( N_noxref_10_c_2330_n N_noxref_16_M5_noxref_s ) capacitor \
 c=0.00538829f //x=8.13 //y=0.915 //x2=7.775 //y2=0.375
cc_1578 ( N_noxref_10_c_2332_n N_noxref_16_M5_noxref_s ) capacitor \
 c=0.00538829f //x=8.13 //y=1.57 //x2=7.775 //y2=0.375
cc_1579 ( N_noxref_10_c_2373_n N_noxref_16_M5_noxref_s ) capacitor \
 c=0.0143002f //x=8.66 //y=0.915 //x2=7.775 //y2=0.375
cc_1580 ( N_noxref_10_c_2374_n N_noxref_16_M5_noxref_s ) capacitor \
 c=0.00290153f //x=8.66 //y=1.26 //x2=7.775 //y2=0.375
cc_1581 ( N_noxref_10_c_2210_n N_noxref_18_c_3027_n ) capacitor c=0.0020642f \
 //x=12.95 //y=2.08 //x2=13.605 //y2=0.54
cc_1582 ( N_noxref_10_c_2291_n N_noxref_18_c_3027_n ) capacitor c=0.0194423f \
 //x=12.94 //y=0.915 //x2=13.605 //y2=0.54
cc_1583 ( N_noxref_10_c_2297_n N_noxref_18_c_3027_n ) capacitor c=0.00656458f \
 //x=13.47 //y=0.915 //x2=13.605 //y2=0.54
cc_1584 ( N_noxref_10_c_2300_n N_noxref_18_c_3027_n ) capacitor c=2.20712e-19 \
 //x=12.95 //y=2.08 //x2=13.605 //y2=0.54
cc_1585 ( N_noxref_10_c_2292_n N_noxref_18_c_3038_n ) capacitor c=0.00538829f \
 //x=12.94 //y=1.26 //x2=12.72 //y2=0.995
cc_1586 ( N_noxref_10_c_2291_n N_noxref_18_M8_noxref_s ) capacitor \
 c=0.00538829f //x=12.94 //y=0.915 //x2=12.585 //y2=0.375
cc_1587 ( N_noxref_10_c_2293_n N_noxref_18_M8_noxref_s ) capacitor \
 c=0.00538829f //x=12.94 //y=1.57 //x2=12.585 //y2=0.375
cc_1588 ( N_noxref_10_c_2297_n N_noxref_18_M8_noxref_s ) capacitor \
 c=0.0143002f //x=13.47 //y=0.915 //x2=12.585 //y2=0.375
cc_1589 ( N_noxref_10_c_2298_n N_noxref_18_M8_noxref_s ) capacitor \
 c=0.00290153f //x=13.47 //y=1.26 //x2=12.585 //y2=0.375
cc_1590 ( N_noxref_10_M11_noxref_d N_noxref_19_M9_noxref_s ) capacitor \
 c=0.00309936f //x=17.825 //y=0.915 //x2=14.885 //y2=0.375
cc_1591 ( N_noxref_10_c_2211_n N_noxref_20_c_3131_n ) capacitor c=0.00461497f \
 //x=18.415 //y=1.665 //x2=18.415 //y2=0.54
cc_1592 ( N_noxref_10_M11_noxref_d N_noxref_20_c_3131_n ) capacitor \
 c=0.0116817f //x=17.825 //y=0.915 //x2=18.415 //y2=0.54
cc_1593 ( N_noxref_10_c_2450_n N_noxref_20_c_3156_n ) capacitor c=0.0200405f \
 //x=18.1 //y=1.665 //x2=17.53 //y2=0.995
cc_1594 ( N_noxref_10_M11_noxref_d N_noxref_20_M10_noxref_d ) capacitor \
 c=5.27807e-19 //x=17.825 //y=0.915 //x2=16.29 //y2=0.91
cc_1595 ( N_noxref_10_c_2211_n N_noxref_20_M11_noxref_s ) capacitor \
 c=0.0201579f //x=18.415 //y=1.665 //x2=17.395 //y2=0.375
cc_1596 ( N_noxref_10_M11_noxref_d N_noxref_20_M11_noxref_s ) capacitor \
 c=0.0426368f //x=17.825 //y=0.915 //x2=17.395 //y2=0.375
cc_1597 ( N_noxref_10_c_2211_n N_noxref_21_c_3195_n ) capacitor c=3.84569e-19 \
 //x=18.415 //y=1.665 //x2=19.83 //y2=1.505
cc_1598 ( N_noxref_10_M11_noxref_d N_noxref_21_M12_noxref_s ) capacitor \
 c=2.55333e-19 //x=17.825 //y=0.915 //x2=19.695 //y2=0.375
cc_1599 ( N_noxref_10_c_2212_n N_noxref_24_c_3338_n ) capacitor c=0.00209116f \
 //x=27.38 //y=2.08 //x2=28.035 //y2=0.54
cc_1600 ( N_noxref_10_c_2465_n N_noxref_24_c_3338_n ) capacitor c=0.0194423f \
 //x=27.37 //y=0.915 //x2=28.035 //y2=0.54
cc_1601 ( N_noxref_10_c_2508_p N_noxref_24_c_3338_n ) capacitor c=0.00656458f \
 //x=27.9 //y=0.915 //x2=28.035 //y2=0.54
cc_1602 ( N_noxref_10_c_2475_n N_noxref_24_c_3338_n ) capacitor c=2.20712e-19 \
 //x=27.38 //y=2.08 //x2=28.035 //y2=0.54
cc_1603 ( N_noxref_10_c_2466_n N_noxref_24_c_3361_n ) capacitor c=0.00538829f \
 //x=27.37 //y=1.26 //x2=27.15 //y2=0.995
cc_1604 ( N_noxref_10_c_2465_n N_noxref_24_M17_noxref_s ) capacitor \
 c=0.00538829f //x=27.37 //y=0.915 //x2=27.015 //y2=0.375
cc_1605 ( N_noxref_10_c_2467_n N_noxref_24_M17_noxref_s ) capacitor \
 c=0.00538829f //x=27.37 //y=1.57 //x2=27.015 //y2=0.375
cc_1606 ( N_noxref_10_c_2508_p N_noxref_24_M17_noxref_s ) capacitor \
 c=0.0143002f //x=27.9 //y=0.915 //x2=27.015 //y2=0.375
cc_1607 ( N_noxref_10_c_2498_p N_noxref_24_M17_noxref_s ) capacitor \
 c=0.00290153f //x=27.9 //y=1.26 //x2=27.015 //y2=0.375
cc_1608 ( N_Q_c_2550_n N_noxref_22_c_3235_n ) capacitor c=0.0020642f //x=22.57 \
 //y=2.08 //x2=23.225 //y2=0.54
cc_1609 ( N_Q_c_2598_n N_noxref_22_c_3235_n ) capacitor c=0.0194423f //x=22.56 \
 //y=0.915 //x2=23.225 //y2=0.54
cc_1610 ( N_Q_c_2630_n N_noxref_22_c_3235_n ) capacitor c=0.00656458f \
 //x=23.09 //y=0.915 //x2=23.225 //y2=0.54
cc_1611 ( N_Q_c_2601_n N_noxref_22_c_3235_n ) capacitor c=2.20712e-19 \
 //x=22.57 //y=2.08 //x2=23.225 //y2=0.54
cc_1612 ( N_Q_c_2599_n N_noxref_22_c_3258_n ) capacitor c=0.00538829f \
 //x=22.56 //y=1.26 //x2=22.34 //y2=0.995
cc_1613 ( N_Q_c_2598_n N_noxref_22_M14_noxref_s ) capacitor c=0.00538829f \
 //x=22.56 //y=0.915 //x2=22.205 //y2=0.375
cc_1614 ( N_Q_c_2600_n N_noxref_22_M14_noxref_s ) capacitor c=0.00538829f \
 //x=22.56 //y=1.57 //x2=22.205 //y2=0.375
cc_1615 ( N_Q_c_2630_n N_noxref_22_M14_noxref_s ) capacitor c=0.0143002f \
 //x=23.09 //y=0.915 //x2=22.205 //y2=0.375
cc_1616 ( N_Q_c_2631_n N_noxref_22_M14_noxref_s ) capacitor c=0.00290153f \
 //x=23.09 //y=1.26 //x2=22.205 //y2=0.375
cc_1617 ( N_Q_c_2549_n N_noxref_23_c_3313_n ) capacitor c=0.00104728f \
 //x=28.005 //y=3.7 //x2=26.495 //y2=1.59
cc_1618 ( N_Q_c_2549_n N_noxref_23_M15_noxref_s ) capacitor c=0.00175826f \
 //x=28.005 //y=3.7 //x2=24.505 //y2=0.375
cc_1619 ( N_Q_M17_noxref_d N_noxref_23_M15_noxref_s ) capacitor c=0.00309936f \
 //x=27.445 //y=0.915 //x2=24.505 //y2=0.375
cc_1620 ( N_Q_c_2549_n N_noxref_24_c_3333_n ) capacitor c=0.00250466f \
 //x=28.005 //y=3.7 //x2=27.065 //y2=0.995
cc_1621 ( N_Q_c_2549_n N_noxref_24_c_3338_n ) capacitor c=3.47229e-19 \
 //x=28.005 //y=3.7 //x2=28.035 //y2=0.54
cc_1622 ( N_Q_c_2551_n N_noxref_24_c_3338_n ) capacitor c=0.00467233f \
 //x=28.035 //y=1.665 //x2=28.035 //y2=0.54
cc_1623 ( N_Q_M17_noxref_d N_noxref_24_c_3338_n ) capacitor c=0.0118029f \
 //x=27.445 //y=0.915 //x2=28.035 //y2=0.54
cc_1624 ( N_Q_c_2701_p N_noxref_24_c_3361_n ) capacitor c=0.0200405f //x=27.72 \
 //y=1.665 //x2=27.15 //y2=0.995
cc_1625 ( N_Q_M17_noxref_d N_noxref_24_M16_noxref_d ) capacitor c=5.27807e-19 \
 //x=27.445 //y=0.915 //x2=25.91 //y2=0.91
cc_1626 ( N_Q_c_2549_n N_noxref_24_M17_noxref_s ) capacitor c=0.00188576f \
 //x=28.005 //y=3.7 //x2=27.015 //y2=0.375
cc_1627 ( N_Q_c_2551_n N_noxref_24_M17_noxref_s ) capacitor c=0.0209131f \
 //x=28.035 //y=1.665 //x2=27.015 //y2=0.375
cc_1628 ( N_Q_M17_noxref_d N_noxref_24_M17_noxref_s ) capacitor c=0.0426368f \
 //x=27.445 //y=0.915 //x2=27.015 //y2=0.375
cc_1629 ( N_D_c_2711_n N_noxref_13_c_2790_n ) capacitor c=0.0034165f //x=0.81 \
 //y=1.915 //x2=0.59 //y2=1.505
cc_1630 ( N_D_c_2706_n N_noxref_13_c_2762_n ) capacitor c=0.0122915f //x=1.11 \
 //y=2.08 //x2=1.475 //y2=1.59
cc_1631 ( N_D_c_2710_n N_noxref_13_c_2762_n ) capacitor c=0.00703864f //x=0.81 \
 //y=1.53 //x2=1.475 //y2=1.59
cc_1632 ( N_D_c_2711_n N_noxref_13_c_2762_n ) capacitor c=0.0259045f //x=0.81 \
 //y=1.915 //x2=1.475 //y2=1.59
cc_1633 ( N_D_c_2713_n N_noxref_13_c_2762_n ) capacitor c=0.00708583f \
 //x=1.185 //y=1.375 //x2=1.475 //y2=1.59
cc_1634 ( N_D_c_2716_n N_noxref_13_c_2762_n ) capacitor c=0.00698822f //x=1.34 \
 //y=1.22 //x2=1.475 //y2=1.59
cc_1635 ( N_D_c_2707_n N_noxref_13_M0_noxref_s ) capacitor c=0.0327271f \
 //x=0.81 //y=0.875 //x2=0.455 //y2=0.375
cc_1636 ( N_D_c_2710_n N_noxref_13_M0_noxref_s ) capacitor c=7.99997e-19 \
 //x=0.81 //y=1.53 //x2=0.455 //y2=0.375
cc_1637 ( N_D_c_2711_n N_noxref_13_M0_noxref_s ) capacitor c=0.00122123f \
 //x=0.81 //y=1.915 //x2=0.455 //y2=0.375
cc_1638 ( N_D_c_2714_n N_noxref_13_M0_noxref_s ) capacitor c=0.0121427f \
 //x=1.34 //y=0.875 //x2=0.455 //y2=0.375
cc_1639 ( N_noxref_13_c_2769_n N_noxref_14_c_2808_n ) capacitor c=0.0136048f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_1640 ( N_noxref_13_c_2781_n N_noxref_14_c_2808_n ) capacitor c=0.0102333f \
 //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_1641 ( N_noxref_13_M0_noxref_s N_noxref_14_c_2808_n ) capacitor c=0.023344f \
 //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_1642 ( N_noxref_13_M0_noxref_s N_noxref_14_c_2811_n ) capacitor \
 c=0.0180035f //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_1643 ( N_noxref_13_c_2769_n N_noxref_14_M1_noxref_d ) capacitor \
 c=0.0129526f //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_1644 ( N_noxref_13_c_2781_n N_noxref_14_M1_noxref_d ) capacitor \
 c=0.00912489f //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_1645 ( N_noxref_13_M0_noxref_s N_noxref_14_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_1646 ( N_noxref_13_M0_noxref_s N_noxref_14_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_1647 ( N_noxref_14_c_2817_n N_noxref_15_M3_noxref_s ) capacitor \
 c=0.00191848f //x=4.07 //y=0.625 //x2=5.265 //y2=0.375
cc_1648 ( N_noxref_15_c_2868_n N_noxref_16_c_2913_n ) capacitor c=0.0133829f \
 //x=7.255 //y=0.54 //x2=7.825 //y2=0.995
cc_1649 ( N_noxref_15_c_2888_n N_noxref_16_c_2913_n ) capacitor c=0.0101148f \
 //x=7.255 //y=1.59 //x2=7.825 //y2=0.995
cc_1650 ( N_noxref_15_M3_noxref_s N_noxref_16_c_2913_n ) capacitor \
 c=0.0226294f //x=5.265 //y=0.375 //x2=7.825 //y2=0.995
cc_1651 ( N_noxref_15_M3_noxref_s N_noxref_16_c_2916_n ) capacitor \
 c=0.0180035f //x=5.265 //y=0.375 //x2=7.91 //y2=0.625
cc_1652 ( N_noxref_15_c_2868_n N_noxref_16_M4_noxref_d ) capacitor \
 c=0.0128573f //x=7.255 //y=0.54 //x2=6.67 //y2=0.91
cc_1653 ( N_noxref_15_c_2888_n N_noxref_16_M4_noxref_d ) capacitor \
 c=0.00892105f //x=7.255 //y=1.59 //x2=6.67 //y2=0.91
cc_1654 ( N_noxref_15_M3_noxref_s N_noxref_16_M4_noxref_d ) capacitor \
 c=0.0159202f //x=5.265 //y=0.375 //x2=6.67 //y2=0.91
cc_1655 ( N_noxref_15_M3_noxref_s N_noxref_16_M5_noxref_s ) capacitor \
 c=0.0213553f //x=5.265 //y=0.375 //x2=7.775 //y2=0.375
cc_1656 ( N_noxref_16_c_2922_n N_noxref_17_M6_noxref_s ) capacitor \
 c=0.00191848f //x=8.88 //y=0.625 //x2=10.075 //y2=0.375
cc_1657 ( N_noxref_17_c_2974_n N_noxref_18_c_3021_n ) capacitor c=0.013301f \
 //x=12.065 //y=0.54 //x2=12.635 //y2=0.995
cc_1658 ( N_noxref_17_c_2997_n N_noxref_18_c_3021_n ) capacitor c=0.0100026f \
 //x=12.065 //y=1.59 //x2=12.635 //y2=0.995
cc_1659 ( N_noxref_17_M6_noxref_s N_noxref_18_c_3021_n ) capacitor \
 c=0.0224457f //x=10.075 //y=0.375 //x2=12.635 //y2=0.995
cc_1660 ( N_noxref_17_M6_noxref_s N_noxref_18_c_3024_n ) capacitor \
 c=0.0180035f //x=10.075 //y=0.375 //x2=12.72 //y2=0.625
cc_1661 ( N_noxref_17_c_2974_n N_noxref_18_M7_noxref_d ) capacitor \
 c=0.0128591f //x=12.065 //y=0.54 //x2=11.48 //y2=0.91
cc_1662 ( N_noxref_17_c_2997_n N_noxref_18_M7_noxref_d ) capacitor \
 c=0.00891456f //x=12.065 //y=1.59 //x2=11.48 //y2=0.91
cc_1663 ( N_noxref_17_M6_noxref_s N_noxref_18_M7_noxref_d ) capacitor \
 c=0.0159202f //x=10.075 //y=0.375 //x2=11.48 //y2=0.91
cc_1664 ( N_noxref_17_M6_noxref_s N_noxref_18_M8_noxref_s ) capacitor \
 c=0.0213553f //x=10.075 //y=0.375 //x2=12.585 //y2=0.375
cc_1665 ( N_noxref_18_c_3030_n N_noxref_19_M9_noxref_s ) capacitor \
 c=0.00191848f //x=13.69 //y=0.625 //x2=14.885 //y2=0.375
cc_1666 ( N_noxref_19_c_3082_n N_noxref_20_c_3125_n ) capacitor c=0.0133059f \
 //x=16.875 //y=0.54 //x2=17.445 //y2=0.995
cc_1667 ( N_noxref_19_c_3105_n N_noxref_20_c_3125_n ) capacitor c=0.0100097f \
 //x=16.875 //y=1.59 //x2=17.445 //y2=0.995
cc_1668 ( N_noxref_19_M9_noxref_s N_noxref_20_c_3125_n ) capacitor \
 c=0.0224457f //x=14.885 //y=0.375 //x2=17.445 //y2=0.995
cc_1669 ( N_noxref_19_M9_noxref_s N_noxref_20_c_3128_n ) capacitor \
 c=0.0180035f //x=14.885 //y=0.375 //x2=17.53 //y2=0.625
cc_1670 ( N_noxref_19_c_3082_n N_noxref_20_M10_noxref_d ) capacitor \
 c=0.0128027f //x=16.875 //y=0.54 //x2=16.29 //y2=0.91
cc_1671 ( N_noxref_19_c_3105_n N_noxref_20_M10_noxref_d ) capacitor \
 c=0.00879751f //x=16.875 //y=1.59 //x2=16.29 //y2=0.91
cc_1672 ( N_noxref_19_M9_noxref_s N_noxref_20_M10_noxref_d ) capacitor \
 c=0.0159202f //x=14.885 //y=0.375 //x2=16.29 //y2=0.91
cc_1673 ( N_noxref_19_M9_noxref_s N_noxref_20_M11_noxref_s ) capacitor \
 c=0.0213553f //x=14.885 //y=0.375 //x2=17.395 //y2=0.375
cc_1674 ( N_noxref_20_c_3134_n N_noxref_21_M12_noxref_s ) capacitor \
 c=0.00191848f //x=18.5 //y=0.625 //x2=19.695 //y2=0.375
cc_1675 ( N_noxref_21_c_3186_n N_noxref_22_c_3229_n ) capacitor c=0.0133059f \
 //x=21.685 //y=0.54 //x2=22.255 //y2=0.995
cc_1676 ( N_noxref_21_c_3207_n N_noxref_22_c_3229_n ) capacitor c=0.0100097f \
 //x=21.685 //y=1.59 //x2=22.255 //y2=0.995
cc_1677 ( N_noxref_21_M12_noxref_s N_noxref_22_c_3229_n ) capacitor \
 c=0.0224457f //x=19.695 //y=0.375 //x2=22.255 //y2=0.995
cc_1678 ( N_noxref_21_M12_noxref_s N_noxref_22_c_3232_n ) capacitor \
 c=0.0180035f //x=19.695 //y=0.375 //x2=22.34 //y2=0.625
cc_1679 ( N_noxref_21_c_3186_n N_noxref_22_M13_noxref_d ) capacitor \
 c=0.0128027f //x=21.685 //y=0.54 //x2=21.1 //y2=0.91
cc_1680 ( N_noxref_21_c_3207_n N_noxref_22_M13_noxref_d ) capacitor \
 c=0.00879751f //x=21.685 //y=1.59 //x2=21.1 //y2=0.91
cc_1681 ( N_noxref_21_M12_noxref_s N_noxref_22_M13_noxref_d ) capacitor \
 c=0.0159202f //x=19.695 //y=0.375 //x2=21.1 //y2=0.91
cc_1682 ( N_noxref_21_M12_noxref_s N_noxref_22_M14_noxref_s ) capacitor \
 c=0.0213553f //x=19.695 //y=0.375 //x2=22.205 //y2=0.375
cc_1683 ( N_noxref_22_c_3238_n N_noxref_23_M15_noxref_s ) capacitor \
 c=0.00191848f //x=23.31 //y=0.625 //x2=24.505 //y2=0.375
cc_1684 ( N_noxref_23_c_3290_n N_noxref_24_c_3333_n ) capacitor c=0.0133434f \
 //x=26.495 //y=0.54 //x2=27.065 //y2=0.995
cc_1685 ( N_noxref_23_c_3313_n N_noxref_24_c_3333_n ) capacitor c=0.0100618f \
 //x=26.495 //y=1.59 //x2=27.065 //y2=0.995
cc_1686 ( N_noxref_23_M15_noxref_s N_noxref_24_c_3333_n ) capacitor \
 c=0.0228195f //x=24.505 //y=0.375 //x2=27.065 //y2=0.995
cc_1687 ( N_noxref_23_M15_noxref_s N_noxref_24_c_3335_n ) capacitor \
 c=0.0180035f //x=24.505 //y=0.375 //x2=27.15 //y2=0.625
cc_1688 ( N_noxref_23_c_3290_n N_noxref_24_M16_noxref_d ) capacitor \
 c=0.0128018f //x=26.495 //y=0.54 //x2=25.91 //y2=0.91
cc_1689 ( N_noxref_23_c_3313_n N_noxref_24_M16_noxref_d ) capacitor \
 c=0.00879464f //x=26.495 //y=1.59 //x2=25.91 //y2=0.91
cc_1690 ( N_noxref_23_M15_noxref_s N_noxref_24_M16_noxref_d ) capacitor \
 c=0.0159202f //x=24.505 //y=0.375 //x2=25.91 //y2=0.91
cc_1691 ( N_noxref_23_M15_noxref_s N_noxref_24_M17_noxref_s ) capacitor \
 c=0.0213553f //x=24.505 //y=0.375 //x2=27.015 //y2=0.375
