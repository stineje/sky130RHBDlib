magic
tech sky130A
magscale 1 2
timestamp 1648061425
<< nmos >>
tri 144 223 160 239 se
rect 160 223 190 276
tri 54 193 84 223 se
rect 84 193 190 223
rect 54 92 84 193
tri 84 177 100 193 nw
tri 144 177 160 193 ne
tri 84 92 100 108 sw
tri 144 92 160 108 se
rect 160 92 190 193
tri 54 62 84 92 ne
rect 84 62 160 92
tri 160 62 190 92 nw
<< ndiff >>
rect 0 260 160 276
rect 0 226 8 260
rect 42 239 160 260
rect 42 226 144 239
rect 0 223 144 226
tri 144 223 160 239 nw
rect 190 260 246 276
rect 190 226 202 260
rect 236 226 246 260
rect 0 188 54 223
tri 54 193 84 223 nw
rect 0 154 8 188
rect 42 154 54 188
rect 0 120 54 154
rect 0 86 8 120
rect 42 86 54 120
tri 84 177 100 193 se
rect 100 177 144 193
tri 144 177 160 193 sw
rect 84 144 160 177
rect 84 110 106 144
rect 140 110 160 144
rect 84 108 160 110
tri 84 92 100 108 ne
rect 100 92 144 108
tri 144 92 160 108 nw
rect 190 188 246 226
rect 190 154 202 188
rect 236 154 246 188
rect 190 120 246 154
rect 0 62 54 86
tri 54 62 84 92 sw
tri 160 62 190 92 se
rect 190 86 202 120
rect 236 86 246 120
rect 190 62 246 86
rect 0 50 246 62
rect 0 16 8 50
rect 42 16 106 50
rect 140 16 202 50
rect 236 16 246 50
rect 0 0 246 16
<< ndiffc >>
rect 8 226 42 260
rect 202 226 236 260
rect 8 154 42 188
rect 8 86 42 120
rect 106 110 140 144
rect 202 154 236 188
rect 202 86 236 120
rect 8 16 42 50
rect 106 16 140 50
rect 202 16 236 50
<< poly >>
rect 160 276 190 308
<< locali >>
rect 8 260 42 276
rect 8 188 42 226
rect 202 260 236 276
rect 202 188 236 226
rect 8 120 42 154
rect 106 144 140 161
rect 106 94 140 110
rect 202 120 236 154
rect 8 50 42 86
rect 202 50 236 86
rect 42 16 106 50
rect 140 16 202 50
rect 8 0 42 16
rect 202 0 236 16
<< end >>
