magic
tech sky130A
magscale 1 2
timestamp 1648748925
<< nwell >>
rect 55 1505 89 1539
<< psubdiffcont >>
rect 55 13 89 47
<< nsubdiffcont >>
rect 55 1505 89 1539
<< viali >>
rect 55 1505 89 1539
rect 55 13 89 47
<< metal1 >>
rect 1093 945 2952 979
rect 406 871 3486 905
rect 1351 797 4604 831
rect 537 575 1822 609
rect 2461 575 2771 609
rect 2055 501 4381 535
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 888 0 -1 591
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 518 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 370 0 -1 888
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_5
timestamp 1648064633
transform 1 0 0 0 1 0
box -84 0 750 1575
use nand3x1_pcell  nand3x1_pcell_0
timestamp 1648064657
transform 1 0 666 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform -1 0 2072 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform 1 0 1850 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform -1 0 1479 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 1332 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 1110 0 -1 962
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_2
timestamp 1648064657
transform 1 0 1628 0 1 0
box -84 0 1046 1575
use nand2x1_pcell  nand2x1_pcell_2
timestamp 1648064633
transform 1 0 3256 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_18
timestamp 1648061256
transform 1 0 2812 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform -1 0 2442 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 3108 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform 1 0 2294 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform 1 0 2960 0 1 962
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_0
timestamp 1648064633
transform 1 0 2590 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 4366 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_19
timestamp 1648061256
transform 1 0 3478 0 1 888
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_1
timestamp 1648064657
transform 1 0 3922 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform 1 0 4588 0 1 814
box -53 -33 29 33
<< end >>
