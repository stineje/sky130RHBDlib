magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect 122 -30 3550 992
<< pwell >>
rect -36 1052 3501 1138
rect -36 -90 50 1052
rect -36 -176 3493 -90
<< mvpmos >>
rect 356 665 1756 765
rect 1886 665 3286 765
rect 356 509 1756 609
rect 1886 509 3286 609
rect 356 353 1756 453
rect 1886 353 3286 453
rect 356 197 1756 297
rect 1886 197 3286 297
<< mvpdiff >>
rect 356 810 1756 818
rect 356 776 418 810
rect 452 776 486 810
rect 520 776 554 810
rect 588 776 622 810
rect 656 776 690 810
rect 724 776 758 810
rect 792 776 826 810
rect 860 776 894 810
rect 928 776 962 810
rect 996 776 1030 810
rect 1064 776 1098 810
rect 1132 776 1166 810
rect 1200 776 1234 810
rect 1268 776 1302 810
rect 1336 776 1370 810
rect 1404 776 1438 810
rect 1472 776 1506 810
rect 1540 776 1574 810
rect 1608 776 1642 810
rect 1676 776 1710 810
rect 1744 776 1756 810
rect 356 765 1756 776
rect 1886 810 3286 818
rect 1886 776 1948 810
rect 1982 776 2016 810
rect 2050 776 2084 810
rect 2118 776 2152 810
rect 2186 776 2220 810
rect 2254 776 2288 810
rect 2322 776 2356 810
rect 2390 776 2424 810
rect 2458 776 2492 810
rect 2526 776 2560 810
rect 2594 776 2628 810
rect 2662 776 2696 810
rect 2730 776 2764 810
rect 2798 776 2832 810
rect 2866 776 2900 810
rect 2934 776 2968 810
rect 3002 776 3036 810
rect 3070 776 3104 810
rect 3138 776 3172 810
rect 3206 776 3240 810
rect 3274 776 3286 810
rect 1886 765 3286 776
rect 356 654 1756 665
rect 356 620 418 654
rect 452 620 486 654
rect 520 620 554 654
rect 588 620 622 654
rect 656 620 690 654
rect 724 620 758 654
rect 792 620 826 654
rect 860 620 894 654
rect 928 620 962 654
rect 996 620 1030 654
rect 1064 620 1098 654
rect 1132 620 1166 654
rect 1200 620 1234 654
rect 1268 620 1302 654
rect 1336 620 1370 654
rect 1404 620 1438 654
rect 1472 620 1506 654
rect 1540 620 1574 654
rect 1608 620 1642 654
rect 1676 620 1710 654
rect 1744 620 1756 654
rect 356 609 1756 620
rect 1886 654 3286 665
rect 1886 620 1948 654
rect 1982 620 2016 654
rect 2050 620 2084 654
rect 2118 620 2152 654
rect 2186 620 2220 654
rect 2254 620 2288 654
rect 2322 620 2356 654
rect 2390 620 2424 654
rect 2458 620 2492 654
rect 2526 620 2560 654
rect 2594 620 2628 654
rect 2662 620 2696 654
rect 2730 620 2764 654
rect 2798 620 2832 654
rect 2866 620 2900 654
rect 2934 620 2968 654
rect 3002 620 3036 654
rect 3070 620 3104 654
rect 3138 620 3172 654
rect 3206 620 3240 654
rect 3274 620 3286 654
rect 1886 609 3286 620
rect 356 498 1756 509
rect 356 464 418 498
rect 452 464 486 498
rect 520 464 554 498
rect 588 464 622 498
rect 656 464 690 498
rect 724 464 758 498
rect 792 464 826 498
rect 860 464 894 498
rect 928 464 962 498
rect 996 464 1030 498
rect 1064 464 1098 498
rect 1132 464 1166 498
rect 1200 464 1234 498
rect 1268 464 1302 498
rect 1336 464 1370 498
rect 1404 464 1438 498
rect 1472 464 1506 498
rect 1540 464 1574 498
rect 1608 464 1642 498
rect 1676 464 1710 498
rect 1744 464 1756 498
rect 356 453 1756 464
rect 1886 498 3286 509
rect 1886 464 1948 498
rect 1982 464 2016 498
rect 2050 464 2084 498
rect 2118 464 2152 498
rect 2186 464 2220 498
rect 2254 464 2288 498
rect 2322 464 2356 498
rect 2390 464 2424 498
rect 2458 464 2492 498
rect 2526 464 2560 498
rect 2594 464 2628 498
rect 2662 464 2696 498
rect 2730 464 2764 498
rect 2798 464 2832 498
rect 2866 464 2900 498
rect 2934 464 2968 498
rect 3002 464 3036 498
rect 3070 464 3104 498
rect 3138 464 3172 498
rect 3206 464 3240 498
rect 3274 464 3286 498
rect 1886 453 3286 464
rect 356 342 1756 353
rect 356 308 418 342
rect 452 308 486 342
rect 520 308 554 342
rect 588 308 622 342
rect 656 308 690 342
rect 724 308 758 342
rect 792 308 826 342
rect 860 308 894 342
rect 928 308 962 342
rect 996 308 1030 342
rect 1064 308 1098 342
rect 1132 308 1166 342
rect 1200 308 1234 342
rect 1268 308 1302 342
rect 1336 308 1370 342
rect 1404 308 1438 342
rect 1472 308 1506 342
rect 1540 308 1574 342
rect 1608 308 1642 342
rect 1676 308 1710 342
rect 1744 308 1756 342
rect 356 297 1756 308
rect 1886 342 3286 353
rect 1886 308 1948 342
rect 1982 308 2016 342
rect 2050 308 2084 342
rect 2118 308 2152 342
rect 2186 308 2220 342
rect 2254 308 2288 342
rect 2322 308 2356 342
rect 2390 308 2424 342
rect 2458 308 2492 342
rect 2526 308 2560 342
rect 2594 308 2628 342
rect 2662 308 2696 342
rect 2730 308 2764 342
rect 2798 308 2832 342
rect 2866 308 2900 342
rect 2934 308 2968 342
rect 3002 308 3036 342
rect 3070 308 3104 342
rect 3138 308 3172 342
rect 3206 308 3240 342
rect 3274 308 3286 342
rect 1886 297 3286 308
rect 356 186 1756 197
rect 356 152 418 186
rect 452 152 486 186
rect 520 152 554 186
rect 588 152 622 186
rect 656 152 690 186
rect 724 152 758 186
rect 792 152 826 186
rect 860 152 894 186
rect 928 152 962 186
rect 996 152 1030 186
rect 1064 152 1098 186
rect 1132 152 1166 186
rect 1200 152 1234 186
rect 1268 152 1302 186
rect 1336 152 1370 186
rect 1404 152 1438 186
rect 1472 152 1506 186
rect 1540 152 1574 186
rect 1608 152 1642 186
rect 1676 152 1710 186
rect 1744 152 1756 186
rect 356 144 1756 152
rect 1886 186 3286 197
rect 1886 152 1948 186
rect 1982 152 2016 186
rect 2050 152 2084 186
rect 2118 152 2152 186
rect 2186 152 2220 186
rect 2254 152 2288 186
rect 2322 152 2356 186
rect 2390 152 2424 186
rect 2458 152 2492 186
rect 2526 152 2560 186
rect 2594 152 2628 186
rect 2662 152 2696 186
rect 2730 152 2764 186
rect 2798 152 2832 186
rect 2866 152 2900 186
rect 2934 152 2968 186
rect 3002 152 3036 186
rect 3070 152 3104 186
rect 3138 152 3172 186
rect 3206 152 3240 186
rect 3274 152 3286 186
rect 1886 144 3286 152
<< mvpdiffc >>
rect 418 776 452 810
rect 486 776 520 810
rect 554 776 588 810
rect 622 776 656 810
rect 690 776 724 810
rect 758 776 792 810
rect 826 776 860 810
rect 894 776 928 810
rect 962 776 996 810
rect 1030 776 1064 810
rect 1098 776 1132 810
rect 1166 776 1200 810
rect 1234 776 1268 810
rect 1302 776 1336 810
rect 1370 776 1404 810
rect 1438 776 1472 810
rect 1506 776 1540 810
rect 1574 776 1608 810
rect 1642 776 1676 810
rect 1710 776 1744 810
rect 1948 776 1982 810
rect 2016 776 2050 810
rect 2084 776 2118 810
rect 2152 776 2186 810
rect 2220 776 2254 810
rect 2288 776 2322 810
rect 2356 776 2390 810
rect 2424 776 2458 810
rect 2492 776 2526 810
rect 2560 776 2594 810
rect 2628 776 2662 810
rect 2696 776 2730 810
rect 2764 776 2798 810
rect 2832 776 2866 810
rect 2900 776 2934 810
rect 2968 776 3002 810
rect 3036 776 3070 810
rect 3104 776 3138 810
rect 3172 776 3206 810
rect 3240 776 3274 810
rect 418 620 452 654
rect 486 620 520 654
rect 554 620 588 654
rect 622 620 656 654
rect 690 620 724 654
rect 758 620 792 654
rect 826 620 860 654
rect 894 620 928 654
rect 962 620 996 654
rect 1030 620 1064 654
rect 1098 620 1132 654
rect 1166 620 1200 654
rect 1234 620 1268 654
rect 1302 620 1336 654
rect 1370 620 1404 654
rect 1438 620 1472 654
rect 1506 620 1540 654
rect 1574 620 1608 654
rect 1642 620 1676 654
rect 1710 620 1744 654
rect 1948 620 1982 654
rect 2016 620 2050 654
rect 2084 620 2118 654
rect 2152 620 2186 654
rect 2220 620 2254 654
rect 2288 620 2322 654
rect 2356 620 2390 654
rect 2424 620 2458 654
rect 2492 620 2526 654
rect 2560 620 2594 654
rect 2628 620 2662 654
rect 2696 620 2730 654
rect 2764 620 2798 654
rect 2832 620 2866 654
rect 2900 620 2934 654
rect 2968 620 3002 654
rect 3036 620 3070 654
rect 3104 620 3138 654
rect 3172 620 3206 654
rect 3240 620 3274 654
rect 418 464 452 498
rect 486 464 520 498
rect 554 464 588 498
rect 622 464 656 498
rect 690 464 724 498
rect 758 464 792 498
rect 826 464 860 498
rect 894 464 928 498
rect 962 464 996 498
rect 1030 464 1064 498
rect 1098 464 1132 498
rect 1166 464 1200 498
rect 1234 464 1268 498
rect 1302 464 1336 498
rect 1370 464 1404 498
rect 1438 464 1472 498
rect 1506 464 1540 498
rect 1574 464 1608 498
rect 1642 464 1676 498
rect 1710 464 1744 498
rect 1948 464 1982 498
rect 2016 464 2050 498
rect 2084 464 2118 498
rect 2152 464 2186 498
rect 2220 464 2254 498
rect 2288 464 2322 498
rect 2356 464 2390 498
rect 2424 464 2458 498
rect 2492 464 2526 498
rect 2560 464 2594 498
rect 2628 464 2662 498
rect 2696 464 2730 498
rect 2764 464 2798 498
rect 2832 464 2866 498
rect 2900 464 2934 498
rect 2968 464 3002 498
rect 3036 464 3070 498
rect 3104 464 3138 498
rect 3172 464 3206 498
rect 3240 464 3274 498
rect 418 308 452 342
rect 486 308 520 342
rect 554 308 588 342
rect 622 308 656 342
rect 690 308 724 342
rect 758 308 792 342
rect 826 308 860 342
rect 894 308 928 342
rect 962 308 996 342
rect 1030 308 1064 342
rect 1098 308 1132 342
rect 1166 308 1200 342
rect 1234 308 1268 342
rect 1302 308 1336 342
rect 1370 308 1404 342
rect 1438 308 1472 342
rect 1506 308 1540 342
rect 1574 308 1608 342
rect 1642 308 1676 342
rect 1710 308 1744 342
rect 1948 308 1982 342
rect 2016 308 2050 342
rect 2084 308 2118 342
rect 2152 308 2186 342
rect 2220 308 2254 342
rect 2288 308 2322 342
rect 2356 308 2390 342
rect 2424 308 2458 342
rect 2492 308 2526 342
rect 2560 308 2594 342
rect 2628 308 2662 342
rect 2696 308 2730 342
rect 2764 308 2798 342
rect 2832 308 2866 342
rect 2900 308 2934 342
rect 2968 308 3002 342
rect 3036 308 3070 342
rect 3104 308 3138 342
rect 3172 308 3206 342
rect 3240 308 3274 342
rect 418 152 452 186
rect 486 152 520 186
rect 554 152 588 186
rect 622 152 656 186
rect 690 152 724 186
rect 758 152 792 186
rect 826 152 860 186
rect 894 152 928 186
rect 962 152 996 186
rect 1030 152 1064 186
rect 1098 152 1132 186
rect 1166 152 1200 186
rect 1234 152 1268 186
rect 1302 152 1336 186
rect 1370 152 1404 186
rect 1438 152 1472 186
rect 1506 152 1540 186
rect 1574 152 1608 186
rect 1642 152 1676 186
rect 1710 152 1744 186
rect 1948 152 1982 186
rect 2016 152 2050 186
rect 2084 152 2118 186
rect 2152 152 2186 186
rect 2220 152 2254 186
rect 2288 152 2322 186
rect 2356 152 2390 186
rect 2424 152 2458 186
rect 2492 152 2526 186
rect 2560 152 2594 186
rect 2628 152 2662 186
rect 2696 152 2730 186
rect 2764 152 2798 186
rect 2832 152 2866 186
rect 2900 152 2934 186
rect 2968 152 3002 186
rect 3036 152 3070 186
rect 3104 152 3138 186
rect 3172 152 3206 186
rect 3240 152 3274 186
<< mvpsubdiff >>
rect -10 1088 69 1112
rect 24 1078 69 1088
rect 103 1078 137 1112
rect 171 1078 205 1112
rect 239 1078 273 1112
rect 307 1078 341 1112
rect 375 1078 409 1112
rect 443 1078 477 1112
rect 511 1078 545 1112
rect 579 1078 613 1112
rect 647 1078 681 1112
rect 715 1078 749 1112
rect 783 1078 817 1112
rect 851 1078 885 1112
rect 919 1078 953 1112
rect 987 1078 1021 1112
rect 1055 1078 1089 1112
rect 1123 1078 1157 1112
rect 1191 1078 1225 1112
rect 1259 1078 1293 1112
rect 1327 1078 1361 1112
rect 1395 1078 1429 1112
rect 1463 1078 1497 1112
rect 1531 1078 1565 1112
rect 1599 1078 1633 1112
rect 1667 1078 1701 1112
rect 1735 1078 1769 1112
rect 1803 1078 1837 1112
rect 1871 1078 1905 1112
rect 1939 1078 1973 1112
rect 2007 1078 2041 1112
rect 2075 1078 2109 1112
rect 2143 1078 2177 1112
rect 2211 1078 2245 1112
rect 2279 1078 2313 1112
rect 2347 1078 2381 1112
rect 2415 1078 2449 1112
rect 2483 1078 2517 1112
rect 2551 1078 2585 1112
rect 2619 1078 2653 1112
rect 2687 1078 2721 1112
rect 2755 1078 2789 1112
rect 2823 1078 2857 1112
rect 2891 1078 2925 1112
rect 2959 1078 2993 1112
rect 3027 1078 3061 1112
rect 3095 1078 3129 1112
rect 3163 1078 3197 1112
rect 3231 1078 3265 1112
rect 3299 1078 3333 1112
rect 3367 1078 3401 1112
rect 3435 1078 3475 1112
rect -10 1020 24 1054
rect -10 952 24 986
rect -10 884 24 918
rect -10 816 24 850
rect -10 748 24 782
rect -10 680 24 714
rect -10 612 24 646
rect -10 544 24 578
rect -10 476 24 510
rect -10 408 24 442
rect -10 340 24 374
rect -10 272 24 306
rect -10 204 24 238
rect -10 136 24 170
rect -10 68 24 102
rect -10 0 24 34
rect -10 -116 24 -34
rect -10 -150 14 -116
rect 48 -150 82 -116
rect 116 -150 150 -116
rect 184 -150 218 -116
rect 252 -150 286 -116
rect 320 -150 354 -116
rect 388 -150 422 -116
rect 456 -150 490 -116
rect 524 -150 558 -116
rect 592 -150 626 -116
rect 660 -150 694 -116
rect 728 -150 762 -116
rect 796 -150 830 -116
rect 864 -150 898 -116
rect 932 -150 966 -116
rect 1000 -150 1034 -116
rect 1068 -150 1102 -116
rect 1136 -150 1170 -116
rect 1204 -150 1238 -116
rect 1272 -150 1306 -116
rect 1340 -150 1374 -116
rect 1408 -150 1442 -116
rect 1476 -150 1510 -116
rect 1544 -150 1578 -116
rect 1612 -150 1646 -116
rect 1680 -150 1714 -116
rect 1748 -150 1782 -116
rect 1816 -150 1850 -116
rect 1884 -150 1918 -116
rect 1952 -150 1986 -116
rect 2020 -150 2054 -116
rect 2088 -150 2122 -116
rect 2156 -150 2190 -116
rect 2224 -150 2258 -116
rect 2292 -150 2326 -116
rect 2360 -150 2394 -116
rect 2428 -150 2462 -116
rect 2496 -150 2530 -116
rect 2564 -150 2598 -116
rect 2632 -150 2666 -116
rect 2700 -150 2734 -116
rect 2768 -150 2802 -116
rect 2836 -150 2870 -116
rect 2904 -150 2938 -116
rect 2972 -150 3006 -116
rect 3040 -150 3074 -116
rect 3108 -150 3142 -116
rect 3176 -150 3210 -116
rect 3244 -150 3278 -116
rect 3312 -150 3346 -116
rect 3380 -150 3467 -116
<< mvnsubdiff >>
rect 188 892 256 926
rect 290 892 326 926
rect 360 892 396 926
rect 430 892 466 926
rect 500 892 536 926
rect 570 892 606 926
rect 640 892 676 926
rect 710 892 746 926
rect 780 892 816 926
rect 850 892 886 926
rect 920 892 956 926
rect 990 892 1026 926
rect 1060 892 1096 926
rect 1130 892 1166 926
rect 1200 892 1236 926
rect 1270 892 1306 926
rect 1340 892 1376 926
rect 1410 892 1446 926
rect 1480 892 1516 926
rect 1550 892 1586 926
rect 1620 892 1656 926
rect 1690 892 1725 926
rect 1759 892 1794 926
rect 1828 892 1863 926
rect 1897 892 1932 926
rect 1966 892 2001 926
rect 2035 892 2070 926
rect 2104 892 2139 926
rect 2173 892 2208 926
rect 2242 892 2277 926
rect 2311 892 2346 926
rect 2380 892 2415 926
rect 2449 892 2484 926
rect 2518 892 2553 926
rect 2587 892 2622 926
rect 2656 892 2691 926
rect 2725 892 2760 926
rect 2794 892 2829 926
rect 2863 892 2898 926
rect 2932 892 2967 926
rect 3001 892 3036 926
rect 3070 892 3105 926
rect 3139 892 3174 926
rect 3208 892 3243 926
rect 3277 892 3312 926
rect 3346 892 3381 926
rect 3415 892 3484 926
rect 188 827 222 892
rect 188 706 222 793
rect 188 638 222 672
rect 188 570 222 604
rect 188 502 222 536
rect 188 434 222 468
rect 188 366 222 400
rect 188 298 222 332
rect 188 230 222 264
rect 188 162 222 196
rect 188 94 222 128
rect 3450 70 3484 892
rect 222 60 286 70
rect 188 36 286 60
rect 320 36 354 70
rect 388 36 422 70
rect 456 36 490 70
rect 524 36 558 70
rect 592 36 626 70
rect 660 36 694 70
rect 728 36 762 70
rect 796 36 830 70
rect 864 36 898 70
rect 932 36 966 70
rect 1000 36 1034 70
rect 1068 36 1102 70
rect 1136 36 1170 70
rect 1204 36 1238 70
rect 1272 36 1306 70
rect 1340 36 1374 70
rect 1408 36 1442 70
rect 1476 36 1510 70
rect 1544 36 1578 70
rect 1612 36 1646 70
rect 1680 36 1714 70
rect 1748 36 1782 70
rect 1816 36 1850 70
rect 1884 36 1918 70
rect 1952 36 1986 70
rect 2020 36 2054 70
rect 2088 36 2122 70
rect 2156 36 2190 70
rect 2224 36 2258 70
rect 2292 36 2326 70
rect 2360 36 2394 70
rect 2428 36 2462 70
rect 2496 36 2530 70
rect 2564 36 2598 70
rect 2632 36 2666 70
rect 2700 36 2734 70
rect 2768 36 2802 70
rect 2836 36 2870 70
rect 2904 36 2938 70
rect 2972 36 3006 70
rect 3040 36 3074 70
rect 3108 36 3142 70
rect 3176 36 3210 70
rect 3244 36 3278 70
rect 3312 36 3346 70
rect 3380 36 3484 70
<< mvpsubdiffcont >>
rect -10 1054 24 1088
rect 69 1078 103 1112
rect 137 1078 171 1112
rect 205 1078 239 1112
rect 273 1078 307 1112
rect 341 1078 375 1112
rect 409 1078 443 1112
rect 477 1078 511 1112
rect 545 1078 579 1112
rect 613 1078 647 1112
rect 681 1078 715 1112
rect 749 1078 783 1112
rect 817 1078 851 1112
rect 885 1078 919 1112
rect 953 1078 987 1112
rect 1021 1078 1055 1112
rect 1089 1078 1123 1112
rect 1157 1078 1191 1112
rect 1225 1078 1259 1112
rect 1293 1078 1327 1112
rect 1361 1078 1395 1112
rect 1429 1078 1463 1112
rect 1497 1078 1531 1112
rect 1565 1078 1599 1112
rect 1633 1078 1667 1112
rect 1701 1078 1735 1112
rect 1769 1078 1803 1112
rect 1837 1078 1871 1112
rect 1905 1078 1939 1112
rect 1973 1078 2007 1112
rect 2041 1078 2075 1112
rect 2109 1078 2143 1112
rect 2177 1078 2211 1112
rect 2245 1078 2279 1112
rect 2313 1078 2347 1112
rect 2381 1078 2415 1112
rect 2449 1078 2483 1112
rect 2517 1078 2551 1112
rect 2585 1078 2619 1112
rect 2653 1078 2687 1112
rect 2721 1078 2755 1112
rect 2789 1078 2823 1112
rect 2857 1078 2891 1112
rect 2925 1078 2959 1112
rect 2993 1078 3027 1112
rect 3061 1078 3095 1112
rect 3129 1078 3163 1112
rect 3197 1078 3231 1112
rect 3265 1078 3299 1112
rect 3333 1078 3367 1112
rect 3401 1078 3435 1112
rect -10 986 24 1020
rect -10 918 24 952
rect -10 850 24 884
rect -10 782 24 816
rect -10 714 24 748
rect -10 646 24 680
rect -10 578 24 612
rect -10 510 24 544
rect -10 442 24 476
rect -10 374 24 408
rect -10 306 24 340
rect -10 238 24 272
rect -10 170 24 204
rect -10 102 24 136
rect -10 34 24 68
rect -10 -34 24 0
rect 14 -150 48 -116
rect 82 -150 116 -116
rect 150 -150 184 -116
rect 218 -150 252 -116
rect 286 -150 320 -116
rect 354 -150 388 -116
rect 422 -150 456 -116
rect 490 -150 524 -116
rect 558 -150 592 -116
rect 626 -150 660 -116
rect 694 -150 728 -116
rect 762 -150 796 -116
rect 830 -150 864 -116
rect 898 -150 932 -116
rect 966 -150 1000 -116
rect 1034 -150 1068 -116
rect 1102 -150 1136 -116
rect 1170 -150 1204 -116
rect 1238 -150 1272 -116
rect 1306 -150 1340 -116
rect 1374 -150 1408 -116
rect 1442 -150 1476 -116
rect 1510 -150 1544 -116
rect 1578 -150 1612 -116
rect 1646 -150 1680 -116
rect 1714 -150 1748 -116
rect 1782 -150 1816 -116
rect 1850 -150 1884 -116
rect 1918 -150 1952 -116
rect 1986 -150 2020 -116
rect 2054 -150 2088 -116
rect 2122 -150 2156 -116
rect 2190 -150 2224 -116
rect 2258 -150 2292 -116
rect 2326 -150 2360 -116
rect 2394 -150 2428 -116
rect 2462 -150 2496 -116
rect 2530 -150 2564 -116
rect 2598 -150 2632 -116
rect 2666 -150 2700 -116
rect 2734 -150 2768 -116
rect 2802 -150 2836 -116
rect 2870 -150 2904 -116
rect 2938 -150 2972 -116
rect 3006 -150 3040 -116
rect 3074 -150 3108 -116
rect 3142 -150 3176 -116
rect 3210 -150 3244 -116
rect 3278 -150 3312 -116
rect 3346 -150 3380 -116
<< mvnsubdiffcont >>
rect 256 892 290 926
rect 326 892 360 926
rect 396 892 430 926
rect 466 892 500 926
rect 536 892 570 926
rect 606 892 640 926
rect 676 892 710 926
rect 746 892 780 926
rect 816 892 850 926
rect 886 892 920 926
rect 956 892 990 926
rect 1026 892 1060 926
rect 1096 892 1130 926
rect 1166 892 1200 926
rect 1236 892 1270 926
rect 1306 892 1340 926
rect 1376 892 1410 926
rect 1446 892 1480 926
rect 1516 892 1550 926
rect 1586 892 1620 926
rect 1656 892 1690 926
rect 1725 892 1759 926
rect 1794 892 1828 926
rect 1863 892 1897 926
rect 1932 892 1966 926
rect 2001 892 2035 926
rect 2070 892 2104 926
rect 2139 892 2173 926
rect 2208 892 2242 926
rect 2277 892 2311 926
rect 2346 892 2380 926
rect 2415 892 2449 926
rect 2484 892 2518 926
rect 2553 892 2587 926
rect 2622 892 2656 926
rect 2691 892 2725 926
rect 2760 892 2794 926
rect 2829 892 2863 926
rect 2898 892 2932 926
rect 2967 892 3001 926
rect 3036 892 3070 926
rect 3105 892 3139 926
rect 3174 892 3208 926
rect 3243 892 3277 926
rect 3312 892 3346 926
rect 3381 892 3415 926
rect 188 793 222 827
rect 188 672 222 706
rect 188 604 222 638
rect 188 536 222 570
rect 188 468 222 502
rect 188 400 222 434
rect 188 332 222 366
rect 188 264 222 298
rect 188 196 222 230
rect 188 128 222 162
rect 188 60 222 94
rect 286 36 320 70
rect 354 36 388 70
rect 422 36 456 70
rect 490 36 524 70
rect 558 36 592 70
rect 626 36 660 70
rect 694 36 728 70
rect 762 36 796 70
rect 830 36 864 70
rect 898 36 932 70
rect 966 36 1000 70
rect 1034 36 1068 70
rect 1102 36 1136 70
rect 1170 36 1204 70
rect 1238 36 1272 70
rect 1306 36 1340 70
rect 1374 36 1408 70
rect 1442 36 1476 70
rect 1510 36 1544 70
rect 1578 36 1612 70
rect 1646 36 1680 70
rect 1714 36 1748 70
rect 1782 36 1816 70
rect 1850 36 1884 70
rect 1918 36 1952 70
rect 1986 36 2020 70
rect 2054 36 2088 70
rect 2122 36 2156 70
rect 2190 36 2224 70
rect 2258 36 2292 70
rect 2326 36 2360 70
rect 2394 36 2428 70
rect 2462 36 2496 70
rect 2530 36 2564 70
rect 2598 36 2632 70
rect 2666 36 2700 70
rect 2734 36 2768 70
rect 2802 36 2836 70
rect 2870 36 2904 70
rect 2938 36 2972 70
rect 3006 36 3040 70
rect 3074 36 3108 70
rect 3142 36 3176 70
rect 3210 36 3244 70
rect 3278 36 3312 70
rect 3346 36 3380 70
<< poly >>
rect 252 749 356 765
rect 252 715 274 749
rect 308 715 356 749
rect 252 677 356 715
rect 252 643 274 677
rect 308 665 356 677
rect 1756 726 1886 765
rect 1756 692 1804 726
rect 1838 692 1886 726
rect 1756 665 1886 692
rect 3286 746 3390 765
rect 3286 712 3334 746
rect 3368 712 3390 746
rect 3286 674 3390 712
rect 3286 665 3334 674
rect 308 643 330 665
rect 252 609 330 643
rect 1782 657 1860 665
rect 1782 623 1804 657
rect 1838 623 1860 657
rect 1782 609 1860 623
rect 3312 640 3334 665
rect 3368 640 3390 674
rect 3312 609 3390 640
rect 252 605 356 609
rect 252 571 274 605
rect 308 571 356 605
rect 252 533 356 571
rect 252 499 274 533
rect 308 509 356 533
rect 1756 588 1886 609
rect 1756 554 1804 588
rect 1838 554 1886 588
rect 1756 519 1886 554
rect 1756 509 1804 519
rect 308 499 330 509
rect 252 461 330 499
rect 252 427 274 461
rect 308 453 330 461
rect 1782 485 1804 509
rect 1838 509 1886 519
rect 3286 602 3390 609
rect 3286 568 3334 602
rect 3368 568 3390 602
rect 3286 531 3390 568
rect 3286 509 3334 531
rect 1838 485 1860 509
rect 1782 453 1860 485
rect 3312 497 3334 509
rect 3368 497 3390 531
rect 3312 460 3390 497
rect 3312 453 3334 460
rect 308 427 356 453
rect 252 389 356 427
rect 252 355 274 389
rect 308 355 356 389
rect 252 353 356 355
rect 1756 451 1886 453
rect 1756 417 1804 451
rect 1838 417 1886 451
rect 1756 383 1886 417
rect 1756 353 1804 383
rect 252 318 330 353
rect 252 284 274 318
rect 308 297 330 318
rect 1782 349 1804 353
rect 1838 353 1886 383
rect 3286 426 3334 453
rect 3368 426 3390 460
rect 3286 389 3390 426
rect 3286 355 3334 389
rect 3368 355 3390 389
rect 3286 353 3390 355
rect 1838 349 1860 353
rect 1782 315 1860 349
rect 1782 297 1804 315
rect 308 284 356 297
rect 252 247 356 284
rect 252 213 274 247
rect 308 213 356 247
rect 252 197 356 213
rect 1756 281 1804 297
rect 1838 297 1860 315
rect 3312 318 3390 353
rect 3312 297 3334 318
rect 1838 281 1886 297
rect 1756 247 1886 281
rect 1756 213 1804 247
rect 1838 213 1886 247
rect 1756 197 1886 213
rect 3286 284 3334 297
rect 3368 284 3390 318
rect 3286 247 3390 284
rect 3286 213 3334 247
rect 3368 213 3390 247
rect 3286 197 3390 213
<< polycont >>
rect 274 715 308 749
rect 274 643 308 677
rect 1804 692 1838 726
rect 3334 712 3368 746
rect 1804 623 1838 657
rect 3334 640 3368 674
rect 274 571 308 605
rect 274 499 308 533
rect 1804 554 1838 588
rect 274 427 308 461
rect 1804 485 1838 519
rect 3334 568 3368 602
rect 3334 497 3368 531
rect 274 355 308 389
rect 1804 417 1838 451
rect 274 284 308 318
rect 1804 349 1838 383
rect 3334 426 3368 460
rect 3334 355 3368 389
rect 274 213 308 247
rect 1804 281 1838 315
rect 1804 213 1838 247
rect 3334 284 3368 318
rect 3334 213 3368 247
<< locali >>
rect -10 1100 69 1112
rect 24 1078 69 1100
rect 135 1078 137 1112
rect 171 1078 173 1112
rect 239 1078 245 1112
rect 307 1078 317 1112
rect 375 1078 389 1112
rect 443 1078 461 1112
rect 511 1078 533 1112
rect 579 1078 605 1112
rect 647 1078 677 1112
rect 715 1078 749 1112
rect 783 1078 817 1112
rect 855 1078 885 1112
rect 927 1078 953 1112
rect 999 1078 1021 1112
rect 1071 1078 1089 1112
rect 1143 1078 1157 1112
rect 1215 1078 1225 1112
rect 1287 1078 1293 1112
rect 1359 1078 1361 1112
rect 1395 1078 1397 1112
rect 1463 1078 1469 1112
rect 1531 1078 1541 1112
rect 1599 1078 1613 1112
rect 1667 1078 1685 1112
rect 1735 1078 1757 1112
rect 1803 1078 1829 1112
rect 1871 1078 1901 1112
rect 1939 1078 1973 1112
rect 2007 1078 2041 1112
rect 2079 1078 2109 1112
rect 2151 1078 2177 1112
rect 2223 1078 2245 1112
rect 2295 1078 2313 1112
rect 2367 1078 2381 1112
rect 2439 1078 2449 1112
rect 2511 1078 2517 1112
rect 2583 1078 2585 1112
rect 2619 1078 2621 1112
rect 2687 1078 2693 1112
rect 2755 1078 2765 1112
rect 2823 1078 2837 1112
rect 2891 1078 2909 1112
rect 2959 1078 2981 1112
rect 3027 1078 3053 1112
rect 3095 1078 3125 1112
rect 3163 1078 3197 1112
rect 3231 1078 3265 1112
rect 3303 1078 3333 1112
rect 3375 1078 3401 1112
rect 3447 1078 3475 1112
rect -10 1028 24 1054
rect -10 956 24 986
rect -10 884 24 918
rect -10 816 24 850
rect -10 748 24 778
rect -10 680 24 706
rect -10 612 24 634
rect -10 544 24 562
rect -10 476 24 490
rect -10 408 24 418
rect -10 340 24 346
rect -10 272 24 274
rect -10 236 24 238
rect -10 164 24 170
rect -10 92 24 102
rect 188 892 256 926
rect 290 892 326 926
rect 360 892 396 926
rect 430 892 466 926
rect 500 892 536 926
rect 570 892 606 926
rect 640 892 676 926
rect 710 892 746 926
rect 780 892 816 926
rect 850 892 886 926
rect 920 892 956 926
rect 990 892 1026 926
rect 1060 892 1096 926
rect 1130 892 1166 926
rect 1200 892 1236 926
rect 1270 892 1306 926
rect 1340 892 1376 926
rect 1410 892 1446 926
rect 1480 892 1516 926
rect 1550 892 1586 926
rect 1620 892 1656 926
rect 1690 892 1725 926
rect 1759 892 1794 926
rect 1828 892 1863 926
rect 1897 892 1932 926
rect 1966 892 2001 926
rect 2035 892 2070 926
rect 2104 892 2139 926
rect 2173 892 2208 926
rect 2242 892 2277 926
rect 2311 892 2346 926
rect 2380 892 2415 926
rect 2449 892 2484 926
rect 2518 892 2553 926
rect 2587 892 2622 926
rect 2656 892 2691 926
rect 2725 892 2760 926
rect 2794 892 2829 926
rect 2863 892 2898 926
rect 2932 892 2967 926
rect 3001 892 3036 926
rect 3070 892 3105 926
rect 3139 892 3174 926
rect 3208 892 3243 926
rect 3277 892 3312 926
rect 3346 892 3381 926
rect 3415 892 3484 926
rect 188 827 3484 892
rect 222 810 3484 827
rect 222 799 358 810
rect 188 730 222 793
rect 392 776 418 810
rect 464 776 486 810
rect 536 776 554 810
rect 608 776 622 810
rect 680 776 690 810
rect 752 776 758 810
rect 824 776 826 810
rect 860 776 862 810
rect 928 776 934 810
rect 996 776 1006 810
rect 1064 776 1078 810
rect 1132 776 1150 810
rect 1200 776 1222 810
rect 1268 776 1294 810
rect 1336 776 1366 810
rect 1404 776 1438 810
rect 1472 776 1506 810
rect 1544 776 1574 810
rect 1616 776 1642 810
rect 1688 776 1710 810
rect 1760 776 1888 810
rect 1922 776 1948 810
rect 1994 776 2016 810
rect 2066 776 2084 810
rect 2138 776 2152 810
rect 2210 776 2220 810
rect 2282 776 2288 810
rect 2354 776 2356 810
rect 2390 776 2392 810
rect 2458 776 2464 810
rect 2526 776 2536 810
rect 2594 776 2608 810
rect 2662 776 2680 810
rect 2730 776 2752 810
rect 2798 776 2824 810
rect 2866 776 2896 810
rect 2934 776 2968 810
rect 3002 776 3036 810
rect 3074 776 3104 810
rect 3146 776 3172 810
rect 3218 776 3240 810
rect 3290 804 3484 810
rect 3290 798 3450 804
rect 3290 776 3294 798
rect 3420 776 3450 798
rect 188 658 222 672
rect 188 586 222 604
rect 188 514 222 536
rect 188 442 222 468
rect 188 370 222 400
rect 188 298 222 332
rect 188 230 222 264
rect 274 749 308 765
rect 3334 746 3368 762
rect 274 677 308 715
rect 1804 726 1838 742
rect 1804 657 1838 692
rect 274 605 308 643
rect 392 620 418 654
rect 464 620 486 654
rect 536 620 554 654
rect 608 620 622 654
rect 680 620 690 654
rect 752 620 758 654
rect 824 620 826 654
rect 860 620 862 654
rect 928 620 934 654
rect 996 620 1006 654
rect 1064 620 1078 654
rect 1132 620 1150 654
rect 1200 620 1222 654
rect 1268 620 1294 654
rect 1336 620 1366 654
rect 1404 620 1438 654
rect 1472 620 1506 654
rect 1544 620 1574 654
rect 1616 620 1642 654
rect 1688 620 1710 654
rect 3334 674 3368 712
rect 1804 588 1838 623
rect 1922 620 1948 654
rect 1994 620 2016 654
rect 2066 620 2084 654
rect 2138 620 2152 654
rect 2210 620 2220 654
rect 2282 620 2288 654
rect 2354 620 2356 654
rect 2390 620 2392 654
rect 2458 620 2464 654
rect 2526 620 2536 654
rect 2594 620 2608 654
rect 2662 620 2680 654
rect 2730 620 2752 654
rect 2798 620 2824 654
rect 2866 620 2896 654
rect 2934 620 2968 654
rect 3002 620 3036 654
rect 3074 620 3104 654
rect 3146 620 3172 654
rect 3218 620 3240 654
rect 3334 602 3368 640
rect 274 541 286 571
rect 320 541 358 575
rect 1838 554 1863 575
rect 1825 541 1863 554
rect 3295 541 3333 575
rect 3367 541 3368 568
rect 274 533 308 541
rect 274 461 308 499
rect 1804 519 1838 541
rect 392 464 418 498
rect 464 464 486 498
rect 536 464 554 498
rect 608 464 622 498
rect 680 464 690 498
rect 752 464 758 498
rect 824 464 826 498
rect 860 464 862 498
rect 928 464 934 498
rect 996 464 1006 498
rect 1064 464 1078 498
rect 1132 464 1150 498
rect 1200 464 1222 498
rect 1268 464 1294 498
rect 1336 464 1366 498
rect 1404 464 1438 498
rect 1472 464 1506 498
rect 1544 464 1574 498
rect 1616 464 1642 498
rect 1688 464 1710 498
rect 3334 531 3368 541
rect 274 389 308 427
rect 274 318 308 355
rect 1804 451 1838 485
rect 1922 464 1948 498
rect 1994 464 2016 498
rect 2066 464 2084 498
rect 2138 464 2152 498
rect 2210 464 2220 498
rect 2282 464 2288 498
rect 2354 464 2356 498
rect 2390 464 2392 498
rect 2458 464 2464 498
rect 2526 464 2536 498
rect 2594 464 2608 498
rect 2662 464 2680 498
rect 2730 464 2752 498
rect 2798 464 2824 498
rect 2866 464 2896 498
rect 2934 464 2968 498
rect 3002 464 3036 498
rect 3074 464 3104 498
rect 3146 464 3172 498
rect 3218 464 3240 498
rect 1804 383 1838 417
rect 392 308 418 342
rect 464 308 486 342
rect 536 308 554 342
rect 608 308 622 342
rect 680 308 690 342
rect 752 308 758 342
rect 824 308 826 342
rect 860 308 862 342
rect 928 308 934 342
rect 996 308 1006 342
rect 1064 308 1078 342
rect 1132 308 1150 342
rect 1200 308 1222 342
rect 1268 308 1294 342
rect 1336 308 1366 342
rect 1404 308 1438 342
rect 1472 308 1506 342
rect 1544 308 1574 342
rect 1616 308 1642 342
rect 1688 308 1710 342
rect 1804 315 1838 349
rect 3334 460 3368 497
rect 3334 389 3368 426
rect 274 247 308 284
rect 274 197 308 213
rect 1922 308 1948 342
rect 1994 308 2016 342
rect 2066 308 2084 342
rect 2138 308 2152 342
rect 2210 308 2220 342
rect 2282 308 2288 342
rect 2354 308 2356 342
rect 2390 308 2392 342
rect 2458 308 2464 342
rect 2526 308 2536 342
rect 2594 308 2608 342
rect 2662 308 2680 342
rect 2730 308 2752 342
rect 2798 308 2824 342
rect 2866 308 2896 342
rect 2934 308 2968 342
rect 3002 308 3036 342
rect 3074 308 3104 342
rect 3146 308 3172 342
rect 3218 308 3240 342
rect 3334 318 3368 355
rect 1804 247 1838 281
rect 1804 197 1838 213
rect 3334 247 3368 284
rect 3334 197 3368 213
rect 3450 732 3484 770
rect 3450 660 3484 698
rect 3450 588 3484 626
rect 3450 516 3484 554
rect 3450 444 3484 482
rect 3450 372 3484 410
rect 3450 300 3484 338
rect 3450 228 3484 266
rect 188 162 222 192
rect 392 152 418 186
rect 464 152 486 186
rect 536 152 554 186
rect 608 152 622 186
rect 680 152 690 186
rect 752 152 758 186
rect 824 152 826 186
rect 860 152 862 186
rect 928 152 934 186
rect 996 152 1006 186
rect 1064 152 1078 186
rect 1132 152 1150 186
rect 1200 152 1222 186
rect 1268 152 1294 186
rect 1336 152 1366 186
rect 1404 152 1438 186
rect 1472 152 1506 186
rect 1544 152 1574 186
rect 1616 152 1642 186
rect 1688 152 1710 186
rect 1922 152 1948 186
rect 1994 152 2016 186
rect 2066 152 2084 186
rect 2138 152 2152 186
rect 2210 152 2220 186
rect 2282 152 2288 186
rect 2354 152 2356 186
rect 2390 152 2392 186
rect 2458 152 2464 186
rect 2526 152 2536 186
rect 2594 152 2608 186
rect 2662 152 2680 186
rect 2730 152 2752 186
rect 2798 152 2824 186
rect 2866 152 2896 186
rect 2934 152 2968 186
rect 3002 152 3036 186
rect 3074 152 3104 186
rect 3146 152 3172 186
rect 3218 152 3240 186
rect 3450 155 3484 194
rect 188 94 222 120
rect 3450 82 3484 121
rect 222 48 286 70
rect 188 36 286 48
rect 320 36 322 70
rect 388 36 394 70
rect 456 36 466 70
rect 524 36 538 70
rect 592 36 610 70
rect 660 36 682 70
rect 728 36 754 70
rect 796 36 826 70
rect 864 36 898 70
rect 932 36 966 70
rect 1004 36 1034 70
rect 1076 36 1102 70
rect 1148 36 1170 70
rect 1220 36 1238 70
rect 1292 36 1306 70
rect 1364 36 1374 70
rect 1436 36 1442 70
rect 1508 36 1510 70
rect 1544 36 1546 70
rect 1612 36 1618 70
rect 1680 36 1690 70
rect 1748 36 1762 70
rect 1816 36 1834 70
rect 1884 36 1906 70
rect 1952 36 1978 70
rect 2020 36 2050 70
rect 2088 36 2122 70
rect 2156 36 2190 70
rect 2228 36 2258 70
rect 2300 36 2326 70
rect 2372 36 2394 70
rect 2444 36 2462 70
rect 2516 36 2530 70
rect 2588 36 2598 70
rect 2660 36 2666 70
rect 2732 36 2734 70
rect 2768 36 2770 70
rect 2836 36 2842 70
rect 2904 36 2914 70
rect 2972 36 2986 70
rect 3040 36 3058 70
rect 3108 36 3130 70
rect 3176 36 3202 70
rect 3244 36 3274 70
rect 3312 36 3346 70
rect 3380 48 3450 70
rect 3380 36 3484 48
rect -10 20 24 34
rect -10 -116 24 -34
rect 1214 -116 1254 -104
rect 1288 -116 1328 -104
rect 1362 -116 1402 -104
rect 1436 -116 1476 -104
rect -10 -150 2 -116
rect 48 -150 74 -116
rect 116 -150 146 -116
rect 184 -150 218 -116
rect 252 -150 286 -116
rect 324 -150 354 -116
rect 396 -150 422 -116
rect 468 -150 490 -116
rect 540 -150 558 -116
rect 612 -150 626 -116
rect 684 -150 694 -116
rect 756 -150 762 -116
rect 828 -150 830 -116
rect 864 -150 866 -116
rect 932 -150 938 -116
rect 1000 -150 1010 -116
rect 1068 -150 1082 -116
rect 1136 -150 1170 -116
rect 1214 -138 1238 -116
rect 1288 -138 1306 -116
rect 1362 -138 1374 -116
rect 1436 -138 1442 -116
rect 1204 -150 1238 -138
rect 1272 -150 1306 -138
rect 1340 -150 1374 -138
rect 1408 -150 1442 -138
rect 1510 -116 1550 -104
rect 1584 -116 1624 -104
rect 1658 -116 1698 -104
rect 1732 -116 1772 -104
rect 1806 -116 1846 -104
rect 1880 -116 1920 -104
rect 1954 -116 1994 -104
rect 2028 -116 2068 -104
rect 2102 -116 2142 -104
rect 2176 -116 2216 -104
rect 2250 -116 2290 -104
rect 2324 -116 2364 -104
rect 2398 -116 2438 -104
rect 2472 -116 2512 -104
rect 2546 -116 2586 -104
rect 2620 -116 2660 -104
rect 2694 -116 2734 -104
rect 2768 -116 2808 -104
rect 2842 -116 2882 -104
rect 2916 -116 2956 -104
rect 2990 -116 3030 -104
rect 3064 -116 3104 -104
rect 3138 -116 3178 -104
rect 3212 -116 3252 -104
rect 3286 -116 3326 -104
rect 3360 -116 3400 -104
rect 1476 -150 1510 -138
rect 1544 -138 1550 -116
rect 1612 -138 1624 -116
rect 1680 -138 1698 -116
rect 1748 -138 1772 -116
rect 1816 -138 1846 -116
rect 1544 -150 1578 -138
rect 1612 -150 1646 -138
rect 1680 -150 1714 -138
rect 1748 -150 1782 -138
rect 1816 -150 1850 -138
rect 1884 -150 1918 -116
rect 1954 -138 1986 -116
rect 2028 -138 2054 -116
rect 2102 -138 2122 -116
rect 2176 -138 2190 -116
rect 2250 -138 2258 -116
rect 2324 -138 2326 -116
rect 1952 -150 1986 -138
rect 2020 -150 2054 -138
rect 2088 -150 2122 -138
rect 2156 -150 2190 -138
rect 2224 -150 2258 -138
rect 2292 -150 2326 -138
rect 2360 -138 2364 -116
rect 2428 -138 2438 -116
rect 2496 -138 2512 -116
rect 2564 -138 2586 -116
rect 2632 -138 2660 -116
rect 2360 -150 2394 -138
rect 2428 -150 2462 -138
rect 2496 -150 2530 -138
rect 2564 -150 2598 -138
rect 2632 -150 2666 -138
rect 2700 -150 2734 -116
rect 2768 -150 2802 -116
rect 2842 -138 2870 -116
rect 2916 -138 2938 -116
rect 2990 -138 3006 -116
rect 3064 -138 3074 -116
rect 3138 -138 3142 -116
rect 2836 -150 2870 -138
rect 2904 -150 2938 -138
rect 2972 -150 3006 -138
rect 3040 -150 3074 -138
rect 3108 -150 3142 -138
rect 3176 -138 3178 -116
rect 3244 -138 3252 -116
rect 3312 -138 3326 -116
rect 3380 -138 3400 -116
rect 3434 -138 3467 -116
rect 3176 -150 3210 -138
rect 3244 -150 3278 -138
rect 3312 -150 3346 -138
rect 3380 -150 3467 -138
<< viali >>
rect -10 1088 24 1100
rect -10 1066 24 1088
rect 101 1078 103 1112
rect 103 1078 135 1112
rect 173 1078 205 1112
rect 205 1078 207 1112
rect 245 1078 273 1112
rect 273 1078 279 1112
rect 317 1078 341 1112
rect 341 1078 351 1112
rect 389 1078 409 1112
rect 409 1078 423 1112
rect 461 1078 477 1112
rect 477 1078 495 1112
rect 533 1078 545 1112
rect 545 1078 567 1112
rect 605 1078 613 1112
rect 613 1078 639 1112
rect 677 1078 681 1112
rect 681 1078 711 1112
rect 749 1078 783 1112
rect 821 1078 851 1112
rect 851 1078 855 1112
rect 893 1078 919 1112
rect 919 1078 927 1112
rect 965 1078 987 1112
rect 987 1078 999 1112
rect 1037 1078 1055 1112
rect 1055 1078 1071 1112
rect 1109 1078 1123 1112
rect 1123 1078 1143 1112
rect 1181 1078 1191 1112
rect 1191 1078 1215 1112
rect 1253 1078 1259 1112
rect 1259 1078 1287 1112
rect 1325 1078 1327 1112
rect 1327 1078 1359 1112
rect 1397 1078 1429 1112
rect 1429 1078 1431 1112
rect 1469 1078 1497 1112
rect 1497 1078 1503 1112
rect 1541 1078 1565 1112
rect 1565 1078 1575 1112
rect 1613 1078 1633 1112
rect 1633 1078 1647 1112
rect 1685 1078 1701 1112
rect 1701 1078 1719 1112
rect 1757 1078 1769 1112
rect 1769 1078 1791 1112
rect 1829 1078 1837 1112
rect 1837 1078 1863 1112
rect 1901 1078 1905 1112
rect 1905 1078 1935 1112
rect 1973 1078 2007 1112
rect 2045 1078 2075 1112
rect 2075 1078 2079 1112
rect 2117 1078 2143 1112
rect 2143 1078 2151 1112
rect 2189 1078 2211 1112
rect 2211 1078 2223 1112
rect 2261 1078 2279 1112
rect 2279 1078 2295 1112
rect 2333 1078 2347 1112
rect 2347 1078 2367 1112
rect 2405 1078 2415 1112
rect 2415 1078 2439 1112
rect 2477 1078 2483 1112
rect 2483 1078 2511 1112
rect 2549 1078 2551 1112
rect 2551 1078 2583 1112
rect 2621 1078 2653 1112
rect 2653 1078 2655 1112
rect 2693 1078 2721 1112
rect 2721 1078 2727 1112
rect 2765 1078 2789 1112
rect 2789 1078 2799 1112
rect 2837 1078 2857 1112
rect 2857 1078 2871 1112
rect 2909 1078 2925 1112
rect 2925 1078 2943 1112
rect 2981 1078 2993 1112
rect 2993 1078 3015 1112
rect 3053 1078 3061 1112
rect 3061 1078 3087 1112
rect 3125 1078 3129 1112
rect 3129 1078 3159 1112
rect 3197 1078 3231 1112
rect 3269 1078 3299 1112
rect 3299 1078 3303 1112
rect 3341 1078 3367 1112
rect 3367 1078 3375 1112
rect 3413 1078 3435 1112
rect 3435 1078 3447 1112
rect -10 1020 24 1028
rect -10 994 24 1020
rect -10 952 24 956
rect -10 922 24 952
rect -10 850 24 884
rect -10 782 24 812
rect -10 778 24 782
rect -10 714 24 740
rect -10 706 24 714
rect -10 646 24 668
rect -10 634 24 646
rect -10 578 24 596
rect -10 562 24 578
rect -10 510 24 524
rect -10 490 24 510
rect -10 442 24 452
rect -10 418 24 442
rect -10 374 24 380
rect -10 346 24 374
rect -10 306 24 308
rect -10 274 24 306
rect -10 204 24 236
rect -10 202 24 204
rect -10 136 24 164
rect -10 130 24 136
rect -10 68 24 92
rect -10 58 24 68
rect 358 776 392 810
rect 430 776 452 810
rect 452 776 464 810
rect 502 776 520 810
rect 520 776 536 810
rect 574 776 588 810
rect 588 776 608 810
rect 646 776 656 810
rect 656 776 680 810
rect 718 776 724 810
rect 724 776 752 810
rect 790 776 792 810
rect 792 776 824 810
rect 862 776 894 810
rect 894 776 896 810
rect 934 776 962 810
rect 962 776 968 810
rect 1006 776 1030 810
rect 1030 776 1040 810
rect 1078 776 1098 810
rect 1098 776 1112 810
rect 1150 776 1166 810
rect 1166 776 1184 810
rect 1222 776 1234 810
rect 1234 776 1256 810
rect 1294 776 1302 810
rect 1302 776 1328 810
rect 1366 776 1370 810
rect 1370 776 1400 810
rect 1438 776 1472 810
rect 1510 776 1540 810
rect 1540 776 1544 810
rect 1582 776 1608 810
rect 1608 776 1616 810
rect 1654 776 1676 810
rect 1676 776 1688 810
rect 1726 776 1744 810
rect 1744 776 1760 810
rect 1888 776 1922 810
rect 1960 776 1982 810
rect 1982 776 1994 810
rect 2032 776 2050 810
rect 2050 776 2066 810
rect 2104 776 2118 810
rect 2118 776 2138 810
rect 2176 776 2186 810
rect 2186 776 2210 810
rect 2248 776 2254 810
rect 2254 776 2282 810
rect 2320 776 2322 810
rect 2322 776 2354 810
rect 2392 776 2424 810
rect 2424 776 2426 810
rect 2464 776 2492 810
rect 2492 776 2498 810
rect 2536 776 2560 810
rect 2560 776 2570 810
rect 2608 776 2628 810
rect 2628 776 2642 810
rect 2680 776 2696 810
rect 2696 776 2714 810
rect 2752 776 2764 810
rect 2764 776 2786 810
rect 2824 776 2832 810
rect 2832 776 2858 810
rect 2896 776 2900 810
rect 2900 776 2930 810
rect 2968 776 3002 810
rect 3040 776 3070 810
rect 3070 776 3074 810
rect 3112 776 3138 810
rect 3138 776 3146 810
rect 3184 776 3206 810
rect 3206 776 3218 810
rect 3256 776 3274 810
rect 3274 776 3290 810
rect 3450 770 3484 804
rect 188 706 222 730
rect 188 696 222 706
rect 188 638 222 658
rect 188 624 222 638
rect 188 570 222 586
rect 188 552 222 570
rect 188 502 222 514
rect 188 480 222 502
rect 188 434 222 442
rect 188 408 222 434
rect 188 366 222 370
rect 188 336 222 366
rect 188 264 222 298
rect 188 196 222 226
rect 358 620 392 654
rect 430 620 452 654
rect 452 620 464 654
rect 502 620 520 654
rect 520 620 536 654
rect 574 620 588 654
rect 588 620 608 654
rect 646 620 656 654
rect 656 620 680 654
rect 718 620 724 654
rect 724 620 752 654
rect 790 620 792 654
rect 792 620 824 654
rect 862 620 894 654
rect 894 620 896 654
rect 934 620 962 654
rect 962 620 968 654
rect 1006 620 1030 654
rect 1030 620 1040 654
rect 1078 620 1098 654
rect 1098 620 1112 654
rect 1150 620 1166 654
rect 1166 620 1184 654
rect 1222 620 1234 654
rect 1234 620 1256 654
rect 1294 620 1302 654
rect 1302 620 1328 654
rect 1366 620 1370 654
rect 1370 620 1400 654
rect 1438 620 1472 654
rect 1510 620 1540 654
rect 1540 620 1544 654
rect 1582 620 1608 654
rect 1608 620 1616 654
rect 1654 620 1676 654
rect 1676 620 1688 654
rect 1726 620 1744 654
rect 1744 620 1760 654
rect 1888 620 1922 654
rect 1960 620 1982 654
rect 1982 620 1994 654
rect 2032 620 2050 654
rect 2050 620 2066 654
rect 2104 620 2118 654
rect 2118 620 2138 654
rect 2176 620 2186 654
rect 2186 620 2210 654
rect 2248 620 2254 654
rect 2254 620 2282 654
rect 2320 620 2322 654
rect 2322 620 2354 654
rect 2392 620 2424 654
rect 2424 620 2426 654
rect 2464 620 2492 654
rect 2492 620 2498 654
rect 2536 620 2560 654
rect 2560 620 2570 654
rect 2608 620 2628 654
rect 2628 620 2642 654
rect 2680 620 2696 654
rect 2696 620 2714 654
rect 2752 620 2764 654
rect 2764 620 2786 654
rect 2824 620 2832 654
rect 2832 620 2858 654
rect 2896 620 2900 654
rect 2900 620 2930 654
rect 2968 620 3002 654
rect 3040 620 3070 654
rect 3070 620 3074 654
rect 3112 620 3138 654
rect 3138 620 3146 654
rect 3184 620 3206 654
rect 3206 620 3218 654
rect 3256 620 3274 654
rect 3274 620 3290 654
rect 286 571 308 575
rect 308 571 320 575
rect 286 541 320 571
rect 358 541 392 575
rect 1791 554 1804 575
rect 1804 554 1825 575
rect 1791 541 1825 554
rect 1863 541 1897 575
rect 3261 541 3295 575
rect 3333 568 3334 575
rect 3334 568 3367 575
rect 3333 541 3367 568
rect 358 464 392 498
rect 430 464 452 498
rect 452 464 464 498
rect 502 464 520 498
rect 520 464 536 498
rect 574 464 588 498
rect 588 464 608 498
rect 646 464 656 498
rect 656 464 680 498
rect 718 464 724 498
rect 724 464 752 498
rect 790 464 792 498
rect 792 464 824 498
rect 862 464 894 498
rect 894 464 896 498
rect 934 464 962 498
rect 962 464 968 498
rect 1006 464 1030 498
rect 1030 464 1040 498
rect 1078 464 1098 498
rect 1098 464 1112 498
rect 1150 464 1166 498
rect 1166 464 1184 498
rect 1222 464 1234 498
rect 1234 464 1256 498
rect 1294 464 1302 498
rect 1302 464 1328 498
rect 1366 464 1370 498
rect 1370 464 1400 498
rect 1438 464 1472 498
rect 1510 464 1540 498
rect 1540 464 1544 498
rect 1582 464 1608 498
rect 1608 464 1616 498
rect 1654 464 1676 498
rect 1676 464 1688 498
rect 1726 464 1744 498
rect 1744 464 1760 498
rect 1888 464 1922 498
rect 1960 464 1982 498
rect 1982 464 1994 498
rect 2032 464 2050 498
rect 2050 464 2066 498
rect 2104 464 2118 498
rect 2118 464 2138 498
rect 2176 464 2186 498
rect 2186 464 2210 498
rect 2248 464 2254 498
rect 2254 464 2282 498
rect 2320 464 2322 498
rect 2322 464 2354 498
rect 2392 464 2424 498
rect 2424 464 2426 498
rect 2464 464 2492 498
rect 2492 464 2498 498
rect 2536 464 2560 498
rect 2560 464 2570 498
rect 2608 464 2628 498
rect 2628 464 2642 498
rect 2680 464 2696 498
rect 2696 464 2714 498
rect 2752 464 2764 498
rect 2764 464 2786 498
rect 2824 464 2832 498
rect 2832 464 2858 498
rect 2896 464 2900 498
rect 2900 464 2930 498
rect 2968 464 3002 498
rect 3040 464 3070 498
rect 3070 464 3074 498
rect 3112 464 3138 498
rect 3138 464 3146 498
rect 3184 464 3206 498
rect 3206 464 3218 498
rect 3256 464 3274 498
rect 3274 464 3290 498
rect 358 308 392 342
rect 430 308 452 342
rect 452 308 464 342
rect 502 308 520 342
rect 520 308 536 342
rect 574 308 588 342
rect 588 308 608 342
rect 646 308 656 342
rect 656 308 680 342
rect 718 308 724 342
rect 724 308 752 342
rect 790 308 792 342
rect 792 308 824 342
rect 862 308 894 342
rect 894 308 896 342
rect 934 308 962 342
rect 962 308 968 342
rect 1006 308 1030 342
rect 1030 308 1040 342
rect 1078 308 1098 342
rect 1098 308 1112 342
rect 1150 308 1166 342
rect 1166 308 1184 342
rect 1222 308 1234 342
rect 1234 308 1256 342
rect 1294 308 1302 342
rect 1302 308 1328 342
rect 1366 308 1370 342
rect 1370 308 1400 342
rect 1438 308 1472 342
rect 1510 308 1540 342
rect 1540 308 1544 342
rect 1582 308 1608 342
rect 1608 308 1616 342
rect 1654 308 1676 342
rect 1676 308 1688 342
rect 1726 308 1744 342
rect 1744 308 1760 342
rect 1888 308 1922 342
rect 1960 308 1982 342
rect 1982 308 1994 342
rect 2032 308 2050 342
rect 2050 308 2066 342
rect 2104 308 2118 342
rect 2118 308 2138 342
rect 2176 308 2186 342
rect 2186 308 2210 342
rect 2248 308 2254 342
rect 2254 308 2282 342
rect 2320 308 2322 342
rect 2322 308 2354 342
rect 2392 308 2424 342
rect 2424 308 2426 342
rect 2464 308 2492 342
rect 2492 308 2498 342
rect 2536 308 2560 342
rect 2560 308 2570 342
rect 2608 308 2628 342
rect 2628 308 2642 342
rect 2680 308 2696 342
rect 2696 308 2714 342
rect 2752 308 2764 342
rect 2764 308 2786 342
rect 2824 308 2832 342
rect 2832 308 2858 342
rect 2896 308 2900 342
rect 2900 308 2930 342
rect 2968 308 3002 342
rect 3040 308 3070 342
rect 3070 308 3074 342
rect 3112 308 3138 342
rect 3138 308 3146 342
rect 3184 308 3206 342
rect 3206 308 3218 342
rect 3256 308 3274 342
rect 3274 308 3290 342
rect 3450 698 3484 732
rect 3450 626 3484 660
rect 3450 554 3484 588
rect 3450 482 3484 516
rect 3450 410 3484 444
rect 3450 338 3484 372
rect 3450 266 3484 300
rect 188 192 222 196
rect 3450 194 3484 228
rect 188 128 222 154
rect 358 152 392 186
rect 430 152 452 186
rect 452 152 464 186
rect 502 152 520 186
rect 520 152 536 186
rect 574 152 588 186
rect 588 152 608 186
rect 646 152 656 186
rect 656 152 680 186
rect 718 152 724 186
rect 724 152 752 186
rect 790 152 792 186
rect 792 152 824 186
rect 862 152 894 186
rect 894 152 896 186
rect 934 152 962 186
rect 962 152 968 186
rect 1006 152 1030 186
rect 1030 152 1040 186
rect 1078 152 1098 186
rect 1098 152 1112 186
rect 1150 152 1166 186
rect 1166 152 1184 186
rect 1222 152 1234 186
rect 1234 152 1256 186
rect 1294 152 1302 186
rect 1302 152 1328 186
rect 1366 152 1370 186
rect 1370 152 1400 186
rect 1438 152 1472 186
rect 1510 152 1540 186
rect 1540 152 1544 186
rect 1582 152 1608 186
rect 1608 152 1616 186
rect 1654 152 1676 186
rect 1676 152 1688 186
rect 1726 152 1744 186
rect 1744 152 1760 186
rect 1888 152 1922 186
rect 1960 152 1982 186
rect 1982 152 1994 186
rect 2032 152 2050 186
rect 2050 152 2066 186
rect 2104 152 2118 186
rect 2118 152 2138 186
rect 2176 152 2186 186
rect 2186 152 2210 186
rect 2248 152 2254 186
rect 2254 152 2282 186
rect 2320 152 2322 186
rect 2322 152 2354 186
rect 2392 152 2424 186
rect 2424 152 2426 186
rect 2464 152 2492 186
rect 2492 152 2498 186
rect 2536 152 2560 186
rect 2560 152 2570 186
rect 2608 152 2628 186
rect 2628 152 2642 186
rect 2680 152 2696 186
rect 2696 152 2714 186
rect 2752 152 2764 186
rect 2764 152 2786 186
rect 2824 152 2832 186
rect 2832 152 2858 186
rect 2896 152 2900 186
rect 2900 152 2930 186
rect 2968 152 3002 186
rect 3040 152 3070 186
rect 3070 152 3074 186
rect 3112 152 3138 186
rect 3138 152 3146 186
rect 3184 152 3206 186
rect 3206 152 3218 186
rect 3256 152 3274 186
rect 3274 152 3290 186
rect 188 120 222 128
rect 188 60 222 82
rect 3450 121 3484 155
rect 188 48 222 60
rect 322 36 354 70
rect 354 36 356 70
rect 394 36 422 70
rect 422 36 428 70
rect 466 36 490 70
rect 490 36 500 70
rect 538 36 558 70
rect 558 36 572 70
rect 610 36 626 70
rect 626 36 644 70
rect 682 36 694 70
rect 694 36 716 70
rect 754 36 762 70
rect 762 36 788 70
rect 826 36 830 70
rect 830 36 860 70
rect 898 36 932 70
rect 970 36 1000 70
rect 1000 36 1004 70
rect 1042 36 1068 70
rect 1068 36 1076 70
rect 1114 36 1136 70
rect 1136 36 1148 70
rect 1186 36 1204 70
rect 1204 36 1220 70
rect 1258 36 1272 70
rect 1272 36 1292 70
rect 1330 36 1340 70
rect 1340 36 1364 70
rect 1402 36 1408 70
rect 1408 36 1436 70
rect 1474 36 1476 70
rect 1476 36 1508 70
rect 1546 36 1578 70
rect 1578 36 1580 70
rect 1618 36 1646 70
rect 1646 36 1652 70
rect 1690 36 1714 70
rect 1714 36 1724 70
rect 1762 36 1782 70
rect 1782 36 1796 70
rect 1834 36 1850 70
rect 1850 36 1868 70
rect 1906 36 1918 70
rect 1918 36 1940 70
rect 1978 36 1986 70
rect 1986 36 2012 70
rect 2050 36 2054 70
rect 2054 36 2084 70
rect 2122 36 2156 70
rect 2194 36 2224 70
rect 2224 36 2228 70
rect 2266 36 2292 70
rect 2292 36 2300 70
rect 2338 36 2360 70
rect 2360 36 2372 70
rect 2410 36 2428 70
rect 2428 36 2444 70
rect 2482 36 2496 70
rect 2496 36 2516 70
rect 2554 36 2564 70
rect 2564 36 2588 70
rect 2626 36 2632 70
rect 2632 36 2660 70
rect 2698 36 2700 70
rect 2700 36 2732 70
rect 2770 36 2802 70
rect 2802 36 2804 70
rect 2842 36 2870 70
rect 2870 36 2876 70
rect 2914 36 2938 70
rect 2938 36 2948 70
rect 2986 36 3006 70
rect 3006 36 3020 70
rect 3058 36 3074 70
rect 3074 36 3092 70
rect 3130 36 3142 70
rect 3142 36 3164 70
rect 3202 36 3210 70
rect 3210 36 3236 70
rect 3274 36 3278 70
rect 3278 36 3308 70
rect 3346 36 3380 70
rect 3450 48 3484 82
rect -10 0 24 20
rect -10 -14 24 0
rect 1180 -116 1214 -104
rect 1254 -116 1288 -104
rect 1328 -116 1362 -104
rect 1402 -116 1436 -104
rect 2 -150 14 -116
rect 14 -150 36 -116
rect 74 -150 82 -116
rect 82 -150 108 -116
rect 146 -150 150 -116
rect 150 -150 180 -116
rect 218 -150 252 -116
rect 290 -150 320 -116
rect 320 -150 324 -116
rect 362 -150 388 -116
rect 388 -150 396 -116
rect 434 -150 456 -116
rect 456 -150 468 -116
rect 506 -150 524 -116
rect 524 -150 540 -116
rect 578 -150 592 -116
rect 592 -150 612 -116
rect 650 -150 660 -116
rect 660 -150 684 -116
rect 722 -150 728 -116
rect 728 -150 756 -116
rect 794 -150 796 -116
rect 796 -150 828 -116
rect 866 -150 898 -116
rect 898 -150 900 -116
rect 938 -150 966 -116
rect 966 -150 972 -116
rect 1010 -150 1034 -116
rect 1034 -150 1044 -116
rect 1082 -150 1102 -116
rect 1102 -150 1116 -116
rect 1180 -138 1204 -116
rect 1204 -138 1214 -116
rect 1254 -138 1272 -116
rect 1272 -138 1288 -116
rect 1328 -138 1340 -116
rect 1340 -138 1362 -116
rect 1402 -138 1408 -116
rect 1408 -138 1436 -116
rect 1476 -138 1510 -104
rect 1550 -116 1584 -104
rect 1624 -116 1658 -104
rect 1698 -116 1732 -104
rect 1772 -116 1806 -104
rect 1846 -116 1880 -104
rect 1920 -116 1954 -104
rect 1994 -116 2028 -104
rect 2068 -116 2102 -104
rect 2142 -116 2176 -104
rect 2216 -116 2250 -104
rect 2290 -116 2324 -104
rect 2364 -116 2398 -104
rect 2438 -116 2472 -104
rect 2512 -116 2546 -104
rect 2586 -116 2620 -104
rect 2660 -116 2694 -104
rect 2734 -116 2768 -104
rect 2808 -116 2842 -104
rect 2882 -116 2916 -104
rect 2956 -116 2990 -104
rect 3030 -116 3064 -104
rect 3104 -116 3138 -104
rect 3178 -116 3212 -104
rect 3252 -116 3286 -104
rect 3326 -116 3360 -104
rect 1550 -138 1578 -116
rect 1578 -138 1584 -116
rect 1624 -138 1646 -116
rect 1646 -138 1658 -116
rect 1698 -138 1714 -116
rect 1714 -138 1732 -116
rect 1772 -138 1782 -116
rect 1782 -138 1806 -116
rect 1846 -138 1850 -116
rect 1850 -138 1880 -116
rect 1920 -138 1952 -116
rect 1952 -138 1954 -116
rect 1994 -138 2020 -116
rect 2020 -138 2028 -116
rect 2068 -138 2088 -116
rect 2088 -138 2102 -116
rect 2142 -138 2156 -116
rect 2156 -138 2176 -116
rect 2216 -138 2224 -116
rect 2224 -138 2250 -116
rect 2290 -138 2292 -116
rect 2292 -138 2324 -116
rect 2364 -138 2394 -116
rect 2394 -138 2398 -116
rect 2438 -138 2462 -116
rect 2462 -138 2472 -116
rect 2512 -138 2530 -116
rect 2530 -138 2546 -116
rect 2586 -138 2598 -116
rect 2598 -138 2620 -116
rect 2660 -138 2666 -116
rect 2666 -138 2694 -116
rect 2734 -138 2768 -116
rect 2808 -138 2836 -116
rect 2836 -138 2842 -116
rect 2882 -138 2904 -116
rect 2904 -138 2916 -116
rect 2956 -138 2972 -116
rect 2972 -138 2990 -116
rect 3030 -138 3040 -116
rect 3040 -138 3064 -116
rect 3104 -138 3108 -116
rect 3108 -138 3138 -116
rect 3178 -138 3210 -116
rect 3210 -138 3212 -116
rect 3252 -138 3278 -116
rect 3278 -138 3286 -116
rect 3326 -138 3346 -116
rect 3346 -138 3360 -116
rect 3400 -138 3434 -104
<< metal1 >>
rect -22 1112 3467 1143
rect -22 1100 101 1112
rect -22 1066 -10 1100
rect 24 1078 101 1100
rect 135 1078 173 1112
rect 207 1078 245 1112
rect 279 1078 317 1112
rect 351 1078 389 1112
rect 423 1078 461 1112
rect 495 1078 533 1112
rect 567 1078 605 1112
rect 639 1078 677 1112
rect 711 1078 749 1112
rect 783 1078 821 1112
rect 855 1078 893 1112
rect 927 1078 965 1112
rect 999 1078 1037 1112
rect 1071 1078 1109 1112
rect 1143 1078 1181 1112
rect 1215 1078 1253 1112
rect 1287 1078 1325 1112
rect 1359 1078 1397 1112
rect 1431 1078 1469 1112
rect 1503 1078 1541 1112
rect 1575 1078 1613 1112
rect 1647 1078 1685 1112
rect 1719 1078 1757 1112
rect 1791 1078 1829 1112
rect 1863 1078 1901 1112
rect 1935 1078 1973 1112
rect 2007 1078 2045 1112
rect 2079 1078 2117 1112
rect 2151 1078 2189 1112
rect 2223 1078 2261 1112
rect 2295 1078 2333 1112
rect 2367 1078 2405 1112
rect 2439 1078 2477 1112
rect 2511 1078 2549 1112
rect 2583 1078 2621 1112
rect 2655 1078 2693 1112
rect 2727 1078 2765 1112
rect 2799 1078 2837 1112
rect 2871 1078 2909 1112
rect 2943 1078 2981 1112
rect 3015 1078 3053 1112
rect 3087 1078 3125 1112
rect 3159 1078 3197 1112
rect 3231 1078 3269 1112
rect 3303 1078 3341 1112
rect 3375 1078 3413 1112
rect 3447 1078 3467 1112
rect 24 1066 3467 1078
rect -22 1028 36 1066
rect -22 994 -10 1028
rect 24 994 36 1028
rect -22 956 36 994
rect -22 922 -10 956
rect 24 922 36 956
rect -22 884 36 922
tri 36 918 184 1066 nw
rect -22 850 -10 884
rect 24 850 36 884
rect -22 812 36 850
rect -22 778 -10 812
rect 24 778 36 812
rect -22 740 36 778
rect -22 706 -10 740
rect 24 706 36 740
rect -22 668 36 706
rect -22 634 -10 668
rect 24 634 36 668
rect -22 596 36 634
rect -22 562 -10 596
rect 24 562 36 596
rect -22 524 36 562
rect -22 490 -10 524
rect 24 490 36 524
rect -22 452 36 490
rect -22 418 -10 452
rect 24 418 36 452
rect -22 380 36 418
rect -22 346 -10 380
rect 24 346 36 380
rect -22 308 36 346
rect -22 274 -10 308
rect 24 274 36 308
rect -22 236 36 274
rect -22 202 -10 236
rect 24 202 36 236
rect -22 164 36 202
rect -22 130 -10 164
rect 24 130 36 164
rect -22 92 36 130
rect -22 58 -10 92
rect 24 58 36 92
rect -22 20 36 58
rect 176 810 3438 816
rect 176 776 358 810
rect 392 776 430 810
rect 464 776 502 810
rect 536 776 574 810
rect 608 776 646 810
rect 680 776 718 810
rect 752 776 790 810
rect 824 776 862 810
rect 896 776 934 810
rect 968 776 1006 810
rect 1040 776 1078 810
rect 1112 776 1150 810
rect 1184 776 1222 810
rect 1256 776 1294 810
rect 1328 776 1366 810
rect 1400 776 1438 810
rect 1472 776 1510 810
rect 1544 776 1582 810
rect 1616 776 1654 810
rect 1688 776 1726 810
rect 1760 776 1888 810
rect 1922 776 1960 810
rect 1994 776 2032 810
rect 2066 776 2104 810
rect 2138 776 2176 810
rect 2210 776 2248 810
rect 2282 776 2320 810
rect 2354 776 2392 810
rect 2426 776 2464 810
rect 2498 776 2536 810
rect 2570 776 2608 810
rect 2642 776 2680 810
rect 2714 776 2752 810
rect 2786 776 2824 810
rect 2858 776 2896 810
rect 2930 776 2968 810
rect 3002 776 3040 810
rect 3074 776 3112 810
rect 3146 776 3184 810
rect 3218 776 3256 810
rect 3290 805 3438 810
rect 3444 805 3490 816
rect 3290 804 3496 805
rect 3290 776 3450 804
rect 176 770 3450 776
rect 3484 770 3496 804
rect 176 730 234 770
tri 234 744 260 770 nw
tri 3379 744 3405 770 ne
rect 3405 744 3496 770
tri 3405 733 3416 744 ne
rect 3416 733 3496 744
rect 176 696 188 730
rect 222 696 234 730
rect 176 658 234 696
rect 176 624 188 658
rect 222 624 234 658
rect 176 586 234 624
rect 346 654 3302 733
tri 3416 732 3417 733 ne
rect 3417 732 3496 733
tri 3417 711 3438 732 ne
rect 346 620 358 654
rect 392 620 430 654
rect 464 620 502 654
rect 536 620 574 654
rect 608 620 646 654
rect 680 620 718 654
rect 752 620 790 654
rect 824 620 862 654
rect 896 620 934 654
rect 968 620 1006 654
rect 1040 620 1078 654
rect 1112 620 1150 654
rect 1184 620 1222 654
rect 1256 620 1294 654
rect 1328 620 1366 654
rect 1400 620 1438 654
rect 1472 620 1510 654
rect 1544 620 1582 654
rect 1616 620 1654 654
rect 1688 620 1726 654
rect 1760 620 1888 654
rect 1922 620 1960 654
rect 1994 620 2032 654
rect 2066 620 2104 654
rect 2138 620 2176 654
rect 2210 620 2248 654
rect 2282 620 2320 654
rect 2354 620 2392 654
rect 2426 620 2464 654
rect 2498 620 2536 654
rect 2570 620 2608 654
rect 2642 620 2680 654
rect 2714 620 2752 654
rect 2786 620 2824 654
rect 2858 620 2896 654
rect 2930 620 2968 654
rect 3002 620 3040 654
rect 3074 620 3112 654
rect 3146 620 3184 654
rect 3218 620 3256 654
rect 3290 620 3302 654
rect 346 614 3302 620
rect 3438 698 3450 732
rect 3484 698 3496 732
rect 3438 660 3496 698
rect 3438 626 3450 660
rect 3484 626 3496 660
rect 176 552 188 586
rect 222 552 234 586
rect 3438 588 3496 626
rect 176 516 234 552
rect 274 575 3379 581
rect 274 541 286 575
rect 320 541 358 575
rect 392 541 1791 575
rect 1825 541 1863 575
rect 1897 541 3261 575
rect 3295 541 3333 575
rect 3367 541 3379 575
rect 3438 554 3450 588
rect 3484 554 3496 588
rect 274 535 3379 541
tri 3422 535 3438 551 se
rect 3438 535 3496 554
tri 3420 533 3422 535 se
rect 3422 533 3496 535
tri 234 516 251 533 sw
tri 3403 516 3420 533 se
rect 3420 516 3496 533
rect 176 514 251 516
rect 176 480 188 514
rect 222 504 251 514
tri 251 504 263 516 sw
tri 3391 504 3403 516 se
rect 3403 504 3450 516
rect 222 498 3450 504
rect 222 480 358 498
rect 176 464 358 480
rect 392 464 430 498
rect 464 464 502 498
rect 536 464 574 498
rect 608 464 646 498
rect 680 464 718 498
rect 752 464 790 498
rect 824 464 862 498
rect 896 464 934 498
rect 968 464 1006 498
rect 1040 464 1078 498
rect 1112 464 1150 498
rect 1184 464 1222 498
rect 1256 464 1294 498
rect 1328 464 1366 498
rect 1400 464 1438 498
rect 1472 464 1510 498
rect 1544 464 1582 498
rect 1616 464 1654 498
rect 1688 464 1726 498
rect 1760 464 1888 498
rect 1922 464 1960 498
rect 1994 464 2032 498
rect 2066 464 2104 498
rect 2138 464 2176 498
rect 2210 464 2248 498
rect 2282 464 2320 498
rect 2354 464 2392 498
rect 2426 464 2464 498
rect 2498 464 2536 498
rect 2570 464 2608 498
rect 2642 464 2680 498
rect 2714 464 2752 498
rect 2786 464 2824 498
rect 2858 464 2896 498
rect 2930 464 2968 498
rect 3002 464 3040 498
rect 3074 464 3112 498
rect 3146 464 3184 498
rect 3218 464 3256 498
rect 3290 482 3450 498
rect 3484 482 3496 516
rect 3290 464 3496 482
rect 176 444 3496 464
rect 176 442 3450 444
rect 176 408 188 442
rect 222 410 3450 442
rect 3484 410 3496 444
rect 222 408 3496 410
rect 176 385 3496 408
rect 176 372 252 385
tri 252 372 265 385 nw
tri 3388 372 3401 385 ne
rect 3401 372 3496 385
rect 176 370 234 372
rect 176 336 188 370
rect 222 336 234 370
tri 234 354 252 372 nw
tri 3401 354 3419 372 ne
rect 3419 354 3450 372
tri 3419 348 3425 354 ne
rect 3425 348 3450 354
rect 176 298 234 336
rect 176 264 188 298
rect 222 264 234 298
rect 176 228 234 264
rect 346 342 3302 348
rect 346 308 358 342
rect 392 308 430 342
rect 464 308 502 342
rect 536 308 574 342
rect 608 308 646 342
rect 680 308 718 342
rect 752 308 790 342
rect 824 308 862 342
rect 896 308 934 342
rect 968 308 1006 342
rect 1040 308 1078 342
rect 1112 308 1150 342
rect 1184 308 1222 342
rect 1256 308 1294 342
rect 1328 308 1366 342
rect 1400 308 1438 342
rect 1472 308 1510 342
rect 1544 308 1582 342
rect 1616 308 1654 342
rect 1688 308 1726 342
rect 1760 308 1888 342
rect 1922 308 1960 342
rect 1994 308 2032 342
rect 2066 308 2104 342
rect 2138 308 2176 342
rect 2210 308 2248 342
rect 2282 308 2320 342
rect 2354 308 2392 342
rect 2426 308 2464 342
rect 2498 308 2536 342
rect 2570 308 2608 342
rect 2642 308 2680 342
rect 2714 308 2752 342
rect 2786 308 2824 342
rect 2858 308 2896 342
rect 2930 308 2968 342
rect 3002 308 3040 342
rect 3074 308 3112 342
rect 3146 308 3184 342
rect 3218 308 3256 342
rect 3290 308 3302 342
tri 3425 338 3435 348 ne
rect 3435 338 3450 348
rect 3484 338 3496 372
tri 3435 335 3438 338 ne
rect 346 229 3302 308
rect 3438 300 3496 338
rect 3438 266 3450 300
rect 3484 266 3496 300
tri 3414 229 3438 253 se
rect 3438 229 3496 266
tri 234 228 235 229 sw
tri 3413 228 3414 229 se
rect 3414 228 3496 229
rect 176 226 235 228
rect 176 192 188 226
rect 222 194 235 226
tri 235 194 269 228 sw
tri 3379 194 3413 228 se
rect 3413 194 3450 228
rect 3484 194 3496 228
rect 222 192 269 194
tri 269 192 271 194 sw
tri 3377 192 3379 194 se
rect 3379 192 3496 194
rect 176 186 3496 192
rect 176 154 358 186
rect 176 120 188 154
rect 222 152 358 154
rect 392 152 430 186
rect 464 152 502 186
rect 536 152 574 186
rect 608 152 646 186
rect 680 152 718 186
rect 752 152 790 186
rect 824 152 862 186
rect 896 152 934 186
rect 968 152 1006 186
rect 1040 152 1078 186
rect 1112 152 1150 186
rect 1184 152 1222 186
rect 1256 152 1294 186
rect 1328 152 1366 186
rect 1400 152 1438 186
rect 1472 152 1510 186
rect 1544 152 1582 186
rect 1616 152 1654 186
rect 1688 152 1726 186
rect 1760 152 1888 186
rect 1922 152 1960 186
rect 1994 152 2032 186
rect 2066 152 2104 186
rect 2138 152 2176 186
rect 2210 152 2248 186
rect 2282 152 2320 186
rect 2354 152 2392 186
rect 2426 152 2464 186
rect 2498 152 2536 186
rect 2570 152 2608 186
rect 2642 152 2680 186
rect 2714 152 2752 186
rect 2786 152 2824 186
rect 2858 152 2896 186
rect 2930 152 2968 186
rect 3002 152 3040 186
rect 3074 152 3112 186
rect 3146 152 3184 186
rect 3218 152 3256 186
rect 3290 155 3496 186
rect 3290 152 3450 155
rect 222 121 3450 152
rect 3484 121 3496 155
rect 222 120 3496 121
rect 176 98 3496 120
rect 176 82 3519 98
rect 176 48 188 82
rect 222 70 3450 82
rect 222 48 322 70
rect 176 36 322 48
rect 356 36 394 70
rect 428 36 466 70
rect 500 36 538 70
rect 572 36 610 70
rect 644 36 682 70
rect 716 36 754 70
rect 788 36 826 70
rect 860 36 898 70
rect 932 36 970 70
rect 1004 36 1042 70
rect 1076 36 1114 70
rect 1148 36 1186 70
rect 1220 36 1258 70
rect 1292 36 1330 70
rect 1364 36 1402 70
rect 1436 36 1474 70
rect 1508 36 1546 70
rect 1580 36 1618 70
rect 1652 36 1690 70
rect 1724 36 1762 70
rect 1796 36 1834 70
rect 1868 36 1906 70
rect 1940 36 1978 70
rect 2012 36 2050 70
rect 2084 36 2122 70
rect 2156 36 2194 70
rect 2228 36 2266 70
rect 2300 36 2338 70
rect 2372 36 2410 70
rect 2444 36 2482 70
rect 2516 36 2554 70
rect 2588 36 2626 70
rect 2660 36 2698 70
rect 2732 36 2770 70
rect 2804 36 2842 70
rect 2876 36 2914 70
rect 2948 36 2986 70
rect 3020 36 3058 70
rect 3092 36 3130 70
rect 3164 36 3202 70
rect 3236 36 3274 70
rect 3308 36 3346 70
rect 3380 48 3450 70
rect 3484 48 3519 82
rect 3380 36 3519 48
rect 176 24 3519 36
rect -22 -14 -10 20
rect 24 -14 36 20
rect -22 -104 36 -14
tri 36 -104 102 -38 sw
tri 1162 -104 1168 -98 se
rect 1168 -104 3488 -98
rect -22 -116 1180 -104
rect -22 -150 2 -116
rect 36 -150 74 -116
rect 108 -150 146 -116
rect 180 -150 218 -116
rect 252 -150 290 -116
rect 324 -150 362 -116
rect 396 -150 434 -116
rect 468 -150 506 -116
rect 540 -150 578 -116
rect 612 -150 650 -116
rect 684 -150 722 -116
rect 756 -150 794 -116
rect 828 -150 866 -116
rect 900 -150 938 -116
rect 972 -150 1010 -116
rect 1044 -150 1082 -116
rect 1116 -138 1180 -116
rect 1214 -138 1254 -104
rect 1288 -138 1328 -104
rect 1362 -138 1402 -104
rect 1436 -138 1476 -104
rect 1510 -138 1550 -104
rect 1584 -138 1624 -104
rect 1658 -138 1698 -104
rect 1732 -138 1772 -104
rect 1806 -138 1846 -104
rect 1880 -138 1920 -104
rect 1954 -138 1994 -104
rect 2028 -138 2068 -104
rect 2102 -138 2142 -104
rect 2176 -138 2216 -104
rect 2250 -138 2290 -104
rect 2324 -138 2364 -104
rect 2398 -138 2438 -104
rect 2472 -138 2512 -104
rect 2546 -138 2586 -104
rect 2620 -138 2660 -104
rect 2694 -138 2734 -104
rect 2768 -138 2808 -104
rect 2842 -138 2882 -104
rect 2916 -138 2956 -104
rect 2990 -138 3030 -104
rect 3064 -138 3104 -104
rect 3138 -138 3178 -104
rect 3212 -138 3252 -104
rect 3286 -138 3326 -104
rect 3360 -138 3400 -104
rect 3434 -138 3488 -104
rect 1116 -144 3488 -138
rect 1116 -150 1168 -144
rect -22 -162 1168 -150
tri 1168 -162 1186 -144 nw
use sky130_fd_pr__pfet_01v8__example_55959141808654  sky130_fd_pr__pfet_01v8__example_55959141808654_0
timestamp 1645210163
transform 0 -1 1756 1 0 197
box -28 0 596 697
use sky130_fd_pr__pfet_01v8__example_55959141808654  sky130_fd_pr__pfet_01v8__example_55959141808654_1
timestamp 1645210163
transform 0 -1 3286 1 0 197
box -28 0 596 697
<< labels >>
flabel metal1 s 274 535 320 581 7 FreeSans 200 180 0 0 PU_H_N
port 1 nsew
flabel metal1 s 347 648 393 700 7 FreeSans 200 180 0 0 PAD
port 2 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 5685224
string GDS_START 5653446
<< end >>
