// File: nmos_top_trim1.spi.NMOS_TOP_TRIM1.pxi
// Created: Tue Oct 15 15:58:57 2024
// 
simulator lang=spectre
cc_1 ( noxref_1 noxref_2 ) capacitor c=0.0463663f //x=0.43 //y=0.54 //x2=0 \
 //y2=0
cc_2 ( noxref_1 noxref_3 ) capacitor c=0.016062f //x=0.43 //y=0.54 //x2=0.62 \
 //y2=0.965
cc_3 ( noxref_2 noxref_3 ) capacitor c=0.0805399f //x=0 //y=0 //x2=0.62 \
 //y2=0.965
