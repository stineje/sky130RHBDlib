* SPICE3 file created from TMRDFFRNQNX1.ext - technology: sky130A

.subckt TMRDFFRNQNX1 QN D CLK RN VDD GND
M1000 a_5779_989.t1 RN.t0 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_9009_1050.t4 a_9331_989.t5 VDD.t39 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_5457_1050.t1 CLK.t0 VDD.t95 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 GND a_9331_989.t7 a_16318_101.t0 nshort w=-1.605u l=1.765u
+  ad=3.7611p pd=32.97u as=0p ps=0u
M1004 a_15757_1051.t4 a_9331_989.t6 a_16421_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD.t97 a_14511_989.t5 a_14189_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VDD.t5 RN.t1 a_147_187.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 GND a_5457_1050.t7 a_8823_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t32 a_147_187.t8 a_4151_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VDD.t28 a_5327_187.t7 a_7321_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_16421_1051.t1 a_4151_989.t5 QN.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_14511_989.t4 a_14189_1050.t7 VDD.t83 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_12501_1050.t1 a_10959_989.t8 VDD.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 GND a_5457_1050.t8 a_6233_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t8 RN.t3 a_10959_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 QN a_14511_989.t8 a_16984_101.t0 nshort w=-1.83u l=2.06u
+  ad=0.5373p pd=4.72u as=0p ps=0u
M1016 a_5457_1050.t3 a_5779_989.t7 VDD.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_5327_187.t3 RN.t5 VDD.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 GND a_9009_1050.t8 a_9806_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 VDD.t64 a_147_187.t9 a_277_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_15757_1051.t7 a_4151_989.t6 a_16421_1051.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t96 a_10507_187.t9 a_10637_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t3 a_12501_1050.t5 a_10507_187.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 GND a_5779_989.t9 a_7216_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 VDD.t17 RN.t6 a_10507_187.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 GND a_147_187.t10 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_14189_1050.t5 a_10637_1050.t7 VDD.t40 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 GND a_7321_1050.t5 a_7861_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_10959_989.t6 a_10637_1050.t8 VDD.t91 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_599_989.t6 D.t1 VDD.t49 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_16421_1051.t0 a_14511_989.t7 QN.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 GND a_5327_187.t9 a_5271_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_5327_187.t1 CLK.t3 VDD.t86 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 VDD.t74 a_599_989.t8 a_2141_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_9331_989.t4 a_9009_1050.t7 VDD.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 VDD.t78 CLK.t4 a_277_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 VDD.t94 a_5457_1050.t9 a_5779_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VDD.t93 a_5457_1050.t10 a_9009_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VDD.t35 a_277_1050.t7 a_3829_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VDD.t36 CLK.t5 a_10507_187.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 VDD.t11 RN.t8 a_5779_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VDD.t38 a_9331_989.t8 a_9009_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VDD.t65 CLK.t6 a_10637_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_9331_989.t2 a_5327_187.t8 VDD.t54 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_14189_1050.t1 RN.t9 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_10959_989.t3 D.t2 VDD.t77 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_599_989.t1 RN.t10 VDD.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_3829_1050.t5 a_4151_989.t7 VDD.t68 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_10637_1050.t5 a_10507_187.t10 VDD.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 VDD.t0 a_14511_989.t9 a_15757_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_147_187.t5 CLK.t7 VDD.t88 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 GND a_12501_1050.t6 a_13041_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1052 QN a_4151_989.t10 a_16318_101.t0 nshort w=-1.235u l=1.535u
+  ad=0p pd=0u as=0p ps=0u
M1053 GND a_277_1050.t8 a_3643_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_4151_989.t4 a_3829_1050.t7 VDD.t33 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_9009_1050.t5 a_5457_1050.t11 VDD.t85 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_15757_1051.t2 a_9331_989.t9 VDD.t72 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 VDD.t82 a_14189_1050.t8 a_14511_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 VDD.t25 a_10959_989.t9 a_12501_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 VDD.t52 a_147_187.t11 a_2141_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 VDD.t45 a_599_989.t9 a_277_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 VDD.t20 RN.t12 a_9009_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 VDD.t30 D.t4 a_5779_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 VDD.t70 a_2141_1050.t5 a_147_187.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 VDD.t90 a_5327_187.t11 a_5457_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 VDD.t51 a_7321_1050.t6 a_5327_187.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 GND a_3829_1050.t8 a_4626_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_14189_1050.t2 a_14511_989.t11 VDD.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_10959_989.t5 RN.t13 VDD.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 GND a_599_989.t10 a_2036_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_147_187.t0 RN.t14 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 GND a_10637_1050.t9 a_14003_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1072 GND a_2141_1050.t6 a_2681_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1073 a_4151_989.t1 a_147_187.t12 VDD.t53 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 a_7321_1050.t2 a_5327_187.t12 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 QN.t5 a_4151_989.t9 a_16421_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 VDD.t24 a_10959_989.t10 a_10637_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 a_15757_1051.t6 a_14511_989.t12 VDD.t58 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 VDD.t79 a_10507_187.t12 a_14511_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VDD.t59 a_10507_187.t13 a_12501_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 GND a_9331_989.t10 a_15652_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1081 GND a_14189_1050.t9 a_14986_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1082 a_277_1050.t2 a_147_187.t13 VDD.t46 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_16421_1051.t4 a_4151_989.t11 a_15757_1051.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 VDD.t41 a_9009_1050.t9 a_9331_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_10507_187.t6 a_12501_1050.t7 VDD.t55 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_10507_187.t3 RN.t15 VDD.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 a_10637_1050.t2 a_10959_989.t11 VDD.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_7321_1050.t1 a_5779_989.t10 VDD.t69 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 VDD.t71 a_277_1050.t9 a_599_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 QN.t3 a_14511_989.t13 a_16421_1051.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 VDD.t89 a_4151_989.t12 a_3829_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 VDD.t13 RN.t17 a_599_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 GND a_277_1050.t11 a_1053_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_2141_1050.t3 a_599_989.t11 VDD.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 VDD.t43 a_5779_989.t11 a_5457_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 VDD.t14 RN.t19 a_5327_187.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_16421_1051.t2 a_9331_989.t11 a_15757_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_277_1050.t0 CLK.t11 VDD.t26 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 a_3829_1050.t2 a_277_1050.t10 VDD.t92 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_5779_989.t5 a_5457_1050.t12 VDD.t80 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 GND a_4151_989.t13 a_16984_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_10507_187.t0 CLK.t12 VDD.t81 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_10637_1050.t0 CLK.t13 VDD.t76 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 VDD.t63 a_10637_1050.t10 a_14189_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 VDD.t61 a_10637_1050.t11 a_10959_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 GND a_10637_1050.t12 a_11413_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1107 VDD.t48 D.t5 a_599_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 VDD.t21 RN.t21 a_3829_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 a_599_989.t3 a_277_1050.t12 VDD.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 VDD.t99 CLK.t15 a_5327_187.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 VDD.t87 CLK.t16 a_5457_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1112 a_2141_1050.t0 a_147_187.t14 VDD.t47 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 GND a_10959_989.t7 a_12396_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1114 a_277_1050.t6 a_599_989.t12 VDD.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 a_3829_1050.t0 RN.t23 VDD.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 a_5779_989.t4 D.t6 VDD.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_9009_1050.t0 RN.t24 VDD.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_5457_1050.t5 a_5327_187.t14 VDD.t50 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_5327_187.t6 a_7321_1050.t7 VDD.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 VDD.t67 a_5327_187.t15 a_9331_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 a_147_187.t6 a_2141_1050.t7 VDD.t98 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 GND a_10507_187.t7 a_10451_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1123 VDD.t19 RN.t25 a_14189_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1124 VDD.t37 D.t7 a_10959_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1125 QN a_14511_989.t6 a_15652_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1126 VDD.t57 CLK.t17 a_147_187.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1127 VDD.t1 a_3829_1050.t9 a_4151_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1128 VDD.t44 a_5779_989.t12 a_7321_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1129 VDD.t42 a_9331_989.t13 a_15757_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1130 a_14511_989.t0 a_10507_187.t14 VDD.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1131 a_12501_1050.t2 a_10507_187.t15 VDD.t60 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD CLK 1.71fF
C1 VDD D 0.15fF
C2 CLK D 0.45fF
C3 VDD RN 0.50fF
C4 CLK RN 1.13fF
C5 VDD QN 0.29fF
C6 D RN 12.60fF
R0 a_10959_989.n5 a_10959_989.t9 480.392
R1 a_10959_989.n7 a_10959_989.t11 454.685
R2 a_10959_989.n7 a_10959_989.t10 428.979
R3 a_10959_989.n5 a_10959_989.t8 403.272
R4 a_10959_989.n6 a_10959_989.t7 283.48
R5 a_10959_989.n8 a_10959_989.t12 237.959
R6 a_10959_989.n12 a_10959_989.n10 219.626
R7 a_10959_989.n10 a_10959_989.n4 170.799
R8 a_10959_989.n8 a_10959_989.n7 98.447
R9 a_10959_989.n6 a_10959_989.n5 98.447
R10 a_10959_989.n9 a_10959_989.n8 80.035
R11 a_10959_989.n3 a_10959_989.n2 79.232
R12 a_10959_989.n9 a_10959_989.n6 77.315
R13 a_10959_989.n10 a_10959_989.n9 76
R14 a_10959_989.n4 a_10959_989.n3 63.152
R15 a_10959_989.n4 a_10959_989.n0 16.08
R16 a_10959_989.n3 a_10959_989.n1 16.08
R17 a_10959_989.n12 a_10959_989.n11 15.218
R18 a_10959_989.n0 a_10959_989.t4 14.282
R19 a_10959_989.n0 a_10959_989.t5 14.282
R20 a_10959_989.n1 a_10959_989.t0 14.282
R21 a_10959_989.n1 a_10959_989.t3 14.282
R22 a_10959_989.n2 a_10959_989.t1 14.282
R23 a_10959_989.n2 a_10959_989.t6 14.282
R24 a_10959_989.n13 a_10959_989.n12 12.014
R25 a_12396_101.n10 a_12396_101.n9 93.333
R26 a_12396_101.n2 a_12396_101.n1 41.622
R27 a_12396_101.n13 a_12396_101.n12 26.667
R28 a_12396_101.n6 a_12396_101.n5 24.977
R29 a_12396_101.t0 a_12396_101.n2 21.209
R30 a_12396_101.t0 a_12396_101.n3 11.595
R31 a_12396_101.t1 a_12396_101.n8 8.137
R32 a_12396_101.t0 a_12396_101.n0 6.109
R33 a_12396_101.t1 a_12396_101.n7 4.864
R34 a_12396_101.t0 a_12396_101.n4 3.871
R35 a_12396_101.t0 a_12396_101.n13 2.535
R36 a_12396_101.n13 a_12396_101.t1 1.145
R37 a_12396_101.n7 a_12396_101.n6 1.13
R38 a_12396_101.t1 a_12396_101.n11 0.804
R39 a_12396_101.n11 a_12396_101.n10 0.136
R40 GND.n26 GND.n24 219.745
R41 GND.n56 GND.n54 219.745
R42 GND.n432 GND.n431 219.745
R43 GND.n474 GND.n472 219.745
R44 GND.n507 GND.n505 219.745
R45 GND.n549 GND.n547 219.745
R46 GND.n591 GND.n589 219.745
R47 GND.n621 GND.n619 219.745
R48 GND.n663 GND.n661 219.745
R49 GND.n705 GND.n703 219.745
R50 GND.n735 GND.n733 219.745
R51 GND.n387 GND.n385 219.745
R52 GND.n347 GND.n345 219.745
R53 GND.n317 GND.n315 219.745
R54 GND.n275 GND.n273 219.745
R55 GND.n230 GND.n228 219.745
R56 GND.n200 GND.n198 219.745
R57 GND.n158 GND.n156 219.745
R58 GND.n116 GND.n114 219.745
R59 GND.n86 GND.n85 219.745
R60 GND.n147 GND.n146 85.559
R61 GND.n189 GND.n188 85.559
R62 GND.n306 GND.n305 85.559
R63 GND.n378 GND.n377 85.559
R64 GND.n744 GND.n743 85.559
R65 GND.n672 GND.n671 85.559
R66 GND.n630 GND.n629 85.559
R67 GND.n558 GND.n557 85.559
R68 GND.n516 GND.n515 85.559
R69 GND.n441 GND.n440 85.559
R70 GND.n399 GND.n398 85.559
R71 GND.n26 GND.n25 85.529
R72 GND.n56 GND.n55 85.529
R73 GND.n432 GND.n430 85.529
R74 GND.n474 GND.n473 85.529
R75 GND.n507 GND.n506 85.529
R76 GND.n549 GND.n548 85.529
R77 GND.n591 GND.n590 85.529
R78 GND.n621 GND.n620 85.529
R79 GND.n663 GND.n662 85.529
R80 GND.n705 GND.n704 85.529
R81 GND.n735 GND.n734 85.529
R82 GND.n387 GND.n386 85.529
R83 GND.n347 GND.n346 85.529
R84 GND.n317 GND.n316 85.529
R85 GND.n275 GND.n274 85.529
R86 GND.n230 GND.n229 85.529
R87 GND.n200 GND.n199 85.529
R88 GND.n158 GND.n157 85.529
R89 GND.n116 GND.n115 85.529
R90 GND.n86 GND.n84 85.529
R91 GND.n44 GND.n43 84.842
R92 GND.n74 GND.n73 84.842
R93 GND.n104 GND.n103 84.842
R94 GND.n218 GND.n217 84.842
R95 GND.n335 GND.n334 84.842
R96 GND.n713 GND.n712 84.842
R97 GND.n599 GND.n598 84.842
R98 GND.n14 GND.n13 84.842
R99 GND.n393 GND.n392 76
R100 GND.n39 GND.n38 76
R101 GND.n42 GND.n41 76
R102 GND.n47 GND.n46 76
R103 GND.n50 GND.n49 76
R104 GND.n53 GND.n52 76
R105 GND.n60 GND.n59 76
R106 GND.n63 GND.n62 76
R107 GND.n66 GND.n65 76
R108 GND.n69 GND.n68 76
R109 GND.n72 GND.n71 76
R110 GND.n77 GND.n76 76
R111 GND.n80 GND.n79 76
R112 GND.n83 GND.n82 76
R113 GND.n90 GND.n89 76
R114 GND.n93 GND.n92 76
R115 GND.n96 GND.n95 76
R116 GND.n99 GND.n98 76
R117 GND.n102 GND.n101 76
R118 GND.n107 GND.n106 76
R119 GND.n110 GND.n109 76
R120 GND.n113 GND.n112 76
R121 GND.n120 GND.n119 76
R122 GND.n123 GND.n122 76
R123 GND.n126 GND.n125 76
R124 GND.n129 GND.n128 76
R125 GND.n132 GND.n131 76
R126 GND.n135 GND.n134 76
R127 GND.n138 GND.n137 76
R128 GND.n141 GND.n140 76
R129 GND.n144 GND.n143 76
R130 GND.n149 GND.n148 76
R131 GND.n152 GND.n151 76
R132 GND.n155 GND.n154 76
R133 GND.n162 GND.n161 76
R134 GND.n165 GND.n164 76
R135 GND.n168 GND.n167 76
R136 GND.n171 GND.n170 76
R137 GND.n174 GND.n173 76
R138 GND.n177 GND.n176 76
R139 GND.n180 GND.n179 76
R140 GND.n183 GND.n182 76
R141 GND.n186 GND.n185 76
R142 GND.n191 GND.n190 76
R143 GND.n194 GND.n193 76
R144 GND.n197 GND.n196 76
R145 GND.n204 GND.n203 76
R146 GND.n207 GND.n206 76
R147 GND.n210 GND.n209 76
R148 GND.n213 GND.n212 76
R149 GND.n216 GND.n215 76
R150 GND.n221 GND.n220 76
R151 GND.n224 GND.n223 76
R152 GND.n227 GND.n226 76
R153 GND.n234 GND.n233 76
R154 GND.n237 GND.n236 76
R155 GND.n240 GND.n239 76
R156 GND.n243 GND.n242 76
R157 GND.n246 GND.n245 76
R158 GND.n249 GND.n248 76
R159 GND.n252 GND.n251 76
R160 GND.n255 GND.n254 76
R161 GND.n258 GND.n257 76
R162 GND.n266 GND.n265 76
R163 GND.n269 GND.n268 76
R164 GND.n272 GND.n271 76
R165 GND.n279 GND.n278 76
R166 GND.n282 GND.n281 76
R167 GND.n285 GND.n284 76
R168 GND.n288 GND.n287 76
R169 GND.n291 GND.n290 76
R170 GND.n294 GND.n293 76
R171 GND.n297 GND.n296 76
R172 GND.n300 GND.n299 76
R173 GND.n303 GND.n302 76
R174 GND.n308 GND.n307 76
R175 GND.n311 GND.n310 76
R176 GND.n314 GND.n313 76
R177 GND.n321 GND.n320 76
R178 GND.n324 GND.n323 76
R179 GND.n327 GND.n326 76
R180 GND.n330 GND.n329 76
R181 GND.n333 GND.n332 76
R182 GND.n338 GND.n337 76
R183 GND.n341 GND.n340 76
R184 GND.n344 GND.n343 76
R185 GND.n351 GND.n350 76
R186 GND.n354 GND.n353 76
R187 GND.n357 GND.n356 76
R188 GND.n360 GND.n359 76
R189 GND.n363 GND.n362 76
R190 GND.n366 GND.n365 76
R191 GND.n369 GND.n368 76
R192 GND.n372 GND.n371 76
R193 GND.n375 GND.n374 76
R194 GND.n380 GND.n379 76
R195 GND.n383 GND.n382 76
R196 GND.n390 GND.n389 76
R197 GND.n773 GND.n772 76
R198 GND.n770 GND.n769 76
R199 GND.n767 GND.n766 76
R200 GND.n764 GND.n763 76
R201 GND.n761 GND.n760 76
R202 GND.n758 GND.n757 76
R203 GND.n755 GND.n754 76
R204 GND.n752 GND.n751 76
R205 GND.n749 GND.n748 76
R206 GND.n746 GND.n745 76
R207 GND.n741 GND.n740 76
R208 GND.n738 GND.n737 76
R209 GND.n731 GND.n730 76
R210 GND.n728 GND.n727 76
R211 GND.n725 GND.n724 76
R212 GND.n722 GND.n721 76
R213 GND.n719 GND.n718 76
R214 GND.n716 GND.n715 76
R215 GND.n711 GND.n710 76
R216 GND.n708 GND.n707 76
R217 GND.n701 GND.n700 76
R218 GND.n698 GND.n697 76
R219 GND.n695 GND.n694 76
R220 GND.n692 GND.n691 76
R221 GND.n689 GND.n688 76
R222 GND.n686 GND.n685 76
R223 GND.n683 GND.n682 76
R224 GND.n680 GND.n679 76
R225 GND.n677 GND.n676 76
R226 GND.n674 GND.n673 76
R227 GND.n669 GND.n668 76
R228 GND.n666 GND.n665 76
R229 GND.n659 GND.n658 76
R230 GND.n656 GND.n655 76
R231 GND.n653 GND.n652 76
R232 GND.n650 GND.n649 76
R233 GND.n647 GND.n646 76
R234 GND.n644 GND.n643 76
R235 GND.n641 GND.n640 76
R236 GND.n638 GND.n637 76
R237 GND.n635 GND.n634 76
R238 GND.n632 GND.n631 76
R239 GND.n627 GND.n626 76
R240 GND.n624 GND.n623 76
R241 GND.n617 GND.n616 76
R242 GND.n614 GND.n613 76
R243 GND.n611 GND.n610 76
R244 GND.n608 GND.n607 76
R245 GND.n605 GND.n604 76
R246 GND.n602 GND.n601 76
R247 GND.n597 GND.n596 76
R248 GND.n594 GND.n593 76
R249 GND.n587 GND.n586 76
R250 GND.n584 GND.n583 76
R251 GND.n581 GND.n580 76
R252 GND.n578 GND.n577 76
R253 GND.n575 GND.n574 76
R254 GND.n572 GND.n571 76
R255 GND.n569 GND.n568 76
R256 GND.n566 GND.n565 76
R257 GND.n563 GND.n562 76
R258 GND.n560 GND.n559 76
R259 GND.n555 GND.n554 76
R260 GND.n552 GND.n551 76
R261 GND.n545 GND.n544 76
R262 GND.n542 GND.n541 76
R263 GND.n539 GND.n538 76
R264 GND.n536 GND.n535 76
R265 GND.n533 GND.n532 76
R266 GND.n530 GND.n529 76
R267 GND.n527 GND.n526 76
R268 GND.n524 GND.n523 76
R269 GND.n521 GND.n520 76
R270 GND.n518 GND.n517 76
R271 GND.n513 GND.n512 76
R272 GND.n510 GND.n509 76
R273 GND.n503 GND.n502 76
R274 GND.n500 GND.n499 76
R275 GND.n497 GND.n496 76
R276 GND.n494 GND.n493 76
R277 GND.n491 GND.n490 76
R278 GND.n488 GND.n487 76
R279 GND.n480 GND.n479 76
R280 GND.n477 GND.n476 76
R281 GND.n470 GND.n469 76
R282 GND.n467 GND.n466 76
R283 GND.n464 GND.n463 76
R284 GND.n461 GND.n460 76
R285 GND.n458 GND.n457 76
R286 GND.n455 GND.n454 76
R287 GND.n452 GND.n451 76
R288 GND.n449 GND.n448 76
R289 GND.n446 GND.n445 76
R290 GND.n443 GND.n442 76
R291 GND.n438 GND.n437 76
R292 GND.n435 GND.n434 76
R293 GND.n428 GND.n427 76
R294 GND.n425 GND.n424 76
R295 GND.n422 GND.n421 76
R296 GND.n419 GND.n418 76
R297 GND.n416 GND.n415 76
R298 GND.n413 GND.n412 76
R299 GND.n410 GND.n409 76
R300 GND.n407 GND.n406 76
R301 GND.n404 GND.n403 76
R302 GND.n401 GND.n400 76
R303 GND.n396 GND.n395 76
R304 GND.n12 GND.n11 76
R305 GND.n17 GND.n16 76
R306 GND.n20 GND.n19 76
R307 GND.n23 GND.n22 76
R308 GND.n30 GND.n29 76
R309 GND.n33 GND.n32 76
R310 GND.n36 GND.n35 76
R311 GND.n264 GND.n263 64.552
R312 GND.n485 GND.n484 63.835
R313 GND.n8 GND.n7 34.942
R314 GND.n263 GND.n262 28.421
R315 GND.n484 GND.n483 28.421
R316 GND.n263 GND.n261 25.263
R317 GND.n484 GND.n482 25.263
R318 GND.n261 GND.n260 24.383
R319 GND.n482 GND.n481 24.383
R320 GND.n5 GND.n4 14.167
R321 GND.n4 GND.n2 14.167
R322 GND.n29 GND.n27 14.167
R323 GND.n59 GND.n57 14.167
R324 GND.n89 GND.n87 14.167
R325 GND.n119 GND.n117 14.167
R326 GND.n161 GND.n159 14.167
R327 GND.n203 GND.n201 14.167
R328 GND.n233 GND.n231 14.167
R329 GND.n278 GND.n276 14.167
R330 GND.n320 GND.n318 14.167
R331 GND.n350 GND.n348 14.167
R332 GND.n389 GND.n388 14.167
R333 GND.n737 GND.n736 14.167
R334 GND.n707 GND.n706 14.167
R335 GND.n665 GND.n664 14.167
R336 GND.n623 GND.n622 14.167
R337 GND.n593 GND.n592 14.167
R338 GND.n551 GND.n550 14.167
R339 GND.n509 GND.n508 14.167
R340 GND.n476 GND.n475 14.167
R341 GND.n434 GND.n433 14.167
R342 GND.n395 GND.n394 13.653
R343 GND.n400 GND.n397 13.653
R344 GND.n403 GND.n402 13.653
R345 GND.n406 GND.n405 13.653
R346 GND.n409 GND.n408 13.653
R347 GND.n412 GND.n411 13.653
R348 GND.n415 GND.n414 13.653
R349 GND.n418 GND.n417 13.653
R350 GND.n421 GND.n420 13.653
R351 GND.n424 GND.n423 13.653
R352 GND.n427 GND.n426 13.653
R353 GND.n434 GND.n429 13.653
R354 GND.n437 GND.n436 13.653
R355 GND.n442 GND.n439 13.653
R356 GND.n445 GND.n444 13.653
R357 GND.n448 GND.n447 13.653
R358 GND.n451 GND.n450 13.653
R359 GND.n454 GND.n453 13.653
R360 GND.n457 GND.n456 13.653
R361 GND.n460 GND.n459 13.653
R362 GND.n463 GND.n462 13.653
R363 GND.n466 GND.n465 13.653
R364 GND.n469 GND.n468 13.653
R365 GND.n476 GND.n471 13.653
R366 GND.n479 GND.n478 13.653
R367 GND.n487 GND.n486 13.653
R368 GND.n490 GND.n489 13.653
R369 GND.n493 GND.n492 13.653
R370 GND.n496 GND.n495 13.653
R371 GND.n499 GND.n498 13.653
R372 GND.n502 GND.n501 13.653
R373 GND.n509 GND.n504 13.653
R374 GND.n512 GND.n511 13.653
R375 GND.n517 GND.n514 13.653
R376 GND.n520 GND.n519 13.653
R377 GND.n523 GND.n522 13.653
R378 GND.n526 GND.n525 13.653
R379 GND.n529 GND.n528 13.653
R380 GND.n532 GND.n531 13.653
R381 GND.n535 GND.n534 13.653
R382 GND.n538 GND.n537 13.653
R383 GND.n541 GND.n540 13.653
R384 GND.n544 GND.n543 13.653
R385 GND.n551 GND.n546 13.653
R386 GND.n554 GND.n553 13.653
R387 GND.n559 GND.n556 13.653
R388 GND.n562 GND.n561 13.653
R389 GND.n565 GND.n564 13.653
R390 GND.n568 GND.n567 13.653
R391 GND.n571 GND.n570 13.653
R392 GND.n574 GND.n573 13.653
R393 GND.n577 GND.n576 13.653
R394 GND.n580 GND.n579 13.653
R395 GND.n583 GND.n582 13.653
R396 GND.n586 GND.n585 13.653
R397 GND.n593 GND.n588 13.653
R398 GND.n596 GND.n595 13.653
R399 GND.n601 GND.n600 13.653
R400 GND.n604 GND.n603 13.653
R401 GND.n607 GND.n606 13.653
R402 GND.n610 GND.n609 13.653
R403 GND.n613 GND.n612 13.653
R404 GND.n616 GND.n615 13.653
R405 GND.n623 GND.n618 13.653
R406 GND.n626 GND.n625 13.653
R407 GND.n631 GND.n628 13.653
R408 GND.n634 GND.n633 13.653
R409 GND.n637 GND.n636 13.653
R410 GND.n640 GND.n639 13.653
R411 GND.n643 GND.n642 13.653
R412 GND.n646 GND.n645 13.653
R413 GND.n649 GND.n648 13.653
R414 GND.n652 GND.n651 13.653
R415 GND.n655 GND.n654 13.653
R416 GND.n658 GND.n657 13.653
R417 GND.n665 GND.n660 13.653
R418 GND.n668 GND.n667 13.653
R419 GND.n673 GND.n670 13.653
R420 GND.n676 GND.n675 13.653
R421 GND.n679 GND.n678 13.653
R422 GND.n682 GND.n681 13.653
R423 GND.n685 GND.n684 13.653
R424 GND.n688 GND.n687 13.653
R425 GND.n691 GND.n690 13.653
R426 GND.n694 GND.n693 13.653
R427 GND.n697 GND.n696 13.653
R428 GND.n700 GND.n699 13.653
R429 GND.n707 GND.n702 13.653
R430 GND.n710 GND.n709 13.653
R431 GND.n715 GND.n714 13.653
R432 GND.n718 GND.n717 13.653
R433 GND.n721 GND.n720 13.653
R434 GND.n724 GND.n723 13.653
R435 GND.n727 GND.n726 13.653
R436 GND.n730 GND.n729 13.653
R437 GND.n737 GND.n732 13.653
R438 GND.n740 GND.n739 13.653
R439 GND.n745 GND.n742 13.653
R440 GND.n748 GND.n747 13.653
R441 GND.n751 GND.n750 13.653
R442 GND.n754 GND.n753 13.653
R443 GND.n757 GND.n756 13.653
R444 GND.n760 GND.n759 13.653
R445 GND.n763 GND.n762 13.653
R446 GND.n766 GND.n765 13.653
R447 GND.n769 GND.n768 13.653
R448 GND.n772 GND.n771 13.653
R449 GND.n389 GND.n384 13.653
R450 GND.n382 GND.n381 13.653
R451 GND.n379 GND.n376 13.653
R452 GND.n374 GND.n373 13.653
R453 GND.n371 GND.n370 13.653
R454 GND.n368 GND.n367 13.653
R455 GND.n365 GND.n364 13.653
R456 GND.n362 GND.n361 13.653
R457 GND.n359 GND.n358 13.653
R458 GND.n356 GND.n355 13.653
R459 GND.n353 GND.n352 13.653
R460 GND.n350 GND.n349 13.653
R461 GND.n343 GND.n342 13.653
R462 GND.n340 GND.n339 13.653
R463 GND.n337 GND.n336 13.653
R464 GND.n332 GND.n331 13.653
R465 GND.n329 GND.n328 13.653
R466 GND.n326 GND.n325 13.653
R467 GND.n323 GND.n322 13.653
R468 GND.n320 GND.n319 13.653
R469 GND.n313 GND.n312 13.653
R470 GND.n310 GND.n309 13.653
R471 GND.n307 GND.n304 13.653
R472 GND.n302 GND.n301 13.653
R473 GND.n299 GND.n298 13.653
R474 GND.n296 GND.n295 13.653
R475 GND.n293 GND.n292 13.653
R476 GND.n290 GND.n289 13.653
R477 GND.n287 GND.n286 13.653
R478 GND.n284 GND.n283 13.653
R479 GND.n281 GND.n280 13.653
R480 GND.n278 GND.n277 13.653
R481 GND.n271 GND.n270 13.653
R482 GND.n268 GND.n267 13.653
R483 GND.n265 GND.n259 13.653
R484 GND.n257 GND.n256 13.653
R485 GND.n254 GND.n253 13.653
R486 GND.n251 GND.n250 13.653
R487 GND.n248 GND.n247 13.653
R488 GND.n245 GND.n244 13.653
R489 GND.n242 GND.n241 13.653
R490 GND.n239 GND.n238 13.653
R491 GND.n236 GND.n235 13.653
R492 GND.n233 GND.n232 13.653
R493 GND.n226 GND.n225 13.653
R494 GND.n223 GND.n222 13.653
R495 GND.n220 GND.n219 13.653
R496 GND.n215 GND.n214 13.653
R497 GND.n212 GND.n211 13.653
R498 GND.n209 GND.n208 13.653
R499 GND.n206 GND.n205 13.653
R500 GND.n203 GND.n202 13.653
R501 GND.n196 GND.n195 13.653
R502 GND.n193 GND.n192 13.653
R503 GND.n190 GND.n187 13.653
R504 GND.n185 GND.n184 13.653
R505 GND.n182 GND.n181 13.653
R506 GND.n179 GND.n178 13.653
R507 GND.n176 GND.n175 13.653
R508 GND.n173 GND.n172 13.653
R509 GND.n170 GND.n169 13.653
R510 GND.n167 GND.n166 13.653
R511 GND.n164 GND.n163 13.653
R512 GND.n161 GND.n160 13.653
R513 GND.n154 GND.n153 13.653
R514 GND.n151 GND.n150 13.653
R515 GND.n148 GND.n145 13.653
R516 GND.n143 GND.n142 13.653
R517 GND.n140 GND.n139 13.653
R518 GND.n137 GND.n136 13.653
R519 GND.n134 GND.n133 13.653
R520 GND.n131 GND.n130 13.653
R521 GND.n128 GND.n127 13.653
R522 GND.n125 GND.n124 13.653
R523 GND.n122 GND.n121 13.653
R524 GND.n119 GND.n118 13.653
R525 GND.n112 GND.n111 13.653
R526 GND.n109 GND.n108 13.653
R527 GND.n106 GND.n105 13.653
R528 GND.n101 GND.n100 13.653
R529 GND.n98 GND.n97 13.653
R530 GND.n95 GND.n94 13.653
R531 GND.n92 GND.n91 13.653
R532 GND.n89 GND.n88 13.653
R533 GND.n82 GND.n81 13.653
R534 GND.n79 GND.n78 13.653
R535 GND.n76 GND.n75 13.653
R536 GND.n71 GND.n70 13.653
R537 GND.n68 GND.n67 13.653
R538 GND.n65 GND.n64 13.653
R539 GND.n62 GND.n61 13.653
R540 GND.n59 GND.n58 13.653
R541 GND.n52 GND.n51 13.653
R542 GND.n49 GND.n48 13.653
R543 GND.n46 GND.n45 13.653
R544 GND.n41 GND.n40 13.653
R545 GND.n38 GND.n37 13.653
R546 GND.n5 GND.n0 13.653
R547 GND.n4 GND.n3 13.653
R548 GND.n2 GND.n1 13.653
R549 GND.n11 GND.n10 13.653
R550 GND.n16 GND.n15 13.653
R551 GND.n19 GND.n18 13.653
R552 GND.n22 GND.n21 13.653
R553 GND.n29 GND.n28 13.653
R554 GND.n32 GND.n31 13.653
R555 GND.n35 GND.n34 13.653
R556 GND.n27 GND.n26 7.312
R557 GND.n57 GND.n56 7.312
R558 GND.n433 GND.n432 7.312
R559 GND.n475 GND.n474 7.312
R560 GND.n508 GND.n507 7.312
R561 GND.n550 GND.n549 7.312
R562 GND.n592 GND.n591 7.312
R563 GND.n622 GND.n621 7.312
R564 GND.n664 GND.n663 7.312
R565 GND.n706 GND.n705 7.312
R566 GND.n736 GND.n735 7.312
R567 GND.n388 GND.n387 7.312
R568 GND.n348 GND.n347 7.312
R569 GND.n318 GND.n317 7.312
R570 GND.n276 GND.n275 7.312
R571 GND.n231 GND.n230 7.312
R572 GND.n201 GND.n200 7.312
R573 GND.n159 GND.n158 7.312
R574 GND.n117 GND.n116 7.312
R575 GND.n87 GND.n86 7.312
R576 GND.n7 GND.n6 7.084
R577 GND.n7 GND.n5 6.475
R578 GND.n16 GND.n14 3.935
R579 GND.n46 GND.n44 3.935
R580 GND.n76 GND.n74 3.935
R581 GND.n106 GND.n104 3.935
R582 GND.n220 GND.n218 3.935
R583 GND.n337 GND.n335 3.935
R584 GND.n715 GND.n713 3.935
R585 GND.n601 GND.n599 3.935
R586 GND.n487 GND.n485 3.935
R587 GND.n392 GND.n391 0.596
R588 GND.n30 GND.n23 0.29
R589 GND.n60 GND.n53 0.29
R590 GND.n90 GND.n83 0.29
R591 GND.n120 GND.n113 0.29
R592 GND.n162 GND.n155 0.29
R593 GND.n204 GND.n197 0.29
R594 GND.n234 GND.n227 0.29
R595 GND.n279 GND.n272 0.29
R596 GND.n321 GND.n314 0.29
R597 GND.n351 GND.n344 0.29
R598 GND.n738 GND.n731 0.29
R599 GND.n708 GND.n701 0.29
R600 GND.n666 GND.n659 0.29
R601 GND.n624 GND.n617 0.29
R602 GND.n594 GND.n587 0.29
R603 GND.n552 GND.n545 0.29
R604 GND.n510 GND.n503 0.29
R605 GND.n477 GND.n470 0.29
R606 GND.n435 GND.n428 0.29
R607 GND GND.n773 0.219
R608 GND.n393 GND 0.207
R609 GND.n138 GND.n135 0.197
R610 GND.n180 GND.n177 0.197
R611 GND.n252 GND.n249 0.197
R612 GND.n297 GND.n294 0.197
R613 GND.n369 GND.n366 0.197
R614 GND.n758 GND.n755 0.197
R615 GND.n686 GND.n683 0.197
R616 GND.n644 GND.n641 0.197
R617 GND.n572 GND.n569 0.197
R618 GND.n530 GND.n527 0.197
R619 GND.n455 GND.n452 0.197
R620 GND.n413 GND.n410 0.197
R621 GND.n148 GND.n147 0.196
R622 GND.n190 GND.n189 0.196
R623 GND.n265 GND.n264 0.196
R624 GND.n307 GND.n306 0.196
R625 GND.n379 GND.n378 0.196
R626 GND.n745 GND.n744 0.196
R627 GND.n673 GND.n672 0.196
R628 GND.n631 GND.n630 0.196
R629 GND.n559 GND.n558 0.196
R630 GND.n517 GND.n516 0.196
R631 GND.n442 GND.n441 0.196
R632 GND.n400 GND.n399 0.196
R633 GND.n12 GND.n9 0.181
R634 GND.n42 GND.n39 0.181
R635 GND.n72 GND.n69 0.181
R636 GND.n102 GND.n99 0.181
R637 GND.n216 GND.n213 0.181
R638 GND.n333 GND.n330 0.181
R639 GND.n722 GND.n719 0.181
R640 GND.n608 GND.n605 0.181
R641 GND.n494 GND.n491 0.181
R642 GND.n9 GND.n8 0.145
R643 GND.n17 GND.n12 0.145
R644 GND.n20 GND.n17 0.145
R645 GND.n23 GND.n20 0.145
R646 GND.n33 GND.n30 0.145
R647 GND.n36 GND.n33 0.145
R648 GND.n39 GND.n36 0.145
R649 GND.n47 GND.n42 0.145
R650 GND.n50 GND.n47 0.145
R651 GND.n53 GND.n50 0.145
R652 GND.n63 GND.n60 0.145
R653 GND.n66 GND.n63 0.145
R654 GND.n69 GND.n66 0.145
R655 GND.n77 GND.n72 0.145
R656 GND.n80 GND.n77 0.145
R657 GND.n83 GND.n80 0.145
R658 GND.n93 GND.n90 0.145
R659 GND.n96 GND.n93 0.145
R660 GND.n99 GND.n96 0.145
R661 GND.n107 GND.n102 0.145
R662 GND.n110 GND.n107 0.145
R663 GND.n113 GND.n110 0.145
R664 GND.n123 GND.n120 0.145
R665 GND.n126 GND.n123 0.145
R666 GND.n129 GND.n126 0.145
R667 GND.n132 GND.n129 0.145
R668 GND.n135 GND.n132 0.145
R669 GND.n141 GND.n138 0.145
R670 GND.n144 GND.n141 0.145
R671 GND.n149 GND.n144 0.145
R672 GND.n152 GND.n149 0.145
R673 GND.n155 GND.n152 0.145
R674 GND.n165 GND.n162 0.145
R675 GND.n168 GND.n165 0.145
R676 GND.n171 GND.n168 0.145
R677 GND.n174 GND.n171 0.145
R678 GND.n177 GND.n174 0.145
R679 GND.n183 GND.n180 0.145
R680 GND.n186 GND.n183 0.145
R681 GND.n191 GND.n186 0.145
R682 GND.n194 GND.n191 0.145
R683 GND.n197 GND.n194 0.145
R684 GND.n207 GND.n204 0.145
R685 GND.n210 GND.n207 0.145
R686 GND.n213 GND.n210 0.145
R687 GND.n221 GND.n216 0.145
R688 GND.n224 GND.n221 0.145
R689 GND.n227 GND.n224 0.145
R690 GND.n237 GND.n234 0.145
R691 GND.n240 GND.n237 0.145
R692 GND.n243 GND.n240 0.145
R693 GND.n246 GND.n243 0.145
R694 GND.n249 GND.n246 0.145
R695 GND.n255 GND.n252 0.145
R696 GND.n258 GND.n255 0.145
R697 GND.n266 GND.n258 0.145
R698 GND.n269 GND.n266 0.145
R699 GND.n272 GND.n269 0.145
R700 GND.n282 GND.n279 0.145
R701 GND.n285 GND.n282 0.145
R702 GND.n288 GND.n285 0.145
R703 GND.n291 GND.n288 0.145
R704 GND.n294 GND.n291 0.145
R705 GND.n300 GND.n297 0.145
R706 GND.n303 GND.n300 0.145
R707 GND.n308 GND.n303 0.145
R708 GND.n311 GND.n308 0.145
R709 GND.n314 GND.n311 0.145
R710 GND.n324 GND.n321 0.145
R711 GND.n327 GND.n324 0.145
R712 GND.n330 GND.n327 0.145
R713 GND.n338 GND.n333 0.145
R714 GND.n341 GND.n338 0.145
R715 GND.n344 GND.n341 0.145
R716 GND.n354 GND.n351 0.145
R717 GND.n357 GND.n354 0.145
R718 GND.n360 GND.n357 0.145
R719 GND.n363 GND.n360 0.145
R720 GND.n366 GND.n363 0.145
R721 GND.n372 GND.n369 0.145
R722 GND.n375 GND.n372 0.145
R723 GND.n380 GND.n375 0.145
R724 GND.n383 GND.n380 0.145
R725 GND.n390 GND.n383 0.145
R726 GND.n773 GND.n770 0.145
R727 GND.n770 GND.n767 0.145
R728 GND.n767 GND.n764 0.145
R729 GND.n764 GND.n761 0.145
R730 GND.n761 GND.n758 0.145
R731 GND.n755 GND.n752 0.145
R732 GND.n752 GND.n749 0.145
R733 GND.n749 GND.n746 0.145
R734 GND.n746 GND.n741 0.145
R735 GND.n741 GND.n738 0.145
R736 GND.n731 GND.n728 0.145
R737 GND.n728 GND.n725 0.145
R738 GND.n725 GND.n722 0.145
R739 GND.n719 GND.n716 0.145
R740 GND.n716 GND.n711 0.145
R741 GND.n711 GND.n708 0.145
R742 GND.n701 GND.n698 0.145
R743 GND.n698 GND.n695 0.145
R744 GND.n695 GND.n692 0.145
R745 GND.n692 GND.n689 0.145
R746 GND.n689 GND.n686 0.145
R747 GND.n683 GND.n680 0.145
R748 GND.n680 GND.n677 0.145
R749 GND.n677 GND.n674 0.145
R750 GND.n674 GND.n669 0.145
R751 GND.n669 GND.n666 0.145
R752 GND.n659 GND.n656 0.145
R753 GND.n656 GND.n653 0.145
R754 GND.n653 GND.n650 0.145
R755 GND.n650 GND.n647 0.145
R756 GND.n647 GND.n644 0.145
R757 GND.n641 GND.n638 0.145
R758 GND.n638 GND.n635 0.145
R759 GND.n635 GND.n632 0.145
R760 GND.n632 GND.n627 0.145
R761 GND.n627 GND.n624 0.145
R762 GND.n617 GND.n614 0.145
R763 GND.n614 GND.n611 0.145
R764 GND.n611 GND.n608 0.145
R765 GND.n605 GND.n602 0.145
R766 GND.n602 GND.n597 0.145
R767 GND.n597 GND.n594 0.145
R768 GND.n587 GND.n584 0.145
R769 GND.n584 GND.n581 0.145
R770 GND.n581 GND.n578 0.145
R771 GND.n578 GND.n575 0.145
R772 GND.n575 GND.n572 0.145
R773 GND.n569 GND.n566 0.145
R774 GND.n566 GND.n563 0.145
R775 GND.n563 GND.n560 0.145
R776 GND.n560 GND.n555 0.145
R777 GND.n555 GND.n552 0.145
R778 GND.n545 GND.n542 0.145
R779 GND.n542 GND.n539 0.145
R780 GND.n539 GND.n536 0.145
R781 GND.n536 GND.n533 0.145
R782 GND.n533 GND.n530 0.145
R783 GND.n527 GND.n524 0.145
R784 GND.n524 GND.n521 0.145
R785 GND.n521 GND.n518 0.145
R786 GND.n518 GND.n513 0.145
R787 GND.n513 GND.n510 0.145
R788 GND.n503 GND.n500 0.145
R789 GND.n500 GND.n497 0.145
R790 GND.n497 GND.n494 0.145
R791 GND.n491 GND.n488 0.145
R792 GND.n488 GND.n480 0.145
R793 GND.n480 GND.n477 0.145
R794 GND.n470 GND.n467 0.145
R795 GND.n467 GND.n464 0.145
R796 GND.n464 GND.n461 0.145
R797 GND.n461 GND.n458 0.145
R798 GND.n458 GND.n455 0.145
R799 GND.n452 GND.n449 0.145
R800 GND.n449 GND.n446 0.145
R801 GND.n446 GND.n443 0.145
R802 GND.n443 GND.n438 0.145
R803 GND.n438 GND.n435 0.145
R804 GND.n428 GND.n425 0.145
R805 GND.n425 GND.n422 0.145
R806 GND.n422 GND.n419 0.145
R807 GND.n419 GND.n416 0.145
R808 GND.n416 GND.n413 0.145
R809 GND.n410 GND.n407 0.145
R810 GND.n407 GND.n404 0.145
R811 GND.n404 GND.n401 0.145
R812 GND.n401 GND.n396 0.145
R813 GND.n396 GND.n393 0.145
R814 GND GND.n390 0.07
R815 RN.n17 RN.t21 479.223
R816 RN.n8 RN.t12 479.223
R817 RN.n0 RN.t25 479.223
R818 RN.n23 RN.t10 454.685
R819 RN.n20 RN.t14 454.685
R820 RN.n14 RN.t0 454.685
R821 RN.n11 RN.t5 454.685
R822 RN.n5 RN.t13 454.685
R823 RN.n2 RN.t15 454.685
R824 RN.n23 RN.t17 428.979
R825 RN.n20 RN.t1 428.979
R826 RN.n14 RN.t8 428.979
R827 RN.n11 RN.t19 428.979
R828 RN.n5 RN.t3 428.979
R829 RN.n2 RN.t6 428.979
R830 RN.n17 RN.t23 375.52
R831 RN.n8 RN.t24 375.52
R832 RN.n0 RN.t9 375.52
R833 RN.n24 RN.n23 178.106
R834 RN.n21 RN.n20 178.106
R835 RN.n15 RN.n14 178.106
R836 RN.n12 RN.n11 178.106
R837 RN.n6 RN.n5 178.106
R838 RN.n3 RN.n2 178.106
R839 RN.n18 RN.n17 175.429
R840 RN.n9 RN.n8 175.429
R841 RN.n1 RN.n0 175.429
R842 RN.n18 RN.t18 162.048
R843 RN.n9 RN.t4 162.048
R844 RN.n1 RN.t22 162.048
R845 RN.n24 RN.t16 158.3
R846 RN.n21 RN.t7 158.3
R847 RN.n15 RN.t2 158.3
R848 RN.n12 RN.t26 158.3
R849 RN.n6 RN.t20 158.3
R850 RN.n3 RN.t11 158.3
R851 RN.n4 RN.n1 78.675
R852 RN.n4 RN.n3 76
R853 RN.n7 RN.n6 76
R854 RN.n10 RN.n9 76
R855 RN.n13 RN.n12 76
R856 RN.n16 RN.n15 76
R857 RN.n19 RN.n18 76
R858 RN.n22 RN.n21 76
R859 RN.n25 RN.n24 76
R860 RN.n10 RN.n7 10.293
R861 RN.n19 RN.n16 10.293
R862 RN.n7 RN.n4 5.94
R863 RN.n16 RN.n13 5.94
R864 RN.n25 RN.n22 5.94
R865 RN.n13 RN.n10 2.675
R866 RN.n22 RN.n19 2.675
R867 RN.n25 RN 0.046
R868 VDD.n880 VDD.n878 144.705
R869 VDD.n961 VDD.n959 144.705
R870 VDD.n1022 VDD.n1020 144.705
R871 VDD.n1103 VDD.n1101 144.705
R872 VDD.n1184 VDD.n1182 144.705
R873 VDD.n1245 VDD.n1243 144.705
R874 VDD.n1326 VDD.n1324 144.705
R875 VDD.n1407 VDD.n1405 144.705
R876 VDD.n1468 VDD.n1466 144.705
R877 VDD.n698 VDD.n696 144.705
R878 VDD.n775 VDD.n773 144.705
R879 VDD.n637 VDD.n635 144.705
R880 VDD.n556 VDD.n554 144.705
R881 VDD.n475 VDD.n473 144.705
R882 VDD.n414 VDD.n412 144.705
R883 VDD.n333 VDD.n331 144.705
R884 VDD.n252 VDD.n250 144.705
R885 VDD.n191 VDD.n189 144.705
R886 VDD.n130 VDD.n128 144.705
R887 VDD.n76 VDD.n74 144.705
R888 VDD.n39 VDD.n38 76
R889 VDD.n43 VDD.n42 76
R890 VDD.n47 VDD.n46 76
R891 VDD.n51 VDD.n50 76
R892 VDD.n78 VDD.n77 76
R893 VDD.n82 VDD.n81 76
R894 VDD.n86 VDD.n85 76
R895 VDD.n90 VDD.n89 76
R896 VDD.n94 VDD.n93 76
R897 VDD.n98 VDD.n97 76
R898 VDD.n102 VDD.n101 76
R899 VDD.n106 VDD.n105 76
R900 VDD.n132 VDD.n131 76
R901 VDD.n137 VDD.n136 76
R902 VDD.n142 VDD.n141 76
R903 VDD.n148 VDD.n147 76
R904 VDD.n153 VDD.n152 76
R905 VDD.n158 VDD.n157 76
R906 VDD.n163 VDD.n162 76
R907 VDD.n167 VDD.n166 76
R908 VDD.n193 VDD.n192 76
R909 VDD.n198 VDD.n197 76
R910 VDD.n203 VDD.n202 76
R911 VDD.n209 VDD.n208 76
R912 VDD.n214 VDD.n213 76
R913 VDD.n219 VDD.n218 76
R914 VDD.n224 VDD.n223 76
R915 VDD.n228 VDD.n227 76
R916 VDD.n254 VDD.n253 76
R917 VDD.n258 VDD.n257 76
R918 VDD.n262 VDD.n261 76
R919 VDD.n267 VDD.n266 76
R920 VDD.n274 VDD.n273 76
R921 VDD.n279 VDD.n278 76
R922 VDD.n284 VDD.n283 76
R923 VDD.n291 VDD.n290 76
R924 VDD.n296 VDD.n295 76
R925 VDD.n301 VDD.n300 76
R926 VDD.n305 VDD.n304 76
R927 VDD.n309 VDD.n308 76
R928 VDD.n335 VDD.n334 76
R929 VDD.n339 VDD.n338 76
R930 VDD.n343 VDD.n342 76
R931 VDD.n348 VDD.n347 76
R932 VDD.n355 VDD.n354 76
R933 VDD.n360 VDD.n359 76
R934 VDD.n365 VDD.n364 76
R935 VDD.n372 VDD.n371 76
R936 VDD.n377 VDD.n376 76
R937 VDD.n382 VDD.n381 76
R938 VDD.n386 VDD.n385 76
R939 VDD.n390 VDD.n389 76
R940 VDD.n416 VDD.n415 76
R941 VDD.n421 VDD.n420 76
R942 VDD.n426 VDD.n425 76
R943 VDD.n432 VDD.n431 76
R944 VDD.n437 VDD.n436 76
R945 VDD.n442 VDD.n441 76
R946 VDD.n447 VDD.n446 76
R947 VDD.n451 VDD.n450 76
R948 VDD.n477 VDD.n476 76
R949 VDD.n481 VDD.n480 76
R950 VDD.n485 VDD.n484 76
R951 VDD.n490 VDD.n489 76
R952 VDD.n497 VDD.n496 76
R953 VDD.n502 VDD.n501 76
R954 VDD.n507 VDD.n506 76
R955 VDD.n514 VDD.n513 76
R956 VDD.n519 VDD.n518 76
R957 VDD.n524 VDD.n523 76
R958 VDD.n528 VDD.n527 76
R959 VDD.n532 VDD.n531 76
R960 VDD.n558 VDD.n557 76
R961 VDD.n562 VDD.n561 76
R962 VDD.n566 VDD.n565 76
R963 VDD.n571 VDD.n570 76
R964 VDD.n578 VDD.n577 76
R965 VDD.n583 VDD.n582 76
R966 VDD.n588 VDD.n587 76
R967 VDD.n595 VDD.n594 76
R968 VDD.n600 VDD.n599 76
R969 VDD.n605 VDD.n604 76
R970 VDD.n609 VDD.n608 76
R971 VDD.n613 VDD.n612 76
R972 VDD.n639 VDD.n638 76
R973 VDD.n644 VDD.n643 76
R974 VDD.n649 VDD.n648 76
R975 VDD.n655 VDD.n654 76
R976 VDD.n660 VDD.n659 76
R977 VDD.n665 VDD.n664 76
R978 VDD.n670 VDD.n669 76
R979 VDD.n674 VDD.n673 76
R980 VDD.n700 VDD.n699 76
R981 VDD.n704 VDD.n703 76
R982 VDD.n708 VDD.n707 76
R983 VDD.n713 VDD.n712 76
R984 VDD.n720 VDD.n719 76
R985 VDD.n725 VDD.n724 76
R986 VDD.n730 VDD.n729 76
R987 VDD.n737 VDD.n736 76
R988 VDD.n742 VDD.n741 76
R989 VDD.n747 VDD.n746 76
R990 VDD.n751 VDD.n750 76
R991 VDD.n777 VDD.n776 76
R992 VDD.n1525 VDD.n1524 76
R993 VDD.n1521 VDD.n1520 76
R994 VDD.n1517 VDD.n1516 76
R995 VDD.n1513 VDD.n1512 76
R996 VDD.n1508 VDD.n1507 76
R997 VDD.n1501 VDD.n1500 76
R998 VDD.n1496 VDD.n1495 76
R999 VDD.n1491 VDD.n1490 76
R1000 VDD.n1484 VDD.n1483 76
R1001 VDD.n1479 VDD.n1478 76
R1002 VDD.n1474 VDD.n1473 76
R1003 VDD.n1470 VDD.n1469 76
R1004 VDD.n1444 VDD.n1443 76
R1005 VDD.n1440 VDD.n1439 76
R1006 VDD.n1435 VDD.n1434 76
R1007 VDD.n1430 VDD.n1429 76
R1008 VDD.n1424 VDD.n1423 76
R1009 VDD.n1419 VDD.n1418 76
R1010 VDD.n1414 VDD.n1413 76
R1011 VDD.n1409 VDD.n1408 76
R1012 VDD.n1383 VDD.n1382 76
R1013 VDD.n1379 VDD.n1378 76
R1014 VDD.n1375 VDD.n1374 76
R1015 VDD.n1371 VDD.n1370 76
R1016 VDD.n1366 VDD.n1365 76
R1017 VDD.n1359 VDD.n1358 76
R1018 VDD.n1354 VDD.n1353 76
R1019 VDD.n1349 VDD.n1348 76
R1020 VDD.n1342 VDD.n1341 76
R1021 VDD.n1337 VDD.n1336 76
R1022 VDD.n1332 VDD.n1331 76
R1023 VDD.n1328 VDD.n1327 76
R1024 VDD.n1302 VDD.n1301 76
R1025 VDD.n1298 VDD.n1297 76
R1026 VDD.n1294 VDD.n1293 76
R1027 VDD.n1290 VDD.n1289 76
R1028 VDD.n1285 VDD.n1284 76
R1029 VDD.n1278 VDD.n1277 76
R1030 VDD.n1273 VDD.n1272 76
R1031 VDD.n1268 VDD.n1267 76
R1032 VDD.n1261 VDD.n1260 76
R1033 VDD.n1256 VDD.n1255 76
R1034 VDD.n1251 VDD.n1250 76
R1035 VDD.n1247 VDD.n1246 76
R1036 VDD.n1221 VDD.n1220 76
R1037 VDD.n1217 VDD.n1216 76
R1038 VDD.n1212 VDD.n1211 76
R1039 VDD.n1207 VDD.n1206 76
R1040 VDD.n1201 VDD.n1200 76
R1041 VDD.n1196 VDD.n1195 76
R1042 VDD.n1191 VDD.n1190 76
R1043 VDD.n1186 VDD.n1185 76
R1044 VDD.n1160 VDD.n1159 76
R1045 VDD.n1156 VDD.n1155 76
R1046 VDD.n1152 VDD.n1151 76
R1047 VDD.n1148 VDD.n1147 76
R1048 VDD.n1143 VDD.n1142 76
R1049 VDD.n1136 VDD.n1135 76
R1050 VDD.n1131 VDD.n1130 76
R1051 VDD.n1126 VDD.n1125 76
R1052 VDD.n1119 VDD.n1118 76
R1053 VDD.n1114 VDD.n1113 76
R1054 VDD.n1109 VDD.n1108 76
R1055 VDD.n1105 VDD.n1104 76
R1056 VDD.n1079 VDD.n1078 76
R1057 VDD.n1075 VDD.n1074 76
R1058 VDD.n1071 VDD.n1070 76
R1059 VDD.n1067 VDD.n1066 76
R1060 VDD.n1062 VDD.n1061 76
R1061 VDD.n1055 VDD.n1054 76
R1062 VDD.n1050 VDD.n1049 76
R1063 VDD.n1045 VDD.n1044 76
R1064 VDD.n1038 VDD.n1037 76
R1065 VDD.n1033 VDD.n1032 76
R1066 VDD.n1028 VDD.n1027 76
R1067 VDD.n1024 VDD.n1023 76
R1068 VDD.n998 VDD.n997 76
R1069 VDD.n994 VDD.n993 76
R1070 VDD.n989 VDD.n988 76
R1071 VDD.n984 VDD.n983 76
R1072 VDD.n978 VDD.n977 76
R1073 VDD.n973 VDD.n972 76
R1074 VDD.n968 VDD.n967 76
R1075 VDD.n963 VDD.n962 76
R1076 VDD.n937 VDD.n936 76
R1077 VDD.n933 VDD.n932 76
R1078 VDD.n929 VDD.n928 76
R1079 VDD.n925 VDD.n924 76
R1080 VDD.n920 VDD.n919 76
R1081 VDD.n913 VDD.n912 76
R1082 VDD.n908 VDD.n907 76
R1083 VDD.n903 VDD.n902 76
R1084 VDD.n896 VDD.n895 76
R1085 VDD.n891 VDD.n890 76
R1086 VDD.n886 VDD.n885 76
R1087 VDD.n882 VDD.n881 76
R1088 VDD.n855 VDD.n854 76
R1089 VDD.n851 VDD.n850 76
R1090 VDD.n847 VDD.n846 76
R1091 VDD.n843 VDD.n842 76
R1092 VDD.n838 VDD.n837 76
R1093 VDD.n831 VDD.n830 76
R1094 VDD.n826 VDD.n825 76
R1095 VDD.n821 VDD.n820 76
R1096 VDD.n814 VDD.n813 76
R1097 VDD.n809 VDD.n808 76
R1098 VDD.n804 VDD.n803 76
R1099 VDD.n800 VDD.n799 76
R1100 VDD.n264 VDD.n263 64.064
R1101 VDD.n345 VDD.n344 64.064
R1102 VDD.n487 VDD.n486 64.064
R1103 VDD.n568 VDD.n567 64.064
R1104 VDD.n710 VDD.n709 64.064
R1105 VDD.n1510 VDD.n1509 64.064
R1106 VDD.n1368 VDD.n1367 64.064
R1107 VDD.n1287 VDD.n1286 64.064
R1108 VDD.n1145 VDD.n1144 64.064
R1109 VDD.n1064 VDD.n1063 64.064
R1110 VDD.n922 VDD.n921 64.064
R1111 VDD.n840 VDD.n839 64.064
R1112 VDD.n293 VDD.n292 59.488
R1113 VDD.n374 VDD.n373 59.488
R1114 VDD.n516 VDD.n515 59.488
R1115 VDD.n597 VDD.n596 59.488
R1116 VDD.n739 VDD.n738 59.488
R1117 VDD.n1481 VDD.n1480 59.488
R1118 VDD.n1339 VDD.n1338 59.488
R1119 VDD.n1258 VDD.n1257 59.488
R1120 VDD.n1116 VDD.n1115 59.488
R1121 VDD.n1035 VDD.n1034 59.488
R1122 VDD.n893 VDD.n892 59.488
R1123 VDD.n811 VDD.n810 59.488
R1124 VDD.n159 VDD.t72 55.465
R1125 VDD.n133 VDD.t0 55.465
R1126 VDD.n805 VDD.t46 55.106
R1127 VDD.n887 VDD.t34 55.106
R1128 VDD.n964 VDD.t62 55.106
R1129 VDD.n1029 VDD.t98 55.106
R1130 VDD.n1110 VDD.t92 55.106
R1131 VDD.n1187 VDD.t33 55.106
R1132 VDD.n1252 VDD.t50 55.106
R1133 VDD.n1333 VDD.t80 55.106
R1134 VDD.n1410 VDD.t69 55.106
R1135 VDD.n1475 VDD.t66 55.106
R1136 VDD.n743 VDD.t85 55.106
R1137 VDD.n666 VDD.t84 55.106
R1138 VDD.n601 VDD.t75 55.106
R1139 VDD.n520 VDD.t91 55.106
R1140 VDD.n443 VDD.t23 55.106
R1141 VDD.n378 VDD.t55 55.106
R1142 VDD.n297 VDD.t40 55.106
R1143 VDD.n220 VDD.t83 55.106
R1144 VDD.n846 VDD.t45 55.106
R1145 VDD.n928 VDD.t13 55.106
R1146 VDD.n1070 VDD.t5 55.106
R1147 VDD.n1151 VDD.t89 55.106
R1148 VDD.n1293 VDD.t43 55.106
R1149 VDD.n1374 VDD.t11 55.106
R1150 VDD.n1516 VDD.t14 55.106
R1151 VDD.n707 VDD.t38 55.106
R1152 VDD.n565 VDD.t24 55.106
R1153 VDD.n484 VDD.t8 55.106
R1154 VDD.n342 VDD.t17 55.106
R1155 VDD.n261 VDD.t97 55.106
R1156 VDD.n990 VDD.t52 55.106
R1157 VDD.n1213 VDD.t32 55.106
R1158 VDD.n1436 VDD.t28 55.106
R1159 VDD.n640 VDD.t67 55.106
R1160 VDD.n417 VDD.t59 55.106
R1161 VDD.n194 VDD.t79 55.106
R1162 VDD.n144 VDD.n143 41.183
R1163 VDD.n816 VDD.n815 40.824
R1164 VDD.n836 VDD.n835 40.824
R1165 VDD.n898 VDD.n897 40.824
R1166 VDD.n918 VDD.n917 40.824
R1167 VDD.n980 VDD.n979 40.824
R1168 VDD.n1040 VDD.n1039 40.824
R1169 VDD.n1060 VDD.n1059 40.824
R1170 VDD.n1121 VDD.n1120 40.824
R1171 VDD.n1141 VDD.n1140 40.824
R1172 VDD.n1203 VDD.n1202 40.824
R1173 VDD.n1263 VDD.n1262 40.824
R1174 VDD.n1283 VDD.n1282 40.824
R1175 VDD.n1344 VDD.n1343 40.824
R1176 VDD.n1364 VDD.n1363 40.824
R1177 VDD.n1426 VDD.n1425 40.824
R1178 VDD.n1486 VDD.n1485 40.824
R1179 VDD.n1506 VDD.n1505 40.824
R1180 VDD.n732 VDD.n731 40.824
R1181 VDD.n718 VDD.n717 40.824
R1182 VDD.n651 VDD.n650 40.824
R1183 VDD.n590 VDD.n589 40.824
R1184 VDD.n576 VDD.n575 40.824
R1185 VDD.n509 VDD.n508 40.824
R1186 VDD.n495 VDD.n494 40.824
R1187 VDD.n428 VDD.n427 40.824
R1188 VDD.n367 VDD.n366 40.824
R1189 VDD.n353 VDD.n352 40.824
R1190 VDD.n286 VDD.n285 40.824
R1191 VDD.n272 VDD.n271 40.824
R1192 VDD.n205 VDD.n204 40.824
R1193 VDD.n942 VDD.n941 36.774
R1194 VDD.n1003 VDD.n1002 36.774
R1195 VDD.n1084 VDD.n1083 36.774
R1196 VDD.n1165 VDD.n1164 36.774
R1197 VDD.n1226 VDD.n1225 36.774
R1198 VDD.n1307 VDD.n1306 36.774
R1199 VDD.n1388 VDD.n1387 36.774
R1200 VDD.n1449 VDD.n1448 36.774
R1201 VDD.n756 VDD.n755 36.774
R1202 VDD.n679 VDD.n678 36.774
R1203 VDD.n618 VDD.n617 36.774
R1204 VDD.n537 VDD.n536 36.774
R1205 VDD.n456 VDD.n455 36.774
R1206 VDD.n395 VDD.n394 36.774
R1207 VDD.n314 VDD.n313 36.774
R1208 VDD.n233 VDD.n232 36.774
R1209 VDD.n172 VDD.n171 36.774
R1210 VDD.n111 VDD.n110 36.774
R1211 VDD.n56 VDD.n55 36.774
R1212 VDD.n871 VDD.n870 36.774
R1213 VDD.n139 VDD.n138 36.608
R1214 VDD.n200 VDD.n199 36.608
R1215 VDD.n423 VDD.n422 36.608
R1216 VDD.n646 VDD.n645 36.608
R1217 VDD.n1432 VDD.n1431 36.608
R1218 VDD.n1209 VDD.n1208 36.608
R1219 VDD.n986 VDD.n985 36.608
R1220 VDD.n34 VDD.n33 34.942
R1221 VDD.n155 VDD.n154 32.032
R1222 VDD.n216 VDD.n215 32.032
R1223 VDD.n439 VDD.n438 32.032
R1224 VDD.n662 VDD.n661 32.032
R1225 VDD.n1416 VDD.n1415 32.032
R1226 VDD.n1193 VDD.n1192 32.032
R1227 VDD.n970 VDD.n969 32.032
R1228 VDD.n269 VDD.n268 27.456
R1229 VDD.n350 VDD.n349 27.456
R1230 VDD.n492 VDD.n491 27.456
R1231 VDD.n573 VDD.n572 27.456
R1232 VDD.n715 VDD.n714 27.456
R1233 VDD.n1503 VDD.n1502 27.456
R1234 VDD.n1361 VDD.n1360 27.456
R1235 VDD.n1280 VDD.n1279 27.456
R1236 VDD.n1138 VDD.n1137 27.456
R1237 VDD.n1057 VDD.n1056 27.456
R1238 VDD.n915 VDD.n914 27.456
R1239 VDD.n833 VDD.n832 27.456
R1240 VDD.n288 VDD.n287 22.88
R1241 VDD.n369 VDD.n368 22.88
R1242 VDD.n511 VDD.n510 22.88
R1243 VDD.n592 VDD.n591 22.88
R1244 VDD.n734 VDD.n733 22.88
R1245 VDD.n1488 VDD.n1487 22.88
R1246 VDD.n1346 VDD.n1345 22.88
R1247 VDD.n1265 VDD.n1264 22.88
R1248 VDD.n1123 VDD.n1122 22.88
R1249 VDD.n1042 VDD.n1041 22.88
R1250 VDD.n900 VDD.n899 22.88
R1251 VDD.n818 VDD.n817 22.88
R1252 VDD.n799 VDD.n796 21.841
R1253 VDD.n23 VDD.n20 21.841
R1254 VDD.n815 VDD.t26 14.282
R1255 VDD.n815 VDD.t64 14.282
R1256 VDD.n835 VDD.t73 14.282
R1257 VDD.n835 VDD.t78 14.282
R1258 VDD.n897 VDD.t49 14.282
R1259 VDD.n897 VDD.t71 14.282
R1260 VDD.n917 VDD.t10 14.282
R1261 VDD.n917 VDD.t48 14.282
R1262 VDD.n979 VDD.t47 14.282
R1263 VDD.n979 VDD.t74 14.282
R1264 VDD.n1039 VDD.t88 14.282
R1265 VDD.n1039 VDD.t70 14.282
R1266 VDD.n1059 VDD.t4 14.282
R1267 VDD.n1059 VDD.t57 14.282
R1268 VDD.n1120 VDD.t15 14.282
R1269 VDD.n1120 VDD.t35 14.282
R1270 VDD.n1140 VDD.t68 14.282
R1271 VDD.n1140 VDD.t21 14.282
R1272 VDD.n1202 VDD.t53 14.282
R1273 VDD.n1202 VDD.t1 14.282
R1274 VDD.n1262 VDD.t95 14.282
R1275 VDD.n1262 VDD.t90 14.282
R1276 VDD.n1282 VDD.t29 14.282
R1277 VDD.n1282 VDD.t87 14.282
R1278 VDD.n1343 VDD.t31 14.282
R1279 VDD.n1343 VDD.t94 14.282
R1280 VDD.n1363 VDD.t12 14.282
R1281 VDD.n1363 VDD.t30 14.282
R1282 VDD.n1425 VDD.t2 14.282
R1283 VDD.n1425 VDD.t44 14.282
R1284 VDD.n1485 VDD.t86 14.282
R1285 VDD.n1485 VDD.t51 14.282
R1286 VDD.n1505 VDD.t9 14.282
R1287 VDD.n1505 VDD.t99 14.282
R1288 VDD.n731 VDD.t16 14.282
R1289 VDD.n731 VDD.t93 14.282
R1290 VDD.n717 VDD.t39 14.282
R1291 VDD.n717 VDD.t20 14.282
R1292 VDD.n650 VDD.t54 14.282
R1293 VDD.n650 VDD.t41 14.282
R1294 VDD.n589 VDD.t76 14.282
R1295 VDD.n589 VDD.t96 14.282
R1296 VDD.n575 VDD.t22 14.282
R1297 VDD.n575 VDD.t65 14.282
R1298 VDD.n508 VDD.t77 14.282
R1299 VDD.n508 VDD.t61 14.282
R1300 VDD.n494 VDD.t7 14.282
R1301 VDD.n494 VDD.t37 14.282
R1302 VDD.n427 VDD.t60 14.282
R1303 VDD.n427 VDD.t25 14.282
R1304 VDD.n366 VDD.t81 14.282
R1305 VDD.n366 VDD.t3 14.282
R1306 VDD.n352 VDD.t6 14.282
R1307 VDD.n352 VDD.t36 14.282
R1308 VDD.n285 VDD.t18 14.282
R1309 VDD.n285 VDD.t63 14.282
R1310 VDD.n271 VDD.t27 14.282
R1311 VDD.n271 VDD.t19 14.282
R1312 VDD.n204 VDD.t56 14.282
R1313 VDD.n204 VDD.t82 14.282
R1314 VDD.n143 VDD.t58 14.282
R1315 VDD.n143 VDD.t42 14.282
R1316 VDD.n796 VDD.n779 14.167
R1317 VDD.n779 VDD.n778 14.167
R1318 VDD.n957 VDD.n939 14.167
R1319 VDD.n939 VDD.n938 14.167
R1320 VDD.n1018 VDD.n1000 14.167
R1321 VDD.n1000 VDD.n999 14.167
R1322 VDD.n1099 VDD.n1081 14.167
R1323 VDD.n1081 VDD.n1080 14.167
R1324 VDD.n1180 VDD.n1162 14.167
R1325 VDD.n1162 VDD.n1161 14.167
R1326 VDD.n1241 VDD.n1223 14.167
R1327 VDD.n1223 VDD.n1222 14.167
R1328 VDD.n1322 VDD.n1304 14.167
R1329 VDD.n1304 VDD.n1303 14.167
R1330 VDD.n1403 VDD.n1385 14.167
R1331 VDD.n1385 VDD.n1384 14.167
R1332 VDD.n1464 VDD.n1446 14.167
R1333 VDD.n1446 VDD.n1445 14.167
R1334 VDD.n771 VDD.n753 14.167
R1335 VDD.n753 VDD.n752 14.167
R1336 VDD.n694 VDD.n676 14.167
R1337 VDD.n676 VDD.n675 14.167
R1338 VDD.n633 VDD.n615 14.167
R1339 VDD.n615 VDD.n614 14.167
R1340 VDD.n552 VDD.n534 14.167
R1341 VDD.n534 VDD.n533 14.167
R1342 VDD.n471 VDD.n453 14.167
R1343 VDD.n453 VDD.n452 14.167
R1344 VDD.n410 VDD.n392 14.167
R1345 VDD.n392 VDD.n391 14.167
R1346 VDD.n329 VDD.n311 14.167
R1347 VDD.n311 VDD.n310 14.167
R1348 VDD.n248 VDD.n230 14.167
R1349 VDD.n230 VDD.n229 14.167
R1350 VDD.n187 VDD.n169 14.167
R1351 VDD.n169 VDD.n168 14.167
R1352 VDD.n126 VDD.n108 14.167
R1353 VDD.n108 VDD.n107 14.167
R1354 VDD.n72 VDD.n53 14.167
R1355 VDD.n53 VDD.n52 14.167
R1356 VDD.n876 VDD.n857 14.167
R1357 VDD.n857 VDD.n856 14.167
R1358 VDD.n20 VDD.n19 14.167
R1359 VDD.n19 VDD.n17 14.167
R1360 VDD.n32 VDD.n29 14.167
R1361 VDD.n29 VDD.n28 14.167
R1362 VDD.n77 VDD.n73 14.167
R1363 VDD.n131 VDD.n127 14.167
R1364 VDD.n192 VDD.n188 14.167
R1365 VDD.n253 VDD.n249 14.167
R1366 VDD.n334 VDD.n330 14.167
R1367 VDD.n415 VDD.n411 14.167
R1368 VDD.n476 VDD.n472 14.167
R1369 VDD.n557 VDD.n553 14.167
R1370 VDD.n638 VDD.n634 14.167
R1371 VDD.n699 VDD.n695 14.167
R1372 VDD.n776 VDD.n772 14.167
R1373 VDD.n1469 VDD.n1465 14.167
R1374 VDD.n1408 VDD.n1404 14.167
R1375 VDD.n1327 VDD.n1323 14.167
R1376 VDD.n1246 VDD.n1242 14.167
R1377 VDD.n1185 VDD.n1181 14.167
R1378 VDD.n1104 VDD.n1100 14.167
R1379 VDD.n1023 VDD.n1019 14.167
R1380 VDD.n962 VDD.n958 14.167
R1381 VDD.n881 VDD.n877 14.167
R1382 VDD.n281 VDD.n280 13.728
R1383 VDD.n362 VDD.n361 13.728
R1384 VDD.n504 VDD.n503 13.728
R1385 VDD.n585 VDD.n584 13.728
R1386 VDD.n727 VDD.n726 13.728
R1387 VDD.n1493 VDD.n1492 13.728
R1388 VDD.n1351 VDD.n1350 13.728
R1389 VDD.n1270 VDD.n1269 13.728
R1390 VDD.n1128 VDD.n1127 13.728
R1391 VDD.n1047 VDD.n1046 13.728
R1392 VDD.n905 VDD.n904 13.728
R1393 VDD.n823 VDD.n822 13.728
R1394 VDD.n23 VDD.n22 13.653
R1395 VDD.n22 VDD.n21 13.653
R1396 VDD.n32 VDD.n31 13.653
R1397 VDD.n31 VDD.n30 13.653
R1398 VDD.n29 VDD.n25 13.653
R1399 VDD.n25 VDD.n24 13.653
R1400 VDD.n28 VDD.n27 13.653
R1401 VDD.n27 VDD.n26 13.653
R1402 VDD.n38 VDD.n37 13.653
R1403 VDD.n37 VDD.n36 13.653
R1404 VDD.n42 VDD.n41 13.653
R1405 VDD.n41 VDD.n40 13.653
R1406 VDD.n46 VDD.n45 13.653
R1407 VDD.n45 VDD.n44 13.653
R1408 VDD.n50 VDD.n49 13.653
R1409 VDD.n49 VDD.n48 13.653
R1410 VDD.n77 VDD.n76 13.653
R1411 VDD.n76 VDD.n75 13.653
R1412 VDD.n81 VDD.n80 13.653
R1413 VDD.n80 VDD.n79 13.653
R1414 VDD.n85 VDD.n84 13.653
R1415 VDD.n84 VDD.n83 13.653
R1416 VDD.n89 VDD.n88 13.653
R1417 VDD.n88 VDD.n87 13.653
R1418 VDD.n93 VDD.n92 13.653
R1419 VDD.n92 VDD.n91 13.653
R1420 VDD.n97 VDD.n96 13.653
R1421 VDD.n96 VDD.n95 13.653
R1422 VDD.n101 VDD.n100 13.653
R1423 VDD.n100 VDD.n99 13.653
R1424 VDD.n105 VDD.n104 13.653
R1425 VDD.n104 VDD.n103 13.653
R1426 VDD.n131 VDD.n130 13.653
R1427 VDD.n130 VDD.n129 13.653
R1428 VDD.n136 VDD.n135 13.653
R1429 VDD.n135 VDD.n134 13.653
R1430 VDD.n141 VDD.n140 13.653
R1431 VDD.n140 VDD.n139 13.653
R1432 VDD.n147 VDD.n146 13.653
R1433 VDD.n146 VDD.n145 13.653
R1434 VDD.n152 VDD.n151 13.653
R1435 VDD.n151 VDD.n150 13.653
R1436 VDD.n157 VDD.n156 13.653
R1437 VDD.n156 VDD.n155 13.653
R1438 VDD.n162 VDD.n161 13.653
R1439 VDD.n161 VDD.n160 13.653
R1440 VDD.n166 VDD.n165 13.653
R1441 VDD.n165 VDD.n164 13.653
R1442 VDD.n192 VDD.n191 13.653
R1443 VDD.n191 VDD.n190 13.653
R1444 VDD.n197 VDD.n196 13.653
R1445 VDD.n196 VDD.n195 13.653
R1446 VDD.n202 VDD.n201 13.653
R1447 VDD.n201 VDD.n200 13.653
R1448 VDD.n208 VDD.n207 13.653
R1449 VDD.n207 VDD.n206 13.653
R1450 VDD.n213 VDD.n212 13.653
R1451 VDD.n212 VDD.n211 13.653
R1452 VDD.n218 VDD.n217 13.653
R1453 VDD.n217 VDD.n216 13.653
R1454 VDD.n223 VDD.n222 13.653
R1455 VDD.n222 VDD.n221 13.653
R1456 VDD.n227 VDD.n226 13.653
R1457 VDD.n226 VDD.n225 13.653
R1458 VDD.n253 VDD.n252 13.653
R1459 VDD.n252 VDD.n251 13.653
R1460 VDD.n257 VDD.n256 13.653
R1461 VDD.n256 VDD.n255 13.653
R1462 VDD.n261 VDD.n260 13.653
R1463 VDD.n260 VDD.n259 13.653
R1464 VDD.n266 VDD.n265 13.653
R1465 VDD.n265 VDD.n264 13.653
R1466 VDD.n273 VDD.n270 13.653
R1467 VDD.n270 VDD.n269 13.653
R1468 VDD.n278 VDD.n277 13.653
R1469 VDD.n277 VDD.n276 13.653
R1470 VDD.n283 VDD.n282 13.653
R1471 VDD.n282 VDD.n281 13.653
R1472 VDD.n290 VDD.n289 13.653
R1473 VDD.n289 VDD.n288 13.653
R1474 VDD.n295 VDD.n294 13.653
R1475 VDD.n294 VDD.n293 13.653
R1476 VDD.n300 VDD.n299 13.653
R1477 VDD.n299 VDD.n298 13.653
R1478 VDD.n304 VDD.n303 13.653
R1479 VDD.n303 VDD.n302 13.653
R1480 VDD.n308 VDD.n307 13.653
R1481 VDD.n307 VDD.n306 13.653
R1482 VDD.n334 VDD.n333 13.653
R1483 VDD.n333 VDD.n332 13.653
R1484 VDD.n338 VDD.n337 13.653
R1485 VDD.n337 VDD.n336 13.653
R1486 VDD.n342 VDD.n341 13.653
R1487 VDD.n341 VDD.n340 13.653
R1488 VDD.n347 VDD.n346 13.653
R1489 VDD.n346 VDD.n345 13.653
R1490 VDD.n354 VDD.n351 13.653
R1491 VDD.n351 VDD.n350 13.653
R1492 VDD.n359 VDD.n358 13.653
R1493 VDD.n358 VDD.n357 13.653
R1494 VDD.n364 VDD.n363 13.653
R1495 VDD.n363 VDD.n362 13.653
R1496 VDD.n371 VDD.n370 13.653
R1497 VDD.n370 VDD.n369 13.653
R1498 VDD.n376 VDD.n375 13.653
R1499 VDD.n375 VDD.n374 13.653
R1500 VDD.n381 VDD.n380 13.653
R1501 VDD.n380 VDD.n379 13.653
R1502 VDD.n385 VDD.n384 13.653
R1503 VDD.n384 VDD.n383 13.653
R1504 VDD.n389 VDD.n388 13.653
R1505 VDD.n388 VDD.n387 13.653
R1506 VDD.n415 VDD.n414 13.653
R1507 VDD.n414 VDD.n413 13.653
R1508 VDD.n420 VDD.n419 13.653
R1509 VDD.n419 VDD.n418 13.653
R1510 VDD.n425 VDD.n424 13.653
R1511 VDD.n424 VDD.n423 13.653
R1512 VDD.n431 VDD.n430 13.653
R1513 VDD.n430 VDD.n429 13.653
R1514 VDD.n436 VDD.n435 13.653
R1515 VDD.n435 VDD.n434 13.653
R1516 VDD.n441 VDD.n440 13.653
R1517 VDD.n440 VDD.n439 13.653
R1518 VDD.n446 VDD.n445 13.653
R1519 VDD.n445 VDD.n444 13.653
R1520 VDD.n450 VDD.n449 13.653
R1521 VDD.n449 VDD.n448 13.653
R1522 VDD.n476 VDD.n475 13.653
R1523 VDD.n475 VDD.n474 13.653
R1524 VDD.n480 VDD.n479 13.653
R1525 VDD.n479 VDD.n478 13.653
R1526 VDD.n484 VDD.n483 13.653
R1527 VDD.n483 VDD.n482 13.653
R1528 VDD.n489 VDD.n488 13.653
R1529 VDD.n488 VDD.n487 13.653
R1530 VDD.n496 VDD.n493 13.653
R1531 VDD.n493 VDD.n492 13.653
R1532 VDD.n501 VDD.n500 13.653
R1533 VDD.n500 VDD.n499 13.653
R1534 VDD.n506 VDD.n505 13.653
R1535 VDD.n505 VDD.n504 13.653
R1536 VDD.n513 VDD.n512 13.653
R1537 VDD.n512 VDD.n511 13.653
R1538 VDD.n518 VDD.n517 13.653
R1539 VDD.n517 VDD.n516 13.653
R1540 VDD.n523 VDD.n522 13.653
R1541 VDD.n522 VDD.n521 13.653
R1542 VDD.n527 VDD.n526 13.653
R1543 VDD.n526 VDD.n525 13.653
R1544 VDD.n531 VDD.n530 13.653
R1545 VDD.n530 VDD.n529 13.653
R1546 VDD.n557 VDD.n556 13.653
R1547 VDD.n556 VDD.n555 13.653
R1548 VDD.n561 VDD.n560 13.653
R1549 VDD.n560 VDD.n559 13.653
R1550 VDD.n565 VDD.n564 13.653
R1551 VDD.n564 VDD.n563 13.653
R1552 VDD.n570 VDD.n569 13.653
R1553 VDD.n569 VDD.n568 13.653
R1554 VDD.n577 VDD.n574 13.653
R1555 VDD.n574 VDD.n573 13.653
R1556 VDD.n582 VDD.n581 13.653
R1557 VDD.n581 VDD.n580 13.653
R1558 VDD.n587 VDD.n586 13.653
R1559 VDD.n586 VDD.n585 13.653
R1560 VDD.n594 VDD.n593 13.653
R1561 VDD.n593 VDD.n592 13.653
R1562 VDD.n599 VDD.n598 13.653
R1563 VDD.n598 VDD.n597 13.653
R1564 VDD.n604 VDD.n603 13.653
R1565 VDD.n603 VDD.n602 13.653
R1566 VDD.n608 VDD.n607 13.653
R1567 VDD.n607 VDD.n606 13.653
R1568 VDD.n612 VDD.n611 13.653
R1569 VDD.n611 VDD.n610 13.653
R1570 VDD.n638 VDD.n637 13.653
R1571 VDD.n637 VDD.n636 13.653
R1572 VDD.n643 VDD.n642 13.653
R1573 VDD.n642 VDD.n641 13.653
R1574 VDD.n648 VDD.n647 13.653
R1575 VDD.n647 VDD.n646 13.653
R1576 VDD.n654 VDD.n653 13.653
R1577 VDD.n653 VDD.n652 13.653
R1578 VDD.n659 VDD.n658 13.653
R1579 VDD.n658 VDD.n657 13.653
R1580 VDD.n664 VDD.n663 13.653
R1581 VDD.n663 VDD.n662 13.653
R1582 VDD.n669 VDD.n668 13.653
R1583 VDD.n668 VDD.n667 13.653
R1584 VDD.n673 VDD.n672 13.653
R1585 VDD.n672 VDD.n671 13.653
R1586 VDD.n699 VDD.n698 13.653
R1587 VDD.n698 VDD.n697 13.653
R1588 VDD.n703 VDD.n702 13.653
R1589 VDD.n702 VDD.n701 13.653
R1590 VDD.n707 VDD.n706 13.653
R1591 VDD.n706 VDD.n705 13.653
R1592 VDD.n712 VDD.n711 13.653
R1593 VDD.n711 VDD.n710 13.653
R1594 VDD.n719 VDD.n716 13.653
R1595 VDD.n716 VDD.n715 13.653
R1596 VDD.n724 VDD.n723 13.653
R1597 VDD.n723 VDD.n722 13.653
R1598 VDD.n729 VDD.n728 13.653
R1599 VDD.n728 VDD.n727 13.653
R1600 VDD.n736 VDD.n735 13.653
R1601 VDD.n735 VDD.n734 13.653
R1602 VDD.n741 VDD.n740 13.653
R1603 VDD.n740 VDD.n739 13.653
R1604 VDD.n746 VDD.n745 13.653
R1605 VDD.n745 VDD.n744 13.653
R1606 VDD.n750 VDD.n749 13.653
R1607 VDD.n749 VDD.n748 13.653
R1608 VDD.n776 VDD.n775 13.653
R1609 VDD.n775 VDD.n774 13.653
R1610 VDD.n1524 VDD.n1523 13.653
R1611 VDD.n1523 VDD.n1522 13.653
R1612 VDD.n1520 VDD.n1519 13.653
R1613 VDD.n1519 VDD.n1518 13.653
R1614 VDD.n1516 VDD.n1515 13.653
R1615 VDD.n1515 VDD.n1514 13.653
R1616 VDD.n1512 VDD.n1511 13.653
R1617 VDD.n1511 VDD.n1510 13.653
R1618 VDD.n1507 VDD.n1504 13.653
R1619 VDD.n1504 VDD.n1503 13.653
R1620 VDD.n1500 VDD.n1499 13.653
R1621 VDD.n1499 VDD.n1498 13.653
R1622 VDD.n1495 VDD.n1494 13.653
R1623 VDD.n1494 VDD.n1493 13.653
R1624 VDD.n1490 VDD.n1489 13.653
R1625 VDD.n1489 VDD.n1488 13.653
R1626 VDD.n1483 VDD.n1482 13.653
R1627 VDD.n1482 VDD.n1481 13.653
R1628 VDD.n1478 VDD.n1477 13.653
R1629 VDD.n1477 VDD.n1476 13.653
R1630 VDD.n1473 VDD.n1472 13.653
R1631 VDD.n1472 VDD.n1471 13.653
R1632 VDD.n1469 VDD.n1468 13.653
R1633 VDD.n1468 VDD.n1467 13.653
R1634 VDD.n1443 VDD.n1442 13.653
R1635 VDD.n1442 VDD.n1441 13.653
R1636 VDD.n1439 VDD.n1438 13.653
R1637 VDD.n1438 VDD.n1437 13.653
R1638 VDD.n1434 VDD.n1433 13.653
R1639 VDD.n1433 VDD.n1432 13.653
R1640 VDD.n1429 VDD.n1428 13.653
R1641 VDD.n1428 VDD.n1427 13.653
R1642 VDD.n1423 VDD.n1422 13.653
R1643 VDD.n1422 VDD.n1421 13.653
R1644 VDD.n1418 VDD.n1417 13.653
R1645 VDD.n1417 VDD.n1416 13.653
R1646 VDD.n1413 VDD.n1412 13.653
R1647 VDD.n1412 VDD.n1411 13.653
R1648 VDD.n1408 VDD.n1407 13.653
R1649 VDD.n1407 VDD.n1406 13.653
R1650 VDD.n1382 VDD.n1381 13.653
R1651 VDD.n1381 VDD.n1380 13.653
R1652 VDD.n1378 VDD.n1377 13.653
R1653 VDD.n1377 VDD.n1376 13.653
R1654 VDD.n1374 VDD.n1373 13.653
R1655 VDD.n1373 VDD.n1372 13.653
R1656 VDD.n1370 VDD.n1369 13.653
R1657 VDD.n1369 VDD.n1368 13.653
R1658 VDD.n1365 VDD.n1362 13.653
R1659 VDD.n1362 VDD.n1361 13.653
R1660 VDD.n1358 VDD.n1357 13.653
R1661 VDD.n1357 VDD.n1356 13.653
R1662 VDD.n1353 VDD.n1352 13.653
R1663 VDD.n1352 VDD.n1351 13.653
R1664 VDD.n1348 VDD.n1347 13.653
R1665 VDD.n1347 VDD.n1346 13.653
R1666 VDD.n1341 VDD.n1340 13.653
R1667 VDD.n1340 VDD.n1339 13.653
R1668 VDD.n1336 VDD.n1335 13.653
R1669 VDD.n1335 VDD.n1334 13.653
R1670 VDD.n1331 VDD.n1330 13.653
R1671 VDD.n1330 VDD.n1329 13.653
R1672 VDD.n1327 VDD.n1326 13.653
R1673 VDD.n1326 VDD.n1325 13.653
R1674 VDD.n1301 VDD.n1300 13.653
R1675 VDD.n1300 VDD.n1299 13.653
R1676 VDD.n1297 VDD.n1296 13.653
R1677 VDD.n1296 VDD.n1295 13.653
R1678 VDD.n1293 VDD.n1292 13.653
R1679 VDD.n1292 VDD.n1291 13.653
R1680 VDD.n1289 VDD.n1288 13.653
R1681 VDD.n1288 VDD.n1287 13.653
R1682 VDD.n1284 VDD.n1281 13.653
R1683 VDD.n1281 VDD.n1280 13.653
R1684 VDD.n1277 VDD.n1276 13.653
R1685 VDD.n1276 VDD.n1275 13.653
R1686 VDD.n1272 VDD.n1271 13.653
R1687 VDD.n1271 VDD.n1270 13.653
R1688 VDD.n1267 VDD.n1266 13.653
R1689 VDD.n1266 VDD.n1265 13.653
R1690 VDD.n1260 VDD.n1259 13.653
R1691 VDD.n1259 VDD.n1258 13.653
R1692 VDD.n1255 VDD.n1254 13.653
R1693 VDD.n1254 VDD.n1253 13.653
R1694 VDD.n1250 VDD.n1249 13.653
R1695 VDD.n1249 VDD.n1248 13.653
R1696 VDD.n1246 VDD.n1245 13.653
R1697 VDD.n1245 VDD.n1244 13.653
R1698 VDD.n1220 VDD.n1219 13.653
R1699 VDD.n1219 VDD.n1218 13.653
R1700 VDD.n1216 VDD.n1215 13.653
R1701 VDD.n1215 VDD.n1214 13.653
R1702 VDD.n1211 VDD.n1210 13.653
R1703 VDD.n1210 VDD.n1209 13.653
R1704 VDD.n1206 VDD.n1205 13.653
R1705 VDD.n1205 VDD.n1204 13.653
R1706 VDD.n1200 VDD.n1199 13.653
R1707 VDD.n1199 VDD.n1198 13.653
R1708 VDD.n1195 VDD.n1194 13.653
R1709 VDD.n1194 VDD.n1193 13.653
R1710 VDD.n1190 VDD.n1189 13.653
R1711 VDD.n1189 VDD.n1188 13.653
R1712 VDD.n1185 VDD.n1184 13.653
R1713 VDD.n1184 VDD.n1183 13.653
R1714 VDD.n1159 VDD.n1158 13.653
R1715 VDD.n1158 VDD.n1157 13.653
R1716 VDD.n1155 VDD.n1154 13.653
R1717 VDD.n1154 VDD.n1153 13.653
R1718 VDD.n1151 VDD.n1150 13.653
R1719 VDD.n1150 VDD.n1149 13.653
R1720 VDD.n1147 VDD.n1146 13.653
R1721 VDD.n1146 VDD.n1145 13.653
R1722 VDD.n1142 VDD.n1139 13.653
R1723 VDD.n1139 VDD.n1138 13.653
R1724 VDD.n1135 VDD.n1134 13.653
R1725 VDD.n1134 VDD.n1133 13.653
R1726 VDD.n1130 VDD.n1129 13.653
R1727 VDD.n1129 VDD.n1128 13.653
R1728 VDD.n1125 VDD.n1124 13.653
R1729 VDD.n1124 VDD.n1123 13.653
R1730 VDD.n1118 VDD.n1117 13.653
R1731 VDD.n1117 VDD.n1116 13.653
R1732 VDD.n1113 VDD.n1112 13.653
R1733 VDD.n1112 VDD.n1111 13.653
R1734 VDD.n1108 VDD.n1107 13.653
R1735 VDD.n1107 VDD.n1106 13.653
R1736 VDD.n1104 VDD.n1103 13.653
R1737 VDD.n1103 VDD.n1102 13.653
R1738 VDD.n1078 VDD.n1077 13.653
R1739 VDD.n1077 VDD.n1076 13.653
R1740 VDD.n1074 VDD.n1073 13.653
R1741 VDD.n1073 VDD.n1072 13.653
R1742 VDD.n1070 VDD.n1069 13.653
R1743 VDD.n1069 VDD.n1068 13.653
R1744 VDD.n1066 VDD.n1065 13.653
R1745 VDD.n1065 VDD.n1064 13.653
R1746 VDD.n1061 VDD.n1058 13.653
R1747 VDD.n1058 VDD.n1057 13.653
R1748 VDD.n1054 VDD.n1053 13.653
R1749 VDD.n1053 VDD.n1052 13.653
R1750 VDD.n1049 VDD.n1048 13.653
R1751 VDD.n1048 VDD.n1047 13.653
R1752 VDD.n1044 VDD.n1043 13.653
R1753 VDD.n1043 VDD.n1042 13.653
R1754 VDD.n1037 VDD.n1036 13.653
R1755 VDD.n1036 VDD.n1035 13.653
R1756 VDD.n1032 VDD.n1031 13.653
R1757 VDD.n1031 VDD.n1030 13.653
R1758 VDD.n1027 VDD.n1026 13.653
R1759 VDD.n1026 VDD.n1025 13.653
R1760 VDD.n1023 VDD.n1022 13.653
R1761 VDD.n1022 VDD.n1021 13.653
R1762 VDD.n997 VDD.n996 13.653
R1763 VDD.n996 VDD.n995 13.653
R1764 VDD.n993 VDD.n992 13.653
R1765 VDD.n992 VDD.n991 13.653
R1766 VDD.n988 VDD.n987 13.653
R1767 VDD.n987 VDD.n986 13.653
R1768 VDD.n983 VDD.n982 13.653
R1769 VDD.n982 VDD.n981 13.653
R1770 VDD.n977 VDD.n976 13.653
R1771 VDD.n976 VDD.n975 13.653
R1772 VDD.n972 VDD.n971 13.653
R1773 VDD.n971 VDD.n970 13.653
R1774 VDD.n967 VDD.n966 13.653
R1775 VDD.n966 VDD.n965 13.653
R1776 VDD.n962 VDD.n961 13.653
R1777 VDD.n961 VDD.n960 13.653
R1778 VDD.n936 VDD.n935 13.653
R1779 VDD.n935 VDD.n934 13.653
R1780 VDD.n932 VDD.n931 13.653
R1781 VDD.n931 VDD.n930 13.653
R1782 VDD.n928 VDD.n927 13.653
R1783 VDD.n927 VDD.n926 13.653
R1784 VDD.n924 VDD.n923 13.653
R1785 VDD.n923 VDD.n922 13.653
R1786 VDD.n919 VDD.n916 13.653
R1787 VDD.n916 VDD.n915 13.653
R1788 VDD.n912 VDD.n911 13.653
R1789 VDD.n911 VDD.n910 13.653
R1790 VDD.n907 VDD.n906 13.653
R1791 VDD.n906 VDD.n905 13.653
R1792 VDD.n902 VDD.n901 13.653
R1793 VDD.n901 VDD.n900 13.653
R1794 VDD.n895 VDD.n894 13.653
R1795 VDD.n894 VDD.n893 13.653
R1796 VDD.n890 VDD.n889 13.653
R1797 VDD.n889 VDD.n888 13.653
R1798 VDD.n885 VDD.n884 13.653
R1799 VDD.n884 VDD.n883 13.653
R1800 VDD.n881 VDD.n880 13.653
R1801 VDD.n880 VDD.n879 13.653
R1802 VDD.n854 VDD.n853 13.653
R1803 VDD.n853 VDD.n852 13.653
R1804 VDD.n850 VDD.n849 13.653
R1805 VDD.n849 VDD.n848 13.653
R1806 VDD.n846 VDD.n845 13.653
R1807 VDD.n845 VDD.n844 13.653
R1808 VDD.n842 VDD.n841 13.653
R1809 VDD.n841 VDD.n840 13.653
R1810 VDD.n837 VDD.n834 13.653
R1811 VDD.n834 VDD.n833 13.653
R1812 VDD.n830 VDD.n829 13.653
R1813 VDD.n829 VDD.n828 13.653
R1814 VDD.n825 VDD.n824 13.653
R1815 VDD.n824 VDD.n823 13.653
R1816 VDD.n820 VDD.n819 13.653
R1817 VDD.n819 VDD.n818 13.653
R1818 VDD.n813 VDD.n812 13.653
R1819 VDD.n812 VDD.n811 13.653
R1820 VDD.n808 VDD.n807 13.653
R1821 VDD.n807 VDD.n806 13.653
R1822 VDD.n803 VDD.n802 13.653
R1823 VDD.n802 VDD.n801 13.653
R1824 VDD.n799 VDD.n798 13.653
R1825 VDD.n798 VDD.n797 13.653
R1826 VDD.n4 VDD.n2 12.915
R1827 VDD.n4 VDD.n3 12.66
R1828 VDD.n12 VDD.n11 12.343
R1829 VDD.n10 VDD.n9 12.343
R1830 VDD.n7 VDD.n6 12.343
R1831 VDD.n276 VDD.n275 9.152
R1832 VDD.n357 VDD.n356 9.152
R1833 VDD.n499 VDD.n498 9.152
R1834 VDD.n580 VDD.n579 9.152
R1835 VDD.n722 VDD.n721 9.152
R1836 VDD.n1498 VDD.n1497 9.152
R1837 VDD.n1356 VDD.n1355 9.152
R1838 VDD.n1275 VDD.n1274 9.152
R1839 VDD.n1133 VDD.n1132 9.152
R1840 VDD.n1052 VDD.n1051 9.152
R1841 VDD.n910 VDD.n909 9.152
R1842 VDD.n828 VDD.n827 9.152
R1843 VDD.n147 VDD.n144 8.658
R1844 VDD.n208 VDD.n205 8.658
R1845 VDD.n431 VDD.n428 8.658
R1846 VDD.n654 VDD.n651 8.658
R1847 VDD.n1429 VDD.n1426 8.658
R1848 VDD.n1206 VDD.n1203 8.658
R1849 VDD.n983 VDD.n980 8.658
R1850 VDD.n958 VDD.n957 7.674
R1851 VDD.n1019 VDD.n1018 7.674
R1852 VDD.n1100 VDD.n1099 7.674
R1853 VDD.n1181 VDD.n1180 7.674
R1854 VDD.n1242 VDD.n1241 7.674
R1855 VDD.n1323 VDD.n1322 7.674
R1856 VDD.n1404 VDD.n1403 7.674
R1857 VDD.n1465 VDD.n1464 7.674
R1858 VDD.n772 VDD.n771 7.674
R1859 VDD.n695 VDD.n694 7.674
R1860 VDD.n634 VDD.n633 7.674
R1861 VDD.n553 VDD.n552 7.674
R1862 VDD.n472 VDD.n471 7.674
R1863 VDD.n411 VDD.n410 7.674
R1864 VDD.n330 VDD.n329 7.674
R1865 VDD.n249 VDD.n248 7.674
R1866 VDD.n188 VDD.n187 7.674
R1867 VDD.n127 VDD.n126 7.674
R1868 VDD.n73 VDD.n72 7.674
R1869 VDD.n877 VDD.n876 7.674
R1870 VDD.n67 VDD.n66 7.5
R1871 VDD.n61 VDD.n60 7.5
R1872 VDD.n63 VDD.n62 7.5
R1873 VDD.n58 VDD.n57 7.5
R1874 VDD.n72 VDD.n71 7.5
R1875 VDD.n121 VDD.n120 7.5
R1876 VDD.n115 VDD.n114 7.5
R1877 VDD.n117 VDD.n116 7.5
R1878 VDD.n123 VDD.n113 7.5
R1879 VDD.n123 VDD.n111 7.5
R1880 VDD.n126 VDD.n125 7.5
R1881 VDD.n182 VDD.n181 7.5
R1882 VDD.n176 VDD.n175 7.5
R1883 VDD.n178 VDD.n177 7.5
R1884 VDD.n184 VDD.n174 7.5
R1885 VDD.n184 VDD.n172 7.5
R1886 VDD.n187 VDD.n186 7.5
R1887 VDD.n243 VDD.n242 7.5
R1888 VDD.n237 VDD.n236 7.5
R1889 VDD.n239 VDD.n238 7.5
R1890 VDD.n245 VDD.n235 7.5
R1891 VDD.n245 VDD.n233 7.5
R1892 VDD.n248 VDD.n247 7.5
R1893 VDD.n324 VDD.n323 7.5
R1894 VDD.n318 VDD.n317 7.5
R1895 VDD.n320 VDD.n319 7.5
R1896 VDD.n326 VDD.n316 7.5
R1897 VDD.n326 VDD.n314 7.5
R1898 VDD.n329 VDD.n328 7.5
R1899 VDD.n405 VDD.n404 7.5
R1900 VDD.n399 VDD.n398 7.5
R1901 VDD.n401 VDD.n400 7.5
R1902 VDD.n407 VDD.n397 7.5
R1903 VDD.n407 VDD.n395 7.5
R1904 VDD.n410 VDD.n409 7.5
R1905 VDD.n466 VDD.n465 7.5
R1906 VDD.n460 VDD.n459 7.5
R1907 VDD.n462 VDD.n461 7.5
R1908 VDD.n468 VDD.n458 7.5
R1909 VDD.n468 VDD.n456 7.5
R1910 VDD.n471 VDD.n470 7.5
R1911 VDD.n547 VDD.n546 7.5
R1912 VDD.n541 VDD.n540 7.5
R1913 VDD.n543 VDD.n542 7.5
R1914 VDD.n549 VDD.n539 7.5
R1915 VDD.n549 VDD.n537 7.5
R1916 VDD.n552 VDD.n551 7.5
R1917 VDD.n628 VDD.n627 7.5
R1918 VDD.n622 VDD.n621 7.5
R1919 VDD.n624 VDD.n623 7.5
R1920 VDD.n630 VDD.n620 7.5
R1921 VDD.n630 VDD.n618 7.5
R1922 VDD.n633 VDD.n632 7.5
R1923 VDD.n689 VDD.n688 7.5
R1924 VDD.n683 VDD.n682 7.5
R1925 VDD.n685 VDD.n684 7.5
R1926 VDD.n691 VDD.n681 7.5
R1927 VDD.n691 VDD.n679 7.5
R1928 VDD.n694 VDD.n693 7.5
R1929 VDD.n766 VDD.n765 7.5
R1930 VDD.n760 VDD.n759 7.5
R1931 VDD.n762 VDD.n761 7.5
R1932 VDD.n768 VDD.n758 7.5
R1933 VDD.n768 VDD.n756 7.5
R1934 VDD.n771 VDD.n770 7.5
R1935 VDD.n1459 VDD.n1458 7.5
R1936 VDD.n1453 VDD.n1452 7.5
R1937 VDD.n1455 VDD.n1454 7.5
R1938 VDD.n1461 VDD.n1451 7.5
R1939 VDD.n1461 VDD.n1449 7.5
R1940 VDD.n1464 VDD.n1463 7.5
R1941 VDD.n1398 VDD.n1397 7.5
R1942 VDD.n1392 VDD.n1391 7.5
R1943 VDD.n1394 VDD.n1393 7.5
R1944 VDD.n1400 VDD.n1390 7.5
R1945 VDD.n1400 VDD.n1388 7.5
R1946 VDD.n1403 VDD.n1402 7.5
R1947 VDD.n1317 VDD.n1316 7.5
R1948 VDD.n1311 VDD.n1310 7.5
R1949 VDD.n1313 VDD.n1312 7.5
R1950 VDD.n1319 VDD.n1309 7.5
R1951 VDD.n1319 VDD.n1307 7.5
R1952 VDD.n1322 VDD.n1321 7.5
R1953 VDD.n1236 VDD.n1235 7.5
R1954 VDD.n1230 VDD.n1229 7.5
R1955 VDD.n1232 VDD.n1231 7.5
R1956 VDD.n1238 VDD.n1228 7.5
R1957 VDD.n1238 VDD.n1226 7.5
R1958 VDD.n1241 VDD.n1240 7.5
R1959 VDD.n1175 VDD.n1174 7.5
R1960 VDD.n1169 VDD.n1168 7.5
R1961 VDD.n1171 VDD.n1170 7.5
R1962 VDD.n1177 VDD.n1167 7.5
R1963 VDD.n1177 VDD.n1165 7.5
R1964 VDD.n1180 VDD.n1179 7.5
R1965 VDD.n1094 VDD.n1093 7.5
R1966 VDD.n1088 VDD.n1087 7.5
R1967 VDD.n1090 VDD.n1089 7.5
R1968 VDD.n1096 VDD.n1086 7.5
R1969 VDD.n1096 VDD.n1084 7.5
R1970 VDD.n1099 VDD.n1098 7.5
R1971 VDD.n1013 VDD.n1012 7.5
R1972 VDD.n1007 VDD.n1006 7.5
R1973 VDD.n1009 VDD.n1008 7.5
R1974 VDD.n1015 VDD.n1005 7.5
R1975 VDD.n1015 VDD.n1003 7.5
R1976 VDD.n1018 VDD.n1017 7.5
R1977 VDD.n952 VDD.n951 7.5
R1978 VDD.n946 VDD.n945 7.5
R1979 VDD.n948 VDD.n947 7.5
R1980 VDD.n954 VDD.n944 7.5
R1981 VDD.n954 VDD.n942 7.5
R1982 VDD.n957 VDD.n956 7.5
R1983 VDD.n861 VDD.n860 7.5
R1984 VDD.n864 VDD.n863 7.5
R1985 VDD.n866 VDD.n865 7.5
R1986 VDD.n869 VDD.n868 7.5
R1987 VDD.n876 VDD.n875 7.5
R1988 VDD.n791 VDD.n790 7.5
R1989 VDD.n785 VDD.n784 7.5
R1990 VDD.n787 VDD.n786 7.5
R1991 VDD.n793 VDD.n783 7.5
R1992 VDD.n793 VDD.n781 7.5
R1993 VDD.n796 VDD.n795 7.5
R1994 VDD.n20 VDD.n16 7.5
R1995 VDD.n2 VDD.n1 7.5
R1996 VDD.n6 VDD.n5 7.5
R1997 VDD.n9 VDD.n8 7.5
R1998 VDD.n19 VDD.n18 7.5
R1999 VDD.n14 VDD.n0 7.5
R2000 VDD.n59 VDD.n56 6.772
R2001 VDD.n70 VDD.n54 6.772
R2002 VDD.n68 VDD.n65 6.772
R2003 VDD.n64 VDD.n61 6.772
R2004 VDD.n124 VDD.n109 6.772
R2005 VDD.n122 VDD.n119 6.772
R2006 VDD.n118 VDD.n115 6.772
R2007 VDD.n185 VDD.n170 6.772
R2008 VDD.n183 VDD.n180 6.772
R2009 VDD.n179 VDD.n176 6.772
R2010 VDD.n246 VDD.n231 6.772
R2011 VDD.n244 VDD.n241 6.772
R2012 VDD.n240 VDD.n237 6.772
R2013 VDD.n327 VDD.n312 6.772
R2014 VDD.n325 VDD.n322 6.772
R2015 VDD.n321 VDD.n318 6.772
R2016 VDD.n408 VDD.n393 6.772
R2017 VDD.n406 VDD.n403 6.772
R2018 VDD.n402 VDD.n399 6.772
R2019 VDD.n469 VDD.n454 6.772
R2020 VDD.n467 VDD.n464 6.772
R2021 VDD.n463 VDD.n460 6.772
R2022 VDD.n550 VDD.n535 6.772
R2023 VDD.n548 VDD.n545 6.772
R2024 VDD.n544 VDD.n541 6.772
R2025 VDD.n631 VDD.n616 6.772
R2026 VDD.n629 VDD.n626 6.772
R2027 VDD.n625 VDD.n622 6.772
R2028 VDD.n692 VDD.n677 6.772
R2029 VDD.n690 VDD.n687 6.772
R2030 VDD.n686 VDD.n683 6.772
R2031 VDD.n769 VDD.n754 6.772
R2032 VDD.n767 VDD.n764 6.772
R2033 VDD.n763 VDD.n760 6.772
R2034 VDD.n1462 VDD.n1447 6.772
R2035 VDD.n1460 VDD.n1457 6.772
R2036 VDD.n1456 VDD.n1453 6.772
R2037 VDD.n1401 VDD.n1386 6.772
R2038 VDD.n1399 VDD.n1396 6.772
R2039 VDD.n1395 VDD.n1392 6.772
R2040 VDD.n1320 VDD.n1305 6.772
R2041 VDD.n1318 VDD.n1315 6.772
R2042 VDD.n1314 VDD.n1311 6.772
R2043 VDD.n1239 VDD.n1224 6.772
R2044 VDD.n1237 VDD.n1234 6.772
R2045 VDD.n1233 VDD.n1230 6.772
R2046 VDD.n1178 VDD.n1163 6.772
R2047 VDD.n1176 VDD.n1173 6.772
R2048 VDD.n1172 VDD.n1169 6.772
R2049 VDD.n1097 VDD.n1082 6.772
R2050 VDD.n1095 VDD.n1092 6.772
R2051 VDD.n1091 VDD.n1088 6.772
R2052 VDD.n1016 VDD.n1001 6.772
R2053 VDD.n1014 VDD.n1011 6.772
R2054 VDD.n1010 VDD.n1007 6.772
R2055 VDD.n955 VDD.n940 6.772
R2056 VDD.n953 VDD.n950 6.772
R2057 VDD.n949 VDD.n946 6.772
R2058 VDD.n794 VDD.n780 6.772
R2059 VDD.n792 VDD.n789 6.772
R2060 VDD.n788 VDD.n785 6.772
R2061 VDD.n59 VDD.n58 6.772
R2062 VDD.n64 VDD.n63 6.772
R2063 VDD.n68 VDD.n67 6.772
R2064 VDD.n71 VDD.n70 6.772
R2065 VDD.n118 VDD.n117 6.772
R2066 VDD.n122 VDD.n121 6.772
R2067 VDD.n125 VDD.n124 6.772
R2068 VDD.n179 VDD.n178 6.772
R2069 VDD.n183 VDD.n182 6.772
R2070 VDD.n186 VDD.n185 6.772
R2071 VDD.n240 VDD.n239 6.772
R2072 VDD.n244 VDD.n243 6.772
R2073 VDD.n247 VDD.n246 6.772
R2074 VDD.n321 VDD.n320 6.772
R2075 VDD.n325 VDD.n324 6.772
R2076 VDD.n328 VDD.n327 6.772
R2077 VDD.n402 VDD.n401 6.772
R2078 VDD.n406 VDD.n405 6.772
R2079 VDD.n409 VDD.n408 6.772
R2080 VDD.n463 VDD.n462 6.772
R2081 VDD.n467 VDD.n466 6.772
R2082 VDD.n470 VDD.n469 6.772
R2083 VDD.n544 VDD.n543 6.772
R2084 VDD.n548 VDD.n547 6.772
R2085 VDD.n551 VDD.n550 6.772
R2086 VDD.n625 VDD.n624 6.772
R2087 VDD.n629 VDD.n628 6.772
R2088 VDD.n632 VDD.n631 6.772
R2089 VDD.n686 VDD.n685 6.772
R2090 VDD.n690 VDD.n689 6.772
R2091 VDD.n693 VDD.n692 6.772
R2092 VDD.n763 VDD.n762 6.772
R2093 VDD.n767 VDD.n766 6.772
R2094 VDD.n770 VDD.n769 6.772
R2095 VDD.n1456 VDD.n1455 6.772
R2096 VDD.n1460 VDD.n1459 6.772
R2097 VDD.n1463 VDD.n1462 6.772
R2098 VDD.n1395 VDD.n1394 6.772
R2099 VDD.n1399 VDD.n1398 6.772
R2100 VDD.n1402 VDD.n1401 6.772
R2101 VDD.n1314 VDD.n1313 6.772
R2102 VDD.n1318 VDD.n1317 6.772
R2103 VDD.n1321 VDD.n1320 6.772
R2104 VDD.n1233 VDD.n1232 6.772
R2105 VDD.n1237 VDD.n1236 6.772
R2106 VDD.n1240 VDD.n1239 6.772
R2107 VDD.n1172 VDD.n1171 6.772
R2108 VDD.n1176 VDD.n1175 6.772
R2109 VDD.n1179 VDD.n1178 6.772
R2110 VDD.n1091 VDD.n1090 6.772
R2111 VDD.n1095 VDD.n1094 6.772
R2112 VDD.n1098 VDD.n1097 6.772
R2113 VDD.n1010 VDD.n1009 6.772
R2114 VDD.n1014 VDD.n1013 6.772
R2115 VDD.n1017 VDD.n1016 6.772
R2116 VDD.n949 VDD.n948 6.772
R2117 VDD.n953 VDD.n952 6.772
R2118 VDD.n956 VDD.n955 6.772
R2119 VDD.n788 VDD.n787 6.772
R2120 VDD.n792 VDD.n791 6.772
R2121 VDD.n795 VDD.n794 6.772
R2122 VDD.n875 VDD.n874 6.772
R2123 VDD.n862 VDD.n859 6.772
R2124 VDD.n867 VDD.n864 6.772
R2125 VDD.n872 VDD.n869 6.772
R2126 VDD.n872 VDD.n871 6.772
R2127 VDD.n867 VDD.n866 6.772
R2128 VDD.n862 VDD.n861 6.772
R2129 VDD.n874 VDD.n858 6.772
R2130 VDD.n290 VDD.n286 6.69
R2131 VDD.n371 VDD.n367 6.69
R2132 VDD.n513 VDD.n509 6.69
R2133 VDD.n594 VDD.n590 6.69
R2134 VDD.n736 VDD.n732 6.69
R2135 VDD.n1490 VDD.n1486 6.69
R2136 VDD.n1348 VDD.n1344 6.69
R2137 VDD.n1267 VDD.n1263 6.69
R2138 VDD.n1125 VDD.n1121 6.69
R2139 VDD.n1044 VDD.n1040 6.69
R2140 VDD.n902 VDD.n898 6.69
R2141 VDD.n820 VDD.n816 6.69
R2142 VDD.n33 VDD.n23 6.487
R2143 VDD.n33 VDD.n32 6.475
R2144 VDD.n16 VDD.n15 6.458
R2145 VDD.n273 VDD.n272 6.296
R2146 VDD.n354 VDD.n353 6.296
R2147 VDD.n496 VDD.n495 6.296
R2148 VDD.n577 VDD.n576 6.296
R2149 VDD.n719 VDD.n718 6.296
R2150 VDD.n1507 VDD.n1506 6.296
R2151 VDD.n1365 VDD.n1364 6.296
R2152 VDD.n1284 VDD.n1283 6.296
R2153 VDD.n1142 VDD.n1141 6.296
R2154 VDD.n1061 VDD.n1060 6.296
R2155 VDD.n919 VDD.n918 6.296
R2156 VDD.n837 VDD.n836 6.296
R2157 VDD.n113 VDD.n112 6.202
R2158 VDD.n174 VDD.n173 6.202
R2159 VDD.n235 VDD.n234 6.202
R2160 VDD.n316 VDD.n315 6.202
R2161 VDD.n397 VDD.n396 6.202
R2162 VDD.n458 VDD.n457 6.202
R2163 VDD.n539 VDD.n538 6.202
R2164 VDD.n620 VDD.n619 6.202
R2165 VDD.n681 VDD.n680 6.202
R2166 VDD.n758 VDD.n757 6.202
R2167 VDD.n1451 VDD.n1450 6.202
R2168 VDD.n1390 VDD.n1389 6.202
R2169 VDD.n1309 VDD.n1308 6.202
R2170 VDD.n1228 VDD.n1227 6.202
R2171 VDD.n1167 VDD.n1166 6.202
R2172 VDD.n1086 VDD.n1085 6.202
R2173 VDD.n1005 VDD.n1004 6.202
R2174 VDD.n944 VDD.n943 6.202
R2175 VDD.n783 VDD.n782 6.202
R2176 VDD.n150 VDD.n149 4.576
R2177 VDD.n211 VDD.n210 4.576
R2178 VDD.n434 VDD.n433 4.576
R2179 VDD.n657 VDD.n656 4.576
R2180 VDD.n1421 VDD.n1420 4.576
R2181 VDD.n1198 VDD.n1197 4.576
R2182 VDD.n975 VDD.n974 4.576
R2183 VDD.n162 VDD.n159 2.754
R2184 VDD.n223 VDD.n220 2.754
R2185 VDD.n446 VDD.n443 2.754
R2186 VDD.n669 VDD.n666 2.754
R2187 VDD.n1413 VDD.n1410 2.754
R2188 VDD.n1190 VDD.n1187 2.754
R2189 VDD.n967 VDD.n964 2.754
R2190 VDD.n136 VDD.n133 2.361
R2191 VDD.n197 VDD.n194 2.361
R2192 VDD.n420 VDD.n417 2.361
R2193 VDD.n643 VDD.n640 2.361
R2194 VDD.n1439 VDD.n1436 2.361
R2195 VDD.n1216 VDD.n1213 2.361
R2196 VDD.n993 VDD.n990 2.361
R2197 VDD.n14 VDD.n7 1.329
R2198 VDD.n14 VDD.n10 1.329
R2199 VDD.n14 VDD.n12 1.329
R2200 VDD.n14 VDD.n13 1.329
R2201 VDD.n15 VDD.n14 0.696
R2202 VDD.n14 VDD.n4 0.696
R2203 VDD.n300 VDD.n297 0.393
R2204 VDD.n381 VDD.n378 0.393
R2205 VDD.n523 VDD.n520 0.393
R2206 VDD.n604 VDD.n601 0.393
R2207 VDD.n746 VDD.n743 0.393
R2208 VDD.n1478 VDD.n1475 0.393
R2209 VDD.n1336 VDD.n1333 0.393
R2210 VDD.n1255 VDD.n1252 0.393
R2211 VDD.n1113 VDD.n1110 0.393
R2212 VDD.n1032 VDD.n1029 0.393
R2213 VDD.n890 VDD.n887 0.393
R2214 VDD.n808 VDD.n805 0.393
R2215 VDD.n69 VDD.n68 0.365
R2216 VDD.n69 VDD.n64 0.365
R2217 VDD.n69 VDD.n59 0.365
R2218 VDD.n70 VDD.n69 0.365
R2219 VDD.n123 VDD.n122 0.365
R2220 VDD.n123 VDD.n118 0.365
R2221 VDD.n124 VDD.n123 0.365
R2222 VDD.n184 VDD.n183 0.365
R2223 VDD.n184 VDD.n179 0.365
R2224 VDD.n185 VDD.n184 0.365
R2225 VDD.n245 VDD.n244 0.365
R2226 VDD.n245 VDD.n240 0.365
R2227 VDD.n246 VDD.n245 0.365
R2228 VDD.n326 VDD.n325 0.365
R2229 VDD.n326 VDD.n321 0.365
R2230 VDD.n327 VDD.n326 0.365
R2231 VDD.n407 VDD.n406 0.365
R2232 VDD.n407 VDD.n402 0.365
R2233 VDD.n408 VDD.n407 0.365
R2234 VDD.n468 VDD.n467 0.365
R2235 VDD.n468 VDD.n463 0.365
R2236 VDD.n469 VDD.n468 0.365
R2237 VDD.n549 VDD.n548 0.365
R2238 VDD.n549 VDD.n544 0.365
R2239 VDD.n550 VDD.n549 0.365
R2240 VDD.n630 VDD.n629 0.365
R2241 VDD.n630 VDD.n625 0.365
R2242 VDD.n631 VDD.n630 0.365
R2243 VDD.n691 VDD.n690 0.365
R2244 VDD.n691 VDD.n686 0.365
R2245 VDD.n692 VDD.n691 0.365
R2246 VDD.n768 VDD.n767 0.365
R2247 VDD.n768 VDD.n763 0.365
R2248 VDD.n769 VDD.n768 0.365
R2249 VDD.n1461 VDD.n1460 0.365
R2250 VDD.n1461 VDD.n1456 0.365
R2251 VDD.n1462 VDD.n1461 0.365
R2252 VDD.n1400 VDD.n1399 0.365
R2253 VDD.n1400 VDD.n1395 0.365
R2254 VDD.n1401 VDD.n1400 0.365
R2255 VDD.n1319 VDD.n1318 0.365
R2256 VDD.n1319 VDD.n1314 0.365
R2257 VDD.n1320 VDD.n1319 0.365
R2258 VDD.n1238 VDD.n1237 0.365
R2259 VDD.n1238 VDD.n1233 0.365
R2260 VDD.n1239 VDD.n1238 0.365
R2261 VDD.n1177 VDD.n1176 0.365
R2262 VDD.n1177 VDD.n1172 0.365
R2263 VDD.n1178 VDD.n1177 0.365
R2264 VDD.n1096 VDD.n1095 0.365
R2265 VDD.n1096 VDD.n1091 0.365
R2266 VDD.n1097 VDD.n1096 0.365
R2267 VDD.n1015 VDD.n1014 0.365
R2268 VDD.n1015 VDD.n1010 0.365
R2269 VDD.n1016 VDD.n1015 0.365
R2270 VDD.n954 VDD.n953 0.365
R2271 VDD.n954 VDD.n949 0.365
R2272 VDD.n955 VDD.n954 0.365
R2273 VDD.n793 VDD.n792 0.365
R2274 VDD.n793 VDD.n788 0.365
R2275 VDD.n794 VDD.n793 0.365
R2276 VDD.n873 VDD.n872 0.365
R2277 VDD.n873 VDD.n867 0.365
R2278 VDD.n873 VDD.n862 0.365
R2279 VDD.n874 VDD.n873 0.365
R2280 VDD.n78 VDD.n51 0.29
R2281 VDD.n132 VDD.n106 0.29
R2282 VDD.n193 VDD.n167 0.29
R2283 VDD.n254 VDD.n228 0.29
R2284 VDD.n335 VDD.n309 0.29
R2285 VDD.n416 VDD.n390 0.29
R2286 VDD.n477 VDD.n451 0.29
R2287 VDD.n558 VDD.n532 0.29
R2288 VDD.n639 VDD.n613 0.29
R2289 VDD.n700 VDD.n674 0.29
R2290 VDD.n1470 VDD.n1444 0.29
R2291 VDD.n1409 VDD.n1383 0.29
R2292 VDD.n1328 VDD.n1302 0.29
R2293 VDD.n1247 VDD.n1221 0.29
R2294 VDD.n1186 VDD.n1160 0.29
R2295 VDD.n1105 VDD.n1079 0.29
R2296 VDD.n1024 VDD.n998 0.29
R2297 VDD.n963 VDD.n937 0.29
R2298 VDD.n882 VDD.n855 0.29
R2299 VDD VDD.n1525 0.219
R2300 VDD.n800 VDD 0.207
R2301 VDD.n284 VDD.n279 0.197
R2302 VDD.n365 VDD.n360 0.197
R2303 VDD.n507 VDD.n502 0.197
R2304 VDD.n588 VDD.n583 0.197
R2305 VDD.n730 VDD.n725 0.197
R2306 VDD.n1501 VDD.n1496 0.197
R2307 VDD.n1359 VDD.n1354 0.197
R2308 VDD.n1278 VDD.n1273 0.197
R2309 VDD.n1136 VDD.n1131 0.197
R2310 VDD.n1055 VDD.n1050 0.197
R2311 VDD.n913 VDD.n908 0.197
R2312 VDD.n831 VDD.n826 0.197
R2313 VDD.n39 VDD.n35 0.181
R2314 VDD.n94 VDD.n90 0.181
R2315 VDD.n153 VDD.n148 0.181
R2316 VDD.n214 VDD.n209 0.181
R2317 VDD.n437 VDD.n432 0.181
R2318 VDD.n660 VDD.n655 0.181
R2319 VDD.n1430 VDD.n1424 0.181
R2320 VDD.n1207 VDD.n1201 0.181
R2321 VDD.n984 VDD.n978 0.181
R2322 VDD.n35 VDD.n34 0.145
R2323 VDD.n43 VDD.n39 0.145
R2324 VDD.n47 VDD.n43 0.145
R2325 VDD.n51 VDD.n47 0.145
R2326 VDD.n82 VDD.n78 0.145
R2327 VDD.n86 VDD.n82 0.145
R2328 VDD.n90 VDD.n86 0.145
R2329 VDD.n98 VDD.n94 0.145
R2330 VDD.n102 VDD.n98 0.145
R2331 VDD.n106 VDD.n102 0.145
R2332 VDD.n137 VDD.n132 0.145
R2333 VDD.n142 VDD.n137 0.145
R2334 VDD.n148 VDD.n142 0.145
R2335 VDD.n158 VDD.n153 0.145
R2336 VDD.n163 VDD.n158 0.145
R2337 VDD.n167 VDD.n163 0.145
R2338 VDD.n198 VDD.n193 0.145
R2339 VDD.n203 VDD.n198 0.145
R2340 VDD.n209 VDD.n203 0.145
R2341 VDD.n219 VDD.n214 0.145
R2342 VDD.n224 VDD.n219 0.145
R2343 VDD.n228 VDD.n224 0.145
R2344 VDD.n258 VDD.n254 0.145
R2345 VDD.n262 VDD.n258 0.145
R2346 VDD.n267 VDD.n262 0.145
R2347 VDD.n274 VDD.n267 0.145
R2348 VDD.n279 VDD.n274 0.145
R2349 VDD.n291 VDD.n284 0.145
R2350 VDD.n296 VDD.n291 0.145
R2351 VDD.n301 VDD.n296 0.145
R2352 VDD.n305 VDD.n301 0.145
R2353 VDD.n309 VDD.n305 0.145
R2354 VDD.n339 VDD.n335 0.145
R2355 VDD.n343 VDD.n339 0.145
R2356 VDD.n348 VDD.n343 0.145
R2357 VDD.n355 VDD.n348 0.145
R2358 VDD.n360 VDD.n355 0.145
R2359 VDD.n372 VDD.n365 0.145
R2360 VDD.n377 VDD.n372 0.145
R2361 VDD.n382 VDD.n377 0.145
R2362 VDD.n386 VDD.n382 0.145
R2363 VDD.n390 VDD.n386 0.145
R2364 VDD.n421 VDD.n416 0.145
R2365 VDD.n426 VDD.n421 0.145
R2366 VDD.n432 VDD.n426 0.145
R2367 VDD.n442 VDD.n437 0.145
R2368 VDD.n447 VDD.n442 0.145
R2369 VDD.n451 VDD.n447 0.145
R2370 VDD.n481 VDD.n477 0.145
R2371 VDD.n485 VDD.n481 0.145
R2372 VDD.n490 VDD.n485 0.145
R2373 VDD.n497 VDD.n490 0.145
R2374 VDD.n502 VDD.n497 0.145
R2375 VDD.n514 VDD.n507 0.145
R2376 VDD.n519 VDD.n514 0.145
R2377 VDD.n524 VDD.n519 0.145
R2378 VDD.n528 VDD.n524 0.145
R2379 VDD.n532 VDD.n528 0.145
R2380 VDD.n562 VDD.n558 0.145
R2381 VDD.n566 VDD.n562 0.145
R2382 VDD.n571 VDD.n566 0.145
R2383 VDD.n578 VDD.n571 0.145
R2384 VDD.n583 VDD.n578 0.145
R2385 VDD.n595 VDD.n588 0.145
R2386 VDD.n600 VDD.n595 0.145
R2387 VDD.n605 VDD.n600 0.145
R2388 VDD.n609 VDD.n605 0.145
R2389 VDD.n613 VDD.n609 0.145
R2390 VDD.n644 VDD.n639 0.145
R2391 VDD.n649 VDD.n644 0.145
R2392 VDD.n655 VDD.n649 0.145
R2393 VDD.n665 VDD.n660 0.145
R2394 VDD.n670 VDD.n665 0.145
R2395 VDD.n674 VDD.n670 0.145
R2396 VDD.n704 VDD.n700 0.145
R2397 VDD.n708 VDD.n704 0.145
R2398 VDD.n713 VDD.n708 0.145
R2399 VDD.n720 VDD.n713 0.145
R2400 VDD.n725 VDD.n720 0.145
R2401 VDD.n737 VDD.n730 0.145
R2402 VDD.n742 VDD.n737 0.145
R2403 VDD.n747 VDD.n742 0.145
R2404 VDD.n751 VDD.n747 0.145
R2405 VDD.n777 VDD.n751 0.145
R2406 VDD.n1525 VDD.n1521 0.145
R2407 VDD.n1521 VDD.n1517 0.145
R2408 VDD.n1517 VDD.n1513 0.145
R2409 VDD.n1513 VDD.n1508 0.145
R2410 VDD.n1508 VDD.n1501 0.145
R2411 VDD.n1496 VDD.n1491 0.145
R2412 VDD.n1491 VDD.n1484 0.145
R2413 VDD.n1484 VDD.n1479 0.145
R2414 VDD.n1479 VDD.n1474 0.145
R2415 VDD.n1474 VDD.n1470 0.145
R2416 VDD.n1444 VDD.n1440 0.145
R2417 VDD.n1440 VDD.n1435 0.145
R2418 VDD.n1435 VDD.n1430 0.145
R2419 VDD.n1424 VDD.n1419 0.145
R2420 VDD.n1419 VDD.n1414 0.145
R2421 VDD.n1414 VDD.n1409 0.145
R2422 VDD.n1383 VDD.n1379 0.145
R2423 VDD.n1379 VDD.n1375 0.145
R2424 VDD.n1375 VDD.n1371 0.145
R2425 VDD.n1371 VDD.n1366 0.145
R2426 VDD.n1366 VDD.n1359 0.145
R2427 VDD.n1354 VDD.n1349 0.145
R2428 VDD.n1349 VDD.n1342 0.145
R2429 VDD.n1342 VDD.n1337 0.145
R2430 VDD.n1337 VDD.n1332 0.145
R2431 VDD.n1332 VDD.n1328 0.145
R2432 VDD.n1302 VDD.n1298 0.145
R2433 VDD.n1298 VDD.n1294 0.145
R2434 VDD.n1294 VDD.n1290 0.145
R2435 VDD.n1290 VDD.n1285 0.145
R2436 VDD.n1285 VDD.n1278 0.145
R2437 VDD.n1273 VDD.n1268 0.145
R2438 VDD.n1268 VDD.n1261 0.145
R2439 VDD.n1261 VDD.n1256 0.145
R2440 VDD.n1256 VDD.n1251 0.145
R2441 VDD.n1251 VDD.n1247 0.145
R2442 VDD.n1221 VDD.n1217 0.145
R2443 VDD.n1217 VDD.n1212 0.145
R2444 VDD.n1212 VDD.n1207 0.145
R2445 VDD.n1201 VDD.n1196 0.145
R2446 VDD.n1196 VDD.n1191 0.145
R2447 VDD.n1191 VDD.n1186 0.145
R2448 VDD.n1160 VDD.n1156 0.145
R2449 VDD.n1156 VDD.n1152 0.145
R2450 VDD.n1152 VDD.n1148 0.145
R2451 VDD.n1148 VDD.n1143 0.145
R2452 VDD.n1143 VDD.n1136 0.145
R2453 VDD.n1131 VDD.n1126 0.145
R2454 VDD.n1126 VDD.n1119 0.145
R2455 VDD.n1119 VDD.n1114 0.145
R2456 VDD.n1114 VDD.n1109 0.145
R2457 VDD.n1109 VDD.n1105 0.145
R2458 VDD.n1079 VDD.n1075 0.145
R2459 VDD.n1075 VDD.n1071 0.145
R2460 VDD.n1071 VDD.n1067 0.145
R2461 VDD.n1067 VDD.n1062 0.145
R2462 VDD.n1062 VDD.n1055 0.145
R2463 VDD.n1050 VDD.n1045 0.145
R2464 VDD.n1045 VDD.n1038 0.145
R2465 VDD.n1038 VDD.n1033 0.145
R2466 VDD.n1033 VDD.n1028 0.145
R2467 VDD.n1028 VDD.n1024 0.145
R2468 VDD.n998 VDD.n994 0.145
R2469 VDD.n994 VDD.n989 0.145
R2470 VDD.n989 VDD.n984 0.145
R2471 VDD.n978 VDD.n973 0.145
R2472 VDD.n973 VDD.n968 0.145
R2473 VDD.n968 VDD.n963 0.145
R2474 VDD.n937 VDD.n933 0.145
R2475 VDD.n933 VDD.n929 0.145
R2476 VDD.n929 VDD.n925 0.145
R2477 VDD.n925 VDD.n920 0.145
R2478 VDD.n920 VDD.n913 0.145
R2479 VDD.n908 VDD.n903 0.145
R2480 VDD.n903 VDD.n896 0.145
R2481 VDD.n896 VDD.n891 0.145
R2482 VDD.n891 VDD.n886 0.145
R2483 VDD.n886 VDD.n882 0.145
R2484 VDD.n855 VDD.n851 0.145
R2485 VDD.n851 VDD.n847 0.145
R2486 VDD.n847 VDD.n843 0.145
R2487 VDD.n843 VDD.n838 0.145
R2488 VDD.n838 VDD.n831 0.145
R2489 VDD.n826 VDD.n821 0.145
R2490 VDD.n821 VDD.n814 0.145
R2491 VDD.n814 VDD.n809 0.145
R2492 VDD.n809 VDD.n804 0.145
R2493 VDD.n804 VDD.n800 0.145
R2494 VDD VDD.n777 0.07
R2495 a_5779_989.n0 a_5779_989.t12 480.392
R2496 a_5779_989.n2 a_5779_989.t7 454.685
R2497 a_5779_989.n2 a_5779_989.t11 428.979
R2498 a_5779_989.n0 a_5779_989.t10 403.272
R2499 a_5779_989.n1 a_5779_989.t9 283.48
R2500 a_5779_989.n3 a_5779_989.t8 237.959
R2501 a_5779_989.n9 a_5779_989.n8 213.104
R2502 a_5779_989.n13 a_5779_989.n9 170.799
R2503 a_5779_989.n3 a_5779_989.n2 98.447
R2504 a_5779_989.n1 a_5779_989.n0 98.447
R2505 a_5779_989.n4 a_5779_989.n3 80.035
R2506 a_5779_989.n12 a_5779_989.n11 79.232
R2507 a_5779_989.n4 a_5779_989.n1 77.315
R2508 a_5779_989.n9 a_5779_989.n4 76
R2509 a_5779_989.n13 a_5779_989.n12 63.152
R2510 a_5779_989.n8 a_5779_989.n7 30
R2511 a_5779_989.n6 a_5779_989.n5 24.383
R2512 a_5779_989.n8 a_5779_989.n6 23.684
R2513 a_5779_989.n12 a_5779_989.n10 16.08
R2514 a_5779_989.n14 a_5779_989.n13 16.078
R2515 a_5779_989.n10 a_5779_989.t3 14.282
R2516 a_5779_989.n10 a_5779_989.t4 14.282
R2517 a_5779_989.n11 a_5779_989.t6 14.282
R2518 a_5779_989.n11 a_5779_989.t5 14.282
R2519 a_5779_989.n14 a_5779_989.t0 14.282
R2520 a_5779_989.t1 a_5779_989.n14 14.282
R2521 a_9331_989.n5 a_9331_989.t13 512.525
R2522 a_9331_989.n3 a_9331_989.t6 477.179
R2523 a_9331_989.n8 a_9331_989.t5 454.685
R2524 a_9331_989.n8 a_9331_989.t8 428.979
R2525 a_9331_989.n3 a_9331_989.t11 406.485
R2526 a_9331_989.n5 a_9331_989.t9 371.139
R2527 a_9331_989.n4 a_9331_989.t7 363.924
R2528 a_9331_989.n7 a_9331_989.t10 250.5
R2529 a_9331_989.n9 a_9331_989.t12 211.406
R2530 a_9331_989.n13 a_9331_989.n11 190.561
R2531 a_9331_989.n11 a_9331_989.n2 179.052
R2532 a_9331_989.n9 a_9331_989.n8 125
R2533 a_9331_989.n7 a_9331_989.n6 106.997
R2534 a_9331_989.n6 a_9331_989.n4 101.359
R2535 a_9331_989.n10 a_9331_989.n7 96.087
R2536 a_9331_989.n10 a_9331_989.n9 78.947
R2537 a_9331_989.n2 a_9331_989.n1 76.002
R2538 a_9331_989.n11 a_9331_989.n10 76
R2539 a_9331_989.n6 a_9331_989.n5 71.88
R2540 a_9331_989.n4 a_9331_989.n3 15.776
R2541 a_9331_989.n13 a_9331_989.n12 15.218
R2542 a_9331_989.n0 a_9331_989.t3 14.282
R2543 a_9331_989.n0 a_9331_989.t2 14.282
R2544 a_9331_989.n1 a_9331_989.t0 14.282
R2545 a_9331_989.n1 a_9331_989.t4 14.282
R2546 a_9331_989.n2 a_9331_989.n0 12.85
R2547 a_9331_989.n14 a_9331_989.n13 12.014
R2548 a_9009_1050.n1 a_9009_1050.t9 480.392
R2549 a_9009_1050.n1 a_9009_1050.t7 403.272
R2550 a_9009_1050.n2 a_9009_1050.t8 310.033
R2551 a_9009_1050.n7 a_9009_1050.n6 239.657
R2552 a_9009_1050.n7 a_9009_1050.n2 153.315
R2553 a_9009_1050.n8 a_9009_1050.n7 144.246
R2554 a_9009_1050.n10 a_9009_1050.n9 79.232
R2555 a_9009_1050.n2 a_9009_1050.n1 71.894
R2556 a_9009_1050.n10 a_9009_1050.n8 63.152
R2557 a_9009_1050.n6 a_9009_1050.n5 30
R2558 a_9009_1050.n4 a_9009_1050.n3 24.383
R2559 a_9009_1050.n6 a_9009_1050.n4 23.684
R2560 a_9009_1050.n8 a_9009_1050.n0 16.08
R2561 a_9009_1050.n11 a_9009_1050.n10 16.078
R2562 a_9009_1050.n0 a_9009_1050.t3 14.282
R2563 a_9009_1050.n0 a_9009_1050.t4 14.282
R2564 a_9009_1050.n9 a_9009_1050.t6 14.282
R2565 a_9009_1050.n9 a_9009_1050.t5 14.282
R2566 a_9009_1050.t1 a_9009_1050.n11 14.282
R2567 a_9009_1050.n11 a_9009_1050.t0 14.282
R2568 a_147_187.n4 a_147_187.t9 512.525
R2569 a_147_187.n2 a_147_187.t11 472.359
R2570 a_147_187.n0 a_147_187.t8 472.359
R2571 a_147_187.n2 a_147_187.t14 384.527
R2572 a_147_187.n0 a_147_187.t12 384.527
R2573 a_147_187.n4 a_147_187.t13 371.139
R2574 a_147_187.n5 a_147_187.t10 340.774
R2575 a_147_187.n3 a_147_187.t7 294.278
R2576 a_147_187.n1 a_147_187.t15 294.278
R2577 a_147_187.n12 a_147_187.n11 266.21
R2578 a_147_187.n16 a_147_187.n12 117.693
R2579 a_147_187.n5 a_147_187.n4 109.607
R2580 a_147_187.n6 a_147_187.n5 83.572
R2581 a_147_187.n7 a_147_187.n1 81.396
R2582 a_147_187.n15 a_147_187.n14 79.232
R2583 a_147_187.n6 a_147_187.n3 76
R2584 a_147_187.n12 a_147_187.n7 76
R2585 a_147_187.n16 a_147_187.n15 63.152
R2586 a_147_187.n3 a_147_187.n2 56.954
R2587 a_147_187.n1 a_147_187.n0 56.954
R2588 a_147_187.n11 a_147_187.n10 30
R2589 a_147_187.n9 a_147_187.n8 24.383
R2590 a_147_187.n11 a_147_187.n9 23.684
R2591 a_147_187.n15 a_147_187.n13 16.08
R2592 a_147_187.n17 a_147_187.n16 16.078
R2593 a_147_187.n13 a_147_187.t3 14.282
R2594 a_147_187.n13 a_147_187.t5 14.282
R2595 a_147_187.n14 a_147_187.t4 14.282
R2596 a_147_187.n14 a_147_187.t6 14.282
R2597 a_147_187.t1 a_147_187.n17 14.282
R2598 a_147_187.n17 a_147_187.t0 14.282
R2599 a_147_187.n7 a_147_187.n6 4.035
R2600 a_2036_101.t0 a_2036_101.n1 34.62
R2601 a_2036_101.t0 a_2036_101.n0 8.137
R2602 a_2036_101.t0 a_2036_101.n2 4.69
R2603 a_2141_1050.n0 a_2141_1050.t5 512.525
R2604 a_2141_1050.n0 a_2141_1050.t7 371.139
R2605 a_2141_1050.n1 a_2141_1050.t6 287.668
R2606 a_2141_1050.n3 a_2141_1050.n2 232.331
R2607 a_2141_1050.n1 a_2141_1050.n0 162.713
R2608 a_2141_1050.n3 a_2141_1050.n1 153.315
R2609 a_2141_1050.n5 a_2141_1050.n3 152.499
R2610 a_2141_1050.n5 a_2141_1050.n4 76.002
R2611 a_2141_1050.n4 a_2141_1050.t4 14.282
R2612 a_2141_1050.n4 a_2141_1050.t3 14.282
R2613 a_2141_1050.t1 a_2141_1050.n6 14.282
R2614 a_2141_1050.n6 a_2141_1050.t0 14.282
R2615 a_2141_1050.n6 a_2141_1050.n5 12.848
R2616 CLK.n14 CLK.t4 459.505
R2617 CLK.n11 CLK.t17 459.505
R2618 CLK.n8 CLK.t16 459.505
R2619 CLK.n5 CLK.t15 459.505
R2620 CLK.n2 CLK.t6 459.505
R2621 CLK.n0 CLK.t5 459.505
R2622 CLK.n14 CLK.t11 384.527
R2623 CLK.n11 CLK.t7 384.527
R2624 CLK.n8 CLK.t0 384.527
R2625 CLK.n5 CLK.t3 384.527
R2626 CLK.n2 CLK.t13 384.527
R2627 CLK.n0 CLK.t12 384.527
R2628 CLK.n15 CLK.t8 322.152
R2629 CLK.n12 CLK.t14 322.151
R2630 CLK.n9 CLK.t9 322.151
R2631 CLK.n6 CLK.t2 322.151
R2632 CLK.n3 CLK.t1 322.151
R2633 CLK.n1 CLK.t10 322.151
R2634 CLK.n4 CLK.n1 58.818
R2635 CLK.n16 CLK.n15 49.342
R2636 CLK.n4 CLK.n3 49.342
R2637 CLK.n7 CLK.n6 49.342
R2638 CLK.n10 CLK.n9 49.342
R2639 CLK.n13 CLK.n12 49.342
R2640 CLK.n15 CLK.n14 27.599
R2641 CLK.n1 CLK.n0 27.599
R2642 CLK.n3 CLK.n2 27.599
R2643 CLK.n6 CLK.n5 27.599
R2644 CLK.n9 CLK.n8 27.599
R2645 CLK.n12 CLK.n11 27.599
R2646 CLK.n7 CLK.n4 9.476
R2647 CLK.n10 CLK.n7 9.476
R2648 CLK.n13 CLK.n10 9.476
R2649 CLK.n16 CLK.n13 9.476
R2650 CLK.n16 CLK 0.046
R2651 a_5457_1050.n3 a_5457_1050.t9 512.525
R2652 a_5457_1050.n1 a_5457_1050.t10 512.525
R2653 a_5457_1050.n3 a_5457_1050.t12 371.139
R2654 a_5457_1050.n1 a_5457_1050.t11 371.139
R2655 a_5457_1050.n4 a_5457_1050.t8 314.221
R2656 a_5457_1050.n2 a_5457_1050.t7 314.221
R2657 a_5457_1050.n10 a_5457_1050.n9 239.657
R2658 a_5457_1050.n11 a_5457_1050.n10 144.246
R2659 a_5457_1050.n4 a_5457_1050.n3 136.16
R2660 a_5457_1050.n2 a_5457_1050.n1 136.16
R2661 a_5457_1050.n5 a_5457_1050.n2 85.476
R2662 a_5457_1050.n13 a_5457_1050.n12 79.232
R2663 a_5457_1050.n10 a_5457_1050.n5 77.315
R2664 a_5457_1050.n5 a_5457_1050.n4 76
R2665 a_5457_1050.n13 a_5457_1050.n11 63.152
R2666 a_5457_1050.n9 a_5457_1050.n8 30
R2667 a_5457_1050.n7 a_5457_1050.n6 24.383
R2668 a_5457_1050.n9 a_5457_1050.n7 23.684
R2669 a_5457_1050.n11 a_5457_1050.n0 16.08
R2670 a_5457_1050.n14 a_5457_1050.n13 16.078
R2671 a_5457_1050.n0 a_5457_1050.t2 14.282
R2672 a_5457_1050.n0 a_5457_1050.t3 14.282
R2673 a_5457_1050.n12 a_5457_1050.t6 14.282
R2674 a_5457_1050.n12 a_5457_1050.t5 14.282
R2675 a_5457_1050.n14 a_5457_1050.t0 14.282
R2676 a_5457_1050.t1 a_5457_1050.n14 14.282
R2677 a_10507_187.n5 a_10507_187.t9 512.525
R2678 a_10507_187.n3 a_10507_187.t13 472.359
R2679 a_10507_187.n1 a_10507_187.t12 472.359
R2680 a_10507_187.n3 a_10507_187.t15 384.527
R2681 a_10507_187.n1 a_10507_187.t14 384.527
R2682 a_10507_187.n5 a_10507_187.t10 371.139
R2683 a_10507_187.n6 a_10507_187.t7 340.774
R2684 a_10507_187.n4 a_10507_187.t11 294.278
R2685 a_10507_187.n2 a_10507_187.t8 294.278
R2686 a_10507_187.n13 a_10507_187.n12 266.21
R2687 a_10507_187.n14 a_10507_187.n13 117.693
R2688 a_10507_187.n6 a_10507_187.n5 109.607
R2689 a_10507_187.n7 a_10507_187.n6 83.572
R2690 a_10507_187.n8 a_10507_187.n2 81.396
R2691 a_10507_187.n16 a_10507_187.n15 79.232
R2692 a_10507_187.n7 a_10507_187.n4 76
R2693 a_10507_187.n13 a_10507_187.n8 76
R2694 a_10507_187.n16 a_10507_187.n14 63.152
R2695 a_10507_187.n4 a_10507_187.n3 56.954
R2696 a_10507_187.n2 a_10507_187.n1 56.954
R2697 a_10507_187.n12 a_10507_187.n11 30
R2698 a_10507_187.n10 a_10507_187.n9 24.383
R2699 a_10507_187.n12 a_10507_187.n10 23.684
R2700 a_10507_187.n14 a_10507_187.n0 16.08
R2701 a_10507_187.n17 a_10507_187.n16 16.078
R2702 a_10507_187.n0 a_10507_187.t4 14.282
R2703 a_10507_187.n0 a_10507_187.t3 14.282
R2704 a_10507_187.n15 a_10507_187.t2 14.282
R2705 a_10507_187.n15 a_10507_187.t6 14.282
R2706 a_10507_187.t1 a_10507_187.n17 14.282
R2707 a_10507_187.n17 a_10507_187.t0 14.282
R2708 a_10507_187.n8 a_10507_187.n7 4.035
R2709 a_10451_103.n1 a_10451_103.n0 25.576
R2710 a_10451_103.n3 a_10451_103.n2 9.111
R2711 a_10451_103.n7 a_10451_103.n5 7.859
R2712 a_10451_103.t0 a_10451_103.n7 3.034
R2713 a_10451_103.n5 a_10451_103.n3 1.964
R2714 a_10451_103.n5 a_10451_103.n4 1.964
R2715 a_10451_103.t0 a_10451_103.n1 1.871
R2716 a_10451_103.n7 a_10451_103.n6 0.443
R2717 a_16421_1051.n4 a_16421_1051.n3 196.002
R2718 a_16421_1051.t0 a_16421_1051.n5 89.556
R2719 a_16421_1051.n3 a_16421_1051.n2 75.271
R2720 a_16421_1051.n5 a_16421_1051.n4 75.214
R2721 a_16421_1051.n3 a_16421_1051.n1 36.52
R2722 a_16421_1051.n4 a_16421_1051.t6 14.338
R2723 a_16421_1051.n1 a_16421_1051.t7 14.282
R2724 a_16421_1051.n1 a_16421_1051.t4 14.282
R2725 a_16421_1051.n2 a_16421_1051.t3 14.282
R2726 a_16421_1051.n2 a_16421_1051.t2 14.282
R2727 a_16421_1051.n0 a_16421_1051.t5 14.282
R2728 a_16421_1051.n0 a_16421_1051.t1 14.282
R2729 a_16421_1051.n5 a_16421_1051.n0 12.119
R2730 a_15757_1051.n4 a_15757_1051.n3 195.987
R2731 a_15757_1051.n2 a_15757_1051.t7 89.553
R2732 a_15757_1051.n5 a_15757_1051.n4 75.27
R2733 a_15757_1051.n3 a_15757_1051.n2 75.214
R2734 a_15757_1051.n4 a_15757_1051.n0 36.519
R2735 a_15757_1051.n3 a_15757_1051.t3 14.338
R2736 a_15757_1051.n0 a_15757_1051.t0 14.282
R2737 a_15757_1051.n0 a_15757_1051.t6 14.282
R2738 a_15757_1051.n1 a_15757_1051.t5 14.282
R2739 a_15757_1051.n1 a_15757_1051.t4 14.282
R2740 a_15757_1051.n5 a_15757_1051.t1 14.282
R2741 a_15757_1051.t2 a_15757_1051.n5 14.282
R2742 a_15757_1051.n2 a_15757_1051.n1 12.119
R2743 a_14511_989.n1 a_14511_989.t7 475.572
R2744 a_14511_989.n0 a_14511_989.t9 469.145
R2745 a_14511_989.n5 a_14511_989.t11 454.685
R2746 a_14511_989.n5 a_14511_989.t5 428.979
R2747 a_14511_989.n1 a_14511_989.t13 384.527
R2748 a_14511_989.n0 a_14511_989.t12 384.527
R2749 a_14511_989.n2 a_14511_989.t8 294.278
R2750 a_14511_989.n4 a_14511_989.t6 241.172
R2751 a_14511_989.n6 a_14511_989.t10 237.959
R2752 a_14511_989.n12 a_14511_989.n11 210.592
R2753 a_14511_989.n3 a_14511_989.n2 156.851
R2754 a_14511_989.n14 a_14511_989.n12 152.499
R2755 a_14511_989.n6 a_14511_989.n5 98.447
R2756 a_14511_989.n7 a_14511_989.n6 78.947
R2757 a_14511_989.n7 a_14511_989.n4 77.859
R2758 a_14511_989.n14 a_14511_989.n13 76.002
R2759 a_14511_989.n12 a_14511_989.n7 76
R2760 a_14511_989.n2 a_14511_989.n1 57.842
R2761 a_14511_989.n3 a_14511_989.n0 56.833
R2762 a_14511_989.n4 a_14511_989.n3 53.105
R2763 a_14511_989.n11 a_14511_989.n10 30
R2764 a_14511_989.n9 a_14511_989.n8 24.383
R2765 a_14511_989.n11 a_14511_989.n9 23.684
R2766 a_14511_989.n13 a_14511_989.t3 14.282
R2767 a_14511_989.n13 a_14511_989.t4 14.282
R2768 a_14511_989.t1 a_14511_989.n15 14.282
R2769 a_14511_989.n15 a_14511_989.t0 14.282
R2770 a_14511_989.n15 a_14511_989.n14 12.848
R2771 a_14189_1050.n1 a_14189_1050.t8 480.392
R2772 a_14189_1050.n1 a_14189_1050.t7 403.272
R2773 a_14189_1050.n2 a_14189_1050.t9 310.033
R2774 a_14189_1050.n7 a_14189_1050.n6 239.657
R2775 a_14189_1050.n7 a_14189_1050.n2 153.315
R2776 a_14189_1050.n8 a_14189_1050.n7 144.246
R2777 a_14189_1050.n10 a_14189_1050.n9 79.232
R2778 a_14189_1050.n2 a_14189_1050.n1 71.894
R2779 a_14189_1050.n10 a_14189_1050.n8 63.152
R2780 a_14189_1050.n6 a_14189_1050.n5 30
R2781 a_14189_1050.n4 a_14189_1050.n3 24.383
R2782 a_14189_1050.n6 a_14189_1050.n4 23.684
R2783 a_14189_1050.n8 a_14189_1050.n0 16.08
R2784 a_14189_1050.n11 a_14189_1050.n10 16.078
R2785 a_14189_1050.n0 a_14189_1050.t3 14.282
R2786 a_14189_1050.n0 a_14189_1050.t2 14.282
R2787 a_14189_1050.n9 a_14189_1050.t6 14.282
R2788 a_14189_1050.n9 a_14189_1050.t5 14.282
R2789 a_14189_1050.n11 a_14189_1050.t0 14.282
R2790 a_14189_1050.t1 a_14189_1050.n11 14.282
R2791 a_15652_101.n1 a_15652_101.n0 32.249
R2792 a_15652_101.t0 a_15652_101.n5 7.911
R2793 a_15652_101.n4 a_15652_101.n2 4.032
R2794 a_15652_101.n4 a_15652_101.n3 3.644
R2795 a_15652_101.t0 a_15652_101.n1 2.534
R2796 a_15652_101.t0 a_15652_101.n4 1.099
R2797 QN.n12 QN.n11 216.728
R2798 QN.n12 QN.n2 126.664
R2799 QN.n7 QN.n6 120.24
R2800 QN.n7 QN.n5 111.94
R2801 QN.n10 QN.n8 80.526
R2802 QN.n11 QN.n7 78.403
R2803 QN.n13 QN.n12 76
R2804 QN.n2 QN.n1 75.271
R2805 QN.n10 QN.n9 30
R2806 QN.n5 QN.n4 22.578
R2807 QN.n11 QN.n10 20.417
R2808 QN.n0 QN.t4 14.282
R2809 QN.n0 QN.t3 14.282
R2810 QN.n1 QN.t0 14.282
R2811 QN.n1 QN.t5 14.282
R2812 QN.n2 QN.n0 12.119
R2813 QN.n5 QN.n3 8.58
R2814 QN.n13 QN 0.046
R2815 a_6514_210.n10 a_6514_210.n8 82.852
R2816 a_6514_210.n11 a_6514_210.n0 49.6
R2817 a_6514_210.n7 a_6514_210.n6 32.833
R2818 a_6514_210.n8 a_6514_210.t1 32.416
R2819 a_6514_210.n10 a_6514_210.n9 27.2
R2820 a_6514_210.n3 a_6514_210.n2 23.284
R2821 a_6514_210.n11 a_6514_210.n10 22.4
R2822 a_6514_210.n7 a_6514_210.n4 19.017
R2823 a_6514_210.n6 a_6514_210.n5 13.494
R2824 a_6514_210.t1 a_6514_210.n1 7.04
R2825 a_6514_210.t1 a_6514_210.n3 5.727
R2826 a_6514_210.n8 a_6514_210.n7 1.435
R2827 a_4151_989.n1 a_4151_989.t5 512.525
R2828 a_4151_989.n0 a_4151_989.t11 512.525
R2829 a_4151_989.n5 a_4151_989.t7 454.685
R2830 a_4151_989.n5 a_4151_989.t12 428.979
R2831 a_4151_989.n1 a_4151_989.t9 371.139
R2832 a_4151_989.n0 a_4151_989.t6 371.139
R2833 a_4151_989.n2 a_4151_989.n1 265.439
R2834 a_4151_989.n4 a_4151_989.n0 212.333
R2835 a_4151_989.n14 a_4151_989.n12 205.605
R2836 a_4151_989.n2 a_4151_989.t13 176.995
R2837 a_4151_989.n6 a_4151_989.t8 173.606
R2838 a_4151_989.n3 a_4151_989.t10 170.569
R2839 a_4151_989.n12 a_4151_989.n11 157.486
R2840 a_4151_989.n3 a_4151_989.n2 153.043
R2841 a_4151_989.n6 a_4151_989.n5 151.553
R2842 a_4151_989.n7 a_4151_989.n4 118.94
R2843 a_4151_989.n7 a_4151_989.n6 78.947
R2844 a_4151_989.n14 a_4151_989.n13 76.002
R2845 a_4151_989.n12 a_4151_989.n7 76
R2846 a_4151_989.n4 a_4151_989.n3 53.105
R2847 a_4151_989.n11 a_4151_989.n10 30
R2848 a_4151_989.n9 a_4151_989.n8 24.383
R2849 a_4151_989.n11 a_4151_989.n9 23.684
R2850 a_4151_989.n13 a_4151_989.t0 14.282
R2851 a_4151_989.n13 a_4151_989.t4 14.282
R2852 a_4151_989.t2 a_4151_989.n15 14.282
R2853 a_4151_989.n15 a_4151_989.t1 14.282
R2854 a_4151_989.n15 a_4151_989.n14 12.848
R2855 a_5327_187.n5 a_5327_187.t11 512.525
R2856 a_5327_187.n3 a_5327_187.t7 472.359
R2857 a_5327_187.n1 a_5327_187.t15 472.359
R2858 a_5327_187.n3 a_5327_187.t12 384.527
R2859 a_5327_187.n1 a_5327_187.t8 384.527
R2860 a_5327_187.n5 a_5327_187.t14 371.139
R2861 a_5327_187.n6 a_5327_187.t9 340.774
R2862 a_5327_187.n4 a_5327_187.t13 294.278
R2863 a_5327_187.n2 a_5327_187.t10 294.278
R2864 a_5327_187.n13 a_5327_187.n12 266.21
R2865 a_5327_187.n14 a_5327_187.n13 117.693
R2866 a_5327_187.n6 a_5327_187.n5 109.607
R2867 a_5327_187.n7 a_5327_187.n6 83.572
R2868 a_5327_187.n8 a_5327_187.n2 81.396
R2869 a_5327_187.n16 a_5327_187.n15 79.232
R2870 a_5327_187.n7 a_5327_187.n4 76
R2871 a_5327_187.n13 a_5327_187.n8 76
R2872 a_5327_187.n16 a_5327_187.n14 63.152
R2873 a_5327_187.n4 a_5327_187.n3 56.954
R2874 a_5327_187.n2 a_5327_187.n1 56.954
R2875 a_5327_187.n12 a_5327_187.n11 30
R2876 a_5327_187.n10 a_5327_187.n9 24.383
R2877 a_5327_187.n12 a_5327_187.n10 23.684
R2878 a_5327_187.n14 a_5327_187.n0 16.08
R2879 a_5327_187.n17 a_5327_187.n16 16.078
R2880 a_5327_187.n0 a_5327_187.t2 14.282
R2881 a_5327_187.n0 a_5327_187.t3 14.282
R2882 a_5327_187.n15 a_5327_187.t5 14.282
R2883 a_5327_187.n15 a_5327_187.t6 14.282
R2884 a_5327_187.n17 a_5327_187.t0 14.282
R2885 a_5327_187.t1 a_5327_187.n17 14.282
R2886 a_5327_187.n8 a_5327_187.n7 4.035
R2887 a_7321_1050.n1 a_7321_1050.t6 512.525
R2888 a_7321_1050.n1 a_7321_1050.t7 371.139
R2889 a_7321_1050.n2 a_7321_1050.t5 287.668
R2890 a_7321_1050.n7 a_7321_1050.n6 210.592
R2891 a_7321_1050.n2 a_7321_1050.n1 162.713
R2892 a_7321_1050.n7 a_7321_1050.n2 153.315
R2893 a_7321_1050.n8 a_7321_1050.n7 152.499
R2894 a_7321_1050.n9 a_7321_1050.n8 76.001
R2895 a_7321_1050.n6 a_7321_1050.n5 30
R2896 a_7321_1050.n4 a_7321_1050.n3 24.383
R2897 a_7321_1050.n6 a_7321_1050.n4 23.684
R2898 a_7321_1050.n0 a_7321_1050.t3 14.282
R2899 a_7321_1050.n0 a_7321_1050.t2 14.282
R2900 a_7321_1050.n9 a_7321_1050.t0 14.282
R2901 a_7321_1050.t1 a_7321_1050.n9 14.282
R2902 a_7321_1050.n8 a_7321_1050.n0 12.85
R2903 D.n5 D.t5 479.223
R2904 D.n2 D.t4 479.223
R2905 D.n0 D.t7 479.223
R2906 D.n5 D.t1 375.52
R2907 D.n2 D.t6 375.52
R2908 D.n0 D.t2 375.52
R2909 D.n6 D.n5 201.982
R2910 D.n3 D.n2 201.982
R2911 D.n1 D.n0 201.982
R2912 D.n6 D.t8 141.649
R2913 D.n3 D.t3 141.649
R2914 D.n1 D.t0 141.649
R2915 D.n4 D.n1 94.999
R2916 D.n4 D.n3 76
R2917 D.n7 D.n6 76
R2918 D.n7 D.n4 18.999
R2919 D.n7 D 0.046
R2920 a_11413_103.n1 a_11413_103.n0 25.576
R2921 a_11413_103.n3 a_11413_103.n2 9.111
R2922 a_11413_103.n7 a_11413_103.n5 7.859
R2923 a_11413_103.t0 a_11413_103.n7 3.034
R2924 a_11413_103.n5 a_11413_103.n3 1.964
R2925 a_11413_103.n5 a_11413_103.n4 1.964
R2926 a_11413_103.t0 a_11413_103.n1 1.871
R2927 a_11413_103.n7 a_11413_103.n6 0.443
R2928 a_11694_210.n8 a_11694_210.n6 96.467
R2929 a_11694_210.n3 a_11694_210.n1 44.628
R2930 a_11694_210.t0 a_11694_210.n8 32.417
R2931 a_11694_210.n3 a_11694_210.n2 23.284
R2932 a_11694_210.n6 a_11694_210.n5 22.349
R2933 a_11694_210.t0 a_11694_210.n10 20.241
R2934 a_11694_210.n10 a_11694_210.n9 13.494
R2935 a_11694_210.n6 a_11694_210.n4 8.443
R2936 a_11694_210.t0 a_11694_210.n0 8.137
R2937 a_11694_210.t0 a_11694_210.n3 5.727
R2938 a_11694_210.n8 a_11694_210.n7 1.435
R2939 a_14986_101.n12 a_14986_101.n11 26.811
R2940 a_14986_101.n6 a_14986_101.n5 24.977
R2941 a_14986_101.n2 a_14986_101.n1 24.877
R2942 a_14986_101.t0 a_14986_101.n2 12.677
R2943 a_14986_101.t0 a_14986_101.n3 11.595
R2944 a_14986_101.t1 a_14986_101.n8 8.137
R2945 a_14986_101.t0 a_14986_101.n4 7.273
R2946 a_14986_101.t0 a_14986_101.n0 6.109
R2947 a_14986_101.t1 a_14986_101.n7 4.864
R2948 a_14986_101.t0 a_14986_101.n12 2.074
R2949 a_14986_101.n7 a_14986_101.n6 1.13
R2950 a_14986_101.n12 a_14986_101.t1 0.937
R2951 a_14986_101.t1 a_14986_101.n10 0.804
R2952 a_14986_101.n10 a_14986_101.n9 0.136
R2953 a_12501_1050.n1 a_12501_1050.t5 512.525
R2954 a_12501_1050.n1 a_12501_1050.t7 371.139
R2955 a_12501_1050.n2 a_12501_1050.t6 287.668
R2956 a_12501_1050.n4 a_12501_1050.n3 232.331
R2957 a_12501_1050.n2 a_12501_1050.n1 162.713
R2958 a_12501_1050.n4 a_12501_1050.n2 153.315
R2959 a_12501_1050.n5 a_12501_1050.n4 152.499
R2960 a_12501_1050.n6 a_12501_1050.n5 76.001
R2961 a_12501_1050.n0 a_12501_1050.t3 14.282
R2962 a_12501_1050.n0 a_12501_1050.t2 14.282
R2963 a_12501_1050.n6 a_12501_1050.t0 14.282
R2964 a_12501_1050.t1 a_12501_1050.n6 14.282
R2965 a_12501_1050.n5 a_12501_1050.n0 12.85
R2966 a_8823_103.n4 a_8823_103.n3 19.724
R2967 a_8823_103.t0 a_8823_103.n5 11.595
R2968 a_8823_103.t0 a_8823_103.n4 9.207
R2969 a_8823_103.n2 a_8823_103.n0 8.543
R2970 a_8823_103.t0 a_8823_103.n2 3.034
R2971 a_8823_103.n2 a_8823_103.n1 0.443
R2972 a_9104_210.n10 a_9104_210.n8 82.852
R2973 a_9104_210.n11 a_9104_210.n0 49.6
R2974 a_9104_210.n7 a_9104_210.n6 32.833
R2975 a_9104_210.n8 a_9104_210.t1 32.416
R2976 a_9104_210.n10 a_9104_210.n9 27.2
R2977 a_9104_210.n3 a_9104_210.n2 23.284
R2978 a_9104_210.n11 a_9104_210.n10 22.4
R2979 a_9104_210.n7 a_9104_210.n4 19.017
R2980 a_9104_210.n6 a_9104_210.n5 13.494
R2981 a_9104_210.t1 a_9104_210.n1 7.04
R2982 a_9104_210.t1 a_9104_210.n3 5.727
R2983 a_9104_210.n8 a_9104_210.n7 1.435
R2984 a_277_1050.n3 a_277_1050.t9 512.525
R2985 a_277_1050.n1 a_277_1050.t7 512.525
R2986 a_277_1050.n3 a_277_1050.t12 371.139
R2987 a_277_1050.n1 a_277_1050.t10 371.139
R2988 a_277_1050.n4 a_277_1050.t11 314.221
R2989 a_277_1050.n2 a_277_1050.t8 314.221
R2990 a_277_1050.n7 a_277_1050.n6 261.396
R2991 a_277_1050.n8 a_277_1050.n7 144.246
R2992 a_277_1050.n4 a_277_1050.n3 136.16
R2993 a_277_1050.n2 a_277_1050.n1 136.16
R2994 a_277_1050.n5 a_277_1050.n2 85.476
R2995 a_277_1050.n10 a_277_1050.n9 79.232
R2996 a_277_1050.n7 a_277_1050.n5 77.315
R2997 a_277_1050.n5 a_277_1050.n4 76
R2998 a_277_1050.n10 a_277_1050.n8 63.152
R2999 a_277_1050.n8 a_277_1050.n0 16.08
R3000 a_277_1050.n11 a_277_1050.n10 16.078
R3001 a_277_1050.n0 a_277_1050.t4 14.282
R3002 a_277_1050.n0 a_277_1050.t6 14.282
R3003 a_277_1050.n9 a_277_1050.t3 14.282
R3004 a_277_1050.n9 a_277_1050.t2 14.282
R3005 a_277_1050.t1 a_277_1050.n11 14.282
R3006 a_277_1050.n11 a_277_1050.t0 14.282
R3007 a_16318_101.t0 a_16318_101.n0 34.602
R3008 a_16318_101.t0 a_16318_101.n1 2.138
R3009 a_10637_1050.n3 a_10637_1050.t11 512.525
R3010 a_10637_1050.n1 a_10637_1050.t10 512.525
R3011 a_10637_1050.n3 a_10637_1050.t8 371.139
R3012 a_10637_1050.n1 a_10637_1050.t7 371.139
R3013 a_10637_1050.n4 a_10637_1050.t12 314.221
R3014 a_10637_1050.n2 a_10637_1050.t9 314.221
R3015 a_10637_1050.n10 a_10637_1050.n9 239.657
R3016 a_10637_1050.n11 a_10637_1050.n10 144.246
R3017 a_10637_1050.n4 a_10637_1050.n3 136.16
R3018 a_10637_1050.n2 a_10637_1050.n1 136.16
R3019 a_10637_1050.n5 a_10637_1050.n2 85.476
R3020 a_10637_1050.n13 a_10637_1050.n12 79.232
R3021 a_10637_1050.n10 a_10637_1050.n5 77.315
R3022 a_10637_1050.n5 a_10637_1050.n4 76
R3023 a_10637_1050.n13 a_10637_1050.n11 63.152
R3024 a_10637_1050.n9 a_10637_1050.n8 30
R3025 a_10637_1050.n7 a_10637_1050.n6 24.383
R3026 a_10637_1050.n9 a_10637_1050.n7 23.684
R3027 a_10637_1050.n11 a_10637_1050.n0 16.08
R3028 a_10637_1050.n14 a_10637_1050.n13 16.078
R3029 a_10637_1050.n0 a_10637_1050.t3 14.282
R3030 a_10637_1050.n0 a_10637_1050.t2 14.282
R3031 a_10637_1050.n12 a_10637_1050.t6 14.282
R3032 a_10637_1050.n12 a_10637_1050.t5 14.282
R3033 a_10637_1050.t1 a_10637_1050.n14 14.282
R3034 a_10637_1050.n14 a_10637_1050.t0 14.282
R3035 a_599_989.n0 a_599_989.t8 480.392
R3036 a_599_989.n2 a_599_989.t12 454.685
R3037 a_599_989.n2 a_599_989.t9 428.979
R3038 a_599_989.n0 a_599_989.t11 403.272
R3039 a_599_989.n1 a_599_989.t10 283.48
R3040 a_599_989.n3 a_599_989.t7 237.959
R3041 a_599_989.n9 a_599_989.n8 213.104
R3042 a_599_989.n13 a_599_989.n9 170.799
R3043 a_599_989.n3 a_599_989.n2 98.447
R3044 a_599_989.n1 a_599_989.n0 98.447
R3045 a_599_989.n4 a_599_989.n3 80.035
R3046 a_599_989.n12 a_599_989.n11 79.232
R3047 a_599_989.n4 a_599_989.n1 77.315
R3048 a_599_989.n9 a_599_989.n4 76
R3049 a_599_989.n13 a_599_989.n12 63.152
R3050 a_599_989.n8 a_599_989.n7 30
R3051 a_599_989.n6 a_599_989.n5 24.383
R3052 a_599_989.n8 a_599_989.n6 23.684
R3053 a_599_989.n12 a_599_989.n10 16.08
R3054 a_599_989.n14 a_599_989.n13 16.078
R3055 a_599_989.n10 a_599_989.t5 14.282
R3056 a_599_989.n10 a_599_989.t6 14.282
R3057 a_599_989.n11 a_599_989.t4 14.282
R3058 a_599_989.n11 a_599_989.t3 14.282
R3059 a_599_989.n14 a_599_989.t0 14.282
R3060 a_599_989.t1 a_599_989.n14 14.282
R3061 a_372_210.n10 a_372_210.n8 82.852
R3062 a_372_210.n7 a_372_210.n6 32.833
R3063 a_372_210.n8 a_372_210.t1 32.416
R3064 a_372_210.n10 a_372_210.n9 27.2
R3065 a_372_210.n11 a_372_210.n0 23.498
R3066 a_372_210.n3 a_372_210.n2 23.284
R3067 a_372_210.n11 a_372_210.n10 22.4
R3068 a_372_210.n7 a_372_210.n4 19.017
R3069 a_372_210.n6 a_372_210.n5 13.494
R3070 a_372_210.t1 a_372_210.n1 7.04
R3071 a_372_210.t1 a_372_210.n3 5.727
R3072 a_372_210.n8 a_372_210.n7 1.435
R3073 a_10732_210.n10 a_10732_210.n8 82.852
R3074 a_10732_210.n11 a_10732_210.n0 49.6
R3075 a_10732_210.n7 a_10732_210.n6 32.833
R3076 a_10732_210.n8 a_10732_210.t1 32.416
R3077 a_10732_210.n10 a_10732_210.n9 27.2
R3078 a_10732_210.n3 a_10732_210.n2 23.284
R3079 a_10732_210.n11 a_10732_210.n10 22.4
R3080 a_10732_210.n7 a_10732_210.n4 19.017
R3081 a_10732_210.n6 a_10732_210.n5 13.494
R3082 a_10732_210.t1 a_10732_210.n1 7.04
R3083 a_10732_210.t1 a_10732_210.n3 5.727
R3084 a_10732_210.n8 a_10732_210.n7 1.435
R3085 a_6233_103.n5 a_6233_103.n4 19.724
R3086 a_6233_103.t0 a_6233_103.n3 11.595
R3087 a_6233_103.t0 a_6233_103.n5 9.207
R3088 a_6233_103.n2 a_6233_103.n1 2.455
R3089 a_6233_103.n2 a_6233_103.n0 1.32
R3090 a_6233_103.t0 a_6233_103.n2 0.246
R3091 a_5552_210.n10 a_5552_210.n8 82.852
R3092 a_5552_210.n7 a_5552_210.n6 32.833
R3093 a_5552_210.n8 a_5552_210.t1 32.416
R3094 a_5552_210.n10 a_5552_210.n9 27.2
R3095 a_5552_210.n11 a_5552_210.n0 23.498
R3096 a_5552_210.n3 a_5552_210.n2 23.284
R3097 a_5552_210.n11 a_5552_210.n10 22.4
R3098 a_5552_210.n7 a_5552_210.n4 19.017
R3099 a_5552_210.n6 a_5552_210.n5 13.494
R3100 a_5552_210.t1 a_5552_210.n1 7.04
R3101 a_5552_210.t1 a_5552_210.n3 5.727
R3102 a_5552_210.n8 a_5552_210.n7 1.435
R3103 a_16984_101.t0 a_16984_101.n1 34.62
R3104 a_16984_101.t0 a_16984_101.n0 8.137
R3105 a_16984_101.t0 a_16984_101.n2 4.69
R3106 a_2962_210.n10 a_2962_210.n8 82.852
R3107 a_2962_210.n7 a_2962_210.n6 32.833
R3108 a_2962_210.n8 a_2962_210.t1 32.416
R3109 a_2962_210.n10 a_2962_210.n9 27.2
R3110 a_2962_210.n11 a_2962_210.n0 23.498
R3111 a_2962_210.n3 a_2962_210.n2 23.284
R3112 a_2962_210.n11 a_2962_210.n10 22.4
R3113 a_2962_210.n7 a_2962_210.n4 19.017
R3114 a_2962_210.n6 a_2962_210.n5 13.494
R3115 a_2962_210.t1 a_2962_210.n1 7.04
R3116 a_2962_210.t1 a_2962_210.n3 5.727
R3117 a_2962_210.n8 a_2962_210.n7 1.435
R3118 a_7861_103.n1 a_7861_103.n0 25.576
R3119 a_7861_103.n3 a_7861_103.n2 9.111
R3120 a_7861_103.n7 a_7861_103.n5 7.859
R3121 a_7861_103.t0 a_7861_103.n7 3.034
R3122 a_7861_103.n5 a_7861_103.n3 1.964
R3123 a_7861_103.n5 a_7861_103.n4 1.964
R3124 a_7861_103.t0 a_7861_103.n1 1.871
R3125 a_7861_103.n7 a_7861_103.n6 0.443
R3126 a_8142_210.n10 a_8142_210.n8 82.852
R3127 a_8142_210.n11 a_8142_210.n0 49.6
R3128 a_8142_210.n7 a_8142_210.n6 32.833
R3129 a_8142_210.n8 a_8142_210.t1 32.416
R3130 a_8142_210.n10 a_8142_210.n9 27.2
R3131 a_8142_210.n3 a_8142_210.n2 23.284
R3132 a_8142_210.n11 a_8142_210.n10 22.4
R3133 a_8142_210.n7 a_8142_210.n4 19.017
R3134 a_8142_210.n6 a_8142_210.n5 13.494
R3135 a_8142_210.t1 a_8142_210.n1 7.04
R3136 a_8142_210.t1 a_8142_210.n3 5.727
R3137 a_8142_210.n8 a_8142_210.n7 1.435
R3138 a_9806_101.n12 a_9806_101.n11 26.811
R3139 a_9806_101.n6 a_9806_101.n5 24.977
R3140 a_9806_101.n2 a_9806_101.n1 24.877
R3141 a_9806_101.t0 a_9806_101.n2 12.677
R3142 a_9806_101.t0 a_9806_101.n3 11.595
R3143 a_9806_101.t1 a_9806_101.n8 8.137
R3144 a_9806_101.t0 a_9806_101.n4 7.273
R3145 a_9806_101.t0 a_9806_101.n0 6.109
R3146 a_9806_101.t1 a_9806_101.n7 4.864
R3147 a_9806_101.t0 a_9806_101.n12 2.074
R3148 a_9806_101.n7 a_9806_101.n6 1.13
R3149 a_9806_101.n12 a_9806_101.t1 0.937
R3150 a_9806_101.t1 a_9806_101.n10 0.804
R3151 a_9806_101.n10 a_9806_101.n9 0.136
R3152 a_3829_1050.n1 a_3829_1050.t9 480.392
R3153 a_3829_1050.n1 a_3829_1050.t7 403.272
R3154 a_3829_1050.n2 a_3829_1050.t8 310.033
R3155 a_3829_1050.n7 a_3829_1050.n6 239.657
R3156 a_3829_1050.n7 a_3829_1050.n2 153.315
R3157 a_3829_1050.n8 a_3829_1050.n7 144.246
R3158 a_3829_1050.n10 a_3829_1050.n9 79.232
R3159 a_3829_1050.n2 a_3829_1050.n1 71.894
R3160 a_3829_1050.n10 a_3829_1050.n8 63.152
R3161 a_3829_1050.n6 a_3829_1050.n5 30
R3162 a_3829_1050.n4 a_3829_1050.n3 24.383
R3163 a_3829_1050.n6 a_3829_1050.n4 23.684
R3164 a_3829_1050.n8 a_3829_1050.n0 16.08
R3165 a_3829_1050.n11 a_3829_1050.n10 16.078
R3166 a_3829_1050.n0 a_3829_1050.t4 14.282
R3167 a_3829_1050.n0 a_3829_1050.t5 14.282
R3168 a_3829_1050.n9 a_3829_1050.t3 14.282
R3169 a_3829_1050.n9 a_3829_1050.t2 14.282
R3170 a_3829_1050.t1 a_3829_1050.n11 14.282
R3171 a_3829_1050.n11 a_3829_1050.t0 14.282
R3172 a_7216_101.n12 a_7216_101.n11 26.811
R3173 a_7216_101.n6 a_7216_101.n5 24.977
R3174 a_7216_101.n2 a_7216_101.n1 24.877
R3175 a_7216_101.t0 a_7216_101.n2 12.677
R3176 a_7216_101.t0 a_7216_101.n3 11.595
R3177 a_7216_101.t1 a_7216_101.n8 8.137
R3178 a_7216_101.t0 a_7216_101.n4 7.273
R3179 a_7216_101.t0 a_7216_101.n0 6.109
R3180 a_7216_101.t1 a_7216_101.n7 4.864
R3181 a_7216_101.t0 a_7216_101.n12 2.074
R3182 a_7216_101.n7 a_7216_101.n6 1.13
R3183 a_7216_101.n12 a_7216_101.t1 0.937
R3184 a_7216_101.t1 a_7216_101.n10 0.804
R3185 a_7216_101.n10 a_7216_101.n9 0.136
R3186 a_91_103.n1 a_91_103.n0 25.576
R3187 a_91_103.n3 a_91_103.n2 9.111
R3188 a_91_103.n7 a_91_103.n6 2.455
R3189 a_91_103.n5 a_91_103.n3 1.964
R3190 a_91_103.n5 a_91_103.n4 1.964
R3191 a_91_103.t0 a_91_103.n1 1.871
R3192 a_91_103.n7 a_91_103.n5 0.636
R3193 a_91_103.t0 a_91_103.n7 0.246
R3194 a_5271_103.n1 a_5271_103.n0 25.576
R3195 a_5271_103.n3 a_5271_103.n2 9.111
R3196 a_5271_103.n7 a_5271_103.n6 2.455
R3197 a_5271_103.n5 a_5271_103.n3 1.964
R3198 a_5271_103.n5 a_5271_103.n4 1.964
R3199 a_5271_103.t0 a_5271_103.n1 1.871
R3200 a_5271_103.n7 a_5271_103.n5 0.636
R3201 a_5271_103.t0 a_5271_103.n7 0.246
R3202 a_3924_210.n10 a_3924_210.n8 82.852
R3203 a_3924_210.n7 a_3924_210.n6 32.833
R3204 a_3924_210.n8 a_3924_210.t1 32.416
R3205 a_3924_210.n10 a_3924_210.n9 27.2
R3206 a_3924_210.n11 a_3924_210.n0 23.498
R3207 a_3924_210.n3 a_3924_210.n2 23.284
R3208 a_3924_210.n11 a_3924_210.n10 22.4
R3209 a_3924_210.n7 a_3924_210.n4 19.017
R3210 a_3924_210.n6 a_3924_210.n5 13.494
R3211 a_3924_210.t1 a_3924_210.n1 7.04
R3212 a_3924_210.t1 a_3924_210.n3 5.727
R3213 a_3924_210.n8 a_3924_210.n7 1.435
R3214 a_13322_210.n10 a_13322_210.n8 82.852
R3215 a_13322_210.n7 a_13322_210.n6 32.833
R3216 a_13322_210.n8 a_13322_210.t1 32.416
R3217 a_13322_210.n10 a_13322_210.n9 27.2
R3218 a_13322_210.n11 a_13322_210.n0 23.498
R3219 a_13322_210.n3 a_13322_210.n2 23.284
R3220 a_13322_210.n11 a_13322_210.n10 22.4
R3221 a_13322_210.n7 a_13322_210.n4 19.017
R3222 a_13322_210.n6 a_13322_210.n5 13.494
R3223 a_13322_210.t1 a_13322_210.n1 7.04
R3224 a_13322_210.t1 a_13322_210.n3 5.727
R3225 a_13322_210.n8 a_13322_210.n7 1.435
R3226 a_14284_210.n10 a_14284_210.n8 82.852
R3227 a_14284_210.n7 a_14284_210.n6 32.833
R3228 a_14284_210.n8 a_14284_210.t1 32.416
R3229 a_14284_210.n10 a_14284_210.n9 27.2
R3230 a_14284_210.n11 a_14284_210.n0 23.498
R3231 a_14284_210.n3 a_14284_210.n2 23.284
R3232 a_14284_210.n11 a_14284_210.n10 22.4
R3233 a_14284_210.n7 a_14284_210.n4 19.017
R3234 a_14284_210.n6 a_14284_210.n5 13.494
R3235 a_14284_210.t1 a_14284_210.n1 7.04
R3236 a_14284_210.t1 a_14284_210.n3 5.727
R3237 a_14284_210.n8 a_14284_210.n7 1.435
R3238 a_13041_103.n1 a_13041_103.n0 25.576
R3239 a_13041_103.n3 a_13041_103.n2 9.111
R3240 a_13041_103.n7 a_13041_103.n6 2.455
R3241 a_13041_103.n5 a_13041_103.n3 1.964
R3242 a_13041_103.n5 a_13041_103.n4 1.964
R3243 a_13041_103.t0 a_13041_103.n1 1.871
R3244 a_13041_103.n7 a_13041_103.n5 0.636
R3245 a_13041_103.t0 a_13041_103.n7 0.246
R3246 a_3643_103.n1 a_3643_103.n0 25.576
R3247 a_3643_103.n3 a_3643_103.n2 9.111
R3248 a_3643_103.n7 a_3643_103.n6 2.455
R3249 a_3643_103.n5 a_3643_103.n3 1.964
R3250 a_3643_103.n5 a_3643_103.n4 1.964
R3251 a_3643_103.t0 a_3643_103.n1 1.871
R3252 a_3643_103.n7 a_3643_103.n5 0.636
R3253 a_3643_103.t0 a_3643_103.n7 0.246
R3254 a_4626_101.t0 a_4626_101.n1 34.62
R3255 a_4626_101.t0 a_4626_101.n0 8.137
R3256 a_4626_101.t0 a_4626_101.n2 4.69
R3257 a_14003_103.n1 a_14003_103.n0 25.576
R3258 a_14003_103.n3 a_14003_103.n2 9.111
R3259 a_14003_103.n7 a_14003_103.n6 2.455
R3260 a_14003_103.n5 a_14003_103.n3 1.964
R3261 a_14003_103.n5 a_14003_103.n4 1.964
R3262 a_14003_103.t0 a_14003_103.n1 1.871
R3263 a_14003_103.n7 a_14003_103.n5 0.636
R3264 a_14003_103.t0 a_14003_103.n7 0.246
R3265 a_2681_103.n1 a_2681_103.n0 25.576
R3266 a_2681_103.n3 a_2681_103.n2 9.111
R3267 a_2681_103.n7 a_2681_103.n6 2.455
R3268 a_2681_103.n5 a_2681_103.n3 1.964
R3269 a_2681_103.n5 a_2681_103.n4 1.964
R3270 a_2681_103.t0 a_2681_103.n1 1.871
R3271 a_2681_103.n7 a_2681_103.n5 0.636
R3272 a_2681_103.t0 a_2681_103.n7 0.246
R3273 a_1334_210.n9 a_1334_210.n7 82.852
R3274 a_1334_210.n3 a_1334_210.n1 44.628
R3275 a_1334_210.t0 a_1334_210.n9 32.417
R3276 a_1334_210.n7 a_1334_210.n6 27.2
R3277 a_1334_210.n5 a_1334_210.n4 23.498
R3278 a_1334_210.n3 a_1334_210.n2 23.284
R3279 a_1334_210.n7 a_1334_210.n5 22.4
R3280 a_1334_210.t0 a_1334_210.n11 20.241
R3281 a_1334_210.n11 a_1334_210.n10 13.494
R3282 a_1334_210.t0 a_1334_210.n0 8.137
R3283 a_1334_210.t0 a_1334_210.n3 5.727
R3284 a_1334_210.n9 a_1334_210.n8 1.435
R3285 a_1053_103.n5 a_1053_103.n4 19.724
R3286 a_1053_103.t0 a_1053_103.n3 11.595
R3287 a_1053_103.t0 a_1053_103.n5 9.207
R3288 a_1053_103.n2 a_1053_103.n1 2.455
R3289 a_1053_103.n2 a_1053_103.n0 1.32
R3290 a_1053_103.t0 a_1053_103.n2 0.246
C7 RN GND 10.14fF
C8 VDD GND 63.35fF
C9 a_1053_103.n0 GND 0.10fF
C10 a_1053_103.n1 GND 0.04fF
C11 a_1053_103.n2 GND 0.03fF
C12 a_1053_103.n3 GND 0.07fF
C13 a_1053_103.n4 GND 0.08fF
C14 a_1053_103.n5 GND 0.06fF
C15 a_1334_210.n0 GND 0.07fF
C16 a_1334_210.n1 GND 0.09fF
C17 a_1334_210.n2 GND 0.13fF
C18 a_1334_210.n3 GND 0.11fF
C19 a_1334_210.n4 GND 0.02fF
C20 a_1334_210.n5 GND 0.03fF
C21 a_1334_210.n6 GND 0.02fF
C22 a_1334_210.n7 GND 0.05fF
C23 a_1334_210.n8 GND 0.03fF
C24 a_1334_210.n9 GND 0.11fF
C25 a_1334_210.n10 GND 0.06fF
C26 a_1334_210.n11 GND 0.01fF
C27 a_1334_210.t0 GND 0.33fF
C28 a_2681_103.n0 GND 0.09fF
C29 a_2681_103.n1 GND 0.10fF
C30 a_2681_103.n2 GND 0.05fF
C31 a_2681_103.n3 GND 0.03fF
C32 a_2681_103.n4 GND 0.04fF
C33 a_2681_103.n5 GND 0.03fF
C34 a_2681_103.n6 GND 0.04fF
C35 a_14003_103.n0 GND 0.09fF
C36 a_14003_103.n1 GND 0.10fF
C37 a_14003_103.n2 GND 0.05fF
C38 a_14003_103.n3 GND 0.03fF
C39 a_14003_103.n4 GND 0.04fF
C40 a_14003_103.n5 GND 0.03fF
C41 a_14003_103.n6 GND 0.04fF
C42 a_4626_101.n0 GND 0.05fF
C43 a_4626_101.n1 GND 0.12fF
C44 a_4626_101.n2 GND 0.04fF
C45 a_3643_103.n0 GND 0.09fF
C46 a_3643_103.n1 GND 0.10fF
C47 a_3643_103.n2 GND 0.05fF
C48 a_3643_103.n3 GND 0.03fF
C49 a_3643_103.n4 GND 0.04fF
C50 a_3643_103.n5 GND 0.03fF
C51 a_3643_103.n6 GND 0.04fF
C52 a_13041_103.n0 GND 0.09fF
C53 a_13041_103.n1 GND 0.10fF
C54 a_13041_103.n2 GND 0.05fF
C55 a_13041_103.n3 GND 0.03fF
C56 a_13041_103.n4 GND 0.04fF
C57 a_13041_103.n5 GND 0.03fF
C58 a_13041_103.n6 GND 0.04fF
C59 a_14284_210.n0 GND 0.02fF
C60 a_14284_210.n1 GND 0.09fF
C61 a_14284_210.n2 GND 0.13fF
C62 a_14284_210.n3 GND 0.11fF
C63 a_14284_210.t1 GND 0.30fF
C64 a_14284_210.n4 GND 0.09fF
C65 a_14284_210.n5 GND 0.06fF
C66 a_14284_210.n6 GND 0.01fF
C67 a_14284_210.n7 GND 0.03fF
C68 a_14284_210.n8 GND 0.11fF
C69 a_14284_210.n9 GND 0.02fF
C70 a_14284_210.n10 GND 0.05fF
C71 a_14284_210.n11 GND 0.03fF
C72 a_13322_210.n0 GND 0.02fF
C73 a_13322_210.n1 GND 0.09fF
C74 a_13322_210.n2 GND 0.13fF
C75 a_13322_210.n3 GND 0.11fF
C76 a_13322_210.t1 GND 0.30fF
C77 a_13322_210.n4 GND 0.09fF
C78 a_13322_210.n5 GND 0.06fF
C79 a_13322_210.n6 GND 0.01fF
C80 a_13322_210.n7 GND 0.03fF
C81 a_13322_210.n8 GND 0.11fF
C82 a_13322_210.n9 GND 0.02fF
C83 a_13322_210.n10 GND 0.05fF
C84 a_13322_210.n11 GND 0.03fF
C85 a_3924_210.n0 GND 0.02fF
C86 a_3924_210.n1 GND 0.09fF
C87 a_3924_210.n2 GND 0.13fF
C88 a_3924_210.n3 GND 0.11fF
C89 a_3924_210.t1 GND 0.30fF
C90 a_3924_210.n4 GND 0.09fF
C91 a_3924_210.n5 GND 0.06fF
C92 a_3924_210.n6 GND 0.01fF
C93 a_3924_210.n7 GND 0.03fF
C94 a_3924_210.n8 GND 0.11fF
C95 a_3924_210.n9 GND 0.02fF
C96 a_3924_210.n10 GND 0.05fF
C97 a_3924_210.n11 GND 0.03fF
C98 a_5271_103.n0 GND 0.09fF
C99 a_5271_103.n1 GND 0.10fF
C100 a_5271_103.n2 GND 0.05fF
C101 a_5271_103.n3 GND 0.03fF
C102 a_5271_103.n4 GND 0.04fF
C103 a_5271_103.n5 GND 0.03fF
C104 a_5271_103.n6 GND 0.04fF
C105 a_91_103.n0 GND 0.09fF
C106 a_91_103.n1 GND 0.09fF
C107 a_91_103.n2 GND 0.04fF
C108 a_91_103.n3 GND 0.03fF
C109 a_91_103.n4 GND 0.04fF
C110 a_91_103.n5 GND 0.03fF
C111 a_91_103.n6 GND 0.04fF
C112 a_7216_101.n0 GND 0.02fF
C113 a_7216_101.n1 GND 0.10fF
C114 a_7216_101.n2 GND 0.06fF
C115 a_7216_101.n3 GND 0.06fF
C116 a_7216_101.n4 GND 0.00fF
C117 a_7216_101.n5 GND 0.04fF
C118 a_7216_101.n6 GND 0.05fF
C119 a_7216_101.n7 GND 0.02fF
C120 a_7216_101.n8 GND 0.05fF
C121 a_7216_101.n9 GND 0.08fF
C122 a_7216_101.n10 GND 0.17fF
C123 a_7216_101.t1 GND 0.23fF
C124 a_7216_101.n11 GND 0.09fF
C125 a_7216_101.n12 GND 0.00fF
C126 a_3829_1050.n0 GND 0.50fF
C127 a_3829_1050.n1 GND 0.32fF
C128 a_3829_1050.n2 GND 0.54fF
C129 a_3829_1050.n3 GND 0.04fF
C130 a_3829_1050.n4 GND 0.05fF
C131 a_3829_1050.n5 GND 0.03fF
C132 a_3829_1050.n6 GND 0.31fF
C133 a_3829_1050.n7 GND 0.59fF
C134 a_3829_1050.n8 GND 0.26fF
C135 a_3829_1050.n9 GND 0.59fF
C136 a_3829_1050.n10 GND 0.19fF
C137 a_3829_1050.n11 GND 0.50fF
C138 a_9806_101.n0 GND 0.02fF
C139 a_9806_101.n1 GND 0.10fF
C140 a_9806_101.n2 GND 0.06fF
C141 a_9806_101.n3 GND 0.06fF
C142 a_9806_101.n4 GND 0.00fF
C143 a_9806_101.n5 GND 0.04fF
C144 a_9806_101.n6 GND 0.05fF
C145 a_9806_101.n7 GND 0.02fF
C146 a_9806_101.n8 GND 0.05fF
C147 a_9806_101.n9 GND 0.08fF
C148 a_9806_101.n10 GND 0.17fF
C149 a_9806_101.t1 GND 0.23fF
C150 a_9806_101.n11 GND 0.09fF
C151 a_9806_101.n12 GND 0.00fF
C152 a_8142_210.n0 GND 0.02fF
C153 a_8142_210.n1 GND 0.09fF
C154 a_8142_210.n2 GND 0.13fF
C155 a_8142_210.n3 GND 0.11fF
C156 a_8142_210.t1 GND 0.30fF
C157 a_8142_210.n4 GND 0.09fF
C158 a_8142_210.n5 GND 0.06fF
C159 a_8142_210.n6 GND 0.01fF
C160 a_8142_210.n7 GND 0.03fF
C161 a_8142_210.n8 GND 0.11fF
C162 a_8142_210.n9 GND 0.02fF
C163 a_8142_210.n10 GND 0.05fF
C164 a_8142_210.n11 GND 0.02fF
C165 a_7861_103.n0 GND 0.09fF
C166 a_7861_103.n1 GND 0.10fF
C167 a_7861_103.n2 GND 0.05fF
C168 a_7861_103.n3 GND 0.03fF
C169 a_7861_103.n4 GND 0.04fF
C170 a_7861_103.n5 GND 0.11fF
C171 a_7861_103.n6 GND 0.04fF
C172 a_2962_210.n0 GND 0.02fF
C173 a_2962_210.n1 GND 0.09fF
C174 a_2962_210.n2 GND 0.13fF
C175 a_2962_210.n3 GND 0.11fF
C176 a_2962_210.t1 GND 0.30fF
C177 a_2962_210.n4 GND 0.09fF
C178 a_2962_210.n5 GND 0.06fF
C179 a_2962_210.n6 GND 0.01fF
C180 a_2962_210.n7 GND 0.03fF
C181 a_2962_210.n8 GND 0.11fF
C182 a_2962_210.n9 GND 0.02fF
C183 a_2962_210.n10 GND 0.05fF
C184 a_2962_210.n11 GND 0.03fF
C185 a_16984_101.n0 GND 0.06fF
C186 a_16984_101.n1 GND 0.13fF
C187 a_16984_101.n2 GND 0.04fF
C188 a_5552_210.n0 GND 0.02fF
C189 a_5552_210.n1 GND 0.09fF
C190 a_5552_210.n2 GND 0.13fF
C191 a_5552_210.n3 GND 0.11fF
C192 a_5552_210.t1 GND 0.30fF
C193 a_5552_210.n4 GND 0.09fF
C194 a_5552_210.n5 GND 0.06fF
C195 a_5552_210.n6 GND 0.01fF
C196 a_5552_210.n7 GND 0.03fF
C197 a_5552_210.n8 GND 0.11fF
C198 a_5552_210.n9 GND 0.02fF
C199 a_5552_210.n10 GND 0.05fF
C200 a_5552_210.n11 GND 0.03fF
C201 a_6233_103.n0 GND 0.10fF
C202 a_6233_103.n1 GND 0.04fF
C203 a_6233_103.n2 GND 0.03fF
C204 a_6233_103.n3 GND 0.07fF
C205 a_6233_103.n4 GND 0.08fF
C206 a_6233_103.n5 GND 0.06fF
C207 a_10732_210.n0 GND 0.02fF
C208 a_10732_210.n1 GND 0.09fF
C209 a_10732_210.n2 GND 0.13fF
C210 a_10732_210.n3 GND 0.11fF
C211 a_10732_210.t1 GND 0.30fF
C212 a_10732_210.n4 GND 0.09fF
C213 a_10732_210.n5 GND 0.06fF
C214 a_10732_210.n6 GND 0.01fF
C215 a_10732_210.n7 GND 0.03fF
C216 a_10732_210.n8 GND 0.11fF
C217 a_10732_210.n9 GND 0.02fF
C218 a_10732_210.n10 GND 0.05fF
C219 a_10732_210.n11 GND 0.02fF
C220 a_372_210.n0 GND 0.02fF
C221 a_372_210.n1 GND 0.09fF
C222 a_372_210.n2 GND 0.13fF
C223 a_372_210.n3 GND 0.11fF
C224 a_372_210.t1 GND 0.30fF
C225 a_372_210.n4 GND 0.09fF
C226 a_372_210.n5 GND 0.06fF
C227 a_372_210.n6 GND 0.01fF
C228 a_372_210.n7 GND 0.03fF
C229 a_372_210.n8 GND 0.11fF
C230 a_372_210.n9 GND 0.02fF
C231 a_372_210.n10 GND 0.05fF
C232 a_372_210.n11 GND 0.03fF
C233 a_599_989.n0 GND 0.40fF
C234 a_599_989.n1 GND 0.43fF
C235 a_599_989.n2 GND 0.40fF
C236 a_599_989.t7 GND 0.57fF
C237 a_599_989.n3 GND 0.42fF
C238 a_599_989.n4 GND 1.34fF
C239 a_599_989.n5 GND 0.04fF
C240 a_599_989.n6 GND 0.06fF
C241 a_599_989.n7 GND 0.04fF
C242 a_599_989.n8 GND 0.32fF
C243 a_599_989.n9 GND 0.48fF
C244 a_599_989.n10 GND 0.58fF
C245 a_599_989.n11 GND 0.68fF
C246 a_599_989.n12 GND 0.21fF
C247 a_599_989.n13 GND 0.33fF
C248 a_599_989.n14 GND 0.58fF
C249 a_10637_1050.n0 GND 0.87fF
C250 a_10637_1050.n1 GND 0.50fF
C251 a_10637_1050.n2 GND 0.98fF
C252 a_10637_1050.n3 GND 0.50fF
C253 a_10637_1050.n4 GND 0.78fF
C254 a_10637_1050.n5 GND 3.83fF
C255 a_10637_1050.n6 GND 0.07fF
C256 a_10637_1050.n7 GND 0.09fF
C257 a_10637_1050.n8 GND 0.06fF
C258 a_10637_1050.n9 GND 0.54fF
C259 a_10637_1050.n10 GND 0.74fF
C260 a_10637_1050.n11 GND 0.45fF
C261 a_10637_1050.n12 GND 1.02fF
C262 a_10637_1050.n13 GND 0.32fF
C263 a_10637_1050.n14 GND 0.87fF
C264 a_16318_101.n0 GND 0.13fF
C265 a_16318_101.n1 GND 0.13fF
C266 a_277_1050.n0 GND 0.78fF
C267 a_277_1050.n1 GND 0.44fF
C268 a_277_1050.n2 GND 0.87fF
C269 a_277_1050.n3 GND 0.44fF
C270 a_277_1050.n4 GND 0.70fF
C271 a_277_1050.n5 GND 3.41fF
C272 a_277_1050.n6 GND 0.62fF
C273 a_277_1050.n7 GND 0.70fF
C274 a_277_1050.n8 GND 0.40fF
C275 a_277_1050.n9 GND 0.91fF
C276 a_277_1050.n10 GND 0.29fF
C277 a_277_1050.n11 GND 0.78fF
C278 a_9104_210.n0 GND 0.02fF
C279 a_9104_210.n1 GND 0.09fF
C280 a_9104_210.n2 GND 0.13fF
C281 a_9104_210.n3 GND 0.11fF
C282 a_9104_210.t1 GND 0.30fF
C283 a_9104_210.n4 GND 0.09fF
C284 a_9104_210.n5 GND 0.06fF
C285 a_9104_210.n6 GND 0.01fF
C286 a_9104_210.n7 GND 0.03fF
C287 a_9104_210.n8 GND 0.11fF
C288 a_9104_210.n9 GND 0.02fF
C289 a_9104_210.n10 GND 0.05fF
C290 a_9104_210.n11 GND 0.02fF
C291 a_8823_103.n0 GND 0.20fF
C292 a_8823_103.n1 GND 0.04fF
C293 a_8823_103.n2 GND 0.01fF
C294 a_8823_103.n3 GND 0.08fF
C295 a_8823_103.n4 GND 0.06fF
C296 a_8823_103.n5 GND 0.07fF
C297 a_12501_1050.n0 GND 0.60fF
C298 a_12501_1050.n1 GND 0.38fF
C299 a_12501_1050.n2 GND 0.75fF
C300 a_12501_1050.n3 GND 0.45fF
C301 a_12501_1050.n4 GND 0.72fF
C302 a_12501_1050.n5 GND 0.35fF
C303 a_12501_1050.n6 GND 0.71fF
C304 a_14986_101.n0 GND 0.02fF
C305 a_14986_101.n1 GND 0.10fF
C306 a_14986_101.n2 GND 0.06fF
C307 a_14986_101.n3 GND 0.06fF
C308 a_14986_101.n4 GND 0.00fF
C309 a_14986_101.n5 GND 0.04fF
C310 a_14986_101.n6 GND 0.05fF
C311 a_14986_101.n7 GND 0.02fF
C312 a_14986_101.n8 GND 0.05fF
C313 a_14986_101.n9 GND 0.08fF
C314 a_14986_101.n10 GND 0.17fF
C315 a_14986_101.t1 GND 0.23fF
C316 a_14986_101.n11 GND 0.09fF
C317 a_14986_101.n12 GND 0.00fF
C318 a_11694_210.n0 GND 0.07fF
C319 a_11694_210.n1 GND 0.09fF
C320 a_11694_210.n2 GND 0.13fF
C321 a_11694_210.n3 GND 0.11fF
C322 a_11694_210.n4 GND 0.02fF
C323 a_11694_210.n5 GND 0.03fF
C324 a_11694_210.n6 GND 0.06fF
C325 a_11694_210.n7 GND 0.03fF
C326 a_11694_210.n8 GND 0.12fF
C327 a_11694_210.n9 GND 0.06fF
C328 a_11694_210.n10 GND 0.01fF
C329 a_11694_210.t0 GND 0.33fF
C330 a_11413_103.n0 GND 0.09fF
C331 a_11413_103.n1 GND 0.10fF
C332 a_11413_103.n2 GND 0.05fF
C333 a_11413_103.n3 GND 0.03fF
C334 a_11413_103.n4 GND 0.04fF
C335 a_11413_103.n5 GND 0.11fF
C336 a_11413_103.n6 GND 0.04fF
C337 a_7321_1050.n0 GND 0.56fF
C338 a_7321_1050.n1 GND 0.36fF
C339 a_7321_1050.n2 GND 0.70fF
C340 a_7321_1050.n3 GND 0.04fF
C341 a_7321_1050.n4 GND 0.06fF
C342 a_7321_1050.n5 GND 0.04fF
C343 a_7321_1050.n6 GND 0.32fF
C344 a_7321_1050.n7 GND 0.64fF
C345 a_7321_1050.n8 GND 0.33fF
C346 a_7321_1050.n9 GND 0.67fF
C347 a_5327_187.n0 GND 0.89fF
C348 a_5327_187.n1 GND 0.46fF
C349 a_5327_187.t10 GND 0.98fF
C350 a_5327_187.n2 GND 0.70fF
C351 a_5327_187.n3 GND 0.46fF
C352 a_5327_187.t13 GND 0.98fF
C353 a_5327_187.n4 GND 0.63fF
C354 a_5327_187.n5 GND 0.45fF
C355 a_5327_187.n6 GND 0.94fF
C356 a_5327_187.n7 GND 3.49fF
C357 a_5327_187.n8 GND 2.75fF
C358 a_5327_187.n9 GND 0.07fF
C359 a_5327_187.n10 GND 0.09fF
C360 a_5327_187.n11 GND 0.06fF
C361 a_5327_187.n12 GND 0.60fF
C362 a_5327_187.n13 GND 0.75fF
C363 a_5327_187.n14 GND 0.41fF
C364 a_5327_187.n15 GND 1.05fF
C365 a_5327_187.n16 GND 0.33fF
C366 a_5327_187.n17 GND 0.89fF
C367 a_4151_989.n0 GND 0.92fF
C368 a_4151_989.n1 GND 1.06fF
C369 a_4151_989.n2 GND 1.30fF
C370 a_4151_989.n3 GND 0.74fF
C371 a_4151_989.n4 GND 4.56fF
C372 a_4151_989.n5 GND 0.98fF
C373 a_4151_989.t8 GND 1.07fF
C374 a_4151_989.n6 GND 0.83fF
C375 a_4151_989.n7 GND 19.06fF
C376 a_4151_989.n8 GND 0.09fF
C377 a_4151_989.n9 GND 0.12fF
C378 a_4151_989.n10 GND 0.08fF
C379 a_4151_989.n11 GND 0.53fF
C380 a_4151_989.n12 GND 0.96fF
C381 a_4151_989.n13 GND 1.40fF
C382 a_4151_989.n14 GND 0.82fF
C383 a_4151_989.n15 GND 1.19fF
C384 a_6514_210.n0 GND 0.02fF
C385 a_6514_210.n1 GND 0.09fF
C386 a_6514_210.n2 GND 0.13fF
C387 a_6514_210.n3 GND 0.11fF
C388 a_6514_210.t1 GND 0.30fF
C389 a_6514_210.n4 GND 0.09fF
C390 a_6514_210.n5 GND 0.06fF
C391 a_6514_210.n6 GND 0.01fF
C392 a_6514_210.n7 GND 0.03fF
C393 a_6514_210.n8 GND 0.11fF
C394 a_6514_210.n9 GND 0.02fF
C395 a_6514_210.n10 GND 0.05fF
C396 a_6514_210.n11 GND 0.02fF
C397 QN.n0 GND 0.42fF
C398 QN.n1 GND 0.51fF
C399 QN.n2 GND 0.25fF
C400 QN.n3 GND 0.04fF
C401 QN.n4 GND 0.05fF
C402 QN.n5 GND 0.11fF
C403 QN.n6 GND 0.20fF
C404 QN.n7 GND 1.11fF
C405 QN.n8 GND 0.06fF
C406 QN.n9 GND 0.03fF
C407 QN.n10 GND 0.08fF
C408 QN.n11 GND 0.28fF
C409 QN.n12 GND 0.37fF
C410 QN.n13 GND 0.01fF
C411 a_15652_101.n0 GND 0.11fF
C412 a_15652_101.n1 GND 0.09fF
C413 a_15652_101.n2 GND 0.08fF
C414 a_15652_101.n3 GND 0.02fF
C415 a_15652_101.n4 GND 0.01fF
C416 a_15652_101.n5 GND 0.06fF
C417 a_14189_1050.n0 GND 0.53fF
C418 a_14189_1050.n1 GND 0.34fF
C419 a_14189_1050.n2 GND 0.56fF
C420 a_14189_1050.n3 GND 0.04fF
C421 a_14189_1050.n4 GND 0.05fF
C422 a_14189_1050.n5 GND 0.03fF
C423 a_14189_1050.n6 GND 0.33fF
C424 a_14189_1050.n7 GND 0.61fF
C425 a_14189_1050.n8 GND 0.27fF
C426 a_14189_1050.n9 GND 0.62fF
C427 a_14189_1050.n10 GND 0.19fF
C428 a_14189_1050.n11 GND 0.53fF
C429 a_14511_989.n0 GND 0.30fF
C430 a_14511_989.n1 GND 0.34fF
C431 a_14511_989.n2 GND 1.06fF
C432 a_14511_989.n3 GND 0.76fF
C433 a_14511_989.n4 GND 0.35fF
C434 a_14511_989.n5 GND 0.41fF
C435 a_14511_989.t10 GND 0.58fF
C436 a_14511_989.n6 GND 0.42fF
C437 a_14511_989.n7 GND 1.24fF
C438 a_14511_989.n8 GND 0.04fF
C439 a_14511_989.n9 GND 0.06fF
C440 a_14511_989.n10 GND 0.04fF
C441 a_14511_989.n11 GND 0.33fF
C442 a_14511_989.n12 GND 0.46fF
C443 a_14511_989.n13 GND 0.69fF
C444 a_14511_989.n14 GND 0.33fF
C445 a_14511_989.n15 GND 0.58fF
C446 a_15757_1051.n0 GND 0.37fF
C447 a_15757_1051.n1 GND 0.33fF
C448 a_15757_1051.n2 GND 0.23fF
C449 a_15757_1051.n3 GND 0.62fF
C450 a_15757_1051.n4 GND 0.28fF
C451 a_15757_1051.n5 GND 0.41fF
C452 a_16421_1051.n0 GND 0.28fF
C453 a_16421_1051.n1 GND 0.27fF
C454 a_16421_1051.n2 GND 0.35fF
C455 a_16421_1051.n3 GND 0.24fF
C456 a_16421_1051.n4 GND 0.55fF
C457 a_16421_1051.n5 GND 0.20fF
C458 a_10451_103.n0 GND 0.09fF
C459 a_10451_103.n1 GND 0.10fF
C460 a_10451_103.n2 GND 0.05fF
C461 a_10451_103.n3 GND 0.03fF
C462 a_10451_103.n4 GND 0.04fF
C463 a_10451_103.n5 GND 0.11fF
C464 a_10451_103.n6 GND 0.04fF
C465 a_10507_187.n0 GND 0.84fF
C466 a_10507_187.n1 GND 0.44fF
C467 a_10507_187.t8 GND 0.93fF
C468 a_10507_187.n2 GND 0.67fF
C469 a_10507_187.n3 GND 0.44fF
C470 a_10507_187.t11 GND 0.93fF
C471 a_10507_187.n4 GND 0.60fF
C472 a_10507_187.n5 GND 0.43fF
C473 a_10507_187.n6 GND 0.89fF
C474 a_10507_187.n7 GND 3.31fF
C475 a_10507_187.n8 GND 2.61fF
C476 a_10507_187.n9 GND 0.06fF
C477 a_10507_187.n10 GND 0.08fF
C478 a_10507_187.n11 GND 0.05fF
C479 a_10507_187.n12 GND 0.57fF
C480 a_10507_187.n13 GND 0.71fF
C481 a_10507_187.n14 GND 0.38fF
C482 a_10507_187.n15 GND 0.99fF
C483 a_10507_187.n16 GND 0.31fF
C484 a_10507_187.n17 GND 0.84fF
C485 a_5457_1050.n0 GND 0.84fF
C486 a_5457_1050.n1 GND 0.48fF
C487 a_5457_1050.n2 GND 0.94fF
C488 a_5457_1050.n3 GND 0.48fF
C489 a_5457_1050.n4 GND 0.76fF
C490 a_5457_1050.n5 GND 3.70fF
C491 a_5457_1050.n6 GND 0.06fF
C492 a_5457_1050.n7 GND 0.08fF
C493 a_5457_1050.n8 GND 0.05fF
C494 a_5457_1050.n9 GND 0.52fF
C495 a_5457_1050.n10 GND 0.71fF
C496 a_5457_1050.n11 GND 0.43fF
C497 a_5457_1050.n12 GND 0.99fF
C498 a_5457_1050.n13 GND 0.31fF
C499 a_5457_1050.n14 GND 0.84fF
C500 a_2141_1050.n0 GND 0.34fF
C501 a_2141_1050.n1 GND 0.67fF
C502 a_2141_1050.n2 GND 0.40fF
C503 a_2141_1050.n3 GND 0.64fF
C504 a_2141_1050.n4 GND 0.64fF
C505 a_2141_1050.n5 GND 0.31fF
C506 a_2141_1050.n6 GND 0.54fF
C507 a_2036_101.n0 GND 0.05fF
C508 a_2036_101.n1 GND 0.12fF
C509 a_2036_101.n2 GND 0.04fF
C510 a_147_187.n0 GND 0.42fF
C511 a_147_187.t15 GND 0.90fF
C512 a_147_187.n1 GND 0.65fF
C513 a_147_187.n2 GND 0.42fF
C514 a_147_187.t7 GND 0.90fF
C515 a_147_187.n3 GND 0.58fF
C516 a_147_187.n4 GND 0.42fF
C517 a_147_187.n5 GND 0.87fF
C518 a_147_187.n6 GND 3.22fF
C519 a_147_187.n7 GND 2.54fF
C520 a_147_187.n8 GND 0.06fF
C521 a_147_187.n9 GND 0.08fF
C522 a_147_187.n10 GND 0.05fF
C523 a_147_187.n11 GND 0.56fF
C524 a_147_187.n12 GND 0.69fF
C525 a_147_187.n13 GND 0.82fF
C526 a_147_187.n14 GND 0.96fF
C527 a_147_187.n15 GND 0.30fF
C528 a_147_187.n16 GND 0.37fF
C529 a_147_187.n17 GND 0.82fF
C530 a_9009_1050.n0 GND 0.53fF
C531 a_9009_1050.n1 GND 0.34fF
C532 a_9009_1050.n2 GND 0.56fF
C533 a_9009_1050.n3 GND 0.04fF
C534 a_9009_1050.n4 GND 0.05fF
C535 a_9009_1050.n5 GND 0.03fF
C536 a_9009_1050.n6 GND 0.33fF
C537 a_9009_1050.n7 GND 0.61fF
C538 a_9009_1050.n8 GND 0.27fF
C539 a_9009_1050.n9 GND 0.62fF
C540 a_9009_1050.n10 GND 0.19fF
C541 a_9009_1050.n11 GND 0.53fF
C542 a_9331_989.n0 GND 1.05fF
C543 a_9331_989.n1 GND 1.25fF
C544 a_9331_989.n2 GND 0.67fF
C545 a_9331_989.n3 GND 0.55fF
C546 a_9331_989.n4 GND 1.47fF
C547 a_9331_989.n5 GND 0.49fF
C548 a_9331_989.n6 GND 1.11fF
C549 a_9331_989.n7 GND 1.66fF
C550 a_9331_989.n8 GND 0.81fF
C551 a_9331_989.t12 GND 1.00fF
C552 a_9331_989.n9 GND 0.75fF
C553 a_9331_989.n10 GND 9.37fF
C554 a_9331_989.n11 GND 0.87fF
C555 a_9331_989.n12 GND 0.17fF
C556 a_9331_989.n13 GND 0.51fF
C557 a_9331_989.n14 GND 0.09fF
C558 a_5779_989.n0 GND 0.46fF
C559 a_5779_989.n1 GND 0.48fF
C560 a_5779_989.n2 GND 0.46fF
C561 a_5779_989.t8 GND 0.65fF
C562 a_5779_989.n3 GND 0.48fF
C563 a_5779_989.n4 GND 1.51fF
C564 a_5779_989.n5 GND 0.05fF
C565 a_5779_989.n6 GND 0.07fF
C566 a_5779_989.n7 GND 0.04fF
C567 a_5779_989.n8 GND 0.37fF
C568 a_5779_989.n9 GND 0.55fF
C569 a_5779_989.n10 GND 0.65fF
C570 a_5779_989.n11 GND 0.76fF
C571 a_5779_989.n12 GND 0.24fF
C572 a_5779_989.n13 GND 0.37fF
C573 a_5779_989.n14 GND 0.65fF
C574 VDD.n0 GND 0.16fF
C575 VDD.n1 GND 0.03fF
C576 VDD.n2 GND 0.02fF
C577 VDD.n3 GND 0.05fF
C578 VDD.n4 GND 0.01fF
C579 VDD.n5 GND 0.02fF
C580 VDD.n6 GND 0.02fF
C581 VDD.n8 GND 0.02fF
C582 VDD.n9 GND 0.02fF
C583 VDD.n11 GND 0.02fF
C584 VDD.n14 GND 0.46fF
C585 VDD.n16 GND 0.03fF
C586 VDD.n17 GND 0.02fF
C587 VDD.n18 GND 0.02fF
C588 VDD.n19 GND 0.02fF
C589 VDD.n20 GND 0.04fF
C590 VDD.n21 GND 0.28fF
C591 VDD.n22 GND 0.02fF
C592 VDD.n23 GND 0.03fF
C593 VDD.n24 GND 0.28fF
C594 VDD.n25 GND 0.01fF
C595 VDD.n26 GND 0.31fF
C596 VDD.n27 GND 0.01fF
C597 VDD.n28 GND 0.03fF
C598 VDD.n29 GND 0.02fF
C599 VDD.n30 GND 0.28fF
C600 VDD.n31 GND 0.01fF
C601 VDD.n32 GND 0.02fF
C602 VDD.n33 GND 0.00fF
C603 VDD.n34 GND 0.09fF
C604 VDD.n35 GND 0.03fF
C605 VDD.n36 GND 0.31fF
C606 VDD.n37 GND 0.01fF
C607 VDD.n38 GND 0.03fF
C608 VDD.n39 GND 0.03fF
C609 VDD.n40 GND 0.28fF
C610 VDD.n41 GND 0.01fF
C611 VDD.n42 GND 0.02fF
C612 VDD.n43 GND 0.02fF
C613 VDD.n44 GND 0.28fF
C614 VDD.n45 GND 0.01fF
C615 VDD.n46 GND 0.02fF
C616 VDD.n47 GND 0.02fF
C617 VDD.n48 GND 0.28fF
C618 VDD.n49 GND 0.01fF
C619 VDD.n50 GND 0.02fF
C620 VDD.n51 GND 0.03fF
C621 VDD.n52 GND 0.02fF
C622 VDD.n53 GND 0.02fF
C623 VDD.n54 GND 0.02fF
C624 VDD.n55 GND 0.22fF
C625 VDD.n56 GND 0.04fF
C626 VDD.n57 GND 0.04fF
C627 VDD.n58 GND 0.02fF
C628 VDD.n60 GND 0.02fF
C629 VDD.n61 GND 0.02fF
C630 VDD.n62 GND 0.02fF
C631 VDD.n63 GND 0.02fF
C632 VDD.n65 GND 0.02fF
C633 VDD.n66 GND 0.02fF
C634 VDD.n67 GND 0.02fF
C635 VDD.n69 GND 0.28fF
C636 VDD.n71 GND 0.02fF
C637 VDD.n72 GND 0.02fF
C638 VDD.n73 GND 0.03fF
C639 VDD.n74 GND 0.02fF
C640 VDD.n75 GND 0.28fF
C641 VDD.n76 GND 0.01fF
C642 VDD.n77 GND 0.02fF
C643 VDD.n78 GND 0.03fF
C644 VDD.n79 GND 0.28fF
C645 VDD.n80 GND 0.01fF
C646 VDD.n81 GND 0.02fF
C647 VDD.n82 GND 0.02fF
C648 VDD.n83 GND 0.28fF
C649 VDD.n84 GND 0.01fF
C650 VDD.n85 GND 0.02fF
C651 VDD.n86 GND 0.02fF
C652 VDD.n87 GND 0.31fF
C653 VDD.n88 GND 0.01fF
C654 VDD.n89 GND 0.03fF
C655 VDD.n90 GND 0.03fF
C656 VDD.n91 GND 0.31fF
C657 VDD.n92 GND 0.01fF
C658 VDD.n93 GND 0.03fF
C659 VDD.n94 GND 0.03fF
C660 VDD.n95 GND 0.28fF
C661 VDD.n96 GND 0.01fF
C662 VDD.n97 GND 0.02fF
C663 VDD.n98 GND 0.02fF
C664 VDD.n99 GND 0.28fF
C665 VDD.n100 GND 0.01fF
C666 VDD.n101 GND 0.02fF
C667 VDD.n102 GND 0.02fF
C668 VDD.n103 GND 0.28fF
C669 VDD.n104 GND 0.01fF
C670 VDD.n105 GND 0.02fF
C671 VDD.n106 GND 0.03fF
C672 VDD.n107 GND 0.02fF
C673 VDD.n108 GND 0.02fF
C674 VDD.n109 GND 0.02fF
C675 VDD.n110 GND 0.22fF
C676 VDD.n111 GND 0.04fF
C677 VDD.n112 GND 0.03fF
C678 VDD.n113 GND 0.02fF
C679 VDD.n114 GND 0.02fF
C680 VDD.n115 GND 0.02fF
C681 VDD.n116 GND 0.03fF
C682 VDD.n117 GND 0.02fF
C683 VDD.n119 GND 0.02fF
C684 VDD.n120 GND 0.02fF
C685 VDD.n121 GND 0.02fF
C686 VDD.n123 GND 0.28fF
C687 VDD.n125 GND 0.02fF
C688 VDD.n126 GND 0.02fF
C689 VDD.n127 GND 0.03fF
C690 VDD.n128 GND 0.02fF
C691 VDD.n129 GND 0.28fF
C692 VDD.n130 GND 0.01fF
C693 VDD.n131 GND 0.02fF
C694 VDD.n132 GND 0.03fF
C695 VDD.n133 GND 0.06fF
C696 VDD.n134 GND 0.25fF
C697 VDD.n135 GND 0.01fF
C698 VDD.n136 GND 0.01fF
C699 VDD.n137 GND 0.02fF
C700 VDD.n138 GND 0.14fF
C701 VDD.n139 GND 0.17fF
C702 VDD.n140 GND 0.01fF
C703 VDD.n141 GND 0.02fF
C704 VDD.n142 GND 0.02fF
C705 VDD.n143 GND 0.11fF
C706 VDD.n144 GND 0.03fF
C707 VDD.n145 GND 0.31fF
C708 VDD.n146 GND 0.01fF
C709 VDD.n147 GND 0.02fF
C710 VDD.n148 GND 0.03fF
C711 VDD.n149 GND 0.17fF
C712 VDD.n150 GND 0.14fF
C713 VDD.n151 GND 0.01fF
C714 VDD.n152 GND 0.02fF
C715 VDD.n153 GND 0.03fF
C716 VDD.n154 GND 0.14fF
C717 VDD.n155 GND 0.16fF
C718 VDD.n156 GND 0.01fF
C719 VDD.n157 GND 0.02fF
C720 VDD.n158 GND 0.02fF
C721 VDD.n159 GND 0.06fF
C722 VDD.n160 GND 0.25fF
C723 VDD.n161 GND 0.01fF
C724 VDD.n162 GND 0.01fF
C725 VDD.n163 GND 0.02fF
C726 VDD.n164 GND 0.28fF
C727 VDD.n165 GND 0.01fF
C728 VDD.n166 GND 0.02fF
C729 VDD.n167 GND 0.03fF
C730 VDD.n168 GND 0.02fF
C731 VDD.n169 GND 0.02fF
C732 VDD.n170 GND 0.02fF
C733 VDD.n171 GND 0.22fF
C734 VDD.n172 GND 0.04fF
C735 VDD.n173 GND 0.03fF
C736 VDD.n174 GND 0.02fF
C737 VDD.n175 GND 0.02fF
C738 VDD.n176 GND 0.02fF
C739 VDD.n177 GND 0.03fF
C740 VDD.n178 GND 0.02fF
C741 VDD.n180 GND 0.02fF
C742 VDD.n181 GND 0.02fF
C743 VDD.n182 GND 0.02fF
C744 VDD.n184 GND 0.28fF
C745 VDD.n186 GND 0.02fF
C746 VDD.n187 GND 0.02fF
C747 VDD.n188 GND 0.03fF
C748 VDD.n189 GND 0.02fF
C749 VDD.n190 GND 0.28fF
C750 VDD.n191 GND 0.01fF
C751 VDD.n192 GND 0.02fF
C752 VDD.n193 GND 0.03fF
C753 VDD.n194 GND 0.06fF
C754 VDD.n195 GND 0.25fF
C755 VDD.n196 GND 0.01fF
C756 VDD.n197 GND 0.01fF
C757 VDD.n198 GND 0.02fF
C758 VDD.n199 GND 0.14fF
C759 VDD.n200 GND 0.17fF
C760 VDD.n201 GND 0.01fF
C761 VDD.n202 GND 0.02fF
C762 VDD.n203 GND 0.02fF
C763 VDD.n204 GND 0.11fF
C764 VDD.n205 GND 0.03fF
C765 VDD.n206 GND 0.31fF
C766 VDD.n207 GND 0.01fF
C767 VDD.n208 GND 0.02fF
C768 VDD.n209 GND 0.03fF
C769 VDD.n210 GND 0.17fF
C770 VDD.n211 GND 0.14fF
C771 VDD.n212 GND 0.01fF
C772 VDD.n213 GND 0.02fF
C773 VDD.n214 GND 0.03fF
C774 VDD.n215 GND 0.14fF
C775 VDD.n216 GND 0.16fF
C776 VDD.n217 GND 0.01fF
C777 VDD.n218 GND 0.02fF
C778 VDD.n219 GND 0.02fF
C779 VDD.n220 GND 0.06fF
C780 VDD.n221 GND 0.25fF
C781 VDD.n222 GND 0.01fF
C782 VDD.n223 GND 0.01fF
C783 VDD.n224 GND 0.02fF
C784 VDD.n225 GND 0.28fF
C785 VDD.n226 GND 0.01fF
C786 VDD.n227 GND 0.02fF
C787 VDD.n228 GND 0.03fF
C788 VDD.n229 GND 0.02fF
C789 VDD.n230 GND 0.02fF
C790 VDD.n231 GND 0.02fF
C791 VDD.n232 GND 0.26fF
C792 VDD.n233 GND 0.04fF
C793 VDD.n234 GND 0.03fF
C794 VDD.n235 GND 0.02fF
C795 VDD.n236 GND 0.02fF
C796 VDD.n237 GND 0.02fF
C797 VDD.n238 GND 0.03fF
C798 VDD.n239 GND 0.02fF
C799 VDD.n241 GND 0.02fF
C800 VDD.n242 GND 0.02fF
C801 VDD.n243 GND 0.02fF
C802 VDD.n245 GND 0.28fF
C803 VDD.n247 GND 0.02fF
C804 VDD.n248 GND 0.02fF
C805 VDD.n249 GND 0.03fF
C806 VDD.n250 GND 0.02fF
C807 VDD.n251 GND 0.28fF
C808 VDD.n252 GND 0.01fF
C809 VDD.n253 GND 0.02fF
C810 VDD.n254 GND 0.03fF
C811 VDD.n255 GND 0.28fF
C812 VDD.n256 GND 0.01fF
C813 VDD.n257 GND 0.02fF
C814 VDD.n258 GND 0.02fF
C815 VDD.n259 GND 0.22fF
C816 VDD.n260 GND 0.01fF
C817 VDD.n261 GND 0.07fF
C818 VDD.n262 GND 0.02fF
C819 VDD.n263 GND 0.14fF
C820 VDD.n264 GND 0.17fF
C821 VDD.n265 GND 0.01fF
C822 VDD.n266 GND 0.02fF
C823 VDD.n267 GND 0.02fF
C824 VDD.n268 GND 0.14fF
C825 VDD.n269 GND 0.16fF
C826 VDD.n270 GND 0.01fF
C827 VDD.n271 GND 0.11fF
C828 VDD.n272 GND 0.02fF
C829 VDD.n273 GND 0.02fF
C830 VDD.n274 GND 0.02fF
C831 VDD.n275 GND 0.18fF
C832 VDD.n276 GND 0.15fF
C833 VDD.n277 GND 0.01fF
C834 VDD.n278 GND 0.02fF
C835 VDD.n279 GND 0.03fF
C836 VDD.n280 GND 0.18fF
C837 VDD.n281 GND 0.15fF
C838 VDD.n282 GND 0.01fF
C839 VDD.n283 GND 0.02fF
C840 VDD.n284 GND 0.03fF
C841 VDD.n285 GND 0.11fF
C842 VDD.n286 GND 0.02fF
C843 VDD.n287 GND 0.14fF
C844 VDD.n288 GND 0.16fF
C845 VDD.n289 GND 0.01fF
C846 VDD.n290 GND 0.02fF
C847 VDD.n291 GND 0.02fF
C848 VDD.n292 GND 0.14fF
C849 VDD.n293 GND 0.17fF
C850 VDD.n294 GND 0.01fF
C851 VDD.n295 GND 0.02fF
C852 VDD.n296 GND 0.02fF
C853 VDD.n297 GND 0.06fF
C854 VDD.n298 GND 0.23fF
C855 VDD.n299 GND 0.01fF
C856 VDD.n300 GND 0.01fF
C857 VDD.n301 GND 0.02fF
C858 VDD.n302 GND 0.28fF
C859 VDD.n303 GND 0.01fF
C860 VDD.n304 GND 0.02fF
C861 VDD.n305 GND 0.02fF
C862 VDD.n306 GND 0.28fF
C863 VDD.n307 GND 0.01fF
C864 VDD.n308 GND 0.02fF
C865 VDD.n309 GND 0.03fF
C866 VDD.n310 GND 0.02fF
C867 VDD.n311 GND 0.02fF
C868 VDD.n312 GND 0.02fF
C869 VDD.n313 GND 0.31fF
C870 VDD.n314 GND 0.04fF
C871 VDD.n315 GND 0.03fF
C872 VDD.n316 GND 0.02fF
C873 VDD.n317 GND 0.02fF
C874 VDD.n318 GND 0.02fF
C875 VDD.n319 GND 0.03fF
C876 VDD.n320 GND 0.02fF
C877 VDD.n322 GND 0.02fF
C878 VDD.n323 GND 0.02fF
C879 VDD.n324 GND 0.02fF
C880 VDD.n326 GND 0.28fF
C881 VDD.n328 GND 0.02fF
C882 VDD.n329 GND 0.02fF
C883 VDD.n330 GND 0.03fF
C884 VDD.n331 GND 0.02fF
C885 VDD.n332 GND 0.28fF
C886 VDD.n333 GND 0.01fF
C887 VDD.n334 GND 0.02fF
C888 VDD.n335 GND 0.03fF
C889 VDD.n336 GND 0.28fF
C890 VDD.n337 GND 0.01fF
C891 VDD.n338 GND 0.02fF
C892 VDD.n339 GND 0.02fF
C893 VDD.n340 GND 0.22fF
C894 VDD.n341 GND 0.01fF
C895 VDD.n342 GND 0.07fF
C896 VDD.n343 GND 0.02fF
C897 VDD.n344 GND 0.14fF
C898 VDD.n345 GND 0.17fF
C899 VDD.n346 GND 0.01fF
C900 VDD.n347 GND 0.02fF
C901 VDD.n348 GND 0.02fF
C902 VDD.n349 GND 0.14fF
C903 VDD.n350 GND 0.16fF
C904 VDD.n351 GND 0.01fF
C905 VDD.n352 GND 0.11fF
C906 VDD.n353 GND 0.02fF
C907 VDD.n354 GND 0.02fF
C908 VDD.n355 GND 0.02fF
C909 VDD.n356 GND 0.18fF
C910 VDD.n357 GND 0.15fF
C911 VDD.n358 GND 0.01fF
C912 VDD.n359 GND 0.02fF
C913 VDD.n360 GND 0.03fF
C914 VDD.n361 GND 0.18fF
C915 VDD.n362 GND 0.15fF
C916 VDD.n363 GND 0.01fF
C917 VDD.n364 GND 0.02fF
C918 VDD.n365 GND 0.03fF
C919 VDD.n366 GND 0.11fF
C920 VDD.n367 GND 0.02fF
C921 VDD.n368 GND 0.14fF
C922 VDD.n369 GND 0.16fF
C923 VDD.n370 GND 0.01fF
C924 VDD.n371 GND 0.02fF
C925 VDD.n372 GND 0.02fF
C926 VDD.n373 GND 0.14fF
C927 VDD.n374 GND 0.17fF
C928 VDD.n375 GND 0.01fF
C929 VDD.n376 GND 0.02fF
C930 VDD.n377 GND 0.02fF
C931 VDD.n378 GND 0.06fF
C932 VDD.n379 GND 0.23fF
C933 VDD.n380 GND 0.01fF
C934 VDD.n381 GND 0.01fF
C935 VDD.n382 GND 0.02fF
C936 VDD.n383 GND 0.28fF
C937 VDD.n384 GND 0.01fF
C938 VDD.n385 GND 0.02fF
C939 VDD.n386 GND 0.02fF
C940 VDD.n387 GND 0.28fF
C941 VDD.n388 GND 0.01fF
C942 VDD.n389 GND 0.02fF
C943 VDD.n390 GND 0.03fF
C944 VDD.n391 GND 0.02fF
C945 VDD.n392 GND 0.02fF
C946 VDD.n393 GND 0.02fF
C947 VDD.n394 GND 0.26fF
C948 VDD.n395 GND 0.04fF
C949 VDD.n396 GND 0.03fF
C950 VDD.n397 GND 0.02fF
C951 VDD.n398 GND 0.02fF
C952 VDD.n399 GND 0.02fF
C953 VDD.n400 GND 0.03fF
C954 VDD.n401 GND 0.02fF
C955 VDD.n403 GND 0.02fF
C956 VDD.n404 GND 0.02fF
C957 VDD.n405 GND 0.02fF
C958 VDD.n407 GND 0.28fF
C959 VDD.n409 GND 0.02fF
C960 VDD.n410 GND 0.02fF
C961 VDD.n411 GND 0.03fF
C962 VDD.n412 GND 0.02fF
C963 VDD.n413 GND 0.28fF
C964 VDD.n414 GND 0.01fF
C965 VDD.n415 GND 0.02fF
C966 VDD.n416 GND 0.03fF
C967 VDD.n417 GND 0.06fF
C968 VDD.n418 GND 0.25fF
C969 VDD.n419 GND 0.01fF
C970 VDD.n420 GND 0.01fF
C971 VDD.n421 GND 0.02fF
C972 VDD.n422 GND 0.14fF
C973 VDD.n423 GND 0.17fF
C974 VDD.n424 GND 0.01fF
C975 VDD.n425 GND 0.02fF
C976 VDD.n426 GND 0.02fF
C977 VDD.n427 GND 0.11fF
C978 VDD.n428 GND 0.03fF
C979 VDD.n429 GND 0.31fF
C980 VDD.n430 GND 0.01fF
C981 VDD.n431 GND 0.02fF
C982 VDD.n432 GND 0.03fF
C983 VDD.n433 GND 0.17fF
C984 VDD.n434 GND 0.14fF
C985 VDD.n435 GND 0.01fF
C986 VDD.n436 GND 0.02fF
C987 VDD.n437 GND 0.03fF
C988 VDD.n438 GND 0.14fF
C989 VDD.n439 GND 0.16fF
C990 VDD.n440 GND 0.01fF
C991 VDD.n441 GND 0.02fF
C992 VDD.n442 GND 0.02fF
C993 VDD.n443 GND 0.06fF
C994 VDD.n444 GND 0.25fF
C995 VDD.n445 GND 0.01fF
C996 VDD.n446 GND 0.01fF
C997 VDD.n447 GND 0.02fF
C998 VDD.n448 GND 0.28fF
C999 VDD.n449 GND 0.01fF
C1000 VDD.n450 GND 0.02fF
C1001 VDD.n451 GND 0.03fF
C1002 VDD.n452 GND 0.02fF
C1003 VDD.n453 GND 0.02fF
C1004 VDD.n454 GND 0.02fF
C1005 VDD.n455 GND 0.26fF
C1006 VDD.n456 GND 0.04fF
C1007 VDD.n457 GND 0.03fF
C1008 VDD.n458 GND 0.02fF
C1009 VDD.n459 GND 0.02fF
C1010 VDD.n460 GND 0.02fF
C1011 VDD.n461 GND 0.03fF
C1012 VDD.n462 GND 0.02fF
C1013 VDD.n464 GND 0.02fF
C1014 VDD.n465 GND 0.02fF
C1015 VDD.n466 GND 0.02fF
C1016 VDD.n468 GND 0.28fF
C1017 VDD.n470 GND 0.02fF
C1018 VDD.n471 GND 0.02fF
C1019 VDD.n472 GND 0.03fF
C1020 VDD.n473 GND 0.02fF
C1021 VDD.n474 GND 0.28fF
C1022 VDD.n475 GND 0.01fF
C1023 VDD.n476 GND 0.02fF
C1024 VDD.n477 GND 0.03fF
C1025 VDD.n478 GND 0.28fF
C1026 VDD.n479 GND 0.01fF
C1027 VDD.n480 GND 0.02fF
C1028 VDD.n481 GND 0.02fF
C1029 VDD.n482 GND 0.22fF
C1030 VDD.n483 GND 0.01fF
C1031 VDD.n484 GND 0.07fF
C1032 VDD.n485 GND 0.02fF
C1033 VDD.n486 GND 0.14fF
C1034 VDD.n487 GND 0.17fF
C1035 VDD.n488 GND 0.01fF
C1036 VDD.n489 GND 0.02fF
C1037 VDD.n490 GND 0.02fF
C1038 VDD.n491 GND 0.14fF
C1039 VDD.n492 GND 0.16fF
C1040 VDD.n493 GND 0.01fF
C1041 VDD.n494 GND 0.11fF
C1042 VDD.n495 GND 0.02fF
C1043 VDD.n496 GND 0.02fF
C1044 VDD.n497 GND 0.02fF
C1045 VDD.n498 GND 0.18fF
C1046 VDD.n499 GND 0.15fF
C1047 VDD.n500 GND 0.01fF
C1048 VDD.n501 GND 0.02fF
C1049 VDD.n502 GND 0.03fF
C1050 VDD.n503 GND 0.18fF
C1051 VDD.n504 GND 0.15fF
C1052 VDD.n505 GND 0.01fF
C1053 VDD.n506 GND 0.02fF
C1054 VDD.n507 GND 0.03fF
C1055 VDD.n508 GND 0.11fF
C1056 VDD.n509 GND 0.02fF
C1057 VDD.n510 GND 0.14fF
C1058 VDD.n511 GND 0.16fF
C1059 VDD.n512 GND 0.01fF
C1060 VDD.n513 GND 0.02fF
C1061 VDD.n514 GND 0.02fF
C1062 VDD.n515 GND 0.14fF
C1063 VDD.n516 GND 0.17fF
C1064 VDD.n517 GND 0.01fF
C1065 VDD.n518 GND 0.02fF
C1066 VDD.n519 GND 0.02fF
C1067 VDD.n520 GND 0.06fF
C1068 VDD.n521 GND 0.23fF
C1069 VDD.n522 GND 0.01fF
C1070 VDD.n523 GND 0.01fF
C1071 VDD.n524 GND 0.02fF
C1072 VDD.n525 GND 0.28fF
C1073 VDD.n526 GND 0.01fF
C1074 VDD.n527 GND 0.02fF
C1075 VDD.n528 GND 0.02fF
C1076 VDD.n529 GND 0.28fF
C1077 VDD.n530 GND 0.01fF
C1078 VDD.n531 GND 0.02fF
C1079 VDD.n532 GND 0.03fF
C1080 VDD.n533 GND 0.02fF
C1081 VDD.n534 GND 0.02fF
C1082 VDD.n535 GND 0.02fF
C1083 VDD.n536 GND 0.31fF
C1084 VDD.n537 GND 0.04fF
C1085 VDD.n538 GND 0.03fF
C1086 VDD.n539 GND 0.02fF
C1087 VDD.n540 GND 0.02fF
C1088 VDD.n541 GND 0.02fF
C1089 VDD.n542 GND 0.03fF
C1090 VDD.n543 GND 0.02fF
C1091 VDD.n545 GND 0.02fF
C1092 VDD.n546 GND 0.02fF
C1093 VDD.n547 GND 0.02fF
C1094 VDD.n549 GND 0.28fF
C1095 VDD.n551 GND 0.02fF
C1096 VDD.n552 GND 0.02fF
C1097 VDD.n553 GND 0.03fF
C1098 VDD.n554 GND 0.02fF
C1099 VDD.n555 GND 0.28fF
C1100 VDD.n556 GND 0.01fF
C1101 VDD.n557 GND 0.02fF
C1102 VDD.n558 GND 0.03fF
C1103 VDD.n559 GND 0.28fF
C1104 VDD.n560 GND 0.01fF
C1105 VDD.n561 GND 0.02fF
C1106 VDD.n562 GND 0.02fF
C1107 VDD.n563 GND 0.22fF
C1108 VDD.n564 GND 0.01fF
C1109 VDD.n565 GND 0.07fF
C1110 VDD.n566 GND 0.02fF
C1111 VDD.n567 GND 0.14fF
C1112 VDD.n568 GND 0.17fF
C1113 VDD.n569 GND 0.01fF
C1114 VDD.n570 GND 0.02fF
C1115 VDD.n571 GND 0.02fF
C1116 VDD.n572 GND 0.14fF
C1117 VDD.n573 GND 0.16fF
C1118 VDD.n574 GND 0.01fF
C1119 VDD.n575 GND 0.11fF
C1120 VDD.n576 GND 0.02fF
C1121 VDD.n577 GND 0.02fF
C1122 VDD.n578 GND 0.02fF
C1123 VDD.n579 GND 0.18fF
C1124 VDD.n580 GND 0.15fF
C1125 VDD.n581 GND 0.01fF
C1126 VDD.n582 GND 0.02fF
C1127 VDD.n583 GND 0.03fF
C1128 VDD.n584 GND 0.18fF
C1129 VDD.n585 GND 0.15fF
C1130 VDD.n586 GND 0.01fF
C1131 VDD.n587 GND 0.02fF
C1132 VDD.n588 GND 0.03fF
C1133 VDD.n589 GND 0.11fF
C1134 VDD.n590 GND 0.02fF
C1135 VDD.n591 GND 0.14fF
C1136 VDD.n592 GND 0.16fF
C1137 VDD.n593 GND 0.01fF
C1138 VDD.n594 GND 0.02fF
C1139 VDD.n595 GND 0.02fF
C1140 VDD.n596 GND 0.14fF
C1141 VDD.n597 GND 0.17fF
C1142 VDD.n598 GND 0.01fF
C1143 VDD.n599 GND 0.02fF
C1144 VDD.n600 GND 0.02fF
C1145 VDD.n601 GND 0.06fF
C1146 VDD.n602 GND 0.23fF
C1147 VDD.n603 GND 0.01fF
C1148 VDD.n604 GND 0.01fF
C1149 VDD.n605 GND 0.02fF
C1150 VDD.n606 GND 0.28fF
C1151 VDD.n607 GND 0.01fF
C1152 VDD.n608 GND 0.02fF
C1153 VDD.n609 GND 0.02fF
C1154 VDD.n610 GND 0.28fF
C1155 VDD.n611 GND 0.01fF
C1156 VDD.n612 GND 0.02fF
C1157 VDD.n613 GND 0.03fF
C1158 VDD.n614 GND 0.02fF
C1159 VDD.n615 GND 0.02fF
C1160 VDD.n616 GND 0.02fF
C1161 VDD.n617 GND 0.26fF
C1162 VDD.n618 GND 0.04fF
C1163 VDD.n619 GND 0.03fF
C1164 VDD.n620 GND 0.02fF
C1165 VDD.n621 GND 0.02fF
C1166 VDD.n622 GND 0.02fF
C1167 VDD.n623 GND 0.03fF
C1168 VDD.n624 GND 0.02fF
C1169 VDD.n626 GND 0.02fF
C1170 VDD.n627 GND 0.02fF
C1171 VDD.n628 GND 0.02fF
C1172 VDD.n630 GND 0.28fF
C1173 VDD.n632 GND 0.02fF
C1174 VDD.n633 GND 0.02fF
C1175 VDD.n634 GND 0.03fF
C1176 VDD.n635 GND 0.02fF
C1177 VDD.n636 GND 0.28fF
C1178 VDD.n637 GND 0.01fF
C1179 VDD.n638 GND 0.02fF
C1180 VDD.n639 GND 0.03fF
C1181 VDD.n640 GND 0.06fF
C1182 VDD.n641 GND 0.25fF
C1183 VDD.n642 GND 0.01fF
C1184 VDD.n643 GND 0.01fF
C1185 VDD.n644 GND 0.02fF
C1186 VDD.n645 GND 0.14fF
C1187 VDD.n646 GND 0.17fF
C1188 VDD.n647 GND 0.01fF
C1189 VDD.n648 GND 0.02fF
C1190 VDD.n649 GND 0.02fF
C1191 VDD.n650 GND 0.11fF
C1192 VDD.n651 GND 0.03fF
C1193 VDD.n652 GND 0.31fF
C1194 VDD.n653 GND 0.01fF
C1195 VDD.n654 GND 0.02fF
C1196 VDD.n655 GND 0.03fF
C1197 VDD.n656 GND 0.17fF
C1198 VDD.n657 GND 0.14fF
C1199 VDD.n658 GND 0.01fF
C1200 VDD.n659 GND 0.02fF
C1201 VDD.n660 GND 0.03fF
C1202 VDD.n661 GND 0.14fF
C1203 VDD.n662 GND 0.16fF
C1204 VDD.n663 GND 0.01fF
C1205 VDD.n664 GND 0.02fF
C1206 VDD.n665 GND 0.02fF
C1207 VDD.n666 GND 0.06fF
C1208 VDD.n667 GND 0.25fF
C1209 VDD.n668 GND 0.01fF
C1210 VDD.n669 GND 0.01fF
C1211 VDD.n670 GND 0.02fF
C1212 VDD.n671 GND 0.28fF
C1213 VDD.n672 GND 0.01fF
C1214 VDD.n673 GND 0.02fF
C1215 VDD.n674 GND 0.03fF
C1216 VDD.n675 GND 0.02fF
C1217 VDD.n676 GND 0.02fF
C1218 VDD.n677 GND 0.02fF
C1219 VDD.n678 GND 0.26fF
C1220 VDD.n679 GND 0.04fF
C1221 VDD.n680 GND 0.03fF
C1222 VDD.n681 GND 0.02fF
C1223 VDD.n682 GND 0.02fF
C1224 VDD.n683 GND 0.02fF
C1225 VDD.n684 GND 0.03fF
C1226 VDD.n685 GND 0.02fF
C1227 VDD.n687 GND 0.02fF
C1228 VDD.n688 GND 0.02fF
C1229 VDD.n689 GND 0.02fF
C1230 VDD.n691 GND 0.28fF
C1231 VDD.n693 GND 0.02fF
C1232 VDD.n694 GND 0.02fF
C1233 VDD.n695 GND 0.03fF
C1234 VDD.n696 GND 0.02fF
C1235 VDD.n697 GND 0.28fF
C1236 VDD.n698 GND 0.01fF
C1237 VDD.n699 GND 0.02fF
C1238 VDD.n700 GND 0.03fF
C1239 VDD.n701 GND 0.28fF
C1240 VDD.n702 GND 0.01fF
C1241 VDD.n703 GND 0.02fF
C1242 VDD.n704 GND 0.02fF
C1243 VDD.n705 GND 0.22fF
C1244 VDD.n706 GND 0.01fF
C1245 VDD.n707 GND 0.07fF
C1246 VDD.n708 GND 0.02fF
C1247 VDD.n709 GND 0.14fF
C1248 VDD.n710 GND 0.17fF
C1249 VDD.n711 GND 0.01fF
C1250 VDD.n712 GND 0.02fF
C1251 VDD.n713 GND 0.02fF
C1252 VDD.n714 GND 0.14fF
C1253 VDD.n715 GND 0.16fF
C1254 VDD.n716 GND 0.01fF
C1255 VDD.n717 GND 0.11fF
C1256 VDD.n718 GND 0.02fF
C1257 VDD.n719 GND 0.02fF
C1258 VDD.n720 GND 0.02fF
C1259 VDD.n721 GND 0.18fF
C1260 VDD.n722 GND 0.15fF
C1261 VDD.n723 GND 0.01fF
C1262 VDD.n724 GND 0.02fF
C1263 VDD.n725 GND 0.03fF
C1264 VDD.n726 GND 0.18fF
C1265 VDD.n727 GND 0.15fF
C1266 VDD.n728 GND 0.01fF
C1267 VDD.n729 GND 0.02fF
C1268 VDD.n730 GND 0.03fF
C1269 VDD.n731 GND 0.11fF
C1270 VDD.n732 GND 0.02fF
C1271 VDD.n733 GND 0.14fF
C1272 VDD.n734 GND 0.16fF
C1273 VDD.n735 GND 0.01fF
C1274 VDD.n736 GND 0.02fF
C1275 VDD.n737 GND 0.02fF
C1276 VDD.n738 GND 0.14fF
C1277 VDD.n739 GND 0.17fF
C1278 VDD.n740 GND 0.01fF
C1279 VDD.n741 GND 0.02fF
C1280 VDD.n742 GND 0.02fF
C1281 VDD.n743 GND 0.06fF
C1282 VDD.n744 GND 0.23fF
C1283 VDD.n745 GND 0.01fF
C1284 VDD.n746 GND 0.01fF
C1285 VDD.n747 GND 0.02fF
C1286 VDD.n748 GND 0.28fF
C1287 VDD.n749 GND 0.01fF
C1288 VDD.n750 GND 0.02fF
C1289 VDD.n751 GND 0.02fF
C1290 VDD.n752 GND 0.02fF
C1291 VDD.n753 GND 0.02fF
C1292 VDD.n754 GND 0.02fF
C1293 VDD.n755 GND 0.31fF
C1294 VDD.n756 GND 0.04fF
C1295 VDD.n757 GND 0.03fF
C1296 VDD.n758 GND 0.02fF
C1297 VDD.n759 GND 0.02fF
C1298 VDD.n760 GND 0.02fF
C1299 VDD.n761 GND 0.03fF
C1300 VDD.n762 GND 0.02fF
C1301 VDD.n764 GND 0.02fF
C1302 VDD.n765 GND 0.02fF
C1303 VDD.n766 GND 0.02fF
C1304 VDD.n768 GND 0.28fF
C1305 VDD.n770 GND 0.02fF
C1306 VDD.n771 GND 0.02fF
C1307 VDD.n772 GND 0.03fF
C1308 VDD.n773 GND 0.02fF
C1309 VDD.n774 GND 0.28fF
C1310 VDD.n775 GND 0.01fF
C1311 VDD.n776 GND 0.02fF
C1312 VDD.n777 GND 0.02fF
C1313 VDD.n778 GND 0.02fF
C1314 VDD.n779 GND 0.02fF
C1315 VDD.n780 GND 0.02fF
C1316 VDD.n781 GND 0.20fF
C1317 VDD.n782 GND 0.03fF
C1318 VDD.n783 GND 0.02fF
C1319 VDD.n784 GND 0.02fF
C1320 VDD.n785 GND 0.02fF
C1321 VDD.n786 GND 0.03fF
C1322 VDD.n787 GND 0.02fF
C1323 VDD.n789 GND 0.02fF
C1324 VDD.n790 GND 0.02fF
C1325 VDD.n791 GND 0.02fF
C1326 VDD.n793 GND 0.46fF
C1327 VDD.n795 GND 0.03fF
C1328 VDD.n796 GND 0.04fF
C1329 VDD.n797 GND 0.28fF
C1330 VDD.n798 GND 0.02fF
C1331 VDD.n799 GND 0.03fF
C1332 VDD.n800 GND 0.03fF
C1333 VDD.n801 GND 0.28fF
C1334 VDD.n802 GND 0.01fF
C1335 VDD.n803 GND 0.02fF
C1336 VDD.n804 GND 0.02fF
C1337 VDD.n805 GND 0.06fF
C1338 VDD.n806 GND 0.23fF
C1339 VDD.n807 GND 0.01fF
C1340 VDD.n808 GND 0.01fF
C1341 VDD.n809 GND 0.02fF
C1342 VDD.n810 GND 0.14fF
C1343 VDD.n811 GND 0.17fF
C1344 VDD.n812 GND 0.01fF
C1345 VDD.n813 GND 0.02fF
C1346 VDD.n814 GND 0.02fF
C1347 VDD.n815 GND 0.11fF
C1348 VDD.n816 GND 0.02fF
C1349 VDD.n817 GND 0.14fF
C1350 VDD.n818 GND 0.16fF
C1351 VDD.n819 GND 0.01fF
C1352 VDD.n820 GND 0.02fF
C1353 VDD.n821 GND 0.02fF
C1354 VDD.n822 GND 0.18fF
C1355 VDD.n823 GND 0.15fF
C1356 VDD.n824 GND 0.01fF
C1357 VDD.n825 GND 0.02fF
C1358 VDD.n826 GND 0.03fF
C1359 VDD.n827 GND 0.18fF
C1360 VDD.n828 GND 0.15fF
C1361 VDD.n829 GND 0.01fF
C1362 VDD.n830 GND 0.02fF
C1363 VDD.n831 GND 0.03fF
C1364 VDD.n832 GND 0.14fF
C1365 VDD.n833 GND 0.16fF
C1366 VDD.n834 GND 0.01fF
C1367 VDD.n835 GND 0.11fF
C1368 VDD.n836 GND 0.02fF
C1369 VDD.n837 GND 0.02fF
C1370 VDD.n838 GND 0.02fF
C1371 VDD.n839 GND 0.14fF
C1372 VDD.n840 GND 0.17fF
C1373 VDD.n841 GND 0.01fF
C1374 VDD.n842 GND 0.02fF
C1375 VDD.n843 GND 0.02fF
C1376 VDD.n844 GND 0.22fF
C1377 VDD.n845 GND 0.01fF
C1378 VDD.n846 GND 0.07fF
C1379 VDD.n847 GND 0.02fF
C1380 VDD.n848 GND 0.28fF
C1381 VDD.n849 GND 0.01fF
C1382 VDD.n850 GND 0.02fF
C1383 VDD.n851 GND 0.02fF
C1384 VDD.n852 GND 0.28fF
C1385 VDD.n853 GND 0.01fF
C1386 VDD.n854 GND 0.02fF
C1387 VDD.n855 GND 0.03fF
C1388 VDD.n856 GND 0.02fF
C1389 VDD.n857 GND 0.02fF
C1390 VDD.n858 GND 0.02fF
C1391 VDD.n859 GND 0.02fF
C1392 VDD.n860 GND 0.02fF
C1393 VDD.n861 GND 0.02fF
C1394 VDD.n863 GND 0.02fF
C1395 VDD.n864 GND 0.02fF
C1396 VDD.n865 GND 0.02fF
C1397 VDD.n866 GND 0.02fF
C1398 VDD.n868 GND 0.04fF
C1399 VDD.n869 GND 0.02fF
C1400 VDD.n870 GND 0.31fF
C1401 VDD.n871 GND 0.04fF
C1402 VDD.n873 GND 0.28fF
C1403 VDD.n875 GND 0.02fF
C1404 VDD.n876 GND 0.02fF
C1405 VDD.n877 GND 0.03fF
C1406 VDD.n878 GND 0.02fF
C1407 VDD.n879 GND 0.28fF
C1408 VDD.n880 GND 0.01fF
C1409 VDD.n881 GND 0.02fF
C1410 VDD.n882 GND 0.03fF
C1411 VDD.n883 GND 0.28fF
C1412 VDD.n884 GND 0.01fF
C1413 VDD.n885 GND 0.02fF
C1414 VDD.n886 GND 0.02fF
C1415 VDD.n887 GND 0.06fF
C1416 VDD.n888 GND 0.23fF
C1417 VDD.n889 GND 0.01fF
C1418 VDD.n890 GND 0.01fF
C1419 VDD.n891 GND 0.02fF
C1420 VDD.n892 GND 0.14fF
C1421 VDD.n893 GND 0.17fF
C1422 VDD.n894 GND 0.01fF
C1423 VDD.n895 GND 0.02fF
C1424 VDD.n896 GND 0.02fF
C1425 VDD.n897 GND 0.11fF
C1426 VDD.n898 GND 0.02fF
C1427 VDD.n899 GND 0.14fF
C1428 VDD.n900 GND 0.16fF
C1429 VDD.n901 GND 0.01fF
C1430 VDD.n902 GND 0.02fF
C1431 VDD.n903 GND 0.02fF
C1432 VDD.n904 GND 0.18fF
C1433 VDD.n905 GND 0.15fF
C1434 VDD.n906 GND 0.01fF
C1435 VDD.n907 GND 0.02fF
C1436 VDD.n908 GND 0.03fF
C1437 VDD.n909 GND 0.18fF
C1438 VDD.n910 GND 0.15fF
C1439 VDD.n911 GND 0.01fF
C1440 VDD.n912 GND 0.02fF
C1441 VDD.n913 GND 0.03fF
C1442 VDD.n914 GND 0.14fF
C1443 VDD.n915 GND 0.16fF
C1444 VDD.n916 GND 0.01fF
C1445 VDD.n917 GND 0.11fF
C1446 VDD.n918 GND 0.02fF
C1447 VDD.n919 GND 0.02fF
C1448 VDD.n920 GND 0.02fF
C1449 VDD.n921 GND 0.14fF
C1450 VDD.n922 GND 0.17fF
C1451 VDD.n923 GND 0.01fF
C1452 VDD.n924 GND 0.02fF
C1453 VDD.n925 GND 0.02fF
C1454 VDD.n926 GND 0.22fF
C1455 VDD.n927 GND 0.01fF
C1456 VDD.n928 GND 0.07fF
C1457 VDD.n929 GND 0.02fF
C1458 VDD.n930 GND 0.28fF
C1459 VDD.n931 GND 0.01fF
C1460 VDD.n932 GND 0.02fF
C1461 VDD.n933 GND 0.02fF
C1462 VDD.n934 GND 0.28fF
C1463 VDD.n935 GND 0.01fF
C1464 VDD.n936 GND 0.02fF
C1465 VDD.n937 GND 0.03fF
C1466 VDD.n938 GND 0.02fF
C1467 VDD.n939 GND 0.02fF
C1468 VDD.n940 GND 0.02fF
C1469 VDD.n941 GND 0.26fF
C1470 VDD.n942 GND 0.04fF
C1471 VDD.n943 GND 0.03fF
C1472 VDD.n944 GND 0.02fF
C1473 VDD.n945 GND 0.02fF
C1474 VDD.n946 GND 0.02fF
C1475 VDD.n947 GND 0.03fF
C1476 VDD.n948 GND 0.02fF
C1477 VDD.n950 GND 0.02fF
C1478 VDD.n951 GND 0.02fF
C1479 VDD.n952 GND 0.02fF
C1480 VDD.n954 GND 0.28fF
C1481 VDD.n956 GND 0.02fF
C1482 VDD.n957 GND 0.02fF
C1483 VDD.n958 GND 0.03fF
C1484 VDD.n959 GND 0.02fF
C1485 VDD.n960 GND 0.28fF
C1486 VDD.n961 GND 0.01fF
C1487 VDD.n962 GND 0.02fF
C1488 VDD.n963 GND 0.03fF
C1489 VDD.n964 GND 0.06fF
C1490 VDD.n965 GND 0.25fF
C1491 VDD.n966 GND 0.01fF
C1492 VDD.n967 GND 0.01fF
C1493 VDD.n968 GND 0.02fF
C1494 VDD.n969 GND 0.14fF
C1495 VDD.n970 GND 0.16fF
C1496 VDD.n971 GND 0.01fF
C1497 VDD.n972 GND 0.02fF
C1498 VDD.n973 GND 0.02fF
C1499 VDD.n974 GND 0.17fF
C1500 VDD.n975 GND 0.14fF
C1501 VDD.n976 GND 0.01fF
C1502 VDD.n977 GND 0.02fF
C1503 VDD.n978 GND 0.03fF
C1504 VDD.n979 GND 0.11fF
C1505 VDD.n980 GND 0.03fF
C1506 VDD.n981 GND 0.31fF
C1507 VDD.n982 GND 0.01fF
C1508 VDD.n983 GND 0.02fF
C1509 VDD.n984 GND 0.03fF
C1510 VDD.n985 GND 0.14fF
C1511 VDD.n986 GND 0.17fF
C1512 VDD.n987 GND 0.01fF
C1513 VDD.n988 GND 0.02fF
C1514 VDD.n989 GND 0.02fF
C1515 VDD.n990 GND 0.06fF
C1516 VDD.n991 GND 0.25fF
C1517 VDD.n992 GND 0.01fF
C1518 VDD.n993 GND 0.01fF
C1519 VDD.n994 GND 0.02fF
C1520 VDD.n995 GND 0.28fF
C1521 VDD.n996 GND 0.01fF
C1522 VDD.n997 GND 0.02fF
C1523 VDD.n998 GND 0.03fF
C1524 VDD.n999 GND 0.02fF
C1525 VDD.n1000 GND 0.02fF
C1526 VDD.n1001 GND 0.02fF
C1527 VDD.n1002 GND 0.26fF
C1528 VDD.n1003 GND 0.04fF
C1529 VDD.n1004 GND 0.03fF
C1530 VDD.n1005 GND 0.02fF
C1531 VDD.n1006 GND 0.02fF
C1532 VDD.n1007 GND 0.02fF
C1533 VDD.n1008 GND 0.03fF
C1534 VDD.n1009 GND 0.02fF
C1535 VDD.n1011 GND 0.02fF
C1536 VDD.n1012 GND 0.02fF
C1537 VDD.n1013 GND 0.02fF
C1538 VDD.n1015 GND 0.28fF
C1539 VDD.n1017 GND 0.02fF
C1540 VDD.n1018 GND 0.02fF
C1541 VDD.n1019 GND 0.03fF
C1542 VDD.n1020 GND 0.02fF
C1543 VDD.n1021 GND 0.28fF
C1544 VDD.n1022 GND 0.01fF
C1545 VDD.n1023 GND 0.02fF
C1546 VDD.n1024 GND 0.03fF
C1547 VDD.n1025 GND 0.28fF
C1548 VDD.n1026 GND 0.01fF
C1549 VDD.n1027 GND 0.02fF
C1550 VDD.n1028 GND 0.02fF
C1551 VDD.n1029 GND 0.06fF
C1552 VDD.n1030 GND 0.23fF
C1553 VDD.n1031 GND 0.01fF
C1554 VDD.n1032 GND 0.01fF
C1555 VDD.n1033 GND 0.02fF
C1556 VDD.n1034 GND 0.14fF
C1557 VDD.n1035 GND 0.17fF
C1558 VDD.n1036 GND 0.01fF
C1559 VDD.n1037 GND 0.02fF
C1560 VDD.n1038 GND 0.02fF
C1561 VDD.n1039 GND 0.11fF
C1562 VDD.n1040 GND 0.02fF
C1563 VDD.n1041 GND 0.14fF
C1564 VDD.n1042 GND 0.16fF
C1565 VDD.n1043 GND 0.01fF
C1566 VDD.n1044 GND 0.02fF
C1567 VDD.n1045 GND 0.02fF
C1568 VDD.n1046 GND 0.18fF
C1569 VDD.n1047 GND 0.15fF
C1570 VDD.n1048 GND 0.01fF
C1571 VDD.n1049 GND 0.02fF
C1572 VDD.n1050 GND 0.03fF
C1573 VDD.n1051 GND 0.18fF
C1574 VDD.n1052 GND 0.15fF
C1575 VDD.n1053 GND 0.01fF
C1576 VDD.n1054 GND 0.02fF
C1577 VDD.n1055 GND 0.03fF
C1578 VDD.n1056 GND 0.14fF
C1579 VDD.n1057 GND 0.16fF
C1580 VDD.n1058 GND 0.01fF
C1581 VDD.n1059 GND 0.11fF
C1582 VDD.n1060 GND 0.02fF
C1583 VDD.n1061 GND 0.02fF
C1584 VDD.n1062 GND 0.02fF
C1585 VDD.n1063 GND 0.14fF
C1586 VDD.n1064 GND 0.17fF
C1587 VDD.n1065 GND 0.01fF
C1588 VDD.n1066 GND 0.02fF
C1589 VDD.n1067 GND 0.02fF
C1590 VDD.n1068 GND 0.22fF
C1591 VDD.n1069 GND 0.01fF
C1592 VDD.n1070 GND 0.07fF
C1593 VDD.n1071 GND 0.02fF
C1594 VDD.n1072 GND 0.28fF
C1595 VDD.n1073 GND 0.01fF
C1596 VDD.n1074 GND 0.02fF
C1597 VDD.n1075 GND 0.02fF
C1598 VDD.n1076 GND 0.28fF
C1599 VDD.n1077 GND 0.01fF
C1600 VDD.n1078 GND 0.02fF
C1601 VDD.n1079 GND 0.03fF
C1602 VDD.n1080 GND 0.02fF
C1603 VDD.n1081 GND 0.02fF
C1604 VDD.n1082 GND 0.02fF
C1605 VDD.n1083 GND 0.31fF
C1606 VDD.n1084 GND 0.04fF
C1607 VDD.n1085 GND 0.03fF
C1608 VDD.n1086 GND 0.02fF
C1609 VDD.n1087 GND 0.02fF
C1610 VDD.n1088 GND 0.02fF
C1611 VDD.n1089 GND 0.03fF
C1612 VDD.n1090 GND 0.02fF
C1613 VDD.n1092 GND 0.02fF
C1614 VDD.n1093 GND 0.02fF
C1615 VDD.n1094 GND 0.02fF
C1616 VDD.n1096 GND 0.28fF
C1617 VDD.n1098 GND 0.02fF
C1618 VDD.n1099 GND 0.02fF
C1619 VDD.n1100 GND 0.03fF
C1620 VDD.n1101 GND 0.02fF
C1621 VDD.n1102 GND 0.28fF
C1622 VDD.n1103 GND 0.01fF
C1623 VDD.n1104 GND 0.02fF
C1624 VDD.n1105 GND 0.03fF
C1625 VDD.n1106 GND 0.28fF
C1626 VDD.n1107 GND 0.01fF
C1627 VDD.n1108 GND 0.02fF
C1628 VDD.n1109 GND 0.02fF
C1629 VDD.n1110 GND 0.06fF
C1630 VDD.n1111 GND 0.23fF
C1631 VDD.n1112 GND 0.01fF
C1632 VDD.n1113 GND 0.01fF
C1633 VDD.n1114 GND 0.02fF
C1634 VDD.n1115 GND 0.14fF
C1635 VDD.n1116 GND 0.17fF
C1636 VDD.n1117 GND 0.01fF
C1637 VDD.n1118 GND 0.02fF
C1638 VDD.n1119 GND 0.02fF
C1639 VDD.n1120 GND 0.11fF
C1640 VDD.n1121 GND 0.02fF
C1641 VDD.n1122 GND 0.14fF
C1642 VDD.n1123 GND 0.16fF
C1643 VDD.n1124 GND 0.01fF
C1644 VDD.n1125 GND 0.02fF
C1645 VDD.n1126 GND 0.02fF
C1646 VDD.n1127 GND 0.18fF
C1647 VDD.n1128 GND 0.15fF
C1648 VDD.n1129 GND 0.01fF
C1649 VDD.n1130 GND 0.02fF
C1650 VDD.n1131 GND 0.03fF
C1651 VDD.n1132 GND 0.18fF
C1652 VDD.n1133 GND 0.15fF
C1653 VDD.n1134 GND 0.01fF
C1654 VDD.n1135 GND 0.02fF
C1655 VDD.n1136 GND 0.03fF
C1656 VDD.n1137 GND 0.14fF
C1657 VDD.n1138 GND 0.16fF
C1658 VDD.n1139 GND 0.01fF
C1659 VDD.n1140 GND 0.11fF
C1660 VDD.n1141 GND 0.02fF
C1661 VDD.n1142 GND 0.02fF
C1662 VDD.n1143 GND 0.02fF
C1663 VDD.n1144 GND 0.14fF
C1664 VDD.n1145 GND 0.17fF
C1665 VDD.n1146 GND 0.01fF
C1666 VDD.n1147 GND 0.02fF
C1667 VDD.n1148 GND 0.02fF
C1668 VDD.n1149 GND 0.22fF
C1669 VDD.n1150 GND 0.01fF
C1670 VDD.n1151 GND 0.07fF
C1671 VDD.n1152 GND 0.02fF
C1672 VDD.n1153 GND 0.28fF
C1673 VDD.n1154 GND 0.01fF
C1674 VDD.n1155 GND 0.02fF
C1675 VDD.n1156 GND 0.02fF
C1676 VDD.n1157 GND 0.28fF
C1677 VDD.n1158 GND 0.01fF
C1678 VDD.n1159 GND 0.02fF
C1679 VDD.n1160 GND 0.03fF
C1680 VDD.n1161 GND 0.02fF
C1681 VDD.n1162 GND 0.02fF
C1682 VDD.n1163 GND 0.02fF
C1683 VDD.n1164 GND 0.26fF
C1684 VDD.n1165 GND 0.04fF
C1685 VDD.n1166 GND 0.03fF
C1686 VDD.n1167 GND 0.02fF
C1687 VDD.n1168 GND 0.02fF
C1688 VDD.n1169 GND 0.02fF
C1689 VDD.n1170 GND 0.03fF
C1690 VDD.n1171 GND 0.02fF
C1691 VDD.n1173 GND 0.02fF
C1692 VDD.n1174 GND 0.02fF
C1693 VDD.n1175 GND 0.02fF
C1694 VDD.n1177 GND 0.28fF
C1695 VDD.n1179 GND 0.02fF
C1696 VDD.n1180 GND 0.02fF
C1697 VDD.n1181 GND 0.03fF
C1698 VDD.n1182 GND 0.02fF
C1699 VDD.n1183 GND 0.28fF
C1700 VDD.n1184 GND 0.01fF
C1701 VDD.n1185 GND 0.02fF
C1702 VDD.n1186 GND 0.03fF
C1703 VDD.n1187 GND 0.06fF
C1704 VDD.n1188 GND 0.25fF
C1705 VDD.n1189 GND 0.01fF
C1706 VDD.n1190 GND 0.01fF
C1707 VDD.n1191 GND 0.02fF
C1708 VDD.n1192 GND 0.14fF
C1709 VDD.n1193 GND 0.16fF
C1710 VDD.n1194 GND 0.01fF
C1711 VDD.n1195 GND 0.02fF
C1712 VDD.n1196 GND 0.02fF
C1713 VDD.n1197 GND 0.17fF
C1714 VDD.n1198 GND 0.14fF
C1715 VDD.n1199 GND 0.01fF
C1716 VDD.n1200 GND 0.02fF
C1717 VDD.n1201 GND 0.03fF
C1718 VDD.n1202 GND 0.11fF
C1719 VDD.n1203 GND 0.03fF
C1720 VDD.n1204 GND 0.31fF
C1721 VDD.n1205 GND 0.01fF
C1722 VDD.n1206 GND 0.02fF
C1723 VDD.n1207 GND 0.03fF
C1724 VDD.n1208 GND 0.14fF
C1725 VDD.n1209 GND 0.17fF
C1726 VDD.n1210 GND 0.01fF
C1727 VDD.n1211 GND 0.02fF
C1728 VDD.n1212 GND 0.02fF
C1729 VDD.n1213 GND 0.06fF
C1730 VDD.n1214 GND 0.25fF
C1731 VDD.n1215 GND 0.01fF
C1732 VDD.n1216 GND 0.01fF
C1733 VDD.n1217 GND 0.02fF
C1734 VDD.n1218 GND 0.28fF
C1735 VDD.n1219 GND 0.01fF
C1736 VDD.n1220 GND 0.02fF
C1737 VDD.n1221 GND 0.03fF
C1738 VDD.n1222 GND 0.02fF
C1739 VDD.n1223 GND 0.02fF
C1740 VDD.n1224 GND 0.02fF
C1741 VDD.n1225 GND 0.26fF
C1742 VDD.n1226 GND 0.04fF
C1743 VDD.n1227 GND 0.03fF
C1744 VDD.n1228 GND 0.02fF
C1745 VDD.n1229 GND 0.02fF
C1746 VDD.n1230 GND 0.02fF
C1747 VDD.n1231 GND 0.03fF
C1748 VDD.n1232 GND 0.02fF
C1749 VDD.n1234 GND 0.02fF
C1750 VDD.n1235 GND 0.02fF
C1751 VDD.n1236 GND 0.02fF
C1752 VDD.n1238 GND 0.28fF
C1753 VDD.n1240 GND 0.02fF
C1754 VDD.n1241 GND 0.02fF
C1755 VDD.n1242 GND 0.03fF
C1756 VDD.n1243 GND 0.02fF
C1757 VDD.n1244 GND 0.28fF
C1758 VDD.n1245 GND 0.01fF
C1759 VDD.n1246 GND 0.02fF
C1760 VDD.n1247 GND 0.03fF
C1761 VDD.n1248 GND 0.28fF
C1762 VDD.n1249 GND 0.01fF
C1763 VDD.n1250 GND 0.02fF
C1764 VDD.n1251 GND 0.02fF
C1765 VDD.n1252 GND 0.06fF
C1766 VDD.n1253 GND 0.23fF
C1767 VDD.n1254 GND 0.01fF
C1768 VDD.n1255 GND 0.01fF
C1769 VDD.n1256 GND 0.02fF
C1770 VDD.n1257 GND 0.14fF
C1771 VDD.n1258 GND 0.17fF
C1772 VDD.n1259 GND 0.01fF
C1773 VDD.n1260 GND 0.02fF
C1774 VDD.n1261 GND 0.02fF
C1775 VDD.n1262 GND 0.11fF
C1776 VDD.n1263 GND 0.02fF
C1777 VDD.n1264 GND 0.14fF
C1778 VDD.n1265 GND 0.16fF
C1779 VDD.n1266 GND 0.01fF
C1780 VDD.n1267 GND 0.02fF
C1781 VDD.n1268 GND 0.02fF
C1782 VDD.n1269 GND 0.18fF
C1783 VDD.n1270 GND 0.15fF
C1784 VDD.n1271 GND 0.01fF
C1785 VDD.n1272 GND 0.02fF
C1786 VDD.n1273 GND 0.03fF
C1787 VDD.n1274 GND 0.18fF
C1788 VDD.n1275 GND 0.15fF
C1789 VDD.n1276 GND 0.01fF
C1790 VDD.n1277 GND 0.02fF
C1791 VDD.n1278 GND 0.03fF
C1792 VDD.n1279 GND 0.14fF
C1793 VDD.n1280 GND 0.16fF
C1794 VDD.n1281 GND 0.01fF
C1795 VDD.n1282 GND 0.11fF
C1796 VDD.n1283 GND 0.02fF
C1797 VDD.n1284 GND 0.02fF
C1798 VDD.n1285 GND 0.02fF
C1799 VDD.n1286 GND 0.14fF
C1800 VDD.n1287 GND 0.17fF
C1801 VDD.n1288 GND 0.01fF
C1802 VDD.n1289 GND 0.02fF
C1803 VDD.n1290 GND 0.02fF
C1804 VDD.n1291 GND 0.22fF
C1805 VDD.n1292 GND 0.01fF
C1806 VDD.n1293 GND 0.07fF
C1807 VDD.n1294 GND 0.02fF
C1808 VDD.n1295 GND 0.28fF
C1809 VDD.n1296 GND 0.01fF
C1810 VDD.n1297 GND 0.02fF
C1811 VDD.n1298 GND 0.02fF
C1812 VDD.n1299 GND 0.28fF
C1813 VDD.n1300 GND 0.01fF
C1814 VDD.n1301 GND 0.02fF
C1815 VDD.n1302 GND 0.03fF
C1816 VDD.n1303 GND 0.02fF
C1817 VDD.n1304 GND 0.02fF
C1818 VDD.n1305 GND 0.02fF
C1819 VDD.n1306 GND 0.31fF
C1820 VDD.n1307 GND 0.04fF
C1821 VDD.n1308 GND 0.03fF
C1822 VDD.n1309 GND 0.02fF
C1823 VDD.n1310 GND 0.02fF
C1824 VDD.n1311 GND 0.02fF
C1825 VDD.n1312 GND 0.03fF
C1826 VDD.n1313 GND 0.02fF
C1827 VDD.n1315 GND 0.02fF
C1828 VDD.n1316 GND 0.02fF
C1829 VDD.n1317 GND 0.02fF
C1830 VDD.n1319 GND 0.28fF
C1831 VDD.n1321 GND 0.02fF
C1832 VDD.n1322 GND 0.02fF
C1833 VDD.n1323 GND 0.03fF
C1834 VDD.n1324 GND 0.02fF
C1835 VDD.n1325 GND 0.28fF
C1836 VDD.n1326 GND 0.01fF
C1837 VDD.n1327 GND 0.02fF
C1838 VDD.n1328 GND 0.03fF
C1839 VDD.n1329 GND 0.28fF
C1840 VDD.n1330 GND 0.01fF
C1841 VDD.n1331 GND 0.02fF
C1842 VDD.n1332 GND 0.02fF
C1843 VDD.n1333 GND 0.06fF
C1844 VDD.n1334 GND 0.23fF
C1845 VDD.n1335 GND 0.01fF
C1846 VDD.n1336 GND 0.01fF
C1847 VDD.n1337 GND 0.02fF
C1848 VDD.n1338 GND 0.14fF
C1849 VDD.n1339 GND 0.17fF
C1850 VDD.n1340 GND 0.01fF
C1851 VDD.n1341 GND 0.02fF
C1852 VDD.n1342 GND 0.02fF
C1853 VDD.n1343 GND 0.11fF
C1854 VDD.n1344 GND 0.02fF
C1855 VDD.n1345 GND 0.14fF
C1856 VDD.n1346 GND 0.16fF
C1857 VDD.n1347 GND 0.01fF
C1858 VDD.n1348 GND 0.02fF
C1859 VDD.n1349 GND 0.02fF
C1860 VDD.n1350 GND 0.18fF
C1861 VDD.n1351 GND 0.15fF
C1862 VDD.n1352 GND 0.01fF
C1863 VDD.n1353 GND 0.02fF
C1864 VDD.n1354 GND 0.03fF
C1865 VDD.n1355 GND 0.18fF
C1866 VDD.n1356 GND 0.15fF
C1867 VDD.n1357 GND 0.01fF
C1868 VDD.n1358 GND 0.02fF
C1869 VDD.n1359 GND 0.03fF
C1870 VDD.n1360 GND 0.14fF
C1871 VDD.n1361 GND 0.16fF
C1872 VDD.n1362 GND 0.01fF
C1873 VDD.n1363 GND 0.11fF
C1874 VDD.n1364 GND 0.02fF
C1875 VDD.n1365 GND 0.02fF
C1876 VDD.n1366 GND 0.02fF
C1877 VDD.n1367 GND 0.14fF
C1878 VDD.n1368 GND 0.17fF
C1879 VDD.n1369 GND 0.01fF
C1880 VDD.n1370 GND 0.02fF
C1881 VDD.n1371 GND 0.02fF
C1882 VDD.n1372 GND 0.22fF
C1883 VDD.n1373 GND 0.01fF
C1884 VDD.n1374 GND 0.07fF
C1885 VDD.n1375 GND 0.02fF
C1886 VDD.n1376 GND 0.28fF
C1887 VDD.n1377 GND 0.01fF
C1888 VDD.n1378 GND 0.02fF
C1889 VDD.n1379 GND 0.02fF
C1890 VDD.n1380 GND 0.28fF
C1891 VDD.n1381 GND 0.01fF
C1892 VDD.n1382 GND 0.02fF
C1893 VDD.n1383 GND 0.03fF
C1894 VDD.n1384 GND 0.02fF
C1895 VDD.n1385 GND 0.02fF
C1896 VDD.n1386 GND 0.02fF
C1897 VDD.n1387 GND 0.26fF
C1898 VDD.n1388 GND 0.04fF
C1899 VDD.n1389 GND 0.03fF
C1900 VDD.n1390 GND 0.02fF
C1901 VDD.n1391 GND 0.02fF
C1902 VDD.n1392 GND 0.02fF
C1903 VDD.n1393 GND 0.03fF
C1904 VDD.n1394 GND 0.02fF
C1905 VDD.n1396 GND 0.02fF
C1906 VDD.n1397 GND 0.02fF
C1907 VDD.n1398 GND 0.02fF
C1908 VDD.n1400 GND 0.28fF
C1909 VDD.n1402 GND 0.02fF
C1910 VDD.n1403 GND 0.02fF
C1911 VDD.n1404 GND 0.03fF
C1912 VDD.n1405 GND 0.02fF
C1913 VDD.n1406 GND 0.28fF
C1914 VDD.n1407 GND 0.01fF
C1915 VDD.n1408 GND 0.02fF
C1916 VDD.n1409 GND 0.03fF
C1917 VDD.n1410 GND 0.06fF
C1918 VDD.n1411 GND 0.25fF
C1919 VDD.n1412 GND 0.01fF
C1920 VDD.n1413 GND 0.01fF
C1921 VDD.n1414 GND 0.02fF
C1922 VDD.n1415 GND 0.14fF
C1923 VDD.n1416 GND 0.16fF
C1924 VDD.n1417 GND 0.01fF
C1925 VDD.n1418 GND 0.02fF
C1926 VDD.n1419 GND 0.02fF
C1927 VDD.n1420 GND 0.17fF
C1928 VDD.n1421 GND 0.14fF
C1929 VDD.n1422 GND 0.01fF
C1930 VDD.n1423 GND 0.02fF
C1931 VDD.n1424 GND 0.03fF
C1932 VDD.n1425 GND 0.11fF
C1933 VDD.n1426 GND 0.03fF
C1934 VDD.n1427 GND 0.31fF
C1935 VDD.n1428 GND 0.01fF
C1936 VDD.n1429 GND 0.02fF
C1937 VDD.n1430 GND 0.03fF
C1938 VDD.n1431 GND 0.14fF
C1939 VDD.n1432 GND 0.17fF
C1940 VDD.n1433 GND 0.01fF
C1941 VDD.n1434 GND 0.02fF
C1942 VDD.n1435 GND 0.02fF
C1943 VDD.n1436 GND 0.06fF
C1944 VDD.n1437 GND 0.25fF
C1945 VDD.n1438 GND 0.01fF
C1946 VDD.n1439 GND 0.01fF
C1947 VDD.n1440 GND 0.02fF
C1948 VDD.n1441 GND 0.28fF
C1949 VDD.n1442 GND 0.01fF
C1950 VDD.n1443 GND 0.02fF
C1951 VDD.n1444 GND 0.03fF
C1952 VDD.n1445 GND 0.02fF
C1953 VDD.n1446 GND 0.02fF
C1954 VDD.n1447 GND 0.02fF
C1955 VDD.n1448 GND 0.26fF
C1956 VDD.n1449 GND 0.04fF
C1957 VDD.n1450 GND 0.03fF
C1958 VDD.n1451 GND 0.02fF
C1959 VDD.n1452 GND 0.02fF
C1960 VDD.n1453 GND 0.02fF
C1961 VDD.n1454 GND 0.03fF
C1962 VDD.n1455 GND 0.02fF
C1963 VDD.n1457 GND 0.02fF
C1964 VDD.n1458 GND 0.02fF
C1965 VDD.n1459 GND 0.02fF
C1966 VDD.n1461 GND 0.28fF
C1967 VDD.n1463 GND 0.02fF
C1968 VDD.n1464 GND 0.02fF
C1969 VDD.n1465 GND 0.03fF
C1970 VDD.n1466 GND 0.02fF
C1971 VDD.n1467 GND 0.28fF
C1972 VDD.n1468 GND 0.01fF
C1973 VDD.n1469 GND 0.02fF
C1974 VDD.n1470 GND 0.03fF
C1975 VDD.n1471 GND 0.28fF
C1976 VDD.n1472 GND 0.01fF
C1977 VDD.n1473 GND 0.02fF
C1978 VDD.n1474 GND 0.02fF
C1979 VDD.n1475 GND 0.06fF
C1980 VDD.n1476 GND 0.23fF
C1981 VDD.n1477 GND 0.01fF
C1982 VDD.n1478 GND 0.01fF
C1983 VDD.n1479 GND 0.02fF
C1984 VDD.n1480 GND 0.14fF
C1985 VDD.n1481 GND 0.17fF
C1986 VDD.n1482 GND 0.01fF
C1987 VDD.n1483 GND 0.02fF
C1988 VDD.n1484 GND 0.02fF
C1989 VDD.n1485 GND 0.11fF
C1990 VDD.n1486 GND 0.02fF
C1991 VDD.n1487 GND 0.14fF
C1992 VDD.n1488 GND 0.16fF
C1993 VDD.n1489 GND 0.01fF
C1994 VDD.n1490 GND 0.02fF
C1995 VDD.n1491 GND 0.02fF
C1996 VDD.n1492 GND 0.18fF
C1997 VDD.n1493 GND 0.15fF
C1998 VDD.n1494 GND 0.01fF
C1999 VDD.n1495 GND 0.02fF
C2000 VDD.n1496 GND 0.03fF
C2001 VDD.n1497 GND 0.18fF
C2002 VDD.n1498 GND 0.15fF
C2003 VDD.n1499 GND 0.01fF
C2004 VDD.n1500 GND 0.02fF
C2005 VDD.n1501 GND 0.03fF
C2006 VDD.n1502 GND 0.14fF
C2007 VDD.n1503 GND 0.16fF
C2008 VDD.n1504 GND 0.01fF
C2009 VDD.n1505 GND 0.11fF
C2010 VDD.n1506 GND 0.02fF
C2011 VDD.n1507 GND 0.02fF
C2012 VDD.n1508 GND 0.02fF
C2013 VDD.n1509 GND 0.14fF
C2014 VDD.n1510 GND 0.17fF
C2015 VDD.n1511 GND 0.01fF
C2016 VDD.n1512 GND 0.02fF
C2017 VDD.n1513 GND 0.02fF
C2018 VDD.n1514 GND 0.22fF
C2019 VDD.n1515 GND 0.01fF
C2020 VDD.n1516 GND 0.07fF
C2021 VDD.n1517 GND 0.02fF
C2022 VDD.n1518 GND 0.28fF
C2023 VDD.n1519 GND 0.01fF
C2024 VDD.n1520 GND 0.02fF
C2025 VDD.n1521 GND 0.02fF
C2026 VDD.n1522 GND 0.28fF
C2027 VDD.n1523 GND 0.01fF
C2028 VDD.n1524 GND 0.02fF
C2029 VDD.n1525 GND 0.03fF
C2030 RN.n0 GND 0.89fF
C2031 RN.t22 GND 0.81fF
C2032 RN.n1 GND 0.68fF
C2033 RN.n2 GND 0.86fF
C2034 RN.t11 GND 0.82fF
C2035 RN.n3 GND 0.66fF
C2036 RN.n4 GND 2.38fF
C2037 RN.n5 GND 0.86fF
C2038 RN.t20 GND 0.83fF
C2039 RN.n6 GND 0.66fF
C2040 RN.n7 GND 3.35fF
C2041 RN.n8 GND 0.89fF
C2042 RN.t4 GND 0.81fF
C2043 RN.n9 GND 0.66fF
C2044 RN.n10 GND 2.69fF
C2045 RN.n11 GND 0.86fF
C2046 RN.t26 GND 0.82fF
C2047 RN.n12 GND 0.66fF
C2048 RN.n13 GND 1.80fF
C2049 RN.n14 GND 0.86fF
C2050 RN.t2 GND 0.83fF
C2051 RN.n15 GND 0.66fF
C2052 RN.n16 GND 3.35fF
C2053 RN.n17 GND 0.89fF
C2054 RN.t18 GND 0.81fF
C2055 RN.n18 GND 0.66fF
C2056 RN.n19 GND 2.69fF
C2057 RN.n20 GND 0.86fF
C2058 RN.t7 GND 0.82fF
C2059 RN.n21 GND 0.66fF
C2060 RN.n22 GND 1.80fF
C2061 RN.n23 GND 0.86fF
C2062 RN.t16 GND 0.83fF
C2063 RN.n24 GND 0.66fF
C2064 RN.n25 GND 1.25fF
C2065 a_12396_101.n0 GND 0.02fF
C2066 a_12396_101.n1 GND 0.10fF
C2067 a_12396_101.n2 GND 0.07fF
C2068 a_12396_101.n3 GND 0.05fF
C2069 a_12396_101.n4 GND 0.00fF
C2070 a_12396_101.n5 GND 0.04fF
C2071 a_12396_101.n6 GND 0.05fF
C2072 a_12396_101.n7 GND 0.02fF
C2073 a_12396_101.n8 GND 0.05fF
C2074 a_12396_101.n9 GND 0.02fF
C2075 a_12396_101.n10 GND 0.08fF
C2076 a_12396_101.n11 GND 0.17fF
C2077 a_12396_101.t1 GND 0.23fF
C2078 a_12396_101.n12 GND 0.09fF
C2079 a_12396_101.n13 GND 0.00fF
C2080 a_10959_989.n0 GND 0.75fF
C2081 a_10959_989.n1 GND 0.75fF
C2082 a_10959_989.n2 GND 0.88fF
C2083 a_10959_989.n3 GND 0.28fF
C2084 a_10959_989.n4 GND 0.43fF
C2085 a_10959_989.n5 GND 0.53fF
C2086 a_10959_989.n6 GND 0.55fF
C2087 a_10959_989.n7 GND 0.53fF
C2088 a_10959_989.t12 GND 0.75fF
C2089 a_10959_989.n8 GND 0.55fF
C2090 a_10959_989.n9 GND 1.75fF
C2091 a_10959_989.n10 GND 0.64fF
C2092 a_10959_989.n11 GND 0.12fF
C2093 a_10959_989.n12 GND 0.41fF
C2094 a_10959_989.n13 GND 0.06fF
.ends
