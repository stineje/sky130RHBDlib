// File: bufx1.spi.pex
// Created: Tue Oct 15 15:55:38 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_BUFX1\%noxref_1 ( 9 21 25 47 51 62 65 76 88 89 )
c60 ( 89 0 ) capacitor c=0.0597349f //x=2.715 //y=0.37
c61 ( 88 0 ) capacitor c=0.0585876f //x=0.495 //y=0.37
c62 ( 76 0 ) capacitor c=0.0969492f //x=2.22 //y=0
c63 ( 65 0 ) capacitor c=0.192508f //x=0.63 //y=0
c64 ( 62 0 ) capacitor c=0.197741f //x=4.07 //y=0
c65 ( 60 0 ) capacitor c=0.0360484f //x=3.905 //y=0
c66 ( 54 0 ) capacitor c=0.00587411f //x=3.82 //y=0.45
c67 ( 51 0 ) capacitor c=0.00542558f //x=3.735 //y=0.535
c68 ( 50 0 ) capacitor c=0.00479856f //x=3.335 //y=0.45
c69 ( 47 0 ) capacitor c=0.00690112f //x=3.25 //y=0.535
c70 ( 42 0 ) capacitor c=0.00592191f //x=2.85 //y=0.45
c71 ( 39 0 ) capacitor c=0.0190475f //x=2.765 //y=0
c72 ( 34 0 ) capacitor c=0.0360484f //x=1.685 //y=0
c73 ( 33 0 ) capacitor c=0.0184787f //x=2.05 //y=0
c74 ( 28 0 ) capacitor c=0.00587411f //x=1.6 //y=0.45
c75 ( 25 0 ) capacitor c=0.00535892f //x=1.515 //y=0.535
c76 ( 24 0 ) capacitor c=0.00479856f //x=1.115 //y=0.45
c77 ( 21 0 ) capacitor c=0.00707849f //x=1.03 //y=0.535
c78 ( 16 0 ) capacitor c=0.00592191f //x=0.63 //y=0.45
c79 ( 9 0 ) capacitor c=0.190722f //x=4.07 //y=0
r80 (  80 81 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.335 //y=0 //x2=3.82 //y2=0
r81 (  79 80 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=3.33 //y=0 //x2=3.335 //y2=0
r82 (  77 79 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=2.85 //y=0 //x2=3.33 //y2=0
r83 (  68 69 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.115 //y=0 //x2=1.6 //y2=0
r84 (  67 68 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.115 //y2=0
r85 (  65 67 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=0.63 //y=0 //x2=0.74 //y2=0
r86 (  60 81 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.905 //y=0 //x2=3.82 //y2=0
r87 (  60 62 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=3.905 //y=0 //x2=4.07 //y2=0
r88 (  55 89 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.82 //y=0.62 //x2=3.82 //y2=0.535
r89 (  55 89 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=3.82 //y=0.62 //x2=3.82 //y2=1.225
r90 (  54 89 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.82 //y=0.45 //x2=3.82 //y2=0.535
r91 (  53 81 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.82 //y=0.17 //x2=3.82 //y2=0
r92 (  53 54 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=3.82 //y=0.17 //x2=3.82 //y2=0.45
r93 (  52 89 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.42 //y=0.535 //x2=3.335 //y2=0.535
r94 (  51 89 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.735 //y=0.535 //x2=3.82 //y2=0.535
r95 (  51 52 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.735 //y=0.535 //x2=3.42 //y2=0.535
r96 (  50 89 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.335 //y=0.45 //x2=3.335 //y2=0.535
r97 (  49 80 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.335 //y=0.17 //x2=3.335 //y2=0
r98 (  49 50 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=3.335 //y=0.17 //x2=3.335 //y2=0.45
r99 (  48 89 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=0.535 //x2=2.85 //y2=0.535
r100 (  47 89 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.25 //y=0.535 //x2=3.335 //y2=0.535
r101 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.25 //y=0.535 //x2=2.935 //y2=0.535
r102 (  43 89 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.62 //x2=2.85 //y2=0.535
r103 (  43 89 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.62 //x2=2.85 //y2=1.225
r104 (  42 89 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.45 //x2=2.85 //y2=0.535
r105 (  41 77 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.17 //x2=2.85 //y2=0
r106 (  41 42 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.17 //x2=2.85 //y2=0.45
r107 (  40 76 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.39 //y=0 //x2=2.22 //y2=0
r108 (  39 77 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=0 //x2=2.85 //y2=0
r109 (  39 40 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=2.765 //y=0 //x2=2.39 //y2=0
r110 (  34 69 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.6 //y2=0
r111 (  34 36 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.85 //y2=0
r112 (  33 76 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.05 //y=0 //x2=2.22 //y2=0
r113 (  33 36 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=1.85 //y2=0
r114 (  29 88 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=0.535
r115 (  29 88 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=1.225
r116 (  28 88 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.45 //x2=1.6 //y2=0.535
r117 (  27 69 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0
r118 (  27 28 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0.45
r119 (  26 88 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.2 //y=0.535 //x2=1.115 //y2=0.535
r120 (  25 88 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.6 //y2=0.535
r121 (  25 26 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.2 //y2=0.535
r122 (  24 88 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.45 //x2=1.115 //y2=0.535
r123 (  23 68 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0
r124 (  23 24 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0.45
r125 (  22 88 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.715 //y=0.535 //x2=0.63 //y2=0.535
r126 (  21 88 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=1.115 //y2=0.535
r127 (  21 22 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=0.715 //y2=0.535
r128 (  17 88 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=0.535
r129 (  17 88 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=1.225
r130 (  16 88 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.45 //x2=0.63 //y2=0.535
r131 (  15 65 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0
r132 (  15 16 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0.45
r133 (  9 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r134 (  7 79 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=0 //x2=3.33 //y2=0
r135 (  7 9 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=0 //x2=4.07 //y2=0
r136 (  5 36 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r137 (  5 7 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=3.33 //y2=0
r138 (  2 67 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r139 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_BUFX1\%noxref_1

subckt PM_BUFX1\%noxref_2 ( 9 21 43 56 60 62 65 66 67 68 )
c47 ( 68 0 ) capacitor c=0.0451925f //x=3.63 //y=5.02
c48 ( 67 0 ) capacitor c=0.0427416f //x=2.76 //y=5.02
c49 ( 66 0 ) capacitor c=0.0451925f //x=1.41 //y=5.02
c50 ( 65 0 ) capacitor c=0.0427416f //x=0.54 //y=5.02
c51 ( 64 0 ) capacitor c=0.00591168f //x=3.775 //y=7.4
c52 ( 63 0 ) capacitor c=0.00591168f //x=2.895 //y=7.4
c53 ( 62 0 ) capacitor c=0.109185f //x=2.22 //y=7.4
c54 ( 61 0 ) capacitor c=0.00591168f //x=1.555 //y=7.4
c55 ( 60 0 ) capacitor c=0.233263f //x=0.74 //y=7.4
c56 ( 56 0 ) capacitor c=0.228884f //x=4.07 //y=7.4
c57 ( 43 0 ) capacitor c=0.028745f //x=3.69 //y=7.4
c58 ( 35 0 ) capacitor c=0.0216067f //x=2.81 //y=7.4
c59 ( 29 0 ) capacitor c=0.0210379f //x=2.05 //y=7.4
c60 ( 21 0 ) capacitor c=0.028745f //x=1.47 //y=7.4
c61 ( 9 0 ) capacitor c=0.191847f //x=4.07 //y=7.4
r62 (  54 64 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.86 //y=7.4 //x2=3.775 //y2=7.4
r63 (  54 56 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=3.86 //y=7.4 //x2=4.07 //y2=7.4
r64 (  47 64 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.775 //y=7.23 //x2=3.775 //y2=7.4
r65 (  47 68 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=3.775 //y=7.23 //x2=3.775 //y2=6.405
r66 (  44 63 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.98 //y=7.4 //x2=2.895 //y2=7.4
r67 (  44 46 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li //thickness=0.1 \
 //x=2.98 //y=7.4 //x2=3.33 //y2=7.4
r68 (  43 64 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.69 //y=7.4 //x2=3.775 //y2=7.4
r69 (  43 46 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=3.69 //y=7.4 //x2=3.33 //y2=7.4
r70 (  37 63 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.895 //y=7.23 //x2=2.895 //y2=7.4
r71 (  37 67 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=2.895 //y=7.23 //x2=2.895 //y2=6.405
r72 (  36 62 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.39 //y=7.4 //x2=2.22 //y2=7.4
r73 (  35 63 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.81 //y=7.4 //x2=2.895 //y2=7.4
r74 (  35 36 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=2.81 //y=7.4 //x2=2.39 //y2=7.4
r75 (  30 61 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.555 //y2=7.4
r76 (  30 32 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.85 //y2=7.4
r77 (  29 62 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.05 //y=7.4 //x2=2.22 //y2=7.4
r78 (  29 32 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li //thickness=0.1 \
 //x=2.05 //y=7.4 //x2=1.85 //y2=7.4
r79 (  23 61 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.555 //y=7.23 //x2=1.555 //y2=7.4
r80 (  23 66 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=6.405
r81 (  22 60 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.76 //y=7.4 //x2=0.675 //y2=7.4
r82 (  21 61 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=1.555 //y2=7.4
r83 (  21 22 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=0.76 //y2=7.4
r84 (  15 60 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=0.675 //y=7.23 //x2=0.675 //y2=7.4
r85 (  15 65 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=6.405
r86 (  9 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=4.07 \
 //y=7.4 //x2=4.07 //y2=7.4
r87 (  7 46 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=3.33 \
 //y=7.4 //x2=3.33 //y2=7.4
r88 (  7 9 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=7.4 //x2=4.07 //y2=7.4
r89 (  5 32 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=1.85 \
 //y=7.4 //x2=1.85 //y2=7.4
r90 (  5 7 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=3.33 //y2=7.4
r91 (  2 60 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=7.4 //x2=0.74 //y2=7.4
r92 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_BUFX1\%noxref_2

subckt PM_BUFX1\%noxref_3 ( 1 2 17 18 19 20 24 26 33 34 35 36 37 38 39 43 44 \
 45 47 53 54 56 64 66 )
c102 ( 66 0 ) capacitor c=0.028734f //x=0.97 //y=5.02
c103 ( 64 0 ) capacitor c=0.0173218f //x=0.925 //y=0.91
c104 ( 56 0 ) capacitor c=0.0517753f //x=2.96 //y=2.085
c105 ( 54 0 ) capacitor c=0.0435629f //x=3.6 //y=1.255
c106 ( 53 0 ) capacitor c=0.0200386f //x=3.6 //y=0.91
c107 ( 47 0 ) capacitor c=0.0152946f //x=3.445 //y=1.41
c108 ( 45 0 ) capacitor c=0.0157804f //x=3.445 //y=0.755
c109 ( 44 0 ) capacitor c=0.0525175f //x=3.19 //y=4.79
c110 ( 43 0 ) capacitor c=0.0322983f //x=3.48 //y=4.79
c111 ( 39 0 ) capacitor c=0.0290017f //x=3.07 //y=1.92
c112 ( 38 0 ) capacitor c=0.0250027f //x=3.07 //y=1.565
c113 ( 37 0 ) capacitor c=0.0234316f //x=3.07 //y=1.255
c114 ( 36 0 ) capacitor c=0.0200596f //x=3.07 //y=0.91
c115 ( 35 0 ) capacitor c=0.154218f //x=3.555 //y=6.02
c116 ( 34 0 ) capacitor c=0.154243f //x=3.115 //y=6.02
c117 ( 26 0 ) capacitor c=0.0948753f //x=2.96 //y=2.085
c118 ( 24 0 ) capacitor c=0.0858431f //x=1.48 //y=2.59
c119 ( 20 0 ) capacitor c=0.00575887f //x=1.2 //y=4.58
c120 ( 19 0 ) capacitor c=0.0146153f //x=1.395 //y=4.58
c121 ( 18 0 ) capacitor c=0.00636159f //x=1.195 //y=2.08
c122 ( 17 0 ) capacitor c=0.0136204f //x=1.395 //y=2.08
c123 ( 2 0 ) capacitor c=0.0171827f //x=1.595 //y=2.59
c124 ( 1 0 ) capacitor c=0.0922367f //x=2.845 //y=2.59
r125 (  56 57 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.96 //y=2.085 //x2=3.07 //y2=2.085
r126 (  54 63 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.6 //y=1.255 //x2=3.56 //y2=1.41
r127 (  53 62 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.6 //y=0.91 //x2=3.56 //y2=0.755
r128 (  53 54 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.6 //y=0.91 //x2=3.6 //y2=1.255
r129 (  48 61 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.225 //y=1.41 //x2=3.11 //y2=1.41
r130 (  47 63 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.445 //y=1.41 //x2=3.56 //y2=1.41
r131 (  46 60 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.225 //y=0.755 //x2=3.11 //y2=0.755
r132 (  45 62 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.445 //y=0.755 //x2=3.56 //y2=0.755
r133 (  45 46 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.445 //y=0.755 //x2=3.225 //y2=0.755
r134 (  43 50 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=3.48 //y=4.79 //x2=3.555 //y2=4.865
r135 (  43 44 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=3.48 //y=4.79 //x2=3.19 //y2=4.79
r136 (  40 44 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=3.115 //y=4.865 //x2=3.19 //y2=4.79
r137 (  40 59 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=3.115 //y=4.865 //x2=2.96 //y2=4.7
r138 (  39 57 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.07 //y=1.92 //x2=3.07 //y2=2.085
r139 (  38 61 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.07 //y=1.565 //x2=3.11 //y2=1.41
r140 (  38 39 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=3.07 //y=1.565 //x2=3.07 //y2=1.92
r141 (  37 61 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.07 //y=1.255 //x2=3.11 //y2=1.41
r142 (  36 60 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.07 //y=0.91 //x2=3.11 //y2=0.755
r143 (  36 37 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.07 //y=0.91 //x2=3.07 //y2=1.255
r144 (  35 50 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.555 //y=6.02 //x2=3.555 //y2=4.865
r145 (  34 40 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.115 //y=6.02 //x2=3.115 //y2=4.865
r146 (  33 47 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.335 //y=1.41 //x2=3.445 //y2=1.41
r147 (  33 48 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.335 //y=1.41 //x2=3.225 //y2=1.41
r148 (  31 59 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.96 //y=4.7 //x2=2.96 //y2=4.7
r149 (  29 31 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=2.59 //x2=2.96 //y2=4.7
r150 (  26 56 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.96 //y=2.085 //x2=2.96 //y2=2.085
r151 (  26 29 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=2.96 //y=2.085 //x2=2.96 //y2=2.59
r152 (  22 24 ) resistor r=130.396 //w=0.187 //l=1.905 //layer=li \
 //thickness=0.1 //x=1.48 //y=4.495 //x2=1.48 //y2=2.59
r153 (  21 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.48 //y=2.165 //x2=1.48 //y2=2.59
r154 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.48 //y2=4.495
r155 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.2 //y2=4.58
r156 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.48 //y2=2.165
r157 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.195 //y2=2.08
r158 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.2 //y2=4.58
r159 (  11 66 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.115 //y2=5.725
r160 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.195 //y2=2.08
r161 (  7 64 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.11 //y2=1.005
r162 (  6 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.96 //y=2.59 //x2=2.96 //y2=2.59
r163 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.48 //y=2.59 //x2=1.48 //y2=2.59
r164 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.595 //y=2.59 //x2=1.48 //y2=2.59
r165 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.845 //y=2.59 //x2=2.96 //y2=2.59
r166 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=2.845 //y=2.59 //x2=1.595 //y2=2.59
ends PM_BUFX1\%noxref_3

subckt PM_BUFX1\%noxref_4 ( 2 7 8 9 10 11 12 13 17 18 19 21 27 28 30 )
c48 ( 30 0 ) capacitor c=0.0537799f //x=0.74 //y=2.085
c49 ( 28 0 ) capacitor c=0.0435629f //x=1.38 //y=1.255
c50 ( 27 0 ) capacitor c=0.0200386f //x=1.38 //y=0.91
c51 ( 21 0 ) capacitor c=0.0152946f //x=1.225 //y=1.41
c52 ( 19 0 ) capacitor c=0.0157804f //x=1.225 //y=0.755
c53 ( 18 0 ) capacitor c=0.0524167f //x=0.97 //y=4.79
c54 ( 17 0 ) capacitor c=0.0323991f //x=1.26 //y=4.79
c55 ( 13 0 ) capacitor c=0.0290017f //x=0.85 //y=1.92
c56 ( 12 0 ) capacitor c=0.0250027f //x=0.85 //y=1.565
c57 ( 11 0 ) capacitor c=0.0234316f //x=0.85 //y=1.255
c58 ( 10 0 ) capacitor c=0.0200596f //x=0.85 //y=0.91
c59 ( 9 0 ) capacitor c=0.154218f //x=1.335 //y=6.02
c60 ( 8 0 ) capacitor c=0.154243f //x=0.895 //y=6.02
c61 ( 2 0 ) capacitor c=0.114635f //x=0.74 //y=2.085
r62 (  30 31 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=0.74 //y=2.085 //x2=0.85 //y2=2.085
r63 (  28 37 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=1.255 //x2=1.34 //y2=1.41
r64 (  27 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.34 //y2=0.755
r65 (  27 28 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.38 //y2=1.255
r66 (  22 35 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=1.41 //x2=0.89 //y2=1.41
r67 (  21 37 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=1.41 //x2=1.34 //y2=1.41
r68 (  20 34 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=0.755 //x2=0.89 //y2=0.755
r69 (  19 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.34 //y2=0.755
r70 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.005 //y2=0.755
r71 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=1.335 //y2=4.865
r72 (  17 18 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=0.97 //y2=4.79
r73 (  14 18 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.97 //y2=4.79
r74 (  14 33 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.74 //y2=4.7
r75 (  13 31 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.92 //x2=0.85 //y2=2.085
r76 (  12 35 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.89 //y2=1.41
r77 (  12 13 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.85 //y2=1.92
r78 (  11 35 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.255 //x2=0.89 //y2=1.41
r79 (  10 34 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.89 //y2=0.755
r80 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.85 //y2=1.255
r81 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.335 //y=6.02 //x2=1.335 //y2=4.865
r82 (  8 14 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.895 //y=6.02 //x2=0.895 //y2=4.865
r83 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.225 //y2=1.41
r84 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.005 //y2=1.41
r85 (  5 33 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.7 //x2=0.74 //y2=4.7
r86 (  2 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=2.085
r87 (  2 5 ) resistor r=178.995 //w=0.187 //l=2.615 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=4.7
ends PM_BUFX1\%noxref_4

subckt PM_BUFX1\%noxref_5 ( 11 12 13 14 16 17 19 )
c43 ( 19 0 ) capacitor c=0.028734f //x=3.19 //y=5.02
c44 ( 17 0 ) capacitor c=0.0173218f //x=3.145 //y=0.91
c45 ( 16 0 ) capacitor c=0.105613f //x=3.7 //y=4.495
c46 ( 14 0 ) capacitor c=0.00575887f //x=3.42 //y=4.58
c47 ( 13 0 ) capacitor c=0.0146395f //x=3.615 //y=4.58
c48 ( 12 0 ) capacitor c=0.00636159f //x=3.415 //y=2.08
c49 ( 11 0 ) capacitor c=0.0141837f //x=3.615 //y=2.08
r50 (  15 16 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=3.7 //y=2.165 //x2=3.7 //y2=4.495
r51 (  13 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.615 //y=4.58 //x2=3.7 //y2=4.495
r52 (  13 14 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=3.615 //y=4.58 //x2=3.42 //y2=4.58
r53 (  11 15 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.615 //y=2.08 //x2=3.7 //y2=2.165
r54 (  11 12 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=3.615 //y=2.08 //x2=3.415 //y2=2.08
r55 (  5 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.335 //y=4.665 //x2=3.42 //y2=4.58
r56 (  5 19 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li //thickness=0.1 \
 //x=3.335 //y=4.665 //x2=3.335 //y2=5.725
r57 (  1 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.33 //y=1.995 //x2=3.415 //y2=2.08
r58 (  1 17 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=3.33 //y=1.995 //x2=3.33 //y2=1.005
ends PM_BUFX1\%noxref_5

