* SPICE3 file created from FILL1.ext - technology: sky130A

.subckt FILL1 VPWR VGND VPB VNB
.ends
