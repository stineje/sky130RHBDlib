* SPICE3 file created from DFFRNQX1.ext - technology: sky130A

.subckt DFFRNQX1 Q D CLK RN VDD VSS
X0 a_599_989 D VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.00124 ps=1.004 w=2 l=0.15 M=2
X1 VDD CLK a_277_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X2 VDD a_599_989 a_2141_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X3 VDD a_277_1050 a_3829_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X4 a_1334_210 D a_1053_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X5 Q a_147_187 a_4626_101 VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
X6 a_2141_1050 a_147_187 a_2036_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X7 a_599_989 RN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X8 a_147_187 CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X9 a_3829_1050 Q VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X10 Q a_3829_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.00116 pd=9.16 as=0 ps=0 w=2 l=0.15 M=2
X11 VDD a_599_989 a_277_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X12 VDD a_147_187 a_2141_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X13 VDD a_2141_1050 a_147_187 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X14 a_147_187 RN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X15 Q a_147_187 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X16 a_277_1050 a_599_989 a_372_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X17 a_147_187 RN a_2962_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X18 a_277_1050 a_147_187 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X19 VDD a_277_1050 a_599_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X20 VSS a_147_187 a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0.0010746 pd=9.42 as=0 ps=0 w=3 l=0.15
X21 a_3829_1050 Q a_3924_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X22 VDD RN a_3829_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X23 a_372_210 CLK a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X24 VSS a_277_1050 a_3643_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X25 VSS a_599_989 a_2036_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X26 VSS a_3829_1050 a_4626_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X27 a_599_989 RN a_1334_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X28 VSS a_2141_1050 a_2681_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X29 a_3924_210 RN a_3643_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X30 VSS a_277_1050 a_1053_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X31 a_2962_210 CLK a_2681_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 a_147_187 VDD 7.74f
C1 Q VDD 2.14f
C2 a_277_1050 a_599_989 2.02f
C3 a_277_1050 a_147_187 3.69f
C4 a_3829_1050 VDD 2.82f
C5 a_2141_1050 VDD 2.17f
C6 a_147_187 CLK 3.44f
C7 a_599_989 VDD 3.11f
C8 a_277_1050 VDD 3.23f
C9 VDD VSS 8.51f
.ends
