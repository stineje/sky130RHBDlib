magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 29 -17 63 21
<< locali >>
rect 35 325 69 493
rect 430 325 627 333
rect 35 299 627 325
rect 35 291 460 299
rect 17 215 87 257
rect 123 215 211 257
rect 245 215 339 257
rect 34 147 247 181
rect 34 51 69 147
rect 213 101 247 147
rect 283 135 339 215
rect 389 215 455 257
rect 389 135 440 215
rect 494 199 551 265
rect 585 165 627 299
rect 476 131 627 165
rect 476 101 516 131
rect 213 51 516 101
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 103 459 337 493
rect 103 359 153 459
rect 271 451 337 459
rect 375 443 441 527
rect 203 409 248 425
rect 475 409 525 493
rect 203 367 525 409
rect 559 375 625 527
rect 203 359 405 367
rect 103 17 169 113
rect 550 17 616 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 389 135 440 215 6 A1
port 1 nsew signal input
rlabel locali s 389 215 455 257 6 A1
port 1 nsew signal input
rlabel locali s 494 199 551 265 6 A2
port 2 nsew signal input
rlabel locali s 283 135 339 215 6 B1
port 3 nsew signal input
rlabel locali s 245 215 339 257 6 B1
port 3 nsew signal input
rlabel locali s 123 215 211 257 6 B2
port 4 nsew signal input
rlabel locali s 17 215 87 257 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 643 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 213 51 516 101 6 Y
port 10 nsew signal output
rlabel locali s 476 101 516 131 6 Y
port 10 nsew signal output
rlabel locali s 476 131 627 165 6 Y
port 10 nsew signal output
rlabel locali s 213 101 247 147 6 Y
port 10 nsew signal output
rlabel locali s 34 51 69 147 6 Y
port 10 nsew signal output
rlabel locali s 585 165 627 299 6 Y
port 10 nsew signal output
rlabel locali s 34 147 247 181 6 Y
port 10 nsew signal output
rlabel locali s 35 291 460 299 6 Y
port 10 nsew signal output
rlabel locali s 35 299 627 325 6 Y
port 10 nsew signal output
rlabel locali s 430 325 627 333 6 Y
port 10 nsew signal output
rlabel locali s 35 325 69 493 6 Y
port 10 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3657942
string GDS_START 3651372
<< end >>
