* SPICE3 file created from TMRDFFSNRNQNX1.ext - technology: sky130A

.subckt TMRDFFSNRNQNX1 SN RN D CLK Q VPB VNB
M1000 a_4447_943.t5 SN VPB.t37 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VPB.t55 CLK a_6371_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_7333_943.t5 RN VPB.t86 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t91 D a_6049_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VNB a_6049_1004.t8 a_6825_75.t0 nshort w=-1.605u l=1.765u
+  ad=3.7611p pd=32.97u as=0p ps=0u
M1005 a_7973_1004.t1 SN VPB.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_18197_1005.t6 a_9897_1004.t7 Q.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t105 a_4125_1004.t7 a_17533_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VNB a_4125_1004.t11 a_4901_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPB.t95 D a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t90 D a_11821_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VNB a_4125_1004.t15 a_17428_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t78 RN a_15669_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_599_943.t2 CLK VPB.t59 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPB.t85 RN a_9897_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPB.t63 CLK a_1561_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_11821_1004.t6 a_12143_943.t8 VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t34 a_13105_943.t7 a_13745_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_15669_1004.t7 a_18094_73.t0 nshort w=-1.235u l=1.535u
+  ad=0.5373p pd=4.72u as=0p ps=0u
M1019 VNB D a_11635_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPB.t13 a_277_1004.t7 a_2201_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_7333_943.t3 CLK VPB.t58 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_10219_943.t1 SN VPB.t41 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPB.t104 a_7333_943.t7 a_6371_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPB.t61 CLK a_12143_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_13105_943.t6 RN VPB.t82 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VNB a_6049_1004.t10 a_7787_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1027 VNB a_6371_943.t10 a_9711_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1028 VNB D a_5863_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB.t80 RN a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_6371_943.t3 a_6049_1004.t7 VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPB.t51 a_7973_1004.t7 a_7333_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPB.t50 a_9897_1004.t8 a_10219_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_17533_1005.t1 a_4125_1004.t8 VPB.t68 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_12143_943.t3 CLK VPB.t57 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_599_943.t6 a_1561_943.t8 VPB.t109 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_15991_943.t3 a_15669_1004.t9 VPB.t99 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPB.t83 RN a_1561_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_9897_1004.t4 a_6371_943.t7 VPB.t100 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VNB a_11821_1004.t9 a_12597_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_4125_1004.t0 a_599_943.t7 VPB.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPB.t38 SN a_2201_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VNB a_13745_1004.t9 a_14521_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_4125_1004.t3 a_4447_943.t8 VPB.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 VNB a_9897_1004.t14 a_10673_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPB.t8 a_6371_943.t8 a_6049_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_18197_1005.t3 a_4125_1004.t9 a_17533_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_1561_943.t2 CLK VPB.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 VNB a_7973_1004.t9 a_8749_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPB.t21 a_599_943.t8 a_277_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 VNB D a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_13745_1004.t1 SN VPB.t46 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 a_17533_1005.t6 a_9897_1004.t9 VPB.t98 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_12143_943.t6 a_11821_1004.t7 VPB.t106 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 VPB.t33 a_13745_1004.t7 a_13105_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_15991_943.t1 SN VPB.t47 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_15669_1004.t5 a_12143_943.t10 VPB.t64 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_4125_1004.t6 RN VPB.t79 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 VNB a_11821_1004.t12 a_13559_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1059 VPB.t102 a_1561_943.t11 a_2201_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 VPB.t76 RN a_6049_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 a_7333_943.t0 a_7973_1004.t8 VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_7973_1004.t5 a_7333_943.t10 VPB.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_9897_1004.t1 a_10219_943.t8 VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 VPB.t5 a_13105_943.t8 a_15991_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 VNB a_12143_943.t7 a_15483_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_1561_943.t1 a_2201_1004.t8 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_18197_1005.t7 a_15669_1004.t10 a_17533_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 VPB.t30 a_4125_1004.t10 a_4447_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_6371_943.t4 CLK VPB.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 VPB.t52 CLK a_7333_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_6049_1004.t5 D VPB.t92 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 Q a_9897_1004.t10 a_17428_73.t1 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1073 Q.t2 a_9897_1004.t11 a_18197_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 a_277_1004.t5 D VPB.t93 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 VPB.t53 CLK a_13105_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 a_15991_943.t5 a_13105_943.t10 VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 VNB a_15669_1004.t8 a_16445_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1078 VPB.t70 a_11821_1004.t8 a_13745_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 a_10219_943.t6 a_7333_943.t12 VPB.t32 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_15669_1004.t0 RN VPB.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 VPB.t10 a_13105_943.t11 a_12143_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 VPB.t29 a_277_1004.t10 a_599_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_9897_1004.t5 RN VPB.t87 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 VPB.t89 RN a_11821_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 VPB.t108 a_1561_943.t12 a_599_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_13745_1004.t4 a_13105_943.t12 VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 VPB.t42 SN a_4447_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_18197_1005.t2 a_15669_1004.t11 Q.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 VPB.t96 a_15991_943.t7 a_15669_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 a_6371_943.t0 a_7333_943.t13 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 VPB.t72 RN a_7333_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 VPB.t44 SN a_7973_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_277_1004.t3 RN VPB.t88 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_11821_1004.t0 RN VPB.t74 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 VNB a_277_1004.t8 a_2015_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1096 VPB.t43 SN a_13745_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_10219_943.t2 a_9897_1004.t12 VPB.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 VPB.t60 CLK a_599_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 VPB.t103 a_12143_943.t11 a_11821_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_1561_943.t5 RN VPB.t81 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 VPB.t101 a_1561_943.t13 a_4447_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_2201_1004.t0 SN VPB.t39 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 VPB.t77 RN a_4125_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_12143_943.t2 a_13105_943.t14 VPB.t36 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 VPB.t19 a_6049_1004.t9 a_7973_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VPB.t73 RN a_13105_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 a_599_943.t3 a_277_1004.t11 VPB.t110 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 a_277_1004.t2 a_599_943.t10 VPB.t26 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 a_11821_1004.t2 D VPB.t94 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 VNB a_2201_1004.t7 a_2977_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1111 VNB a_15669_1004.t12 a_18760_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1112 VNB a_4125_1004.t12 a_18094_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1113 a_13105_943.t1 a_13745_1004.t8 VPB.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1114 VPB.t4 a_15669_1004.t13 a_15991_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 VNB a_277_1004.t9 a_1053_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1116 a_7973_1004.t2 a_6049_1004.t11 VPB.t67 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1117 VPB.t0 a_6371_943.t11 a_9897_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_2201_1004.t2 a_277_1004.t12 VPB.t97 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 VPB.t23 a_7333_943.t14 a_10219_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 a_2201_1004.t5 a_1561_943.t14 VPB.t107 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 VPB.t49 a_599_943.t12 a_4125_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 VPB.t15 a_4447_943.t9 a_4125_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 a_6049_1004.t3 RN VPB.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1124 a_17533_1005.t3 a_4125_1004.t13 a_18197_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1125 a_4447_943.t1 a_4125_1004.t14 VPB.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1126 VPB.t16 a_6049_1004.t12 a_6371_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1127 a_4447_943.t2 a_1561_943.t15 VPB.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1128 Q a_9897_1004.t13 a_18760_73.t0 nshort w=-1.83u l=2.06u
+  ad=0p pd=0u as=0p ps=0u
M1129 VNB a_599_943.t9 a_3939_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1130 a_15669_1004.t6 a_15991_943.t9 VPB.t111 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1131 VPB.t69 a_11821_1004.t10 a_12143_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1132 VPB.t18 a_9897_1004.t15 a_17533_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1133 a_13105_943.t2 CLK VPB.t54 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1134 VPB.t48 SN a_15991_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1135 VPB.t40 SN a_10219_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1136 a_13745_1004.t2 a_11821_1004.t11 VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1137 VPB.t22 a_12143_943.t12 a_15669_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1138 a_6049_1004.t1 a_6371_943.t12 VPB.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1139 VPB.t65 a_7333_943.t15 a_7973_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1140 VPB.t6 a_10219_943.t9 a_9897_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1141 VPB.t11 a_2201_1004.t9 a_1561_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1142 Q.t1 a_15669_1004.t14 a_18197_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1143 a_17533_1005.t0 a_15669_1004.t15 a_18197_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u











R0 VPB VPB.n1682 126.832
R1 VPB.n40 VPB.n38 94.117
R2 VPB.n1604 VPB.n1602 94.117
R3 VPB.n1521 VPB.n1519 94.117
R4 VPB.n1438 VPB.n1436 94.117
R5 VPB.n1355 VPB.n1353 94.117
R6 VPB.n1272 VPB.n1270 94.117
R7 VPB.n1189 VPB.n1187 94.117
R8 VPB.n1106 VPB.n1104 94.117
R9 VPB.n1023 VPB.n1021 94.117
R10 VPB.n940 VPB.n938 94.117
R11 VPB.n129 VPB.n127 94.117
R12 VPB.n863 VPB.n861 94.117
R13 VPB.n780 VPB.n778 94.117
R14 VPB.n697 VPB.n695 94.117
R15 VPB.n614 VPB.n612 94.117
R16 VPB.n531 VPB.n529 94.117
R17 VPB.n448 VPB.n446 94.117
R18 VPB.n365 VPB.n363 94.117
R19 VPB.n302 VPB.n300 94.117
R20 VPB.n247 VPB.n245 94.117
R21 VPB.n378 VPB.n377 80.104
R22 VPB.n461 VPB.n460 80.104
R23 VPB.n544 VPB.n543 80.104
R24 VPB.n627 VPB.n626 80.104
R25 VPB.n710 VPB.n709 80.104
R26 VPB.n793 VPB.n792 80.104
R27 VPB.n876 VPB.n875 80.104
R28 VPB.n139 VPB.n138 80.104
R29 VPB.n953 VPB.n952 80.104
R30 VPB.n1036 VPB.n1035 80.104
R31 VPB.n1119 VPB.n1118 80.104
R32 VPB.n1202 VPB.n1201 80.104
R33 VPB.n1285 VPB.n1284 80.104
R34 VPB.n1368 VPB.n1367 80.104
R35 VPB.n1451 VPB.n1450 80.104
R36 VPB.n1534 VPB.n1533 80.104
R37 VPB.n1617 VPB.n1616 80.104
R38 VPB.n50 VPB.n49 80.104
R39 VPB.n210 VPB.n209 76
R40 VPB.n214 VPB.n213 76
R41 VPB.n218 VPB.n217 76
R42 VPB.n222 VPB.n221 76
R43 VPB.n249 VPB.n248 76
R44 VPB.n253 VPB.n252 76
R45 VPB.n257 VPB.n256 76
R46 VPB.n261 VPB.n260 76
R47 VPB.n265 VPB.n264 76
R48 VPB.n269 VPB.n268 76
R49 VPB.n273 VPB.n272 76
R50 VPB.n277 VPB.n276 76
R51 VPB.n304 VPB.n303 76
R52 VPB.n309 VPB.n308 76
R53 VPB.n314 VPB.n313 76
R54 VPB.n321 VPB.n320 76
R55 VPB.n326 VPB.n325 76
R56 VPB.n331 VPB.n330 76
R57 VPB.n336 VPB.n335 76
R58 VPB.n340 VPB.n339 76
R59 VPB.n367 VPB.n366 76
R60 VPB.n371 VPB.n370 76
R61 VPB.n376 VPB.n375 76
R62 VPB.n381 VPB.n380 76
R63 VPB.n388 VPB.n387 76
R64 VPB.n393 VPB.n392 76
R65 VPB.n398 VPB.n397 76
R66 VPB.n405 VPB.n404 76
R67 VPB.n410 VPB.n409 76
R68 VPB.n415 VPB.n414 76
R69 VPB.n419 VPB.n418 76
R70 VPB.n423 VPB.n422 76
R71 VPB.n450 VPB.n449 76
R72 VPB.n454 VPB.n453 76
R73 VPB.n459 VPB.n458 76
R74 VPB.n464 VPB.n463 76
R75 VPB.n471 VPB.n470 76
R76 VPB.n476 VPB.n475 76
R77 VPB.n481 VPB.n480 76
R78 VPB.n488 VPB.n487 76
R79 VPB.n493 VPB.n492 76
R80 VPB.n498 VPB.n497 76
R81 VPB.n502 VPB.n501 76
R82 VPB.n506 VPB.n505 76
R83 VPB.n533 VPB.n532 76
R84 VPB.n537 VPB.n536 76
R85 VPB.n542 VPB.n541 76
R86 VPB.n547 VPB.n546 76
R87 VPB.n554 VPB.n553 76
R88 VPB.n559 VPB.n558 76
R89 VPB.n564 VPB.n563 76
R90 VPB.n571 VPB.n570 76
R91 VPB.n576 VPB.n575 76
R92 VPB.n581 VPB.n580 76
R93 VPB.n585 VPB.n584 76
R94 VPB.n589 VPB.n588 76
R95 VPB.n616 VPB.n615 76
R96 VPB.n620 VPB.n619 76
R97 VPB.n625 VPB.n624 76
R98 VPB.n630 VPB.n629 76
R99 VPB.n637 VPB.n636 76
R100 VPB.n642 VPB.n641 76
R101 VPB.n647 VPB.n646 76
R102 VPB.n654 VPB.n653 76
R103 VPB.n659 VPB.n658 76
R104 VPB.n664 VPB.n663 76
R105 VPB.n668 VPB.n667 76
R106 VPB.n672 VPB.n671 76
R107 VPB.n699 VPB.n698 76
R108 VPB.n703 VPB.n702 76
R109 VPB.n708 VPB.n707 76
R110 VPB.n713 VPB.n712 76
R111 VPB.n720 VPB.n719 76
R112 VPB.n725 VPB.n724 76
R113 VPB.n730 VPB.n729 76
R114 VPB.n737 VPB.n736 76
R115 VPB.n742 VPB.n741 76
R116 VPB.n747 VPB.n746 76
R117 VPB.n751 VPB.n750 76
R118 VPB.n755 VPB.n754 76
R119 VPB.n782 VPB.n781 76
R120 VPB.n786 VPB.n785 76
R121 VPB.n791 VPB.n790 76
R122 VPB.n796 VPB.n795 76
R123 VPB.n803 VPB.n802 76
R124 VPB.n808 VPB.n807 76
R125 VPB.n813 VPB.n812 76
R126 VPB.n820 VPB.n819 76
R127 VPB.n825 VPB.n824 76
R128 VPB.n830 VPB.n829 76
R129 VPB.n834 VPB.n833 76
R130 VPB.n838 VPB.n837 76
R131 VPB.n865 VPB.n864 76
R132 VPB.n869 VPB.n868 76
R133 VPB.n874 VPB.n873 76
R134 VPB.n879 VPB.n878 76
R135 VPB.n886 VPB.n885 76
R136 VPB.n891 VPB.n890 76
R137 VPB.n896 VPB.n895 76
R138 VPB.n903 VPB.n902 76
R139 VPB.n908 VPB.n907 76
R140 VPB.n913 VPB.n912 76
R141 VPB.n917 VPB.n916 76
R142 VPB.n921 VPB.n920 76
R143 VPB.n936 VPB.n933 76
R144 VPB.n942 VPB.n941 76
R145 VPB.n946 VPB.n945 76
R146 VPB.n951 VPB.n950 76
R147 VPB.n956 VPB.n955 76
R148 VPB.n963 VPB.n962 76
R149 VPB.n968 VPB.n967 76
R150 VPB.n973 VPB.n972 76
R151 VPB.n980 VPB.n979 76
R152 VPB.n985 VPB.n984 76
R153 VPB.n990 VPB.n989 76
R154 VPB.n994 VPB.n993 76
R155 VPB.n998 VPB.n997 76
R156 VPB.n1025 VPB.n1024 76
R157 VPB.n1029 VPB.n1028 76
R158 VPB.n1034 VPB.n1033 76
R159 VPB.n1039 VPB.n1038 76
R160 VPB.n1046 VPB.n1045 76
R161 VPB.n1051 VPB.n1050 76
R162 VPB.n1056 VPB.n1055 76
R163 VPB.n1063 VPB.n1062 76
R164 VPB.n1068 VPB.n1067 76
R165 VPB.n1073 VPB.n1072 76
R166 VPB.n1077 VPB.n1076 76
R167 VPB.n1081 VPB.n1080 76
R168 VPB.n1108 VPB.n1107 76
R169 VPB.n1112 VPB.n1111 76
R170 VPB.n1117 VPB.n1116 76
R171 VPB.n1122 VPB.n1121 76
R172 VPB.n1129 VPB.n1128 76
R173 VPB.n1134 VPB.n1133 76
R174 VPB.n1139 VPB.n1138 76
R175 VPB.n1146 VPB.n1145 76
R176 VPB.n1151 VPB.n1150 76
R177 VPB.n1156 VPB.n1155 76
R178 VPB.n1160 VPB.n1159 76
R179 VPB.n1164 VPB.n1163 76
R180 VPB.n1191 VPB.n1190 76
R181 VPB.n1195 VPB.n1194 76
R182 VPB.n1200 VPB.n1199 76
R183 VPB.n1205 VPB.n1204 76
R184 VPB.n1212 VPB.n1211 76
R185 VPB.n1217 VPB.n1216 76
R186 VPB.n1222 VPB.n1221 76
R187 VPB.n1229 VPB.n1228 76
R188 VPB.n1234 VPB.n1233 76
R189 VPB.n1239 VPB.n1238 76
R190 VPB.n1243 VPB.n1242 76
R191 VPB.n1247 VPB.n1246 76
R192 VPB.n1274 VPB.n1273 76
R193 VPB.n1278 VPB.n1277 76
R194 VPB.n1283 VPB.n1282 76
R195 VPB.n1288 VPB.n1287 76
R196 VPB.n1295 VPB.n1294 76
R197 VPB.n1300 VPB.n1299 76
R198 VPB.n1305 VPB.n1304 76
R199 VPB.n1312 VPB.n1311 76
R200 VPB.n1317 VPB.n1316 76
R201 VPB.n1322 VPB.n1321 76
R202 VPB.n1326 VPB.n1325 76
R203 VPB.n1330 VPB.n1329 76
R204 VPB.n1357 VPB.n1356 76
R205 VPB.n1361 VPB.n1360 76
R206 VPB.n1366 VPB.n1365 76
R207 VPB.n1371 VPB.n1370 76
R208 VPB.n1378 VPB.n1377 76
R209 VPB.n1383 VPB.n1382 76
R210 VPB.n1388 VPB.n1387 76
R211 VPB.n1395 VPB.n1394 76
R212 VPB.n1400 VPB.n1399 76
R213 VPB.n1405 VPB.n1404 76
R214 VPB.n1409 VPB.n1408 76
R215 VPB.n1413 VPB.n1412 76
R216 VPB.n1440 VPB.n1439 76
R217 VPB.n1444 VPB.n1443 76
R218 VPB.n1449 VPB.n1448 76
R219 VPB.n1454 VPB.n1453 76
R220 VPB.n1461 VPB.n1460 76
R221 VPB.n1466 VPB.n1465 76
R222 VPB.n1471 VPB.n1470 76
R223 VPB.n1478 VPB.n1477 76
R224 VPB.n1483 VPB.n1482 76
R225 VPB.n1488 VPB.n1487 76
R226 VPB.n1492 VPB.n1491 76
R227 VPB.n1496 VPB.n1495 76
R228 VPB.n1523 VPB.n1522 76
R229 VPB.n1527 VPB.n1526 76
R230 VPB.n1532 VPB.n1531 76
R231 VPB.n1537 VPB.n1536 76
R232 VPB.n1544 VPB.n1543 76
R233 VPB.n1549 VPB.n1548 76
R234 VPB.n1554 VPB.n1553 76
R235 VPB.n1561 VPB.n1560 76
R236 VPB.n1566 VPB.n1565 76
R237 VPB.n1571 VPB.n1570 76
R238 VPB.n1575 VPB.n1574 76
R239 VPB.n1579 VPB.n1578 76
R240 VPB.n1606 VPB.n1605 76
R241 VPB.n1610 VPB.n1609 76
R242 VPB.n1615 VPB.n1614 76
R243 VPB.n1620 VPB.n1619 76
R244 VPB.n1627 VPB.n1626 76
R245 VPB.n1632 VPB.n1631 76
R246 VPB.n1637 VPB.n1636 76
R247 VPB.n1644 VPB.n1643 76
R248 VPB.n1649 VPB.n1648 76
R249 VPB.n1654 VPB.n1653 76
R250 VPB.n1658 VPB.n1657 76
R251 VPB.n1662 VPB.n1661 76
R252 VPB.n1675 VPB.n1674 76
R253 VPB.n407 VPB.n406 75.654
R254 VPB.n490 VPB.n489 75.654
R255 VPB.n573 VPB.n572 75.654
R256 VPB.n656 VPB.n655 75.654
R257 VPB.n739 VPB.n738 75.654
R258 VPB.n822 VPB.n821 75.654
R259 VPB.n905 VPB.n904 75.654
R260 VPB.n161 VPB.n160 75.654
R261 VPB.n982 VPB.n981 75.654
R262 VPB.n1065 VPB.n1064 75.654
R263 VPB.n1148 VPB.n1147 75.654
R264 VPB.n1231 VPB.n1230 75.654
R265 VPB.n1314 VPB.n1313 75.654
R266 VPB.n1397 VPB.n1396 75.654
R267 VPB.n1480 VPB.n1479 75.654
R268 VPB.n1563 VPB.n1562 75.654
R269 VPB.n1646 VPB.n1645 75.654
R270 VPB.n72 VPB.n71 75.654
R271 VPB.n22 VPB.n21 61.764
R272 VPB.n1586 VPB.n1585 61.764
R273 VPB.n1503 VPB.n1502 61.764
R274 VPB.n1420 VPB.n1419 61.764
R275 VPB.n1337 VPB.n1336 61.764
R276 VPB.n1254 VPB.n1253 61.764
R277 VPB.n1171 VPB.n1170 61.764
R278 VPB.n1088 VPB.n1087 61.764
R279 VPB.n1005 VPB.n1004 61.764
R280 VPB.n88 VPB.n87 61.764
R281 VPB.n111 VPB.n110 61.764
R282 VPB.n845 VPB.n844 61.764
R283 VPB.n762 VPB.n761 61.764
R284 VPB.n679 VPB.n678 61.764
R285 VPB.n596 VPB.n595 61.764
R286 VPB.n513 VPB.n512 61.764
R287 VPB.n430 VPB.n429 61.764
R288 VPB.n347 VPB.n346 61.764
R289 VPB.n284 VPB.n283 61.764
R290 VPB.n229 VPB.n228 61.764
R291 VPB.n332 VPB.t68 55.465
R292 VPB.n305 VPB.t18 55.465
R293 VPB.n78 VPB.t93 55.106
R294 VPB.n1650 VPB.t110 55.106
R295 VPB.n1567 VPB.t97 55.106
R296 VPB.n1484 VPB.t12 55.106
R297 VPB.n1401 VPB.t27 55.106
R298 VPB.n1318 VPB.t24 55.106
R299 VPB.n1235 VPB.t92 55.106
R300 VPB.n1152 VPB.t17 55.106
R301 VPB.n1069 VPB.t67 55.106
R302 VPB.n986 VPB.t14 55.106
R303 VPB.n167 VPB.t100 55.106
R304 VPB.n909 VPB.t28 55.106
R305 VPB.n826 VPB.t94 55.106
R306 VPB.n743 VPB.t106 55.106
R307 VPB.n660 VPB.t3 55.106
R308 VPB.n577 VPB.t35 55.106
R309 VPB.n494 VPB.t64 55.106
R310 VPB.n411 VPB.t99 55.106
R311 VPB.n45 VPB.t21 55.106
R312 VPB.n1611 VPB.t108 55.106
R313 VPB.n1528 VPB.t102 55.106
R314 VPB.n1445 VPB.t83 55.106
R315 VPB.n1362 VPB.t15 55.106
R316 VPB.n1279 VPB.t101 55.106
R317 VPB.n1196 VPB.t8 55.106
R318 VPB.n1113 VPB.t104 55.106
R319 VPB.n1030 VPB.t65 55.106
R320 VPB.n947 VPB.t72 55.106
R321 VPB.n134 VPB.t6 55.106
R322 VPB.n870 VPB.t23 55.106
R323 VPB.n787 VPB.t103 55.106
R324 VPB.n704 VPB.t10 55.106
R325 VPB.n621 VPB.t34 55.106
R326 VPB.n538 VPB.t73 55.106
R327 VPB.n455 VPB.t96 55.106
R328 VPB.n372 VPB.t5 55.106
R329 VPB.n311 VPB.n310 48.952
R330 VPB.n385 VPB.n384 48.952
R331 VPB.n468 VPB.n467 48.952
R332 VPB.n551 VPB.n550 48.952
R333 VPB.n634 VPB.n633 48.952
R334 VPB.n717 VPB.n716 48.952
R335 VPB.n800 VPB.n799 48.952
R336 VPB.n883 VPB.n882 48.952
R337 VPB.n143 VPB.n142 48.952
R338 VPB.n960 VPB.n959 48.952
R339 VPB.n1043 VPB.n1042 48.952
R340 VPB.n1126 VPB.n1125 48.952
R341 VPB.n1209 VPB.n1208 48.952
R342 VPB.n1292 VPB.n1291 48.952
R343 VPB.n1375 VPB.n1374 48.952
R344 VPB.n1458 VPB.n1457 48.952
R345 VPB.n1541 VPB.n1540 48.952
R346 VPB.n1624 VPB.n1623 48.952
R347 VPB.n54 VPB.n53 48.952
R348 VPB.n328 VPB.n327 44.502
R349 VPB.n402 VPB.n401 44.502
R350 VPB.n485 VPB.n484 44.502
R351 VPB.n568 VPB.n567 44.502
R352 VPB.n651 VPB.n650 44.502
R353 VPB.n734 VPB.n733 44.502
R354 VPB.n817 VPB.n816 44.502
R355 VPB.n900 VPB.n899 44.502
R356 VPB.n157 VPB.n156 44.502
R357 VPB.n977 VPB.n976 44.502
R358 VPB.n1060 VPB.n1059 44.502
R359 VPB.n1143 VPB.n1142 44.502
R360 VPB.n1226 VPB.n1225 44.502
R361 VPB.n1309 VPB.n1308 44.502
R362 VPB.n1392 VPB.n1391 44.502
R363 VPB.n1475 VPB.n1474 44.502
R364 VPB.n1558 VPB.n1557 44.502
R365 VPB.n1641 VPB.n1640 44.502
R366 VPB.n68 VPB.n67 44.502
R367 VPB.n316 VPB.n315 41.183
R368 VPB.n66 VPB.n14 40.824
R369 VPB.n57 VPB.n15 40.824
R370 VPB.n1639 VPB.n1638 40.824
R371 VPB.n1622 VPB.n1621 40.824
R372 VPB.n1556 VPB.n1555 40.824
R373 VPB.n1539 VPB.n1538 40.824
R374 VPB.n1473 VPB.n1472 40.824
R375 VPB.n1456 VPB.n1455 40.824
R376 VPB.n1390 VPB.n1389 40.824
R377 VPB.n1373 VPB.n1372 40.824
R378 VPB.n1307 VPB.n1306 40.824
R379 VPB.n1290 VPB.n1289 40.824
R380 VPB.n1224 VPB.n1223 40.824
R381 VPB.n1207 VPB.n1206 40.824
R382 VPB.n1141 VPB.n1140 40.824
R383 VPB.n1124 VPB.n1123 40.824
R384 VPB.n1058 VPB.n1057 40.824
R385 VPB.n1041 VPB.n1040 40.824
R386 VPB.n975 VPB.n974 40.824
R387 VPB.n958 VPB.n957 40.824
R388 VPB.n155 VPB.n103 40.824
R389 VPB.n146 VPB.n104 40.824
R390 VPB.n898 VPB.n897 40.824
R391 VPB.n881 VPB.n880 40.824
R392 VPB.n815 VPB.n814 40.824
R393 VPB.n798 VPB.n797 40.824
R394 VPB.n732 VPB.n731 40.824
R395 VPB.n715 VPB.n714 40.824
R396 VPB.n649 VPB.n648 40.824
R397 VPB.n632 VPB.n631 40.824
R398 VPB.n566 VPB.n565 40.824
R399 VPB.n549 VPB.n548 40.824
R400 VPB.n483 VPB.n482 40.824
R401 VPB.n466 VPB.n465 40.824
R402 VPB.n400 VPB.n399 40.824
R403 VPB.n383 VPB.n382 40.824
R404 VPB.n205 VPB.n204 35.118
R405 VPB.n1679 VPB.n1675 20.452
R406 VPB.n194 VPB.n191 20.452
R407 VPB.n318 VPB.n317 17.801
R408 VPB.n390 VPB.n389 17.801
R409 VPB.n473 VPB.n472 17.801
R410 VPB.n556 VPB.n555 17.801
R411 VPB.n639 VPB.n638 17.801
R412 VPB.n722 VPB.n721 17.801
R413 VPB.n805 VPB.n804 17.801
R414 VPB.n888 VPB.n887 17.801
R415 VPB.n148 VPB.n147 17.801
R416 VPB.n965 VPB.n964 17.801
R417 VPB.n1048 VPB.n1047 17.801
R418 VPB.n1131 VPB.n1130 17.801
R419 VPB.n1214 VPB.n1213 17.801
R420 VPB.n1297 VPB.n1296 17.801
R421 VPB.n1380 VPB.n1379 17.801
R422 VPB.n1463 VPB.n1462 17.801
R423 VPB.n1546 VPB.n1545 17.801
R424 VPB.n1629 VPB.n1628 17.801
R425 VPB.n59 VPB.n58 17.801
R426 VPB.n14 VPB.t88 14.282
R427 VPB.n14 VPB.t95 14.282
R428 VPB.n15 VPB.t26 14.282
R429 VPB.n15 VPB.t80 14.282
R430 VPB.n1638 VPB.t59 14.282
R431 VPB.n1638 VPB.t29 14.282
R432 VPB.n1621 VPB.t109 14.282
R433 VPB.n1621 VPB.t60 14.282
R434 VPB.n1555 VPB.t39 14.282
R435 VPB.n1555 VPB.t13 14.282
R436 VPB.n1538 VPB.t107 14.282
R437 VPB.n1538 VPB.t38 14.282
R438 VPB.n1472 VPB.t62 14.282
R439 VPB.n1472 VPB.t11 14.282
R440 VPB.n1455 VPB.t81 14.282
R441 VPB.n1455 VPB.t63 14.282
R442 VPB.n1389 VPB.t79 14.282
R443 VPB.n1389 VPB.t49 14.282
R444 VPB.n1372 VPB.t66 14.282
R445 VPB.n1372 VPB.t77 14.282
R446 VPB.n1306 VPB.t37 14.282
R447 VPB.n1306 VPB.t30 14.282
R448 VPB.n1289 VPB.t25 14.282
R449 VPB.n1289 VPB.t42 14.282
R450 VPB.n1223 VPB.t75 14.282
R451 VPB.n1223 VPB.t91 14.282
R452 VPB.n1206 VPB.t71 14.282
R453 VPB.n1206 VPB.t76 14.282
R454 VPB.n1140 VPB.t56 14.282
R455 VPB.n1140 VPB.t16 14.282
R456 VPB.n1123 VPB.t1 14.282
R457 VPB.n1123 VPB.t55 14.282
R458 VPB.n1057 VPB.t45 14.282
R459 VPB.n1057 VPB.t19 14.282
R460 VPB.n1040 VPB.t31 14.282
R461 VPB.n1040 VPB.t44 14.282
R462 VPB.n974 VPB.t58 14.282
R463 VPB.n974 VPB.t51 14.282
R464 VPB.n957 VPB.t86 14.282
R465 VPB.n957 VPB.t52 14.282
R466 VPB.n103 VPB.t87 14.282
R467 VPB.n103 VPB.t0 14.282
R468 VPB.n104 VPB.t7 14.282
R469 VPB.n104 VPB.t85 14.282
R470 VPB.n897 VPB.t41 14.282
R471 VPB.n897 VPB.t50 14.282
R472 VPB.n880 VPB.t32 14.282
R473 VPB.n880 VPB.t40 14.282
R474 VPB.n814 VPB.t74 14.282
R475 VPB.n814 VPB.t90 14.282
R476 VPB.n797 VPB.t20 14.282
R477 VPB.n797 VPB.t89 14.282
R478 VPB.n731 VPB.t57 14.282
R479 VPB.n731 VPB.t69 14.282
R480 VPB.n714 VPB.t36 14.282
R481 VPB.n714 VPB.t61 14.282
R482 VPB.n648 VPB.t46 14.282
R483 VPB.n648 VPB.t70 14.282
R484 VPB.n631 VPB.t9 14.282
R485 VPB.n631 VPB.t43 14.282
R486 VPB.n565 VPB.t54 14.282
R487 VPB.n565 VPB.t33 14.282
R488 VPB.n548 VPB.t82 14.282
R489 VPB.n548 VPB.t53 14.282
R490 VPB.n482 VPB.t84 14.282
R491 VPB.n482 VPB.t22 14.282
R492 VPB.n465 VPB.t111 14.282
R493 VPB.n465 VPB.t78 14.282
R494 VPB.n399 VPB.t47 14.282
R495 VPB.n399 VPB.t4 14.282
R496 VPB.n382 VPB.t2 14.282
R497 VPB.n382 VPB.t48 14.282
R498 VPB.n315 VPB.t98 14.282
R499 VPB.n315 VPB.t105 14.282
R500 VPB.n194 VPB.n193 13.653
R501 VPB.n193 VPB.n192 13.653
R502 VPB.n203 VPB.n202 13.653
R503 VPB.n202 VPB.n201 13.653
R504 VPB.n200 VPB.n199 13.653
R505 VPB.n199 VPB.n198 13.653
R506 VPB.n197 VPB.n196 13.653
R507 VPB.n196 VPB.n195 13.653
R508 VPB.n209 VPB.n208 13.653
R509 VPB.n208 VPB.n207 13.653
R510 VPB.n213 VPB.n212 13.653
R511 VPB.n212 VPB.n211 13.653
R512 VPB.n217 VPB.n216 13.653
R513 VPB.n216 VPB.n215 13.653
R514 VPB.n221 VPB.n220 13.653
R515 VPB.n220 VPB.n219 13.653
R516 VPB.n248 VPB.n247 13.653
R517 VPB.n247 VPB.n246 13.653
R518 VPB.n252 VPB.n251 13.653
R519 VPB.n251 VPB.n250 13.653
R520 VPB.n256 VPB.n255 13.653
R521 VPB.n255 VPB.n254 13.653
R522 VPB.n260 VPB.n259 13.653
R523 VPB.n259 VPB.n258 13.653
R524 VPB.n264 VPB.n263 13.653
R525 VPB.n263 VPB.n262 13.653
R526 VPB.n268 VPB.n267 13.653
R527 VPB.n267 VPB.n266 13.653
R528 VPB.n272 VPB.n271 13.653
R529 VPB.n271 VPB.n270 13.653
R530 VPB.n276 VPB.n275 13.653
R531 VPB.n275 VPB.n274 13.653
R532 VPB.n303 VPB.n302 13.653
R533 VPB.n302 VPB.n301 13.653
R534 VPB.n308 VPB.n307 13.653
R535 VPB.n307 VPB.n306 13.653
R536 VPB.n313 VPB.n312 13.653
R537 VPB.n312 VPB.n311 13.653
R538 VPB.n320 VPB.n319 13.653
R539 VPB.n319 VPB.n318 13.653
R540 VPB.n325 VPB.n324 13.653
R541 VPB.n324 VPB.n323 13.653
R542 VPB.n330 VPB.n329 13.653
R543 VPB.n329 VPB.n328 13.653
R544 VPB.n335 VPB.n334 13.653
R545 VPB.n334 VPB.n333 13.653
R546 VPB.n339 VPB.n338 13.653
R547 VPB.n338 VPB.n337 13.653
R548 VPB.n366 VPB.n365 13.653
R549 VPB.n365 VPB.n364 13.653
R550 VPB.n370 VPB.n369 13.653
R551 VPB.n369 VPB.n368 13.653
R552 VPB.n375 VPB.n374 13.653
R553 VPB.n374 VPB.n373 13.653
R554 VPB.n380 VPB.n379 13.653
R555 VPB.n379 VPB.n378 13.653
R556 VPB.n387 VPB.n386 13.653
R557 VPB.n386 VPB.n385 13.653
R558 VPB.n392 VPB.n391 13.653
R559 VPB.n391 VPB.n390 13.653
R560 VPB.n397 VPB.n396 13.653
R561 VPB.n396 VPB.n395 13.653
R562 VPB.n404 VPB.n403 13.653
R563 VPB.n403 VPB.n402 13.653
R564 VPB.n409 VPB.n408 13.653
R565 VPB.n408 VPB.n407 13.653
R566 VPB.n414 VPB.n413 13.653
R567 VPB.n413 VPB.n412 13.653
R568 VPB.n418 VPB.n417 13.653
R569 VPB.n417 VPB.n416 13.653
R570 VPB.n422 VPB.n421 13.653
R571 VPB.n421 VPB.n420 13.653
R572 VPB.n449 VPB.n448 13.653
R573 VPB.n448 VPB.n447 13.653
R574 VPB.n453 VPB.n452 13.653
R575 VPB.n452 VPB.n451 13.653
R576 VPB.n458 VPB.n457 13.653
R577 VPB.n457 VPB.n456 13.653
R578 VPB.n463 VPB.n462 13.653
R579 VPB.n462 VPB.n461 13.653
R580 VPB.n470 VPB.n469 13.653
R581 VPB.n469 VPB.n468 13.653
R582 VPB.n475 VPB.n474 13.653
R583 VPB.n474 VPB.n473 13.653
R584 VPB.n480 VPB.n479 13.653
R585 VPB.n479 VPB.n478 13.653
R586 VPB.n487 VPB.n486 13.653
R587 VPB.n486 VPB.n485 13.653
R588 VPB.n492 VPB.n491 13.653
R589 VPB.n491 VPB.n490 13.653
R590 VPB.n497 VPB.n496 13.653
R591 VPB.n496 VPB.n495 13.653
R592 VPB.n501 VPB.n500 13.653
R593 VPB.n500 VPB.n499 13.653
R594 VPB.n505 VPB.n504 13.653
R595 VPB.n504 VPB.n503 13.653
R596 VPB.n532 VPB.n531 13.653
R597 VPB.n531 VPB.n530 13.653
R598 VPB.n536 VPB.n535 13.653
R599 VPB.n535 VPB.n534 13.653
R600 VPB.n541 VPB.n540 13.653
R601 VPB.n540 VPB.n539 13.653
R602 VPB.n546 VPB.n545 13.653
R603 VPB.n545 VPB.n544 13.653
R604 VPB.n553 VPB.n552 13.653
R605 VPB.n552 VPB.n551 13.653
R606 VPB.n558 VPB.n557 13.653
R607 VPB.n557 VPB.n556 13.653
R608 VPB.n563 VPB.n562 13.653
R609 VPB.n562 VPB.n561 13.653
R610 VPB.n570 VPB.n569 13.653
R611 VPB.n569 VPB.n568 13.653
R612 VPB.n575 VPB.n574 13.653
R613 VPB.n574 VPB.n573 13.653
R614 VPB.n580 VPB.n579 13.653
R615 VPB.n579 VPB.n578 13.653
R616 VPB.n584 VPB.n583 13.653
R617 VPB.n583 VPB.n582 13.653
R618 VPB.n588 VPB.n587 13.653
R619 VPB.n587 VPB.n586 13.653
R620 VPB.n615 VPB.n614 13.653
R621 VPB.n614 VPB.n613 13.653
R622 VPB.n619 VPB.n618 13.653
R623 VPB.n618 VPB.n617 13.653
R624 VPB.n624 VPB.n623 13.653
R625 VPB.n623 VPB.n622 13.653
R626 VPB.n629 VPB.n628 13.653
R627 VPB.n628 VPB.n627 13.653
R628 VPB.n636 VPB.n635 13.653
R629 VPB.n635 VPB.n634 13.653
R630 VPB.n641 VPB.n640 13.653
R631 VPB.n640 VPB.n639 13.653
R632 VPB.n646 VPB.n645 13.653
R633 VPB.n645 VPB.n644 13.653
R634 VPB.n653 VPB.n652 13.653
R635 VPB.n652 VPB.n651 13.653
R636 VPB.n658 VPB.n657 13.653
R637 VPB.n657 VPB.n656 13.653
R638 VPB.n663 VPB.n662 13.653
R639 VPB.n662 VPB.n661 13.653
R640 VPB.n667 VPB.n666 13.653
R641 VPB.n666 VPB.n665 13.653
R642 VPB.n671 VPB.n670 13.653
R643 VPB.n670 VPB.n669 13.653
R644 VPB.n698 VPB.n697 13.653
R645 VPB.n697 VPB.n696 13.653
R646 VPB.n702 VPB.n701 13.653
R647 VPB.n701 VPB.n700 13.653
R648 VPB.n707 VPB.n706 13.653
R649 VPB.n706 VPB.n705 13.653
R650 VPB.n712 VPB.n711 13.653
R651 VPB.n711 VPB.n710 13.653
R652 VPB.n719 VPB.n718 13.653
R653 VPB.n718 VPB.n717 13.653
R654 VPB.n724 VPB.n723 13.653
R655 VPB.n723 VPB.n722 13.653
R656 VPB.n729 VPB.n728 13.653
R657 VPB.n728 VPB.n727 13.653
R658 VPB.n736 VPB.n735 13.653
R659 VPB.n735 VPB.n734 13.653
R660 VPB.n741 VPB.n740 13.653
R661 VPB.n740 VPB.n739 13.653
R662 VPB.n746 VPB.n745 13.653
R663 VPB.n745 VPB.n744 13.653
R664 VPB.n750 VPB.n749 13.653
R665 VPB.n749 VPB.n748 13.653
R666 VPB.n754 VPB.n753 13.653
R667 VPB.n753 VPB.n752 13.653
R668 VPB.n781 VPB.n780 13.653
R669 VPB.n780 VPB.n779 13.653
R670 VPB.n785 VPB.n784 13.653
R671 VPB.n784 VPB.n783 13.653
R672 VPB.n790 VPB.n789 13.653
R673 VPB.n789 VPB.n788 13.653
R674 VPB.n795 VPB.n794 13.653
R675 VPB.n794 VPB.n793 13.653
R676 VPB.n802 VPB.n801 13.653
R677 VPB.n801 VPB.n800 13.653
R678 VPB.n807 VPB.n806 13.653
R679 VPB.n806 VPB.n805 13.653
R680 VPB.n812 VPB.n811 13.653
R681 VPB.n811 VPB.n810 13.653
R682 VPB.n819 VPB.n818 13.653
R683 VPB.n818 VPB.n817 13.653
R684 VPB.n824 VPB.n823 13.653
R685 VPB.n823 VPB.n822 13.653
R686 VPB.n829 VPB.n828 13.653
R687 VPB.n828 VPB.n827 13.653
R688 VPB.n833 VPB.n832 13.653
R689 VPB.n832 VPB.n831 13.653
R690 VPB.n837 VPB.n836 13.653
R691 VPB.n836 VPB.n835 13.653
R692 VPB.n864 VPB.n863 13.653
R693 VPB.n863 VPB.n862 13.653
R694 VPB.n868 VPB.n867 13.653
R695 VPB.n867 VPB.n866 13.653
R696 VPB.n873 VPB.n872 13.653
R697 VPB.n872 VPB.n871 13.653
R698 VPB.n878 VPB.n877 13.653
R699 VPB.n877 VPB.n876 13.653
R700 VPB.n885 VPB.n884 13.653
R701 VPB.n884 VPB.n883 13.653
R702 VPB.n890 VPB.n889 13.653
R703 VPB.n889 VPB.n888 13.653
R704 VPB.n895 VPB.n894 13.653
R705 VPB.n894 VPB.n893 13.653
R706 VPB.n902 VPB.n901 13.653
R707 VPB.n901 VPB.n900 13.653
R708 VPB.n907 VPB.n906 13.653
R709 VPB.n906 VPB.n905 13.653
R710 VPB.n912 VPB.n911 13.653
R711 VPB.n911 VPB.n910 13.653
R712 VPB.n916 VPB.n915 13.653
R713 VPB.n915 VPB.n914 13.653
R714 VPB.n920 VPB.n919 13.653
R715 VPB.n919 VPB.n918 13.653
R716 VPB.n130 VPB.n129 13.653
R717 VPB.n129 VPB.n128 13.653
R718 VPB.n133 VPB.n132 13.653
R719 VPB.n132 VPB.n131 13.653
R720 VPB.n137 VPB.n136 13.653
R721 VPB.n136 VPB.n135 13.653
R722 VPB.n141 VPB.n140 13.653
R723 VPB.n140 VPB.n139 13.653
R724 VPB.n145 VPB.n144 13.653
R725 VPB.n144 VPB.n143 13.653
R726 VPB.n150 VPB.n149 13.653
R727 VPB.n149 VPB.n148 13.653
R728 VPB.n154 VPB.n153 13.653
R729 VPB.n153 VPB.n152 13.653
R730 VPB.n159 VPB.n158 13.653
R731 VPB.n158 VPB.n157 13.653
R732 VPB.n163 VPB.n162 13.653
R733 VPB.n162 VPB.n161 13.653
R734 VPB.n166 VPB.n165 13.653
R735 VPB.n165 VPB.n164 13.653
R736 VPB.n170 VPB.n169 13.653
R737 VPB.n169 VPB.n168 13.653
R738 VPB.n936 VPB.n935 13.653
R739 VPB.n935 VPB.n934 13.653
R740 VPB.n941 VPB.n940 13.653
R741 VPB.n940 VPB.n939 13.653
R742 VPB.n945 VPB.n944 13.653
R743 VPB.n944 VPB.n943 13.653
R744 VPB.n950 VPB.n949 13.653
R745 VPB.n949 VPB.n948 13.653
R746 VPB.n955 VPB.n954 13.653
R747 VPB.n954 VPB.n953 13.653
R748 VPB.n962 VPB.n961 13.653
R749 VPB.n961 VPB.n960 13.653
R750 VPB.n967 VPB.n966 13.653
R751 VPB.n966 VPB.n965 13.653
R752 VPB.n972 VPB.n971 13.653
R753 VPB.n971 VPB.n970 13.653
R754 VPB.n979 VPB.n978 13.653
R755 VPB.n978 VPB.n977 13.653
R756 VPB.n984 VPB.n983 13.653
R757 VPB.n983 VPB.n982 13.653
R758 VPB.n989 VPB.n988 13.653
R759 VPB.n988 VPB.n987 13.653
R760 VPB.n993 VPB.n992 13.653
R761 VPB.n992 VPB.n991 13.653
R762 VPB.n997 VPB.n996 13.653
R763 VPB.n996 VPB.n995 13.653
R764 VPB.n1024 VPB.n1023 13.653
R765 VPB.n1023 VPB.n1022 13.653
R766 VPB.n1028 VPB.n1027 13.653
R767 VPB.n1027 VPB.n1026 13.653
R768 VPB.n1033 VPB.n1032 13.653
R769 VPB.n1032 VPB.n1031 13.653
R770 VPB.n1038 VPB.n1037 13.653
R771 VPB.n1037 VPB.n1036 13.653
R772 VPB.n1045 VPB.n1044 13.653
R773 VPB.n1044 VPB.n1043 13.653
R774 VPB.n1050 VPB.n1049 13.653
R775 VPB.n1049 VPB.n1048 13.653
R776 VPB.n1055 VPB.n1054 13.653
R777 VPB.n1054 VPB.n1053 13.653
R778 VPB.n1062 VPB.n1061 13.653
R779 VPB.n1061 VPB.n1060 13.653
R780 VPB.n1067 VPB.n1066 13.653
R781 VPB.n1066 VPB.n1065 13.653
R782 VPB.n1072 VPB.n1071 13.653
R783 VPB.n1071 VPB.n1070 13.653
R784 VPB.n1076 VPB.n1075 13.653
R785 VPB.n1075 VPB.n1074 13.653
R786 VPB.n1080 VPB.n1079 13.653
R787 VPB.n1079 VPB.n1078 13.653
R788 VPB.n1107 VPB.n1106 13.653
R789 VPB.n1106 VPB.n1105 13.653
R790 VPB.n1111 VPB.n1110 13.653
R791 VPB.n1110 VPB.n1109 13.653
R792 VPB.n1116 VPB.n1115 13.653
R793 VPB.n1115 VPB.n1114 13.653
R794 VPB.n1121 VPB.n1120 13.653
R795 VPB.n1120 VPB.n1119 13.653
R796 VPB.n1128 VPB.n1127 13.653
R797 VPB.n1127 VPB.n1126 13.653
R798 VPB.n1133 VPB.n1132 13.653
R799 VPB.n1132 VPB.n1131 13.653
R800 VPB.n1138 VPB.n1137 13.653
R801 VPB.n1137 VPB.n1136 13.653
R802 VPB.n1145 VPB.n1144 13.653
R803 VPB.n1144 VPB.n1143 13.653
R804 VPB.n1150 VPB.n1149 13.653
R805 VPB.n1149 VPB.n1148 13.653
R806 VPB.n1155 VPB.n1154 13.653
R807 VPB.n1154 VPB.n1153 13.653
R808 VPB.n1159 VPB.n1158 13.653
R809 VPB.n1158 VPB.n1157 13.653
R810 VPB.n1163 VPB.n1162 13.653
R811 VPB.n1162 VPB.n1161 13.653
R812 VPB.n1190 VPB.n1189 13.653
R813 VPB.n1189 VPB.n1188 13.653
R814 VPB.n1194 VPB.n1193 13.653
R815 VPB.n1193 VPB.n1192 13.653
R816 VPB.n1199 VPB.n1198 13.653
R817 VPB.n1198 VPB.n1197 13.653
R818 VPB.n1204 VPB.n1203 13.653
R819 VPB.n1203 VPB.n1202 13.653
R820 VPB.n1211 VPB.n1210 13.653
R821 VPB.n1210 VPB.n1209 13.653
R822 VPB.n1216 VPB.n1215 13.653
R823 VPB.n1215 VPB.n1214 13.653
R824 VPB.n1221 VPB.n1220 13.653
R825 VPB.n1220 VPB.n1219 13.653
R826 VPB.n1228 VPB.n1227 13.653
R827 VPB.n1227 VPB.n1226 13.653
R828 VPB.n1233 VPB.n1232 13.653
R829 VPB.n1232 VPB.n1231 13.653
R830 VPB.n1238 VPB.n1237 13.653
R831 VPB.n1237 VPB.n1236 13.653
R832 VPB.n1242 VPB.n1241 13.653
R833 VPB.n1241 VPB.n1240 13.653
R834 VPB.n1246 VPB.n1245 13.653
R835 VPB.n1245 VPB.n1244 13.653
R836 VPB.n1273 VPB.n1272 13.653
R837 VPB.n1272 VPB.n1271 13.653
R838 VPB.n1277 VPB.n1276 13.653
R839 VPB.n1276 VPB.n1275 13.653
R840 VPB.n1282 VPB.n1281 13.653
R841 VPB.n1281 VPB.n1280 13.653
R842 VPB.n1287 VPB.n1286 13.653
R843 VPB.n1286 VPB.n1285 13.653
R844 VPB.n1294 VPB.n1293 13.653
R845 VPB.n1293 VPB.n1292 13.653
R846 VPB.n1299 VPB.n1298 13.653
R847 VPB.n1298 VPB.n1297 13.653
R848 VPB.n1304 VPB.n1303 13.653
R849 VPB.n1303 VPB.n1302 13.653
R850 VPB.n1311 VPB.n1310 13.653
R851 VPB.n1310 VPB.n1309 13.653
R852 VPB.n1316 VPB.n1315 13.653
R853 VPB.n1315 VPB.n1314 13.653
R854 VPB.n1321 VPB.n1320 13.653
R855 VPB.n1320 VPB.n1319 13.653
R856 VPB.n1325 VPB.n1324 13.653
R857 VPB.n1324 VPB.n1323 13.653
R858 VPB.n1329 VPB.n1328 13.653
R859 VPB.n1328 VPB.n1327 13.653
R860 VPB.n1356 VPB.n1355 13.653
R861 VPB.n1355 VPB.n1354 13.653
R862 VPB.n1360 VPB.n1359 13.653
R863 VPB.n1359 VPB.n1358 13.653
R864 VPB.n1365 VPB.n1364 13.653
R865 VPB.n1364 VPB.n1363 13.653
R866 VPB.n1370 VPB.n1369 13.653
R867 VPB.n1369 VPB.n1368 13.653
R868 VPB.n1377 VPB.n1376 13.653
R869 VPB.n1376 VPB.n1375 13.653
R870 VPB.n1382 VPB.n1381 13.653
R871 VPB.n1381 VPB.n1380 13.653
R872 VPB.n1387 VPB.n1386 13.653
R873 VPB.n1386 VPB.n1385 13.653
R874 VPB.n1394 VPB.n1393 13.653
R875 VPB.n1393 VPB.n1392 13.653
R876 VPB.n1399 VPB.n1398 13.653
R877 VPB.n1398 VPB.n1397 13.653
R878 VPB.n1404 VPB.n1403 13.653
R879 VPB.n1403 VPB.n1402 13.653
R880 VPB.n1408 VPB.n1407 13.653
R881 VPB.n1407 VPB.n1406 13.653
R882 VPB.n1412 VPB.n1411 13.653
R883 VPB.n1411 VPB.n1410 13.653
R884 VPB.n1439 VPB.n1438 13.653
R885 VPB.n1438 VPB.n1437 13.653
R886 VPB.n1443 VPB.n1442 13.653
R887 VPB.n1442 VPB.n1441 13.653
R888 VPB.n1448 VPB.n1447 13.653
R889 VPB.n1447 VPB.n1446 13.653
R890 VPB.n1453 VPB.n1452 13.653
R891 VPB.n1452 VPB.n1451 13.653
R892 VPB.n1460 VPB.n1459 13.653
R893 VPB.n1459 VPB.n1458 13.653
R894 VPB.n1465 VPB.n1464 13.653
R895 VPB.n1464 VPB.n1463 13.653
R896 VPB.n1470 VPB.n1469 13.653
R897 VPB.n1469 VPB.n1468 13.653
R898 VPB.n1477 VPB.n1476 13.653
R899 VPB.n1476 VPB.n1475 13.653
R900 VPB.n1482 VPB.n1481 13.653
R901 VPB.n1481 VPB.n1480 13.653
R902 VPB.n1487 VPB.n1486 13.653
R903 VPB.n1486 VPB.n1485 13.653
R904 VPB.n1491 VPB.n1490 13.653
R905 VPB.n1490 VPB.n1489 13.653
R906 VPB.n1495 VPB.n1494 13.653
R907 VPB.n1494 VPB.n1493 13.653
R908 VPB.n1522 VPB.n1521 13.653
R909 VPB.n1521 VPB.n1520 13.653
R910 VPB.n1526 VPB.n1525 13.653
R911 VPB.n1525 VPB.n1524 13.653
R912 VPB.n1531 VPB.n1530 13.653
R913 VPB.n1530 VPB.n1529 13.653
R914 VPB.n1536 VPB.n1535 13.653
R915 VPB.n1535 VPB.n1534 13.653
R916 VPB.n1543 VPB.n1542 13.653
R917 VPB.n1542 VPB.n1541 13.653
R918 VPB.n1548 VPB.n1547 13.653
R919 VPB.n1547 VPB.n1546 13.653
R920 VPB.n1553 VPB.n1552 13.653
R921 VPB.n1552 VPB.n1551 13.653
R922 VPB.n1560 VPB.n1559 13.653
R923 VPB.n1559 VPB.n1558 13.653
R924 VPB.n1565 VPB.n1564 13.653
R925 VPB.n1564 VPB.n1563 13.653
R926 VPB.n1570 VPB.n1569 13.653
R927 VPB.n1569 VPB.n1568 13.653
R928 VPB.n1574 VPB.n1573 13.653
R929 VPB.n1573 VPB.n1572 13.653
R930 VPB.n1578 VPB.n1577 13.653
R931 VPB.n1577 VPB.n1576 13.653
R932 VPB.n1605 VPB.n1604 13.653
R933 VPB.n1604 VPB.n1603 13.653
R934 VPB.n1609 VPB.n1608 13.653
R935 VPB.n1608 VPB.n1607 13.653
R936 VPB.n1614 VPB.n1613 13.653
R937 VPB.n1613 VPB.n1612 13.653
R938 VPB.n1619 VPB.n1618 13.653
R939 VPB.n1618 VPB.n1617 13.653
R940 VPB.n1626 VPB.n1625 13.653
R941 VPB.n1625 VPB.n1624 13.653
R942 VPB.n1631 VPB.n1630 13.653
R943 VPB.n1630 VPB.n1629 13.653
R944 VPB.n1636 VPB.n1635 13.653
R945 VPB.n1635 VPB.n1634 13.653
R946 VPB.n1643 VPB.n1642 13.653
R947 VPB.n1642 VPB.n1641 13.653
R948 VPB.n1648 VPB.n1647 13.653
R949 VPB.n1647 VPB.n1646 13.653
R950 VPB.n1653 VPB.n1652 13.653
R951 VPB.n1652 VPB.n1651 13.653
R952 VPB.n1657 VPB.n1656 13.653
R953 VPB.n1656 VPB.n1655 13.653
R954 VPB.n1661 VPB.n1660 13.653
R955 VPB.n1660 VPB.n1659 13.653
R956 VPB.n41 VPB.n40 13.653
R957 VPB.n40 VPB.n39 13.653
R958 VPB.n44 VPB.n43 13.653
R959 VPB.n43 VPB.n42 13.653
R960 VPB.n48 VPB.n47 13.653
R961 VPB.n47 VPB.n46 13.653
R962 VPB.n52 VPB.n51 13.653
R963 VPB.n51 VPB.n50 13.653
R964 VPB.n56 VPB.n55 13.653
R965 VPB.n55 VPB.n54 13.653
R966 VPB.n61 VPB.n60 13.653
R967 VPB.n60 VPB.n59 13.653
R968 VPB.n65 VPB.n64 13.653
R969 VPB.n64 VPB.n63 13.653
R970 VPB.n70 VPB.n69 13.653
R971 VPB.n69 VPB.n68 13.653
R972 VPB.n74 VPB.n73 13.653
R973 VPB.n73 VPB.n72 13.653
R974 VPB.n77 VPB.n76 13.653
R975 VPB.n76 VPB.n75 13.653
R976 VPB.n81 VPB.n80 13.653
R977 VPB.n80 VPB.n79 13.653
R978 VPB.n1675 VPB.n0 13.653
R979 VPB VPB.n0 13.653
R980 VPB.n323 VPB.n322 13.35
R981 VPB.n395 VPB.n394 13.35
R982 VPB.n478 VPB.n477 13.35
R983 VPB.n561 VPB.n560 13.35
R984 VPB.n644 VPB.n643 13.35
R985 VPB.n727 VPB.n726 13.35
R986 VPB.n810 VPB.n809 13.35
R987 VPB.n893 VPB.n892 13.35
R988 VPB.n152 VPB.n151 13.35
R989 VPB.n970 VPB.n969 13.35
R990 VPB.n1053 VPB.n1052 13.35
R991 VPB.n1136 VPB.n1135 13.35
R992 VPB.n1219 VPB.n1218 13.35
R993 VPB.n1302 VPB.n1301 13.35
R994 VPB.n1385 VPB.n1384 13.35
R995 VPB.n1468 VPB.n1467 13.35
R996 VPB.n1551 VPB.n1550 13.35
R997 VPB.n1634 VPB.n1633 13.35
R998 VPB.n63 VPB.n62 13.35
R999 VPB.n1679 VPB.n1678 13.276
R1000 VPB.n1678 VPB.n1676 13.276
R1001 VPB.n36 VPB.n18 13.276
R1002 VPB.n18 VPB.n16 13.276
R1003 VPB.n1600 VPB.n1582 13.276
R1004 VPB.n1582 VPB.n1580 13.276
R1005 VPB.n1517 VPB.n1499 13.276
R1006 VPB.n1499 VPB.n1497 13.276
R1007 VPB.n1434 VPB.n1416 13.276
R1008 VPB.n1416 VPB.n1414 13.276
R1009 VPB.n1351 VPB.n1333 13.276
R1010 VPB.n1333 VPB.n1331 13.276
R1011 VPB.n1268 VPB.n1250 13.276
R1012 VPB.n1250 VPB.n1248 13.276
R1013 VPB.n1185 VPB.n1167 13.276
R1014 VPB.n1167 VPB.n1165 13.276
R1015 VPB.n1102 VPB.n1084 13.276
R1016 VPB.n1084 VPB.n1082 13.276
R1017 VPB.n1019 VPB.n1001 13.276
R1018 VPB.n1001 VPB.n999 13.276
R1019 VPB.n102 VPB.n84 13.276
R1020 VPB.n84 VPB.n82 13.276
R1021 VPB.n125 VPB.n107 13.276
R1022 VPB.n107 VPB.n105 13.276
R1023 VPB.n859 VPB.n841 13.276
R1024 VPB.n841 VPB.n839 13.276
R1025 VPB.n776 VPB.n758 13.276
R1026 VPB.n758 VPB.n756 13.276
R1027 VPB.n693 VPB.n675 13.276
R1028 VPB.n675 VPB.n673 13.276
R1029 VPB.n610 VPB.n592 13.276
R1030 VPB.n592 VPB.n590 13.276
R1031 VPB.n527 VPB.n509 13.276
R1032 VPB.n509 VPB.n507 13.276
R1033 VPB.n444 VPB.n426 13.276
R1034 VPB.n426 VPB.n424 13.276
R1035 VPB.n361 VPB.n343 13.276
R1036 VPB.n343 VPB.n341 13.276
R1037 VPB.n298 VPB.n280 13.276
R1038 VPB.n280 VPB.n278 13.276
R1039 VPB.n243 VPB.n225 13.276
R1040 VPB.n225 VPB.n223 13.276
R1041 VPB.n203 VPB.n200 13.276
R1042 VPB.n200 VPB.n197 13.276
R1043 VPB.n248 VPB.n244 13.276
R1044 VPB.n303 VPB.n299 13.276
R1045 VPB.n366 VPB.n362 13.276
R1046 VPB.n449 VPB.n445 13.276
R1047 VPB.n532 VPB.n528 13.276
R1048 VPB.n615 VPB.n611 13.276
R1049 VPB.n698 VPB.n694 13.276
R1050 VPB.n781 VPB.n777 13.276
R1051 VPB.n864 VPB.n860 13.276
R1052 VPB.n130 VPB.n126 13.276
R1053 VPB.n133 VPB.n130 13.276
R1054 VPB.n141 VPB.n137 13.276
R1055 VPB.n145 VPB.n141 13.276
R1056 VPB.n154 VPB.n150 13.276
R1057 VPB.n163 VPB.n159 13.276
R1058 VPB.n166 VPB.n163 13.276
R1059 VPB.n936 VPB.n170 13.276
R1060 VPB.n937 VPB.n936 13.276
R1061 VPB.n941 VPB.n937 13.276
R1062 VPB.n1024 VPB.n1020 13.276
R1063 VPB.n1107 VPB.n1103 13.276
R1064 VPB.n1190 VPB.n1186 13.276
R1065 VPB.n1273 VPB.n1269 13.276
R1066 VPB.n1356 VPB.n1352 13.276
R1067 VPB.n1439 VPB.n1435 13.276
R1068 VPB.n1522 VPB.n1518 13.276
R1069 VPB.n1605 VPB.n1601 13.276
R1070 VPB.n41 VPB.n37 13.276
R1071 VPB.n44 VPB.n41 13.276
R1072 VPB.n52 VPB.n48 13.276
R1073 VPB.n56 VPB.n52 13.276
R1074 VPB.n65 VPB.n61 13.276
R1075 VPB.n74 VPB.n70 13.276
R1076 VPB.n77 VPB.n74 13.276
R1077 VPB.n1675 VPB.n81 13.276
R1078 VPB.n191 VPB.n173 13.276
R1079 VPB.n173 VPB.n171 13.276
R1080 VPB.n178 VPB.n176 12.796
R1081 VPB.n178 VPB.n177 12.564
R1082 VPB.n170 VPB.n167 12.558
R1083 VPB.n81 VPB.n78 12.558
R1084 VPB.n134 VPB.n133 12.2
R1085 VPB.n45 VPB.n44 12.2
R1086 VPB.n186 VPB.n185 12.198
R1087 VPB.n184 VPB.n183 12.198
R1088 VPB.n181 VPB.n180 12.198
R1089 VPB.n150 VPB.n146 9.329
R1090 VPB.n61 VPB.n57 9.329
R1091 VPB.n155 VPB.n154 8.97
R1092 VPB.n66 VPB.n65 8.97
R1093 VPB.n191 VPB.n190 7.5
R1094 VPB.n176 VPB.n175 7.5
R1095 VPB.n180 VPB.n179 7.5
R1096 VPB.n183 VPB.n182 7.5
R1097 VPB.n173 VPB.n172 7.5
R1098 VPB.n188 VPB.n174 7.5
R1099 VPB.n225 VPB.n224 7.5
R1100 VPB.n238 VPB.n237 7.5
R1101 VPB.n232 VPB.n231 7.5
R1102 VPB.n234 VPB.n233 7.5
R1103 VPB.n227 VPB.n226 7.5
R1104 VPB.n243 VPB.n242 7.5
R1105 VPB.n280 VPB.n279 7.5
R1106 VPB.n293 VPB.n292 7.5
R1107 VPB.n287 VPB.n286 7.5
R1108 VPB.n289 VPB.n288 7.5
R1109 VPB.n282 VPB.n281 7.5
R1110 VPB.n298 VPB.n297 7.5
R1111 VPB.n343 VPB.n342 7.5
R1112 VPB.n356 VPB.n355 7.5
R1113 VPB.n350 VPB.n349 7.5
R1114 VPB.n352 VPB.n351 7.5
R1115 VPB.n345 VPB.n344 7.5
R1116 VPB.n361 VPB.n360 7.5
R1117 VPB.n426 VPB.n425 7.5
R1118 VPB.n439 VPB.n438 7.5
R1119 VPB.n433 VPB.n432 7.5
R1120 VPB.n435 VPB.n434 7.5
R1121 VPB.n428 VPB.n427 7.5
R1122 VPB.n444 VPB.n443 7.5
R1123 VPB.n509 VPB.n508 7.5
R1124 VPB.n522 VPB.n521 7.5
R1125 VPB.n516 VPB.n515 7.5
R1126 VPB.n518 VPB.n517 7.5
R1127 VPB.n511 VPB.n510 7.5
R1128 VPB.n527 VPB.n526 7.5
R1129 VPB.n592 VPB.n591 7.5
R1130 VPB.n605 VPB.n604 7.5
R1131 VPB.n599 VPB.n598 7.5
R1132 VPB.n601 VPB.n600 7.5
R1133 VPB.n594 VPB.n593 7.5
R1134 VPB.n610 VPB.n609 7.5
R1135 VPB.n675 VPB.n674 7.5
R1136 VPB.n688 VPB.n687 7.5
R1137 VPB.n682 VPB.n681 7.5
R1138 VPB.n684 VPB.n683 7.5
R1139 VPB.n677 VPB.n676 7.5
R1140 VPB.n693 VPB.n692 7.5
R1141 VPB.n758 VPB.n757 7.5
R1142 VPB.n771 VPB.n770 7.5
R1143 VPB.n765 VPB.n764 7.5
R1144 VPB.n767 VPB.n766 7.5
R1145 VPB.n760 VPB.n759 7.5
R1146 VPB.n776 VPB.n775 7.5
R1147 VPB.n841 VPB.n840 7.5
R1148 VPB.n854 VPB.n853 7.5
R1149 VPB.n848 VPB.n847 7.5
R1150 VPB.n850 VPB.n849 7.5
R1151 VPB.n843 VPB.n842 7.5
R1152 VPB.n859 VPB.n858 7.5
R1153 VPB.n107 VPB.n106 7.5
R1154 VPB.n120 VPB.n119 7.5
R1155 VPB.n114 VPB.n113 7.5
R1156 VPB.n116 VPB.n115 7.5
R1157 VPB.n109 VPB.n108 7.5
R1158 VPB.n125 VPB.n124 7.5
R1159 VPB.n84 VPB.n83 7.5
R1160 VPB.n97 VPB.n96 7.5
R1161 VPB.n91 VPB.n90 7.5
R1162 VPB.n93 VPB.n92 7.5
R1163 VPB.n86 VPB.n85 7.5
R1164 VPB.n102 VPB.n101 7.5
R1165 VPB.n1001 VPB.n1000 7.5
R1166 VPB.n1014 VPB.n1013 7.5
R1167 VPB.n1008 VPB.n1007 7.5
R1168 VPB.n1010 VPB.n1009 7.5
R1169 VPB.n1003 VPB.n1002 7.5
R1170 VPB.n1019 VPB.n1018 7.5
R1171 VPB.n1084 VPB.n1083 7.5
R1172 VPB.n1097 VPB.n1096 7.5
R1173 VPB.n1091 VPB.n1090 7.5
R1174 VPB.n1093 VPB.n1092 7.5
R1175 VPB.n1086 VPB.n1085 7.5
R1176 VPB.n1102 VPB.n1101 7.5
R1177 VPB.n1167 VPB.n1166 7.5
R1178 VPB.n1180 VPB.n1179 7.5
R1179 VPB.n1174 VPB.n1173 7.5
R1180 VPB.n1176 VPB.n1175 7.5
R1181 VPB.n1169 VPB.n1168 7.5
R1182 VPB.n1185 VPB.n1184 7.5
R1183 VPB.n1250 VPB.n1249 7.5
R1184 VPB.n1263 VPB.n1262 7.5
R1185 VPB.n1257 VPB.n1256 7.5
R1186 VPB.n1259 VPB.n1258 7.5
R1187 VPB.n1252 VPB.n1251 7.5
R1188 VPB.n1268 VPB.n1267 7.5
R1189 VPB.n1333 VPB.n1332 7.5
R1190 VPB.n1346 VPB.n1345 7.5
R1191 VPB.n1340 VPB.n1339 7.5
R1192 VPB.n1342 VPB.n1341 7.5
R1193 VPB.n1335 VPB.n1334 7.5
R1194 VPB.n1351 VPB.n1350 7.5
R1195 VPB.n1416 VPB.n1415 7.5
R1196 VPB.n1429 VPB.n1428 7.5
R1197 VPB.n1423 VPB.n1422 7.5
R1198 VPB.n1425 VPB.n1424 7.5
R1199 VPB.n1418 VPB.n1417 7.5
R1200 VPB.n1434 VPB.n1433 7.5
R1201 VPB.n1499 VPB.n1498 7.5
R1202 VPB.n1512 VPB.n1511 7.5
R1203 VPB.n1506 VPB.n1505 7.5
R1204 VPB.n1508 VPB.n1507 7.5
R1205 VPB.n1501 VPB.n1500 7.5
R1206 VPB.n1517 VPB.n1516 7.5
R1207 VPB.n1582 VPB.n1581 7.5
R1208 VPB.n1595 VPB.n1594 7.5
R1209 VPB.n1589 VPB.n1588 7.5
R1210 VPB.n1591 VPB.n1590 7.5
R1211 VPB.n1584 VPB.n1583 7.5
R1212 VPB.n1600 VPB.n1599 7.5
R1213 VPB.n18 VPB.n17 7.5
R1214 VPB.n31 VPB.n30 7.5
R1215 VPB.n25 VPB.n24 7.5
R1216 VPB.n27 VPB.n26 7.5
R1217 VPB.n20 VPB.n19 7.5
R1218 VPB.n36 VPB.n35 7.5
R1219 VPB.n1678 VPB.n1677 7.5
R1220 VPB.n12 VPB.n11 7.5
R1221 VPB.n6 VPB.n5 7.5
R1222 VPB.n8 VPB.n7 7.5
R1223 VPB.n2 VPB.n1 7.5
R1224 VPB.n1680 VPB.n1679 7.5
R1225 VPB.n37 VPB.n36 7.176
R1226 VPB.n1601 VPB.n1600 7.176
R1227 VPB.n1518 VPB.n1517 7.176
R1228 VPB.n1435 VPB.n1434 7.176
R1229 VPB.n1352 VPB.n1351 7.176
R1230 VPB.n1269 VPB.n1268 7.176
R1231 VPB.n1186 VPB.n1185 7.176
R1232 VPB.n1103 VPB.n1102 7.176
R1233 VPB.n1020 VPB.n1019 7.176
R1234 VPB.n937 VPB.n102 7.176
R1235 VPB.n126 VPB.n125 7.176
R1236 VPB.n860 VPB.n859 7.176
R1237 VPB.n777 VPB.n776 7.176
R1238 VPB.n694 VPB.n693 7.176
R1239 VPB.n611 VPB.n610 7.176
R1240 VPB.n528 VPB.n527 7.176
R1241 VPB.n445 VPB.n444 7.176
R1242 VPB.n362 VPB.n361 7.176
R1243 VPB.n299 VPB.n298 7.176
R1244 VPB.n244 VPB.n243 7.176
R1245 VPB.n239 VPB.n236 6.729
R1246 VPB.n235 VPB.n232 6.729
R1247 VPB.n230 VPB.n227 6.729
R1248 VPB.n294 VPB.n291 6.729
R1249 VPB.n290 VPB.n287 6.729
R1250 VPB.n285 VPB.n282 6.729
R1251 VPB.n357 VPB.n354 6.729
R1252 VPB.n353 VPB.n350 6.729
R1253 VPB.n348 VPB.n345 6.729
R1254 VPB.n440 VPB.n437 6.729
R1255 VPB.n436 VPB.n433 6.729
R1256 VPB.n431 VPB.n428 6.729
R1257 VPB.n523 VPB.n520 6.729
R1258 VPB.n519 VPB.n516 6.729
R1259 VPB.n514 VPB.n511 6.729
R1260 VPB.n606 VPB.n603 6.729
R1261 VPB.n602 VPB.n599 6.729
R1262 VPB.n597 VPB.n594 6.729
R1263 VPB.n689 VPB.n686 6.729
R1264 VPB.n685 VPB.n682 6.729
R1265 VPB.n680 VPB.n677 6.729
R1266 VPB.n772 VPB.n769 6.729
R1267 VPB.n768 VPB.n765 6.729
R1268 VPB.n763 VPB.n760 6.729
R1269 VPB.n855 VPB.n852 6.729
R1270 VPB.n851 VPB.n848 6.729
R1271 VPB.n846 VPB.n843 6.729
R1272 VPB.n121 VPB.n118 6.729
R1273 VPB.n117 VPB.n114 6.729
R1274 VPB.n112 VPB.n109 6.729
R1275 VPB.n98 VPB.n95 6.729
R1276 VPB.n94 VPB.n91 6.729
R1277 VPB.n89 VPB.n86 6.729
R1278 VPB.n1015 VPB.n1012 6.729
R1279 VPB.n1011 VPB.n1008 6.729
R1280 VPB.n1006 VPB.n1003 6.729
R1281 VPB.n1098 VPB.n1095 6.729
R1282 VPB.n1094 VPB.n1091 6.729
R1283 VPB.n1089 VPB.n1086 6.729
R1284 VPB.n1181 VPB.n1178 6.729
R1285 VPB.n1177 VPB.n1174 6.729
R1286 VPB.n1172 VPB.n1169 6.729
R1287 VPB.n1264 VPB.n1261 6.729
R1288 VPB.n1260 VPB.n1257 6.729
R1289 VPB.n1255 VPB.n1252 6.729
R1290 VPB.n1347 VPB.n1344 6.729
R1291 VPB.n1343 VPB.n1340 6.729
R1292 VPB.n1338 VPB.n1335 6.729
R1293 VPB.n1430 VPB.n1427 6.729
R1294 VPB.n1426 VPB.n1423 6.729
R1295 VPB.n1421 VPB.n1418 6.729
R1296 VPB.n1513 VPB.n1510 6.729
R1297 VPB.n1509 VPB.n1506 6.729
R1298 VPB.n1504 VPB.n1501 6.729
R1299 VPB.n1596 VPB.n1593 6.729
R1300 VPB.n1592 VPB.n1589 6.729
R1301 VPB.n1587 VPB.n1584 6.729
R1302 VPB.n32 VPB.n29 6.729
R1303 VPB.n28 VPB.n25 6.729
R1304 VPB.n23 VPB.n20 6.729
R1305 VPB.n13 VPB.n10 6.729
R1306 VPB.n9 VPB.n6 6.729
R1307 VPB.n4 VPB.n2 6.729
R1308 VPB.n230 VPB.n229 6.728
R1309 VPB.n235 VPB.n234 6.728
R1310 VPB.n239 VPB.n238 6.728
R1311 VPB.n242 VPB.n241 6.728
R1312 VPB.n285 VPB.n284 6.728
R1313 VPB.n290 VPB.n289 6.728
R1314 VPB.n294 VPB.n293 6.728
R1315 VPB.n297 VPB.n296 6.728
R1316 VPB.n348 VPB.n347 6.728
R1317 VPB.n353 VPB.n352 6.728
R1318 VPB.n357 VPB.n356 6.728
R1319 VPB.n360 VPB.n359 6.728
R1320 VPB.n431 VPB.n430 6.728
R1321 VPB.n436 VPB.n435 6.728
R1322 VPB.n440 VPB.n439 6.728
R1323 VPB.n443 VPB.n442 6.728
R1324 VPB.n514 VPB.n513 6.728
R1325 VPB.n519 VPB.n518 6.728
R1326 VPB.n523 VPB.n522 6.728
R1327 VPB.n526 VPB.n525 6.728
R1328 VPB.n597 VPB.n596 6.728
R1329 VPB.n602 VPB.n601 6.728
R1330 VPB.n606 VPB.n605 6.728
R1331 VPB.n609 VPB.n608 6.728
R1332 VPB.n680 VPB.n679 6.728
R1333 VPB.n685 VPB.n684 6.728
R1334 VPB.n689 VPB.n688 6.728
R1335 VPB.n692 VPB.n691 6.728
R1336 VPB.n763 VPB.n762 6.728
R1337 VPB.n768 VPB.n767 6.728
R1338 VPB.n772 VPB.n771 6.728
R1339 VPB.n775 VPB.n774 6.728
R1340 VPB.n846 VPB.n845 6.728
R1341 VPB.n851 VPB.n850 6.728
R1342 VPB.n855 VPB.n854 6.728
R1343 VPB.n858 VPB.n857 6.728
R1344 VPB.n112 VPB.n111 6.728
R1345 VPB.n117 VPB.n116 6.728
R1346 VPB.n121 VPB.n120 6.728
R1347 VPB.n124 VPB.n123 6.728
R1348 VPB.n89 VPB.n88 6.728
R1349 VPB.n94 VPB.n93 6.728
R1350 VPB.n98 VPB.n97 6.728
R1351 VPB.n101 VPB.n100 6.728
R1352 VPB.n1006 VPB.n1005 6.728
R1353 VPB.n1011 VPB.n1010 6.728
R1354 VPB.n1015 VPB.n1014 6.728
R1355 VPB.n1018 VPB.n1017 6.728
R1356 VPB.n1089 VPB.n1088 6.728
R1357 VPB.n1094 VPB.n1093 6.728
R1358 VPB.n1098 VPB.n1097 6.728
R1359 VPB.n1101 VPB.n1100 6.728
R1360 VPB.n1172 VPB.n1171 6.728
R1361 VPB.n1177 VPB.n1176 6.728
R1362 VPB.n1181 VPB.n1180 6.728
R1363 VPB.n1184 VPB.n1183 6.728
R1364 VPB.n1255 VPB.n1254 6.728
R1365 VPB.n1260 VPB.n1259 6.728
R1366 VPB.n1264 VPB.n1263 6.728
R1367 VPB.n1267 VPB.n1266 6.728
R1368 VPB.n1338 VPB.n1337 6.728
R1369 VPB.n1343 VPB.n1342 6.728
R1370 VPB.n1347 VPB.n1346 6.728
R1371 VPB.n1350 VPB.n1349 6.728
R1372 VPB.n1421 VPB.n1420 6.728
R1373 VPB.n1426 VPB.n1425 6.728
R1374 VPB.n1430 VPB.n1429 6.728
R1375 VPB.n1433 VPB.n1432 6.728
R1376 VPB.n1504 VPB.n1503 6.728
R1377 VPB.n1509 VPB.n1508 6.728
R1378 VPB.n1513 VPB.n1512 6.728
R1379 VPB.n1516 VPB.n1515 6.728
R1380 VPB.n1587 VPB.n1586 6.728
R1381 VPB.n1592 VPB.n1591 6.728
R1382 VPB.n1596 VPB.n1595 6.728
R1383 VPB.n1599 VPB.n1598 6.728
R1384 VPB.n23 VPB.n22 6.728
R1385 VPB.n28 VPB.n27 6.728
R1386 VPB.n32 VPB.n31 6.728
R1387 VPB.n35 VPB.n34 6.728
R1388 VPB.n4 VPB.n3 6.728
R1389 VPB.n9 VPB.n8 6.728
R1390 VPB.n13 VPB.n12 6.728
R1391 VPB.n1681 VPB.n1680 6.728
R1392 VPB.n320 VPB.n316 6.458
R1393 VPB.n190 VPB.n189 6.398
R1394 VPB.n204 VPB.n194 6.112
R1395 VPB.n204 VPB.n203 6.101
R1396 VPB.n404 VPB.n400 4.305
R1397 VPB.n487 VPB.n483 4.305
R1398 VPB.n570 VPB.n566 4.305
R1399 VPB.n653 VPB.n649 4.305
R1400 VPB.n736 VPB.n732 4.305
R1401 VPB.n819 VPB.n815 4.305
R1402 VPB.n902 VPB.n898 4.305
R1403 VPB.n159 VPB.n155 4.305
R1404 VPB.n979 VPB.n975 4.305
R1405 VPB.n1062 VPB.n1058 4.305
R1406 VPB.n1145 VPB.n1141 4.305
R1407 VPB.n1228 VPB.n1224 4.305
R1408 VPB.n1311 VPB.n1307 4.305
R1409 VPB.n1394 VPB.n1390 4.305
R1410 VPB.n1477 VPB.n1473 4.305
R1411 VPB.n1560 VPB.n1556 4.305
R1412 VPB.n1643 VPB.n1639 4.305
R1413 VPB.n70 VPB.n66 4.305
R1414 VPB.n387 VPB.n383 3.947
R1415 VPB.n470 VPB.n466 3.947
R1416 VPB.n553 VPB.n549 3.947
R1417 VPB.n636 VPB.n632 3.947
R1418 VPB.n719 VPB.n715 3.947
R1419 VPB.n802 VPB.n798 3.947
R1420 VPB.n885 VPB.n881 3.947
R1421 VPB.n146 VPB.n145 3.947
R1422 VPB.n962 VPB.n958 3.947
R1423 VPB.n1045 VPB.n1041 3.947
R1424 VPB.n1128 VPB.n1124 3.947
R1425 VPB.n1211 VPB.n1207 3.947
R1426 VPB.n1294 VPB.n1290 3.947
R1427 VPB.n1377 VPB.n1373 3.947
R1428 VPB.n1460 VPB.n1456 3.947
R1429 VPB.n1543 VPB.n1539 3.947
R1430 VPB.n1626 VPB.n1622 3.947
R1431 VPB.n57 VPB.n56 3.947
R1432 VPB.n335 VPB.n332 1.794
R1433 VPB.n308 VPB.n305 1.435
R1434 VPB.n188 VPB.n181 1.402
R1435 VPB.n188 VPB.n184 1.402
R1436 VPB.n188 VPB.n186 1.402
R1437 VPB.n188 VPB.n187 1.402
R1438 VPB.n375 VPB.n372 1.076
R1439 VPB.n458 VPB.n455 1.076
R1440 VPB.n541 VPB.n538 1.076
R1441 VPB.n624 VPB.n621 1.076
R1442 VPB.n707 VPB.n704 1.076
R1443 VPB.n790 VPB.n787 1.076
R1444 VPB.n873 VPB.n870 1.076
R1445 VPB.n137 VPB.n134 1.076
R1446 VPB.n950 VPB.n947 1.076
R1447 VPB.n1033 VPB.n1030 1.076
R1448 VPB.n1116 VPB.n1113 1.076
R1449 VPB.n1199 VPB.n1196 1.076
R1450 VPB.n1282 VPB.n1279 1.076
R1451 VPB.n1365 VPB.n1362 1.076
R1452 VPB.n1448 VPB.n1445 1.076
R1453 VPB.n1531 VPB.n1528 1.076
R1454 VPB.n1614 VPB.n1611 1.076
R1455 VPB.n48 VPB.n45 1.076
R1456 VPB.n189 VPB.n188 0.735
R1457 VPB.n188 VPB.n178 0.735
R1458 VPB.n414 VPB.n411 0.717
R1459 VPB.n497 VPB.n494 0.717
R1460 VPB.n580 VPB.n577 0.717
R1461 VPB.n663 VPB.n660 0.717
R1462 VPB.n746 VPB.n743 0.717
R1463 VPB.n829 VPB.n826 0.717
R1464 VPB.n912 VPB.n909 0.717
R1465 VPB.n167 VPB.n166 0.717
R1466 VPB.n989 VPB.n986 0.717
R1467 VPB.n1072 VPB.n1069 0.717
R1468 VPB.n1155 VPB.n1152 0.717
R1469 VPB.n1238 VPB.n1235 0.717
R1470 VPB.n1321 VPB.n1318 0.717
R1471 VPB.n1404 VPB.n1401 0.717
R1472 VPB.n1487 VPB.n1484 0.717
R1473 VPB.n1570 VPB.n1567 0.717
R1474 VPB.n1653 VPB.n1650 0.717
R1475 VPB.n78 VPB.n77 0.717
R1476 VPB.n240 VPB.n239 0.387
R1477 VPB.n240 VPB.n235 0.387
R1478 VPB.n240 VPB.n230 0.387
R1479 VPB.n241 VPB.n240 0.387
R1480 VPB.n295 VPB.n294 0.387
R1481 VPB.n295 VPB.n290 0.387
R1482 VPB.n295 VPB.n285 0.387
R1483 VPB.n296 VPB.n295 0.387
R1484 VPB.n358 VPB.n357 0.387
R1485 VPB.n358 VPB.n353 0.387
R1486 VPB.n358 VPB.n348 0.387
R1487 VPB.n359 VPB.n358 0.387
R1488 VPB.n441 VPB.n440 0.387
R1489 VPB.n441 VPB.n436 0.387
R1490 VPB.n441 VPB.n431 0.387
R1491 VPB.n442 VPB.n441 0.387
R1492 VPB.n524 VPB.n523 0.387
R1493 VPB.n524 VPB.n519 0.387
R1494 VPB.n524 VPB.n514 0.387
R1495 VPB.n525 VPB.n524 0.387
R1496 VPB.n607 VPB.n606 0.387
R1497 VPB.n607 VPB.n602 0.387
R1498 VPB.n607 VPB.n597 0.387
R1499 VPB.n608 VPB.n607 0.387
R1500 VPB.n690 VPB.n689 0.387
R1501 VPB.n690 VPB.n685 0.387
R1502 VPB.n690 VPB.n680 0.387
R1503 VPB.n691 VPB.n690 0.387
R1504 VPB.n773 VPB.n772 0.387
R1505 VPB.n773 VPB.n768 0.387
R1506 VPB.n773 VPB.n763 0.387
R1507 VPB.n774 VPB.n773 0.387
R1508 VPB.n856 VPB.n855 0.387
R1509 VPB.n856 VPB.n851 0.387
R1510 VPB.n856 VPB.n846 0.387
R1511 VPB.n857 VPB.n856 0.387
R1512 VPB.n122 VPB.n121 0.387
R1513 VPB.n122 VPB.n117 0.387
R1514 VPB.n122 VPB.n112 0.387
R1515 VPB.n123 VPB.n122 0.387
R1516 VPB.n99 VPB.n98 0.387
R1517 VPB.n99 VPB.n94 0.387
R1518 VPB.n99 VPB.n89 0.387
R1519 VPB.n100 VPB.n99 0.387
R1520 VPB.n1016 VPB.n1015 0.387
R1521 VPB.n1016 VPB.n1011 0.387
R1522 VPB.n1016 VPB.n1006 0.387
R1523 VPB.n1017 VPB.n1016 0.387
R1524 VPB.n1099 VPB.n1098 0.387
R1525 VPB.n1099 VPB.n1094 0.387
R1526 VPB.n1099 VPB.n1089 0.387
R1527 VPB.n1100 VPB.n1099 0.387
R1528 VPB.n1182 VPB.n1181 0.387
R1529 VPB.n1182 VPB.n1177 0.387
R1530 VPB.n1182 VPB.n1172 0.387
R1531 VPB.n1183 VPB.n1182 0.387
R1532 VPB.n1265 VPB.n1264 0.387
R1533 VPB.n1265 VPB.n1260 0.387
R1534 VPB.n1265 VPB.n1255 0.387
R1535 VPB.n1266 VPB.n1265 0.387
R1536 VPB.n1348 VPB.n1347 0.387
R1537 VPB.n1348 VPB.n1343 0.387
R1538 VPB.n1348 VPB.n1338 0.387
R1539 VPB.n1349 VPB.n1348 0.387
R1540 VPB.n1431 VPB.n1430 0.387
R1541 VPB.n1431 VPB.n1426 0.387
R1542 VPB.n1431 VPB.n1421 0.387
R1543 VPB.n1432 VPB.n1431 0.387
R1544 VPB.n1514 VPB.n1513 0.387
R1545 VPB.n1514 VPB.n1509 0.387
R1546 VPB.n1514 VPB.n1504 0.387
R1547 VPB.n1515 VPB.n1514 0.387
R1548 VPB.n1597 VPB.n1596 0.387
R1549 VPB.n1597 VPB.n1592 0.387
R1550 VPB.n1597 VPB.n1587 0.387
R1551 VPB.n1598 VPB.n1597 0.387
R1552 VPB.n33 VPB.n32 0.387
R1553 VPB.n33 VPB.n28 0.387
R1554 VPB.n33 VPB.n23 0.387
R1555 VPB.n34 VPB.n33 0.387
R1556 VPB.n1682 VPB.n13 0.387
R1557 VPB.n1682 VPB.n9 0.387
R1558 VPB.n1682 VPB.n4 0.387
R1559 VPB.n1682 VPB.n1681 0.387
R1560 VPB.n249 VPB.n222 0.272
R1561 VPB.n304 VPB.n277 0.272
R1562 VPB.n367 VPB.n340 0.272
R1563 VPB.n450 VPB.n423 0.272
R1564 VPB.n533 VPB.n506 0.272
R1565 VPB.n616 VPB.n589 0.272
R1566 VPB.n699 VPB.n672 0.272
R1567 VPB.n782 VPB.n755 0.272
R1568 VPB.n865 VPB.n838 0.272
R1569 VPB.n922 VPB.n921 0.272
R1570 VPB.n1025 VPB.n998 0.272
R1571 VPB.n1108 VPB.n1081 0.272
R1572 VPB.n1191 VPB.n1164 0.272
R1573 VPB.n1274 VPB.n1247 0.272
R1574 VPB.n1357 VPB.n1330 0.272
R1575 VPB.n1440 VPB.n1413 0.272
R1576 VPB.n1523 VPB.n1496 0.272
R1577 VPB.n1606 VPB.n1579 0.272
R1578 VPB.n1663 VPB.n1662 0.272
R1579 VPB.n942 VPB 0.204
R1580 VPB.n1674 VPB 0.198
R1581 VPB.n206 VPB.n205 0.136
R1582 VPB.n210 VPB.n206 0.136
R1583 VPB.n214 VPB.n210 0.136
R1584 VPB.n218 VPB.n214 0.136
R1585 VPB.n222 VPB.n218 0.136
R1586 VPB.n253 VPB.n249 0.136
R1587 VPB.n257 VPB.n253 0.136
R1588 VPB.n261 VPB.n257 0.136
R1589 VPB.n265 VPB.n261 0.136
R1590 VPB.n269 VPB.n265 0.136
R1591 VPB.n273 VPB.n269 0.136
R1592 VPB.n277 VPB.n273 0.136
R1593 VPB.n309 VPB.n304 0.136
R1594 VPB.n314 VPB.n309 0.136
R1595 VPB.n321 VPB.n314 0.136
R1596 VPB.n326 VPB.n321 0.136
R1597 VPB.n331 VPB.n326 0.136
R1598 VPB.n336 VPB.n331 0.136
R1599 VPB.n340 VPB.n336 0.136
R1600 VPB.n371 VPB.n367 0.136
R1601 VPB.n376 VPB.n371 0.136
R1602 VPB.n381 VPB.n376 0.136
R1603 VPB.n388 VPB.n381 0.136
R1604 VPB.n393 VPB.n388 0.136
R1605 VPB.n398 VPB.n393 0.136
R1606 VPB.n405 VPB.n398 0.136
R1607 VPB.n410 VPB.n405 0.136
R1608 VPB.n415 VPB.n410 0.136
R1609 VPB.n419 VPB.n415 0.136
R1610 VPB.n423 VPB.n419 0.136
R1611 VPB.n454 VPB.n450 0.136
R1612 VPB.n459 VPB.n454 0.136
R1613 VPB.n464 VPB.n459 0.136
R1614 VPB.n471 VPB.n464 0.136
R1615 VPB.n476 VPB.n471 0.136
R1616 VPB.n481 VPB.n476 0.136
R1617 VPB.n488 VPB.n481 0.136
R1618 VPB.n493 VPB.n488 0.136
R1619 VPB.n498 VPB.n493 0.136
R1620 VPB.n502 VPB.n498 0.136
R1621 VPB.n506 VPB.n502 0.136
R1622 VPB.n537 VPB.n533 0.136
R1623 VPB.n542 VPB.n537 0.136
R1624 VPB.n547 VPB.n542 0.136
R1625 VPB.n554 VPB.n547 0.136
R1626 VPB.n559 VPB.n554 0.136
R1627 VPB.n564 VPB.n559 0.136
R1628 VPB.n571 VPB.n564 0.136
R1629 VPB.n576 VPB.n571 0.136
R1630 VPB.n581 VPB.n576 0.136
R1631 VPB.n585 VPB.n581 0.136
R1632 VPB.n589 VPB.n585 0.136
R1633 VPB.n620 VPB.n616 0.136
R1634 VPB.n625 VPB.n620 0.136
R1635 VPB.n630 VPB.n625 0.136
R1636 VPB.n637 VPB.n630 0.136
R1637 VPB.n642 VPB.n637 0.136
R1638 VPB.n647 VPB.n642 0.136
R1639 VPB.n654 VPB.n647 0.136
R1640 VPB.n659 VPB.n654 0.136
R1641 VPB.n664 VPB.n659 0.136
R1642 VPB.n668 VPB.n664 0.136
R1643 VPB.n672 VPB.n668 0.136
R1644 VPB.n703 VPB.n699 0.136
R1645 VPB.n708 VPB.n703 0.136
R1646 VPB.n713 VPB.n708 0.136
R1647 VPB.n720 VPB.n713 0.136
R1648 VPB.n725 VPB.n720 0.136
R1649 VPB.n730 VPB.n725 0.136
R1650 VPB.n737 VPB.n730 0.136
R1651 VPB.n742 VPB.n737 0.136
R1652 VPB.n747 VPB.n742 0.136
R1653 VPB.n751 VPB.n747 0.136
R1654 VPB.n755 VPB.n751 0.136
R1655 VPB.n786 VPB.n782 0.136
R1656 VPB.n791 VPB.n786 0.136
R1657 VPB.n796 VPB.n791 0.136
R1658 VPB.n803 VPB.n796 0.136
R1659 VPB.n808 VPB.n803 0.136
R1660 VPB.n813 VPB.n808 0.136
R1661 VPB.n820 VPB.n813 0.136
R1662 VPB.n825 VPB.n820 0.136
R1663 VPB.n830 VPB.n825 0.136
R1664 VPB.n834 VPB.n830 0.136
R1665 VPB.n838 VPB.n834 0.136
R1666 VPB.n869 VPB.n865 0.136
R1667 VPB.n874 VPB.n869 0.136
R1668 VPB.n879 VPB.n874 0.136
R1669 VPB.n886 VPB.n879 0.136
R1670 VPB.n891 VPB.n886 0.136
R1671 VPB.n896 VPB.n891 0.136
R1672 VPB.n903 VPB.n896 0.136
R1673 VPB.n908 VPB.n903 0.136
R1674 VPB.n913 VPB.n908 0.136
R1675 VPB.n917 VPB.n913 0.136
R1676 VPB.n921 VPB.n917 0.136
R1677 VPB.n923 VPB.n922 0.136
R1678 VPB.n924 VPB.n923 0.136
R1679 VPB.n925 VPB.n924 0.136
R1680 VPB.n926 VPB.n925 0.136
R1681 VPB.n927 VPB.n926 0.136
R1682 VPB.n928 VPB.n927 0.136
R1683 VPB.n929 VPB.n928 0.136
R1684 VPB.n930 VPB.n929 0.136
R1685 VPB.n931 VPB.n930 0.136
R1686 VPB.n932 VPB.n931 0.136
R1687 VPB.n933 VPB.n932 0.136
R1688 VPB.n946 VPB.n942 0.136
R1689 VPB.n951 VPB.n946 0.136
R1690 VPB.n956 VPB.n951 0.136
R1691 VPB.n963 VPB.n956 0.136
R1692 VPB.n968 VPB.n963 0.136
R1693 VPB.n973 VPB.n968 0.136
R1694 VPB.n980 VPB.n973 0.136
R1695 VPB.n985 VPB.n980 0.136
R1696 VPB.n990 VPB.n985 0.136
R1697 VPB.n994 VPB.n990 0.136
R1698 VPB.n998 VPB.n994 0.136
R1699 VPB.n1029 VPB.n1025 0.136
R1700 VPB.n1034 VPB.n1029 0.136
R1701 VPB.n1039 VPB.n1034 0.136
R1702 VPB.n1046 VPB.n1039 0.136
R1703 VPB.n1051 VPB.n1046 0.136
R1704 VPB.n1056 VPB.n1051 0.136
R1705 VPB.n1063 VPB.n1056 0.136
R1706 VPB.n1068 VPB.n1063 0.136
R1707 VPB.n1073 VPB.n1068 0.136
R1708 VPB.n1077 VPB.n1073 0.136
R1709 VPB.n1081 VPB.n1077 0.136
R1710 VPB.n1112 VPB.n1108 0.136
R1711 VPB.n1117 VPB.n1112 0.136
R1712 VPB.n1122 VPB.n1117 0.136
R1713 VPB.n1129 VPB.n1122 0.136
R1714 VPB.n1134 VPB.n1129 0.136
R1715 VPB.n1139 VPB.n1134 0.136
R1716 VPB.n1146 VPB.n1139 0.136
R1717 VPB.n1151 VPB.n1146 0.136
R1718 VPB.n1156 VPB.n1151 0.136
R1719 VPB.n1160 VPB.n1156 0.136
R1720 VPB.n1164 VPB.n1160 0.136
R1721 VPB.n1195 VPB.n1191 0.136
R1722 VPB.n1200 VPB.n1195 0.136
R1723 VPB.n1205 VPB.n1200 0.136
R1724 VPB.n1212 VPB.n1205 0.136
R1725 VPB.n1217 VPB.n1212 0.136
R1726 VPB.n1222 VPB.n1217 0.136
R1727 VPB.n1229 VPB.n1222 0.136
R1728 VPB.n1234 VPB.n1229 0.136
R1729 VPB.n1239 VPB.n1234 0.136
R1730 VPB.n1243 VPB.n1239 0.136
R1731 VPB.n1247 VPB.n1243 0.136
R1732 VPB.n1278 VPB.n1274 0.136
R1733 VPB.n1283 VPB.n1278 0.136
R1734 VPB.n1288 VPB.n1283 0.136
R1735 VPB.n1295 VPB.n1288 0.136
R1736 VPB.n1300 VPB.n1295 0.136
R1737 VPB.n1305 VPB.n1300 0.136
R1738 VPB.n1312 VPB.n1305 0.136
R1739 VPB.n1317 VPB.n1312 0.136
R1740 VPB.n1322 VPB.n1317 0.136
R1741 VPB.n1326 VPB.n1322 0.136
R1742 VPB.n1330 VPB.n1326 0.136
R1743 VPB.n1361 VPB.n1357 0.136
R1744 VPB.n1366 VPB.n1361 0.136
R1745 VPB.n1371 VPB.n1366 0.136
R1746 VPB.n1378 VPB.n1371 0.136
R1747 VPB.n1383 VPB.n1378 0.136
R1748 VPB.n1388 VPB.n1383 0.136
R1749 VPB.n1395 VPB.n1388 0.136
R1750 VPB.n1400 VPB.n1395 0.136
R1751 VPB.n1405 VPB.n1400 0.136
R1752 VPB.n1409 VPB.n1405 0.136
R1753 VPB.n1413 VPB.n1409 0.136
R1754 VPB.n1444 VPB.n1440 0.136
R1755 VPB.n1449 VPB.n1444 0.136
R1756 VPB.n1454 VPB.n1449 0.136
R1757 VPB.n1461 VPB.n1454 0.136
R1758 VPB.n1466 VPB.n1461 0.136
R1759 VPB.n1471 VPB.n1466 0.136
R1760 VPB.n1478 VPB.n1471 0.136
R1761 VPB.n1483 VPB.n1478 0.136
R1762 VPB.n1488 VPB.n1483 0.136
R1763 VPB.n1492 VPB.n1488 0.136
R1764 VPB.n1496 VPB.n1492 0.136
R1765 VPB.n1527 VPB.n1523 0.136
R1766 VPB.n1532 VPB.n1527 0.136
R1767 VPB.n1537 VPB.n1532 0.136
R1768 VPB.n1544 VPB.n1537 0.136
R1769 VPB.n1549 VPB.n1544 0.136
R1770 VPB.n1554 VPB.n1549 0.136
R1771 VPB.n1561 VPB.n1554 0.136
R1772 VPB.n1566 VPB.n1561 0.136
R1773 VPB.n1571 VPB.n1566 0.136
R1774 VPB.n1575 VPB.n1571 0.136
R1775 VPB.n1579 VPB.n1575 0.136
R1776 VPB.n1610 VPB.n1606 0.136
R1777 VPB.n1615 VPB.n1610 0.136
R1778 VPB.n1620 VPB.n1615 0.136
R1779 VPB.n1627 VPB.n1620 0.136
R1780 VPB.n1632 VPB.n1627 0.136
R1781 VPB.n1637 VPB.n1632 0.136
R1782 VPB.n1644 VPB.n1637 0.136
R1783 VPB.n1649 VPB.n1644 0.136
R1784 VPB.n1654 VPB.n1649 0.136
R1785 VPB.n1658 VPB.n1654 0.136
R1786 VPB.n1662 VPB.n1658 0.136
R1787 VPB.n1664 VPB.n1663 0.136
R1788 VPB.n1665 VPB.n1664 0.136
R1789 VPB.n1666 VPB.n1665 0.136
R1790 VPB.n1667 VPB.n1666 0.136
R1791 VPB.n1668 VPB.n1667 0.136
R1792 VPB.n1669 VPB.n1668 0.136
R1793 VPB.n1670 VPB.n1669 0.136
R1794 VPB.n1671 VPB.n1670 0.136
R1795 VPB.n1672 VPB.n1671 0.136
R1796 VPB.n1673 VPB.n1672 0.136
R1797 VPB.n1674 VPB.n1673 0.136
R1798 VPB.n933 VPB 0.068
R1799 a_4447_943.n5 a_4447_943.t8 454.685
R1800 a_4447_943.n5 a_4447_943.t9 428.979
R1801 a_4447_943.n6 a_4447_943.t7 221.453
R1802 a_4447_943.n9 a_4447_943.n7 203.12
R1803 a_4447_943.n7 a_4447_943.n4 180.846
R1804 a_4447_943.n7 a_4447_943.n6 156.035
R1805 a_4447_943.n6 a_4447_943.n5 108.494
R1806 a_4447_943.n3 a_4447_943.n2 79.232
R1807 a_4447_943.n4 a_4447_943.n3 63.152
R1808 a_4447_943.n4 a_4447_943.n0 16.08
R1809 a_4447_943.n3 a_4447_943.n1 16.08
R1810 a_4447_943.n9 a_4447_943.n8 15.218
R1811 a_4447_943.n0 a_4447_943.t6 14.282
R1812 a_4447_943.n0 a_4447_943.t2 14.282
R1813 a_4447_943.n1 a_4447_943.t4 14.282
R1814 a_4447_943.n1 a_4447_943.t5 14.282
R1815 a_4447_943.n2 a_4447_943.t3 14.282
R1816 a_4447_943.n2 a_4447_943.t1 14.282
R1817 a_4447_943.n10 a_4447_943.n9 12.014
R1818 a_6371_943.n5 a_6371_943.t11 512.525
R1819 a_6371_943.n7 a_6371_943.t12 454.685
R1820 a_6371_943.n7 a_6371_943.t8 428.979
R1821 a_6371_943.n5 a_6371_943.t7 371.139
R1822 a_6371_943.n6 a_6371_943.t10 271.162
R1823 a_6371_943.n8 a_6371_943.t9 221.453
R1824 a_6371_943.n12 a_6371_943.n10 203.12
R1825 a_6371_943.n10 a_6371_943.n4 180.846
R1826 a_6371_943.n6 a_6371_943.n5 172.76
R1827 a_6371_943.n8 a_6371_943.n7 108.494
R1828 a_6371_943.n9 a_6371_943.n6 84.388
R1829 a_6371_943.n9 a_6371_943.n8 80.035
R1830 a_6371_943.n3 a_6371_943.n2 79.232
R1831 a_6371_943.n10 a_6371_943.n9 76
R1832 a_6371_943.n4 a_6371_943.n3 63.152
R1833 a_6371_943.n4 a_6371_943.n0 16.08
R1834 a_6371_943.n3 a_6371_943.n1 16.08
R1835 a_6371_943.n12 a_6371_943.n11 15.218
R1836 a_6371_943.n0 a_6371_943.t6 14.282
R1837 a_6371_943.n0 a_6371_943.t0 14.282
R1838 a_6371_943.n1 a_6371_943.t5 14.282
R1839 a_6371_943.n1 a_6371_943.t4 14.282
R1840 a_6371_943.n2 a_6371_943.t2 14.282
R1841 a_6371_943.n2 a_6371_943.t3 14.282
R1842 a_6371_943.n13 a_6371_943.n12 12.014
R1843 a_7333_943.n8 a_7333_943.t10 454.685
R1844 a_7333_943.n10 a_7333_943.t13 454.685
R1845 a_7333_943.n6 a_7333_943.t12 454.685
R1846 a_7333_943.n8 a_7333_943.t15 428.979
R1847 a_7333_943.n10 a_7333_943.t7 428.979
R1848 a_7333_943.n6 a_7333_943.t14 428.979
R1849 a_7333_943.n9 a_7333_943.t9 248.006
R1850 a_7333_943.n11 a_7333_943.t8 248.006
R1851 a_7333_943.n7 a_7333_943.t11 248.006
R1852 a_7333_943.n16 a_7333_943.n14 223.151
R1853 a_7333_943.n14 a_7333_943.n5 154.293
R1854 a_7333_943.n13 a_7333_943.n7 82.484
R1855 a_7333_943.n9 a_7333_943.n8 81.941
R1856 a_7333_943.n11 a_7333_943.n10 81.941
R1857 a_7333_943.n7 a_7333_943.n6 81.941
R1858 a_7333_943.n12 a_7333_943.n11 79.491
R1859 a_7333_943.n4 a_7333_943.n3 79.232
R1860 a_7333_943.n12 a_7333_943.n9 76
R1861 a_7333_943.n14 a_7333_943.n13 76
R1862 a_7333_943.n5 a_7333_943.n4 63.152
R1863 a_7333_943.n16 a_7333_943.n15 30
R1864 a_7333_943.n17 a_7333_943.n0 24.383
R1865 a_7333_943.n17 a_7333_943.n16 23.684
R1866 a_7333_943.n5 a_7333_943.n1 16.08
R1867 a_7333_943.n4 a_7333_943.n2 16.08
R1868 a_7333_943.n1 a_7333_943.t4 14.282
R1869 a_7333_943.n1 a_7333_943.t5 14.282
R1870 a_7333_943.n2 a_7333_943.t2 14.282
R1871 a_7333_943.n2 a_7333_943.t3 14.282
R1872 a_7333_943.n3 a_7333_943.t1 14.282
R1873 a_7333_943.n3 a_7333_943.t0 14.282
R1874 a_7333_943.n13 a_7333_943.n12 4.035
R1875 a_12143_943.n6 a_12143_943.t12 512.525
R1876 a_12143_943.n8 a_12143_943.t8 454.685
R1877 a_12143_943.n8 a_12143_943.t11 428.979
R1878 a_12143_943.n6 a_12143_943.t10 371.139
R1879 a_12143_943.n7 a_12143_943.t7 271.162
R1880 a_12143_943.n9 a_12143_943.t9 221.453
R1881 a_12143_943.n13 a_12143_943.n11 196.598
R1882 a_12143_943.n11 a_12143_943.n5 180.846
R1883 a_12143_943.n7 a_12143_943.n6 172.76
R1884 a_12143_943.n9 a_12143_943.n8 108.494
R1885 a_12143_943.n10 a_12143_943.n7 84.388
R1886 a_12143_943.n10 a_12143_943.n9 80.035
R1887 a_12143_943.n4 a_12143_943.n3 79.232
R1888 a_12143_943.n11 a_12143_943.n10 76
R1889 a_12143_943.n5 a_12143_943.n4 63.152
R1890 a_12143_943.n13 a_12143_943.n12 30
R1891 a_12143_943.n14 a_12143_943.n0 24.383
R1892 a_12143_943.n14 a_12143_943.n13 23.684
R1893 a_12143_943.n5 a_12143_943.n1 16.08
R1894 a_12143_943.n4 a_12143_943.n2 16.08
R1895 a_12143_943.n1 a_12143_943.t1 14.282
R1896 a_12143_943.n1 a_12143_943.t2 14.282
R1897 a_12143_943.n2 a_12143_943.t4 14.282
R1898 a_12143_943.n2 a_12143_943.t3 14.282
R1899 a_12143_943.n3 a_12143_943.t5 14.282
R1900 a_12143_943.n3 a_12143_943.t6 14.282
R1901 a_15483_75.t0 a_15483_75.n0 117.777
R1902 a_15483_75.n2 a_15483_75.n1 55.228
R1903 a_15483_75.n4 a_15483_75.n3 9.111
R1904 a_15483_75.n8 a_15483_75.n6 7.859
R1905 a_15483_75.t0 a_15483_75.n2 4.04
R1906 a_15483_75.t0 a_15483_75.n8 3.034
R1907 a_15483_75.n6 a_15483_75.n4 1.964
R1908 a_15483_75.n6 a_15483_75.n5 1.964
R1909 a_15483_75.n8 a_15483_75.n7 0.443
R1910 VNB VNB.n1425 300.778
R1911 VNB.n198 VNB.n197 199.897
R1912 VNB.n250 VNB.n249 199.897
R1913 VNB.n302 VNB.n301 199.897
R1914 VNB.n370 VNB.n369 199.897
R1915 VNB.n438 VNB.n437 199.897
R1916 VNB.n513 VNB.n512 199.897
R1917 VNB.n581 VNB.n580 199.897
R1918 VNB.n649 VNB.n648 199.897
R1919 VNB.n724 VNB.n723 199.897
R1920 VNB.n94 VNB.n93 199.897
R1921 VNB.n74 VNB.n73 199.897
R1922 VNB.n859 VNB.n858 199.897
R1923 VNB.n927 VNB.n926 199.897
R1924 VNB.n995 VNB.n994 199.897
R1925 VNB.n1070 VNB.n1069 199.897
R1926 VNB.n1138 VNB.n1137 199.897
R1927 VNB.n1206 VNB.n1205 199.897
R1928 VNB.n1274 VNB.n1273 199.897
R1929 VNB.n1342 VNB.n1341 199.897
R1930 VNB.n18 VNB.n17 199.897
R1931 VNB.n207 VNB.n205 154.509
R1932 VNB.n311 VNB.n309 154.509
R1933 VNB.n259 VNB.n257 154.509
R1934 VNB.n447 VNB.n445 154.509
R1935 VNB.n379 VNB.n377 154.509
R1936 VNB.n590 VNB.n588 154.509
R1937 VNB.n522 VNB.n520 154.509
R1938 VNB.n733 VNB.n731 154.509
R1939 VNB.n658 VNB.n656 154.509
R1940 VNB.n800 VNB.n798 154.509
R1941 VNB.n103 VNB.n101 154.509
R1942 VNB.n936 VNB.n934 154.509
R1943 VNB.n868 VNB.n866 154.509
R1944 VNB.n1079 VNB.n1077 154.509
R1945 VNB.n1004 VNB.n1002 154.509
R1946 VNB.n1215 VNB.n1213 154.509
R1947 VNB.n1147 VNB.n1145 154.509
R1948 VNB.n1351 VNB.n1349 154.509
R1949 VNB.n1283 VNB.n1281 154.509
R1950 VNB.n27 VNB.n25 154.509
R1951 VNB.n479 VNB.n478 147.75
R1952 VNB.n690 VNB.n689 147.75
R1953 VNB.n127 VNB.n126 147.75
R1954 VNB.n1036 VNB.n1035 147.75
R1955 VNB.n51 VNB.n50 147.75
R1956 VNB.n491 VNB.n488 121.366
R1957 VNB.n702 VNB.n699 121.366
R1958 VNB.n132 VNB.n130 121.366
R1959 VNB.n1048 VNB.n1045 121.366
R1960 VNB.n56 VNB.n54 121.366
R1961 VNB.n347 VNB.n346 85.559
R1962 VNB.n415 VNB.n414 85.559
R1963 VNB.n558 VNB.n557 85.559
R1964 VNB.n626 VNB.n625 85.559
R1965 VNB.n769 VNB.n768 85.559
R1966 VNB.n836 VNB.n835 85.559
R1967 VNB.n904 VNB.n903 85.559
R1968 VNB.n972 VNB.n971 85.559
R1969 VNB.n1115 VNB.n1114 85.559
R1970 VNB.n1183 VNB.n1182 85.559
R1971 VNB.n1251 VNB.n1250 85.559
R1972 VNB.n1319 VNB.n1318 85.559
R1973 VNB.n1387 VNB.n1386 85.559
R1974 VNB.n175 VNB.n174 84.842
R1975 VNB.n227 VNB.n226 84.842
R1976 VNB.n279 VNB.n278 84.842
R1977 VNB.n1412 VNB.n1411 76
R1978 VNB.n1399 VNB.n1398 76
R1979 VNB.n1395 VNB.n1394 76
R1980 VNB.n1391 VNB.n1390 76
R1981 VNB.n1385 VNB.n1384 76
R1982 VNB.n1381 VNB.n1380 76
R1983 VNB.n1377 VNB.n1376 76
R1984 VNB.n1373 VNB.n1372 76
R1985 VNB.n1369 VNB.n1368 76
R1986 VNB.n1365 VNB.n1364 76
R1987 VNB.n1361 VNB.n1360 76
R1988 VNB.n1357 VNB.n1356 76
R1989 VNB.n1353 VNB.n1352 76
R1990 VNB.n1331 VNB.n1330 76
R1991 VNB.n1327 VNB.n1326 76
R1992 VNB.n1323 VNB.n1322 76
R1993 VNB.n1317 VNB.n1316 76
R1994 VNB.n1313 VNB.n1312 76
R1995 VNB.n1309 VNB.n1308 76
R1996 VNB.n1305 VNB.n1304 76
R1997 VNB.n1301 VNB.n1300 76
R1998 VNB.n1297 VNB.n1296 76
R1999 VNB.n1293 VNB.n1292 76
R2000 VNB.n1289 VNB.n1288 76
R2001 VNB.n1285 VNB.n1284 76
R2002 VNB.n1263 VNB.n1262 76
R2003 VNB.n1259 VNB.n1258 76
R2004 VNB.n1255 VNB.n1254 76
R2005 VNB.n1249 VNB.n1248 76
R2006 VNB.n1245 VNB.n1244 76
R2007 VNB.n1241 VNB.n1240 76
R2008 VNB.n1237 VNB.n1236 76
R2009 VNB.n1233 VNB.n1232 76
R2010 VNB.n1229 VNB.n1228 76
R2011 VNB.n1225 VNB.n1224 76
R2012 VNB.n1221 VNB.n1220 76
R2013 VNB.n1217 VNB.n1216 76
R2014 VNB.n1195 VNB.n1194 76
R2015 VNB.n1191 VNB.n1190 76
R2016 VNB.n1187 VNB.n1186 76
R2017 VNB.n1181 VNB.n1180 76
R2018 VNB.n1177 VNB.n1176 76
R2019 VNB.n1173 VNB.n1172 76
R2020 VNB.n1169 VNB.n1168 76
R2021 VNB.n1165 VNB.n1164 76
R2022 VNB.n1161 VNB.n1160 76
R2023 VNB.n1157 VNB.n1156 76
R2024 VNB.n1153 VNB.n1152 76
R2025 VNB.n1149 VNB.n1148 76
R2026 VNB.n1127 VNB.n1126 76
R2027 VNB.n1123 VNB.n1122 76
R2028 VNB.n1119 VNB.n1118 76
R2029 VNB.n1113 VNB.n1112 76
R2030 VNB.n1109 VNB.n1108 76
R2031 VNB.n1105 VNB.n1104 76
R2032 VNB.n1101 VNB.n1100 76
R2033 VNB.n1097 VNB.n1096 76
R2034 VNB.n1093 VNB.n1092 76
R2035 VNB.n1089 VNB.n1088 76
R2036 VNB.n1085 VNB.n1084 76
R2037 VNB.n1081 VNB.n1080 76
R2038 VNB.n1059 VNB.n1058 76
R2039 VNB.n1055 VNB.n1054 76
R2040 VNB.n1051 VNB.n1050 76
R2041 VNB.n1039 VNB.n1038 76
R2042 VNB.n1034 VNB.n1033 76
R2043 VNB.n1030 VNB.n1029 76
R2044 VNB.n1026 VNB.n1025 76
R2045 VNB.n1022 VNB.n1021 76
R2046 VNB.n1018 VNB.n1017 76
R2047 VNB.n1014 VNB.n1013 76
R2048 VNB.n1010 VNB.n1009 76
R2049 VNB.n1006 VNB.n1005 76
R2050 VNB.n984 VNB.n983 76
R2051 VNB.n980 VNB.n979 76
R2052 VNB.n976 VNB.n975 76
R2053 VNB.n970 VNB.n969 76
R2054 VNB.n966 VNB.n965 76
R2055 VNB.n962 VNB.n961 76
R2056 VNB.n958 VNB.n957 76
R2057 VNB.n954 VNB.n953 76
R2058 VNB.n950 VNB.n949 76
R2059 VNB.n946 VNB.n945 76
R2060 VNB.n942 VNB.n941 76
R2061 VNB.n938 VNB.n937 76
R2062 VNB.n916 VNB.n915 76
R2063 VNB.n912 VNB.n911 76
R2064 VNB.n908 VNB.n907 76
R2065 VNB.n902 VNB.n901 76
R2066 VNB.n898 VNB.n897 76
R2067 VNB.n894 VNB.n893 76
R2068 VNB.n890 VNB.n889 76
R2069 VNB.n886 VNB.n885 76
R2070 VNB.n882 VNB.n881 76
R2071 VNB.n878 VNB.n877 76
R2072 VNB.n874 VNB.n873 76
R2073 VNB.n870 VNB.n869 76
R2074 VNB.n848 VNB.n847 76
R2075 VNB.n844 VNB.n843 76
R2076 VNB.n840 VNB.n839 76
R2077 VNB.n834 VNB.n833 76
R2078 VNB.n830 VNB.n829 76
R2079 VNB.n826 VNB.n825 76
R2080 VNB.n822 VNB.n821 76
R2081 VNB.n818 VNB.n817 76
R2082 VNB.n814 VNB.n813 76
R2083 VNB.n810 VNB.n809 76
R2084 VNB.n806 VNB.n805 76
R2085 VNB.n802 VNB.n801 76
R2086 VNB.n796 VNB.n793 76
R2087 VNB.n781 VNB.n780 76
R2088 VNB.n777 VNB.n776 76
R2089 VNB.n773 VNB.n772 76
R2090 VNB.n767 VNB.n766 76
R2091 VNB.n763 VNB.n762 76
R2092 VNB.n759 VNB.n758 76
R2093 VNB.n755 VNB.n754 76
R2094 VNB.n751 VNB.n750 76
R2095 VNB.n747 VNB.n746 76
R2096 VNB.n743 VNB.n742 76
R2097 VNB.n739 VNB.n738 76
R2098 VNB.n735 VNB.n734 76
R2099 VNB.n713 VNB.n712 76
R2100 VNB.n709 VNB.n708 76
R2101 VNB.n705 VNB.n704 76
R2102 VNB.n693 VNB.n692 76
R2103 VNB.n688 VNB.n687 76
R2104 VNB.n684 VNB.n683 76
R2105 VNB.n680 VNB.n679 76
R2106 VNB.n676 VNB.n675 76
R2107 VNB.n672 VNB.n671 76
R2108 VNB.n668 VNB.n667 76
R2109 VNB.n664 VNB.n663 76
R2110 VNB.n660 VNB.n659 76
R2111 VNB.n638 VNB.n637 76
R2112 VNB.n634 VNB.n633 76
R2113 VNB.n630 VNB.n629 76
R2114 VNB.n624 VNB.n623 76
R2115 VNB.n620 VNB.n619 76
R2116 VNB.n616 VNB.n615 76
R2117 VNB.n612 VNB.n611 76
R2118 VNB.n608 VNB.n607 76
R2119 VNB.n604 VNB.n603 76
R2120 VNB.n600 VNB.n599 76
R2121 VNB.n596 VNB.n595 76
R2122 VNB.n592 VNB.n591 76
R2123 VNB.n570 VNB.n569 76
R2124 VNB.n566 VNB.n565 76
R2125 VNB.n562 VNB.n561 76
R2126 VNB.n556 VNB.n555 76
R2127 VNB.n552 VNB.n551 76
R2128 VNB.n548 VNB.n547 76
R2129 VNB.n544 VNB.n543 76
R2130 VNB.n540 VNB.n539 76
R2131 VNB.n536 VNB.n535 76
R2132 VNB.n532 VNB.n531 76
R2133 VNB.n528 VNB.n527 76
R2134 VNB.n524 VNB.n523 76
R2135 VNB.n502 VNB.n501 76
R2136 VNB.n498 VNB.n497 76
R2137 VNB.n494 VNB.n493 76
R2138 VNB.n482 VNB.n481 76
R2139 VNB.n477 VNB.n476 76
R2140 VNB.n473 VNB.n472 76
R2141 VNB.n469 VNB.n468 76
R2142 VNB.n465 VNB.n464 76
R2143 VNB.n461 VNB.n460 76
R2144 VNB.n457 VNB.n456 76
R2145 VNB.n453 VNB.n452 76
R2146 VNB.n449 VNB.n448 76
R2147 VNB.n427 VNB.n426 76
R2148 VNB.n423 VNB.n422 76
R2149 VNB.n419 VNB.n418 76
R2150 VNB.n413 VNB.n412 76
R2151 VNB.n409 VNB.n408 76
R2152 VNB.n405 VNB.n404 76
R2153 VNB.n401 VNB.n400 76
R2154 VNB.n397 VNB.n396 76
R2155 VNB.n393 VNB.n392 76
R2156 VNB.n389 VNB.n388 76
R2157 VNB.n385 VNB.n384 76
R2158 VNB.n381 VNB.n380 76
R2159 VNB.n359 VNB.n358 76
R2160 VNB.n355 VNB.n354 76
R2161 VNB.n351 VNB.n350 76
R2162 VNB.n345 VNB.n344 76
R2163 VNB.n341 VNB.n340 76
R2164 VNB.n337 VNB.n336 76
R2165 VNB.n333 VNB.n332 76
R2166 VNB.n329 VNB.n328 76
R2167 VNB.n325 VNB.n324 76
R2168 VNB.n321 VNB.n320 76
R2169 VNB.n317 VNB.n316 76
R2170 VNB.n313 VNB.n312 76
R2171 VNB.n291 VNB.n290 76
R2172 VNB.n287 VNB.n286 76
R2173 VNB.n283 VNB.n282 76
R2174 VNB.n277 VNB.n276 76
R2175 VNB.n273 VNB.n272 76
R2176 VNB.n269 VNB.n268 76
R2177 VNB.n265 VNB.n264 76
R2178 VNB.n261 VNB.n260 76
R2179 VNB.n239 VNB.n238 76
R2180 VNB.n235 VNB.n234 76
R2181 VNB.n231 VNB.n230 76
R2182 VNB.n225 VNB.n224 76
R2183 VNB.n221 VNB.n220 76
R2184 VNB.n217 VNB.n216 76
R2185 VNB.n213 VNB.n212 76
R2186 VNB.n209 VNB.n208 76
R2187 VNB.n187 VNB.n186 76
R2188 VNB.n183 VNB.n182 76
R2189 VNB.n179 VNB.n178 76
R2190 VNB.n173 VNB.n172 76
R2191 VNB.n137 VNB.n136 73.875
R2192 VNB.n61 VNB.n60 73.875
R2193 VNB.n487 VNB.n486 64.552
R2194 VNB.n698 VNB.n697 64.552
R2195 VNB.n135 VNB.n83 64.552
R2196 VNB.n1044 VNB.n1043 64.552
R2197 VNB.n59 VNB.n7 64.552
R2198 VNB.n349 VNB.n348 41.971
R2199 VNB.n417 VNB.n416 41.971
R2200 VNB.n560 VNB.n559 41.971
R2201 VNB.n628 VNB.n627 41.971
R2202 VNB.n771 VNB.n770 41.971
R2203 VNB.n838 VNB.n837 41.971
R2204 VNB.n906 VNB.n905 41.971
R2205 VNB.n974 VNB.n973 41.971
R2206 VNB.n1117 VNB.n1116 41.971
R2207 VNB.n1185 VNB.n1184 41.971
R2208 VNB.n1253 VNB.n1252 41.971
R2209 VNB.n1321 VNB.n1320 41.971
R2210 VNB.n1389 VNB.n1388 41.971
R2211 VNB.n491 VNB.n490 36.937
R2212 VNB.n702 VNB.n701 36.937
R2213 VNB.n132 VNB.n131 36.937
R2214 VNB.n1048 VNB.n1047 36.937
R2215 VNB.n56 VNB.n55 36.937
R2216 VNB.n177 VNB.n176 36.678
R2217 VNB.n229 VNB.n228 36.678
R2218 VNB.n281 VNB.n280 36.678
R2219 VNB.n168 VNB.n167 35.118
R2220 VNB.n490 VNB.n489 29.844
R2221 VNB.n701 VNB.n700 29.844
R2222 VNB.n1047 VNB.n1046 29.844
R2223 VNB.n486 VNB.n485 28.421
R2224 VNB.n697 VNB.n696 28.421
R2225 VNB.n83 VNB.n82 28.421
R2226 VNB.n1043 VNB.n1042 28.421
R2227 VNB.n7 VNB.n6 28.421
R2228 VNB.n486 VNB.n484 25.263
R2229 VNB.n697 VNB.n695 25.263
R2230 VNB.n83 VNB.n81 25.263
R2231 VNB.n1043 VNB.n1041 25.263
R2232 VNB.n7 VNB.n5 25.263
R2233 VNB.n484 VNB.n483 24.383
R2234 VNB.n695 VNB.n694 24.383
R2235 VNB.n81 VNB.n80 24.383
R2236 VNB.n1041 VNB.n1040 24.383
R2237 VNB.n5 VNB.n4 24.383
R2238 VNB.n157 VNB.n154 20.452
R2239 VNB.n1413 VNB.n1412 20.452
R2240 VNB.n166 VNB.n165 13.653
R2241 VNB.n165 VNB.n164 13.653
R2242 VNB.n163 VNB.n162 13.653
R2243 VNB.n162 VNB.n161 13.653
R2244 VNB.n160 VNB.n159 13.653
R2245 VNB.n159 VNB.n158 13.653
R2246 VNB.n172 VNB.n171 13.653
R2247 VNB.n171 VNB.n170 13.653
R2248 VNB.n178 VNB.n177 13.653
R2249 VNB.n182 VNB.n181 13.653
R2250 VNB.n181 VNB.n180 13.653
R2251 VNB.n186 VNB.n185 13.653
R2252 VNB.n185 VNB.n184 13.653
R2253 VNB.n208 VNB.n207 13.653
R2254 VNB.n207 VNB.n206 13.653
R2255 VNB.n212 VNB.n211 13.653
R2256 VNB.n211 VNB.n210 13.653
R2257 VNB.n216 VNB.n215 13.653
R2258 VNB.n215 VNB.n214 13.653
R2259 VNB.n220 VNB.n219 13.653
R2260 VNB.n219 VNB.n218 13.653
R2261 VNB.n224 VNB.n223 13.653
R2262 VNB.n223 VNB.n222 13.653
R2263 VNB.n230 VNB.n229 13.653
R2264 VNB.n234 VNB.n233 13.653
R2265 VNB.n233 VNB.n232 13.653
R2266 VNB.n238 VNB.n237 13.653
R2267 VNB.n237 VNB.n236 13.653
R2268 VNB.n260 VNB.n259 13.653
R2269 VNB.n259 VNB.n258 13.653
R2270 VNB.n264 VNB.n263 13.653
R2271 VNB.n263 VNB.n262 13.653
R2272 VNB.n268 VNB.n267 13.653
R2273 VNB.n267 VNB.n266 13.653
R2274 VNB.n272 VNB.n271 13.653
R2275 VNB.n271 VNB.n270 13.653
R2276 VNB.n276 VNB.n275 13.653
R2277 VNB.n275 VNB.n274 13.653
R2278 VNB.n282 VNB.n281 13.653
R2279 VNB.n286 VNB.n285 13.653
R2280 VNB.n285 VNB.n284 13.653
R2281 VNB.n290 VNB.n289 13.653
R2282 VNB.n289 VNB.n288 13.653
R2283 VNB.n312 VNB.n311 13.653
R2284 VNB.n311 VNB.n310 13.653
R2285 VNB.n316 VNB.n315 13.653
R2286 VNB.n315 VNB.n314 13.653
R2287 VNB.n320 VNB.n319 13.653
R2288 VNB.n319 VNB.n318 13.653
R2289 VNB.n324 VNB.n323 13.653
R2290 VNB.n323 VNB.n322 13.653
R2291 VNB.n328 VNB.n327 13.653
R2292 VNB.n327 VNB.n326 13.653
R2293 VNB.n332 VNB.n331 13.653
R2294 VNB.n331 VNB.n330 13.653
R2295 VNB.n336 VNB.n335 13.653
R2296 VNB.n335 VNB.n334 13.653
R2297 VNB.n340 VNB.n339 13.653
R2298 VNB.n339 VNB.n338 13.653
R2299 VNB.n344 VNB.n343 13.653
R2300 VNB.n343 VNB.n342 13.653
R2301 VNB.n350 VNB.n349 13.653
R2302 VNB.n354 VNB.n353 13.653
R2303 VNB.n353 VNB.n352 13.653
R2304 VNB.n358 VNB.n357 13.653
R2305 VNB.n357 VNB.n356 13.653
R2306 VNB.n380 VNB.n379 13.653
R2307 VNB.n379 VNB.n378 13.653
R2308 VNB.n384 VNB.n383 13.653
R2309 VNB.n383 VNB.n382 13.653
R2310 VNB.n388 VNB.n387 13.653
R2311 VNB.n387 VNB.n386 13.653
R2312 VNB.n392 VNB.n391 13.653
R2313 VNB.n391 VNB.n390 13.653
R2314 VNB.n396 VNB.n395 13.653
R2315 VNB.n395 VNB.n394 13.653
R2316 VNB.n400 VNB.n399 13.653
R2317 VNB.n399 VNB.n398 13.653
R2318 VNB.n404 VNB.n403 13.653
R2319 VNB.n403 VNB.n402 13.653
R2320 VNB.n408 VNB.n407 13.653
R2321 VNB.n407 VNB.n406 13.653
R2322 VNB.n412 VNB.n411 13.653
R2323 VNB.n411 VNB.n410 13.653
R2324 VNB.n418 VNB.n417 13.653
R2325 VNB.n422 VNB.n421 13.653
R2326 VNB.n421 VNB.n420 13.653
R2327 VNB.n426 VNB.n425 13.653
R2328 VNB.n425 VNB.n424 13.653
R2329 VNB.n448 VNB.n447 13.653
R2330 VNB.n447 VNB.n446 13.653
R2331 VNB.n452 VNB.n451 13.653
R2332 VNB.n451 VNB.n450 13.653
R2333 VNB.n456 VNB.n455 13.653
R2334 VNB.n455 VNB.n454 13.653
R2335 VNB.n460 VNB.n459 13.653
R2336 VNB.n459 VNB.n458 13.653
R2337 VNB.n464 VNB.n463 13.653
R2338 VNB.n463 VNB.n462 13.653
R2339 VNB.n468 VNB.n467 13.653
R2340 VNB.n467 VNB.n466 13.653
R2341 VNB.n472 VNB.n471 13.653
R2342 VNB.n471 VNB.n470 13.653
R2343 VNB.n476 VNB.n475 13.653
R2344 VNB.n475 VNB.n474 13.653
R2345 VNB.n481 VNB.n480 13.653
R2346 VNB.n480 VNB.n479 13.653
R2347 VNB.n493 VNB.n492 13.653
R2348 VNB.n492 VNB.n491 13.653
R2349 VNB.n497 VNB.n496 13.653
R2350 VNB.n496 VNB.n495 13.653
R2351 VNB.n501 VNB.n500 13.653
R2352 VNB.n500 VNB.n499 13.653
R2353 VNB.n523 VNB.n522 13.653
R2354 VNB.n522 VNB.n521 13.653
R2355 VNB.n527 VNB.n526 13.653
R2356 VNB.n526 VNB.n525 13.653
R2357 VNB.n531 VNB.n530 13.653
R2358 VNB.n530 VNB.n529 13.653
R2359 VNB.n535 VNB.n534 13.653
R2360 VNB.n534 VNB.n533 13.653
R2361 VNB.n539 VNB.n538 13.653
R2362 VNB.n538 VNB.n537 13.653
R2363 VNB.n543 VNB.n542 13.653
R2364 VNB.n542 VNB.n541 13.653
R2365 VNB.n547 VNB.n546 13.653
R2366 VNB.n546 VNB.n545 13.653
R2367 VNB.n551 VNB.n550 13.653
R2368 VNB.n550 VNB.n549 13.653
R2369 VNB.n555 VNB.n554 13.653
R2370 VNB.n554 VNB.n553 13.653
R2371 VNB.n561 VNB.n560 13.653
R2372 VNB.n565 VNB.n564 13.653
R2373 VNB.n564 VNB.n563 13.653
R2374 VNB.n569 VNB.n568 13.653
R2375 VNB.n568 VNB.n567 13.653
R2376 VNB.n591 VNB.n590 13.653
R2377 VNB.n590 VNB.n589 13.653
R2378 VNB.n595 VNB.n594 13.653
R2379 VNB.n594 VNB.n593 13.653
R2380 VNB.n599 VNB.n598 13.653
R2381 VNB.n598 VNB.n597 13.653
R2382 VNB.n603 VNB.n602 13.653
R2383 VNB.n602 VNB.n601 13.653
R2384 VNB.n607 VNB.n606 13.653
R2385 VNB.n606 VNB.n605 13.653
R2386 VNB.n611 VNB.n610 13.653
R2387 VNB.n610 VNB.n609 13.653
R2388 VNB.n615 VNB.n614 13.653
R2389 VNB.n614 VNB.n613 13.653
R2390 VNB.n619 VNB.n618 13.653
R2391 VNB.n618 VNB.n617 13.653
R2392 VNB.n623 VNB.n622 13.653
R2393 VNB.n622 VNB.n621 13.653
R2394 VNB.n629 VNB.n628 13.653
R2395 VNB.n633 VNB.n632 13.653
R2396 VNB.n632 VNB.n631 13.653
R2397 VNB.n637 VNB.n636 13.653
R2398 VNB.n636 VNB.n635 13.653
R2399 VNB.n659 VNB.n658 13.653
R2400 VNB.n658 VNB.n657 13.653
R2401 VNB.n663 VNB.n662 13.653
R2402 VNB.n662 VNB.n661 13.653
R2403 VNB.n667 VNB.n666 13.653
R2404 VNB.n666 VNB.n665 13.653
R2405 VNB.n671 VNB.n670 13.653
R2406 VNB.n670 VNB.n669 13.653
R2407 VNB.n675 VNB.n674 13.653
R2408 VNB.n674 VNB.n673 13.653
R2409 VNB.n679 VNB.n678 13.653
R2410 VNB.n678 VNB.n677 13.653
R2411 VNB.n683 VNB.n682 13.653
R2412 VNB.n682 VNB.n681 13.653
R2413 VNB.n687 VNB.n686 13.653
R2414 VNB.n686 VNB.n685 13.653
R2415 VNB.n692 VNB.n691 13.653
R2416 VNB.n691 VNB.n690 13.653
R2417 VNB.n704 VNB.n703 13.653
R2418 VNB.n703 VNB.n702 13.653
R2419 VNB.n708 VNB.n707 13.653
R2420 VNB.n707 VNB.n706 13.653
R2421 VNB.n712 VNB.n711 13.653
R2422 VNB.n711 VNB.n710 13.653
R2423 VNB.n734 VNB.n733 13.653
R2424 VNB.n733 VNB.n732 13.653
R2425 VNB.n738 VNB.n737 13.653
R2426 VNB.n737 VNB.n736 13.653
R2427 VNB.n742 VNB.n741 13.653
R2428 VNB.n741 VNB.n740 13.653
R2429 VNB.n746 VNB.n745 13.653
R2430 VNB.n745 VNB.n744 13.653
R2431 VNB.n750 VNB.n749 13.653
R2432 VNB.n749 VNB.n748 13.653
R2433 VNB.n754 VNB.n753 13.653
R2434 VNB.n753 VNB.n752 13.653
R2435 VNB.n758 VNB.n757 13.653
R2436 VNB.n757 VNB.n756 13.653
R2437 VNB.n762 VNB.n761 13.653
R2438 VNB.n761 VNB.n760 13.653
R2439 VNB.n766 VNB.n765 13.653
R2440 VNB.n765 VNB.n764 13.653
R2441 VNB.n772 VNB.n771 13.653
R2442 VNB.n776 VNB.n775 13.653
R2443 VNB.n775 VNB.n774 13.653
R2444 VNB.n780 VNB.n779 13.653
R2445 VNB.n779 VNB.n778 13.653
R2446 VNB.n104 VNB.n103 13.653
R2447 VNB.n103 VNB.n102 13.653
R2448 VNB.n107 VNB.n106 13.653
R2449 VNB.n106 VNB.n105 13.653
R2450 VNB.n110 VNB.n109 13.653
R2451 VNB.n109 VNB.n108 13.653
R2452 VNB.n113 VNB.n112 13.653
R2453 VNB.n112 VNB.n111 13.653
R2454 VNB.n116 VNB.n115 13.653
R2455 VNB.n115 VNB.n114 13.653
R2456 VNB.n119 VNB.n118 13.653
R2457 VNB.n118 VNB.n117 13.653
R2458 VNB.n122 VNB.n121 13.653
R2459 VNB.n121 VNB.n120 13.653
R2460 VNB.n125 VNB.n124 13.653
R2461 VNB.n124 VNB.n123 13.653
R2462 VNB.n129 VNB.n128 13.653
R2463 VNB.n128 VNB.n127 13.653
R2464 VNB.n134 VNB.n133 13.653
R2465 VNB.n133 VNB.n132 13.653
R2466 VNB.n139 VNB.n138 13.653
R2467 VNB.n138 VNB.n137 13.653
R2468 VNB.n796 VNB.n795 13.653
R2469 VNB.n795 VNB.n794 13.653
R2470 VNB.n801 VNB.n800 13.653
R2471 VNB.n800 VNB.n799 13.653
R2472 VNB.n805 VNB.n804 13.653
R2473 VNB.n804 VNB.n803 13.653
R2474 VNB.n809 VNB.n808 13.653
R2475 VNB.n808 VNB.n807 13.653
R2476 VNB.n813 VNB.n812 13.653
R2477 VNB.n812 VNB.n811 13.653
R2478 VNB.n817 VNB.n816 13.653
R2479 VNB.n816 VNB.n815 13.653
R2480 VNB.n821 VNB.n820 13.653
R2481 VNB.n820 VNB.n819 13.653
R2482 VNB.n825 VNB.n824 13.653
R2483 VNB.n824 VNB.n823 13.653
R2484 VNB.n829 VNB.n828 13.653
R2485 VNB.n828 VNB.n827 13.653
R2486 VNB.n833 VNB.n832 13.653
R2487 VNB.n832 VNB.n831 13.653
R2488 VNB.n839 VNB.n838 13.653
R2489 VNB.n843 VNB.n842 13.653
R2490 VNB.n842 VNB.n841 13.653
R2491 VNB.n847 VNB.n846 13.653
R2492 VNB.n846 VNB.n845 13.653
R2493 VNB.n869 VNB.n868 13.653
R2494 VNB.n868 VNB.n867 13.653
R2495 VNB.n873 VNB.n872 13.653
R2496 VNB.n872 VNB.n871 13.653
R2497 VNB.n877 VNB.n876 13.653
R2498 VNB.n876 VNB.n875 13.653
R2499 VNB.n881 VNB.n880 13.653
R2500 VNB.n880 VNB.n879 13.653
R2501 VNB.n885 VNB.n884 13.653
R2502 VNB.n884 VNB.n883 13.653
R2503 VNB.n889 VNB.n888 13.653
R2504 VNB.n888 VNB.n887 13.653
R2505 VNB.n893 VNB.n892 13.653
R2506 VNB.n892 VNB.n891 13.653
R2507 VNB.n897 VNB.n896 13.653
R2508 VNB.n896 VNB.n895 13.653
R2509 VNB.n901 VNB.n900 13.653
R2510 VNB.n900 VNB.n899 13.653
R2511 VNB.n907 VNB.n906 13.653
R2512 VNB.n911 VNB.n910 13.653
R2513 VNB.n910 VNB.n909 13.653
R2514 VNB.n915 VNB.n914 13.653
R2515 VNB.n914 VNB.n913 13.653
R2516 VNB.n937 VNB.n936 13.653
R2517 VNB.n936 VNB.n935 13.653
R2518 VNB.n941 VNB.n940 13.653
R2519 VNB.n940 VNB.n939 13.653
R2520 VNB.n945 VNB.n944 13.653
R2521 VNB.n944 VNB.n943 13.653
R2522 VNB.n949 VNB.n948 13.653
R2523 VNB.n948 VNB.n947 13.653
R2524 VNB.n953 VNB.n952 13.653
R2525 VNB.n952 VNB.n951 13.653
R2526 VNB.n957 VNB.n956 13.653
R2527 VNB.n956 VNB.n955 13.653
R2528 VNB.n961 VNB.n960 13.653
R2529 VNB.n960 VNB.n959 13.653
R2530 VNB.n965 VNB.n964 13.653
R2531 VNB.n964 VNB.n963 13.653
R2532 VNB.n969 VNB.n968 13.653
R2533 VNB.n968 VNB.n967 13.653
R2534 VNB.n975 VNB.n974 13.653
R2535 VNB.n979 VNB.n978 13.653
R2536 VNB.n978 VNB.n977 13.653
R2537 VNB.n983 VNB.n982 13.653
R2538 VNB.n982 VNB.n981 13.653
R2539 VNB.n1005 VNB.n1004 13.653
R2540 VNB.n1004 VNB.n1003 13.653
R2541 VNB.n1009 VNB.n1008 13.653
R2542 VNB.n1008 VNB.n1007 13.653
R2543 VNB.n1013 VNB.n1012 13.653
R2544 VNB.n1012 VNB.n1011 13.653
R2545 VNB.n1017 VNB.n1016 13.653
R2546 VNB.n1016 VNB.n1015 13.653
R2547 VNB.n1021 VNB.n1020 13.653
R2548 VNB.n1020 VNB.n1019 13.653
R2549 VNB.n1025 VNB.n1024 13.653
R2550 VNB.n1024 VNB.n1023 13.653
R2551 VNB.n1029 VNB.n1028 13.653
R2552 VNB.n1028 VNB.n1027 13.653
R2553 VNB.n1033 VNB.n1032 13.653
R2554 VNB.n1032 VNB.n1031 13.653
R2555 VNB.n1038 VNB.n1037 13.653
R2556 VNB.n1037 VNB.n1036 13.653
R2557 VNB.n1050 VNB.n1049 13.653
R2558 VNB.n1049 VNB.n1048 13.653
R2559 VNB.n1054 VNB.n1053 13.653
R2560 VNB.n1053 VNB.n1052 13.653
R2561 VNB.n1058 VNB.n1057 13.653
R2562 VNB.n1057 VNB.n1056 13.653
R2563 VNB.n1080 VNB.n1079 13.653
R2564 VNB.n1079 VNB.n1078 13.653
R2565 VNB.n1084 VNB.n1083 13.653
R2566 VNB.n1083 VNB.n1082 13.653
R2567 VNB.n1088 VNB.n1087 13.653
R2568 VNB.n1087 VNB.n1086 13.653
R2569 VNB.n1092 VNB.n1091 13.653
R2570 VNB.n1091 VNB.n1090 13.653
R2571 VNB.n1096 VNB.n1095 13.653
R2572 VNB.n1095 VNB.n1094 13.653
R2573 VNB.n1100 VNB.n1099 13.653
R2574 VNB.n1099 VNB.n1098 13.653
R2575 VNB.n1104 VNB.n1103 13.653
R2576 VNB.n1103 VNB.n1102 13.653
R2577 VNB.n1108 VNB.n1107 13.653
R2578 VNB.n1107 VNB.n1106 13.653
R2579 VNB.n1112 VNB.n1111 13.653
R2580 VNB.n1111 VNB.n1110 13.653
R2581 VNB.n1118 VNB.n1117 13.653
R2582 VNB.n1122 VNB.n1121 13.653
R2583 VNB.n1121 VNB.n1120 13.653
R2584 VNB.n1126 VNB.n1125 13.653
R2585 VNB.n1125 VNB.n1124 13.653
R2586 VNB.n1148 VNB.n1147 13.653
R2587 VNB.n1147 VNB.n1146 13.653
R2588 VNB.n1152 VNB.n1151 13.653
R2589 VNB.n1151 VNB.n1150 13.653
R2590 VNB.n1156 VNB.n1155 13.653
R2591 VNB.n1155 VNB.n1154 13.653
R2592 VNB.n1160 VNB.n1159 13.653
R2593 VNB.n1159 VNB.n1158 13.653
R2594 VNB.n1164 VNB.n1163 13.653
R2595 VNB.n1163 VNB.n1162 13.653
R2596 VNB.n1168 VNB.n1167 13.653
R2597 VNB.n1167 VNB.n1166 13.653
R2598 VNB.n1172 VNB.n1171 13.653
R2599 VNB.n1171 VNB.n1170 13.653
R2600 VNB.n1176 VNB.n1175 13.653
R2601 VNB.n1175 VNB.n1174 13.653
R2602 VNB.n1180 VNB.n1179 13.653
R2603 VNB.n1179 VNB.n1178 13.653
R2604 VNB.n1186 VNB.n1185 13.653
R2605 VNB.n1190 VNB.n1189 13.653
R2606 VNB.n1189 VNB.n1188 13.653
R2607 VNB.n1194 VNB.n1193 13.653
R2608 VNB.n1193 VNB.n1192 13.653
R2609 VNB.n1216 VNB.n1215 13.653
R2610 VNB.n1215 VNB.n1214 13.653
R2611 VNB.n1220 VNB.n1219 13.653
R2612 VNB.n1219 VNB.n1218 13.653
R2613 VNB.n1224 VNB.n1223 13.653
R2614 VNB.n1223 VNB.n1222 13.653
R2615 VNB.n1228 VNB.n1227 13.653
R2616 VNB.n1227 VNB.n1226 13.653
R2617 VNB.n1232 VNB.n1231 13.653
R2618 VNB.n1231 VNB.n1230 13.653
R2619 VNB.n1236 VNB.n1235 13.653
R2620 VNB.n1235 VNB.n1234 13.653
R2621 VNB.n1240 VNB.n1239 13.653
R2622 VNB.n1239 VNB.n1238 13.653
R2623 VNB.n1244 VNB.n1243 13.653
R2624 VNB.n1243 VNB.n1242 13.653
R2625 VNB.n1248 VNB.n1247 13.653
R2626 VNB.n1247 VNB.n1246 13.653
R2627 VNB.n1254 VNB.n1253 13.653
R2628 VNB.n1258 VNB.n1257 13.653
R2629 VNB.n1257 VNB.n1256 13.653
R2630 VNB.n1262 VNB.n1261 13.653
R2631 VNB.n1261 VNB.n1260 13.653
R2632 VNB.n1284 VNB.n1283 13.653
R2633 VNB.n1283 VNB.n1282 13.653
R2634 VNB.n1288 VNB.n1287 13.653
R2635 VNB.n1287 VNB.n1286 13.653
R2636 VNB.n1292 VNB.n1291 13.653
R2637 VNB.n1291 VNB.n1290 13.653
R2638 VNB.n1296 VNB.n1295 13.653
R2639 VNB.n1295 VNB.n1294 13.653
R2640 VNB.n1300 VNB.n1299 13.653
R2641 VNB.n1299 VNB.n1298 13.653
R2642 VNB.n1304 VNB.n1303 13.653
R2643 VNB.n1303 VNB.n1302 13.653
R2644 VNB.n1308 VNB.n1307 13.653
R2645 VNB.n1307 VNB.n1306 13.653
R2646 VNB.n1312 VNB.n1311 13.653
R2647 VNB.n1311 VNB.n1310 13.653
R2648 VNB.n1316 VNB.n1315 13.653
R2649 VNB.n1315 VNB.n1314 13.653
R2650 VNB.n1322 VNB.n1321 13.653
R2651 VNB.n1326 VNB.n1325 13.653
R2652 VNB.n1325 VNB.n1324 13.653
R2653 VNB.n1330 VNB.n1329 13.653
R2654 VNB.n1329 VNB.n1328 13.653
R2655 VNB.n1352 VNB.n1351 13.653
R2656 VNB.n1351 VNB.n1350 13.653
R2657 VNB.n1356 VNB.n1355 13.653
R2658 VNB.n1355 VNB.n1354 13.653
R2659 VNB.n1360 VNB.n1359 13.653
R2660 VNB.n1359 VNB.n1358 13.653
R2661 VNB.n1364 VNB.n1363 13.653
R2662 VNB.n1363 VNB.n1362 13.653
R2663 VNB.n1368 VNB.n1367 13.653
R2664 VNB.n1367 VNB.n1366 13.653
R2665 VNB.n1372 VNB.n1371 13.653
R2666 VNB.n1371 VNB.n1370 13.653
R2667 VNB.n1376 VNB.n1375 13.653
R2668 VNB.n1375 VNB.n1374 13.653
R2669 VNB.n1380 VNB.n1379 13.653
R2670 VNB.n1379 VNB.n1378 13.653
R2671 VNB.n1384 VNB.n1383 13.653
R2672 VNB.n1383 VNB.n1382 13.653
R2673 VNB.n1390 VNB.n1389 13.653
R2674 VNB.n1394 VNB.n1393 13.653
R2675 VNB.n1393 VNB.n1392 13.653
R2676 VNB.n1398 VNB.n1397 13.653
R2677 VNB.n1397 VNB.n1396 13.653
R2678 VNB.n28 VNB.n27 13.653
R2679 VNB.n27 VNB.n26 13.653
R2680 VNB.n31 VNB.n30 13.653
R2681 VNB.n30 VNB.n29 13.653
R2682 VNB.n34 VNB.n33 13.653
R2683 VNB.n33 VNB.n32 13.653
R2684 VNB.n37 VNB.n36 13.653
R2685 VNB.n36 VNB.n35 13.653
R2686 VNB.n40 VNB.n39 13.653
R2687 VNB.n39 VNB.n38 13.653
R2688 VNB.n43 VNB.n42 13.653
R2689 VNB.n42 VNB.n41 13.653
R2690 VNB.n46 VNB.n45 13.653
R2691 VNB.n45 VNB.n44 13.653
R2692 VNB.n49 VNB.n48 13.653
R2693 VNB.n48 VNB.n47 13.653
R2694 VNB.n53 VNB.n52 13.653
R2695 VNB.n52 VNB.n51 13.653
R2696 VNB.n58 VNB.n57 13.653
R2697 VNB.n57 VNB.n56 13.653
R2698 VNB.n63 VNB.n62 13.653
R2699 VNB.n62 VNB.n61 13.653
R2700 VNB.n1412 VNB.n0 13.653
R2701 VNB VNB.n0 13.653
R2702 VNB.n157 VNB.n156 13.653
R2703 VNB.n156 VNB.n155 13.653
R2704 VNB.n1420 VNB.n1417 13.577
R2705 VNB.n142 VNB.n140 13.276
R2706 VNB.n154 VNB.n142 13.276
R2707 VNB.n190 VNB.n188 13.276
R2708 VNB.n203 VNB.n190 13.276
R2709 VNB.n242 VNB.n240 13.276
R2710 VNB.n255 VNB.n242 13.276
R2711 VNB.n294 VNB.n292 13.276
R2712 VNB.n307 VNB.n294 13.276
R2713 VNB.n362 VNB.n360 13.276
R2714 VNB.n375 VNB.n362 13.276
R2715 VNB.n430 VNB.n428 13.276
R2716 VNB.n443 VNB.n430 13.276
R2717 VNB.n505 VNB.n503 13.276
R2718 VNB.n518 VNB.n505 13.276
R2719 VNB.n573 VNB.n571 13.276
R2720 VNB.n586 VNB.n573 13.276
R2721 VNB.n641 VNB.n639 13.276
R2722 VNB.n654 VNB.n641 13.276
R2723 VNB.n716 VNB.n714 13.276
R2724 VNB.n729 VNB.n716 13.276
R2725 VNB.n86 VNB.n84 13.276
R2726 VNB.n99 VNB.n86 13.276
R2727 VNB.n66 VNB.n64 13.276
R2728 VNB.n79 VNB.n66 13.276
R2729 VNB.n851 VNB.n849 13.276
R2730 VNB.n864 VNB.n851 13.276
R2731 VNB.n919 VNB.n917 13.276
R2732 VNB.n932 VNB.n919 13.276
R2733 VNB.n987 VNB.n985 13.276
R2734 VNB.n1000 VNB.n987 13.276
R2735 VNB.n1062 VNB.n1060 13.276
R2736 VNB.n1075 VNB.n1062 13.276
R2737 VNB.n1130 VNB.n1128 13.276
R2738 VNB.n1143 VNB.n1130 13.276
R2739 VNB.n1198 VNB.n1196 13.276
R2740 VNB.n1211 VNB.n1198 13.276
R2741 VNB.n1266 VNB.n1264 13.276
R2742 VNB.n1279 VNB.n1266 13.276
R2743 VNB.n1334 VNB.n1332 13.276
R2744 VNB.n1347 VNB.n1334 13.276
R2745 VNB.n10 VNB.n8 13.276
R2746 VNB.n23 VNB.n10 13.276
R2747 VNB.n166 VNB.n163 13.276
R2748 VNB.n163 VNB.n160 13.276
R2749 VNB.n208 VNB.n204 13.276
R2750 VNB.n260 VNB.n256 13.276
R2751 VNB.n312 VNB.n308 13.276
R2752 VNB.n380 VNB.n376 13.276
R2753 VNB.n448 VNB.n444 13.276
R2754 VNB.n523 VNB.n519 13.276
R2755 VNB.n591 VNB.n587 13.276
R2756 VNB.n659 VNB.n655 13.276
R2757 VNB.n734 VNB.n730 13.276
R2758 VNB.n104 VNB.n100 13.276
R2759 VNB.n107 VNB.n104 13.276
R2760 VNB.n110 VNB.n107 13.276
R2761 VNB.n113 VNB.n110 13.276
R2762 VNB.n116 VNB.n113 13.276
R2763 VNB.n119 VNB.n116 13.276
R2764 VNB.n122 VNB.n119 13.276
R2765 VNB.n125 VNB.n122 13.276
R2766 VNB.n129 VNB.n125 13.276
R2767 VNB.n134 VNB.n129 13.276
R2768 VNB.n796 VNB.n139 13.276
R2769 VNB.n797 VNB.n796 13.276
R2770 VNB.n801 VNB.n797 13.276
R2771 VNB.n869 VNB.n865 13.276
R2772 VNB.n937 VNB.n933 13.276
R2773 VNB.n1005 VNB.n1001 13.276
R2774 VNB.n1080 VNB.n1076 13.276
R2775 VNB.n1148 VNB.n1144 13.276
R2776 VNB.n1216 VNB.n1212 13.276
R2777 VNB.n1284 VNB.n1280 13.276
R2778 VNB.n1352 VNB.n1348 13.276
R2779 VNB.n28 VNB.n24 13.276
R2780 VNB.n31 VNB.n28 13.276
R2781 VNB.n34 VNB.n31 13.276
R2782 VNB.n37 VNB.n34 13.276
R2783 VNB.n40 VNB.n37 13.276
R2784 VNB.n43 VNB.n40 13.276
R2785 VNB.n46 VNB.n43 13.276
R2786 VNB.n49 VNB.n46 13.276
R2787 VNB.n53 VNB.n49 13.276
R2788 VNB.n58 VNB.n53 13.276
R2789 VNB.n1412 VNB.n63 13.276
R2790 VNB.n3 VNB.n1 13.276
R2791 VNB.n1413 VNB.n3 13.276
R2792 VNB.n139 VNB.n135 12.02
R2793 VNB.n63 VNB.n59 12.02
R2794 VNB.n1422 VNB.n1421 7.5
R2795 VNB.n196 VNB.n195 7.5
R2796 VNB.n192 VNB.n191 7.5
R2797 VNB.n190 VNB.n189 7.5
R2798 VNB.n203 VNB.n202 7.5
R2799 VNB.n248 VNB.n247 7.5
R2800 VNB.n244 VNB.n243 7.5
R2801 VNB.n242 VNB.n241 7.5
R2802 VNB.n255 VNB.n254 7.5
R2803 VNB.n300 VNB.n299 7.5
R2804 VNB.n296 VNB.n295 7.5
R2805 VNB.n294 VNB.n293 7.5
R2806 VNB.n307 VNB.n306 7.5
R2807 VNB.n368 VNB.n367 7.5
R2808 VNB.n364 VNB.n363 7.5
R2809 VNB.n362 VNB.n361 7.5
R2810 VNB.n375 VNB.n374 7.5
R2811 VNB.n436 VNB.n435 7.5
R2812 VNB.n432 VNB.n431 7.5
R2813 VNB.n430 VNB.n429 7.5
R2814 VNB.n443 VNB.n442 7.5
R2815 VNB.n511 VNB.n510 7.5
R2816 VNB.n507 VNB.n506 7.5
R2817 VNB.n505 VNB.n504 7.5
R2818 VNB.n518 VNB.n517 7.5
R2819 VNB.n579 VNB.n578 7.5
R2820 VNB.n575 VNB.n574 7.5
R2821 VNB.n573 VNB.n572 7.5
R2822 VNB.n586 VNB.n585 7.5
R2823 VNB.n647 VNB.n646 7.5
R2824 VNB.n643 VNB.n642 7.5
R2825 VNB.n641 VNB.n640 7.5
R2826 VNB.n654 VNB.n653 7.5
R2827 VNB.n722 VNB.n721 7.5
R2828 VNB.n718 VNB.n717 7.5
R2829 VNB.n716 VNB.n715 7.5
R2830 VNB.n729 VNB.n728 7.5
R2831 VNB.n92 VNB.n91 7.5
R2832 VNB.n88 VNB.n87 7.5
R2833 VNB.n86 VNB.n85 7.5
R2834 VNB.n99 VNB.n98 7.5
R2835 VNB.n72 VNB.n71 7.5
R2836 VNB.n68 VNB.n67 7.5
R2837 VNB.n66 VNB.n65 7.5
R2838 VNB.n79 VNB.n78 7.5
R2839 VNB.n857 VNB.n856 7.5
R2840 VNB.n853 VNB.n852 7.5
R2841 VNB.n851 VNB.n850 7.5
R2842 VNB.n864 VNB.n863 7.5
R2843 VNB.n925 VNB.n924 7.5
R2844 VNB.n921 VNB.n920 7.5
R2845 VNB.n919 VNB.n918 7.5
R2846 VNB.n932 VNB.n931 7.5
R2847 VNB.n993 VNB.n992 7.5
R2848 VNB.n989 VNB.n988 7.5
R2849 VNB.n987 VNB.n986 7.5
R2850 VNB.n1000 VNB.n999 7.5
R2851 VNB.n1068 VNB.n1067 7.5
R2852 VNB.n1064 VNB.n1063 7.5
R2853 VNB.n1062 VNB.n1061 7.5
R2854 VNB.n1075 VNB.n1074 7.5
R2855 VNB.n1136 VNB.n1135 7.5
R2856 VNB.n1132 VNB.n1131 7.5
R2857 VNB.n1130 VNB.n1129 7.5
R2858 VNB.n1143 VNB.n1142 7.5
R2859 VNB.n1204 VNB.n1203 7.5
R2860 VNB.n1200 VNB.n1199 7.5
R2861 VNB.n1198 VNB.n1197 7.5
R2862 VNB.n1211 VNB.n1210 7.5
R2863 VNB.n1272 VNB.n1271 7.5
R2864 VNB.n1268 VNB.n1267 7.5
R2865 VNB.n1266 VNB.n1265 7.5
R2866 VNB.n1279 VNB.n1278 7.5
R2867 VNB.n1340 VNB.n1339 7.5
R2868 VNB.n1336 VNB.n1335 7.5
R2869 VNB.n1334 VNB.n1333 7.5
R2870 VNB.n1347 VNB.n1346 7.5
R2871 VNB.n16 VNB.n15 7.5
R2872 VNB.n12 VNB.n11 7.5
R2873 VNB.n10 VNB.n9 7.5
R2874 VNB.n23 VNB.n22 7.5
R2875 VNB.n1414 VNB.n1413 7.5
R2876 VNB.n3 VNB.n2 7.5
R2877 VNB.n1419 VNB.n1418 7.5
R2878 VNB.n148 VNB.n147 7.5
R2879 VNB.n144 VNB.n143 7.5
R2880 VNB.n142 VNB.n141 7.5
R2881 VNB.n154 VNB.n153 7.5
R2882 VNB.n204 VNB.n203 7.176
R2883 VNB.n256 VNB.n255 7.176
R2884 VNB.n308 VNB.n307 7.176
R2885 VNB.n376 VNB.n375 7.176
R2886 VNB.n444 VNB.n443 7.176
R2887 VNB.n519 VNB.n518 7.176
R2888 VNB.n587 VNB.n586 7.176
R2889 VNB.n655 VNB.n654 7.176
R2890 VNB.n730 VNB.n729 7.176
R2891 VNB.n100 VNB.n99 7.176
R2892 VNB.n797 VNB.n79 7.176
R2893 VNB.n865 VNB.n864 7.176
R2894 VNB.n933 VNB.n932 7.176
R2895 VNB.n1001 VNB.n1000 7.176
R2896 VNB.n1076 VNB.n1075 7.176
R2897 VNB.n1144 VNB.n1143 7.176
R2898 VNB.n1212 VNB.n1211 7.176
R2899 VNB.n1280 VNB.n1279 7.176
R2900 VNB.n1348 VNB.n1347 7.176
R2901 VNB.n24 VNB.n23 7.176
R2902 VNB.n1424 VNB.n1422 7.011
R2903 VNB.n199 VNB.n196 7.011
R2904 VNB.n194 VNB.n192 7.011
R2905 VNB.n251 VNB.n248 7.011
R2906 VNB.n246 VNB.n244 7.011
R2907 VNB.n303 VNB.n300 7.011
R2908 VNB.n298 VNB.n296 7.011
R2909 VNB.n371 VNB.n368 7.011
R2910 VNB.n366 VNB.n364 7.011
R2911 VNB.n439 VNB.n436 7.011
R2912 VNB.n434 VNB.n432 7.011
R2913 VNB.n514 VNB.n511 7.011
R2914 VNB.n509 VNB.n507 7.011
R2915 VNB.n582 VNB.n579 7.011
R2916 VNB.n577 VNB.n575 7.011
R2917 VNB.n650 VNB.n647 7.011
R2918 VNB.n645 VNB.n643 7.011
R2919 VNB.n725 VNB.n722 7.011
R2920 VNB.n720 VNB.n718 7.011
R2921 VNB.n95 VNB.n92 7.011
R2922 VNB.n90 VNB.n88 7.011
R2923 VNB.n75 VNB.n72 7.011
R2924 VNB.n70 VNB.n68 7.011
R2925 VNB.n860 VNB.n857 7.011
R2926 VNB.n855 VNB.n853 7.011
R2927 VNB.n928 VNB.n925 7.011
R2928 VNB.n923 VNB.n921 7.011
R2929 VNB.n996 VNB.n993 7.011
R2930 VNB.n991 VNB.n989 7.011
R2931 VNB.n1071 VNB.n1068 7.011
R2932 VNB.n1066 VNB.n1064 7.011
R2933 VNB.n1139 VNB.n1136 7.011
R2934 VNB.n1134 VNB.n1132 7.011
R2935 VNB.n1207 VNB.n1204 7.011
R2936 VNB.n1202 VNB.n1200 7.011
R2937 VNB.n1275 VNB.n1272 7.011
R2938 VNB.n1270 VNB.n1268 7.011
R2939 VNB.n1343 VNB.n1340 7.011
R2940 VNB.n1338 VNB.n1336 7.011
R2941 VNB.n19 VNB.n16 7.011
R2942 VNB.n14 VNB.n12 7.011
R2943 VNB.n150 VNB.n148 7.011
R2944 VNB.n146 VNB.n144 7.011
R2945 VNB.n202 VNB.n201 7.01
R2946 VNB.n194 VNB.n193 7.01
R2947 VNB.n199 VNB.n198 7.01
R2948 VNB.n254 VNB.n253 7.01
R2949 VNB.n246 VNB.n245 7.01
R2950 VNB.n251 VNB.n250 7.01
R2951 VNB.n306 VNB.n305 7.01
R2952 VNB.n298 VNB.n297 7.01
R2953 VNB.n303 VNB.n302 7.01
R2954 VNB.n374 VNB.n373 7.01
R2955 VNB.n366 VNB.n365 7.01
R2956 VNB.n371 VNB.n370 7.01
R2957 VNB.n442 VNB.n441 7.01
R2958 VNB.n434 VNB.n433 7.01
R2959 VNB.n439 VNB.n438 7.01
R2960 VNB.n517 VNB.n516 7.01
R2961 VNB.n509 VNB.n508 7.01
R2962 VNB.n514 VNB.n513 7.01
R2963 VNB.n585 VNB.n584 7.01
R2964 VNB.n577 VNB.n576 7.01
R2965 VNB.n582 VNB.n581 7.01
R2966 VNB.n653 VNB.n652 7.01
R2967 VNB.n645 VNB.n644 7.01
R2968 VNB.n650 VNB.n649 7.01
R2969 VNB.n728 VNB.n727 7.01
R2970 VNB.n720 VNB.n719 7.01
R2971 VNB.n725 VNB.n724 7.01
R2972 VNB.n98 VNB.n97 7.01
R2973 VNB.n90 VNB.n89 7.01
R2974 VNB.n95 VNB.n94 7.01
R2975 VNB.n78 VNB.n77 7.01
R2976 VNB.n70 VNB.n69 7.01
R2977 VNB.n75 VNB.n74 7.01
R2978 VNB.n863 VNB.n862 7.01
R2979 VNB.n855 VNB.n854 7.01
R2980 VNB.n860 VNB.n859 7.01
R2981 VNB.n931 VNB.n930 7.01
R2982 VNB.n923 VNB.n922 7.01
R2983 VNB.n928 VNB.n927 7.01
R2984 VNB.n999 VNB.n998 7.01
R2985 VNB.n991 VNB.n990 7.01
R2986 VNB.n996 VNB.n995 7.01
R2987 VNB.n1074 VNB.n1073 7.01
R2988 VNB.n1066 VNB.n1065 7.01
R2989 VNB.n1071 VNB.n1070 7.01
R2990 VNB.n1142 VNB.n1141 7.01
R2991 VNB.n1134 VNB.n1133 7.01
R2992 VNB.n1139 VNB.n1138 7.01
R2993 VNB.n1210 VNB.n1209 7.01
R2994 VNB.n1202 VNB.n1201 7.01
R2995 VNB.n1207 VNB.n1206 7.01
R2996 VNB.n1278 VNB.n1277 7.01
R2997 VNB.n1270 VNB.n1269 7.01
R2998 VNB.n1275 VNB.n1274 7.01
R2999 VNB.n1346 VNB.n1345 7.01
R3000 VNB.n1338 VNB.n1337 7.01
R3001 VNB.n1343 VNB.n1342 7.01
R3002 VNB.n22 VNB.n21 7.01
R3003 VNB.n14 VNB.n13 7.01
R3004 VNB.n19 VNB.n18 7.01
R3005 VNB.n153 VNB.n152 7.01
R3006 VNB.n146 VNB.n145 7.01
R3007 VNB.n150 VNB.n149 7.01
R3008 VNB.n1424 VNB.n1423 7.01
R3009 VNB.n1420 VNB.n1419 6.788
R3010 VNB.n1415 VNB.n1414 6.788
R3011 VNB.n167 VNB.n157 6.111
R3012 VNB.n167 VNB.n166 6.1
R3013 VNB.n178 VNB.n175 2.511
R3014 VNB.n230 VNB.n227 2.511
R3015 VNB.n282 VNB.n279 2.511
R3016 VNB.n350 VNB.n347 1.255
R3017 VNB.n418 VNB.n415 1.255
R3018 VNB.n493 VNB.n487 1.255
R3019 VNB.n561 VNB.n558 1.255
R3020 VNB.n629 VNB.n626 1.255
R3021 VNB.n704 VNB.n698 1.255
R3022 VNB.n772 VNB.n769 1.255
R3023 VNB.n135 VNB.n134 1.255
R3024 VNB.n839 VNB.n836 1.255
R3025 VNB.n907 VNB.n904 1.255
R3026 VNB.n975 VNB.n972 1.255
R3027 VNB.n1050 VNB.n1044 1.255
R3028 VNB.n1118 VNB.n1115 1.255
R3029 VNB.n1186 VNB.n1183 1.255
R3030 VNB.n1254 VNB.n1251 1.255
R3031 VNB.n1322 VNB.n1319 1.255
R3032 VNB.n1390 VNB.n1387 1.255
R3033 VNB.n59 VNB.n58 1.255
R3034 VNB.n1425 VNB.n1416 0.921
R3035 VNB.n1425 VNB.n1420 0.476
R3036 VNB.n1425 VNB.n1415 0.475
R3037 VNB.n209 VNB.n187 0.272
R3038 VNB.n261 VNB.n239 0.272
R3039 VNB.n313 VNB.n291 0.272
R3040 VNB.n381 VNB.n359 0.272
R3041 VNB.n449 VNB.n427 0.272
R3042 VNB.n524 VNB.n502 0.272
R3043 VNB.n592 VNB.n570 0.272
R3044 VNB.n660 VNB.n638 0.272
R3045 VNB.n735 VNB.n713 0.272
R3046 VNB.n782 VNB.n781 0.272
R3047 VNB.n870 VNB.n848 0.272
R3048 VNB.n938 VNB.n916 0.272
R3049 VNB.n1006 VNB.n984 0.272
R3050 VNB.n1081 VNB.n1059 0.272
R3051 VNB.n1149 VNB.n1127 0.272
R3052 VNB.n1217 VNB.n1195 0.272
R3053 VNB.n1285 VNB.n1263 0.272
R3054 VNB.n1353 VNB.n1331 0.272
R3055 VNB.n1400 VNB.n1399 0.272
R3056 VNB.n200 VNB.n194 0.246
R3057 VNB.n201 VNB.n200 0.246
R3058 VNB.n200 VNB.n199 0.246
R3059 VNB.n252 VNB.n246 0.246
R3060 VNB.n253 VNB.n252 0.246
R3061 VNB.n252 VNB.n251 0.246
R3062 VNB.n304 VNB.n298 0.246
R3063 VNB.n305 VNB.n304 0.246
R3064 VNB.n304 VNB.n303 0.246
R3065 VNB.n372 VNB.n366 0.246
R3066 VNB.n373 VNB.n372 0.246
R3067 VNB.n372 VNB.n371 0.246
R3068 VNB.n440 VNB.n434 0.246
R3069 VNB.n441 VNB.n440 0.246
R3070 VNB.n440 VNB.n439 0.246
R3071 VNB.n515 VNB.n509 0.246
R3072 VNB.n516 VNB.n515 0.246
R3073 VNB.n515 VNB.n514 0.246
R3074 VNB.n583 VNB.n577 0.246
R3075 VNB.n584 VNB.n583 0.246
R3076 VNB.n583 VNB.n582 0.246
R3077 VNB.n651 VNB.n645 0.246
R3078 VNB.n652 VNB.n651 0.246
R3079 VNB.n651 VNB.n650 0.246
R3080 VNB.n726 VNB.n720 0.246
R3081 VNB.n727 VNB.n726 0.246
R3082 VNB.n726 VNB.n725 0.246
R3083 VNB.n96 VNB.n90 0.246
R3084 VNB.n97 VNB.n96 0.246
R3085 VNB.n96 VNB.n95 0.246
R3086 VNB.n76 VNB.n70 0.246
R3087 VNB.n77 VNB.n76 0.246
R3088 VNB.n76 VNB.n75 0.246
R3089 VNB.n861 VNB.n855 0.246
R3090 VNB.n862 VNB.n861 0.246
R3091 VNB.n861 VNB.n860 0.246
R3092 VNB.n929 VNB.n923 0.246
R3093 VNB.n930 VNB.n929 0.246
R3094 VNB.n929 VNB.n928 0.246
R3095 VNB.n997 VNB.n991 0.246
R3096 VNB.n998 VNB.n997 0.246
R3097 VNB.n997 VNB.n996 0.246
R3098 VNB.n1072 VNB.n1066 0.246
R3099 VNB.n1073 VNB.n1072 0.246
R3100 VNB.n1072 VNB.n1071 0.246
R3101 VNB.n1140 VNB.n1134 0.246
R3102 VNB.n1141 VNB.n1140 0.246
R3103 VNB.n1140 VNB.n1139 0.246
R3104 VNB.n1208 VNB.n1202 0.246
R3105 VNB.n1209 VNB.n1208 0.246
R3106 VNB.n1208 VNB.n1207 0.246
R3107 VNB.n1276 VNB.n1270 0.246
R3108 VNB.n1277 VNB.n1276 0.246
R3109 VNB.n1276 VNB.n1275 0.246
R3110 VNB.n1344 VNB.n1338 0.246
R3111 VNB.n1345 VNB.n1344 0.246
R3112 VNB.n1344 VNB.n1343 0.246
R3113 VNB.n20 VNB.n14 0.246
R3114 VNB.n21 VNB.n20 0.246
R3115 VNB.n20 VNB.n19 0.246
R3116 VNB.n151 VNB.n146 0.246
R3117 VNB.n152 VNB.n151 0.246
R3118 VNB.n151 VNB.n150 0.246
R3119 VNB.n1425 VNB.n1424 0.246
R3120 VNB.n802 VNB 0.204
R3121 VNB.n1411 VNB 0.198
R3122 VNB.n169 VNB.n168 0.136
R3123 VNB.n173 VNB.n169 0.136
R3124 VNB.n179 VNB.n173 0.136
R3125 VNB.n183 VNB.n179 0.136
R3126 VNB.n187 VNB.n183 0.136
R3127 VNB.n213 VNB.n209 0.136
R3128 VNB.n217 VNB.n213 0.136
R3129 VNB.n221 VNB.n217 0.136
R3130 VNB.n225 VNB.n221 0.136
R3131 VNB.n231 VNB.n225 0.136
R3132 VNB.n235 VNB.n231 0.136
R3133 VNB.n239 VNB.n235 0.136
R3134 VNB.n265 VNB.n261 0.136
R3135 VNB.n269 VNB.n265 0.136
R3136 VNB.n273 VNB.n269 0.136
R3137 VNB.n277 VNB.n273 0.136
R3138 VNB.n283 VNB.n277 0.136
R3139 VNB.n287 VNB.n283 0.136
R3140 VNB.n291 VNB.n287 0.136
R3141 VNB.n317 VNB.n313 0.136
R3142 VNB.n321 VNB.n317 0.136
R3143 VNB.n325 VNB.n321 0.136
R3144 VNB.n329 VNB.n325 0.136
R3145 VNB.n333 VNB.n329 0.136
R3146 VNB.n337 VNB.n333 0.136
R3147 VNB.n341 VNB.n337 0.136
R3148 VNB.n345 VNB.n341 0.136
R3149 VNB.n351 VNB.n345 0.136
R3150 VNB.n355 VNB.n351 0.136
R3151 VNB.n359 VNB.n355 0.136
R3152 VNB.n385 VNB.n381 0.136
R3153 VNB.n389 VNB.n385 0.136
R3154 VNB.n393 VNB.n389 0.136
R3155 VNB.n397 VNB.n393 0.136
R3156 VNB.n401 VNB.n397 0.136
R3157 VNB.n405 VNB.n401 0.136
R3158 VNB.n409 VNB.n405 0.136
R3159 VNB.n413 VNB.n409 0.136
R3160 VNB.n419 VNB.n413 0.136
R3161 VNB.n423 VNB.n419 0.136
R3162 VNB.n427 VNB.n423 0.136
R3163 VNB.n453 VNB.n449 0.136
R3164 VNB.n457 VNB.n453 0.136
R3165 VNB.n461 VNB.n457 0.136
R3166 VNB.n465 VNB.n461 0.136
R3167 VNB.n469 VNB.n465 0.136
R3168 VNB.n473 VNB.n469 0.136
R3169 VNB.n477 VNB.n473 0.136
R3170 VNB.n482 VNB.n477 0.136
R3171 VNB.n494 VNB.n482 0.136
R3172 VNB.n498 VNB.n494 0.136
R3173 VNB.n502 VNB.n498 0.136
R3174 VNB.n528 VNB.n524 0.136
R3175 VNB.n532 VNB.n528 0.136
R3176 VNB.n536 VNB.n532 0.136
R3177 VNB.n540 VNB.n536 0.136
R3178 VNB.n544 VNB.n540 0.136
R3179 VNB.n548 VNB.n544 0.136
R3180 VNB.n552 VNB.n548 0.136
R3181 VNB.n556 VNB.n552 0.136
R3182 VNB.n562 VNB.n556 0.136
R3183 VNB.n566 VNB.n562 0.136
R3184 VNB.n570 VNB.n566 0.136
R3185 VNB.n596 VNB.n592 0.136
R3186 VNB.n600 VNB.n596 0.136
R3187 VNB.n604 VNB.n600 0.136
R3188 VNB.n608 VNB.n604 0.136
R3189 VNB.n612 VNB.n608 0.136
R3190 VNB.n616 VNB.n612 0.136
R3191 VNB.n620 VNB.n616 0.136
R3192 VNB.n624 VNB.n620 0.136
R3193 VNB.n630 VNB.n624 0.136
R3194 VNB.n634 VNB.n630 0.136
R3195 VNB.n638 VNB.n634 0.136
R3196 VNB.n664 VNB.n660 0.136
R3197 VNB.n668 VNB.n664 0.136
R3198 VNB.n672 VNB.n668 0.136
R3199 VNB.n676 VNB.n672 0.136
R3200 VNB.n680 VNB.n676 0.136
R3201 VNB.n684 VNB.n680 0.136
R3202 VNB.n688 VNB.n684 0.136
R3203 VNB.n693 VNB.n688 0.136
R3204 VNB.n705 VNB.n693 0.136
R3205 VNB.n709 VNB.n705 0.136
R3206 VNB.n713 VNB.n709 0.136
R3207 VNB.n739 VNB.n735 0.136
R3208 VNB.n743 VNB.n739 0.136
R3209 VNB.n747 VNB.n743 0.136
R3210 VNB.n751 VNB.n747 0.136
R3211 VNB.n755 VNB.n751 0.136
R3212 VNB.n759 VNB.n755 0.136
R3213 VNB.n763 VNB.n759 0.136
R3214 VNB.n767 VNB.n763 0.136
R3215 VNB.n773 VNB.n767 0.136
R3216 VNB.n777 VNB.n773 0.136
R3217 VNB.n781 VNB.n777 0.136
R3218 VNB.n783 VNB.n782 0.136
R3219 VNB.n784 VNB.n783 0.136
R3220 VNB.n785 VNB.n784 0.136
R3221 VNB.n786 VNB.n785 0.136
R3222 VNB.n787 VNB.n786 0.136
R3223 VNB.n788 VNB.n787 0.136
R3224 VNB.n789 VNB.n788 0.136
R3225 VNB.n790 VNB.n789 0.136
R3226 VNB.n791 VNB.n790 0.136
R3227 VNB.n792 VNB.n791 0.136
R3228 VNB.n793 VNB.n792 0.136
R3229 VNB.n806 VNB.n802 0.136
R3230 VNB.n810 VNB.n806 0.136
R3231 VNB.n814 VNB.n810 0.136
R3232 VNB.n818 VNB.n814 0.136
R3233 VNB.n822 VNB.n818 0.136
R3234 VNB.n826 VNB.n822 0.136
R3235 VNB.n830 VNB.n826 0.136
R3236 VNB.n834 VNB.n830 0.136
R3237 VNB.n840 VNB.n834 0.136
R3238 VNB.n844 VNB.n840 0.136
R3239 VNB.n848 VNB.n844 0.136
R3240 VNB.n874 VNB.n870 0.136
R3241 VNB.n878 VNB.n874 0.136
R3242 VNB.n882 VNB.n878 0.136
R3243 VNB.n886 VNB.n882 0.136
R3244 VNB.n890 VNB.n886 0.136
R3245 VNB.n894 VNB.n890 0.136
R3246 VNB.n898 VNB.n894 0.136
R3247 VNB.n902 VNB.n898 0.136
R3248 VNB.n908 VNB.n902 0.136
R3249 VNB.n912 VNB.n908 0.136
R3250 VNB.n916 VNB.n912 0.136
R3251 VNB.n942 VNB.n938 0.136
R3252 VNB.n946 VNB.n942 0.136
R3253 VNB.n950 VNB.n946 0.136
R3254 VNB.n954 VNB.n950 0.136
R3255 VNB.n958 VNB.n954 0.136
R3256 VNB.n962 VNB.n958 0.136
R3257 VNB.n966 VNB.n962 0.136
R3258 VNB.n970 VNB.n966 0.136
R3259 VNB.n976 VNB.n970 0.136
R3260 VNB.n980 VNB.n976 0.136
R3261 VNB.n984 VNB.n980 0.136
R3262 VNB.n1010 VNB.n1006 0.136
R3263 VNB.n1014 VNB.n1010 0.136
R3264 VNB.n1018 VNB.n1014 0.136
R3265 VNB.n1022 VNB.n1018 0.136
R3266 VNB.n1026 VNB.n1022 0.136
R3267 VNB.n1030 VNB.n1026 0.136
R3268 VNB.n1034 VNB.n1030 0.136
R3269 VNB.n1039 VNB.n1034 0.136
R3270 VNB.n1051 VNB.n1039 0.136
R3271 VNB.n1055 VNB.n1051 0.136
R3272 VNB.n1059 VNB.n1055 0.136
R3273 VNB.n1085 VNB.n1081 0.136
R3274 VNB.n1089 VNB.n1085 0.136
R3275 VNB.n1093 VNB.n1089 0.136
R3276 VNB.n1097 VNB.n1093 0.136
R3277 VNB.n1101 VNB.n1097 0.136
R3278 VNB.n1105 VNB.n1101 0.136
R3279 VNB.n1109 VNB.n1105 0.136
R3280 VNB.n1113 VNB.n1109 0.136
R3281 VNB.n1119 VNB.n1113 0.136
R3282 VNB.n1123 VNB.n1119 0.136
R3283 VNB.n1127 VNB.n1123 0.136
R3284 VNB.n1153 VNB.n1149 0.136
R3285 VNB.n1157 VNB.n1153 0.136
R3286 VNB.n1161 VNB.n1157 0.136
R3287 VNB.n1165 VNB.n1161 0.136
R3288 VNB.n1169 VNB.n1165 0.136
R3289 VNB.n1173 VNB.n1169 0.136
R3290 VNB.n1177 VNB.n1173 0.136
R3291 VNB.n1181 VNB.n1177 0.136
R3292 VNB.n1187 VNB.n1181 0.136
R3293 VNB.n1191 VNB.n1187 0.136
R3294 VNB.n1195 VNB.n1191 0.136
R3295 VNB.n1221 VNB.n1217 0.136
R3296 VNB.n1225 VNB.n1221 0.136
R3297 VNB.n1229 VNB.n1225 0.136
R3298 VNB.n1233 VNB.n1229 0.136
R3299 VNB.n1237 VNB.n1233 0.136
R3300 VNB.n1241 VNB.n1237 0.136
R3301 VNB.n1245 VNB.n1241 0.136
R3302 VNB.n1249 VNB.n1245 0.136
R3303 VNB.n1255 VNB.n1249 0.136
R3304 VNB.n1259 VNB.n1255 0.136
R3305 VNB.n1263 VNB.n1259 0.136
R3306 VNB.n1289 VNB.n1285 0.136
R3307 VNB.n1293 VNB.n1289 0.136
R3308 VNB.n1297 VNB.n1293 0.136
R3309 VNB.n1301 VNB.n1297 0.136
R3310 VNB.n1305 VNB.n1301 0.136
R3311 VNB.n1309 VNB.n1305 0.136
R3312 VNB.n1313 VNB.n1309 0.136
R3313 VNB.n1317 VNB.n1313 0.136
R3314 VNB.n1323 VNB.n1317 0.136
R3315 VNB.n1327 VNB.n1323 0.136
R3316 VNB.n1331 VNB.n1327 0.136
R3317 VNB.n1357 VNB.n1353 0.136
R3318 VNB.n1361 VNB.n1357 0.136
R3319 VNB.n1365 VNB.n1361 0.136
R3320 VNB.n1369 VNB.n1365 0.136
R3321 VNB.n1373 VNB.n1369 0.136
R3322 VNB.n1377 VNB.n1373 0.136
R3323 VNB.n1381 VNB.n1377 0.136
R3324 VNB.n1385 VNB.n1381 0.136
R3325 VNB.n1391 VNB.n1385 0.136
R3326 VNB.n1395 VNB.n1391 0.136
R3327 VNB.n1399 VNB.n1395 0.136
R3328 VNB.n1401 VNB.n1400 0.136
R3329 VNB.n1402 VNB.n1401 0.136
R3330 VNB.n1403 VNB.n1402 0.136
R3331 VNB.n1404 VNB.n1403 0.136
R3332 VNB.n1405 VNB.n1404 0.136
R3333 VNB.n1406 VNB.n1405 0.136
R3334 VNB.n1407 VNB.n1406 0.136
R3335 VNB.n1408 VNB.n1407 0.136
R3336 VNB.n1409 VNB.n1408 0.136
R3337 VNB.n1410 VNB.n1409 0.136
R3338 VNB.n1411 VNB.n1410 0.136
R3339 VNB.n793 VNB 0.068
R3340 a_6049_1004.n8 a_6049_1004.t12 512.525
R3341 a_6049_1004.n6 a_6049_1004.t9 512.525
R3342 a_6049_1004.n8 a_6049_1004.t7 371.139
R3343 a_6049_1004.n6 a_6049_1004.t11 371.139
R3344 a_6049_1004.n11 a_6049_1004.n5 233.952
R3345 a_6049_1004.n9 a_6049_1004.n8 225.866
R3346 a_6049_1004.n7 a_6049_1004.n6 225.866
R3347 a_6049_1004.n9 a_6049_1004.t8 218.057
R3348 a_6049_1004.n7 a_6049_1004.t10 218.057
R3349 a_6049_1004.n13 a_6049_1004.n11 143.492
R3350 a_6049_1004.n10 a_6049_1004.n7 79.491
R3351 a_6049_1004.n4 a_6049_1004.n3 79.232
R3352 a_6049_1004.n11 a_6049_1004.n10 77.315
R3353 a_6049_1004.n10 a_6049_1004.n9 76
R3354 a_6049_1004.n5 a_6049_1004.n4 63.152
R3355 a_6049_1004.n13 a_6049_1004.n12 30
R3356 a_6049_1004.n14 a_6049_1004.n0 24.383
R3357 a_6049_1004.n14 a_6049_1004.n13 23.684
R3358 a_6049_1004.n5 a_6049_1004.n1 16.08
R3359 a_6049_1004.n4 a_6049_1004.n2 16.08
R3360 a_6049_1004.n1 a_6049_1004.t2 14.282
R3361 a_6049_1004.n1 a_6049_1004.t1 14.282
R3362 a_6049_1004.n2 a_6049_1004.t4 14.282
R3363 a_6049_1004.n2 a_6049_1004.t3 14.282
R3364 a_6049_1004.n3 a_6049_1004.t6 14.282
R3365 a_6049_1004.n3 a_6049_1004.t5 14.282
R3366 a_7973_1004.n6 a_7973_1004.t7 512.525
R3367 a_7973_1004.n6 a_7973_1004.t8 371.139
R3368 a_7973_1004.n8 a_7973_1004.n5 233.952
R3369 a_7973_1004.n7 a_7973_1004.n6 225.866
R3370 a_7973_1004.n7 a_7973_1004.t9 218.057
R3371 a_7973_1004.n8 a_7973_1004.n7 153.315
R3372 a_7973_1004.n10 a_7973_1004.n8 143.492
R3373 a_7973_1004.n4 a_7973_1004.n3 79.232
R3374 a_7973_1004.n5 a_7973_1004.n4 63.152
R3375 a_7973_1004.n10 a_7973_1004.n9 30
R3376 a_7973_1004.n11 a_7973_1004.n0 24.383
R3377 a_7973_1004.n11 a_7973_1004.n10 23.684
R3378 a_7973_1004.n5 a_7973_1004.n1 16.08
R3379 a_7973_1004.n4 a_7973_1004.n2 16.08
R3380 a_7973_1004.n1 a_7973_1004.t4 14.282
R3381 a_7973_1004.n1 a_7973_1004.t5 14.282
R3382 a_7973_1004.n2 a_7973_1004.t0 14.282
R3383 a_7973_1004.n2 a_7973_1004.t1 14.282
R3384 a_7973_1004.n3 a_7973_1004.t3 14.282
R3385 a_7973_1004.n3 a_7973_1004.t2 14.282
R3386 a_9897_1004.n10 a_9897_1004.t8 512.525
R3387 a_9897_1004.n5 a_9897_1004.t7 475.572
R3388 a_9897_1004.n7 a_9897_1004.t15 469.145
R3389 a_9897_1004.n7 a_9897_1004.t9 384.527
R3390 a_9897_1004.n5 a_9897_1004.t11 384.527
R3391 a_9897_1004.n10 a_9897_1004.t12 371.139
R3392 a_9897_1004.n8 a_9897_1004.t10 277.772
R3393 a_9897_1004.n6 a_9897_1004.t13 277.772
R3394 a_9897_1004.n11 a_9897_1004.t14 271.162
R3395 a_9897_1004.n15 a_9897_1004.n13 203.12
R3396 a_9897_1004.n13 a_9897_1004.n4 180.846
R3397 a_9897_1004.n11 a_9897_1004.n10 172.76
R3398 a_9897_1004.n9 a_9897_1004.n6 80.851
R3399 a_9897_1004.n3 a_9897_1004.n2 79.232
R3400 a_9897_1004.n13 a_9897_1004.n12 77.315
R3401 a_9897_1004.n9 a_9897_1004.n8 76
R3402 a_9897_1004.n12 a_9897_1004.n11 76
R3403 a_9897_1004.n6 a_9897_1004.n5 67.889
R3404 a_9897_1004.n8 a_9897_1004.n7 66.88
R3405 a_9897_1004.n4 a_9897_1004.n3 63.152
R3406 a_9897_1004.n12 a_9897_1004.n9 25.549
R3407 a_9897_1004.n4 a_9897_1004.n0 16.08
R3408 a_9897_1004.n3 a_9897_1004.n1 16.08
R3409 a_9897_1004.n15 a_9897_1004.n14 15.218
R3410 a_9897_1004.n0 a_9897_1004.t0 14.282
R3411 a_9897_1004.n0 a_9897_1004.t1 14.282
R3412 a_9897_1004.n1 a_9897_1004.t6 14.282
R3413 a_9897_1004.n1 a_9897_1004.t5 14.282
R3414 a_9897_1004.n2 a_9897_1004.t3 14.282
R3415 a_9897_1004.n2 a_9897_1004.t4 14.282
R3416 a_9897_1004.n16 a_9897_1004.n15 12.014
R3417 Q.n15 Q.n14 226.775
R3418 Q.n10 Q.n5 111.94
R3419 Q.n15 Q.n2 110.158
R3420 Q.n10 Q.n9 98.501
R3421 Q.n13 Q.n11 80.526
R3422 Q.n14 Q.n10 78.403
R3423 Q.n16 Q.n15 76
R3424 Q.n2 Q.n1 75.271
R3425 Q.n9 Q.n8 30
R3426 Q.n13 Q.n12 30
R3427 Q.n7 Q.n6 24.383
R3428 Q.n9 Q.n7 23.684
R3429 Q.n5 Q.n4 22.578
R3430 Q.n14 Q.n13 20.417
R3431 Q.n0 Q.t4 14.282
R3432 Q.n0 Q.t2 14.282
R3433 Q.n1 Q.t0 14.282
R3434 Q.n1 Q.t1 14.282
R3435 Q.n2 Q.n0 12.119
R3436 Q.n5 Q.n3 8.58
R3437 Q.n16 Q 0.046
R3438 a_18197_1005.n4 a_18197_1005.n3 196.002
R3439 a_18197_1005.t6 a_18197_1005.n5 89.556
R3440 a_18197_1005.n3 a_18197_1005.n2 75.271
R3441 a_18197_1005.n5 a_18197_1005.n4 75.214
R3442 a_18197_1005.n3 a_18197_1005.n1 36.52
R3443 a_18197_1005.n4 a_18197_1005.t4 14.338
R3444 a_18197_1005.n1 a_18197_1005.t0 14.282
R3445 a_18197_1005.n1 a_18197_1005.t7 14.282
R3446 a_18197_1005.n2 a_18197_1005.t1 14.282
R3447 a_18197_1005.n2 a_18197_1005.t3 14.282
R3448 a_18197_1005.n0 a_18197_1005.t5 14.282
R3449 a_18197_1005.n0 a_18197_1005.t2 14.282
R3450 a_18197_1005.n5 a_18197_1005.n0 12.119
R3451 a_4125_1004.n8 a_4125_1004.t7 512.525
R3452 a_4125_1004.n12 a_4125_1004.t10 512.525
R3453 a_4125_1004.n6 a_4125_1004.t13 477.179
R3454 a_4125_1004.n6 a_4125_1004.t9 406.485
R3455 a_4125_1004.n8 a_4125_1004.t8 371.139
R3456 a_4125_1004.n12 a_4125_1004.t14 371.139
R3457 a_4125_1004.n7 a_4125_1004.t12 346.633
R3458 a_4125_1004.n9 a_4125_1004.t15 340.206
R3459 a_4125_1004.n13 a_4125_1004.n12 225.866
R3460 a_4125_1004.n13 a_4125_1004.t11 218.057
R3461 a_4125_1004.n14 a_4125_1004.n11 159.317
R3462 a_4125_1004.n14 a_4125_1004.n13 153.315
R3463 a_4125_1004.n16 a_4125_1004.n14 143.492
R3464 a_4125_1004.n11 a_4125_1004.n10 123.155
R3465 a_4125_1004.n9 a_4125_1004.n8 89.615
R3466 a_4125_1004.n4 a_4125_1004.n3 79.232
R3467 a_4125_1004.n10 a_4125_1004.n7 78.675
R3468 a_4125_1004.n10 a_4125_1004.n9 76
R3469 a_4125_1004.n11 a_4125_1004.n5 74.634
R3470 a_4125_1004.n5 a_4125_1004.n4 63.152
R3471 a_4125_1004.n16 a_4125_1004.n15 30
R3472 a_4125_1004.n7 a_4125_1004.n6 29.194
R3473 a_4125_1004.n17 a_4125_1004.n0 24.383
R3474 a_4125_1004.n17 a_4125_1004.n16 23.684
R3475 a_4125_1004.n5 a_4125_1004.n1 16.08
R3476 a_4125_1004.n4 a_4125_1004.n2 16.08
R3477 a_4125_1004.n1 a_4125_1004.t2 14.282
R3478 a_4125_1004.n1 a_4125_1004.t3 14.282
R3479 a_4125_1004.n2 a_4125_1004.t5 14.282
R3480 a_4125_1004.n2 a_4125_1004.t6 14.282
R3481 a_4125_1004.n3 a_4125_1004.t4 14.282
R3482 a_4125_1004.n3 a_4125_1004.t0 14.282
R3483 a_17533_1005.n4 a_17533_1005.n3 195.987
R3484 a_17533_1005.n2 a_17533_1005.t0 89.553
R3485 a_17533_1005.n5 a_17533_1005.n4 75.27
R3486 a_17533_1005.n3 a_17533_1005.n2 75.214
R3487 a_17533_1005.n4 a_17533_1005.n0 36.519
R3488 a_17533_1005.n3 a_17533_1005.t4 14.338
R3489 a_17533_1005.n0 a_17533_1005.t5 14.282
R3490 a_17533_1005.n0 a_17533_1005.t6 14.282
R3491 a_17533_1005.n1 a_17533_1005.t7 14.282
R3492 a_17533_1005.n1 a_17533_1005.t3 14.282
R3493 a_17533_1005.t2 a_17533_1005.n5 14.282
R3494 a_17533_1005.n5 a_17533_1005.t1 14.282
R3495 a_17533_1005.n2 a_17533_1005.n1 12.119
R3496 a_14521_75.n1 a_14521_75.n0 25.576
R3497 a_14521_75.n3 a_14521_75.n2 9.111
R3498 a_14521_75.n7 a_14521_75.n5 7.859
R3499 a_14521_75.t0 a_14521_75.n7 3.034
R3500 a_14521_75.n5 a_14521_75.n3 1.964
R3501 a_14521_75.n5 a_14521_75.n4 1.964
R3502 a_14521_75.t0 a_14521_75.n1 1.871
R3503 a_14521_75.n7 a_14521_75.n6 0.443
R3504 a_14802_182.n12 a_14802_182.n10 82.852
R3505 a_14802_182.n13 a_14802_182.n0 49.6
R3506 a_14802_182.t1 a_14802_182.n2 46.91
R3507 a_14802_182.n7 a_14802_182.n5 34.805
R3508 a_14802_182.n7 a_14802_182.n6 32.622
R3509 a_14802_182.n10 a_14802_182.t1 32.416
R3510 a_14802_182.n12 a_14802_182.n11 27.2
R3511 a_14802_182.n13 a_14802_182.n12 22.4
R3512 a_14802_182.n9 a_14802_182.n7 19.017
R3513 a_14802_182.n2 a_14802_182.n1 17.006
R3514 a_14802_182.n5 a_14802_182.n4 7.5
R3515 a_14802_182.n9 a_14802_182.n8 7.5
R3516 a_14802_182.t1 a_14802_182.n3 7.04
R3517 a_14802_182.n10 a_14802_182.n9 1.435
R3518 a_277_1004.n7 a_277_1004.t10 512.525
R3519 a_277_1004.n5 a_277_1004.t7 512.525
R3520 a_277_1004.n7 a_277_1004.t11 371.139
R3521 a_277_1004.n5 a_277_1004.t12 371.139
R3522 a_277_1004.n10 a_277_1004.n4 233.952
R3523 a_277_1004.n8 a_277_1004.n7 225.866
R3524 a_277_1004.n6 a_277_1004.n5 225.866
R3525 a_277_1004.n8 a_277_1004.t9 218.057
R3526 a_277_1004.n6 a_277_1004.t8 218.057
R3527 a_277_1004.n12 a_277_1004.n10 150.014
R3528 a_277_1004.n9 a_277_1004.n6 79.491
R3529 a_277_1004.n3 a_277_1004.n2 79.232
R3530 a_277_1004.n10 a_277_1004.n9 77.315
R3531 a_277_1004.n9 a_277_1004.n8 76
R3532 a_277_1004.n4 a_277_1004.n3 63.152
R3533 a_277_1004.n4 a_277_1004.n0 16.08
R3534 a_277_1004.n3 a_277_1004.n1 16.08
R3535 a_277_1004.n12 a_277_1004.n11 15.218
R3536 a_277_1004.n0 a_277_1004.t1 14.282
R3537 a_277_1004.n0 a_277_1004.t2 14.282
R3538 a_277_1004.n1 a_277_1004.t4 14.282
R3539 a_277_1004.n1 a_277_1004.t3 14.282
R3540 a_277_1004.n2 a_277_1004.t6 14.282
R3541 a_277_1004.n2 a_277_1004.t5 14.282
R3542 a_277_1004.n13 a_277_1004.n12 12.014
R3543 a_11821_1004.n8 a_11821_1004.t10 512.525
R3544 a_11821_1004.n6 a_11821_1004.t8 512.525
R3545 a_11821_1004.n8 a_11821_1004.t7 371.139
R3546 a_11821_1004.n6 a_11821_1004.t11 371.139
R3547 a_11821_1004.n11 a_11821_1004.n5 233.952
R3548 a_11821_1004.n9 a_11821_1004.n8 225.866
R3549 a_11821_1004.n7 a_11821_1004.n6 225.866
R3550 a_11821_1004.n9 a_11821_1004.t9 218.057
R3551 a_11821_1004.n7 a_11821_1004.t12 218.057
R3552 a_11821_1004.n13 a_11821_1004.n11 143.492
R3553 a_11821_1004.n10 a_11821_1004.n7 79.491
R3554 a_11821_1004.n4 a_11821_1004.n3 79.232
R3555 a_11821_1004.n11 a_11821_1004.n10 77.315
R3556 a_11821_1004.n10 a_11821_1004.n9 76
R3557 a_11821_1004.n5 a_11821_1004.n4 63.152
R3558 a_11821_1004.n13 a_11821_1004.n12 30
R3559 a_11821_1004.n14 a_11821_1004.n0 24.383
R3560 a_11821_1004.n14 a_11821_1004.n13 23.684
R3561 a_11821_1004.n5 a_11821_1004.n1 16.08
R3562 a_11821_1004.n4 a_11821_1004.n2 16.08
R3563 a_11821_1004.n1 a_11821_1004.t5 14.282
R3564 a_11821_1004.n1 a_11821_1004.t6 14.282
R3565 a_11821_1004.n2 a_11821_1004.t1 14.282
R3566 a_11821_1004.n2 a_11821_1004.t0 14.282
R3567 a_11821_1004.n3 a_11821_1004.t3 14.282
R3568 a_11821_1004.n3 a_11821_1004.t2 14.282
R3569 a_15669_1004.n11 a_15669_1004.t13 512.525
R3570 a_15669_1004.n8 a_15669_1004.t10 512.525
R3571 a_15669_1004.n6 a_15669_1004.t11 512.525
R3572 a_15669_1004.n11 a_15669_1004.t9 371.139
R3573 a_15669_1004.n8 a_15669_1004.t15 371.139
R3574 a_15669_1004.n6 a_15669_1004.t14 371.139
R3575 a_15669_1004.n14 a_15669_1004.n5 260.505
R3576 a_15669_1004.n9 a_15669_1004.n8 258.98
R3577 a_15669_1004.n7 a_15669_1004.n6 258.98
R3578 a_15669_1004.n12 a_15669_1004.n11 253.685
R3579 a_15669_1004.n12 a_15669_1004.t8 179.042
R3580 a_15669_1004.n7 a_15669_1004.t12 176.995
R3581 a_15669_1004.n9 a_15669_1004.t7 170.569
R3582 a_15669_1004.n16 a_15669_1004.n14 116.939
R3583 a_15669_1004.n4 a_15669_1004.n3 79.232
R3584 a_15669_1004.n14 a_15669_1004.n13 77.315
R3585 a_15669_1004.n10 a_15669_1004.n7 77.027
R3586 a_15669_1004.n10 a_15669_1004.n9 76
R3587 a_15669_1004.n5 a_15669_1004.n4 63.152
R3588 a_15669_1004.n13 a_15669_1004.n12 49.344
R3589 a_15669_1004.n16 a_15669_1004.n15 30
R3590 a_15669_1004.n17 a_15669_1004.n0 24.383
R3591 a_15669_1004.n17 a_15669_1004.n16 23.684
R3592 a_15669_1004.n5 a_15669_1004.n1 16.08
R3593 a_15669_1004.n4 a_15669_1004.n2 16.08
R3594 a_15669_1004.n1 a_15669_1004.t2 14.282
R3595 a_15669_1004.n1 a_15669_1004.t6 14.282
R3596 a_15669_1004.n2 a_15669_1004.t1 14.282
R3597 a_15669_1004.n2 a_15669_1004.t0 14.282
R3598 a_15669_1004.n3 a_15669_1004.t4 14.282
R3599 a_15669_1004.n3 a_15669_1004.t5 14.282
R3600 a_15669_1004.n13 a_15669_1004.n10 7.002
R3601 a_18094_73.n2 a_18094_73.n0 34.602
R3602 a_18094_73.n2 a_18094_73.n1 2.138
R3603 a_18094_73.t0 a_18094_73.n2 0.069
R3604 a_16445_75.n1 a_16445_75.n0 25.576
R3605 a_16445_75.n3 a_16445_75.n2 9.111
R3606 a_16445_75.n7 a_16445_75.n5 7.859
R3607 a_16445_75.t0 a_16445_75.n7 3.034
R3608 a_16445_75.n5 a_16445_75.n3 1.964
R3609 a_16445_75.n5 a_16445_75.n4 1.964
R3610 a_16445_75.t0 a_16445_75.n1 1.871
R3611 a_16445_75.n7 a_16445_75.n6 0.443
R3612 a_16726_182.n8 a_16726_182.n6 96.467
R3613 a_16726_182.n3 a_16726_182.n1 44.628
R3614 a_16726_182.t0 a_16726_182.n8 32.417
R3615 a_16726_182.n3 a_16726_182.n2 23.284
R3616 a_16726_182.n6 a_16726_182.n5 22.349
R3617 a_16726_182.t0 a_16726_182.n10 20.241
R3618 a_16726_182.n10 a_16726_182.n9 13.494
R3619 a_16726_182.n6 a_16726_182.n4 8.443
R3620 a_16726_182.t0 a_16726_182.n0 8.137
R3621 a_16726_182.t0 a_16726_182.n3 5.727
R3622 a_16726_182.n8 a_16726_182.n7 1.435
R3623 a_10673_75.n1 a_10673_75.n0 25.576
R3624 a_10673_75.n3 a_10673_75.n2 9.111
R3625 a_10673_75.n7 a_10673_75.n5 7.859
R3626 a_10673_75.t0 a_10673_75.n7 3.034
R3627 a_10673_75.n5 a_10673_75.n3 1.964
R3628 a_10673_75.n5 a_10673_75.n4 1.964
R3629 a_10673_75.t0 a_10673_75.n1 1.871
R3630 a_10673_75.n7 a_10673_75.n6 0.443
R3631 a_10954_182.n12 a_10954_182.n10 82.852
R3632 a_10954_182.n13 a_10954_182.n0 49.6
R3633 a_10954_182.t1 a_10954_182.n2 46.91
R3634 a_10954_182.n7 a_10954_182.n5 34.805
R3635 a_10954_182.n7 a_10954_182.n6 32.622
R3636 a_10954_182.n10 a_10954_182.t1 32.416
R3637 a_10954_182.n12 a_10954_182.n11 27.2
R3638 a_10954_182.n13 a_10954_182.n12 22.4
R3639 a_10954_182.n9 a_10954_182.n7 19.017
R3640 a_10954_182.n2 a_10954_182.n1 17.006
R3641 a_10954_182.n5 a_10954_182.n4 7.5
R3642 a_10954_182.n9 a_10954_182.n8 7.5
R3643 a_10954_182.t1 a_10954_182.n3 7.04
R3644 a_10954_182.n10 a_10954_182.n9 1.435
R3645 a_12597_75.n1 a_12597_75.n0 25.576
R3646 a_12597_75.n3 a_12597_75.n2 9.111
R3647 a_12597_75.n7 a_12597_75.n5 7.859
R3648 a_12597_75.t0 a_12597_75.n7 3.034
R3649 a_12597_75.n5 a_12597_75.n3 1.964
R3650 a_12597_75.n5 a_12597_75.n4 1.964
R3651 a_12597_75.t0 a_12597_75.n1 1.871
R3652 a_12597_75.n7 a_12597_75.n6 0.443
R3653 a_12878_182.n8 a_12878_182.n6 96.467
R3654 a_12878_182.n3 a_12878_182.n1 44.628
R3655 a_12878_182.t0 a_12878_182.n8 32.417
R3656 a_12878_182.n3 a_12878_182.n2 23.284
R3657 a_12878_182.n6 a_12878_182.n5 22.349
R3658 a_12878_182.t0 a_12878_182.n10 20.241
R3659 a_12878_182.n10 a_12878_182.n9 13.494
R3660 a_12878_182.n6 a_12878_182.n4 8.443
R3661 a_12878_182.t0 a_12878_182.n0 8.137
R3662 a_12878_182.t0 a_12878_182.n3 5.727
R3663 a_12878_182.n8 a_12878_182.n7 1.435
R3664 a_599_943.n5 a_599_943.t12 512.525
R3665 a_599_943.n7 a_599_943.t10 454.685
R3666 a_599_943.n7 a_599_943.t8 428.979
R3667 a_599_943.n5 a_599_943.t7 371.139
R3668 a_599_943.n6 a_599_943.t9 271.162
R3669 a_599_943.n8 a_599_943.t11 221.453
R3670 a_599_943.n12 a_599_943.n10 203.12
R3671 a_599_943.n10 a_599_943.n4 180.846
R3672 a_599_943.n6 a_599_943.n5 172.76
R3673 a_599_943.n8 a_599_943.n7 108.494
R3674 a_599_943.n9 a_599_943.n6 84.388
R3675 a_599_943.n9 a_599_943.n8 80.035
R3676 a_599_943.n3 a_599_943.n2 79.232
R3677 a_599_943.n10 a_599_943.n9 76
R3678 a_599_943.n4 a_599_943.n3 63.152
R3679 a_599_943.n4 a_599_943.n0 16.08
R3680 a_599_943.n3 a_599_943.n1 16.08
R3681 a_599_943.n12 a_599_943.n11 15.218
R3682 a_599_943.n0 a_599_943.t5 14.282
R3683 a_599_943.n0 a_599_943.t6 14.282
R3684 a_599_943.n1 a_599_943.t1 14.282
R3685 a_599_943.n1 a_599_943.t2 14.282
R3686 a_599_943.n2 a_599_943.t4 14.282
R3687 a_599_943.n2 a_599_943.t3 14.282
R3688 a_599_943.n13 a_599_943.n12 12.014
R3689 a_1561_943.n8 a_1561_943.t14 454.685
R3690 a_1561_943.n10 a_1561_943.t8 454.685
R3691 a_1561_943.n6 a_1561_943.t15 454.685
R3692 a_1561_943.n8 a_1561_943.t11 428.979
R3693 a_1561_943.n10 a_1561_943.t12 428.979
R3694 a_1561_943.n6 a_1561_943.t13 428.979
R3695 a_1561_943.n9 a_1561_943.t7 248.006
R3696 a_1561_943.n11 a_1561_943.t9 248.006
R3697 a_1561_943.n7 a_1561_943.t10 248.006
R3698 a_1561_943.n16 a_1561_943.n14 223.151
R3699 a_1561_943.n14 a_1561_943.n5 154.293
R3700 a_1561_943.n13 a_1561_943.n7 82.484
R3701 a_1561_943.n9 a_1561_943.n8 81.941
R3702 a_1561_943.n11 a_1561_943.n10 81.941
R3703 a_1561_943.n7 a_1561_943.n6 81.941
R3704 a_1561_943.n12 a_1561_943.n11 79.491
R3705 a_1561_943.n4 a_1561_943.n3 79.232
R3706 a_1561_943.n12 a_1561_943.n9 76
R3707 a_1561_943.n14 a_1561_943.n13 76
R3708 a_1561_943.n5 a_1561_943.n4 63.152
R3709 a_1561_943.n16 a_1561_943.n15 30
R3710 a_1561_943.n17 a_1561_943.n0 24.383
R3711 a_1561_943.n17 a_1561_943.n16 23.684
R3712 a_1561_943.n5 a_1561_943.n1 16.08
R3713 a_1561_943.n4 a_1561_943.n2 16.08
R3714 a_1561_943.n1 a_1561_943.t6 14.282
R3715 a_1561_943.n1 a_1561_943.t5 14.282
R3716 a_1561_943.n2 a_1561_943.t3 14.282
R3717 a_1561_943.n2 a_1561_943.t2 14.282
R3718 a_1561_943.n3 a_1561_943.t0 14.282
R3719 a_1561_943.n3 a_1561_943.t1 14.282
R3720 a_1561_943.n13 a_1561_943.n12 4.035
R3721 a_2296_182.n12 a_2296_182.n10 82.852
R3722 a_2296_182.t1 a_2296_182.n2 46.91
R3723 a_2296_182.n7 a_2296_182.n5 34.805
R3724 a_2296_182.n7 a_2296_182.n6 32.622
R3725 a_2296_182.n10 a_2296_182.t1 32.416
R3726 a_2296_182.n12 a_2296_182.n11 27.2
R3727 a_2296_182.n13 a_2296_182.n0 23.498
R3728 a_2296_182.n13 a_2296_182.n12 22.4
R3729 a_2296_182.n9 a_2296_182.n7 19.017
R3730 a_2296_182.n2 a_2296_182.n1 17.006
R3731 a_2296_182.n5 a_2296_182.n4 7.5
R3732 a_2296_182.n9 a_2296_182.n8 7.5
R3733 a_2296_182.t1 a_2296_182.n3 7.04
R3734 a_2296_182.n10 a_2296_182.n9 1.435
R3735 a_2201_1004.n5 a_2201_1004.t9 512.525
R3736 a_2201_1004.n5 a_2201_1004.t8 371.139
R3737 a_2201_1004.n7 a_2201_1004.n4 233.952
R3738 a_2201_1004.n6 a_2201_1004.n5 225.866
R3739 a_2201_1004.n6 a_2201_1004.t7 218.057
R3740 a_2201_1004.n7 a_2201_1004.n6 153.315
R3741 a_2201_1004.n9 a_2201_1004.n7 150.014
R3742 a_2201_1004.n3 a_2201_1004.n2 79.232
R3743 a_2201_1004.n4 a_2201_1004.n3 63.152
R3744 a_2201_1004.n4 a_2201_1004.n0 16.08
R3745 a_2201_1004.n3 a_2201_1004.n1 16.08
R3746 a_2201_1004.n9 a_2201_1004.n8 15.218
R3747 a_2201_1004.n0 a_2201_1004.t6 14.282
R3748 a_2201_1004.n0 a_2201_1004.t5 14.282
R3749 a_2201_1004.n1 a_2201_1004.t1 14.282
R3750 a_2201_1004.n1 a_2201_1004.t0 14.282
R3751 a_2201_1004.n2 a_2201_1004.t3 14.282
R3752 a_2201_1004.n2 a_2201_1004.t2 14.282
R3753 a_2201_1004.n10 a_2201_1004.n9 12.014
R3754 a_91_75.n1 a_91_75.n0 25.576
R3755 a_91_75.n3 a_91_75.n2 9.111
R3756 a_91_75.n7 a_91_75.n5 7.859
R3757 a_91_75.t0 a_91_75.n7 3.034
R3758 a_91_75.n5 a_91_75.n3 1.964
R3759 a_91_75.n5 a_91_75.n4 1.964
R3760 a_91_75.t0 a_91_75.n1 1.871
R3761 a_91_75.n7 a_91_75.n6 0.443
R3762 a_372_182.n8 a_372_182.n6 96.467
R3763 a_372_182.n3 a_372_182.n1 44.628
R3764 a_372_182.t0 a_372_182.n8 32.417
R3765 a_372_182.n3 a_372_182.n2 23.284
R3766 a_372_182.n6 a_372_182.n5 22.349
R3767 a_372_182.t0 a_372_182.n10 20.241
R3768 a_372_182.n10 a_372_182.n9 13.494
R3769 a_372_182.n6 a_372_182.n4 8.443
R3770 a_372_182.t0 a_372_182.n0 8.137
R3771 a_372_182.t0 a_372_182.n3 5.727
R3772 a_372_182.n8 a_372_182.n7 1.435
R3773 a_13105_943.n7 a_13105_943.t12 454.685
R3774 a_13105_943.n9 a_13105_943.t14 454.685
R3775 a_13105_943.n5 a_13105_943.t10 454.685
R3776 a_13105_943.n7 a_13105_943.t7 428.979
R3777 a_13105_943.n9 a_13105_943.t11 428.979
R3778 a_13105_943.n5 a_13105_943.t8 428.979
R3779 a_13105_943.n8 a_13105_943.t13 248.006
R3780 a_13105_943.n10 a_13105_943.t9 248.006
R3781 a_13105_943.n6 a_13105_943.t15 248.006
R3782 a_13105_943.n15 a_13105_943.n13 229.673
R3783 a_13105_943.n13 a_13105_943.n4 154.293
R3784 a_13105_943.n12 a_13105_943.n6 82.484
R3785 a_13105_943.n8 a_13105_943.n7 81.941
R3786 a_13105_943.n10 a_13105_943.n9 81.941
R3787 a_13105_943.n6 a_13105_943.n5 81.941
R3788 a_13105_943.n11 a_13105_943.n10 79.491
R3789 a_13105_943.n3 a_13105_943.n2 79.232
R3790 a_13105_943.n11 a_13105_943.n8 76
R3791 a_13105_943.n13 a_13105_943.n12 76
R3792 a_13105_943.n4 a_13105_943.n3 63.152
R3793 a_13105_943.n4 a_13105_943.n0 16.08
R3794 a_13105_943.n3 a_13105_943.n1 16.08
R3795 a_13105_943.n15 a_13105_943.n14 15.218
R3796 a_13105_943.n0 a_13105_943.t5 14.282
R3797 a_13105_943.n0 a_13105_943.t6 14.282
R3798 a_13105_943.n1 a_13105_943.t3 14.282
R3799 a_13105_943.n1 a_13105_943.t2 14.282
R3800 a_13105_943.n2 a_13105_943.t0 14.282
R3801 a_13105_943.n2 a_13105_943.t1 14.282
R3802 a_13105_943.n16 a_13105_943.n15 12.014
R3803 a_13105_943.n12 a_13105_943.n11 4.035
R3804 a_13745_1004.n6 a_13745_1004.t7 512.525
R3805 a_13745_1004.n6 a_13745_1004.t8 371.139
R3806 a_13745_1004.n8 a_13745_1004.n5 233.952
R3807 a_13745_1004.n7 a_13745_1004.n6 225.866
R3808 a_13745_1004.n7 a_13745_1004.t9 218.057
R3809 a_13745_1004.n8 a_13745_1004.n7 153.315
R3810 a_13745_1004.n10 a_13745_1004.n8 143.492
R3811 a_13745_1004.n4 a_13745_1004.n3 79.232
R3812 a_13745_1004.n5 a_13745_1004.n4 63.152
R3813 a_13745_1004.n10 a_13745_1004.n9 30
R3814 a_13745_1004.n11 a_13745_1004.n0 24.383
R3815 a_13745_1004.n11 a_13745_1004.n10 23.684
R3816 a_13745_1004.n5 a_13745_1004.n1 16.08
R3817 a_13745_1004.n4 a_13745_1004.n2 16.08
R3818 a_13745_1004.n1 a_13745_1004.t5 14.282
R3819 a_13745_1004.n1 a_13745_1004.t4 14.282
R3820 a_13745_1004.n2 a_13745_1004.t0 14.282
R3821 a_13745_1004.n2 a_13745_1004.t1 14.282
R3822 a_13745_1004.n3 a_13745_1004.t3 14.282
R3823 a_13745_1004.n3 a_13745_1004.t2 14.282
R3824 a_10219_943.n5 a_10219_943.t8 454.685
R3825 a_10219_943.n5 a_10219_943.t9 428.979
R3826 a_10219_943.n7 a_10219_943.n4 233.952
R3827 a_10219_943.n6 a_10219_943.t7 168.348
R3828 a_10219_943.n6 a_10219_943.n5 161.6
R3829 a_10219_943.n7 a_10219_943.n6 156.035
R3830 a_10219_943.n9 a_10219_943.n7 150.014
R3831 a_10219_943.n3 a_10219_943.n2 79.232
R3832 a_10219_943.n4 a_10219_943.n3 63.152
R3833 a_10219_943.n4 a_10219_943.n0 16.08
R3834 a_10219_943.n3 a_10219_943.n1 16.08
R3835 a_10219_943.n9 a_10219_943.n8 15.218
R3836 a_10219_943.n0 a_10219_943.t5 14.282
R3837 a_10219_943.n0 a_10219_943.t6 14.282
R3838 a_10219_943.n1 a_10219_943.t0 14.282
R3839 a_10219_943.n1 a_10219_943.t1 14.282
R3840 a_10219_943.n2 a_10219_943.t3 14.282
R3841 a_10219_943.n2 a_10219_943.t2 14.282
R3842 a_10219_943.n10 a_10219_943.n9 12.014
R3843 a_4220_182.n9 a_4220_182.n7 82.852
R3844 a_4220_182.n3 a_4220_182.n1 44.628
R3845 a_4220_182.t0 a_4220_182.n9 32.417
R3846 a_4220_182.n7 a_4220_182.n6 27.2
R3847 a_4220_182.n5 a_4220_182.n4 23.498
R3848 a_4220_182.n3 a_4220_182.n2 23.284
R3849 a_4220_182.n7 a_4220_182.n5 22.4
R3850 a_4220_182.t0 a_4220_182.n11 20.241
R3851 a_4220_182.n11 a_4220_182.n10 13.494
R3852 a_4220_182.t0 a_4220_182.n0 8.137
R3853 a_4220_182.t0 a_4220_182.n3 5.727
R3854 a_4220_182.n9 a_4220_182.n8 1.435
R3855 a_13559_75.n1 a_13559_75.n0 25.576
R3856 a_13559_75.n3 a_13559_75.n2 9.111
R3857 a_13559_75.n7 a_13559_75.n5 7.859
R3858 a_13559_75.t0 a_13559_75.n7 3.034
R3859 a_13559_75.n5 a_13559_75.n3 1.964
R3860 a_13559_75.n5 a_13559_75.n4 1.964
R3861 a_13559_75.t0 a_13559_75.n1 1.871
R3862 a_13559_75.n7 a_13559_75.n6 0.443
R3863 a_13840_182.n10 a_13840_182.n8 82.852
R3864 a_13840_182.n11 a_13840_182.n0 49.6
R3865 a_13840_182.n7 a_13840_182.n6 32.833
R3866 a_13840_182.n8 a_13840_182.t1 32.416
R3867 a_13840_182.n10 a_13840_182.n9 27.2
R3868 a_13840_182.n3 a_13840_182.n2 23.284
R3869 a_13840_182.n11 a_13840_182.n10 22.4
R3870 a_13840_182.n7 a_13840_182.n4 19.017
R3871 a_13840_182.n6 a_13840_182.n5 13.494
R3872 a_13840_182.t1 a_13840_182.n1 7.04
R3873 a_13840_182.t1 a_13840_182.n3 5.727
R3874 a_13840_182.n8 a_13840_182.n7 1.435
R3875 a_15764_182.n10 a_15764_182.n8 82.852
R3876 a_15764_182.n11 a_15764_182.n0 49.6
R3877 a_15764_182.n7 a_15764_182.n6 32.833
R3878 a_15764_182.n8 a_15764_182.t1 32.416
R3879 a_15764_182.n10 a_15764_182.n9 27.2
R3880 a_15764_182.n3 a_15764_182.n2 23.284
R3881 a_15764_182.n11 a_15764_182.n10 22.4
R3882 a_15764_182.n7 a_15764_182.n4 19.017
R3883 a_15764_182.n6 a_15764_182.n5 13.494
R3884 a_15764_182.t1 a_15764_182.n1 7.04
R3885 a_15764_182.t1 a_15764_182.n3 5.727
R3886 a_15764_182.n8 a_15764_182.n7 1.435
R3887 a_7106_182.n10 a_7106_182.n8 82.852
R3888 a_7106_182.n7 a_7106_182.n6 32.833
R3889 a_7106_182.n8 a_7106_182.t1 32.416
R3890 a_7106_182.n10 a_7106_182.n9 27.2
R3891 a_7106_182.n11 a_7106_182.n0 23.498
R3892 a_7106_182.n3 a_7106_182.n2 23.284
R3893 a_7106_182.n11 a_7106_182.n10 22.4
R3894 a_7106_182.n7 a_7106_182.n4 19.017
R3895 a_7106_182.n6 a_7106_182.n5 13.494
R3896 a_7106_182.t1 a_7106_182.n1 7.04
R3897 a_7106_182.t1 a_7106_182.n3 5.727
R3898 a_7106_182.n8 a_7106_182.n7 1.435
R3899 a_2015_75.n1 a_2015_75.n0 25.576
R3900 a_2015_75.n3 a_2015_75.n2 9.111
R3901 a_2015_75.n7 a_2015_75.n6 2.455
R3902 a_2015_75.n5 a_2015_75.n3 1.964
R3903 a_2015_75.n5 a_2015_75.n4 1.964
R3904 a_2015_75.t0 a_2015_75.n1 1.871
R3905 a_2015_75.n7 a_2015_75.n5 0.636
R3906 a_2015_75.t0 a_2015_75.n7 0.246
R3907 a_1334_182.n10 a_1334_182.n8 82.852
R3908 a_1334_182.n7 a_1334_182.n6 32.833
R3909 a_1334_182.n8 a_1334_182.t1 32.416
R3910 a_1334_182.n10 a_1334_182.n9 27.2
R3911 a_1334_182.n11 a_1334_182.n0 23.498
R3912 a_1334_182.n3 a_1334_182.n2 23.284
R3913 a_1334_182.n11 a_1334_182.n10 22.4
R3914 a_1334_182.n7 a_1334_182.n4 19.017
R3915 a_1334_182.n6 a_1334_182.n5 13.494
R3916 a_1334_182.t1 a_1334_182.n1 7.04
R3917 a_1334_182.t1 a_1334_182.n3 5.727
R3918 a_1334_182.n8 a_1334_182.n7 1.435
R3919 a_15991_943.n5 a_15991_943.t9 454.685
R3920 a_15991_943.n5 a_15991_943.t7 428.979
R3921 a_15991_943.n7 a_15991_943.n4 233.952
R3922 a_15991_943.n6 a_15991_943.t8 168.348
R3923 a_15991_943.n6 a_15991_943.n5 161.6
R3924 a_15991_943.n7 a_15991_943.n6 156.035
R3925 a_15991_943.n9 a_15991_943.n7 150.014
R3926 a_15991_943.n3 a_15991_943.n2 79.232
R3927 a_15991_943.n4 a_15991_943.n3 63.152
R3928 a_15991_943.n4 a_15991_943.n0 16.08
R3929 a_15991_943.n3 a_15991_943.n1 16.08
R3930 a_15991_943.n9 a_15991_943.n8 15.218
R3931 a_15991_943.n0 a_15991_943.t6 14.282
R3932 a_15991_943.n0 a_15991_943.t5 14.282
R3933 a_15991_943.n1 a_15991_943.t0 14.282
R3934 a_15991_943.n1 a_15991_943.t1 14.282
R3935 a_15991_943.n2 a_15991_943.t2 14.282
R3936 a_15991_943.n2 a_15991_943.t3 14.282
R3937 a_15991_943.n10 a_15991_943.n9 12.014
R3938 a_3258_182.n10 a_3258_182.n8 82.852
R3939 a_3258_182.n7 a_3258_182.n6 32.833
R3940 a_3258_182.n8 a_3258_182.t1 32.416
R3941 a_3258_182.n10 a_3258_182.n9 27.2
R3942 a_3258_182.n11 a_3258_182.n0 23.498
R3943 a_3258_182.n3 a_3258_182.n2 23.284
R3944 a_3258_182.n11 a_3258_182.n10 22.4
R3945 a_3258_182.n7 a_3258_182.n4 19.017
R3946 a_3258_182.n6 a_3258_182.n5 13.494
R3947 a_3258_182.t1 a_3258_182.n1 7.04
R3948 a_3258_182.t1 a_3258_182.n3 5.727
R3949 a_3258_182.n8 a_3258_182.n7 1.435
R3950 a_5182_182.n10 a_5182_182.n8 82.852
R3951 a_5182_182.n7 a_5182_182.n6 32.833
R3952 a_5182_182.n8 a_5182_182.t1 32.416
R3953 a_5182_182.n10 a_5182_182.n9 27.2
R3954 a_5182_182.n11 a_5182_182.n0 23.498
R3955 a_5182_182.n3 a_5182_182.n2 23.284
R3956 a_5182_182.n11 a_5182_182.n10 22.4
R3957 a_5182_182.n7 a_5182_182.n4 19.017
R3958 a_5182_182.n6 a_5182_182.n5 13.494
R3959 a_5182_182.t1 a_5182_182.n1 7.04
R3960 a_5182_182.t1 a_5182_182.n3 5.727
R3961 a_5182_182.n8 a_5182_182.n7 1.435
R3962 a_11916_182.n10 a_11916_182.n8 82.852
R3963 a_11916_182.n7 a_11916_182.n6 32.833
R3964 a_11916_182.n8 a_11916_182.t1 32.416
R3965 a_11916_182.n10 a_11916_182.n9 27.2
R3966 a_11916_182.n11 a_11916_182.n0 23.498
R3967 a_11916_182.n3 a_11916_182.n2 23.284
R3968 a_11916_182.n11 a_11916_182.n10 22.4
R3969 a_11916_182.n7 a_11916_182.n4 19.017
R3970 a_11916_182.n6 a_11916_182.n5 13.494
R3971 a_11916_182.t1 a_11916_182.n1 7.04
R3972 a_11916_182.t1 a_11916_182.n3 5.727
R3973 a_11916_182.n8 a_11916_182.n7 1.435
R3974 a_17428_73.n13 a_17428_73.n12 26.811
R3975 a_17428_73.n6 a_17428_73.n5 24.977
R3976 a_17428_73.n2 a_17428_73.n1 24.877
R3977 a_17428_73.t0 a_17428_73.n2 12.677
R3978 a_17428_73.t0 a_17428_73.n3 11.595
R3979 a_17428_73.n11 a_17428_73.n10 8.561
R3980 a_17428_73.t0 a_17428_73.n4 7.273
R3981 a_17428_73.n9 a_17428_73.n8 7.066
R3982 a_17428_73.t0 a_17428_73.n0 6.109
R3983 a_17428_73.t1 a_17428_73.n7 4.864
R3984 a_17428_73.t0 a_17428_73.n13 2.074
R3985 a_17428_73.n7 a_17428_73.n6 1.13
R3986 a_17428_73.t1 a_17428_73.n11 0.958
R3987 a_17428_73.n13 a_17428_73.t1 0.937
R3988 a_17428_73.t1 a_17428_73.n9 0.86
R3989 a_9992_182.n9 a_9992_182.n7 82.852
R3990 a_9992_182.n3 a_9992_182.n1 44.628
R3991 a_9992_182.t0 a_9992_182.n9 32.417
R3992 a_9992_182.n7 a_9992_182.n6 27.2
R3993 a_9992_182.n5 a_9992_182.n4 23.498
R3994 a_9992_182.n3 a_9992_182.n2 23.284
R3995 a_9992_182.n7 a_9992_182.n5 22.4
R3996 a_9992_182.t0 a_9992_182.n11 20.241
R3997 a_9992_182.n11 a_9992_182.n10 13.494
R3998 a_9992_182.t0 a_9992_182.n0 8.137
R3999 a_9992_182.t0 a_9992_182.n3 5.727
R4000 a_9992_182.n9 a_9992_182.n8 1.435
R4001 a_6144_182.n9 a_6144_182.n7 82.852
R4002 a_6144_182.n3 a_6144_182.n1 44.628
R4003 a_6144_182.t0 a_6144_182.n9 32.417
R4004 a_6144_182.n7 a_6144_182.n6 27.2
R4005 a_6144_182.n5 a_6144_182.n4 23.498
R4006 a_6144_182.n3 a_6144_182.n2 23.284
R4007 a_6144_182.n7 a_6144_182.n5 22.4
R4008 a_6144_182.t0 a_6144_182.n11 20.241
R4009 a_6144_182.n11 a_6144_182.n10 13.494
R4010 a_6144_182.t0 a_6144_182.n0 8.137
R4011 a_6144_182.t0 a_6144_182.n3 5.727
R4012 a_6144_182.n9 a_6144_182.n8 1.435
R4013 a_8068_182.n10 a_8068_182.n8 82.852
R4014 a_8068_182.n7 a_8068_182.n6 32.833
R4015 a_8068_182.n8 a_8068_182.t1 32.416
R4016 a_8068_182.n10 a_8068_182.n9 27.2
R4017 a_8068_182.n11 a_8068_182.n0 23.498
R4018 a_8068_182.n3 a_8068_182.n2 23.284
R4019 a_8068_182.n11 a_8068_182.n10 22.4
R4020 a_8068_182.n7 a_8068_182.n4 19.017
R4021 a_8068_182.n6 a_8068_182.n5 13.494
R4022 a_8068_182.t1 a_8068_182.n1 7.04
R4023 a_8068_182.t1 a_8068_182.n3 5.727
R4024 a_8068_182.n8 a_8068_182.n7 1.435
R4025 a_2977_75.n1 a_2977_75.n0 25.576
R4026 a_2977_75.n3 a_2977_75.n2 9.111
R4027 a_2977_75.n7 a_2977_75.n6 2.455
R4028 a_2977_75.n5 a_2977_75.n3 1.964
R4029 a_2977_75.n5 a_2977_75.n4 1.964
R4030 a_2977_75.t0 a_2977_75.n1 1.871
R4031 a_2977_75.n7 a_2977_75.n5 0.636
R4032 a_2977_75.t0 a_2977_75.n7 0.246
R4033 a_1053_75.n1 a_1053_75.n0 25.576
R4034 a_1053_75.n3 a_1053_75.n2 9.111
R4035 a_1053_75.n7 a_1053_75.n6 2.455
R4036 a_1053_75.n5 a_1053_75.n3 1.964
R4037 a_1053_75.n5 a_1053_75.n4 1.964
R4038 a_1053_75.t0 a_1053_75.n1 1.871
R4039 a_1053_75.n7 a_1053_75.n5 0.636
R4040 a_1053_75.t0 a_1053_75.n7 0.246
R4041 a_3939_75.n5 a_3939_75.n4 19.724
R4042 a_3939_75.t0 a_3939_75.n3 11.595
R4043 a_3939_75.t0 a_3939_75.n5 9.207
R4044 a_3939_75.n2 a_3939_75.n1 2.455
R4045 a_3939_75.n2 a_3939_75.n0 1.32
R4046 a_3939_75.t0 a_3939_75.n2 0.246
R4047 a_9030_182.n10 a_9030_182.n8 82.852
R4048 a_9030_182.n7 a_9030_182.n6 32.833
R4049 a_9030_182.n8 a_9030_182.t1 32.416
R4050 a_9030_182.n10 a_9030_182.n9 27.2
R4051 a_9030_182.n11 a_9030_182.n0 23.498
R4052 a_9030_182.n3 a_9030_182.n2 23.284
R4053 a_9030_182.n11 a_9030_182.n10 22.4
R4054 a_9030_182.n7 a_9030_182.n4 19.017
R4055 a_9030_182.n6 a_9030_182.n5 13.494
R4056 a_9030_182.t1 a_9030_182.n1 7.04
R4057 a_9030_182.t1 a_9030_182.n3 5.727
R4058 a_9030_182.n8 a_9030_182.n7 1.435
R4059 a_4901_75.n5 a_4901_75.n4 19.724
R4060 a_4901_75.t0 a_4901_75.n3 11.595
R4061 a_4901_75.t0 a_4901_75.n5 9.207
R4062 a_4901_75.n2 a_4901_75.n1 2.455
R4063 a_4901_75.n2 a_4901_75.n0 1.32
R4064 a_4901_75.t0 a_4901_75.n2 0.246
R4065 a_6825_75.n1 a_6825_75.n0 25.576
R4066 a_6825_75.n3 a_6825_75.n2 9.111
R4067 a_6825_75.n7 a_6825_75.n6 2.455
R4068 a_6825_75.n5 a_6825_75.n3 1.964
R4069 a_6825_75.n5 a_6825_75.n4 1.964
R4070 a_6825_75.t0 a_6825_75.n1 1.871
R4071 a_6825_75.n7 a_6825_75.n5 0.636
R4072 a_6825_75.t0 a_6825_75.n7 0.246
R4073 a_18760_73.t0 a_18760_73.n1 34.62
R4074 a_18760_73.t0 a_18760_73.n0 8.137
R4075 a_18760_73.t0 a_18760_73.n2 4.69
R4076 a_11635_75.n1 a_11635_75.n0 25.576
R4077 a_11635_75.n3 a_11635_75.n2 9.111
R4078 a_11635_75.n7 a_11635_75.n6 2.455
R4079 a_11635_75.n5 a_11635_75.n3 1.964
R4080 a_11635_75.n5 a_11635_75.n4 1.964
R4081 a_11635_75.t0 a_11635_75.n1 1.871
R4082 a_11635_75.n7 a_11635_75.n5 0.636
R4083 a_11635_75.t0 a_11635_75.n7 0.246
R4084 a_5863_75.n1 a_5863_75.n0 25.576
R4085 a_5863_75.n3 a_5863_75.n2 9.111
R4086 a_5863_75.n7 a_5863_75.n6 2.455
R4087 a_5863_75.n5 a_5863_75.n3 1.964
R4088 a_5863_75.n5 a_5863_75.n4 1.964
R4089 a_5863_75.t0 a_5863_75.n1 1.871
R4090 a_5863_75.n7 a_5863_75.n5 0.636
R4091 a_5863_75.t0 a_5863_75.n7 0.246
R4092 a_7787_75.n1 a_7787_75.n0 25.576
R4093 a_7787_75.n3 a_7787_75.n2 9.111
R4094 a_7787_75.n7 a_7787_75.n6 2.455
R4095 a_7787_75.n5 a_7787_75.n3 1.964
R4096 a_7787_75.n5 a_7787_75.n4 1.964
R4097 a_7787_75.t0 a_7787_75.n1 1.871
R4098 a_7787_75.n7 a_7787_75.n5 0.636
R4099 a_7787_75.t0 a_7787_75.n7 0.246
R4100 a_9711_75.n5 a_9711_75.n4 19.724
R4101 a_9711_75.t0 a_9711_75.n3 11.595
R4102 a_9711_75.t0 a_9711_75.n5 9.207
R4103 a_9711_75.n2 a_9711_75.n1 2.455
R4104 a_9711_75.n2 a_9711_75.n0 1.32
R4105 a_9711_75.t0 a_9711_75.n2 0.246
R4106 a_8749_75.n1 a_8749_75.n0 25.576
R4107 a_8749_75.n3 a_8749_75.n2 9.111
R4108 a_8749_75.n7 a_8749_75.n6 2.455
R4109 a_8749_75.n5 a_8749_75.n3 1.964
R4110 a_8749_75.n5 a_8749_75.n4 1.964
R4111 a_8749_75.t0 a_8749_75.n1 1.871
R4112 a_8749_75.n7 a_8749_75.n5 0.636
R4113 a_8749_75.t0 a_8749_75.n7 0.246









































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































































.ends
