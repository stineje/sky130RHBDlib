** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/TMRDFFSNRNQNX1.sch
.subckt TMRDFFSNRNQNX1 QN D CLK SN RN VDD GND
*.PININFO QN:O D:I CLK:I SN:I RN:I
x4 QN net3 net2 net1 VDD VSS VOTERN3X1
x1 net3 D CLK SN RN VDD VSS DFFSNRNQX1
x2 net2 D CLK SN RN VDD VSS DFFSNRNQX1
x3 net1 D CLK SN RN VDD VSS DFFSNRNQX1
.ends

* expanding   symbol:  VOTERN3X1.sym # of pins=4
** sym_path: /home/rjridle/OpenRadHardSCL/lib/xschem/VOTERN3X1.sym
** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/VOTERN3X1.sch
.subckt VOTERN3X1  YN A B C  VDD  VSS VDD GND
*.PININFO YN:O A:I B:I C:I
XM2 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM3 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 YN A net2 VSS sky130_fd_pr__nfet_01v8 L=0.15u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM5 net3 B net1 VDD sky130_fd_pr__pfet_01v8 L=0.15u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM6 YN C net3 VDD sky130_fd_pr__pfet_01v8 L=0.15u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM7 net3 C net1 VDD sky130_fd_pr__pfet_01v8 L=0.15u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM10 YN A net3 VDD sky130_fd_pr__pfet_01v8 L=0.15u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM8 net4 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 YN C net4 VSS sky130_fd_pr__nfet_01v8 L=0.15u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 net5 C VSS VSS sky130_fd_pr__nfet_01v8 L=0.15u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 YN A net5 VSS sky130_fd_pr__nfet_01v8 L=0.15u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  DFFSNRNQX1.sym # of pins=5
** sym_path: /home/rjridle/OpenRadHardSCL/lib/xschem/DFFSNRNQX1.sym
** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/DFFSNRNQX1.sch
.subckt DFFSNRNQX1  Q D CLK SN RN  VDD  VSS VDD GND
*.PININFO Q:O D:I CLK:I SN:I RN:I
x1 net3 net1 SN net4 VDD VSS NAND3X1
x3 net2 net1 CLK net4 VDD VSS NAND3X1
x6 Q net5 SN net4 VDD VSS NAND3X1
x2 net1 D RN net2 VDD VSS NAND3X1
x4 net4 net3 CLK RN VDD VSS NAND3X1
x5 net5 net2 RN Q VDD VSS NAND3X1
.ends


* expanding   symbol:  NAND3X1.sym # of pins=4
** sym_path: /home/rjridle/OpenRadHardSCL/lib/xschem/NAND3X1.sym
** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/NAND3X1.sch
.subckt NAND3X1  Y A B C  VDD  VSS VDD GND
*.PININFO Y:O A:I B:I C:I
XM1 net2 A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM3 net1 B net2 VSS sky130_fd_pr__nfet_01v8 L=0.15u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 Y C net1 VSS sky130_fd_pr__nfet_01v8 L=0.15u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Y B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM6 Y C VDD VDD sky130_fd_pr__pfet_01v8 L=0.15u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends

.end
