* SPICE3 file created from DFFSNX1.ext - technology: sky130A

.subckt DFFSNX1 Q QN D CLK SN VDD GND
X0 a_1905_1004 a_217_1004 VDD VDD pshort w=2 l=0.15 M=2
X1 GND a_217_1004 a_757_75 GND nshort w=3 l=0.15
X2 VDD a_343_383 a_217_1004 VDD pshort w=2 l=0.15 M=2
X3 GND D a_112_73 GND nshort w=3 l=0.15
X4 GND a_343_383 a_3368_73 GND nshort w=3 l=0.15
X5 VDD a_217_1004 a_343_383 VDD pshort w=2 l=0.15 M=2
X6 QN Q VDD VDD pshort w=2 l=0.15 M=2
X7 VDD CLK a_343_383 VDD pshort w=2 l=0.15 M=2
X8 VDD a_1905_1004 a_1265_943 VDD pshort w=2 l=0.15 M=2
X9 QN a_343_383 VDD VDD pshort w=2 l=0.15 M=2
X10 GND a_217_1004 a_1719_75 GND nshort w=3 l=0.15
X11 VDD QN Q VDD pshort w=2 l=0.15 M=2
X12 VDD a_1265_943 Q VDD pshort w=2 l=0.15 M=2
X13 VDD a_1265_943 a_343_383 VDD pshort w=2 l=0.15 M=2
X14 a_1038_182 CLK a_757_75 GND nshort w=3 l=0.15
X15 a_217_1004 D VDD VDD pshort w=2 l=0.15 M=2
X16 a_1905_1004 a_1265_943 VDD VDD pshort w=2 l=0.15 M=2
X17 GND a_1905_1004 a_2702_73 GND nshort w=3 l=0.15
X18 a_217_1004 a_343_383 a_112_73 GND nshort w=3 l=0.15
X19 a_2000_182 SN a_1719_75 GND nshort w=3 l=0.15
X20 Q a_1265_943 a_4294_182 GND nshort w=3 l=0.15
X21 VDD SN Q VDD pshort w=2 l=0.15 M=2
X22 QN Q a_3368_73 GND nshort w=3 l=0.15
X23 a_1905_1004 SN VDD VDD pshort w=2 l=0.15 M=2
X24 GND QN a_4013_75 GND nshort w=3 l=0.15
X25 VDD CLK a_1265_943 VDD pshort w=2 l=0.15 M=2
X26 a_1265_943 CLK a_2702_73 GND nshort w=3 l=0.15
X27 a_4294_182 SN a_4013_75 GND nshort w=3 l=0.15
X28 a_1905_1004 a_1265_943 a_2000_182 GND nshort w=3 l=0.15
X29 a_343_383 a_1265_943 a_1038_182 GND nshort w=3 l=0.15
C0 a_343_383 CLK 2.36fF
C1 a_1905_1004 VDD 2.09fF
C2 a_343_383 VDD 3.07fF
C3 a_1265_943 VDD 2.14fF
C4 VDD Q 2.25fF
C5 a_1265_943 a_343_383 2.89fF
C6 VDD GND 11.88fF
.ends
