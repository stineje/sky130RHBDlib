* SPICE3 file created from TMRDFFRNQX1.ext - technology: sky130A

.subckt TMRDFFRNQX1 Q D CLK RN VDD GND
X0 GND m1_4419_797# dffrnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 dffrnx1_pcell_0/m1_867_723# dffrnx1_pcell_0/m1_689_649# dffrnx1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X2 dffrnx1_pcell_0/nand3x1_pcell_0/li_393_182# CLK dffrnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X3 VDD m1_4419_797# dffrnx1_pcell_0/m1_867_723# VDD pshort w=2 l=0.15
X4 VDD CLK dffrnx1_pcell_0/m1_867_723# VDD pshort w=2 l=0.15
X5 VDD dffrnx1_pcell_0/m1_689_649# dffrnx1_pcell_0/m1_867_723# VDD pshort w=2 l=0.15
X6 GND dffrnx1_pcell_0/m1_867_723# dffrnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X7 dffrnx1_pcell_0/m1_689_649# RN dffrnx1_pcell_0/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X8 dffrnx1_pcell_0/nand3x1_pcell_1/li_393_182# D dffrnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X9 VDD dffrnx1_pcell_0/m1_867_723# dffrnx1_pcell_0/m1_689_649# VDD pshort w=2 l=0.15
X10 VDD D dffrnx1_pcell_0/m1_689_649# VDD pshort w=2 l=0.15
X11 VDD RN dffrnx1_pcell_0/m1_689_649# VDD pshort w=2 l=0.15
X12 GND dffrnx1_pcell_0/m1_2461_649# dffrnx1_pcell_0/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X13 m1_4419_797# RN dffrnx1_pcell_0/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X14 dffrnx1_pcell_0/nand3x1_pcell_3/li_393_182# CLK dffrnx1_pcell_0/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X15 VDD dffrnx1_pcell_0/m1_2461_649# m1_4419_797# VDD pshort w=2 l=0.15
X16 VDD CLK m1_4419_797# VDD pshort w=2 l=0.15
X17 VDD RN m1_4419_797# VDD pshort w=2 l=0.15
X18 GND dffrnx1_pcell_0/m1_867_723# dffrnx1_pcell_0/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X19 m1_4419_797# m1_5061_575# dffrnx1_pcell_0/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X20 dffrnx1_pcell_0/nand3x1_pcell_4/li_393_182# RN dffrnx1_pcell_0/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X21 VDD dffrnx1_pcell_0/m1_867_723# m1_4419_797# VDD pshort w=2 l=0.15
X22 VDD m1_5061_575# m1_4419_797# VDD pshort w=2 l=0.15
X23 GND dffrnx1_pcell_0/m1_689_649# dffrnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X24 dffrnx1_pcell_0/m1_2461_649# m1_4419_797# dffrnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X25 VDD dffrnx1_pcell_0/m1_689_649# dffrnx1_pcell_0/m1_2461_649# VDD pshort w=2 l=0.15
X26 VDD m1_4419_797# dffrnx1_pcell_0/m1_2461_649# VDD pshort w=2 l=0.15
X27 GND m1_4419_797# dffrnx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X28 m1_5061_575# m1_4419_797# dffrnx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X29 VDD m1_4419_797# m1_5061_575# VDD pshort w=2 l=0.15
X30 GND dffrnx1_pcell_1/m1_241_797# dffrnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X31 dffrnx1_pcell_1/m1_867_723# dffrnx1_pcell_1/m1_689_649# dffrnx1_pcell_1/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X32 dffrnx1_pcell_1/nand3x1_pcell_0/li_393_182# CLK dffrnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X33 VDD dffrnx1_pcell_1/m1_241_797# dffrnx1_pcell_1/m1_867_723# VDD pshort w=2 l=0.15
X34 VDD CLK dffrnx1_pcell_1/m1_867_723# VDD pshort w=2 l=0.15
X35 VDD dffrnx1_pcell_1/m1_689_649# dffrnx1_pcell_1/m1_867_723# VDD pshort w=2 l=0.15
X36 GND dffrnx1_pcell_1/m1_867_723# dffrnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X37 dffrnx1_pcell_1/m1_689_649# RN dffrnx1_pcell_1/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X38 dffrnx1_pcell_1/nand3x1_pcell_1/li_393_182# D dffrnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X39 VDD dffrnx1_pcell_1/m1_867_723# dffrnx1_pcell_1/m1_689_649# VDD pshort w=2 l=0.15
X40 VDD D dffrnx1_pcell_1/m1_689_649# VDD pshort w=2 l=0.15
X41 VDD RN dffrnx1_pcell_1/m1_689_649# VDD pshort w=2 l=0.15
X42 GND dffrnx1_pcell_1/m1_2461_649# dffrnx1_pcell_1/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X43 dffrnx1_pcell_1/m1_241_797# RN dffrnx1_pcell_1/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X44 dffrnx1_pcell_1/nand3x1_pcell_3/li_393_182# CLK dffrnx1_pcell_1/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X45 VDD dffrnx1_pcell_1/m1_2461_649# dffrnx1_pcell_1/m1_241_797# VDD pshort w=2 l=0.15
X46 VDD CLK dffrnx1_pcell_1/m1_241_797# VDD pshort w=2 l=0.15
X47 VDD RN dffrnx1_pcell_1/m1_241_797# VDD pshort w=2 l=0.15
X48 GND dffrnx1_pcell_1/m1_867_723# dffrnx1_pcell_1/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X49 m1_9599_723# m1_9451_649# dffrnx1_pcell_1/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X50 dffrnx1_pcell_1/nand3x1_pcell_4/li_393_182# RN dffrnx1_pcell_1/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X51 VDD dffrnx1_pcell_1/m1_867_723# m1_9599_723# VDD pshort w=2 l=0.15
X52 VDD RN m1_9599_723# VDD pshort w=2 l=0.15
X53 VDD m1_9451_649# m1_9599_723# VDD pshort w=2 l=0.15
X54 GND dffrnx1_pcell_1/m1_689_649# dffrnx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X55 dffrnx1_pcell_1/m1_2461_649# dffrnx1_pcell_1/m1_241_797# dffrnx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X56 VDD dffrnx1_pcell_1/m1_689_649# dffrnx1_pcell_1/m1_2461_649# VDD pshort w=2 l=0.15
X57 VDD dffrnx1_pcell_1/m1_241_797# dffrnx1_pcell_1/m1_2461_649# VDD pshort w=2 l=0.15
X58 GND m1_9599_723# dffrnx1_pcell_1/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X59 m1_9451_649# dffrnx1_pcell_1/m1_241_797# dffrnx1_pcell_1/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X60 VDD m1_9599_723# m1_9451_649# VDD pshort w=2 l=0.15
X61 VDD dffrnx1_pcell_1/m1_241_797# m1_9451_649# VDD pshort w=2 l=0.15
X62 GND m1_14779_797# dffrnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X63 dffrnx1_pcell_2/m1_867_723# m1_9451_649# dffrnx1_pcell_2/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X64 dffrnx1_pcell_2/nand3x1_pcell_0/li_393_182# CLK dffrnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X65 VDD m1_14779_797# dffrnx1_pcell_2/m1_867_723# VDD pshort w=2 l=0.15
X66 VDD CLK dffrnx1_pcell_2/m1_867_723# VDD pshort w=2 l=0.15
X67 VDD m1_9451_649# dffrnx1_pcell_2/m1_867_723# VDD pshort w=2 l=0.15
X68 GND dffrnx1_pcell_2/m1_867_723# dffrnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X69 m1_9451_649# RN dffrnx1_pcell_2/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X70 dffrnx1_pcell_2/nand3x1_pcell_1/li_393_182# D dffrnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X71 VDD dffrnx1_pcell_2/m1_867_723# m1_9451_649# VDD pshort w=2 l=0.15
X72 VDD D m1_9451_649# VDD pshort w=2 l=0.15
X73 VDD RN m1_9451_649# VDD pshort w=2 l=0.15
X74 GND m1_9451_649# dffrnx1_pcell_2/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X75 m1_14779_797# RN dffrnx1_pcell_2/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X76 dffrnx1_pcell_2/nand3x1_pcell_3/li_393_182# CLK dffrnx1_pcell_2/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X77 VDD m1_9451_649# m1_14779_797# VDD pshort w=2 l=0.15
X78 VDD CLK m1_14779_797# VDD pshort w=2 l=0.15
X79 VDD RN m1_14779_797# VDD pshort w=2 l=0.15
X80 GND dffrnx1_pcell_2/m1_867_723# dffrnx1_pcell_2/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X81 m1_14779_797# m1_15421_723# dffrnx1_pcell_2/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X82 dffrnx1_pcell_2/nand3x1_pcell_4/li_393_182# RN dffrnx1_pcell_2/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X83 VDD dffrnx1_pcell_2/m1_867_723# m1_14779_797# VDD pshort w=2 l=0.15
X84 VDD m1_15421_723# m1_14779_797# VDD pshort w=2 l=0.15
X85 GND m1_9451_649# dffrnx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X86 m1_9451_649# m1_14779_797# dffrnx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X87 VDD m1_9451_649# m1_9451_649# VDD pshort w=2 l=0.15
X88 VDD m1_14779_797# m1_9451_649# VDD pshort w=2 l=0.15
X89 GND m1_14779_797# dffrnx1_pcell_2/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X90 m1_15421_723# m1_14779_797# dffrnx1_pcell_2/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X91 VDD m1_14779_797# m1_15421_723# VDD pshort w=2 l=0.15
X92 GND m1_9451_649# voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X93 GND m1_9451_649# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X94 GND m1_5061_575# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X95 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# m1_9451_649# VDD VDD pshort w=2 l=0.15
X96 voter3x1_pcell_0/m1_1867_797# m1_5061_575# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X97 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# m1_15421_723# VDD VDD pshort w=2 l=0.15
X98 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# m1_5061_575# voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X99 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# m1_9451_649# voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X100 voter3x1_pcell_0/m1_1867_797# m1_5061_575# voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X101 voter3x1_pcell_0/m1_1867_797# m1_15421_723# voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X102 voter3x1_pcell_0/m1_1867_797# m1_15421_723# voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X103 voter3x1_pcell_0/m1_1867_797# m1_15421_723# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X104 Q voter3x1_pcell_0/m1_1867_797# GND GND nshort w=3 l=0.15
X105 VDD voter3x1_pcell_0/m1_1867_797# Q VDD pshort w=2 l=0.15
C0 VDD RN 2.46fF
C1 dffrnx1_pcell_0/m1_867_723# dffrnx1_pcell_0/m1_689_649# 2.07fF
C2 dffrnx1_pcell_1/m1_241_797# dffrnx1_pcell_1/m1_867_723# 3.63fF
C3 m1_5061_575# m1_9451_649# 7.61fF
C4 m1_4419_797# dffrnx1_pcell_0/m1_867_723# 3.69fF
C5 VDD dffrnx1_pcell_1/m1_241_797# 2.85fF
C6 m1_9451_649# m1_14779_797# 2.98fF
C7 m1_4419_797# CLK 5.49fF
C8 m1_14779_797# dffrnx1_pcell_2/m1_867_723# 3.69fF
C9 CLK m1_14779_797# 3.54fF
C10 m1_9451_649# dffrnx1_pcell_2/m1_867_723# 4.14fF
C11 m1_9451_649# m1_15421_723# 2.50fF
C12 dffrnx1_pcell_1/m1_867_723# dffrnx1_pcell_1/m1_689_649# 2.07fF
C13 D RN 11.85fF
C14 VDD m1_4419_797# 4.08fF
C15 m1_5061_575# VDD 2.20fF
C16 m1_5061_575# RN 4.25fF
C17 VDD m1_14779_797# 4.24fF
C18 m1_9451_649# VDD 4.55fF
C19 VDD CLK 6.49fF
C20 CLK RN 2.13fF
C21 VDD m1_15421_723# 2.01fF
C22 VDD voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# 2.07fF
C23 dffrnx1_pcell_1/m1_241_797# CLK 5.65fF
C24 m1_5061_575# D 8.50fF
.ends
