* SPICE3 file created from TMRDFFRNQNX1.ext - technology: sky130A

.subckt TMRDFFRNQNX1 QN D CLK RN VPB VNB
M1000 a_14511_943.t3 a_10507_159.t14 VPB.t65 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_9331_943.t8 a_9331_943.t7 VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VNB a_9009_1004.t9 a_9806_73.t0 nshort w=-1.605u l=1.765u
+  ad=3.7611p pd=32.97u as=0p ps=0u
M1003 VPB.t44 RN a_9331_943.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VNB a_5779_943.t12 a_7216_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1005 VNB a_10507_159.t21 a_10451_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_5457_1004.t3 a_5779_943.t7 VPB.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_5327_159.t3 RN VPB.t41 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t8 a_147_159.t14 a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_15757_1005.t5 a_4151_943.t5 a_16421_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t67 a_10507_159.t15 a_10637_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPB.t4 a_9331_943.t19 a_10507_159.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t55 RN a_10507_159.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_10507_159.t3 a_10637_1004.t7 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_9331_943.t4 a_10637_1004.t8 VPB.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_599_943.t6 D VPB.t79 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_16421_1005.t6 a_14511_943.t6 a_15932_181.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_5327_159.t6 CLK VPB.t92 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPB.t15 a_599_943.t7 a_2141_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_9331_943.t13 a_9009_1004.t7 VPB.t60 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPB.t98 CLK a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPB.t17 a_5457_1004.t7 a_9009_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t85 a_277_1004.t8 a_147_159.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPB.t18 a_5457_1004.t8 a_5779_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPB.t50 RN a_5779_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPB.t69 a_9331_943.t21 a_9009_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPB.t95 CLK a_10507_159.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPB.t90 CLK a_10637_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_9331_943.t2 a_5327_159.t8 VPB.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VNB a_5457_1004.t11 a_8823_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_10507_159.t7 RN VPB.t54 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_9331_943.t18 D VPB.t82 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_599_943.t2 RN VPB.t58 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_147_159.t9 a_4151_943.t7 VPB.t76 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VNB a_5457_1004.t12 a_6233_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPB.t24 a_14511_943.t7 a_15757_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_10637_1004.t3 a_10507_159.t16 VPB.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_147_159.t13 CLK VPB.t87 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_4151_943.t3 a_147_159.t16 VPB.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_9009_1004.t5 a_5457_1004.t9 VPB.t59 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_15757_1005.t1 a_9331_943.t23 VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPB.t68 a_10507_159.t17 a_14511_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPB.t26 a_9331_943.t5 a_9331_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 VNB a_147_159.t15 a_4626_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPB.t0 a_147_159.t17 a_2141_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPB.t16 a_599_943.t9 a_277_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 VNB a_147_159.t24 a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPB.t83 D a_5779_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 VPB.t48 RN a_9009_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 VNB a_599_943.t8 a_2036_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1050 VNB a_7321_1004.t7 a_7861_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1051 VPB.t31 a_5327_159.t10 a_5457_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 VPB.t40 a_7321_1004.t5 a_5327_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 VPB.t36 a_2141_1004.t6 a_147_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_10507_159.t10 a_14511_943.t8 VPB.t72 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 VNB a_5327_159.t14 a_5271_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_9331_943.t10 RN VPB.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_147_159.t7 RN VPB.t57 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_4151_943.t2 a_147_159.t18 VPB.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 a_7321_1004.t1 a_5327_159.t11 VPB.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 a_15932_181.t2 a_4151_943.t8 a_16421_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 VPB.t1 a_9331_943.t26 a_10637_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 VNB a_9331_943.t24 a_15652_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1063 VNB a_10507_159.t18 a_14986_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_15757_1005.t6 a_14511_943.t9 VPB.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 VPB.t64 a_10507_159.t19 a_14511_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 VPB.t63 a_10507_159.t20 a_9331_943.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_277_1004.t3 a_147_159.t19 VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 VPB.t39 a_9009_1004.t8 a_9331_943.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_16421_1005.t5 a_4151_943.t10 a_15757_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 VNB a_9331_943.t20 a_13041_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_10507_159.t1 a_9331_943.t27 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_10507_159.t6 RN VPB.t53 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 a_10637_1004.t0 a_9331_943.t28 VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 VNB a_277_1004.t7 a_3643_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1075 a_7321_1004.t4 a_5779_943.t8 VPB.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 VPB.t86 a_277_1004.t10 a_599_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 a_15932_181.t4 a_14511_943.t10 a_16421_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 VPB.t56 RN a_599_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VPB.t32 a_4151_943.t11 a_147_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 VNB a_4151_943.t9 a_16984_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1081 VPB.t75 a_5779_943.t9 a_5457_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 VPB.t43 RN a_5327_159.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_16421_1005.t0 a_9331_943.t30 a_15757_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_2141_1004.t3 a_599_943.t10 VPB.t99 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_277_1004.t5 CLK VPB.t97 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_147_159.t2 a_277_1004.t11 VPB.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 a_5779_943.t1 a_5457_1004.t10 VPB.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_10507_159.t12 CLK VPB.t94 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_10637_1004.t5 CLK VPB.t96 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 VNB a_10637_1004.t9 a_14003_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1091 VNB a_2141_1004.t5 a_2681_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1092 VPB.t38 a_10637_1004.t11 a_10507_159.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 VPB.t25 a_10637_1004.t12 a_9331_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 VPB.t81 D a_599_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 VPB.t47 RN a_147_159.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 VNB a_9331_943.t29 a_12396_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_599_943.t3 a_277_1004.t12 VPB.t33 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 VPB.t89 CLK a_5457_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 VPB.t91 CLK a_5327_159.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_2141_1004.t0 a_147_159.t22 VPB.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 a_277_1004.t0 a_599_943.t11 VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_147_159.t5 RN VPB.t42 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_5779_943.t5 D VPB.t78 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_9009_1004.t3 RN VPB.t51 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 a_5327_159.t0 a_7321_1004.t6 VPB.t37 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VPB.t29 a_5327_159.t12 a_9331_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 a_147_159.t10 a_2141_1004.t7 VPB.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 a_5457_1004.t0 a_5327_159.t13 VPB.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 VPB.t52 RN a_10507_159.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 VPB.t80 D a_9331_943.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 VNB a_277_1004.t9 a_1053_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1112 VPB.t88 CLK a_147_159.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 VPB.t70 a_5779_943.t10 a_7321_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1114 VPB.t7 a_147_159.t23 a_4151_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 VPB.t20 a_9331_943.t32 a_15757_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 a_14511_943.t0 a_10507_159.t23 VPB.t61 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_9331_943.t14 a_10507_159.t24 VPB.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 VNB a_9331_943.t31 a_16318_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_9009_1004.t0 a_9331_943.t33 VPB.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 a_5779_943.t2 RN VPB.t49 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 VNB a_10637_1004.t10 a_11413_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1122 a_5457_1004.t5 CLK VPB.t93 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 a_15757_1005.t2 a_9331_943.t34 a_16421_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1124 VPB.t11 a_14511_943.t13 a_10507_159.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1125 VPB.t46 RN a_147_159.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1126 VPB.t74 a_147_159.t25 a_4151_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1127 VPB.t77 a_5327_159.t15 a_7321_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1128 a_16421_1005.t4 a_4151_943.t13 a_15932_181.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB D 0.15fF
C1 VPB CLK 3.49fF
C2 VPB RN 0.50fF
C3 D CLK 1.65fF
C4 D RN 12.41fF
C5 CLK RN 1.02fF
R0 a_10507_159.n21 a_10507_159.t15 512.525
R1 a_10507_159.n8 a_10507_159.t17 480.392
R2 a_10507_159.n19 a_10507_159.t20 472.359
R3 a_10507_159.n6 a_10507_159.t19 472.359
R4 a_10507_159.n8 a_10507_159.t14 403.272
R5 a_10507_159.n19 a_10507_159.t24 384.527
R6 a_10507_159.n6 a_10507_159.t23 384.527
R7 a_10507_159.n21 a_10507_159.t16 371.139
R8 a_10507_159.n22 a_10507_159.t21 324.268
R9 a_10507_159.n9 a_10507_159.t18 320.08
R10 a_10507_159.n20 a_10507_159.t25 277.772
R11 a_10507_159.n7 a_10507_159.t22 277.772
R12 a_10507_159.n17 a_10507_159.n16 271.443
R13 a_10507_159.n27 a_10507_159.n25 249.704
R14 a_10507_159.n17 a_10507_159.n15 127.74
R15 a_10507_159.n25 a_10507_159.n5 127.74
R16 a_10507_159.n22 a_10507_159.n21 119.654
R17 a_10507_159.n23 a_10507_159.n22 83.572
R18 a_10507_159.n14 a_10507_159.n13 79.232
R19 a_10507_159.n4 a_10507_159.n3 79.232
R20 a_10507_159.n10 a_10507_159.n7 76.499
R21 a_10507_159.n23 a_10507_159.n20 76
R22 a_10507_159.n10 a_10507_159.n9 76
R23 a_10507_159.n18 a_10507_159.n17 76
R24 a_10507_159.n25 a_10507_159.n24 76
R25 a_10507_159.n20 a_10507_159.n19 67.001
R26 a_10507_159.n7 a_10507_159.n6 67.001
R27 a_10507_159.n15 a_10507_159.n14 63.152
R28 a_10507_159.n5 a_10507_159.n4 63.152
R29 a_10507_159.n9 a_10507_159.n8 55.388
R30 a_10507_159.n27 a_10507_159.n26 30
R31 a_10507_159.n28 a_10507_159.n0 24.383
R32 a_10507_159.n28 a_10507_159.n27 23.684
R33 a_10507_159.n15 a_10507_159.n11 16.08
R34 a_10507_159.n14 a_10507_159.n12 16.08
R35 a_10507_159.n5 a_10507_159.n1 16.08
R36 a_10507_159.n4 a_10507_159.n2 16.08
R37 a_10507_159.n11 a_10507_159.t2 14.282
R38 a_10507_159.n11 a_10507_159.t10 14.282
R39 a_10507_159.n12 a_10507_159.t5 14.282
R40 a_10507_159.n12 a_10507_159.t7 14.282
R41 a_10507_159.n13 a_10507_159.t4 14.282
R42 a_10507_159.n13 a_10507_159.t3 14.282
R43 a_10507_159.n1 a_10507_159.t8 14.282
R44 a_10507_159.n1 a_10507_159.t6 14.282
R45 a_10507_159.n2 a_10507_159.t13 14.282
R46 a_10507_159.n2 a_10507_159.t12 14.282
R47 a_10507_159.n3 a_10507_159.t0 14.282
R48 a_10507_159.n3 a_10507_159.t1 14.282
R49 a_10507_159.n24 a_10507_159.n23 4.035
R50 a_10507_159.n24 a_10507_159.n18 3.491
R51 a_10507_159.n18 a_10507_159.n10 1.315
R52 VPB VPB.n1562 126.832
R53 VPB.n40 VPB.n38 94.117
R54 VPB.n1484 VPB.n1482 94.117
R55 VPB.n1421 VPB.n1419 94.117
R56 VPB.n1338 VPB.n1336 94.117
R57 VPB.n1255 VPB.n1253 94.117
R58 VPB.n1192 VPB.n1190 94.117
R59 VPB.n1109 VPB.n1107 94.117
R60 VPB.n1026 VPB.n1024 94.117
R61 VPB.n963 VPB.n961 94.117
R62 VPB.n880 VPB.n878 94.117
R63 VPB.n129 VPB.n127 94.117
R64 VPB.n823 VPB.n821 94.117
R65 VPB.n740 VPB.n738 94.117
R66 VPB.n657 VPB.n655 94.117
R67 VPB.n594 VPB.n592 94.117
R68 VPB.n511 VPB.n509 94.117
R69 VPB.n428 VPB.n426 94.117
R70 VPB.n365 VPB.n363 94.117
R71 VPB.n302 VPB.n300 94.117
R72 VPB.n247 VPB.n245 94.117
R73 VPB.n441 VPB.n440 80.104
R74 VPB.n524 VPB.n523 80.104
R75 VPB.n670 VPB.n669 80.104
R76 VPB.n753 VPB.n752 80.104
R77 VPB.n139 VPB.n138 80.104
R78 VPB.n893 VPB.n892 80.104
R79 VPB.n1039 VPB.n1038 80.104
R80 VPB.n1122 VPB.n1121 80.104
R81 VPB.n1268 VPB.n1267 80.104
R82 VPB.n1351 VPB.n1350 80.104
R83 VPB.n1497 VPB.n1496 80.104
R84 VPB.n50 VPB.n49 80.104
R85 VPB.n210 VPB.n209 76
R86 VPB.n214 VPB.n213 76
R87 VPB.n218 VPB.n217 76
R88 VPB.n222 VPB.n221 76
R89 VPB.n249 VPB.n248 76
R90 VPB.n253 VPB.n252 76
R91 VPB.n257 VPB.n256 76
R92 VPB.n261 VPB.n260 76
R93 VPB.n265 VPB.n264 76
R94 VPB.n269 VPB.n268 76
R95 VPB.n273 VPB.n272 76
R96 VPB.n277 VPB.n276 76
R97 VPB.n304 VPB.n303 76
R98 VPB.n309 VPB.n308 76
R99 VPB.n314 VPB.n313 76
R100 VPB.n321 VPB.n320 76
R101 VPB.n326 VPB.n325 76
R102 VPB.n331 VPB.n330 76
R103 VPB.n336 VPB.n335 76
R104 VPB.n340 VPB.n339 76
R105 VPB.n367 VPB.n366 76
R106 VPB.n372 VPB.n371 76
R107 VPB.n377 VPB.n376 76
R108 VPB.n384 VPB.n383 76
R109 VPB.n389 VPB.n388 76
R110 VPB.n394 VPB.n393 76
R111 VPB.n399 VPB.n398 76
R112 VPB.n403 VPB.n402 76
R113 VPB.n430 VPB.n429 76
R114 VPB.n434 VPB.n433 76
R115 VPB.n439 VPB.n438 76
R116 VPB.n444 VPB.n443 76
R117 VPB.n451 VPB.n450 76
R118 VPB.n456 VPB.n455 76
R119 VPB.n461 VPB.n460 76
R120 VPB.n468 VPB.n467 76
R121 VPB.n473 VPB.n472 76
R122 VPB.n478 VPB.n477 76
R123 VPB.n482 VPB.n481 76
R124 VPB.n486 VPB.n485 76
R125 VPB.n513 VPB.n512 76
R126 VPB.n517 VPB.n516 76
R127 VPB.n522 VPB.n521 76
R128 VPB.n527 VPB.n526 76
R129 VPB.n534 VPB.n533 76
R130 VPB.n539 VPB.n538 76
R131 VPB.n544 VPB.n543 76
R132 VPB.n551 VPB.n550 76
R133 VPB.n556 VPB.n555 76
R134 VPB.n561 VPB.n560 76
R135 VPB.n565 VPB.n564 76
R136 VPB.n569 VPB.n568 76
R137 VPB.n596 VPB.n595 76
R138 VPB.n601 VPB.n600 76
R139 VPB.n606 VPB.n605 76
R140 VPB.n613 VPB.n612 76
R141 VPB.n618 VPB.n617 76
R142 VPB.n623 VPB.n622 76
R143 VPB.n628 VPB.n627 76
R144 VPB.n632 VPB.n631 76
R145 VPB.n659 VPB.n658 76
R146 VPB.n663 VPB.n662 76
R147 VPB.n668 VPB.n667 76
R148 VPB.n673 VPB.n672 76
R149 VPB.n680 VPB.n679 76
R150 VPB.n685 VPB.n684 76
R151 VPB.n690 VPB.n689 76
R152 VPB.n697 VPB.n696 76
R153 VPB.n702 VPB.n701 76
R154 VPB.n707 VPB.n706 76
R155 VPB.n711 VPB.n710 76
R156 VPB.n715 VPB.n714 76
R157 VPB.n742 VPB.n741 76
R158 VPB.n746 VPB.n745 76
R159 VPB.n751 VPB.n750 76
R160 VPB.n756 VPB.n755 76
R161 VPB.n763 VPB.n762 76
R162 VPB.n768 VPB.n767 76
R163 VPB.n773 VPB.n772 76
R164 VPB.n780 VPB.n779 76
R165 VPB.n785 VPB.n784 76
R166 VPB.n790 VPB.n789 76
R167 VPB.n794 VPB.n793 76
R168 VPB.n798 VPB.n797 76
R169 VPB.n825 VPB.n824 76
R170 VPB.n830 VPB.n829 76
R171 VPB.n835 VPB.n834 76
R172 VPB.n842 VPB.n841 76
R173 VPB.n847 VPB.n846 76
R174 VPB.n852 VPB.n851 76
R175 VPB.n857 VPB.n856 76
R176 VPB.n861 VPB.n860 76
R177 VPB.n876 VPB.n873 76
R178 VPB.n882 VPB.n881 76
R179 VPB.n886 VPB.n885 76
R180 VPB.n891 VPB.n890 76
R181 VPB.n896 VPB.n895 76
R182 VPB.n903 VPB.n902 76
R183 VPB.n908 VPB.n907 76
R184 VPB.n913 VPB.n912 76
R185 VPB.n920 VPB.n919 76
R186 VPB.n925 VPB.n924 76
R187 VPB.n930 VPB.n929 76
R188 VPB.n934 VPB.n933 76
R189 VPB.n938 VPB.n937 76
R190 VPB.n965 VPB.n964 76
R191 VPB.n970 VPB.n969 76
R192 VPB.n975 VPB.n974 76
R193 VPB.n982 VPB.n981 76
R194 VPB.n987 VPB.n986 76
R195 VPB.n992 VPB.n991 76
R196 VPB.n997 VPB.n996 76
R197 VPB.n1001 VPB.n1000 76
R198 VPB.n1028 VPB.n1027 76
R199 VPB.n1032 VPB.n1031 76
R200 VPB.n1037 VPB.n1036 76
R201 VPB.n1042 VPB.n1041 76
R202 VPB.n1049 VPB.n1048 76
R203 VPB.n1054 VPB.n1053 76
R204 VPB.n1059 VPB.n1058 76
R205 VPB.n1066 VPB.n1065 76
R206 VPB.n1071 VPB.n1070 76
R207 VPB.n1076 VPB.n1075 76
R208 VPB.n1080 VPB.n1079 76
R209 VPB.n1084 VPB.n1083 76
R210 VPB.n1111 VPB.n1110 76
R211 VPB.n1115 VPB.n1114 76
R212 VPB.n1120 VPB.n1119 76
R213 VPB.n1125 VPB.n1124 76
R214 VPB.n1132 VPB.n1131 76
R215 VPB.n1137 VPB.n1136 76
R216 VPB.n1142 VPB.n1141 76
R217 VPB.n1149 VPB.n1148 76
R218 VPB.n1154 VPB.n1153 76
R219 VPB.n1159 VPB.n1158 76
R220 VPB.n1163 VPB.n1162 76
R221 VPB.n1167 VPB.n1166 76
R222 VPB.n1194 VPB.n1193 76
R223 VPB.n1199 VPB.n1198 76
R224 VPB.n1204 VPB.n1203 76
R225 VPB.n1211 VPB.n1210 76
R226 VPB.n1216 VPB.n1215 76
R227 VPB.n1221 VPB.n1220 76
R228 VPB.n1226 VPB.n1225 76
R229 VPB.n1230 VPB.n1229 76
R230 VPB.n1257 VPB.n1256 76
R231 VPB.n1261 VPB.n1260 76
R232 VPB.n1266 VPB.n1265 76
R233 VPB.n1271 VPB.n1270 76
R234 VPB.n1278 VPB.n1277 76
R235 VPB.n1283 VPB.n1282 76
R236 VPB.n1288 VPB.n1287 76
R237 VPB.n1295 VPB.n1294 76
R238 VPB.n1300 VPB.n1299 76
R239 VPB.n1305 VPB.n1304 76
R240 VPB.n1309 VPB.n1308 76
R241 VPB.n1313 VPB.n1312 76
R242 VPB.n1340 VPB.n1339 76
R243 VPB.n1344 VPB.n1343 76
R244 VPB.n1349 VPB.n1348 76
R245 VPB.n1354 VPB.n1353 76
R246 VPB.n1361 VPB.n1360 76
R247 VPB.n1366 VPB.n1365 76
R248 VPB.n1371 VPB.n1370 76
R249 VPB.n1378 VPB.n1377 76
R250 VPB.n1383 VPB.n1382 76
R251 VPB.n1388 VPB.n1387 76
R252 VPB.n1392 VPB.n1391 76
R253 VPB.n1396 VPB.n1395 76
R254 VPB.n1423 VPB.n1422 76
R255 VPB.n1428 VPB.n1427 76
R256 VPB.n1433 VPB.n1432 76
R257 VPB.n1440 VPB.n1439 76
R258 VPB.n1445 VPB.n1444 76
R259 VPB.n1450 VPB.n1449 76
R260 VPB.n1455 VPB.n1454 76
R261 VPB.n1459 VPB.n1458 76
R262 VPB.n1486 VPB.n1485 76
R263 VPB.n1490 VPB.n1489 76
R264 VPB.n1495 VPB.n1494 76
R265 VPB.n1500 VPB.n1499 76
R266 VPB.n1507 VPB.n1506 76
R267 VPB.n1512 VPB.n1511 76
R268 VPB.n1517 VPB.n1516 76
R269 VPB.n1524 VPB.n1523 76
R270 VPB.n1529 VPB.n1528 76
R271 VPB.n1534 VPB.n1533 76
R272 VPB.n1538 VPB.n1537 76
R273 VPB.n1542 VPB.n1541 76
R274 VPB.n1555 VPB.n1554 76
R275 VPB.n470 VPB.n469 75.654
R276 VPB.n553 VPB.n552 75.654
R277 VPB.n699 VPB.n698 75.654
R278 VPB.n782 VPB.n781 75.654
R279 VPB.n161 VPB.n160 75.654
R280 VPB.n922 VPB.n921 75.654
R281 VPB.n1068 VPB.n1067 75.654
R282 VPB.n1151 VPB.n1150 75.654
R283 VPB.n1297 VPB.n1296 75.654
R284 VPB.n1380 VPB.n1379 75.654
R285 VPB.n1526 VPB.n1525 75.654
R286 VPB.n72 VPB.n71 75.654
R287 VPB.n22 VPB.n21 61.764
R288 VPB.n1466 VPB.n1465 61.764
R289 VPB.n1403 VPB.n1402 61.764
R290 VPB.n1320 VPB.n1319 61.764
R291 VPB.n1237 VPB.n1236 61.764
R292 VPB.n1174 VPB.n1173 61.764
R293 VPB.n1091 VPB.n1090 61.764
R294 VPB.n1008 VPB.n1007 61.764
R295 VPB.n945 VPB.n944 61.764
R296 VPB.n88 VPB.n87 61.764
R297 VPB.n111 VPB.n110 61.764
R298 VPB.n805 VPB.n804 61.764
R299 VPB.n722 VPB.n721 61.764
R300 VPB.n639 VPB.n638 61.764
R301 VPB.n576 VPB.n575 61.764
R302 VPB.n493 VPB.n492 61.764
R303 VPB.n410 VPB.n409 61.764
R304 VPB.n347 VPB.n346 61.764
R305 VPB.n284 VPB.n283 61.764
R306 VPB.n229 VPB.n228 61.764
R307 VPB.n332 VPB.t9 55.465
R308 VPB.n305 VPB.t24 55.465
R309 VPB.n78 VPB.t5 55.106
R310 VPB.n1530 VPB.t33 55.106
R311 VPB.n1451 VPB.t99 55.106
R312 VPB.n1384 VPB.t84 55.106
R313 VPB.n1301 VPB.t35 55.106
R314 VPB.n1222 VPB.t13 55.106
R315 VPB.n1155 VPB.t27 55.106
R316 VPB.n1072 VPB.t21 55.106
R317 VPB.n993 VPB.t71 55.106
R318 VPB.n926 VPB.t37 55.106
R319 VPB.n167 VPB.t59 55.106
R320 VPB.n853 VPB.t60 55.106
R321 VPB.n786 VPB.t66 55.106
R322 VPB.n703 VPB.t34 55.106
R323 VPB.n624 VPB.t2 55.106
R324 VPB.n557 VPB.t6 55.106
R325 VPB.n474 VPB.t12 55.106
R326 VPB.n395 VPB.t65 55.106
R327 VPB.n45 VPB.t16 55.106
R328 VPB.n1491 VPB.t56 55.106
R329 VPB.n1424 VPB.t0 55.106
R330 VPB.n1345 VPB.t46 55.106
R331 VPB.n1262 VPB.t32 55.106
R332 VPB.n1195 VPB.t74 55.106
R333 VPB.n1116 VPB.t75 55.106
R334 VPB.n1033 VPB.t50 55.106
R335 VPB.n966 VPB.t77 55.106
R336 VPB.n887 VPB.t43 55.106
R337 VPB.n134 VPB.t69 55.106
R338 VPB.n826 VPB.t29 55.106
R339 VPB.n747 VPB.t1 55.106
R340 VPB.n664 VPB.t44 55.106
R341 VPB.n597 VPB.t63 55.106
R342 VPB.n518 VPB.t55 55.106
R343 VPB.n435 VPB.t11 55.106
R344 VPB.n368 VPB.t64 55.106
R345 VPB.n311 VPB.n310 48.952
R346 VPB.n374 VPB.n373 48.952
R347 VPB.n448 VPB.n447 48.952
R348 VPB.n531 VPB.n530 48.952
R349 VPB.n603 VPB.n602 48.952
R350 VPB.n677 VPB.n676 48.952
R351 VPB.n760 VPB.n759 48.952
R352 VPB.n832 VPB.n831 48.952
R353 VPB.n143 VPB.n142 48.952
R354 VPB.n900 VPB.n899 48.952
R355 VPB.n972 VPB.n971 48.952
R356 VPB.n1046 VPB.n1045 48.952
R357 VPB.n1129 VPB.n1128 48.952
R358 VPB.n1201 VPB.n1200 48.952
R359 VPB.n1275 VPB.n1274 48.952
R360 VPB.n1358 VPB.n1357 48.952
R361 VPB.n1430 VPB.n1429 48.952
R362 VPB.n1504 VPB.n1503 48.952
R363 VPB.n54 VPB.n53 48.952
R364 VPB.n328 VPB.n327 44.502
R365 VPB.n391 VPB.n390 44.502
R366 VPB.n465 VPB.n464 44.502
R367 VPB.n548 VPB.n547 44.502
R368 VPB.n620 VPB.n619 44.502
R369 VPB.n694 VPB.n693 44.502
R370 VPB.n777 VPB.n776 44.502
R371 VPB.n849 VPB.n848 44.502
R372 VPB.n157 VPB.n156 44.502
R373 VPB.n917 VPB.n916 44.502
R374 VPB.n989 VPB.n988 44.502
R375 VPB.n1063 VPB.n1062 44.502
R376 VPB.n1146 VPB.n1145 44.502
R377 VPB.n1218 VPB.n1217 44.502
R378 VPB.n1292 VPB.n1291 44.502
R379 VPB.n1375 VPB.n1374 44.502
R380 VPB.n1447 VPB.n1446 44.502
R381 VPB.n1521 VPB.n1520 44.502
R382 VPB.n68 VPB.n67 44.502
R383 VPB.n316 VPB.n315 41.183
R384 VPB.n66 VPB.n14 40.824
R385 VPB.n57 VPB.n15 40.824
R386 VPB.n1519 VPB.n1518 40.824
R387 VPB.n1502 VPB.n1501 40.824
R388 VPB.n1435 VPB.n1434 40.824
R389 VPB.n1373 VPB.n1372 40.824
R390 VPB.n1356 VPB.n1355 40.824
R391 VPB.n1290 VPB.n1289 40.824
R392 VPB.n1273 VPB.n1272 40.824
R393 VPB.n1206 VPB.n1205 40.824
R394 VPB.n1144 VPB.n1143 40.824
R395 VPB.n1127 VPB.n1126 40.824
R396 VPB.n1061 VPB.n1060 40.824
R397 VPB.n1044 VPB.n1043 40.824
R398 VPB.n977 VPB.n976 40.824
R399 VPB.n915 VPB.n914 40.824
R400 VPB.n898 VPB.n897 40.824
R401 VPB.n155 VPB.n103 40.824
R402 VPB.n146 VPB.n104 40.824
R403 VPB.n837 VPB.n836 40.824
R404 VPB.n775 VPB.n774 40.824
R405 VPB.n758 VPB.n757 40.824
R406 VPB.n692 VPB.n691 40.824
R407 VPB.n675 VPB.n674 40.824
R408 VPB.n608 VPB.n607 40.824
R409 VPB.n546 VPB.n545 40.824
R410 VPB.n529 VPB.n528 40.824
R411 VPB.n463 VPB.n462 40.824
R412 VPB.n446 VPB.n445 40.824
R413 VPB.n379 VPB.n378 40.824
R414 VPB.n205 VPB.n204 35.118
R415 VPB.n1559 VPB.n1555 20.452
R416 VPB.n194 VPB.n191 20.452
R417 VPB.n318 VPB.n317 17.801
R418 VPB.n381 VPB.n380 17.801
R419 VPB.n453 VPB.n452 17.801
R420 VPB.n536 VPB.n535 17.801
R421 VPB.n610 VPB.n609 17.801
R422 VPB.n682 VPB.n681 17.801
R423 VPB.n765 VPB.n764 17.801
R424 VPB.n839 VPB.n838 17.801
R425 VPB.n148 VPB.n147 17.801
R426 VPB.n905 VPB.n904 17.801
R427 VPB.n979 VPB.n978 17.801
R428 VPB.n1051 VPB.n1050 17.801
R429 VPB.n1134 VPB.n1133 17.801
R430 VPB.n1208 VPB.n1207 17.801
R431 VPB.n1280 VPB.n1279 17.801
R432 VPB.n1363 VPB.n1362 17.801
R433 VPB.n1437 VPB.n1436 17.801
R434 VPB.n1509 VPB.n1508 17.801
R435 VPB.n59 VPB.n58 17.801
R436 VPB.n14 VPB.t97 14.282
R437 VPB.n14 VPB.t8 14.282
R438 VPB.n15 VPB.t14 14.282
R439 VPB.n15 VPB.t98 14.282
R440 VPB.n1518 VPB.t79 14.282
R441 VPB.n1518 VPB.t86 14.282
R442 VPB.n1501 VPB.t58 14.282
R443 VPB.n1501 VPB.t81 14.282
R444 VPB.n1434 VPB.t73 14.282
R445 VPB.n1434 VPB.t15 14.282
R446 VPB.n1372 VPB.t87 14.282
R447 VPB.n1372 VPB.t36 14.282
R448 VPB.n1355 VPB.t57 14.282
R449 VPB.n1355 VPB.t88 14.282
R450 VPB.n1289 VPB.t42 14.282
R451 VPB.n1289 VPB.t85 14.282
R452 VPB.n1272 VPB.t76 14.282
R453 VPB.n1272 VPB.t47 14.282
R454 VPB.n1205 VPB.t22 14.282
R455 VPB.n1205 VPB.t7 14.282
R456 VPB.n1143 VPB.t93 14.282
R457 VPB.n1143 VPB.t31 14.282
R458 VPB.n1126 VPB.t10 14.282
R459 VPB.n1126 VPB.t89 14.282
R460 VPB.n1060 VPB.t78 14.282
R461 VPB.n1060 VPB.t18 14.282
R462 VPB.n1043 VPB.t49 14.282
R463 VPB.n1043 VPB.t83 14.282
R464 VPB.n976 VPB.t30 14.282
R465 VPB.n976 VPB.t70 14.282
R466 VPB.n914 VPB.t92 14.282
R467 VPB.n914 VPB.t40 14.282
R468 VPB.n897 VPB.t41 14.282
R469 VPB.n897 VPB.t91 14.282
R470 VPB.n103 VPB.t51 14.282
R471 VPB.n103 VPB.t17 14.282
R472 VPB.n104 VPB.t23 14.282
R473 VPB.n104 VPB.t48 14.282
R474 VPB.n836 VPB.t28 14.282
R475 VPB.n836 VPB.t39 14.282
R476 VPB.n774 VPB.t96 14.282
R477 VPB.n774 VPB.t67 14.282
R478 VPB.n757 VPB.t3 14.282
R479 VPB.n757 VPB.t90 14.282
R480 VPB.n691 VPB.t82 14.282
R481 VPB.n691 VPB.t25 14.282
R482 VPB.n674 VPB.t45 14.282
R483 VPB.n674 VPB.t80 14.282
R484 VPB.n607 VPB.t62 14.282
R485 VPB.n607 VPB.t26 14.282
R486 VPB.n545 VPB.t94 14.282
R487 VPB.n545 VPB.t4 14.282
R488 VPB.n528 VPB.t53 14.282
R489 VPB.n528 VPB.t95 14.282
R490 VPB.n462 VPB.t54 14.282
R491 VPB.n462 VPB.t38 14.282
R492 VPB.n445 VPB.t72 14.282
R493 VPB.n445 VPB.t52 14.282
R494 VPB.n378 VPB.t61 14.282
R495 VPB.n378 VPB.t68 14.282
R496 VPB.n315 VPB.t19 14.282
R497 VPB.n315 VPB.t20 14.282
R498 VPB.n194 VPB.n193 13.653
R499 VPB.n193 VPB.n192 13.653
R500 VPB.n203 VPB.n202 13.653
R501 VPB.n202 VPB.n201 13.653
R502 VPB.n200 VPB.n199 13.653
R503 VPB.n199 VPB.n198 13.653
R504 VPB.n197 VPB.n196 13.653
R505 VPB.n196 VPB.n195 13.653
R506 VPB.n209 VPB.n208 13.653
R507 VPB.n208 VPB.n207 13.653
R508 VPB.n213 VPB.n212 13.653
R509 VPB.n212 VPB.n211 13.653
R510 VPB.n217 VPB.n216 13.653
R511 VPB.n216 VPB.n215 13.653
R512 VPB.n221 VPB.n220 13.653
R513 VPB.n220 VPB.n219 13.653
R514 VPB.n248 VPB.n247 13.653
R515 VPB.n247 VPB.n246 13.653
R516 VPB.n252 VPB.n251 13.653
R517 VPB.n251 VPB.n250 13.653
R518 VPB.n256 VPB.n255 13.653
R519 VPB.n255 VPB.n254 13.653
R520 VPB.n260 VPB.n259 13.653
R521 VPB.n259 VPB.n258 13.653
R522 VPB.n264 VPB.n263 13.653
R523 VPB.n263 VPB.n262 13.653
R524 VPB.n268 VPB.n267 13.653
R525 VPB.n267 VPB.n266 13.653
R526 VPB.n272 VPB.n271 13.653
R527 VPB.n271 VPB.n270 13.653
R528 VPB.n276 VPB.n275 13.653
R529 VPB.n275 VPB.n274 13.653
R530 VPB.n303 VPB.n302 13.653
R531 VPB.n302 VPB.n301 13.653
R532 VPB.n308 VPB.n307 13.653
R533 VPB.n307 VPB.n306 13.653
R534 VPB.n313 VPB.n312 13.653
R535 VPB.n312 VPB.n311 13.653
R536 VPB.n320 VPB.n319 13.653
R537 VPB.n319 VPB.n318 13.653
R538 VPB.n325 VPB.n324 13.653
R539 VPB.n324 VPB.n323 13.653
R540 VPB.n330 VPB.n329 13.653
R541 VPB.n329 VPB.n328 13.653
R542 VPB.n335 VPB.n334 13.653
R543 VPB.n334 VPB.n333 13.653
R544 VPB.n339 VPB.n338 13.653
R545 VPB.n338 VPB.n337 13.653
R546 VPB.n366 VPB.n365 13.653
R547 VPB.n365 VPB.n364 13.653
R548 VPB.n371 VPB.n370 13.653
R549 VPB.n370 VPB.n369 13.653
R550 VPB.n376 VPB.n375 13.653
R551 VPB.n375 VPB.n374 13.653
R552 VPB.n383 VPB.n382 13.653
R553 VPB.n382 VPB.n381 13.653
R554 VPB.n388 VPB.n387 13.653
R555 VPB.n387 VPB.n386 13.653
R556 VPB.n393 VPB.n392 13.653
R557 VPB.n392 VPB.n391 13.653
R558 VPB.n398 VPB.n397 13.653
R559 VPB.n397 VPB.n396 13.653
R560 VPB.n402 VPB.n401 13.653
R561 VPB.n401 VPB.n400 13.653
R562 VPB.n429 VPB.n428 13.653
R563 VPB.n428 VPB.n427 13.653
R564 VPB.n433 VPB.n432 13.653
R565 VPB.n432 VPB.n431 13.653
R566 VPB.n438 VPB.n437 13.653
R567 VPB.n437 VPB.n436 13.653
R568 VPB.n443 VPB.n442 13.653
R569 VPB.n442 VPB.n441 13.653
R570 VPB.n450 VPB.n449 13.653
R571 VPB.n449 VPB.n448 13.653
R572 VPB.n455 VPB.n454 13.653
R573 VPB.n454 VPB.n453 13.653
R574 VPB.n460 VPB.n459 13.653
R575 VPB.n459 VPB.n458 13.653
R576 VPB.n467 VPB.n466 13.653
R577 VPB.n466 VPB.n465 13.653
R578 VPB.n472 VPB.n471 13.653
R579 VPB.n471 VPB.n470 13.653
R580 VPB.n477 VPB.n476 13.653
R581 VPB.n476 VPB.n475 13.653
R582 VPB.n481 VPB.n480 13.653
R583 VPB.n480 VPB.n479 13.653
R584 VPB.n485 VPB.n484 13.653
R585 VPB.n484 VPB.n483 13.653
R586 VPB.n512 VPB.n511 13.653
R587 VPB.n511 VPB.n510 13.653
R588 VPB.n516 VPB.n515 13.653
R589 VPB.n515 VPB.n514 13.653
R590 VPB.n521 VPB.n520 13.653
R591 VPB.n520 VPB.n519 13.653
R592 VPB.n526 VPB.n525 13.653
R593 VPB.n525 VPB.n524 13.653
R594 VPB.n533 VPB.n532 13.653
R595 VPB.n532 VPB.n531 13.653
R596 VPB.n538 VPB.n537 13.653
R597 VPB.n537 VPB.n536 13.653
R598 VPB.n543 VPB.n542 13.653
R599 VPB.n542 VPB.n541 13.653
R600 VPB.n550 VPB.n549 13.653
R601 VPB.n549 VPB.n548 13.653
R602 VPB.n555 VPB.n554 13.653
R603 VPB.n554 VPB.n553 13.653
R604 VPB.n560 VPB.n559 13.653
R605 VPB.n559 VPB.n558 13.653
R606 VPB.n564 VPB.n563 13.653
R607 VPB.n563 VPB.n562 13.653
R608 VPB.n568 VPB.n567 13.653
R609 VPB.n567 VPB.n566 13.653
R610 VPB.n595 VPB.n594 13.653
R611 VPB.n594 VPB.n593 13.653
R612 VPB.n600 VPB.n599 13.653
R613 VPB.n599 VPB.n598 13.653
R614 VPB.n605 VPB.n604 13.653
R615 VPB.n604 VPB.n603 13.653
R616 VPB.n612 VPB.n611 13.653
R617 VPB.n611 VPB.n610 13.653
R618 VPB.n617 VPB.n616 13.653
R619 VPB.n616 VPB.n615 13.653
R620 VPB.n622 VPB.n621 13.653
R621 VPB.n621 VPB.n620 13.653
R622 VPB.n627 VPB.n626 13.653
R623 VPB.n626 VPB.n625 13.653
R624 VPB.n631 VPB.n630 13.653
R625 VPB.n630 VPB.n629 13.653
R626 VPB.n658 VPB.n657 13.653
R627 VPB.n657 VPB.n656 13.653
R628 VPB.n662 VPB.n661 13.653
R629 VPB.n661 VPB.n660 13.653
R630 VPB.n667 VPB.n666 13.653
R631 VPB.n666 VPB.n665 13.653
R632 VPB.n672 VPB.n671 13.653
R633 VPB.n671 VPB.n670 13.653
R634 VPB.n679 VPB.n678 13.653
R635 VPB.n678 VPB.n677 13.653
R636 VPB.n684 VPB.n683 13.653
R637 VPB.n683 VPB.n682 13.653
R638 VPB.n689 VPB.n688 13.653
R639 VPB.n688 VPB.n687 13.653
R640 VPB.n696 VPB.n695 13.653
R641 VPB.n695 VPB.n694 13.653
R642 VPB.n701 VPB.n700 13.653
R643 VPB.n700 VPB.n699 13.653
R644 VPB.n706 VPB.n705 13.653
R645 VPB.n705 VPB.n704 13.653
R646 VPB.n710 VPB.n709 13.653
R647 VPB.n709 VPB.n708 13.653
R648 VPB.n714 VPB.n713 13.653
R649 VPB.n713 VPB.n712 13.653
R650 VPB.n741 VPB.n740 13.653
R651 VPB.n740 VPB.n739 13.653
R652 VPB.n745 VPB.n744 13.653
R653 VPB.n744 VPB.n743 13.653
R654 VPB.n750 VPB.n749 13.653
R655 VPB.n749 VPB.n748 13.653
R656 VPB.n755 VPB.n754 13.653
R657 VPB.n754 VPB.n753 13.653
R658 VPB.n762 VPB.n761 13.653
R659 VPB.n761 VPB.n760 13.653
R660 VPB.n767 VPB.n766 13.653
R661 VPB.n766 VPB.n765 13.653
R662 VPB.n772 VPB.n771 13.653
R663 VPB.n771 VPB.n770 13.653
R664 VPB.n779 VPB.n778 13.653
R665 VPB.n778 VPB.n777 13.653
R666 VPB.n784 VPB.n783 13.653
R667 VPB.n783 VPB.n782 13.653
R668 VPB.n789 VPB.n788 13.653
R669 VPB.n788 VPB.n787 13.653
R670 VPB.n793 VPB.n792 13.653
R671 VPB.n792 VPB.n791 13.653
R672 VPB.n797 VPB.n796 13.653
R673 VPB.n796 VPB.n795 13.653
R674 VPB.n824 VPB.n823 13.653
R675 VPB.n823 VPB.n822 13.653
R676 VPB.n829 VPB.n828 13.653
R677 VPB.n828 VPB.n827 13.653
R678 VPB.n834 VPB.n833 13.653
R679 VPB.n833 VPB.n832 13.653
R680 VPB.n841 VPB.n840 13.653
R681 VPB.n840 VPB.n839 13.653
R682 VPB.n846 VPB.n845 13.653
R683 VPB.n845 VPB.n844 13.653
R684 VPB.n851 VPB.n850 13.653
R685 VPB.n850 VPB.n849 13.653
R686 VPB.n856 VPB.n855 13.653
R687 VPB.n855 VPB.n854 13.653
R688 VPB.n860 VPB.n859 13.653
R689 VPB.n859 VPB.n858 13.653
R690 VPB.n130 VPB.n129 13.653
R691 VPB.n129 VPB.n128 13.653
R692 VPB.n133 VPB.n132 13.653
R693 VPB.n132 VPB.n131 13.653
R694 VPB.n137 VPB.n136 13.653
R695 VPB.n136 VPB.n135 13.653
R696 VPB.n141 VPB.n140 13.653
R697 VPB.n140 VPB.n139 13.653
R698 VPB.n145 VPB.n144 13.653
R699 VPB.n144 VPB.n143 13.653
R700 VPB.n150 VPB.n149 13.653
R701 VPB.n149 VPB.n148 13.653
R702 VPB.n154 VPB.n153 13.653
R703 VPB.n153 VPB.n152 13.653
R704 VPB.n159 VPB.n158 13.653
R705 VPB.n158 VPB.n157 13.653
R706 VPB.n163 VPB.n162 13.653
R707 VPB.n162 VPB.n161 13.653
R708 VPB.n166 VPB.n165 13.653
R709 VPB.n165 VPB.n164 13.653
R710 VPB.n170 VPB.n169 13.653
R711 VPB.n169 VPB.n168 13.653
R712 VPB.n876 VPB.n875 13.653
R713 VPB.n875 VPB.n874 13.653
R714 VPB.n881 VPB.n880 13.653
R715 VPB.n880 VPB.n879 13.653
R716 VPB.n885 VPB.n884 13.653
R717 VPB.n884 VPB.n883 13.653
R718 VPB.n890 VPB.n889 13.653
R719 VPB.n889 VPB.n888 13.653
R720 VPB.n895 VPB.n894 13.653
R721 VPB.n894 VPB.n893 13.653
R722 VPB.n902 VPB.n901 13.653
R723 VPB.n901 VPB.n900 13.653
R724 VPB.n907 VPB.n906 13.653
R725 VPB.n906 VPB.n905 13.653
R726 VPB.n912 VPB.n911 13.653
R727 VPB.n911 VPB.n910 13.653
R728 VPB.n919 VPB.n918 13.653
R729 VPB.n918 VPB.n917 13.653
R730 VPB.n924 VPB.n923 13.653
R731 VPB.n923 VPB.n922 13.653
R732 VPB.n929 VPB.n928 13.653
R733 VPB.n928 VPB.n927 13.653
R734 VPB.n933 VPB.n932 13.653
R735 VPB.n932 VPB.n931 13.653
R736 VPB.n937 VPB.n936 13.653
R737 VPB.n936 VPB.n935 13.653
R738 VPB.n964 VPB.n963 13.653
R739 VPB.n963 VPB.n962 13.653
R740 VPB.n969 VPB.n968 13.653
R741 VPB.n968 VPB.n967 13.653
R742 VPB.n974 VPB.n973 13.653
R743 VPB.n973 VPB.n972 13.653
R744 VPB.n981 VPB.n980 13.653
R745 VPB.n980 VPB.n979 13.653
R746 VPB.n986 VPB.n985 13.653
R747 VPB.n985 VPB.n984 13.653
R748 VPB.n991 VPB.n990 13.653
R749 VPB.n990 VPB.n989 13.653
R750 VPB.n996 VPB.n995 13.653
R751 VPB.n995 VPB.n994 13.653
R752 VPB.n1000 VPB.n999 13.653
R753 VPB.n999 VPB.n998 13.653
R754 VPB.n1027 VPB.n1026 13.653
R755 VPB.n1026 VPB.n1025 13.653
R756 VPB.n1031 VPB.n1030 13.653
R757 VPB.n1030 VPB.n1029 13.653
R758 VPB.n1036 VPB.n1035 13.653
R759 VPB.n1035 VPB.n1034 13.653
R760 VPB.n1041 VPB.n1040 13.653
R761 VPB.n1040 VPB.n1039 13.653
R762 VPB.n1048 VPB.n1047 13.653
R763 VPB.n1047 VPB.n1046 13.653
R764 VPB.n1053 VPB.n1052 13.653
R765 VPB.n1052 VPB.n1051 13.653
R766 VPB.n1058 VPB.n1057 13.653
R767 VPB.n1057 VPB.n1056 13.653
R768 VPB.n1065 VPB.n1064 13.653
R769 VPB.n1064 VPB.n1063 13.653
R770 VPB.n1070 VPB.n1069 13.653
R771 VPB.n1069 VPB.n1068 13.653
R772 VPB.n1075 VPB.n1074 13.653
R773 VPB.n1074 VPB.n1073 13.653
R774 VPB.n1079 VPB.n1078 13.653
R775 VPB.n1078 VPB.n1077 13.653
R776 VPB.n1083 VPB.n1082 13.653
R777 VPB.n1082 VPB.n1081 13.653
R778 VPB.n1110 VPB.n1109 13.653
R779 VPB.n1109 VPB.n1108 13.653
R780 VPB.n1114 VPB.n1113 13.653
R781 VPB.n1113 VPB.n1112 13.653
R782 VPB.n1119 VPB.n1118 13.653
R783 VPB.n1118 VPB.n1117 13.653
R784 VPB.n1124 VPB.n1123 13.653
R785 VPB.n1123 VPB.n1122 13.653
R786 VPB.n1131 VPB.n1130 13.653
R787 VPB.n1130 VPB.n1129 13.653
R788 VPB.n1136 VPB.n1135 13.653
R789 VPB.n1135 VPB.n1134 13.653
R790 VPB.n1141 VPB.n1140 13.653
R791 VPB.n1140 VPB.n1139 13.653
R792 VPB.n1148 VPB.n1147 13.653
R793 VPB.n1147 VPB.n1146 13.653
R794 VPB.n1153 VPB.n1152 13.653
R795 VPB.n1152 VPB.n1151 13.653
R796 VPB.n1158 VPB.n1157 13.653
R797 VPB.n1157 VPB.n1156 13.653
R798 VPB.n1162 VPB.n1161 13.653
R799 VPB.n1161 VPB.n1160 13.653
R800 VPB.n1166 VPB.n1165 13.653
R801 VPB.n1165 VPB.n1164 13.653
R802 VPB.n1193 VPB.n1192 13.653
R803 VPB.n1192 VPB.n1191 13.653
R804 VPB.n1198 VPB.n1197 13.653
R805 VPB.n1197 VPB.n1196 13.653
R806 VPB.n1203 VPB.n1202 13.653
R807 VPB.n1202 VPB.n1201 13.653
R808 VPB.n1210 VPB.n1209 13.653
R809 VPB.n1209 VPB.n1208 13.653
R810 VPB.n1215 VPB.n1214 13.653
R811 VPB.n1214 VPB.n1213 13.653
R812 VPB.n1220 VPB.n1219 13.653
R813 VPB.n1219 VPB.n1218 13.653
R814 VPB.n1225 VPB.n1224 13.653
R815 VPB.n1224 VPB.n1223 13.653
R816 VPB.n1229 VPB.n1228 13.653
R817 VPB.n1228 VPB.n1227 13.653
R818 VPB.n1256 VPB.n1255 13.653
R819 VPB.n1255 VPB.n1254 13.653
R820 VPB.n1260 VPB.n1259 13.653
R821 VPB.n1259 VPB.n1258 13.653
R822 VPB.n1265 VPB.n1264 13.653
R823 VPB.n1264 VPB.n1263 13.653
R824 VPB.n1270 VPB.n1269 13.653
R825 VPB.n1269 VPB.n1268 13.653
R826 VPB.n1277 VPB.n1276 13.653
R827 VPB.n1276 VPB.n1275 13.653
R828 VPB.n1282 VPB.n1281 13.653
R829 VPB.n1281 VPB.n1280 13.653
R830 VPB.n1287 VPB.n1286 13.653
R831 VPB.n1286 VPB.n1285 13.653
R832 VPB.n1294 VPB.n1293 13.653
R833 VPB.n1293 VPB.n1292 13.653
R834 VPB.n1299 VPB.n1298 13.653
R835 VPB.n1298 VPB.n1297 13.653
R836 VPB.n1304 VPB.n1303 13.653
R837 VPB.n1303 VPB.n1302 13.653
R838 VPB.n1308 VPB.n1307 13.653
R839 VPB.n1307 VPB.n1306 13.653
R840 VPB.n1312 VPB.n1311 13.653
R841 VPB.n1311 VPB.n1310 13.653
R842 VPB.n1339 VPB.n1338 13.653
R843 VPB.n1338 VPB.n1337 13.653
R844 VPB.n1343 VPB.n1342 13.653
R845 VPB.n1342 VPB.n1341 13.653
R846 VPB.n1348 VPB.n1347 13.653
R847 VPB.n1347 VPB.n1346 13.653
R848 VPB.n1353 VPB.n1352 13.653
R849 VPB.n1352 VPB.n1351 13.653
R850 VPB.n1360 VPB.n1359 13.653
R851 VPB.n1359 VPB.n1358 13.653
R852 VPB.n1365 VPB.n1364 13.653
R853 VPB.n1364 VPB.n1363 13.653
R854 VPB.n1370 VPB.n1369 13.653
R855 VPB.n1369 VPB.n1368 13.653
R856 VPB.n1377 VPB.n1376 13.653
R857 VPB.n1376 VPB.n1375 13.653
R858 VPB.n1382 VPB.n1381 13.653
R859 VPB.n1381 VPB.n1380 13.653
R860 VPB.n1387 VPB.n1386 13.653
R861 VPB.n1386 VPB.n1385 13.653
R862 VPB.n1391 VPB.n1390 13.653
R863 VPB.n1390 VPB.n1389 13.653
R864 VPB.n1395 VPB.n1394 13.653
R865 VPB.n1394 VPB.n1393 13.653
R866 VPB.n1422 VPB.n1421 13.653
R867 VPB.n1421 VPB.n1420 13.653
R868 VPB.n1427 VPB.n1426 13.653
R869 VPB.n1426 VPB.n1425 13.653
R870 VPB.n1432 VPB.n1431 13.653
R871 VPB.n1431 VPB.n1430 13.653
R872 VPB.n1439 VPB.n1438 13.653
R873 VPB.n1438 VPB.n1437 13.653
R874 VPB.n1444 VPB.n1443 13.653
R875 VPB.n1443 VPB.n1442 13.653
R876 VPB.n1449 VPB.n1448 13.653
R877 VPB.n1448 VPB.n1447 13.653
R878 VPB.n1454 VPB.n1453 13.653
R879 VPB.n1453 VPB.n1452 13.653
R880 VPB.n1458 VPB.n1457 13.653
R881 VPB.n1457 VPB.n1456 13.653
R882 VPB.n1485 VPB.n1484 13.653
R883 VPB.n1484 VPB.n1483 13.653
R884 VPB.n1489 VPB.n1488 13.653
R885 VPB.n1488 VPB.n1487 13.653
R886 VPB.n1494 VPB.n1493 13.653
R887 VPB.n1493 VPB.n1492 13.653
R888 VPB.n1499 VPB.n1498 13.653
R889 VPB.n1498 VPB.n1497 13.653
R890 VPB.n1506 VPB.n1505 13.653
R891 VPB.n1505 VPB.n1504 13.653
R892 VPB.n1511 VPB.n1510 13.653
R893 VPB.n1510 VPB.n1509 13.653
R894 VPB.n1516 VPB.n1515 13.653
R895 VPB.n1515 VPB.n1514 13.653
R896 VPB.n1523 VPB.n1522 13.653
R897 VPB.n1522 VPB.n1521 13.653
R898 VPB.n1528 VPB.n1527 13.653
R899 VPB.n1527 VPB.n1526 13.653
R900 VPB.n1533 VPB.n1532 13.653
R901 VPB.n1532 VPB.n1531 13.653
R902 VPB.n1537 VPB.n1536 13.653
R903 VPB.n1536 VPB.n1535 13.653
R904 VPB.n1541 VPB.n1540 13.653
R905 VPB.n1540 VPB.n1539 13.653
R906 VPB.n41 VPB.n40 13.653
R907 VPB.n40 VPB.n39 13.653
R908 VPB.n44 VPB.n43 13.653
R909 VPB.n43 VPB.n42 13.653
R910 VPB.n48 VPB.n47 13.653
R911 VPB.n47 VPB.n46 13.653
R912 VPB.n52 VPB.n51 13.653
R913 VPB.n51 VPB.n50 13.653
R914 VPB.n56 VPB.n55 13.653
R915 VPB.n55 VPB.n54 13.653
R916 VPB.n61 VPB.n60 13.653
R917 VPB.n60 VPB.n59 13.653
R918 VPB.n65 VPB.n64 13.653
R919 VPB.n64 VPB.n63 13.653
R920 VPB.n70 VPB.n69 13.653
R921 VPB.n69 VPB.n68 13.653
R922 VPB.n74 VPB.n73 13.653
R923 VPB.n73 VPB.n72 13.653
R924 VPB.n77 VPB.n76 13.653
R925 VPB.n76 VPB.n75 13.653
R926 VPB.n81 VPB.n80 13.653
R927 VPB.n80 VPB.n79 13.653
R928 VPB.n1555 VPB.n0 13.653
R929 VPB VPB.n0 13.653
R930 VPB.n323 VPB.n322 13.35
R931 VPB.n386 VPB.n385 13.35
R932 VPB.n458 VPB.n457 13.35
R933 VPB.n541 VPB.n540 13.35
R934 VPB.n615 VPB.n614 13.35
R935 VPB.n687 VPB.n686 13.35
R936 VPB.n770 VPB.n769 13.35
R937 VPB.n844 VPB.n843 13.35
R938 VPB.n152 VPB.n151 13.35
R939 VPB.n910 VPB.n909 13.35
R940 VPB.n984 VPB.n983 13.35
R941 VPB.n1056 VPB.n1055 13.35
R942 VPB.n1139 VPB.n1138 13.35
R943 VPB.n1213 VPB.n1212 13.35
R944 VPB.n1285 VPB.n1284 13.35
R945 VPB.n1368 VPB.n1367 13.35
R946 VPB.n1442 VPB.n1441 13.35
R947 VPB.n1514 VPB.n1513 13.35
R948 VPB.n63 VPB.n62 13.35
R949 VPB.n1559 VPB.n1558 13.276
R950 VPB.n1558 VPB.n1556 13.276
R951 VPB.n36 VPB.n18 13.276
R952 VPB.n18 VPB.n16 13.276
R953 VPB.n1480 VPB.n1462 13.276
R954 VPB.n1462 VPB.n1460 13.276
R955 VPB.n1417 VPB.n1399 13.276
R956 VPB.n1399 VPB.n1397 13.276
R957 VPB.n1334 VPB.n1316 13.276
R958 VPB.n1316 VPB.n1314 13.276
R959 VPB.n1251 VPB.n1233 13.276
R960 VPB.n1233 VPB.n1231 13.276
R961 VPB.n1188 VPB.n1170 13.276
R962 VPB.n1170 VPB.n1168 13.276
R963 VPB.n1105 VPB.n1087 13.276
R964 VPB.n1087 VPB.n1085 13.276
R965 VPB.n1022 VPB.n1004 13.276
R966 VPB.n1004 VPB.n1002 13.276
R967 VPB.n959 VPB.n941 13.276
R968 VPB.n941 VPB.n939 13.276
R969 VPB.n102 VPB.n84 13.276
R970 VPB.n84 VPB.n82 13.276
R971 VPB.n125 VPB.n107 13.276
R972 VPB.n107 VPB.n105 13.276
R973 VPB.n819 VPB.n801 13.276
R974 VPB.n801 VPB.n799 13.276
R975 VPB.n736 VPB.n718 13.276
R976 VPB.n718 VPB.n716 13.276
R977 VPB.n653 VPB.n635 13.276
R978 VPB.n635 VPB.n633 13.276
R979 VPB.n590 VPB.n572 13.276
R980 VPB.n572 VPB.n570 13.276
R981 VPB.n507 VPB.n489 13.276
R982 VPB.n489 VPB.n487 13.276
R983 VPB.n424 VPB.n406 13.276
R984 VPB.n406 VPB.n404 13.276
R985 VPB.n361 VPB.n343 13.276
R986 VPB.n343 VPB.n341 13.276
R987 VPB.n298 VPB.n280 13.276
R988 VPB.n280 VPB.n278 13.276
R989 VPB.n243 VPB.n225 13.276
R990 VPB.n225 VPB.n223 13.276
R991 VPB.n203 VPB.n200 13.276
R992 VPB.n200 VPB.n197 13.276
R993 VPB.n248 VPB.n244 13.276
R994 VPB.n303 VPB.n299 13.276
R995 VPB.n366 VPB.n362 13.276
R996 VPB.n429 VPB.n425 13.276
R997 VPB.n512 VPB.n508 13.276
R998 VPB.n595 VPB.n591 13.276
R999 VPB.n658 VPB.n654 13.276
R1000 VPB.n741 VPB.n737 13.276
R1001 VPB.n824 VPB.n820 13.276
R1002 VPB.n130 VPB.n126 13.276
R1003 VPB.n133 VPB.n130 13.276
R1004 VPB.n141 VPB.n137 13.276
R1005 VPB.n145 VPB.n141 13.276
R1006 VPB.n154 VPB.n150 13.276
R1007 VPB.n163 VPB.n159 13.276
R1008 VPB.n166 VPB.n163 13.276
R1009 VPB.n876 VPB.n170 13.276
R1010 VPB.n877 VPB.n876 13.276
R1011 VPB.n881 VPB.n877 13.276
R1012 VPB.n964 VPB.n960 13.276
R1013 VPB.n1027 VPB.n1023 13.276
R1014 VPB.n1110 VPB.n1106 13.276
R1015 VPB.n1193 VPB.n1189 13.276
R1016 VPB.n1256 VPB.n1252 13.276
R1017 VPB.n1339 VPB.n1335 13.276
R1018 VPB.n1422 VPB.n1418 13.276
R1019 VPB.n1485 VPB.n1481 13.276
R1020 VPB.n41 VPB.n37 13.276
R1021 VPB.n44 VPB.n41 13.276
R1022 VPB.n52 VPB.n48 13.276
R1023 VPB.n56 VPB.n52 13.276
R1024 VPB.n65 VPB.n61 13.276
R1025 VPB.n74 VPB.n70 13.276
R1026 VPB.n77 VPB.n74 13.276
R1027 VPB.n1555 VPB.n81 13.276
R1028 VPB.n191 VPB.n173 13.276
R1029 VPB.n173 VPB.n171 13.276
R1030 VPB.n178 VPB.n176 12.796
R1031 VPB.n178 VPB.n177 12.564
R1032 VPB.n170 VPB.n167 12.558
R1033 VPB.n81 VPB.n78 12.558
R1034 VPB.n134 VPB.n133 12.2
R1035 VPB.n45 VPB.n44 12.2
R1036 VPB.n186 VPB.n185 12.198
R1037 VPB.n186 VPB.n183 12.198
R1038 VPB.n181 VPB.n180 12.198
R1039 VPB.n150 VPB.n146 9.329
R1040 VPB.n61 VPB.n57 9.329
R1041 VPB.n155 VPB.n154 8.97
R1042 VPB.n66 VPB.n65 8.97
R1043 VPB.n191 VPB.n190 7.5
R1044 VPB.n176 VPB.n175 7.5
R1045 VPB.n180 VPB.n179 7.5
R1046 VPB.n185 VPB.n184 7.5
R1047 VPB.n173 VPB.n172 7.5
R1048 VPB.n188 VPB.n174 7.5
R1049 VPB.n225 VPB.n224 7.5
R1050 VPB.n238 VPB.n237 7.5
R1051 VPB.n232 VPB.n231 7.5
R1052 VPB.n234 VPB.n233 7.5
R1053 VPB.n227 VPB.n226 7.5
R1054 VPB.n243 VPB.n242 7.5
R1055 VPB.n280 VPB.n279 7.5
R1056 VPB.n293 VPB.n292 7.5
R1057 VPB.n287 VPB.n286 7.5
R1058 VPB.n289 VPB.n288 7.5
R1059 VPB.n282 VPB.n281 7.5
R1060 VPB.n298 VPB.n297 7.5
R1061 VPB.n343 VPB.n342 7.5
R1062 VPB.n356 VPB.n355 7.5
R1063 VPB.n350 VPB.n349 7.5
R1064 VPB.n352 VPB.n351 7.5
R1065 VPB.n345 VPB.n344 7.5
R1066 VPB.n361 VPB.n360 7.5
R1067 VPB.n406 VPB.n405 7.5
R1068 VPB.n419 VPB.n418 7.5
R1069 VPB.n413 VPB.n412 7.5
R1070 VPB.n415 VPB.n414 7.5
R1071 VPB.n408 VPB.n407 7.5
R1072 VPB.n424 VPB.n423 7.5
R1073 VPB.n489 VPB.n488 7.5
R1074 VPB.n502 VPB.n501 7.5
R1075 VPB.n496 VPB.n495 7.5
R1076 VPB.n498 VPB.n497 7.5
R1077 VPB.n491 VPB.n490 7.5
R1078 VPB.n507 VPB.n506 7.5
R1079 VPB.n572 VPB.n571 7.5
R1080 VPB.n585 VPB.n584 7.5
R1081 VPB.n579 VPB.n578 7.5
R1082 VPB.n581 VPB.n580 7.5
R1083 VPB.n574 VPB.n573 7.5
R1084 VPB.n590 VPB.n589 7.5
R1085 VPB.n635 VPB.n634 7.5
R1086 VPB.n648 VPB.n647 7.5
R1087 VPB.n642 VPB.n641 7.5
R1088 VPB.n644 VPB.n643 7.5
R1089 VPB.n637 VPB.n636 7.5
R1090 VPB.n653 VPB.n652 7.5
R1091 VPB.n718 VPB.n717 7.5
R1092 VPB.n731 VPB.n730 7.5
R1093 VPB.n725 VPB.n724 7.5
R1094 VPB.n727 VPB.n726 7.5
R1095 VPB.n720 VPB.n719 7.5
R1096 VPB.n736 VPB.n735 7.5
R1097 VPB.n801 VPB.n800 7.5
R1098 VPB.n814 VPB.n813 7.5
R1099 VPB.n808 VPB.n807 7.5
R1100 VPB.n810 VPB.n809 7.5
R1101 VPB.n803 VPB.n802 7.5
R1102 VPB.n819 VPB.n818 7.5
R1103 VPB.n107 VPB.n106 7.5
R1104 VPB.n120 VPB.n119 7.5
R1105 VPB.n114 VPB.n113 7.5
R1106 VPB.n116 VPB.n115 7.5
R1107 VPB.n109 VPB.n108 7.5
R1108 VPB.n125 VPB.n124 7.5
R1109 VPB.n84 VPB.n83 7.5
R1110 VPB.n97 VPB.n96 7.5
R1111 VPB.n91 VPB.n90 7.5
R1112 VPB.n93 VPB.n92 7.5
R1113 VPB.n86 VPB.n85 7.5
R1114 VPB.n102 VPB.n101 7.5
R1115 VPB.n941 VPB.n940 7.5
R1116 VPB.n954 VPB.n953 7.5
R1117 VPB.n948 VPB.n947 7.5
R1118 VPB.n950 VPB.n949 7.5
R1119 VPB.n943 VPB.n942 7.5
R1120 VPB.n959 VPB.n958 7.5
R1121 VPB.n1004 VPB.n1003 7.5
R1122 VPB.n1017 VPB.n1016 7.5
R1123 VPB.n1011 VPB.n1010 7.5
R1124 VPB.n1013 VPB.n1012 7.5
R1125 VPB.n1006 VPB.n1005 7.5
R1126 VPB.n1022 VPB.n1021 7.5
R1127 VPB.n1087 VPB.n1086 7.5
R1128 VPB.n1100 VPB.n1099 7.5
R1129 VPB.n1094 VPB.n1093 7.5
R1130 VPB.n1096 VPB.n1095 7.5
R1131 VPB.n1089 VPB.n1088 7.5
R1132 VPB.n1105 VPB.n1104 7.5
R1133 VPB.n1170 VPB.n1169 7.5
R1134 VPB.n1183 VPB.n1182 7.5
R1135 VPB.n1177 VPB.n1176 7.5
R1136 VPB.n1179 VPB.n1178 7.5
R1137 VPB.n1172 VPB.n1171 7.5
R1138 VPB.n1188 VPB.n1187 7.5
R1139 VPB.n1233 VPB.n1232 7.5
R1140 VPB.n1246 VPB.n1245 7.5
R1141 VPB.n1240 VPB.n1239 7.5
R1142 VPB.n1242 VPB.n1241 7.5
R1143 VPB.n1235 VPB.n1234 7.5
R1144 VPB.n1251 VPB.n1250 7.5
R1145 VPB.n1316 VPB.n1315 7.5
R1146 VPB.n1329 VPB.n1328 7.5
R1147 VPB.n1323 VPB.n1322 7.5
R1148 VPB.n1325 VPB.n1324 7.5
R1149 VPB.n1318 VPB.n1317 7.5
R1150 VPB.n1334 VPB.n1333 7.5
R1151 VPB.n1399 VPB.n1398 7.5
R1152 VPB.n1412 VPB.n1411 7.5
R1153 VPB.n1406 VPB.n1405 7.5
R1154 VPB.n1408 VPB.n1407 7.5
R1155 VPB.n1401 VPB.n1400 7.5
R1156 VPB.n1417 VPB.n1416 7.5
R1157 VPB.n1462 VPB.n1461 7.5
R1158 VPB.n1475 VPB.n1474 7.5
R1159 VPB.n1469 VPB.n1468 7.5
R1160 VPB.n1471 VPB.n1470 7.5
R1161 VPB.n1464 VPB.n1463 7.5
R1162 VPB.n1480 VPB.n1479 7.5
R1163 VPB.n18 VPB.n17 7.5
R1164 VPB.n31 VPB.n30 7.5
R1165 VPB.n25 VPB.n24 7.5
R1166 VPB.n27 VPB.n26 7.5
R1167 VPB.n20 VPB.n19 7.5
R1168 VPB.n36 VPB.n35 7.5
R1169 VPB.n1558 VPB.n1557 7.5
R1170 VPB.n12 VPB.n11 7.5
R1171 VPB.n6 VPB.n5 7.5
R1172 VPB.n8 VPB.n7 7.5
R1173 VPB.n2 VPB.n1 7.5
R1174 VPB.n1560 VPB.n1559 7.5
R1175 VPB.n37 VPB.n36 7.176
R1176 VPB.n1481 VPB.n1480 7.176
R1177 VPB.n1418 VPB.n1417 7.176
R1178 VPB.n1335 VPB.n1334 7.176
R1179 VPB.n1252 VPB.n1251 7.176
R1180 VPB.n1189 VPB.n1188 7.176
R1181 VPB.n1106 VPB.n1105 7.176
R1182 VPB.n1023 VPB.n1022 7.176
R1183 VPB.n960 VPB.n959 7.176
R1184 VPB.n877 VPB.n102 7.176
R1185 VPB.n126 VPB.n125 7.176
R1186 VPB.n820 VPB.n819 7.176
R1187 VPB.n737 VPB.n736 7.176
R1188 VPB.n654 VPB.n653 7.176
R1189 VPB.n591 VPB.n590 7.176
R1190 VPB.n508 VPB.n507 7.176
R1191 VPB.n425 VPB.n424 7.176
R1192 VPB.n362 VPB.n361 7.176
R1193 VPB.n299 VPB.n298 7.176
R1194 VPB.n244 VPB.n243 7.176
R1195 VPB.n239 VPB.n236 6.729
R1196 VPB.n235 VPB.n232 6.729
R1197 VPB.n230 VPB.n227 6.729
R1198 VPB.n294 VPB.n291 6.729
R1199 VPB.n290 VPB.n287 6.729
R1200 VPB.n285 VPB.n282 6.729
R1201 VPB.n357 VPB.n354 6.729
R1202 VPB.n353 VPB.n350 6.729
R1203 VPB.n348 VPB.n345 6.729
R1204 VPB.n420 VPB.n417 6.729
R1205 VPB.n416 VPB.n413 6.729
R1206 VPB.n411 VPB.n408 6.729
R1207 VPB.n503 VPB.n500 6.729
R1208 VPB.n499 VPB.n496 6.729
R1209 VPB.n494 VPB.n491 6.729
R1210 VPB.n586 VPB.n583 6.729
R1211 VPB.n582 VPB.n579 6.729
R1212 VPB.n577 VPB.n574 6.729
R1213 VPB.n649 VPB.n646 6.729
R1214 VPB.n645 VPB.n642 6.729
R1215 VPB.n640 VPB.n637 6.729
R1216 VPB.n732 VPB.n729 6.729
R1217 VPB.n728 VPB.n725 6.729
R1218 VPB.n723 VPB.n720 6.729
R1219 VPB.n815 VPB.n812 6.729
R1220 VPB.n811 VPB.n808 6.729
R1221 VPB.n806 VPB.n803 6.729
R1222 VPB.n121 VPB.n118 6.729
R1223 VPB.n117 VPB.n114 6.729
R1224 VPB.n112 VPB.n109 6.729
R1225 VPB.n98 VPB.n95 6.729
R1226 VPB.n94 VPB.n91 6.729
R1227 VPB.n89 VPB.n86 6.729
R1228 VPB.n955 VPB.n952 6.729
R1229 VPB.n951 VPB.n948 6.729
R1230 VPB.n946 VPB.n943 6.729
R1231 VPB.n1018 VPB.n1015 6.729
R1232 VPB.n1014 VPB.n1011 6.729
R1233 VPB.n1009 VPB.n1006 6.729
R1234 VPB.n1101 VPB.n1098 6.729
R1235 VPB.n1097 VPB.n1094 6.729
R1236 VPB.n1092 VPB.n1089 6.729
R1237 VPB.n1184 VPB.n1181 6.729
R1238 VPB.n1180 VPB.n1177 6.729
R1239 VPB.n1175 VPB.n1172 6.729
R1240 VPB.n1247 VPB.n1244 6.729
R1241 VPB.n1243 VPB.n1240 6.729
R1242 VPB.n1238 VPB.n1235 6.729
R1243 VPB.n1330 VPB.n1327 6.729
R1244 VPB.n1326 VPB.n1323 6.729
R1245 VPB.n1321 VPB.n1318 6.729
R1246 VPB.n1413 VPB.n1410 6.729
R1247 VPB.n1409 VPB.n1406 6.729
R1248 VPB.n1404 VPB.n1401 6.729
R1249 VPB.n1476 VPB.n1473 6.729
R1250 VPB.n1472 VPB.n1469 6.729
R1251 VPB.n1467 VPB.n1464 6.729
R1252 VPB.n32 VPB.n29 6.729
R1253 VPB.n28 VPB.n25 6.729
R1254 VPB.n23 VPB.n20 6.729
R1255 VPB.n13 VPB.n10 6.729
R1256 VPB.n9 VPB.n6 6.729
R1257 VPB.n4 VPB.n2 6.729
R1258 VPB.n230 VPB.n229 6.728
R1259 VPB.n235 VPB.n234 6.728
R1260 VPB.n239 VPB.n238 6.728
R1261 VPB.n242 VPB.n241 6.728
R1262 VPB.n285 VPB.n284 6.728
R1263 VPB.n290 VPB.n289 6.728
R1264 VPB.n294 VPB.n293 6.728
R1265 VPB.n297 VPB.n296 6.728
R1266 VPB.n348 VPB.n347 6.728
R1267 VPB.n353 VPB.n352 6.728
R1268 VPB.n357 VPB.n356 6.728
R1269 VPB.n360 VPB.n359 6.728
R1270 VPB.n411 VPB.n410 6.728
R1271 VPB.n416 VPB.n415 6.728
R1272 VPB.n420 VPB.n419 6.728
R1273 VPB.n423 VPB.n422 6.728
R1274 VPB.n494 VPB.n493 6.728
R1275 VPB.n499 VPB.n498 6.728
R1276 VPB.n503 VPB.n502 6.728
R1277 VPB.n506 VPB.n505 6.728
R1278 VPB.n577 VPB.n576 6.728
R1279 VPB.n582 VPB.n581 6.728
R1280 VPB.n586 VPB.n585 6.728
R1281 VPB.n589 VPB.n588 6.728
R1282 VPB.n640 VPB.n639 6.728
R1283 VPB.n645 VPB.n644 6.728
R1284 VPB.n649 VPB.n648 6.728
R1285 VPB.n652 VPB.n651 6.728
R1286 VPB.n723 VPB.n722 6.728
R1287 VPB.n728 VPB.n727 6.728
R1288 VPB.n732 VPB.n731 6.728
R1289 VPB.n735 VPB.n734 6.728
R1290 VPB.n806 VPB.n805 6.728
R1291 VPB.n811 VPB.n810 6.728
R1292 VPB.n815 VPB.n814 6.728
R1293 VPB.n818 VPB.n817 6.728
R1294 VPB.n112 VPB.n111 6.728
R1295 VPB.n117 VPB.n116 6.728
R1296 VPB.n121 VPB.n120 6.728
R1297 VPB.n124 VPB.n123 6.728
R1298 VPB.n89 VPB.n88 6.728
R1299 VPB.n94 VPB.n93 6.728
R1300 VPB.n98 VPB.n97 6.728
R1301 VPB.n101 VPB.n100 6.728
R1302 VPB.n946 VPB.n945 6.728
R1303 VPB.n951 VPB.n950 6.728
R1304 VPB.n955 VPB.n954 6.728
R1305 VPB.n958 VPB.n957 6.728
R1306 VPB.n1009 VPB.n1008 6.728
R1307 VPB.n1014 VPB.n1013 6.728
R1308 VPB.n1018 VPB.n1017 6.728
R1309 VPB.n1021 VPB.n1020 6.728
R1310 VPB.n1092 VPB.n1091 6.728
R1311 VPB.n1097 VPB.n1096 6.728
R1312 VPB.n1101 VPB.n1100 6.728
R1313 VPB.n1104 VPB.n1103 6.728
R1314 VPB.n1175 VPB.n1174 6.728
R1315 VPB.n1180 VPB.n1179 6.728
R1316 VPB.n1184 VPB.n1183 6.728
R1317 VPB.n1187 VPB.n1186 6.728
R1318 VPB.n1238 VPB.n1237 6.728
R1319 VPB.n1243 VPB.n1242 6.728
R1320 VPB.n1247 VPB.n1246 6.728
R1321 VPB.n1250 VPB.n1249 6.728
R1322 VPB.n1321 VPB.n1320 6.728
R1323 VPB.n1326 VPB.n1325 6.728
R1324 VPB.n1330 VPB.n1329 6.728
R1325 VPB.n1333 VPB.n1332 6.728
R1326 VPB.n1404 VPB.n1403 6.728
R1327 VPB.n1409 VPB.n1408 6.728
R1328 VPB.n1413 VPB.n1412 6.728
R1329 VPB.n1416 VPB.n1415 6.728
R1330 VPB.n1467 VPB.n1466 6.728
R1331 VPB.n1472 VPB.n1471 6.728
R1332 VPB.n1476 VPB.n1475 6.728
R1333 VPB.n1479 VPB.n1478 6.728
R1334 VPB.n23 VPB.n22 6.728
R1335 VPB.n28 VPB.n27 6.728
R1336 VPB.n32 VPB.n31 6.728
R1337 VPB.n35 VPB.n34 6.728
R1338 VPB.n4 VPB.n3 6.728
R1339 VPB.n9 VPB.n8 6.728
R1340 VPB.n13 VPB.n12 6.728
R1341 VPB.n1561 VPB.n1560 6.728
R1342 VPB.n320 VPB.n316 6.458
R1343 VPB.n383 VPB.n379 6.458
R1344 VPB.n612 VPB.n608 6.458
R1345 VPB.n841 VPB.n837 6.458
R1346 VPB.n981 VPB.n977 6.458
R1347 VPB.n1210 VPB.n1206 6.458
R1348 VPB.n1439 VPB.n1435 6.458
R1349 VPB.n190 VPB.n189 6.398
R1350 VPB.n204 VPB.n194 6.112
R1351 VPB.n204 VPB.n203 6.101
R1352 VPB.n467 VPB.n463 4.305
R1353 VPB.n550 VPB.n546 4.305
R1354 VPB.n696 VPB.n692 4.305
R1355 VPB.n779 VPB.n775 4.305
R1356 VPB.n159 VPB.n155 4.305
R1357 VPB.n919 VPB.n915 4.305
R1358 VPB.n1065 VPB.n1061 4.305
R1359 VPB.n1148 VPB.n1144 4.305
R1360 VPB.n1294 VPB.n1290 4.305
R1361 VPB.n1377 VPB.n1373 4.305
R1362 VPB.n1523 VPB.n1519 4.305
R1363 VPB.n70 VPB.n66 4.305
R1364 VPB.n450 VPB.n446 3.947
R1365 VPB.n533 VPB.n529 3.947
R1366 VPB.n679 VPB.n675 3.947
R1367 VPB.n762 VPB.n758 3.947
R1368 VPB.n146 VPB.n145 3.947
R1369 VPB.n902 VPB.n898 3.947
R1370 VPB.n1048 VPB.n1044 3.947
R1371 VPB.n1131 VPB.n1127 3.947
R1372 VPB.n1277 VPB.n1273 3.947
R1373 VPB.n1360 VPB.n1356 3.947
R1374 VPB.n1506 VPB.n1502 3.947
R1375 VPB.n57 VPB.n56 3.947
R1376 VPB.n335 VPB.n332 1.794
R1377 VPB.n398 VPB.n395 1.794
R1378 VPB.n627 VPB.n624 1.794
R1379 VPB.n856 VPB.n853 1.794
R1380 VPB.n996 VPB.n993 1.794
R1381 VPB.n1225 VPB.n1222 1.794
R1382 VPB.n1454 VPB.n1451 1.794
R1383 VPB.n308 VPB.n305 1.435
R1384 VPB.n371 VPB.n368 1.435
R1385 VPB.n600 VPB.n597 1.435
R1386 VPB.n829 VPB.n826 1.435
R1387 VPB.n969 VPB.n966 1.435
R1388 VPB.n1198 VPB.n1195 1.435
R1389 VPB.n1427 VPB.n1424 1.435
R1390 VPB.n188 VPB.n181 1.402
R1391 VPB.n188 VPB.n182 1.402
R1392 VPB.n188 VPB.n186 1.402
R1393 VPB.n188 VPB.n187 1.402
R1394 VPB.n438 VPB.n435 1.076
R1395 VPB.n521 VPB.n518 1.076
R1396 VPB.n667 VPB.n664 1.076
R1397 VPB.n750 VPB.n747 1.076
R1398 VPB.n137 VPB.n134 1.076
R1399 VPB.n890 VPB.n887 1.076
R1400 VPB.n1036 VPB.n1033 1.076
R1401 VPB.n1119 VPB.n1116 1.076
R1402 VPB.n1265 VPB.n1262 1.076
R1403 VPB.n1348 VPB.n1345 1.076
R1404 VPB.n1494 VPB.n1491 1.076
R1405 VPB.n48 VPB.n45 1.076
R1406 VPB.n189 VPB.n188 0.735
R1407 VPB.n188 VPB.n178 0.735
R1408 VPB.n477 VPB.n474 0.717
R1409 VPB.n560 VPB.n557 0.717
R1410 VPB.n706 VPB.n703 0.717
R1411 VPB.n789 VPB.n786 0.717
R1412 VPB.n167 VPB.n166 0.717
R1413 VPB.n929 VPB.n926 0.717
R1414 VPB.n1075 VPB.n1072 0.717
R1415 VPB.n1158 VPB.n1155 0.717
R1416 VPB.n1304 VPB.n1301 0.717
R1417 VPB.n1387 VPB.n1384 0.717
R1418 VPB.n1533 VPB.n1530 0.717
R1419 VPB.n78 VPB.n77 0.717
R1420 VPB.n240 VPB.n239 0.387
R1421 VPB.n240 VPB.n235 0.387
R1422 VPB.n240 VPB.n230 0.387
R1423 VPB.n241 VPB.n240 0.387
R1424 VPB.n295 VPB.n294 0.387
R1425 VPB.n295 VPB.n290 0.387
R1426 VPB.n295 VPB.n285 0.387
R1427 VPB.n296 VPB.n295 0.387
R1428 VPB.n358 VPB.n357 0.387
R1429 VPB.n358 VPB.n353 0.387
R1430 VPB.n358 VPB.n348 0.387
R1431 VPB.n359 VPB.n358 0.387
R1432 VPB.n421 VPB.n420 0.387
R1433 VPB.n421 VPB.n416 0.387
R1434 VPB.n421 VPB.n411 0.387
R1435 VPB.n422 VPB.n421 0.387
R1436 VPB.n504 VPB.n503 0.387
R1437 VPB.n504 VPB.n499 0.387
R1438 VPB.n504 VPB.n494 0.387
R1439 VPB.n505 VPB.n504 0.387
R1440 VPB.n587 VPB.n586 0.387
R1441 VPB.n587 VPB.n582 0.387
R1442 VPB.n587 VPB.n577 0.387
R1443 VPB.n588 VPB.n587 0.387
R1444 VPB.n650 VPB.n649 0.387
R1445 VPB.n650 VPB.n645 0.387
R1446 VPB.n650 VPB.n640 0.387
R1447 VPB.n651 VPB.n650 0.387
R1448 VPB.n733 VPB.n732 0.387
R1449 VPB.n733 VPB.n728 0.387
R1450 VPB.n733 VPB.n723 0.387
R1451 VPB.n734 VPB.n733 0.387
R1452 VPB.n816 VPB.n815 0.387
R1453 VPB.n816 VPB.n811 0.387
R1454 VPB.n816 VPB.n806 0.387
R1455 VPB.n817 VPB.n816 0.387
R1456 VPB.n122 VPB.n121 0.387
R1457 VPB.n122 VPB.n117 0.387
R1458 VPB.n122 VPB.n112 0.387
R1459 VPB.n123 VPB.n122 0.387
R1460 VPB.n99 VPB.n98 0.387
R1461 VPB.n99 VPB.n94 0.387
R1462 VPB.n99 VPB.n89 0.387
R1463 VPB.n100 VPB.n99 0.387
R1464 VPB.n956 VPB.n955 0.387
R1465 VPB.n956 VPB.n951 0.387
R1466 VPB.n956 VPB.n946 0.387
R1467 VPB.n957 VPB.n956 0.387
R1468 VPB.n1019 VPB.n1018 0.387
R1469 VPB.n1019 VPB.n1014 0.387
R1470 VPB.n1019 VPB.n1009 0.387
R1471 VPB.n1020 VPB.n1019 0.387
R1472 VPB.n1102 VPB.n1101 0.387
R1473 VPB.n1102 VPB.n1097 0.387
R1474 VPB.n1102 VPB.n1092 0.387
R1475 VPB.n1103 VPB.n1102 0.387
R1476 VPB.n1185 VPB.n1184 0.387
R1477 VPB.n1185 VPB.n1180 0.387
R1478 VPB.n1185 VPB.n1175 0.387
R1479 VPB.n1186 VPB.n1185 0.387
R1480 VPB.n1248 VPB.n1247 0.387
R1481 VPB.n1248 VPB.n1243 0.387
R1482 VPB.n1248 VPB.n1238 0.387
R1483 VPB.n1249 VPB.n1248 0.387
R1484 VPB.n1331 VPB.n1330 0.387
R1485 VPB.n1331 VPB.n1326 0.387
R1486 VPB.n1331 VPB.n1321 0.387
R1487 VPB.n1332 VPB.n1331 0.387
R1488 VPB.n1414 VPB.n1413 0.387
R1489 VPB.n1414 VPB.n1409 0.387
R1490 VPB.n1414 VPB.n1404 0.387
R1491 VPB.n1415 VPB.n1414 0.387
R1492 VPB.n1477 VPB.n1476 0.387
R1493 VPB.n1477 VPB.n1472 0.387
R1494 VPB.n1477 VPB.n1467 0.387
R1495 VPB.n1478 VPB.n1477 0.387
R1496 VPB.n33 VPB.n32 0.387
R1497 VPB.n33 VPB.n28 0.387
R1498 VPB.n33 VPB.n23 0.387
R1499 VPB.n34 VPB.n33 0.387
R1500 VPB.n1562 VPB.n13 0.387
R1501 VPB.n1562 VPB.n9 0.387
R1502 VPB.n1562 VPB.n4 0.387
R1503 VPB.n1562 VPB.n1561 0.387
R1504 VPB.n249 VPB.n222 0.272
R1505 VPB.n304 VPB.n277 0.272
R1506 VPB.n367 VPB.n340 0.272
R1507 VPB.n430 VPB.n403 0.272
R1508 VPB.n513 VPB.n486 0.272
R1509 VPB.n596 VPB.n569 0.272
R1510 VPB.n659 VPB.n632 0.272
R1511 VPB.n742 VPB.n715 0.272
R1512 VPB.n825 VPB.n798 0.272
R1513 VPB.n862 VPB.n861 0.272
R1514 VPB.n965 VPB.n938 0.272
R1515 VPB.n1028 VPB.n1001 0.272
R1516 VPB.n1111 VPB.n1084 0.272
R1517 VPB.n1194 VPB.n1167 0.272
R1518 VPB.n1257 VPB.n1230 0.272
R1519 VPB.n1340 VPB.n1313 0.272
R1520 VPB.n1423 VPB.n1396 0.272
R1521 VPB.n1486 VPB.n1459 0.272
R1522 VPB.n1543 VPB.n1542 0.272
R1523 VPB.n882 VPB 0.204
R1524 VPB.n1554 VPB 0.198
R1525 VPB.n206 VPB.n205 0.136
R1526 VPB.n210 VPB.n206 0.136
R1527 VPB.n214 VPB.n210 0.136
R1528 VPB.n218 VPB.n214 0.136
R1529 VPB.n222 VPB.n218 0.136
R1530 VPB.n253 VPB.n249 0.136
R1531 VPB.n257 VPB.n253 0.136
R1532 VPB.n261 VPB.n257 0.136
R1533 VPB.n265 VPB.n261 0.136
R1534 VPB.n269 VPB.n265 0.136
R1535 VPB.n273 VPB.n269 0.136
R1536 VPB.n277 VPB.n273 0.136
R1537 VPB.n309 VPB.n304 0.136
R1538 VPB.n314 VPB.n309 0.136
R1539 VPB.n321 VPB.n314 0.136
R1540 VPB.n326 VPB.n321 0.136
R1541 VPB.n331 VPB.n326 0.136
R1542 VPB.n336 VPB.n331 0.136
R1543 VPB.n340 VPB.n336 0.136
R1544 VPB.n372 VPB.n367 0.136
R1545 VPB.n377 VPB.n372 0.136
R1546 VPB.n384 VPB.n377 0.136
R1547 VPB.n389 VPB.n384 0.136
R1548 VPB.n394 VPB.n389 0.136
R1549 VPB.n399 VPB.n394 0.136
R1550 VPB.n403 VPB.n399 0.136
R1551 VPB.n434 VPB.n430 0.136
R1552 VPB.n439 VPB.n434 0.136
R1553 VPB.n444 VPB.n439 0.136
R1554 VPB.n451 VPB.n444 0.136
R1555 VPB.n456 VPB.n451 0.136
R1556 VPB.n461 VPB.n456 0.136
R1557 VPB.n468 VPB.n461 0.136
R1558 VPB.n473 VPB.n468 0.136
R1559 VPB.n478 VPB.n473 0.136
R1560 VPB.n482 VPB.n478 0.136
R1561 VPB.n486 VPB.n482 0.136
R1562 VPB.n517 VPB.n513 0.136
R1563 VPB.n522 VPB.n517 0.136
R1564 VPB.n527 VPB.n522 0.136
R1565 VPB.n534 VPB.n527 0.136
R1566 VPB.n539 VPB.n534 0.136
R1567 VPB.n544 VPB.n539 0.136
R1568 VPB.n551 VPB.n544 0.136
R1569 VPB.n556 VPB.n551 0.136
R1570 VPB.n561 VPB.n556 0.136
R1571 VPB.n565 VPB.n561 0.136
R1572 VPB.n569 VPB.n565 0.136
R1573 VPB.n601 VPB.n596 0.136
R1574 VPB.n606 VPB.n601 0.136
R1575 VPB.n613 VPB.n606 0.136
R1576 VPB.n618 VPB.n613 0.136
R1577 VPB.n623 VPB.n618 0.136
R1578 VPB.n628 VPB.n623 0.136
R1579 VPB.n632 VPB.n628 0.136
R1580 VPB.n663 VPB.n659 0.136
R1581 VPB.n668 VPB.n663 0.136
R1582 VPB.n673 VPB.n668 0.136
R1583 VPB.n680 VPB.n673 0.136
R1584 VPB.n685 VPB.n680 0.136
R1585 VPB.n690 VPB.n685 0.136
R1586 VPB.n697 VPB.n690 0.136
R1587 VPB.n702 VPB.n697 0.136
R1588 VPB.n707 VPB.n702 0.136
R1589 VPB.n711 VPB.n707 0.136
R1590 VPB.n715 VPB.n711 0.136
R1591 VPB.n746 VPB.n742 0.136
R1592 VPB.n751 VPB.n746 0.136
R1593 VPB.n756 VPB.n751 0.136
R1594 VPB.n763 VPB.n756 0.136
R1595 VPB.n768 VPB.n763 0.136
R1596 VPB.n773 VPB.n768 0.136
R1597 VPB.n780 VPB.n773 0.136
R1598 VPB.n785 VPB.n780 0.136
R1599 VPB.n790 VPB.n785 0.136
R1600 VPB.n794 VPB.n790 0.136
R1601 VPB.n798 VPB.n794 0.136
R1602 VPB.n830 VPB.n825 0.136
R1603 VPB.n835 VPB.n830 0.136
R1604 VPB.n842 VPB.n835 0.136
R1605 VPB.n847 VPB.n842 0.136
R1606 VPB.n852 VPB.n847 0.136
R1607 VPB.n857 VPB.n852 0.136
R1608 VPB.n861 VPB.n857 0.136
R1609 VPB.n863 VPB.n862 0.136
R1610 VPB.n864 VPB.n863 0.136
R1611 VPB.n865 VPB.n864 0.136
R1612 VPB.n866 VPB.n865 0.136
R1613 VPB.n867 VPB.n866 0.136
R1614 VPB.n868 VPB.n867 0.136
R1615 VPB.n869 VPB.n868 0.136
R1616 VPB.n870 VPB.n869 0.136
R1617 VPB.n871 VPB.n870 0.136
R1618 VPB.n872 VPB.n871 0.136
R1619 VPB.n873 VPB.n872 0.136
R1620 VPB.n886 VPB.n882 0.136
R1621 VPB.n891 VPB.n886 0.136
R1622 VPB.n896 VPB.n891 0.136
R1623 VPB.n903 VPB.n896 0.136
R1624 VPB.n908 VPB.n903 0.136
R1625 VPB.n913 VPB.n908 0.136
R1626 VPB.n920 VPB.n913 0.136
R1627 VPB.n925 VPB.n920 0.136
R1628 VPB.n930 VPB.n925 0.136
R1629 VPB.n934 VPB.n930 0.136
R1630 VPB.n938 VPB.n934 0.136
R1631 VPB.n970 VPB.n965 0.136
R1632 VPB.n975 VPB.n970 0.136
R1633 VPB.n982 VPB.n975 0.136
R1634 VPB.n987 VPB.n982 0.136
R1635 VPB.n992 VPB.n987 0.136
R1636 VPB.n997 VPB.n992 0.136
R1637 VPB.n1001 VPB.n997 0.136
R1638 VPB.n1032 VPB.n1028 0.136
R1639 VPB.n1037 VPB.n1032 0.136
R1640 VPB.n1042 VPB.n1037 0.136
R1641 VPB.n1049 VPB.n1042 0.136
R1642 VPB.n1054 VPB.n1049 0.136
R1643 VPB.n1059 VPB.n1054 0.136
R1644 VPB.n1066 VPB.n1059 0.136
R1645 VPB.n1071 VPB.n1066 0.136
R1646 VPB.n1076 VPB.n1071 0.136
R1647 VPB.n1080 VPB.n1076 0.136
R1648 VPB.n1084 VPB.n1080 0.136
R1649 VPB.n1115 VPB.n1111 0.136
R1650 VPB.n1120 VPB.n1115 0.136
R1651 VPB.n1125 VPB.n1120 0.136
R1652 VPB.n1132 VPB.n1125 0.136
R1653 VPB.n1137 VPB.n1132 0.136
R1654 VPB.n1142 VPB.n1137 0.136
R1655 VPB.n1149 VPB.n1142 0.136
R1656 VPB.n1154 VPB.n1149 0.136
R1657 VPB.n1159 VPB.n1154 0.136
R1658 VPB.n1163 VPB.n1159 0.136
R1659 VPB.n1167 VPB.n1163 0.136
R1660 VPB.n1199 VPB.n1194 0.136
R1661 VPB.n1204 VPB.n1199 0.136
R1662 VPB.n1211 VPB.n1204 0.136
R1663 VPB.n1216 VPB.n1211 0.136
R1664 VPB.n1221 VPB.n1216 0.136
R1665 VPB.n1226 VPB.n1221 0.136
R1666 VPB.n1230 VPB.n1226 0.136
R1667 VPB.n1261 VPB.n1257 0.136
R1668 VPB.n1266 VPB.n1261 0.136
R1669 VPB.n1271 VPB.n1266 0.136
R1670 VPB.n1278 VPB.n1271 0.136
R1671 VPB.n1283 VPB.n1278 0.136
R1672 VPB.n1288 VPB.n1283 0.136
R1673 VPB.n1295 VPB.n1288 0.136
R1674 VPB.n1300 VPB.n1295 0.136
R1675 VPB.n1305 VPB.n1300 0.136
R1676 VPB.n1309 VPB.n1305 0.136
R1677 VPB.n1313 VPB.n1309 0.136
R1678 VPB.n1344 VPB.n1340 0.136
R1679 VPB.n1349 VPB.n1344 0.136
R1680 VPB.n1354 VPB.n1349 0.136
R1681 VPB.n1361 VPB.n1354 0.136
R1682 VPB.n1366 VPB.n1361 0.136
R1683 VPB.n1371 VPB.n1366 0.136
R1684 VPB.n1378 VPB.n1371 0.136
R1685 VPB.n1383 VPB.n1378 0.136
R1686 VPB.n1388 VPB.n1383 0.136
R1687 VPB.n1392 VPB.n1388 0.136
R1688 VPB.n1396 VPB.n1392 0.136
R1689 VPB.n1428 VPB.n1423 0.136
R1690 VPB.n1433 VPB.n1428 0.136
R1691 VPB.n1440 VPB.n1433 0.136
R1692 VPB.n1445 VPB.n1440 0.136
R1693 VPB.n1450 VPB.n1445 0.136
R1694 VPB.n1455 VPB.n1450 0.136
R1695 VPB.n1459 VPB.n1455 0.136
R1696 VPB.n1490 VPB.n1486 0.136
R1697 VPB.n1495 VPB.n1490 0.136
R1698 VPB.n1500 VPB.n1495 0.136
R1699 VPB.n1507 VPB.n1500 0.136
R1700 VPB.n1512 VPB.n1507 0.136
R1701 VPB.n1517 VPB.n1512 0.136
R1702 VPB.n1524 VPB.n1517 0.136
R1703 VPB.n1529 VPB.n1524 0.136
R1704 VPB.n1534 VPB.n1529 0.136
R1705 VPB.n1538 VPB.n1534 0.136
R1706 VPB.n1542 VPB.n1538 0.136
R1707 VPB.n1544 VPB.n1543 0.136
R1708 VPB.n1545 VPB.n1544 0.136
R1709 VPB.n1546 VPB.n1545 0.136
R1710 VPB.n1547 VPB.n1546 0.136
R1711 VPB.n1548 VPB.n1547 0.136
R1712 VPB.n1549 VPB.n1548 0.136
R1713 VPB.n1550 VPB.n1549 0.136
R1714 VPB.n1551 VPB.n1550 0.136
R1715 VPB.n1552 VPB.n1551 0.136
R1716 VPB.n1553 VPB.n1552 0.136
R1717 VPB.n1554 VPB.n1553 0.136
R1718 VPB.n873 VPB 0.068
R1719 a_14511_943.n2 a_14511_943.t6 475.572
R1720 a_14511_943.n1 a_14511_943.t7 469.145
R1721 a_14511_943.n6 a_14511_943.t8 454.685
R1722 a_14511_943.n6 a_14511_943.t13 428.979
R1723 a_14511_943.n2 a_14511_943.t10 384.527
R1724 a_14511_943.n1 a_14511_943.t9 384.527
R1725 a_14511_943.n3 a_14511_943.t12 277.772
R1726 a_14511_943.n5 a_14511_943.t11 251.219
R1727 a_14511_943.n7 a_14511_943.t5 248.006
R1728 a_14511_943.n13 a_14511_943.n12 220.639
R1729 a_14511_943.n4 a_14511_943.n3 156.851
R1730 a_14511_943.n14 a_14511_943.n13 135.994
R1731 a_14511_943.n7 a_14511_943.n6 81.941
R1732 a_14511_943.n8 a_14511_943.n7 78.947
R1733 a_14511_943.n8 a_14511_943.n5 77.859
R1734 a_14511_943.n15 a_14511_943.n14 76.001
R1735 a_14511_943.n13 a_14511_943.n8 76
R1736 a_14511_943.n3 a_14511_943.n2 67.889
R1737 a_14511_943.n4 a_14511_943.n1 66.88
R1738 a_14511_943.n12 a_14511_943.n11 30
R1739 a_14511_943.n5 a_14511_943.n4 26.552
R1740 a_14511_943.n10 a_14511_943.n9 24.383
R1741 a_14511_943.n12 a_14511_943.n10 23.684
R1742 a_14511_943.n0 a_14511_943.t1 14.282
R1743 a_14511_943.n0 a_14511_943.t0 14.282
R1744 a_14511_943.n15 a_14511_943.t2 14.282
R1745 a_14511_943.t3 a_14511_943.n15 14.282
R1746 a_14511_943.n14 a_14511_943.n0 12.85
R1747 a_9331_943.n9 a_9331_943.t19 512.525
R1748 a_9331_943.n4 a_9331_943.t32 512.525
R1749 a_9331_943.n21 a_9331_943.t5 480.392
R1750 a_9331_943.n5 a_9331_943.t34 477.179
R1751 a_9331_943.n38 a_9331_943.t33 454.685
R1752 a_9331_943.n35 a_9331_943.t28 454.685
R1753 a_9331_943.n38 a_9331_943.t21 428.979
R1754 a_9331_943.n35 a_9331_943.t26 428.979
R1755 a_9331_943.n5 a_9331_943.t30 406.485
R1756 a_9331_943.n21 a_9331_943.t7 403.272
R1757 a_9331_943.n9 a_9331_943.t27 371.139
R1758 a_9331_943.n4 a_9331_943.t23 371.139
R1759 a_9331_943.n6 a_9331_943.t31 346.633
R1760 a_9331_943.n10 a_9331_943.t20 271.162
R1761 a_9331_943.n22 a_9331_943.t29 266.974
R1762 a_9331_943.n8 a_9331_943.t24 260.547
R1763 a_9331_943.n39 a_9331_943.t25 221.453
R1764 a_9331_943.n36 a_9331_943.t22 221.453
R1765 a_9331_943.n33 a_9331_943.n32 196.598
R1766 a_9331_943.n19 a_9331_943.n18 194.086
R1767 a_9331_943.n43 a_9331_943.n41 194.086
R1768 a_9331_943.n33 a_9331_943.n28 180.846
R1769 a_9331_943.n10 a_9331_943.n9 172.76
R1770 a_9331_943.n19 a_9331_943.n14 162.547
R1771 a_9331_943.n41 a_9331_943.n3 162.547
R1772 a_9331_943.n7 a_9331_943.n6 154.675
R1773 a_9331_943.n39 a_9331_943.n38 108.494
R1774 a_9331_943.n36 a_9331_943.n35 108.494
R1775 a_9331_943.n22 a_9331_943.n21 108.494
R1776 a_9331_943.n7 a_9331_943.n4 89.615
R1777 a_9331_943.n11 a_9331_943.n8 85.204
R1778 a_9331_943.n8 a_9331_943.n7 79.658
R1779 a_9331_943.n27 a_9331_943.n26 79.232
R1780 a_9331_943.n40 a_9331_943.n39 78.947
R1781 a_9331_943.n14 a_9331_943.n13 76.002
R1782 a_9331_943.n3 a_9331_943.n2 76.002
R1783 a_9331_943.n11 a_9331_943.n10 76
R1784 a_9331_943.n20 a_9331_943.n19 76
R1785 a_9331_943.n23 a_9331_943.n22 76
R1786 a_9331_943.n34 a_9331_943.n33 76
R1787 a_9331_943.n37 a_9331_943.n36 76
R1788 a_9331_943.n41 a_9331_943.n40 76
R1789 a_9331_943.n28 a_9331_943.n27 63.152
R1790 a_9331_943.n44 a_9331_943.n0 55.263
R1791 a_9331_943.n32 a_9331_943.n31 30
R1792 a_9331_943.n18 a_9331_943.n17 30
R1793 a_9331_943.n43 a_9331_943.n42 30
R1794 a_9331_943.n6 a_9331_943.n5 29.194
R1795 a_9331_943.n30 a_9331_943.n29 24.383
R1796 a_9331_943.n16 a_9331_943.n15 24.383
R1797 a_9331_943.n32 a_9331_943.n30 23.684
R1798 a_9331_943.n18 a_9331_943.n16 23.684
R1799 a_9331_943.n44 a_9331_943.n43 23.684
R1800 a_9331_943.n28 a_9331_943.n24 16.08
R1801 a_9331_943.n27 a_9331_943.n25 16.08
R1802 a_9331_943.n24 a_9331_943.t11 14.282
R1803 a_9331_943.n24 a_9331_943.t10 14.282
R1804 a_9331_943.n25 a_9331_943.t17 14.282
R1805 a_9331_943.n25 a_9331_943.t18 14.282
R1806 a_9331_943.n26 a_9331_943.t1 14.282
R1807 a_9331_943.n26 a_9331_943.t4 14.282
R1808 a_9331_943.n12 a_9331_943.t15 14.282
R1809 a_9331_943.n12 a_9331_943.t14 14.282
R1810 a_9331_943.n13 a_9331_943.t6 14.282
R1811 a_9331_943.n13 a_9331_943.t8 14.282
R1812 a_9331_943.n1 a_9331_943.t3 14.282
R1813 a_9331_943.n1 a_9331_943.t2 14.282
R1814 a_9331_943.n2 a_9331_943.t9 14.282
R1815 a_9331_943.n2 a_9331_943.t13 14.282
R1816 a_9331_943.n14 a_9331_943.n12 12.85
R1817 a_9331_943.n3 a_9331_943.n1 12.85
R1818 a_9331_943.n37 a_9331_943.n34 4.035
R1819 a_9331_943.n40 a_9331_943.n37 2.947
R1820 a_9331_943.n20 a_9331_943.n11 1.315
R1821 a_9331_943.n34 a_9331_943.n23 1.315
R1822 a_9331_943.n23 a_9331_943.n20 1.043
R1823 a_5327_159.n10 a_5327_159.t10 512.525
R1824 a_5327_159.n8 a_5327_159.t15 472.359
R1825 a_5327_159.n6 a_5327_159.t12 472.359
R1826 a_5327_159.n8 a_5327_159.t11 384.527
R1827 a_5327_159.n6 a_5327_159.t8 384.527
R1828 a_5327_159.n10 a_5327_159.t13 371.139
R1829 a_5327_159.n11 a_5327_159.t14 324.268
R1830 a_5327_159.n9 a_5327_159.t9 277.772
R1831 a_5327_159.n7 a_5327_159.t7 277.772
R1832 a_5327_159.n16 a_5327_159.n14 249.704
R1833 a_5327_159.n14 a_5327_159.n5 127.74
R1834 a_5327_159.n11 a_5327_159.n10 119.654
R1835 a_5327_159.n12 a_5327_159.n11 83.572
R1836 a_5327_159.n13 a_5327_159.n7 81.396
R1837 a_5327_159.n4 a_5327_159.n3 79.232
R1838 a_5327_159.n12 a_5327_159.n9 76
R1839 a_5327_159.n14 a_5327_159.n13 76
R1840 a_5327_159.n9 a_5327_159.n8 67.001
R1841 a_5327_159.n7 a_5327_159.n6 67.001
R1842 a_5327_159.n5 a_5327_159.n4 63.152
R1843 a_5327_159.n16 a_5327_159.n15 30
R1844 a_5327_159.n17 a_5327_159.n0 24.383
R1845 a_5327_159.n17 a_5327_159.n16 23.684
R1846 a_5327_159.n5 a_5327_159.n1 16.08
R1847 a_5327_159.n4 a_5327_159.n2 16.08
R1848 a_5327_159.n1 a_5327_159.t2 14.282
R1849 a_5327_159.n1 a_5327_159.t3 14.282
R1850 a_5327_159.n2 a_5327_159.t5 14.282
R1851 a_5327_159.n2 a_5327_159.t6 14.282
R1852 a_5327_159.n3 a_5327_159.t1 14.282
R1853 a_5327_159.n3 a_5327_159.t0 14.282
R1854 a_5327_159.n13 a_5327_159.n12 4.035
R1855 a_9806_73.t0 a_9806_73.n1 93.333
R1856 a_9806_73.n4 a_9806_73.n2 55.07
R1857 a_9806_73.t0 a_9806_73.n0 8.137
R1858 a_9806_73.n4 a_9806_73.n3 4.619
R1859 a_9806_73.t0 a_9806_73.n4 0.071
R1860 a_6233_75.n4 a_6233_75.n3 19.724
R1861 a_6233_75.t0 a_6233_75.n5 11.595
R1862 a_6233_75.t0 a_6233_75.n4 9.207
R1863 a_6233_75.n2 a_6233_75.n0 8.543
R1864 a_6233_75.t0 a_6233_75.n2 3.034
R1865 a_6233_75.n2 a_6233_75.n1 0.443
R1866 a_6514_182.n12 a_6514_182.n5 96.467
R1867 a_6514_182.t0 a_6514_182.n1 46.91
R1868 a_6514_182.n9 a_6514_182.n7 34.805
R1869 a_6514_182.n9 a_6514_182.n8 32.622
R1870 a_6514_182.t0 a_6514_182.n12 32.417
R1871 a_6514_182.n5 a_6514_182.n4 22.349
R1872 a_6514_182.n11 a_6514_182.n9 19.017
R1873 a_6514_182.n1 a_6514_182.n0 17.006
R1874 a_6514_182.n5 a_6514_182.n3 8.443
R1875 a_6514_182.t0 a_6514_182.n2 8.137
R1876 a_6514_182.n7 a_6514_182.n6 7.5
R1877 a_6514_182.n11 a_6514_182.n10 7.5
R1878 a_6514_182.n12 a_6514_182.n11 1.435
R1879 a_5779_943.n5 a_5779_943.t10 480.392
R1880 a_5779_943.n7 a_5779_943.t7 454.685
R1881 a_5779_943.n7 a_5779_943.t9 428.979
R1882 a_5779_943.n5 a_5779_943.t8 403.272
R1883 a_5779_943.n6 a_5779_943.t12 266.974
R1884 a_5779_943.n8 a_5779_943.t11 221.453
R1885 a_5779_943.n12 a_5779_943.n10 203.12
R1886 a_5779_943.n10 a_5779_943.n4 180.846
R1887 a_5779_943.n8 a_5779_943.n7 108.494
R1888 a_5779_943.n6 a_5779_943.n5 108.494
R1889 a_5779_943.n9 a_5779_943.n8 80.035
R1890 a_5779_943.n3 a_5779_943.n2 79.232
R1891 a_5779_943.n9 a_5779_943.n6 77.315
R1892 a_5779_943.n10 a_5779_943.n9 76
R1893 a_5779_943.n4 a_5779_943.n3 63.152
R1894 a_5779_943.n4 a_5779_943.n0 16.08
R1895 a_5779_943.n3 a_5779_943.n1 16.08
R1896 a_5779_943.n12 a_5779_943.n11 15.218
R1897 a_5779_943.n0 a_5779_943.t3 14.282
R1898 a_5779_943.n0 a_5779_943.t2 14.282
R1899 a_5779_943.n1 a_5779_943.t6 14.282
R1900 a_5779_943.n1 a_5779_943.t5 14.282
R1901 a_5779_943.n2 a_5779_943.t0 14.282
R1902 a_5779_943.n2 a_5779_943.t1 14.282
R1903 a_5779_943.n13 a_5779_943.n12 12.014
R1904 a_5457_1004.n8 a_5457_1004.t8 512.525
R1905 a_5457_1004.n6 a_5457_1004.t7 512.525
R1906 a_5457_1004.n8 a_5457_1004.t10 371.139
R1907 a_5457_1004.n6 a_5457_1004.t9 371.139
R1908 a_5457_1004.n9 a_5457_1004.t12 297.715
R1909 a_5457_1004.n7 a_5457_1004.t11 297.715
R1910 a_5457_1004.n13 a_5457_1004.n11 223.151
R1911 a_5457_1004.n11 a_5457_1004.n5 154.293
R1912 a_5457_1004.n9 a_5457_1004.n8 146.207
R1913 a_5457_1004.n7 a_5457_1004.n6 146.207
R1914 a_5457_1004.n10 a_5457_1004.n7 85.476
R1915 a_5457_1004.n4 a_5457_1004.n3 79.232
R1916 a_5457_1004.n11 a_5457_1004.n10 77.315
R1917 a_5457_1004.n10 a_5457_1004.n9 76
R1918 a_5457_1004.n5 a_5457_1004.n4 63.152
R1919 a_5457_1004.n13 a_5457_1004.n12 30
R1920 a_5457_1004.n14 a_5457_1004.n0 24.383
R1921 a_5457_1004.n14 a_5457_1004.n13 23.684
R1922 a_5457_1004.n5 a_5457_1004.n1 16.08
R1923 a_5457_1004.n4 a_5457_1004.n2 16.08
R1924 a_5457_1004.n1 a_5457_1004.t2 14.282
R1925 a_5457_1004.n1 a_5457_1004.t3 14.282
R1926 a_5457_1004.n2 a_5457_1004.t6 14.282
R1927 a_5457_1004.n2 a_5457_1004.t5 14.282
R1928 a_5457_1004.n3 a_5457_1004.t1 14.282
R1929 a_5457_1004.n3 a_5457_1004.t0 14.282
R1930 a_147_159.n17 a_147_159.t14 512.525
R1931 a_147_159.n2 a_147_159.t23 480.392
R1932 a_147_159.n15 a_147_159.t17 472.359
R1933 a_147_159.n0 a_147_159.t25 472.359
R1934 a_147_159.n2 a_147_159.t16 403.272
R1935 a_147_159.n15 a_147_159.t22 384.527
R1936 a_147_159.n0 a_147_159.t18 384.527
R1937 a_147_159.n17 a_147_159.t19 371.139
R1938 a_147_159.n18 a_147_159.t24 324.268
R1939 a_147_159.n3 a_147_159.t15 320.08
R1940 a_147_159.n16 a_147_159.t21 277.772
R1941 a_147_159.n1 a_147_159.t20 277.772
R1942 a_147_159.n13 a_147_159.n12 265.227
R1943 a_147_159.n25 a_147_159.n24 249.704
R1944 a_147_159.n13 a_147_159.n9 127.74
R1945 a_147_159.n29 a_147_159.n25 127.74
R1946 a_147_159.n18 a_147_159.n17 119.654
R1947 a_147_159.n19 a_147_159.n18 83.572
R1948 a_147_159.n8 a_147_159.n7 79.232
R1949 a_147_159.n28 a_147_159.n27 79.232
R1950 a_147_159.n4 a_147_159.n1 76.499
R1951 a_147_159.n19 a_147_159.n16 76
R1952 a_147_159.n4 a_147_159.n3 76
R1953 a_147_159.n14 a_147_159.n13 76
R1954 a_147_159.n25 a_147_159.n20 76
R1955 a_147_159.n16 a_147_159.n15 67.001
R1956 a_147_159.n1 a_147_159.n0 67.001
R1957 a_147_159.n9 a_147_159.n8 63.152
R1958 a_147_159.n29 a_147_159.n28 63.152
R1959 a_147_159.n3 a_147_159.n2 55.388
R1960 a_147_159.n24 a_147_159.n23 30
R1961 a_147_159.n22 a_147_159.n21 24.383
R1962 a_147_159.n24 a_147_159.n22 23.684
R1963 a_147_159.n12 a_147_159.n11 22.578
R1964 a_147_159.n28 a_147_159.n26 16.08
R1965 a_147_159.n9 a_147_159.n5 16.08
R1966 a_147_159.n8 a_147_159.n6 16.08
R1967 a_147_159.n30 a_147_159.n29 16.078
R1968 a_147_159.n26 a_147_159.t12 14.282
R1969 a_147_159.n26 a_147_159.t13 14.282
R1970 a_147_159.n27 a_147_159.t3 14.282
R1971 a_147_159.n27 a_147_159.t10 14.282
R1972 a_147_159.n5 a_147_159.t1 14.282
R1973 a_147_159.n5 a_147_159.t9 14.282
R1974 a_147_159.n6 a_147_159.t6 14.282
R1975 a_147_159.n6 a_147_159.t5 14.282
R1976 a_147_159.n7 a_147_159.t11 14.282
R1977 a_147_159.n7 a_147_159.t2 14.282
R1978 a_147_159.n30 a_147_159.t4 14.282
R1979 a_147_159.t7 a_147_159.n30 14.282
R1980 a_147_159.n12 a_147_159.n10 8.58
R1981 a_147_159.n20 a_147_159.n19 4.035
R1982 a_147_159.n20 a_147_159.n14 3.491
R1983 a_147_159.n14 a_147_159.n4 1.315
R1984 a_277_1004.n7 a_277_1004.t10 512.525
R1985 a_277_1004.n5 a_277_1004.t8 512.525
R1986 a_277_1004.n7 a_277_1004.t12 371.139
R1987 a_277_1004.n5 a_277_1004.t11 371.139
R1988 a_277_1004.n8 a_277_1004.t9 297.715
R1989 a_277_1004.n6 a_277_1004.t7 297.715
R1990 a_277_1004.n12 a_277_1004.n10 229.673
R1991 a_277_1004.n10 a_277_1004.n4 154.293
R1992 a_277_1004.n8 a_277_1004.n7 146.207
R1993 a_277_1004.n6 a_277_1004.n5 146.207
R1994 a_277_1004.n9 a_277_1004.n6 85.476
R1995 a_277_1004.n3 a_277_1004.n2 79.232
R1996 a_277_1004.n10 a_277_1004.n9 77.315
R1997 a_277_1004.n9 a_277_1004.n8 76
R1998 a_277_1004.n4 a_277_1004.n3 63.152
R1999 a_277_1004.n4 a_277_1004.n0 16.08
R2000 a_277_1004.n3 a_277_1004.n1 16.08
R2001 a_277_1004.n12 a_277_1004.n11 15.218
R2002 a_277_1004.n0 a_277_1004.t2 14.282
R2003 a_277_1004.n0 a_277_1004.t0 14.282
R2004 a_277_1004.n1 a_277_1004.t6 14.282
R2005 a_277_1004.n1 a_277_1004.t5 14.282
R2006 a_277_1004.n2 a_277_1004.t4 14.282
R2007 a_277_1004.n2 a_277_1004.t3 14.282
R2008 a_277_1004.n13 a_277_1004.n12 12.014
R2009 a_4151_943.n2 a_4151_943.t13 512.525
R2010 a_4151_943.n1 a_4151_943.t10 512.525
R2011 a_4151_943.n6 a_4151_943.t7 454.685
R2012 a_4151_943.n6 a_4151_943.t11 428.979
R2013 a_4151_943.n2 a_4151_943.t8 371.139
R2014 a_4151_943.n1 a_4151_943.t5 371.139
R2015 a_4151_943.n3 a_4151_943.n2 258.98
R2016 a_4151_943.n5 a_4151_943.n1 195.827
R2017 a_4151_943.n14 a_4151_943.n13 189.099
R2018 a_4151_943.n7 a_4151_943.t12 183.653
R2019 a_4151_943.n3 a_4151_943.t9 176.995
R2020 a_4151_943.n4 a_4151_943.t6 170.569
R2021 a_4151_943.n13 a_4151_943.n12 167.533
R2022 a_4151_943.n4 a_4151_943.n3 153.043
R2023 a_4151_943.n7 a_4151_943.n6 135.047
R2024 a_4151_943.n8 a_4151_943.n5 118.94
R2025 a_4151_943.n8 a_4151_943.n7 78.947
R2026 a_4151_943.n15 a_4151_943.n14 76.001
R2027 a_4151_943.n13 a_4151_943.n8 76
R2028 a_4151_943.n5 a_4151_943.n4 63.152
R2029 a_4151_943.n12 a_4151_943.n11 30
R2030 a_4151_943.n10 a_4151_943.n9 24.383
R2031 a_4151_943.n12 a_4151_943.n10 23.684
R2032 a_4151_943.n0 a_4151_943.t0 14.282
R2033 a_4151_943.n0 a_4151_943.t2 14.282
R2034 a_4151_943.n15 a_4151_943.t1 14.282
R2035 a_4151_943.t3 a_4151_943.n15 14.282
R2036 a_4151_943.n14 a_4151_943.n0 12.85
R2037 a_16421_1005.n4 a_16421_1005.n3 196.002
R2038 a_16421_1005.n2 a_16421_1005.t6 89.553
R2039 a_16421_1005.n5 a_16421_1005.n4 75.27
R2040 a_16421_1005.n3 a_16421_1005.n2 75.214
R2041 a_16421_1005.n4 a_16421_1005.n0 36.52
R2042 a_16421_1005.n3 a_16421_1005.t3 14.338
R2043 a_16421_1005.n0 a_16421_1005.t2 14.282
R2044 a_16421_1005.n0 a_16421_1005.t5 14.282
R2045 a_16421_1005.n1 a_16421_1005.t7 14.282
R2046 a_16421_1005.n1 a_16421_1005.t4 14.282
R2047 a_16421_1005.n5 a_16421_1005.t1 14.282
R2048 a_16421_1005.t0 a_16421_1005.n5 14.282
R2049 a_16421_1005.n2 a_16421_1005.n1 12.119
R2050 a_15757_1005.n4 a_15757_1005.n3 195.987
R2051 a_15757_1005.n2 a_15757_1005.t5 89.553
R2052 a_15757_1005.n5 a_15757_1005.n4 75.27
R2053 a_15757_1005.n3 a_15757_1005.n2 75.214
R2054 a_15757_1005.n4 a_15757_1005.n0 36.519
R2055 a_15757_1005.n3 a_15757_1005.t3 14.338
R2056 a_15757_1005.n0 a_15757_1005.t7 14.282
R2057 a_15757_1005.n0 a_15757_1005.t6 14.282
R2058 a_15757_1005.n1 a_15757_1005.t4 14.282
R2059 a_15757_1005.n1 a_15757_1005.t2 14.282
R2060 a_15757_1005.n5 a_15757_1005.t0 14.282
R2061 a_15757_1005.t1 a_15757_1005.n5 14.282
R2062 a_15757_1005.n2 a_15757_1005.n1 12.119
R2063 a_10637_1004.n8 a_10637_1004.t12 512.525
R2064 a_10637_1004.n6 a_10637_1004.t11 512.525
R2065 a_10637_1004.n8 a_10637_1004.t8 371.139
R2066 a_10637_1004.n6 a_10637_1004.t7 371.139
R2067 a_10637_1004.n9 a_10637_1004.t10 297.715
R2068 a_10637_1004.n7 a_10637_1004.t9 297.715
R2069 a_10637_1004.n13 a_10637_1004.n11 223.151
R2070 a_10637_1004.n11 a_10637_1004.n5 154.293
R2071 a_10637_1004.n9 a_10637_1004.n8 146.207
R2072 a_10637_1004.n7 a_10637_1004.n6 146.207
R2073 a_10637_1004.n10 a_10637_1004.n7 85.476
R2074 a_10637_1004.n4 a_10637_1004.n3 79.232
R2075 a_10637_1004.n11 a_10637_1004.n10 77.315
R2076 a_10637_1004.n10 a_10637_1004.n9 76
R2077 a_10637_1004.n5 a_10637_1004.n4 63.152
R2078 a_10637_1004.n13 a_10637_1004.n12 30
R2079 a_10637_1004.n14 a_10637_1004.n0 24.383
R2080 a_10637_1004.n14 a_10637_1004.n13 23.684
R2081 a_10637_1004.n5 a_10637_1004.n1 16.08
R2082 a_10637_1004.n4 a_10637_1004.n2 16.08
R2083 a_10637_1004.n1 a_10637_1004.t1 14.282
R2084 a_10637_1004.n1 a_10637_1004.t0 14.282
R2085 a_10637_1004.n2 a_10637_1004.t6 14.282
R2086 a_10637_1004.n2 a_10637_1004.t5 14.282
R2087 a_10637_1004.n3 a_10637_1004.t4 14.282
R2088 a_10637_1004.n3 a_10637_1004.t3 14.282
R2089 a_14284_182.n10 a_14284_182.n8 82.852
R2090 a_14284_182.n7 a_14284_182.n6 32.833
R2091 a_14284_182.n8 a_14284_182.t1 32.416
R2092 a_14284_182.n10 a_14284_182.n9 27.2
R2093 a_14284_182.n11 a_14284_182.n0 23.498
R2094 a_14284_182.n3 a_14284_182.n2 23.284
R2095 a_14284_182.n11 a_14284_182.n10 22.4
R2096 a_14284_182.n7 a_14284_182.n4 19.017
R2097 a_14284_182.n6 a_14284_182.n5 13.494
R2098 a_14284_182.t1 a_14284_182.n1 7.04
R2099 a_14284_182.t1 a_14284_182.n3 5.727
R2100 a_14284_182.n8 a_14284_182.n7 1.435
R2101 a_13041_75.t0 a_13041_75.n3 117.777
R2102 a_13041_75.n6 a_13041_75.n5 45.444
R2103 a_13041_75.t0 a_13041_75.n6 21.213
R2104 a_13041_75.t0 a_13041_75.n4 11.595
R2105 a_13041_75.n2 a_13041_75.n0 8.543
R2106 a_13041_75.t0 a_13041_75.n2 3.034
R2107 a_13041_75.n2 a_13041_75.n1 0.443
R2108 VNB VNB.n1399 300.778
R2109 VNB.n205 VNB.n204 199.897
R2110 VNB.n264 VNB.n263 199.897
R2111 VNB.n323 VNB.n322 199.897
R2112 VNB.n382 VNB.n381 199.897
R2113 VNB.n457 VNB.n456 199.897
R2114 VNB.n525 VNB.n524 199.897
R2115 VNB.n584 VNB.n583 199.897
R2116 VNB.n659 VNB.n658 199.897
R2117 VNB.n734 VNB.n733 199.897
R2118 VNB.n94 VNB.n93 199.897
R2119 VNB.n74 VNB.n73 199.897
R2120 VNB.n853 VNB.n852 199.897
R2121 VNB.n912 VNB.n911 199.897
R2122 VNB.n980 VNB.n979 199.897
R2123 VNB.n1055 VNB.n1054 199.897
R2124 VNB.n1114 VNB.n1113 199.897
R2125 VNB.n1189 VNB.n1188 199.897
R2126 VNB.n1257 VNB.n1256 199.897
R2127 VNB.n1309 VNB.n1308 199.897
R2128 VNB.n18 VNB.n17 199.897
R2129 VNB.n214 VNB.n212 154.509
R2130 VNB.n332 VNB.n330 154.509
R2131 VNB.n273 VNB.n271 154.509
R2132 VNB.n466 VNB.n464 154.509
R2133 VNB.n391 VNB.n389 154.509
R2134 VNB.n593 VNB.n591 154.509
R2135 VNB.n534 VNB.n532 154.509
R2136 VNB.n743 VNB.n741 154.509
R2137 VNB.n668 VNB.n666 154.509
R2138 VNB.n794 VNB.n792 154.509
R2139 VNB.n103 VNB.n101 154.509
R2140 VNB.n921 VNB.n919 154.509
R2141 VNB.n862 VNB.n860 154.509
R2142 VNB.n1064 VNB.n1062 154.509
R2143 VNB.n989 VNB.n987 154.509
R2144 VNB.n1198 VNB.n1196 154.509
R2145 VNB.n1123 VNB.n1121 154.509
R2146 VNB.n1318 VNB.n1316 154.509
R2147 VNB.n1266 VNB.n1264 154.509
R2148 VNB.n27 VNB.n25 154.509
R2149 VNB.n423 VNB.n422 147.75
R2150 VNB.n625 VNB.n624 147.75
R2151 VNB.n700 VNB.n699 147.75
R2152 VNB.n127 VNB.n126 147.75
R2153 VNB.n1021 VNB.n1020 147.75
R2154 VNB.n1155 VNB.n1154 147.75
R2155 VNB.n1350 VNB.n1349 147.75
R2156 VNB.n51 VNB.n50 147.75
R2157 VNB.n171 VNB.n170 121.366
R2158 VNB.n230 VNB.n229 121.366
R2159 VNB.n289 VNB.n288 121.366
R2160 VNB.n348 VNB.n347 121.366
R2161 VNB.n435 VNB.n432 121.366
R2162 VNB.n550 VNB.n549 121.366
R2163 VNB.n637 VNB.n634 121.366
R2164 VNB.n712 VNB.n709 121.366
R2165 VNB.n132 VNB.n130 121.366
R2166 VNB.n878 VNB.n877 121.366
R2167 VNB.n1033 VNB.n1030 121.366
R2168 VNB.n1080 VNB.n1079 121.366
R2169 VNB.n1167 VNB.n1164 121.366
R2170 VNB.n1362 VNB.n1359 121.366
R2171 VNB.n56 VNB.n54 121.366
R2172 VNB.n502 VNB.n501 85.559
R2173 VNB.n830 VNB.n829 85.559
R2174 VNB.n957 VNB.n956 85.559
R2175 VNB.n1234 VNB.n1233 85.559
R2176 VNB.n763 VNB.n762 84.842
R2177 VNB.n1286 VNB.n1285 84.842
R2178 VNB.n1386 VNB.n1385 76
R2179 VNB.n1373 VNB.n1372 76
R2180 VNB.n1369 VNB.n1368 76
R2181 VNB.n1365 VNB.n1364 76
R2182 VNB.n1353 VNB.n1352 76
R2183 VNB.n1348 VNB.n1347 76
R2184 VNB.n1344 VNB.n1343 76
R2185 VNB.n1340 VNB.n1339 76
R2186 VNB.n1336 VNB.n1335 76
R2187 VNB.n1332 VNB.n1331 76
R2188 VNB.n1328 VNB.n1327 76
R2189 VNB.n1324 VNB.n1323 76
R2190 VNB.n1320 VNB.n1319 76
R2191 VNB.n1298 VNB.n1297 76
R2192 VNB.n1294 VNB.n1293 76
R2193 VNB.n1290 VNB.n1289 76
R2194 VNB.n1284 VNB.n1283 76
R2195 VNB.n1280 VNB.n1279 76
R2196 VNB.n1276 VNB.n1275 76
R2197 VNB.n1272 VNB.n1271 76
R2198 VNB.n1268 VNB.n1267 76
R2199 VNB.n1246 VNB.n1245 76
R2200 VNB.n1242 VNB.n1241 76
R2201 VNB.n1238 VNB.n1237 76
R2202 VNB.n1232 VNB.n1231 76
R2203 VNB.n1228 VNB.n1227 76
R2204 VNB.n1224 VNB.n1223 76
R2205 VNB.n1220 VNB.n1219 76
R2206 VNB.n1216 VNB.n1215 76
R2207 VNB.n1212 VNB.n1211 76
R2208 VNB.n1208 VNB.n1207 76
R2209 VNB.n1204 VNB.n1203 76
R2210 VNB.n1200 VNB.n1199 76
R2211 VNB.n1178 VNB.n1177 76
R2212 VNB.n1174 VNB.n1173 76
R2213 VNB.n1170 VNB.n1169 76
R2214 VNB.n1158 VNB.n1157 76
R2215 VNB.n1153 VNB.n1152 76
R2216 VNB.n1149 VNB.n1148 76
R2217 VNB.n1145 VNB.n1144 76
R2218 VNB.n1141 VNB.n1140 76
R2219 VNB.n1137 VNB.n1136 76
R2220 VNB.n1133 VNB.n1132 76
R2221 VNB.n1129 VNB.n1128 76
R2222 VNB.n1125 VNB.n1124 76
R2223 VNB.n1103 VNB.n1102 76
R2224 VNB.n1099 VNB.n1098 76
R2225 VNB.n1095 VNB.n1094 76
R2226 VNB.n1084 VNB.n1083 76
R2227 VNB.n1078 VNB.n1077 76
R2228 VNB.n1074 VNB.n1073 76
R2229 VNB.n1070 VNB.n1069 76
R2230 VNB.n1066 VNB.n1065 76
R2231 VNB.n1044 VNB.n1043 76
R2232 VNB.n1040 VNB.n1039 76
R2233 VNB.n1036 VNB.n1035 76
R2234 VNB.n1024 VNB.n1023 76
R2235 VNB.n1019 VNB.n1018 76
R2236 VNB.n1015 VNB.n1014 76
R2237 VNB.n1011 VNB.n1010 76
R2238 VNB.n1007 VNB.n1006 76
R2239 VNB.n1003 VNB.n1002 76
R2240 VNB.n999 VNB.n998 76
R2241 VNB.n995 VNB.n994 76
R2242 VNB.n991 VNB.n990 76
R2243 VNB.n969 VNB.n968 76
R2244 VNB.n965 VNB.n964 76
R2245 VNB.n961 VNB.n960 76
R2246 VNB.n955 VNB.n954 76
R2247 VNB.n951 VNB.n950 76
R2248 VNB.n947 VNB.n946 76
R2249 VNB.n943 VNB.n942 76
R2250 VNB.n939 VNB.n938 76
R2251 VNB.n935 VNB.n934 76
R2252 VNB.n931 VNB.n930 76
R2253 VNB.n927 VNB.n926 76
R2254 VNB.n923 VNB.n922 76
R2255 VNB.n901 VNB.n900 76
R2256 VNB.n897 VNB.n896 76
R2257 VNB.n893 VNB.n892 76
R2258 VNB.n882 VNB.n881 76
R2259 VNB.n876 VNB.n875 76
R2260 VNB.n872 VNB.n871 76
R2261 VNB.n868 VNB.n867 76
R2262 VNB.n864 VNB.n863 76
R2263 VNB.n842 VNB.n841 76
R2264 VNB.n838 VNB.n837 76
R2265 VNB.n834 VNB.n833 76
R2266 VNB.n828 VNB.n827 76
R2267 VNB.n824 VNB.n823 76
R2268 VNB.n820 VNB.n819 76
R2269 VNB.n816 VNB.n815 76
R2270 VNB.n812 VNB.n811 76
R2271 VNB.n808 VNB.n807 76
R2272 VNB.n804 VNB.n803 76
R2273 VNB.n800 VNB.n799 76
R2274 VNB.n796 VNB.n795 76
R2275 VNB.n790 VNB.n787 76
R2276 VNB.n775 VNB.n774 76
R2277 VNB.n771 VNB.n770 76
R2278 VNB.n767 VNB.n766 76
R2279 VNB.n761 VNB.n760 76
R2280 VNB.n757 VNB.n756 76
R2281 VNB.n753 VNB.n752 76
R2282 VNB.n749 VNB.n748 76
R2283 VNB.n745 VNB.n744 76
R2284 VNB.n723 VNB.n722 76
R2285 VNB.n719 VNB.n718 76
R2286 VNB.n715 VNB.n714 76
R2287 VNB.n703 VNB.n702 76
R2288 VNB.n698 VNB.n697 76
R2289 VNB.n694 VNB.n693 76
R2290 VNB.n690 VNB.n689 76
R2291 VNB.n686 VNB.n685 76
R2292 VNB.n682 VNB.n681 76
R2293 VNB.n678 VNB.n677 76
R2294 VNB.n674 VNB.n673 76
R2295 VNB.n670 VNB.n669 76
R2296 VNB.n648 VNB.n647 76
R2297 VNB.n644 VNB.n643 76
R2298 VNB.n640 VNB.n639 76
R2299 VNB.n628 VNB.n627 76
R2300 VNB.n623 VNB.n622 76
R2301 VNB.n619 VNB.n618 76
R2302 VNB.n615 VNB.n614 76
R2303 VNB.n611 VNB.n610 76
R2304 VNB.n607 VNB.n606 76
R2305 VNB.n603 VNB.n602 76
R2306 VNB.n599 VNB.n598 76
R2307 VNB.n595 VNB.n594 76
R2308 VNB.n573 VNB.n572 76
R2309 VNB.n569 VNB.n568 76
R2310 VNB.n565 VNB.n564 76
R2311 VNB.n554 VNB.n553 76
R2312 VNB.n548 VNB.n547 76
R2313 VNB.n544 VNB.n543 76
R2314 VNB.n540 VNB.n539 76
R2315 VNB.n536 VNB.n535 76
R2316 VNB.n514 VNB.n513 76
R2317 VNB.n510 VNB.n509 76
R2318 VNB.n506 VNB.n505 76
R2319 VNB.n500 VNB.n499 76
R2320 VNB.n496 VNB.n495 76
R2321 VNB.n492 VNB.n491 76
R2322 VNB.n488 VNB.n487 76
R2323 VNB.n484 VNB.n483 76
R2324 VNB.n480 VNB.n479 76
R2325 VNB.n476 VNB.n475 76
R2326 VNB.n472 VNB.n471 76
R2327 VNB.n468 VNB.n467 76
R2328 VNB.n446 VNB.n445 76
R2329 VNB.n442 VNB.n441 76
R2330 VNB.n438 VNB.n437 76
R2331 VNB.n426 VNB.n425 76
R2332 VNB.n421 VNB.n420 76
R2333 VNB.n417 VNB.n416 76
R2334 VNB.n413 VNB.n412 76
R2335 VNB.n409 VNB.n408 76
R2336 VNB.n405 VNB.n404 76
R2337 VNB.n401 VNB.n400 76
R2338 VNB.n397 VNB.n396 76
R2339 VNB.n393 VNB.n392 76
R2340 VNB.n371 VNB.n370 76
R2341 VNB.n367 VNB.n366 76
R2342 VNB.n363 VNB.n362 76
R2343 VNB.n352 VNB.n351 76
R2344 VNB.n346 VNB.n345 76
R2345 VNB.n342 VNB.n341 76
R2346 VNB.n338 VNB.n337 76
R2347 VNB.n334 VNB.n333 76
R2348 VNB.n312 VNB.n311 76
R2349 VNB.n308 VNB.n307 76
R2350 VNB.n304 VNB.n303 76
R2351 VNB.n293 VNB.n292 76
R2352 VNB.n287 VNB.n286 76
R2353 VNB.n283 VNB.n282 76
R2354 VNB.n279 VNB.n278 76
R2355 VNB.n275 VNB.n274 76
R2356 VNB.n253 VNB.n252 76
R2357 VNB.n249 VNB.n248 76
R2358 VNB.n245 VNB.n244 76
R2359 VNB.n234 VNB.n233 76
R2360 VNB.n228 VNB.n227 76
R2361 VNB.n224 VNB.n223 76
R2362 VNB.n220 VNB.n219 76
R2363 VNB.n216 VNB.n215 76
R2364 VNB.n194 VNB.n193 76
R2365 VNB.n190 VNB.n189 76
R2366 VNB.n186 VNB.n185 76
R2367 VNB.n175 VNB.n174 76
R2368 VNB.n137 VNB.n136 73.875
R2369 VNB.n61 VNB.n60 73.875
R2370 VNB.n431 VNB.n430 64.552
R2371 VNB.n633 VNB.n632 64.552
R2372 VNB.n708 VNB.n707 64.552
R2373 VNB.n135 VNB.n83 64.552
R2374 VNB.n1029 VNB.n1028 64.552
R2375 VNB.n1163 VNB.n1162 64.552
R2376 VNB.n1358 VNB.n1357 64.552
R2377 VNB.n59 VNB.n7 64.552
R2378 VNB.n180 VNB.n179 63.835
R2379 VNB.n239 VNB.n238 63.835
R2380 VNB.n298 VNB.n297 63.835
R2381 VNB.n357 VNB.n356 63.835
R2382 VNB.n559 VNB.n558 63.835
R2383 VNB.n887 VNB.n886 63.835
R2384 VNB.n1089 VNB.n1088 63.835
R2385 VNB.n504 VNB.n503 41.971
R2386 VNB.n832 VNB.n831 41.971
R2387 VNB.n959 VNB.n958 41.971
R2388 VNB.n1236 VNB.n1235 41.971
R2389 VNB.n172 VNB.n171 36.937
R2390 VNB.n231 VNB.n230 36.937
R2391 VNB.n290 VNB.n289 36.937
R2392 VNB.n349 VNB.n348 36.937
R2393 VNB.n435 VNB.n434 36.937
R2394 VNB.n551 VNB.n550 36.937
R2395 VNB.n637 VNB.n636 36.937
R2396 VNB.n712 VNB.n711 36.937
R2397 VNB.n132 VNB.n131 36.937
R2398 VNB.n879 VNB.n878 36.937
R2399 VNB.n1033 VNB.n1032 36.937
R2400 VNB.n1081 VNB.n1080 36.937
R2401 VNB.n1167 VNB.n1166 36.937
R2402 VNB.n1362 VNB.n1361 36.937
R2403 VNB.n56 VNB.n55 36.937
R2404 VNB.n765 VNB.n764 36.678
R2405 VNB.n1288 VNB.n1287 36.678
R2406 VNB.n168 VNB.n167 35.118
R2407 VNB.n434 VNB.n433 29.844
R2408 VNB.n636 VNB.n635 29.844
R2409 VNB.n711 VNB.n710 29.844
R2410 VNB.n1032 VNB.n1031 29.844
R2411 VNB.n1166 VNB.n1165 29.844
R2412 VNB.n1361 VNB.n1360 29.844
R2413 VNB.n179 VNB.n178 28.421
R2414 VNB.n238 VNB.n237 28.421
R2415 VNB.n297 VNB.n296 28.421
R2416 VNB.n356 VNB.n355 28.421
R2417 VNB.n430 VNB.n429 28.421
R2418 VNB.n558 VNB.n557 28.421
R2419 VNB.n632 VNB.n631 28.421
R2420 VNB.n707 VNB.n706 28.421
R2421 VNB.n83 VNB.n82 28.421
R2422 VNB.n886 VNB.n885 28.421
R2423 VNB.n1028 VNB.n1027 28.421
R2424 VNB.n1088 VNB.n1087 28.421
R2425 VNB.n1162 VNB.n1161 28.421
R2426 VNB.n1357 VNB.n1356 28.421
R2427 VNB.n7 VNB.n6 28.421
R2428 VNB.n183 VNB.n182 27.855
R2429 VNB.n242 VNB.n241 27.855
R2430 VNB.n301 VNB.n300 27.855
R2431 VNB.n360 VNB.n359 27.855
R2432 VNB.n562 VNB.n561 27.855
R2433 VNB.n890 VNB.n889 27.855
R2434 VNB.n1092 VNB.n1091 27.855
R2435 VNB.n179 VNB.n177 25.263
R2436 VNB.n238 VNB.n236 25.263
R2437 VNB.n297 VNB.n295 25.263
R2438 VNB.n356 VNB.n354 25.263
R2439 VNB.n430 VNB.n428 25.263
R2440 VNB.n558 VNB.n556 25.263
R2441 VNB.n632 VNB.n630 25.263
R2442 VNB.n707 VNB.n705 25.263
R2443 VNB.n83 VNB.n81 25.263
R2444 VNB.n886 VNB.n884 25.263
R2445 VNB.n1028 VNB.n1026 25.263
R2446 VNB.n1088 VNB.n1086 25.263
R2447 VNB.n1162 VNB.n1160 25.263
R2448 VNB.n1357 VNB.n1355 25.263
R2449 VNB.n7 VNB.n5 25.263
R2450 VNB.n177 VNB.n176 24.383
R2451 VNB.n236 VNB.n235 24.383
R2452 VNB.n295 VNB.n294 24.383
R2453 VNB.n354 VNB.n353 24.383
R2454 VNB.n428 VNB.n427 24.383
R2455 VNB.n556 VNB.n555 24.383
R2456 VNB.n630 VNB.n629 24.383
R2457 VNB.n705 VNB.n704 24.383
R2458 VNB.n81 VNB.n80 24.383
R2459 VNB.n884 VNB.n883 24.383
R2460 VNB.n1026 VNB.n1025 24.383
R2461 VNB.n1086 VNB.n1085 24.383
R2462 VNB.n1160 VNB.n1159 24.383
R2463 VNB.n1355 VNB.n1354 24.383
R2464 VNB.n5 VNB.n4 24.383
R2465 VNB.n157 VNB.n154 20.452
R2466 VNB.n1387 VNB.n1386 20.452
R2467 VNB.n184 VNB.n183 16.721
R2468 VNB.n243 VNB.n242 16.721
R2469 VNB.n302 VNB.n301 16.721
R2470 VNB.n361 VNB.n360 16.721
R2471 VNB.n563 VNB.n562 16.721
R2472 VNB.n891 VNB.n890 16.721
R2473 VNB.n1093 VNB.n1092 16.721
R2474 VNB.n166 VNB.n165 13.653
R2475 VNB.n165 VNB.n164 13.653
R2476 VNB.n163 VNB.n162 13.653
R2477 VNB.n162 VNB.n161 13.653
R2478 VNB.n160 VNB.n159 13.653
R2479 VNB.n159 VNB.n158 13.653
R2480 VNB.n174 VNB.n173 13.653
R2481 VNB.n173 VNB.n172 13.653
R2482 VNB.n185 VNB.n184 13.653
R2483 VNB.n189 VNB.n188 13.653
R2484 VNB.n188 VNB.n187 13.653
R2485 VNB.n193 VNB.n192 13.653
R2486 VNB.n192 VNB.n191 13.653
R2487 VNB.n215 VNB.n214 13.653
R2488 VNB.n214 VNB.n213 13.653
R2489 VNB.n219 VNB.n218 13.653
R2490 VNB.n218 VNB.n217 13.653
R2491 VNB.n223 VNB.n222 13.653
R2492 VNB.n222 VNB.n221 13.653
R2493 VNB.n227 VNB.n226 13.653
R2494 VNB.n226 VNB.n225 13.653
R2495 VNB.n233 VNB.n232 13.653
R2496 VNB.n232 VNB.n231 13.653
R2497 VNB.n244 VNB.n243 13.653
R2498 VNB.n248 VNB.n247 13.653
R2499 VNB.n247 VNB.n246 13.653
R2500 VNB.n252 VNB.n251 13.653
R2501 VNB.n251 VNB.n250 13.653
R2502 VNB.n274 VNB.n273 13.653
R2503 VNB.n273 VNB.n272 13.653
R2504 VNB.n278 VNB.n277 13.653
R2505 VNB.n277 VNB.n276 13.653
R2506 VNB.n282 VNB.n281 13.653
R2507 VNB.n281 VNB.n280 13.653
R2508 VNB.n286 VNB.n285 13.653
R2509 VNB.n285 VNB.n284 13.653
R2510 VNB.n292 VNB.n291 13.653
R2511 VNB.n291 VNB.n290 13.653
R2512 VNB.n303 VNB.n302 13.653
R2513 VNB.n307 VNB.n306 13.653
R2514 VNB.n306 VNB.n305 13.653
R2515 VNB.n311 VNB.n310 13.653
R2516 VNB.n310 VNB.n309 13.653
R2517 VNB.n333 VNB.n332 13.653
R2518 VNB.n332 VNB.n331 13.653
R2519 VNB.n337 VNB.n336 13.653
R2520 VNB.n336 VNB.n335 13.653
R2521 VNB.n341 VNB.n340 13.653
R2522 VNB.n340 VNB.n339 13.653
R2523 VNB.n345 VNB.n344 13.653
R2524 VNB.n344 VNB.n343 13.653
R2525 VNB.n351 VNB.n350 13.653
R2526 VNB.n350 VNB.n349 13.653
R2527 VNB.n362 VNB.n361 13.653
R2528 VNB.n366 VNB.n365 13.653
R2529 VNB.n365 VNB.n364 13.653
R2530 VNB.n370 VNB.n369 13.653
R2531 VNB.n369 VNB.n368 13.653
R2532 VNB.n392 VNB.n391 13.653
R2533 VNB.n391 VNB.n390 13.653
R2534 VNB.n396 VNB.n395 13.653
R2535 VNB.n395 VNB.n394 13.653
R2536 VNB.n400 VNB.n399 13.653
R2537 VNB.n399 VNB.n398 13.653
R2538 VNB.n404 VNB.n403 13.653
R2539 VNB.n403 VNB.n402 13.653
R2540 VNB.n408 VNB.n407 13.653
R2541 VNB.n407 VNB.n406 13.653
R2542 VNB.n412 VNB.n411 13.653
R2543 VNB.n411 VNB.n410 13.653
R2544 VNB.n416 VNB.n415 13.653
R2545 VNB.n415 VNB.n414 13.653
R2546 VNB.n420 VNB.n419 13.653
R2547 VNB.n419 VNB.n418 13.653
R2548 VNB.n425 VNB.n424 13.653
R2549 VNB.n424 VNB.n423 13.653
R2550 VNB.n437 VNB.n436 13.653
R2551 VNB.n436 VNB.n435 13.653
R2552 VNB.n441 VNB.n440 13.653
R2553 VNB.n440 VNB.n439 13.653
R2554 VNB.n445 VNB.n444 13.653
R2555 VNB.n444 VNB.n443 13.653
R2556 VNB.n467 VNB.n466 13.653
R2557 VNB.n466 VNB.n465 13.653
R2558 VNB.n471 VNB.n470 13.653
R2559 VNB.n470 VNB.n469 13.653
R2560 VNB.n475 VNB.n474 13.653
R2561 VNB.n474 VNB.n473 13.653
R2562 VNB.n479 VNB.n478 13.653
R2563 VNB.n478 VNB.n477 13.653
R2564 VNB.n483 VNB.n482 13.653
R2565 VNB.n482 VNB.n481 13.653
R2566 VNB.n487 VNB.n486 13.653
R2567 VNB.n486 VNB.n485 13.653
R2568 VNB.n491 VNB.n490 13.653
R2569 VNB.n490 VNB.n489 13.653
R2570 VNB.n495 VNB.n494 13.653
R2571 VNB.n494 VNB.n493 13.653
R2572 VNB.n499 VNB.n498 13.653
R2573 VNB.n498 VNB.n497 13.653
R2574 VNB.n505 VNB.n504 13.653
R2575 VNB.n509 VNB.n508 13.653
R2576 VNB.n508 VNB.n507 13.653
R2577 VNB.n513 VNB.n512 13.653
R2578 VNB.n512 VNB.n511 13.653
R2579 VNB.n535 VNB.n534 13.653
R2580 VNB.n534 VNB.n533 13.653
R2581 VNB.n539 VNB.n538 13.653
R2582 VNB.n538 VNB.n537 13.653
R2583 VNB.n543 VNB.n542 13.653
R2584 VNB.n542 VNB.n541 13.653
R2585 VNB.n547 VNB.n546 13.653
R2586 VNB.n546 VNB.n545 13.653
R2587 VNB.n553 VNB.n552 13.653
R2588 VNB.n552 VNB.n551 13.653
R2589 VNB.n564 VNB.n563 13.653
R2590 VNB.n568 VNB.n567 13.653
R2591 VNB.n567 VNB.n566 13.653
R2592 VNB.n572 VNB.n571 13.653
R2593 VNB.n571 VNB.n570 13.653
R2594 VNB.n594 VNB.n593 13.653
R2595 VNB.n593 VNB.n592 13.653
R2596 VNB.n598 VNB.n597 13.653
R2597 VNB.n597 VNB.n596 13.653
R2598 VNB.n602 VNB.n601 13.653
R2599 VNB.n601 VNB.n600 13.653
R2600 VNB.n606 VNB.n605 13.653
R2601 VNB.n605 VNB.n604 13.653
R2602 VNB.n610 VNB.n609 13.653
R2603 VNB.n609 VNB.n608 13.653
R2604 VNB.n614 VNB.n613 13.653
R2605 VNB.n613 VNB.n612 13.653
R2606 VNB.n618 VNB.n617 13.653
R2607 VNB.n617 VNB.n616 13.653
R2608 VNB.n622 VNB.n621 13.653
R2609 VNB.n621 VNB.n620 13.653
R2610 VNB.n627 VNB.n626 13.653
R2611 VNB.n626 VNB.n625 13.653
R2612 VNB.n639 VNB.n638 13.653
R2613 VNB.n638 VNB.n637 13.653
R2614 VNB.n643 VNB.n642 13.653
R2615 VNB.n642 VNB.n641 13.653
R2616 VNB.n647 VNB.n646 13.653
R2617 VNB.n646 VNB.n645 13.653
R2618 VNB.n669 VNB.n668 13.653
R2619 VNB.n668 VNB.n667 13.653
R2620 VNB.n673 VNB.n672 13.653
R2621 VNB.n672 VNB.n671 13.653
R2622 VNB.n677 VNB.n676 13.653
R2623 VNB.n676 VNB.n675 13.653
R2624 VNB.n681 VNB.n680 13.653
R2625 VNB.n680 VNB.n679 13.653
R2626 VNB.n685 VNB.n684 13.653
R2627 VNB.n684 VNB.n683 13.653
R2628 VNB.n689 VNB.n688 13.653
R2629 VNB.n688 VNB.n687 13.653
R2630 VNB.n693 VNB.n692 13.653
R2631 VNB.n692 VNB.n691 13.653
R2632 VNB.n697 VNB.n696 13.653
R2633 VNB.n696 VNB.n695 13.653
R2634 VNB.n702 VNB.n701 13.653
R2635 VNB.n701 VNB.n700 13.653
R2636 VNB.n714 VNB.n713 13.653
R2637 VNB.n713 VNB.n712 13.653
R2638 VNB.n718 VNB.n717 13.653
R2639 VNB.n717 VNB.n716 13.653
R2640 VNB.n722 VNB.n721 13.653
R2641 VNB.n721 VNB.n720 13.653
R2642 VNB.n744 VNB.n743 13.653
R2643 VNB.n743 VNB.n742 13.653
R2644 VNB.n748 VNB.n747 13.653
R2645 VNB.n747 VNB.n746 13.653
R2646 VNB.n752 VNB.n751 13.653
R2647 VNB.n751 VNB.n750 13.653
R2648 VNB.n756 VNB.n755 13.653
R2649 VNB.n755 VNB.n754 13.653
R2650 VNB.n760 VNB.n759 13.653
R2651 VNB.n759 VNB.n758 13.653
R2652 VNB.n766 VNB.n765 13.653
R2653 VNB.n770 VNB.n769 13.653
R2654 VNB.n769 VNB.n768 13.653
R2655 VNB.n774 VNB.n773 13.653
R2656 VNB.n773 VNB.n772 13.653
R2657 VNB.n104 VNB.n103 13.653
R2658 VNB.n103 VNB.n102 13.653
R2659 VNB.n107 VNB.n106 13.653
R2660 VNB.n106 VNB.n105 13.653
R2661 VNB.n110 VNB.n109 13.653
R2662 VNB.n109 VNB.n108 13.653
R2663 VNB.n113 VNB.n112 13.653
R2664 VNB.n112 VNB.n111 13.653
R2665 VNB.n116 VNB.n115 13.653
R2666 VNB.n115 VNB.n114 13.653
R2667 VNB.n119 VNB.n118 13.653
R2668 VNB.n118 VNB.n117 13.653
R2669 VNB.n122 VNB.n121 13.653
R2670 VNB.n121 VNB.n120 13.653
R2671 VNB.n125 VNB.n124 13.653
R2672 VNB.n124 VNB.n123 13.653
R2673 VNB.n129 VNB.n128 13.653
R2674 VNB.n128 VNB.n127 13.653
R2675 VNB.n134 VNB.n133 13.653
R2676 VNB.n133 VNB.n132 13.653
R2677 VNB.n139 VNB.n138 13.653
R2678 VNB.n138 VNB.n137 13.653
R2679 VNB.n790 VNB.n789 13.653
R2680 VNB.n789 VNB.n788 13.653
R2681 VNB.n795 VNB.n794 13.653
R2682 VNB.n794 VNB.n793 13.653
R2683 VNB.n799 VNB.n798 13.653
R2684 VNB.n798 VNB.n797 13.653
R2685 VNB.n803 VNB.n802 13.653
R2686 VNB.n802 VNB.n801 13.653
R2687 VNB.n807 VNB.n806 13.653
R2688 VNB.n806 VNB.n805 13.653
R2689 VNB.n811 VNB.n810 13.653
R2690 VNB.n810 VNB.n809 13.653
R2691 VNB.n815 VNB.n814 13.653
R2692 VNB.n814 VNB.n813 13.653
R2693 VNB.n819 VNB.n818 13.653
R2694 VNB.n818 VNB.n817 13.653
R2695 VNB.n823 VNB.n822 13.653
R2696 VNB.n822 VNB.n821 13.653
R2697 VNB.n827 VNB.n826 13.653
R2698 VNB.n826 VNB.n825 13.653
R2699 VNB.n833 VNB.n832 13.653
R2700 VNB.n837 VNB.n836 13.653
R2701 VNB.n836 VNB.n835 13.653
R2702 VNB.n841 VNB.n840 13.653
R2703 VNB.n840 VNB.n839 13.653
R2704 VNB.n863 VNB.n862 13.653
R2705 VNB.n862 VNB.n861 13.653
R2706 VNB.n867 VNB.n866 13.653
R2707 VNB.n866 VNB.n865 13.653
R2708 VNB.n871 VNB.n870 13.653
R2709 VNB.n870 VNB.n869 13.653
R2710 VNB.n875 VNB.n874 13.653
R2711 VNB.n874 VNB.n873 13.653
R2712 VNB.n881 VNB.n880 13.653
R2713 VNB.n880 VNB.n879 13.653
R2714 VNB.n892 VNB.n891 13.653
R2715 VNB.n896 VNB.n895 13.653
R2716 VNB.n895 VNB.n894 13.653
R2717 VNB.n900 VNB.n899 13.653
R2718 VNB.n899 VNB.n898 13.653
R2719 VNB.n922 VNB.n921 13.653
R2720 VNB.n921 VNB.n920 13.653
R2721 VNB.n926 VNB.n925 13.653
R2722 VNB.n925 VNB.n924 13.653
R2723 VNB.n930 VNB.n929 13.653
R2724 VNB.n929 VNB.n928 13.653
R2725 VNB.n934 VNB.n933 13.653
R2726 VNB.n933 VNB.n932 13.653
R2727 VNB.n938 VNB.n937 13.653
R2728 VNB.n937 VNB.n936 13.653
R2729 VNB.n942 VNB.n941 13.653
R2730 VNB.n941 VNB.n940 13.653
R2731 VNB.n946 VNB.n945 13.653
R2732 VNB.n945 VNB.n944 13.653
R2733 VNB.n950 VNB.n949 13.653
R2734 VNB.n949 VNB.n948 13.653
R2735 VNB.n954 VNB.n953 13.653
R2736 VNB.n953 VNB.n952 13.653
R2737 VNB.n960 VNB.n959 13.653
R2738 VNB.n964 VNB.n963 13.653
R2739 VNB.n963 VNB.n962 13.653
R2740 VNB.n968 VNB.n967 13.653
R2741 VNB.n967 VNB.n966 13.653
R2742 VNB.n990 VNB.n989 13.653
R2743 VNB.n989 VNB.n988 13.653
R2744 VNB.n994 VNB.n993 13.653
R2745 VNB.n993 VNB.n992 13.653
R2746 VNB.n998 VNB.n997 13.653
R2747 VNB.n997 VNB.n996 13.653
R2748 VNB.n1002 VNB.n1001 13.653
R2749 VNB.n1001 VNB.n1000 13.653
R2750 VNB.n1006 VNB.n1005 13.653
R2751 VNB.n1005 VNB.n1004 13.653
R2752 VNB.n1010 VNB.n1009 13.653
R2753 VNB.n1009 VNB.n1008 13.653
R2754 VNB.n1014 VNB.n1013 13.653
R2755 VNB.n1013 VNB.n1012 13.653
R2756 VNB.n1018 VNB.n1017 13.653
R2757 VNB.n1017 VNB.n1016 13.653
R2758 VNB.n1023 VNB.n1022 13.653
R2759 VNB.n1022 VNB.n1021 13.653
R2760 VNB.n1035 VNB.n1034 13.653
R2761 VNB.n1034 VNB.n1033 13.653
R2762 VNB.n1039 VNB.n1038 13.653
R2763 VNB.n1038 VNB.n1037 13.653
R2764 VNB.n1043 VNB.n1042 13.653
R2765 VNB.n1042 VNB.n1041 13.653
R2766 VNB.n1065 VNB.n1064 13.653
R2767 VNB.n1064 VNB.n1063 13.653
R2768 VNB.n1069 VNB.n1068 13.653
R2769 VNB.n1068 VNB.n1067 13.653
R2770 VNB.n1073 VNB.n1072 13.653
R2771 VNB.n1072 VNB.n1071 13.653
R2772 VNB.n1077 VNB.n1076 13.653
R2773 VNB.n1076 VNB.n1075 13.653
R2774 VNB.n1083 VNB.n1082 13.653
R2775 VNB.n1082 VNB.n1081 13.653
R2776 VNB.n1094 VNB.n1093 13.653
R2777 VNB.n1098 VNB.n1097 13.653
R2778 VNB.n1097 VNB.n1096 13.653
R2779 VNB.n1102 VNB.n1101 13.653
R2780 VNB.n1101 VNB.n1100 13.653
R2781 VNB.n1124 VNB.n1123 13.653
R2782 VNB.n1123 VNB.n1122 13.653
R2783 VNB.n1128 VNB.n1127 13.653
R2784 VNB.n1127 VNB.n1126 13.653
R2785 VNB.n1132 VNB.n1131 13.653
R2786 VNB.n1131 VNB.n1130 13.653
R2787 VNB.n1136 VNB.n1135 13.653
R2788 VNB.n1135 VNB.n1134 13.653
R2789 VNB.n1140 VNB.n1139 13.653
R2790 VNB.n1139 VNB.n1138 13.653
R2791 VNB.n1144 VNB.n1143 13.653
R2792 VNB.n1143 VNB.n1142 13.653
R2793 VNB.n1148 VNB.n1147 13.653
R2794 VNB.n1147 VNB.n1146 13.653
R2795 VNB.n1152 VNB.n1151 13.653
R2796 VNB.n1151 VNB.n1150 13.653
R2797 VNB.n1157 VNB.n1156 13.653
R2798 VNB.n1156 VNB.n1155 13.653
R2799 VNB.n1169 VNB.n1168 13.653
R2800 VNB.n1168 VNB.n1167 13.653
R2801 VNB.n1173 VNB.n1172 13.653
R2802 VNB.n1172 VNB.n1171 13.653
R2803 VNB.n1177 VNB.n1176 13.653
R2804 VNB.n1176 VNB.n1175 13.653
R2805 VNB.n1199 VNB.n1198 13.653
R2806 VNB.n1198 VNB.n1197 13.653
R2807 VNB.n1203 VNB.n1202 13.653
R2808 VNB.n1202 VNB.n1201 13.653
R2809 VNB.n1207 VNB.n1206 13.653
R2810 VNB.n1206 VNB.n1205 13.653
R2811 VNB.n1211 VNB.n1210 13.653
R2812 VNB.n1210 VNB.n1209 13.653
R2813 VNB.n1215 VNB.n1214 13.653
R2814 VNB.n1214 VNB.n1213 13.653
R2815 VNB.n1219 VNB.n1218 13.653
R2816 VNB.n1218 VNB.n1217 13.653
R2817 VNB.n1223 VNB.n1222 13.653
R2818 VNB.n1222 VNB.n1221 13.653
R2819 VNB.n1227 VNB.n1226 13.653
R2820 VNB.n1226 VNB.n1225 13.653
R2821 VNB.n1231 VNB.n1230 13.653
R2822 VNB.n1230 VNB.n1229 13.653
R2823 VNB.n1237 VNB.n1236 13.653
R2824 VNB.n1241 VNB.n1240 13.653
R2825 VNB.n1240 VNB.n1239 13.653
R2826 VNB.n1245 VNB.n1244 13.653
R2827 VNB.n1244 VNB.n1243 13.653
R2828 VNB.n1267 VNB.n1266 13.653
R2829 VNB.n1266 VNB.n1265 13.653
R2830 VNB.n1271 VNB.n1270 13.653
R2831 VNB.n1270 VNB.n1269 13.653
R2832 VNB.n1275 VNB.n1274 13.653
R2833 VNB.n1274 VNB.n1273 13.653
R2834 VNB.n1279 VNB.n1278 13.653
R2835 VNB.n1278 VNB.n1277 13.653
R2836 VNB.n1283 VNB.n1282 13.653
R2837 VNB.n1282 VNB.n1281 13.653
R2838 VNB.n1289 VNB.n1288 13.653
R2839 VNB.n1293 VNB.n1292 13.653
R2840 VNB.n1292 VNB.n1291 13.653
R2841 VNB.n1297 VNB.n1296 13.653
R2842 VNB.n1296 VNB.n1295 13.653
R2843 VNB.n1319 VNB.n1318 13.653
R2844 VNB.n1318 VNB.n1317 13.653
R2845 VNB.n1323 VNB.n1322 13.653
R2846 VNB.n1322 VNB.n1321 13.653
R2847 VNB.n1327 VNB.n1326 13.653
R2848 VNB.n1326 VNB.n1325 13.653
R2849 VNB.n1331 VNB.n1330 13.653
R2850 VNB.n1330 VNB.n1329 13.653
R2851 VNB.n1335 VNB.n1334 13.653
R2852 VNB.n1334 VNB.n1333 13.653
R2853 VNB.n1339 VNB.n1338 13.653
R2854 VNB.n1338 VNB.n1337 13.653
R2855 VNB.n1343 VNB.n1342 13.653
R2856 VNB.n1342 VNB.n1341 13.653
R2857 VNB.n1347 VNB.n1346 13.653
R2858 VNB.n1346 VNB.n1345 13.653
R2859 VNB.n1352 VNB.n1351 13.653
R2860 VNB.n1351 VNB.n1350 13.653
R2861 VNB.n1364 VNB.n1363 13.653
R2862 VNB.n1363 VNB.n1362 13.653
R2863 VNB.n1368 VNB.n1367 13.653
R2864 VNB.n1367 VNB.n1366 13.653
R2865 VNB.n1372 VNB.n1371 13.653
R2866 VNB.n1371 VNB.n1370 13.653
R2867 VNB.n28 VNB.n27 13.653
R2868 VNB.n27 VNB.n26 13.653
R2869 VNB.n31 VNB.n30 13.653
R2870 VNB.n30 VNB.n29 13.653
R2871 VNB.n34 VNB.n33 13.653
R2872 VNB.n33 VNB.n32 13.653
R2873 VNB.n37 VNB.n36 13.653
R2874 VNB.n36 VNB.n35 13.653
R2875 VNB.n40 VNB.n39 13.653
R2876 VNB.n39 VNB.n38 13.653
R2877 VNB.n43 VNB.n42 13.653
R2878 VNB.n42 VNB.n41 13.653
R2879 VNB.n46 VNB.n45 13.653
R2880 VNB.n45 VNB.n44 13.653
R2881 VNB.n49 VNB.n48 13.653
R2882 VNB.n48 VNB.n47 13.653
R2883 VNB.n53 VNB.n52 13.653
R2884 VNB.n52 VNB.n51 13.653
R2885 VNB.n58 VNB.n57 13.653
R2886 VNB.n57 VNB.n56 13.653
R2887 VNB.n63 VNB.n62 13.653
R2888 VNB.n62 VNB.n61 13.653
R2889 VNB.n1386 VNB.n0 13.653
R2890 VNB VNB.n0 13.653
R2891 VNB.n157 VNB.n156 13.653
R2892 VNB.n156 VNB.n155 13.653
R2893 VNB.n1394 VNB.n1391 13.577
R2894 VNB.n142 VNB.n140 13.276
R2895 VNB.n154 VNB.n142 13.276
R2896 VNB.n197 VNB.n195 13.276
R2897 VNB.n210 VNB.n197 13.276
R2898 VNB.n256 VNB.n254 13.276
R2899 VNB.n269 VNB.n256 13.276
R2900 VNB.n315 VNB.n313 13.276
R2901 VNB.n328 VNB.n315 13.276
R2902 VNB.n374 VNB.n372 13.276
R2903 VNB.n387 VNB.n374 13.276
R2904 VNB.n449 VNB.n447 13.276
R2905 VNB.n462 VNB.n449 13.276
R2906 VNB.n517 VNB.n515 13.276
R2907 VNB.n530 VNB.n517 13.276
R2908 VNB.n576 VNB.n574 13.276
R2909 VNB.n589 VNB.n576 13.276
R2910 VNB.n651 VNB.n649 13.276
R2911 VNB.n664 VNB.n651 13.276
R2912 VNB.n726 VNB.n724 13.276
R2913 VNB.n739 VNB.n726 13.276
R2914 VNB.n86 VNB.n84 13.276
R2915 VNB.n99 VNB.n86 13.276
R2916 VNB.n66 VNB.n64 13.276
R2917 VNB.n79 VNB.n66 13.276
R2918 VNB.n845 VNB.n843 13.276
R2919 VNB.n858 VNB.n845 13.276
R2920 VNB.n904 VNB.n902 13.276
R2921 VNB.n917 VNB.n904 13.276
R2922 VNB.n972 VNB.n970 13.276
R2923 VNB.n985 VNB.n972 13.276
R2924 VNB.n1047 VNB.n1045 13.276
R2925 VNB.n1060 VNB.n1047 13.276
R2926 VNB.n1106 VNB.n1104 13.276
R2927 VNB.n1119 VNB.n1106 13.276
R2928 VNB.n1181 VNB.n1179 13.276
R2929 VNB.n1194 VNB.n1181 13.276
R2930 VNB.n1249 VNB.n1247 13.276
R2931 VNB.n1262 VNB.n1249 13.276
R2932 VNB.n1301 VNB.n1299 13.276
R2933 VNB.n1314 VNB.n1301 13.276
R2934 VNB.n10 VNB.n8 13.276
R2935 VNB.n23 VNB.n10 13.276
R2936 VNB.n166 VNB.n163 13.276
R2937 VNB.n163 VNB.n160 13.276
R2938 VNB.n215 VNB.n211 13.276
R2939 VNB.n274 VNB.n270 13.276
R2940 VNB.n333 VNB.n329 13.276
R2941 VNB.n392 VNB.n388 13.276
R2942 VNB.n467 VNB.n463 13.276
R2943 VNB.n535 VNB.n531 13.276
R2944 VNB.n594 VNB.n590 13.276
R2945 VNB.n669 VNB.n665 13.276
R2946 VNB.n744 VNB.n740 13.276
R2947 VNB.n104 VNB.n100 13.276
R2948 VNB.n107 VNB.n104 13.276
R2949 VNB.n110 VNB.n107 13.276
R2950 VNB.n113 VNB.n110 13.276
R2951 VNB.n116 VNB.n113 13.276
R2952 VNB.n119 VNB.n116 13.276
R2953 VNB.n122 VNB.n119 13.276
R2954 VNB.n125 VNB.n122 13.276
R2955 VNB.n129 VNB.n125 13.276
R2956 VNB.n134 VNB.n129 13.276
R2957 VNB.n790 VNB.n139 13.276
R2958 VNB.n791 VNB.n790 13.276
R2959 VNB.n795 VNB.n791 13.276
R2960 VNB.n863 VNB.n859 13.276
R2961 VNB.n922 VNB.n918 13.276
R2962 VNB.n990 VNB.n986 13.276
R2963 VNB.n1065 VNB.n1061 13.276
R2964 VNB.n1124 VNB.n1120 13.276
R2965 VNB.n1199 VNB.n1195 13.276
R2966 VNB.n1267 VNB.n1263 13.276
R2967 VNB.n1319 VNB.n1315 13.276
R2968 VNB.n28 VNB.n24 13.276
R2969 VNB.n31 VNB.n28 13.276
R2970 VNB.n34 VNB.n31 13.276
R2971 VNB.n37 VNB.n34 13.276
R2972 VNB.n40 VNB.n37 13.276
R2973 VNB.n43 VNB.n40 13.276
R2974 VNB.n46 VNB.n43 13.276
R2975 VNB.n49 VNB.n46 13.276
R2976 VNB.n53 VNB.n49 13.276
R2977 VNB.n58 VNB.n53 13.276
R2978 VNB.n1386 VNB.n63 13.276
R2979 VNB.n3 VNB.n1 13.276
R2980 VNB.n1387 VNB.n3 13.276
R2981 VNB.n139 VNB.n135 12.02
R2982 VNB.n63 VNB.n59 12.02
R2983 VNB.n1396 VNB.n1395 7.5
R2984 VNB.n203 VNB.n202 7.5
R2985 VNB.n199 VNB.n198 7.5
R2986 VNB.n197 VNB.n196 7.5
R2987 VNB.n210 VNB.n209 7.5
R2988 VNB.n262 VNB.n261 7.5
R2989 VNB.n258 VNB.n257 7.5
R2990 VNB.n256 VNB.n255 7.5
R2991 VNB.n269 VNB.n268 7.5
R2992 VNB.n321 VNB.n320 7.5
R2993 VNB.n317 VNB.n316 7.5
R2994 VNB.n315 VNB.n314 7.5
R2995 VNB.n328 VNB.n327 7.5
R2996 VNB.n380 VNB.n379 7.5
R2997 VNB.n376 VNB.n375 7.5
R2998 VNB.n374 VNB.n373 7.5
R2999 VNB.n387 VNB.n386 7.5
R3000 VNB.n455 VNB.n454 7.5
R3001 VNB.n451 VNB.n450 7.5
R3002 VNB.n449 VNB.n448 7.5
R3003 VNB.n462 VNB.n461 7.5
R3004 VNB.n523 VNB.n522 7.5
R3005 VNB.n519 VNB.n518 7.5
R3006 VNB.n517 VNB.n516 7.5
R3007 VNB.n530 VNB.n529 7.5
R3008 VNB.n582 VNB.n581 7.5
R3009 VNB.n578 VNB.n577 7.5
R3010 VNB.n576 VNB.n575 7.5
R3011 VNB.n589 VNB.n588 7.5
R3012 VNB.n657 VNB.n656 7.5
R3013 VNB.n653 VNB.n652 7.5
R3014 VNB.n651 VNB.n650 7.5
R3015 VNB.n664 VNB.n663 7.5
R3016 VNB.n732 VNB.n731 7.5
R3017 VNB.n728 VNB.n727 7.5
R3018 VNB.n726 VNB.n725 7.5
R3019 VNB.n739 VNB.n738 7.5
R3020 VNB.n92 VNB.n91 7.5
R3021 VNB.n88 VNB.n87 7.5
R3022 VNB.n86 VNB.n85 7.5
R3023 VNB.n99 VNB.n98 7.5
R3024 VNB.n72 VNB.n71 7.5
R3025 VNB.n68 VNB.n67 7.5
R3026 VNB.n66 VNB.n65 7.5
R3027 VNB.n79 VNB.n78 7.5
R3028 VNB.n851 VNB.n850 7.5
R3029 VNB.n847 VNB.n846 7.5
R3030 VNB.n845 VNB.n844 7.5
R3031 VNB.n858 VNB.n857 7.5
R3032 VNB.n910 VNB.n909 7.5
R3033 VNB.n906 VNB.n905 7.5
R3034 VNB.n904 VNB.n903 7.5
R3035 VNB.n917 VNB.n916 7.5
R3036 VNB.n978 VNB.n977 7.5
R3037 VNB.n974 VNB.n973 7.5
R3038 VNB.n972 VNB.n971 7.5
R3039 VNB.n985 VNB.n984 7.5
R3040 VNB.n1053 VNB.n1052 7.5
R3041 VNB.n1049 VNB.n1048 7.5
R3042 VNB.n1047 VNB.n1046 7.5
R3043 VNB.n1060 VNB.n1059 7.5
R3044 VNB.n1112 VNB.n1111 7.5
R3045 VNB.n1108 VNB.n1107 7.5
R3046 VNB.n1106 VNB.n1105 7.5
R3047 VNB.n1119 VNB.n1118 7.5
R3048 VNB.n1187 VNB.n1186 7.5
R3049 VNB.n1183 VNB.n1182 7.5
R3050 VNB.n1181 VNB.n1180 7.5
R3051 VNB.n1194 VNB.n1193 7.5
R3052 VNB.n1255 VNB.n1254 7.5
R3053 VNB.n1251 VNB.n1250 7.5
R3054 VNB.n1249 VNB.n1248 7.5
R3055 VNB.n1262 VNB.n1261 7.5
R3056 VNB.n1307 VNB.n1306 7.5
R3057 VNB.n1303 VNB.n1302 7.5
R3058 VNB.n1301 VNB.n1300 7.5
R3059 VNB.n1314 VNB.n1313 7.5
R3060 VNB.n16 VNB.n15 7.5
R3061 VNB.n12 VNB.n11 7.5
R3062 VNB.n10 VNB.n9 7.5
R3063 VNB.n23 VNB.n22 7.5
R3064 VNB.n1388 VNB.n1387 7.5
R3065 VNB.n3 VNB.n2 7.5
R3066 VNB.n1393 VNB.n1392 7.5
R3067 VNB.n148 VNB.n147 7.5
R3068 VNB.n144 VNB.n143 7.5
R3069 VNB.n142 VNB.n141 7.5
R3070 VNB.n154 VNB.n153 7.5
R3071 VNB.n211 VNB.n210 7.176
R3072 VNB.n270 VNB.n269 7.176
R3073 VNB.n329 VNB.n328 7.176
R3074 VNB.n388 VNB.n387 7.176
R3075 VNB.n463 VNB.n462 7.176
R3076 VNB.n531 VNB.n530 7.176
R3077 VNB.n590 VNB.n589 7.176
R3078 VNB.n665 VNB.n664 7.176
R3079 VNB.n740 VNB.n739 7.176
R3080 VNB.n100 VNB.n99 7.176
R3081 VNB.n791 VNB.n79 7.176
R3082 VNB.n859 VNB.n858 7.176
R3083 VNB.n918 VNB.n917 7.176
R3084 VNB.n986 VNB.n985 7.176
R3085 VNB.n1061 VNB.n1060 7.176
R3086 VNB.n1120 VNB.n1119 7.176
R3087 VNB.n1195 VNB.n1194 7.176
R3088 VNB.n1263 VNB.n1262 7.176
R3089 VNB.n1315 VNB.n1314 7.176
R3090 VNB.n24 VNB.n23 7.176
R3091 VNB.n1398 VNB.n1396 7.011
R3092 VNB.n206 VNB.n203 7.011
R3093 VNB.n201 VNB.n199 7.011
R3094 VNB.n265 VNB.n262 7.011
R3095 VNB.n260 VNB.n258 7.011
R3096 VNB.n324 VNB.n321 7.011
R3097 VNB.n319 VNB.n317 7.011
R3098 VNB.n383 VNB.n380 7.011
R3099 VNB.n378 VNB.n376 7.011
R3100 VNB.n458 VNB.n455 7.011
R3101 VNB.n453 VNB.n451 7.011
R3102 VNB.n526 VNB.n523 7.011
R3103 VNB.n521 VNB.n519 7.011
R3104 VNB.n585 VNB.n582 7.011
R3105 VNB.n580 VNB.n578 7.011
R3106 VNB.n660 VNB.n657 7.011
R3107 VNB.n655 VNB.n653 7.011
R3108 VNB.n735 VNB.n732 7.011
R3109 VNB.n730 VNB.n728 7.011
R3110 VNB.n95 VNB.n92 7.011
R3111 VNB.n90 VNB.n88 7.011
R3112 VNB.n75 VNB.n72 7.011
R3113 VNB.n70 VNB.n68 7.011
R3114 VNB.n854 VNB.n851 7.011
R3115 VNB.n849 VNB.n847 7.011
R3116 VNB.n913 VNB.n910 7.011
R3117 VNB.n908 VNB.n906 7.011
R3118 VNB.n981 VNB.n978 7.011
R3119 VNB.n976 VNB.n974 7.011
R3120 VNB.n1056 VNB.n1053 7.011
R3121 VNB.n1051 VNB.n1049 7.011
R3122 VNB.n1115 VNB.n1112 7.011
R3123 VNB.n1110 VNB.n1108 7.011
R3124 VNB.n1190 VNB.n1187 7.011
R3125 VNB.n1185 VNB.n1183 7.011
R3126 VNB.n1258 VNB.n1255 7.011
R3127 VNB.n1253 VNB.n1251 7.011
R3128 VNB.n1310 VNB.n1307 7.011
R3129 VNB.n1305 VNB.n1303 7.011
R3130 VNB.n19 VNB.n16 7.011
R3131 VNB.n14 VNB.n12 7.011
R3132 VNB.n150 VNB.n148 7.011
R3133 VNB.n146 VNB.n144 7.011
R3134 VNB.n209 VNB.n208 7.01
R3135 VNB.n201 VNB.n200 7.01
R3136 VNB.n206 VNB.n205 7.01
R3137 VNB.n268 VNB.n267 7.01
R3138 VNB.n260 VNB.n259 7.01
R3139 VNB.n265 VNB.n264 7.01
R3140 VNB.n327 VNB.n326 7.01
R3141 VNB.n319 VNB.n318 7.01
R3142 VNB.n324 VNB.n323 7.01
R3143 VNB.n386 VNB.n385 7.01
R3144 VNB.n378 VNB.n377 7.01
R3145 VNB.n383 VNB.n382 7.01
R3146 VNB.n461 VNB.n460 7.01
R3147 VNB.n453 VNB.n452 7.01
R3148 VNB.n458 VNB.n457 7.01
R3149 VNB.n529 VNB.n528 7.01
R3150 VNB.n521 VNB.n520 7.01
R3151 VNB.n526 VNB.n525 7.01
R3152 VNB.n588 VNB.n587 7.01
R3153 VNB.n580 VNB.n579 7.01
R3154 VNB.n585 VNB.n584 7.01
R3155 VNB.n663 VNB.n662 7.01
R3156 VNB.n655 VNB.n654 7.01
R3157 VNB.n660 VNB.n659 7.01
R3158 VNB.n738 VNB.n737 7.01
R3159 VNB.n730 VNB.n729 7.01
R3160 VNB.n735 VNB.n734 7.01
R3161 VNB.n98 VNB.n97 7.01
R3162 VNB.n90 VNB.n89 7.01
R3163 VNB.n95 VNB.n94 7.01
R3164 VNB.n78 VNB.n77 7.01
R3165 VNB.n70 VNB.n69 7.01
R3166 VNB.n75 VNB.n74 7.01
R3167 VNB.n857 VNB.n856 7.01
R3168 VNB.n849 VNB.n848 7.01
R3169 VNB.n854 VNB.n853 7.01
R3170 VNB.n916 VNB.n915 7.01
R3171 VNB.n908 VNB.n907 7.01
R3172 VNB.n913 VNB.n912 7.01
R3173 VNB.n984 VNB.n983 7.01
R3174 VNB.n976 VNB.n975 7.01
R3175 VNB.n981 VNB.n980 7.01
R3176 VNB.n1059 VNB.n1058 7.01
R3177 VNB.n1051 VNB.n1050 7.01
R3178 VNB.n1056 VNB.n1055 7.01
R3179 VNB.n1118 VNB.n1117 7.01
R3180 VNB.n1110 VNB.n1109 7.01
R3181 VNB.n1115 VNB.n1114 7.01
R3182 VNB.n1193 VNB.n1192 7.01
R3183 VNB.n1185 VNB.n1184 7.01
R3184 VNB.n1190 VNB.n1189 7.01
R3185 VNB.n1261 VNB.n1260 7.01
R3186 VNB.n1253 VNB.n1252 7.01
R3187 VNB.n1258 VNB.n1257 7.01
R3188 VNB.n1313 VNB.n1312 7.01
R3189 VNB.n1305 VNB.n1304 7.01
R3190 VNB.n1310 VNB.n1309 7.01
R3191 VNB.n22 VNB.n21 7.01
R3192 VNB.n14 VNB.n13 7.01
R3193 VNB.n19 VNB.n18 7.01
R3194 VNB.n153 VNB.n152 7.01
R3195 VNB.n146 VNB.n145 7.01
R3196 VNB.n150 VNB.n149 7.01
R3197 VNB.n1398 VNB.n1397 7.01
R3198 VNB.n1394 VNB.n1393 6.788
R3199 VNB.n1389 VNB.n1388 6.788
R3200 VNB.n167 VNB.n157 6.111
R3201 VNB.n167 VNB.n166 6.1
R3202 VNB.n185 VNB.n180 2.511
R3203 VNB.n244 VNB.n239 2.511
R3204 VNB.n303 VNB.n298 2.511
R3205 VNB.n362 VNB.n357 2.511
R3206 VNB.n564 VNB.n559 2.511
R3207 VNB.n766 VNB.n763 2.511
R3208 VNB.n892 VNB.n887 2.511
R3209 VNB.n1094 VNB.n1089 2.511
R3210 VNB.n1289 VNB.n1286 2.511
R3211 VNB.n183 VNB.n181 1.99
R3212 VNB.n242 VNB.n240 1.99
R3213 VNB.n301 VNB.n299 1.99
R3214 VNB.n360 VNB.n358 1.99
R3215 VNB.n562 VNB.n560 1.99
R3216 VNB.n890 VNB.n888 1.99
R3217 VNB.n1092 VNB.n1090 1.99
R3218 VNB.n437 VNB.n431 1.255
R3219 VNB.n505 VNB.n502 1.255
R3220 VNB.n639 VNB.n633 1.255
R3221 VNB.n714 VNB.n708 1.255
R3222 VNB.n135 VNB.n134 1.255
R3223 VNB.n833 VNB.n830 1.255
R3224 VNB.n960 VNB.n957 1.255
R3225 VNB.n1035 VNB.n1029 1.255
R3226 VNB.n1169 VNB.n1163 1.255
R3227 VNB.n1237 VNB.n1234 1.255
R3228 VNB.n1364 VNB.n1358 1.255
R3229 VNB.n59 VNB.n58 1.255
R3230 VNB.n1399 VNB.n1390 0.921
R3231 VNB.n1399 VNB.n1394 0.476
R3232 VNB.n1399 VNB.n1389 0.475
R3233 VNB.n216 VNB.n194 0.272
R3234 VNB.n275 VNB.n253 0.272
R3235 VNB.n334 VNB.n312 0.272
R3236 VNB.n393 VNB.n371 0.272
R3237 VNB.n468 VNB.n446 0.272
R3238 VNB.n536 VNB.n514 0.272
R3239 VNB.n595 VNB.n573 0.272
R3240 VNB.n670 VNB.n648 0.272
R3241 VNB.n745 VNB.n723 0.272
R3242 VNB.n776 VNB.n775 0.272
R3243 VNB.n864 VNB.n842 0.272
R3244 VNB.n923 VNB.n901 0.272
R3245 VNB.n991 VNB.n969 0.272
R3246 VNB.n1066 VNB.n1044 0.272
R3247 VNB.n1125 VNB.n1103 0.272
R3248 VNB.n1200 VNB.n1178 0.272
R3249 VNB.n1268 VNB.n1246 0.272
R3250 VNB.n1320 VNB.n1298 0.272
R3251 VNB.n1374 VNB.n1373 0.272
R3252 VNB.n207 VNB.n201 0.246
R3253 VNB.n208 VNB.n207 0.246
R3254 VNB.n207 VNB.n206 0.246
R3255 VNB.n266 VNB.n260 0.246
R3256 VNB.n267 VNB.n266 0.246
R3257 VNB.n266 VNB.n265 0.246
R3258 VNB.n325 VNB.n319 0.246
R3259 VNB.n326 VNB.n325 0.246
R3260 VNB.n325 VNB.n324 0.246
R3261 VNB.n384 VNB.n378 0.246
R3262 VNB.n385 VNB.n384 0.246
R3263 VNB.n384 VNB.n383 0.246
R3264 VNB.n459 VNB.n453 0.246
R3265 VNB.n460 VNB.n459 0.246
R3266 VNB.n459 VNB.n458 0.246
R3267 VNB.n527 VNB.n521 0.246
R3268 VNB.n528 VNB.n527 0.246
R3269 VNB.n527 VNB.n526 0.246
R3270 VNB.n586 VNB.n580 0.246
R3271 VNB.n587 VNB.n586 0.246
R3272 VNB.n586 VNB.n585 0.246
R3273 VNB.n661 VNB.n655 0.246
R3274 VNB.n662 VNB.n661 0.246
R3275 VNB.n661 VNB.n660 0.246
R3276 VNB.n736 VNB.n730 0.246
R3277 VNB.n737 VNB.n736 0.246
R3278 VNB.n736 VNB.n735 0.246
R3279 VNB.n96 VNB.n90 0.246
R3280 VNB.n97 VNB.n96 0.246
R3281 VNB.n96 VNB.n95 0.246
R3282 VNB.n76 VNB.n70 0.246
R3283 VNB.n77 VNB.n76 0.246
R3284 VNB.n76 VNB.n75 0.246
R3285 VNB.n855 VNB.n849 0.246
R3286 VNB.n856 VNB.n855 0.246
R3287 VNB.n855 VNB.n854 0.246
R3288 VNB.n914 VNB.n908 0.246
R3289 VNB.n915 VNB.n914 0.246
R3290 VNB.n914 VNB.n913 0.246
R3291 VNB.n982 VNB.n976 0.246
R3292 VNB.n983 VNB.n982 0.246
R3293 VNB.n982 VNB.n981 0.246
R3294 VNB.n1057 VNB.n1051 0.246
R3295 VNB.n1058 VNB.n1057 0.246
R3296 VNB.n1057 VNB.n1056 0.246
R3297 VNB.n1116 VNB.n1110 0.246
R3298 VNB.n1117 VNB.n1116 0.246
R3299 VNB.n1116 VNB.n1115 0.246
R3300 VNB.n1191 VNB.n1185 0.246
R3301 VNB.n1192 VNB.n1191 0.246
R3302 VNB.n1191 VNB.n1190 0.246
R3303 VNB.n1259 VNB.n1253 0.246
R3304 VNB.n1260 VNB.n1259 0.246
R3305 VNB.n1259 VNB.n1258 0.246
R3306 VNB.n1311 VNB.n1305 0.246
R3307 VNB.n1312 VNB.n1311 0.246
R3308 VNB.n1311 VNB.n1310 0.246
R3309 VNB.n20 VNB.n14 0.246
R3310 VNB.n21 VNB.n20 0.246
R3311 VNB.n20 VNB.n19 0.246
R3312 VNB.n151 VNB.n146 0.246
R3313 VNB.n152 VNB.n151 0.246
R3314 VNB.n151 VNB.n150 0.246
R3315 VNB.n1399 VNB.n1398 0.246
R3316 VNB.n796 VNB 0.204
R3317 VNB.n1385 VNB 0.198
R3318 VNB.n169 VNB.n168 0.136
R3319 VNB.n175 VNB.n169 0.136
R3320 VNB.n186 VNB.n175 0.136
R3321 VNB.n190 VNB.n186 0.136
R3322 VNB.n194 VNB.n190 0.136
R3323 VNB.n220 VNB.n216 0.136
R3324 VNB.n224 VNB.n220 0.136
R3325 VNB.n228 VNB.n224 0.136
R3326 VNB.n234 VNB.n228 0.136
R3327 VNB.n245 VNB.n234 0.136
R3328 VNB.n249 VNB.n245 0.136
R3329 VNB.n253 VNB.n249 0.136
R3330 VNB.n279 VNB.n275 0.136
R3331 VNB.n283 VNB.n279 0.136
R3332 VNB.n287 VNB.n283 0.136
R3333 VNB.n293 VNB.n287 0.136
R3334 VNB.n304 VNB.n293 0.136
R3335 VNB.n308 VNB.n304 0.136
R3336 VNB.n312 VNB.n308 0.136
R3337 VNB.n338 VNB.n334 0.136
R3338 VNB.n342 VNB.n338 0.136
R3339 VNB.n346 VNB.n342 0.136
R3340 VNB.n352 VNB.n346 0.136
R3341 VNB.n363 VNB.n352 0.136
R3342 VNB.n367 VNB.n363 0.136
R3343 VNB.n371 VNB.n367 0.136
R3344 VNB.n397 VNB.n393 0.136
R3345 VNB.n401 VNB.n397 0.136
R3346 VNB.n405 VNB.n401 0.136
R3347 VNB.n409 VNB.n405 0.136
R3348 VNB.n413 VNB.n409 0.136
R3349 VNB.n417 VNB.n413 0.136
R3350 VNB.n421 VNB.n417 0.136
R3351 VNB.n426 VNB.n421 0.136
R3352 VNB.n438 VNB.n426 0.136
R3353 VNB.n442 VNB.n438 0.136
R3354 VNB.n446 VNB.n442 0.136
R3355 VNB.n472 VNB.n468 0.136
R3356 VNB.n476 VNB.n472 0.136
R3357 VNB.n480 VNB.n476 0.136
R3358 VNB.n484 VNB.n480 0.136
R3359 VNB.n488 VNB.n484 0.136
R3360 VNB.n492 VNB.n488 0.136
R3361 VNB.n496 VNB.n492 0.136
R3362 VNB.n500 VNB.n496 0.136
R3363 VNB.n506 VNB.n500 0.136
R3364 VNB.n510 VNB.n506 0.136
R3365 VNB.n514 VNB.n510 0.136
R3366 VNB.n540 VNB.n536 0.136
R3367 VNB.n544 VNB.n540 0.136
R3368 VNB.n548 VNB.n544 0.136
R3369 VNB.n554 VNB.n548 0.136
R3370 VNB.n565 VNB.n554 0.136
R3371 VNB.n569 VNB.n565 0.136
R3372 VNB.n573 VNB.n569 0.136
R3373 VNB.n599 VNB.n595 0.136
R3374 VNB.n603 VNB.n599 0.136
R3375 VNB.n607 VNB.n603 0.136
R3376 VNB.n611 VNB.n607 0.136
R3377 VNB.n615 VNB.n611 0.136
R3378 VNB.n619 VNB.n615 0.136
R3379 VNB.n623 VNB.n619 0.136
R3380 VNB.n628 VNB.n623 0.136
R3381 VNB.n640 VNB.n628 0.136
R3382 VNB.n644 VNB.n640 0.136
R3383 VNB.n648 VNB.n644 0.136
R3384 VNB.n674 VNB.n670 0.136
R3385 VNB.n678 VNB.n674 0.136
R3386 VNB.n682 VNB.n678 0.136
R3387 VNB.n686 VNB.n682 0.136
R3388 VNB.n690 VNB.n686 0.136
R3389 VNB.n694 VNB.n690 0.136
R3390 VNB.n698 VNB.n694 0.136
R3391 VNB.n703 VNB.n698 0.136
R3392 VNB.n715 VNB.n703 0.136
R3393 VNB.n719 VNB.n715 0.136
R3394 VNB.n723 VNB.n719 0.136
R3395 VNB.n749 VNB.n745 0.136
R3396 VNB.n753 VNB.n749 0.136
R3397 VNB.n757 VNB.n753 0.136
R3398 VNB.n761 VNB.n757 0.136
R3399 VNB.n767 VNB.n761 0.136
R3400 VNB.n771 VNB.n767 0.136
R3401 VNB.n775 VNB.n771 0.136
R3402 VNB.n777 VNB.n776 0.136
R3403 VNB.n778 VNB.n777 0.136
R3404 VNB.n779 VNB.n778 0.136
R3405 VNB.n780 VNB.n779 0.136
R3406 VNB.n781 VNB.n780 0.136
R3407 VNB.n782 VNB.n781 0.136
R3408 VNB.n783 VNB.n782 0.136
R3409 VNB.n784 VNB.n783 0.136
R3410 VNB.n785 VNB.n784 0.136
R3411 VNB.n786 VNB.n785 0.136
R3412 VNB.n787 VNB.n786 0.136
R3413 VNB.n800 VNB.n796 0.136
R3414 VNB.n804 VNB.n800 0.136
R3415 VNB.n808 VNB.n804 0.136
R3416 VNB.n812 VNB.n808 0.136
R3417 VNB.n816 VNB.n812 0.136
R3418 VNB.n820 VNB.n816 0.136
R3419 VNB.n824 VNB.n820 0.136
R3420 VNB.n828 VNB.n824 0.136
R3421 VNB.n834 VNB.n828 0.136
R3422 VNB.n838 VNB.n834 0.136
R3423 VNB.n842 VNB.n838 0.136
R3424 VNB.n868 VNB.n864 0.136
R3425 VNB.n872 VNB.n868 0.136
R3426 VNB.n876 VNB.n872 0.136
R3427 VNB.n882 VNB.n876 0.136
R3428 VNB.n893 VNB.n882 0.136
R3429 VNB.n897 VNB.n893 0.136
R3430 VNB.n901 VNB.n897 0.136
R3431 VNB.n927 VNB.n923 0.136
R3432 VNB.n931 VNB.n927 0.136
R3433 VNB.n935 VNB.n931 0.136
R3434 VNB.n939 VNB.n935 0.136
R3435 VNB.n943 VNB.n939 0.136
R3436 VNB.n947 VNB.n943 0.136
R3437 VNB.n951 VNB.n947 0.136
R3438 VNB.n955 VNB.n951 0.136
R3439 VNB.n961 VNB.n955 0.136
R3440 VNB.n965 VNB.n961 0.136
R3441 VNB.n969 VNB.n965 0.136
R3442 VNB.n995 VNB.n991 0.136
R3443 VNB.n999 VNB.n995 0.136
R3444 VNB.n1003 VNB.n999 0.136
R3445 VNB.n1007 VNB.n1003 0.136
R3446 VNB.n1011 VNB.n1007 0.136
R3447 VNB.n1015 VNB.n1011 0.136
R3448 VNB.n1019 VNB.n1015 0.136
R3449 VNB.n1024 VNB.n1019 0.136
R3450 VNB.n1036 VNB.n1024 0.136
R3451 VNB.n1040 VNB.n1036 0.136
R3452 VNB.n1044 VNB.n1040 0.136
R3453 VNB.n1070 VNB.n1066 0.136
R3454 VNB.n1074 VNB.n1070 0.136
R3455 VNB.n1078 VNB.n1074 0.136
R3456 VNB.n1084 VNB.n1078 0.136
R3457 VNB.n1095 VNB.n1084 0.136
R3458 VNB.n1099 VNB.n1095 0.136
R3459 VNB.n1103 VNB.n1099 0.136
R3460 VNB.n1129 VNB.n1125 0.136
R3461 VNB.n1133 VNB.n1129 0.136
R3462 VNB.n1137 VNB.n1133 0.136
R3463 VNB.n1141 VNB.n1137 0.136
R3464 VNB.n1145 VNB.n1141 0.136
R3465 VNB.n1149 VNB.n1145 0.136
R3466 VNB.n1153 VNB.n1149 0.136
R3467 VNB.n1158 VNB.n1153 0.136
R3468 VNB.n1170 VNB.n1158 0.136
R3469 VNB.n1174 VNB.n1170 0.136
R3470 VNB.n1178 VNB.n1174 0.136
R3471 VNB.n1204 VNB.n1200 0.136
R3472 VNB.n1208 VNB.n1204 0.136
R3473 VNB.n1212 VNB.n1208 0.136
R3474 VNB.n1216 VNB.n1212 0.136
R3475 VNB.n1220 VNB.n1216 0.136
R3476 VNB.n1224 VNB.n1220 0.136
R3477 VNB.n1228 VNB.n1224 0.136
R3478 VNB.n1232 VNB.n1228 0.136
R3479 VNB.n1238 VNB.n1232 0.136
R3480 VNB.n1242 VNB.n1238 0.136
R3481 VNB.n1246 VNB.n1242 0.136
R3482 VNB.n1272 VNB.n1268 0.136
R3483 VNB.n1276 VNB.n1272 0.136
R3484 VNB.n1280 VNB.n1276 0.136
R3485 VNB.n1284 VNB.n1280 0.136
R3486 VNB.n1290 VNB.n1284 0.136
R3487 VNB.n1294 VNB.n1290 0.136
R3488 VNB.n1298 VNB.n1294 0.136
R3489 VNB.n1324 VNB.n1320 0.136
R3490 VNB.n1328 VNB.n1324 0.136
R3491 VNB.n1332 VNB.n1328 0.136
R3492 VNB.n1336 VNB.n1332 0.136
R3493 VNB.n1340 VNB.n1336 0.136
R3494 VNB.n1344 VNB.n1340 0.136
R3495 VNB.n1348 VNB.n1344 0.136
R3496 VNB.n1353 VNB.n1348 0.136
R3497 VNB.n1365 VNB.n1353 0.136
R3498 VNB.n1369 VNB.n1365 0.136
R3499 VNB.n1373 VNB.n1369 0.136
R3500 VNB.n1375 VNB.n1374 0.136
R3501 VNB.n1376 VNB.n1375 0.136
R3502 VNB.n1377 VNB.n1376 0.136
R3503 VNB.n1378 VNB.n1377 0.136
R3504 VNB.n1379 VNB.n1378 0.136
R3505 VNB.n1380 VNB.n1379 0.136
R3506 VNB.n1381 VNB.n1380 0.136
R3507 VNB.n1382 VNB.n1381 0.136
R3508 VNB.n1383 VNB.n1382 0.136
R3509 VNB.n1384 VNB.n1383 0.136
R3510 VNB.n1385 VNB.n1384 0.136
R3511 VNB.n787 VNB 0.068
R3512 a_599_943.n6 a_599_943.t7 480.392
R3513 a_599_943.n8 a_599_943.t11 454.685
R3514 a_599_943.n8 a_599_943.t9 428.979
R3515 a_599_943.n6 a_599_943.t10 403.272
R3516 a_599_943.n7 a_599_943.t8 266.974
R3517 a_599_943.n9 a_599_943.t12 221.453
R3518 a_599_943.n13 a_599_943.n11 196.598
R3519 a_599_943.n11 a_599_943.n5 180.846
R3520 a_599_943.n9 a_599_943.n8 108.494
R3521 a_599_943.n7 a_599_943.n6 108.494
R3522 a_599_943.n10 a_599_943.n9 80.035
R3523 a_599_943.n4 a_599_943.n3 79.232
R3524 a_599_943.n10 a_599_943.n7 77.315
R3525 a_599_943.n11 a_599_943.n10 76
R3526 a_599_943.n5 a_599_943.n4 63.152
R3527 a_599_943.n13 a_599_943.n12 30
R3528 a_599_943.n14 a_599_943.n0 24.383
R3529 a_599_943.n14 a_599_943.n13 23.684
R3530 a_599_943.n5 a_599_943.n1 16.08
R3531 a_599_943.n4 a_599_943.n2 16.08
R3532 a_599_943.n1 a_599_943.t1 14.282
R3533 a_599_943.n1 a_599_943.t2 14.282
R3534 a_599_943.n2 a_599_943.t5 14.282
R3535 a_599_943.n2 a_599_943.t6 14.282
R3536 a_599_943.n3 a_599_943.t4 14.282
R3537 a_599_943.n3 a_599_943.t3 14.282
R3538 a_15932_181.n7 a_15932_181.n3 336.934
R3539 a_15932_181.n12 a_15932_181.n11 98.501
R3540 a_15932_181.n14 a_15932_181.n12 96.417
R3541 a_15932_181.n6 a_15932_181.n4 80.526
R3542 a_15932_181.n12 a_15932_181.n7 78.403
R3543 a_15932_181.n3 a_15932_181.n2 75.271
R3544 a_15932_181.n11 a_15932_181.n10 30
R3545 a_15932_181.n6 a_15932_181.n5 30
R3546 a_15932_181.n14 a_15932_181.n13 30
R3547 a_15932_181.n9 a_15932_181.n8 24.383
R3548 a_15932_181.n15 a_15932_181.n0 24.383
R3549 a_15932_181.n11 a_15932_181.n9 23.684
R3550 a_15932_181.n15 a_15932_181.n14 23.684
R3551 a_15932_181.n7 a_15932_181.n6 20.417
R3552 a_15932_181.n1 a_15932_181.t5 14.282
R3553 a_15932_181.n1 a_15932_181.t4 14.282
R3554 a_15932_181.n2 a_15932_181.t1 14.282
R3555 a_15932_181.n2 a_15932_181.t2 14.282
R3556 a_15932_181.n3 a_15932_181.n1 12.119
R3557 a_3643_75.n1 a_3643_75.n0 25.576
R3558 a_3643_75.n3 a_3643_75.n2 9.111
R3559 a_3643_75.n7 a_3643_75.n5 7.859
R3560 a_3643_75.t0 a_3643_75.n7 3.034
R3561 a_3643_75.n5 a_3643_75.n3 1.964
R3562 a_3643_75.n5 a_3643_75.n4 1.964
R3563 a_3643_75.t0 a_3643_75.n1 1.871
R3564 a_3643_75.n7 a_3643_75.n6 0.443
R3565 a_91_75.n4 a_91_75.n3 19.724
R3566 a_91_75.t0 a_91_75.n5 11.595
R3567 a_91_75.t0 a_91_75.n4 9.207
R3568 a_91_75.n2 a_91_75.n0 8.543
R3569 a_91_75.t0 a_91_75.n2 3.034
R3570 a_91_75.n2 a_91_75.n1 0.443
R3571 a_372_182.n8 a_372_182.n6 96.467
R3572 a_372_182.n3 a_372_182.n1 44.628
R3573 a_372_182.t0 a_372_182.n8 32.417
R3574 a_372_182.n3 a_372_182.n2 23.284
R3575 a_372_182.n6 a_372_182.n5 22.349
R3576 a_372_182.t0 a_372_182.n10 20.241
R3577 a_372_182.n10 a_372_182.n9 13.494
R3578 a_372_182.n6 a_372_182.n4 8.443
R3579 a_372_182.t0 a_372_182.n0 8.137
R3580 a_372_182.t0 a_372_182.n3 5.727
R3581 a_372_182.n8 a_372_182.n7 1.435
R3582 a_5271_75.n4 a_5271_75.n3 19.724
R3583 a_5271_75.t0 a_5271_75.n5 11.595
R3584 a_5271_75.t0 a_5271_75.n4 9.207
R3585 a_5271_75.n2 a_5271_75.n0 8.543
R3586 a_5271_75.t0 a_5271_75.n2 3.034
R3587 a_5271_75.n2 a_5271_75.n1 0.443
R3588 a_5552_182.n8 a_5552_182.n6 96.467
R3589 a_5552_182.n3 a_5552_182.n1 44.628
R3590 a_5552_182.t0 a_5552_182.n8 32.417
R3591 a_5552_182.n3 a_5552_182.n2 23.284
R3592 a_5552_182.n6 a_5552_182.n5 22.349
R3593 a_5552_182.t0 a_5552_182.n10 20.241
R3594 a_5552_182.n10 a_5552_182.n9 13.494
R3595 a_5552_182.n6 a_5552_182.n4 8.443
R3596 a_5552_182.t0 a_5552_182.n0 8.137
R3597 a_5552_182.t0 a_5552_182.n3 5.727
R3598 a_5552_182.n8 a_5552_182.n7 1.435
R3599 a_16318_73.n2 a_16318_73.n0 34.602
R3600 a_16318_73.n2 a_16318_73.n1 2.138
R3601 a_16318_73.t0 a_16318_73.n2 0.069
R3602 a_2141_1004.n4 a_2141_1004.t6 512.525
R3603 a_2141_1004.n4 a_2141_1004.t7 371.139
R3604 a_2141_1004.n5 a_2141_1004.t5 271.162
R3605 a_2141_1004.n8 a_2141_1004.n6 194.086
R3606 a_2141_1004.n5 a_2141_1004.n4 172.76
R3607 a_2141_1004.n6 a_2141_1004.n3 162.547
R3608 a_2141_1004.n6 a_2141_1004.n5 153.315
R3609 a_2141_1004.n3 a_2141_1004.n2 76.002
R3610 a_2141_1004.n8 a_2141_1004.n7 30
R3611 a_2141_1004.n9 a_2141_1004.n0 24.383
R3612 a_2141_1004.n9 a_2141_1004.n8 23.684
R3613 a_2141_1004.n1 a_2141_1004.t1 14.282
R3614 a_2141_1004.n1 a_2141_1004.t0 14.282
R3615 a_2141_1004.n2 a_2141_1004.t4 14.282
R3616 a_2141_1004.n2 a_2141_1004.t3 14.282
R3617 a_2141_1004.n3 a_2141_1004.n1 12.85
R3618 a_9009_1004.n6 a_9009_1004.t8 480.392
R3619 a_9009_1004.n6 a_9009_1004.t7 403.272
R3620 a_9009_1004.n7 a_9009_1004.t9 293.527
R3621 a_9009_1004.n10 a_9009_1004.n8 223.151
R3622 a_9009_1004.n8 a_9009_1004.n5 154.293
R3623 a_9009_1004.n8 a_9009_1004.n7 153.315
R3624 a_9009_1004.n7 a_9009_1004.n6 81.941
R3625 a_9009_1004.n4 a_9009_1004.n3 79.232
R3626 a_9009_1004.n5 a_9009_1004.n4 63.152
R3627 a_9009_1004.n10 a_9009_1004.n9 30
R3628 a_9009_1004.n11 a_9009_1004.n0 24.383
R3629 a_9009_1004.n11 a_9009_1004.n10 23.684
R3630 a_9009_1004.n5 a_9009_1004.n1 16.08
R3631 a_9009_1004.n4 a_9009_1004.n2 16.08
R3632 a_9009_1004.n1 a_9009_1004.t1 14.282
R3633 a_9009_1004.n1 a_9009_1004.t0 14.282
R3634 a_9009_1004.n2 a_9009_1004.t4 14.282
R3635 a_9009_1004.n2 a_9009_1004.t3 14.282
R3636 a_9009_1004.n3 a_9009_1004.t6 14.282
R3637 a_9009_1004.n3 a_9009_1004.t5 14.282
R3638 a_4626_73.t0 a_4626_73.n1 34.62
R3639 a_4626_73.t0 a_4626_73.n0 8.137
R3640 a_4626_73.t0 a_4626_73.n2 4.69
R3641 a_2036_73.t0 a_2036_73.n1 34.62
R3642 a_2036_73.t0 a_2036_73.n0 8.137
R3643 a_2036_73.t0 a_2036_73.n2 4.69
R3644 a_14003_75.n5 a_14003_75.n4 19.724
R3645 a_14003_75.t0 a_14003_75.n3 11.595
R3646 a_14003_75.t0 a_14003_75.n5 9.207
R3647 a_14003_75.n2 a_14003_75.n1 2.455
R3648 a_14003_75.n2 a_14003_75.n0 1.32
R3649 a_14003_75.t0 a_14003_75.n2 0.246
R3650 a_2681_75.n4 a_2681_75.n3 19.724
R3651 a_2681_75.t0 a_2681_75.n5 11.595
R3652 a_2681_75.t0 a_2681_75.n4 9.207
R3653 a_2681_75.n2 a_2681_75.n0 8.543
R3654 a_2681_75.t0 a_2681_75.n2 3.034
R3655 a_2681_75.n2 a_2681_75.n1 0.443
R3656 a_1334_182.n9 a_1334_182.n7 82.852
R3657 a_1334_182.n3 a_1334_182.n1 44.628
R3658 a_1334_182.t0 a_1334_182.n9 32.417
R3659 a_1334_182.n7 a_1334_182.n6 27.2
R3660 a_1334_182.n5 a_1334_182.n4 23.498
R3661 a_1334_182.n3 a_1334_182.n2 23.284
R3662 a_1334_182.n7 a_1334_182.n5 22.4
R3663 a_1334_182.t0 a_1334_182.n11 20.241
R3664 a_1334_182.n11 a_1334_182.n10 13.494
R3665 a_1334_182.t0 a_1334_182.n0 8.137
R3666 a_1334_182.t0 a_1334_182.n3 5.727
R3667 a_1334_182.n9 a_1334_182.n8 1.435
R3668 a_10732_182.n9 a_10732_182.n7 82.852
R3669 a_10732_182.n3 a_10732_182.n1 44.628
R3670 a_10732_182.t0 a_10732_182.n9 32.417
R3671 a_10732_182.n7 a_10732_182.n6 27.2
R3672 a_10732_182.n5 a_10732_182.n4 23.498
R3673 a_10732_182.n3 a_10732_182.n2 23.284
R3674 a_10732_182.n7 a_10732_182.n5 22.4
R3675 a_10732_182.t0 a_10732_182.n11 20.241
R3676 a_10732_182.n11 a_10732_182.n10 13.494
R3677 a_10732_182.t0 a_10732_182.n0 8.137
R3678 a_10732_182.t0 a_10732_182.n3 5.727
R3679 a_10732_182.n9 a_10732_182.n8 1.435
R3680 a_13322_182.n8 a_13322_182.n6 96.467
R3681 a_13322_182.n3 a_13322_182.n1 44.628
R3682 a_13322_182.t0 a_13322_182.n8 32.417
R3683 a_13322_182.n3 a_13322_182.n2 23.284
R3684 a_13322_182.n6 a_13322_182.n5 22.349
R3685 a_13322_182.t0 a_13322_182.n10 20.241
R3686 a_13322_182.n10 a_13322_182.n9 13.494
R3687 a_13322_182.n6 a_13322_182.n4 8.443
R3688 a_13322_182.t0 a_13322_182.n0 8.137
R3689 a_13322_182.t0 a_13322_182.n3 5.727
R3690 a_13322_182.n8 a_13322_182.n7 1.435
R3691 a_3924_182.n10 a_3924_182.n8 82.852
R3692 a_3924_182.n11 a_3924_182.n0 49.6
R3693 a_3924_182.n7 a_3924_182.n6 32.833
R3694 a_3924_182.n8 a_3924_182.t1 32.416
R3695 a_3924_182.n10 a_3924_182.n9 27.2
R3696 a_3924_182.n3 a_3924_182.n2 23.284
R3697 a_3924_182.n11 a_3924_182.n10 22.4
R3698 a_3924_182.n7 a_3924_182.n4 19.017
R3699 a_3924_182.n6 a_3924_182.n5 13.494
R3700 a_3924_182.t1 a_3924_182.n1 7.04
R3701 a_3924_182.t1 a_3924_182.n3 5.727
R3702 a_3924_182.n8 a_3924_182.n7 1.435
R3703 a_7216_73.t0 a_7216_73.n1 34.62
R3704 a_7216_73.t0 a_7216_73.n0 8.137
R3705 a_7216_73.t0 a_7216_73.n2 4.69
R3706 a_7321_1004.n3 a_7321_1004.t5 512.525
R3707 a_7321_1004.n3 a_7321_1004.t6 371.139
R3708 a_7321_1004.n4 a_7321_1004.t7 271.162
R3709 a_7321_1004.n7 a_7321_1004.n5 200.608
R3710 a_7321_1004.n4 a_7321_1004.n3 172.76
R3711 a_7321_1004.n5 a_7321_1004.n2 162.547
R3712 a_7321_1004.n5 a_7321_1004.n4 153.315
R3713 a_7321_1004.n2 a_7321_1004.n1 76.002
R3714 a_7321_1004.n7 a_7321_1004.n6 15.218
R3715 a_7321_1004.n0 a_7321_1004.t0 14.282
R3716 a_7321_1004.n0 a_7321_1004.t1 14.282
R3717 a_7321_1004.n1 a_7321_1004.t3 14.282
R3718 a_7321_1004.n1 a_7321_1004.t4 14.282
R3719 a_7321_1004.n2 a_7321_1004.n0 12.85
R3720 a_7321_1004.n8 a_7321_1004.n7 12.014
R3721 a_15652_73.n13 a_15652_73.n12 26.811
R3722 a_15652_73.n6 a_15652_73.n5 24.977
R3723 a_15652_73.n2 a_15652_73.n1 24.877
R3724 a_15652_73.t0 a_15652_73.n2 12.677
R3725 a_15652_73.t0 a_15652_73.n3 11.595
R3726 a_15652_73.n11 a_15652_73.n10 8.561
R3727 a_15652_73.t0 a_15652_73.n4 7.273
R3728 a_15652_73.n9 a_15652_73.n8 7.066
R3729 a_15652_73.t0 a_15652_73.n0 6.109
R3730 a_15652_73.t1 a_15652_73.n7 4.864
R3731 a_15652_73.t0 a_15652_73.n13 2.074
R3732 a_15652_73.n7 a_15652_73.n6 1.13
R3733 a_15652_73.t1 a_15652_73.n11 0.958
R3734 a_15652_73.n13 a_15652_73.t1 0.937
R3735 a_15652_73.t1 a_15652_73.n9 0.86
R3736 a_14986_73.t0 a_14986_73.n1 34.62
R3737 a_14986_73.t0 a_14986_73.n0 8.137
R3738 a_14986_73.t0 a_14986_73.n2 4.69
R3739 a_11694_182.n9 a_11694_182.n7 82.852
R3740 a_11694_182.n3 a_11694_182.n1 44.628
R3741 a_11694_182.t0 a_11694_182.n9 32.417
R3742 a_11694_182.n7 a_11694_182.n6 27.2
R3743 a_11694_182.n5 a_11694_182.n4 23.498
R3744 a_11694_182.n3 a_11694_182.n2 23.284
R3745 a_11694_182.n7 a_11694_182.n5 22.4
R3746 a_11694_182.t0 a_11694_182.n11 20.241
R3747 a_11694_182.n11 a_11694_182.n10 13.494
R3748 a_11694_182.t0 a_11694_182.n0 8.137
R3749 a_11694_182.t0 a_11694_182.n3 5.727
R3750 a_11694_182.n9 a_11694_182.n8 1.435
R3751 a_9104_182.n9 a_9104_182.n7 82.852
R3752 a_9104_182.n3 a_9104_182.n1 44.628
R3753 a_9104_182.t0 a_9104_182.n9 32.417
R3754 a_9104_182.n7 a_9104_182.n6 27.2
R3755 a_9104_182.n5 a_9104_182.n4 23.498
R3756 a_9104_182.n3 a_9104_182.n2 23.284
R3757 a_9104_182.n7 a_9104_182.n5 22.4
R3758 a_9104_182.t0 a_9104_182.n11 20.241
R3759 a_9104_182.n11 a_9104_182.n10 13.494
R3760 a_9104_182.t0 a_9104_182.n0 8.137
R3761 a_9104_182.t0 a_9104_182.n3 5.727
R3762 a_9104_182.n9 a_9104_182.n8 1.435
R3763 a_1053_75.n5 a_1053_75.n4 19.724
R3764 a_1053_75.t0 a_1053_75.n3 11.595
R3765 a_1053_75.t0 a_1053_75.n5 9.207
R3766 a_1053_75.n2 a_1053_75.n1 2.455
R3767 a_1053_75.n2 a_1053_75.n0 1.32
R3768 a_1053_75.t0 a_1053_75.n2 0.246
R3769 a_2962_182.n8 a_2962_182.n6 96.467
R3770 a_2962_182.n3 a_2962_182.n1 44.628
R3771 a_2962_182.t0 a_2962_182.n8 32.417
R3772 a_2962_182.n3 a_2962_182.n2 23.284
R3773 a_2962_182.n6 a_2962_182.n5 22.349
R3774 a_2962_182.t0 a_2962_182.n10 20.241
R3775 a_2962_182.n10 a_2962_182.n9 13.494
R3776 a_2962_182.n6 a_2962_182.n4 8.443
R3777 a_2962_182.t0 a_2962_182.n0 8.137
R3778 a_2962_182.t0 a_2962_182.n3 5.727
R3779 a_2962_182.n8 a_2962_182.n7 1.435
R3780 a_16984_73.t0 a_16984_73.n1 34.62
R3781 a_16984_73.t0 a_16984_73.n0 8.137
R3782 a_16984_73.t0 a_16984_73.n2 4.69
R3783 a_11413_75.n5 a_11413_75.n4 19.724
R3784 a_11413_75.t0 a_11413_75.n3 11.595
R3785 a_11413_75.t0 a_11413_75.n5 9.207
R3786 a_11413_75.n2 a_11413_75.n1 2.455
R3787 a_11413_75.n2 a_11413_75.n0 1.32
R3788 a_11413_75.t0 a_11413_75.n2 0.246
R3789 a_8142_182.n9 a_8142_182.n7 82.852
R3790 a_8142_182.n3 a_8142_182.n1 44.628
R3791 a_8142_182.t0 a_8142_182.n9 32.417
R3792 a_8142_182.n7 a_8142_182.n6 27.2
R3793 a_8142_182.n5 a_8142_182.n4 23.498
R3794 a_8142_182.n3 a_8142_182.n2 23.284
R3795 a_8142_182.n7 a_8142_182.n5 22.4
R3796 a_8142_182.t0 a_8142_182.n11 20.241
R3797 a_8142_182.n11 a_8142_182.n10 13.494
R3798 a_8142_182.t0 a_8142_182.n0 8.137
R3799 a_8142_182.t0 a_8142_182.n3 5.727
R3800 a_8142_182.n9 a_8142_182.n8 1.435
R3801 a_12396_73.n12 a_12396_73.n11 26.811
R3802 a_12396_73.n6 a_12396_73.n5 24.977
R3803 a_12396_73.n2 a_12396_73.n1 24.877
R3804 a_12396_73.t0 a_12396_73.n2 12.677
R3805 a_12396_73.t0 a_12396_73.n3 11.595
R3806 a_12396_73.t1 a_12396_73.n8 8.137
R3807 a_12396_73.t0 a_12396_73.n4 7.273
R3808 a_12396_73.t0 a_12396_73.n0 6.109
R3809 a_12396_73.t1 a_12396_73.n7 4.864
R3810 a_12396_73.t0 a_12396_73.n12 2.074
R3811 a_12396_73.n7 a_12396_73.n6 1.13
R3812 a_12396_73.n12 a_12396_73.t1 0.937
R3813 a_12396_73.t1 a_12396_73.n10 0.804
R3814 a_12396_73.n10 a_12396_73.n9 0.136
R3815 a_10451_75.n5 a_10451_75.n4 19.724
R3816 a_10451_75.t0 a_10451_75.n3 11.595
R3817 a_10451_75.t0 a_10451_75.n5 9.207
R3818 a_10451_75.n2 a_10451_75.n1 2.455
R3819 a_10451_75.n2 a_10451_75.n0 1.32
R3820 a_10451_75.t0 a_10451_75.n2 0.246
R3821 a_8823_75.n1 a_8823_75.n0 25.576
R3822 a_8823_75.n3 a_8823_75.n2 9.111
R3823 a_8823_75.n7 a_8823_75.n6 2.455
R3824 a_8823_75.n5 a_8823_75.n3 1.964
R3825 a_8823_75.n5 a_8823_75.n4 1.964
R3826 a_8823_75.t0 a_8823_75.n1 1.871
R3827 a_8823_75.n7 a_8823_75.n5 0.636
R3828 a_8823_75.t0 a_8823_75.n7 0.246
R3829 a_7861_75.n5 a_7861_75.n4 19.724
R3830 a_7861_75.t0 a_7861_75.n3 11.595
R3831 a_7861_75.t0 a_7861_75.n5 9.207
R3832 a_7861_75.n2 a_7861_75.n1 2.455
R3833 a_7861_75.n2 a_7861_75.n0 1.32
R3834 a_7861_75.t0 a_7861_75.n2 0.246
C6 VPB VNB 65.08fF
C7 a_7861_75.n0 VNB 0.10fF
C8 a_7861_75.n1 VNB 0.04fF
C9 a_7861_75.n2 VNB 0.03fF
C10 a_7861_75.n3 VNB 0.07fF
C11 a_7861_75.n4 VNB 0.08fF
C12 a_7861_75.n5 VNB 0.06fF
C13 a_8823_75.n0 VNB 0.09fF
C14 a_8823_75.n1 VNB 0.10fF
C15 a_8823_75.n2 VNB 0.05fF
C16 a_8823_75.n3 VNB 0.03fF
C17 a_8823_75.n4 VNB 0.04fF
C18 a_8823_75.n5 VNB 0.03fF
C19 a_8823_75.n6 VNB 0.04fF
C20 a_10451_75.n0 VNB 0.10fF
C21 a_10451_75.n1 VNB 0.04fF
C22 a_10451_75.n2 VNB 0.03fF
C23 a_10451_75.n3 VNB 0.07fF
C24 a_10451_75.n4 VNB 0.08fF
C25 a_10451_75.n5 VNB 0.06fF
C26 a_12396_73.n0 VNB 0.02fF
C27 a_12396_73.n1 VNB 0.10fF
C28 a_12396_73.n2 VNB 0.06fF
C29 a_12396_73.n3 VNB 0.06fF
C30 a_12396_73.n4 VNB 0.00fF
C31 a_12396_73.n5 VNB 0.04fF
C32 a_12396_73.n6 VNB 0.05fF
C33 a_12396_73.n7 VNB 0.02fF
C34 a_12396_73.n8 VNB 0.05fF
C35 a_12396_73.n9 VNB 0.08fF
C36 a_12396_73.n10 VNB 0.17fF
C37 a_12396_73.t1 VNB 0.23fF
C38 a_12396_73.n11 VNB 0.09fF
C39 a_12396_73.n12 VNB 0.00fF
C40 a_8142_182.n0 VNB 0.07fF
C41 a_8142_182.n1 VNB 0.09fF
C42 a_8142_182.n2 VNB 0.13fF
C43 a_8142_182.n3 VNB 0.11fF
C44 a_8142_182.n4 VNB 0.02fF
C45 a_8142_182.n5 VNB 0.03fF
C46 a_8142_182.n6 VNB 0.02fF
C47 a_8142_182.n7 VNB 0.05fF
C48 a_8142_182.n8 VNB 0.03fF
C49 a_8142_182.n9 VNB 0.11fF
C50 a_8142_182.n10 VNB 0.06fF
C51 a_8142_182.n11 VNB 0.01fF
C52 a_8142_182.t0 VNB 0.33fF
C53 a_11413_75.n0 VNB 0.10fF
C54 a_11413_75.n1 VNB 0.04fF
C55 a_11413_75.n2 VNB 0.03fF
C56 a_11413_75.n3 VNB 0.07fF
C57 a_11413_75.n4 VNB 0.08fF
C58 a_11413_75.n5 VNB 0.06fF
C59 a_16984_73.n0 VNB 0.06fF
C60 a_16984_73.n1 VNB 0.13fF
C61 a_16984_73.n2 VNB 0.04fF
C62 a_2962_182.n0 VNB 0.07fF
C63 a_2962_182.n1 VNB 0.09fF
C64 a_2962_182.n2 VNB 0.13fF
C65 a_2962_182.n3 VNB 0.11fF
C66 a_2962_182.n4 VNB 0.02fF
C67 a_2962_182.n5 VNB 0.03fF
C68 a_2962_182.n6 VNB 0.06fF
C69 a_2962_182.n7 VNB 0.03fF
C70 a_2962_182.n8 VNB 0.12fF
C71 a_2962_182.n9 VNB 0.06fF
C72 a_2962_182.n10 VNB 0.01fF
C73 a_2962_182.t0 VNB 0.33fF
C74 a_1053_75.n0 VNB 0.10fF
C75 a_1053_75.n1 VNB 0.04fF
C76 a_1053_75.n2 VNB 0.03fF
C77 a_1053_75.n3 VNB 0.07fF
C78 a_1053_75.n4 VNB 0.08fF
C79 a_1053_75.n5 VNB 0.06fF
C80 a_9104_182.n0 VNB 0.07fF
C81 a_9104_182.n1 VNB 0.09fF
C82 a_9104_182.n2 VNB 0.13fF
C83 a_9104_182.n3 VNB 0.11fF
C84 a_9104_182.n4 VNB 0.02fF
C85 a_9104_182.n5 VNB 0.03fF
C86 a_9104_182.n6 VNB 0.02fF
C87 a_9104_182.n7 VNB 0.05fF
C88 a_9104_182.n8 VNB 0.03fF
C89 a_9104_182.n9 VNB 0.11fF
C90 a_9104_182.n10 VNB 0.06fF
C91 a_9104_182.n11 VNB 0.01fF
C92 a_9104_182.t0 VNB 0.33fF
C93 a_11694_182.n0 VNB 0.07fF
C94 a_11694_182.n1 VNB 0.09fF
C95 a_11694_182.n2 VNB 0.13fF
C96 a_11694_182.n3 VNB 0.11fF
C97 a_11694_182.n4 VNB 0.02fF
C98 a_11694_182.n5 VNB 0.03fF
C99 a_11694_182.n6 VNB 0.02fF
C100 a_11694_182.n7 VNB 0.05fF
C101 a_11694_182.n8 VNB 0.03fF
C102 a_11694_182.n9 VNB 0.11fF
C103 a_11694_182.n10 VNB 0.06fF
C104 a_11694_182.n11 VNB 0.01fF
C105 a_11694_182.t0 VNB 0.33fF
C106 a_14986_73.n0 VNB 0.05fF
C107 a_14986_73.n1 VNB 0.12fF
C108 a_14986_73.n2 VNB 0.04fF
C109 a_15652_73.n0 VNB 0.02fF
C110 a_15652_73.n1 VNB 0.09fF
C111 a_15652_73.n2 VNB 0.05fF
C112 a_15652_73.n3 VNB 0.06fF
C113 a_15652_73.n4 VNB 0.00fF
C114 a_15652_73.n5 VNB 0.04fF
C115 a_15652_73.n6 VNB 0.05fF
C116 a_15652_73.n7 VNB 0.02fF
C117 a_15652_73.n8 VNB 0.05fF
C118 a_15652_73.n9 VNB 0.09fF
C119 a_15652_73.n10 VNB 0.21fF
C120 a_15652_73.n11 VNB 0.07fF
C121 a_15652_73.t1 VNB 0.14fF
C122 a_15652_73.n12 VNB 0.04fF
C123 a_15652_73.n13 VNB 0.00fF
C124 a_7321_1004.n0 VNB 0.61fF
C125 a_7321_1004.n1 VNB 0.72fF
C126 a_7321_1004.n2 VNB 0.36fF
C127 a_7321_1004.n3 VNB 0.40fF
C128 a_7321_1004.n4 VNB 0.74fF
C129 a_7321_1004.n5 VNB 0.69fF
C130 a_7321_1004.n6 VNB 0.10fF
C131 a_7321_1004.n7 VNB 0.31fF
C132 a_7321_1004.n8 VNB 0.05fF
C133 a_7216_73.n0 VNB 0.05fF
C134 a_7216_73.n1 VNB 0.12fF
C135 a_7216_73.n2 VNB 0.04fF
C136 a_3924_182.n0 VNB 0.02fF
C137 a_3924_182.n1 VNB 0.09fF
C138 a_3924_182.n2 VNB 0.13fF
C139 a_3924_182.n3 VNB 0.11fF
C140 a_3924_182.t1 VNB 0.30fF
C141 a_3924_182.n4 VNB 0.09fF
C142 a_3924_182.n5 VNB 0.06fF
C143 a_3924_182.n6 VNB 0.01fF
C144 a_3924_182.n7 VNB 0.03fF
C145 a_3924_182.n8 VNB 0.11fF
C146 a_3924_182.n9 VNB 0.02fF
C147 a_3924_182.n10 VNB 0.05fF
C148 a_3924_182.n11 VNB 0.02fF
C149 a_13322_182.n0 VNB 0.07fF
C150 a_13322_182.n1 VNB 0.09fF
C151 a_13322_182.n2 VNB 0.13fF
C152 a_13322_182.n3 VNB 0.11fF
C153 a_13322_182.n4 VNB 0.02fF
C154 a_13322_182.n5 VNB 0.03fF
C155 a_13322_182.n6 VNB 0.06fF
C156 a_13322_182.n7 VNB 0.03fF
C157 a_13322_182.n8 VNB 0.12fF
C158 a_13322_182.n9 VNB 0.06fF
C159 a_13322_182.n10 VNB 0.01fF
C160 a_13322_182.t0 VNB 0.33fF
C161 a_10732_182.n0 VNB 0.07fF
C162 a_10732_182.n1 VNB 0.09fF
C163 a_10732_182.n2 VNB 0.13fF
C164 a_10732_182.n3 VNB 0.11fF
C165 a_10732_182.n4 VNB 0.02fF
C166 a_10732_182.n5 VNB 0.03fF
C167 a_10732_182.n6 VNB 0.02fF
C168 a_10732_182.n7 VNB 0.05fF
C169 a_10732_182.n8 VNB 0.03fF
C170 a_10732_182.n9 VNB 0.11fF
C171 a_10732_182.n10 VNB 0.06fF
C172 a_10732_182.n11 VNB 0.01fF
C173 a_10732_182.t0 VNB 0.33fF
C174 a_1334_182.n0 VNB 0.07fF
C175 a_1334_182.n1 VNB 0.09fF
C176 a_1334_182.n2 VNB 0.13fF
C177 a_1334_182.n3 VNB 0.11fF
C178 a_1334_182.n4 VNB 0.02fF
C179 a_1334_182.n5 VNB 0.03fF
C180 a_1334_182.n6 VNB 0.02fF
C181 a_1334_182.n7 VNB 0.05fF
C182 a_1334_182.n8 VNB 0.03fF
C183 a_1334_182.n9 VNB 0.11fF
C184 a_1334_182.n10 VNB 0.06fF
C185 a_1334_182.n11 VNB 0.01fF
C186 a_1334_182.t0 VNB 0.33fF
C187 a_2681_75.n0 VNB 0.20fF
C188 a_2681_75.n1 VNB 0.04fF
C189 a_2681_75.n2 VNB 0.01fF
C190 a_2681_75.n3 VNB 0.08fF
C191 a_2681_75.n4 VNB 0.06fF
C192 a_2681_75.n5 VNB 0.07fF
C193 a_14003_75.n0 VNB 0.10fF
C194 a_14003_75.n1 VNB 0.04fF
C195 a_14003_75.n2 VNB 0.03fF
C196 a_14003_75.n3 VNB 0.07fF
C197 a_14003_75.n4 VNB 0.08fF
C198 a_14003_75.n5 VNB 0.06fF
C199 a_2036_73.n0 VNB 0.05fF
C200 a_2036_73.n1 VNB 0.12fF
C201 a_2036_73.n2 VNB 0.04fF
C202 a_4626_73.n0 VNB 0.05fF
C203 a_4626_73.n1 VNB 0.12fF
C204 a_4626_73.n2 VNB 0.04fF
C205 a_9009_1004.n0 VNB 0.04fF
C206 a_9009_1004.n1 VNB 0.56fF
C207 a_9009_1004.n2 VNB 0.56fF
C208 a_9009_1004.n3 VNB 0.66fF
C209 a_9009_1004.n4 VNB 0.21fF
C210 a_9009_1004.n5 VNB 0.30fF
C211 a_9009_1004.n6 VNB 0.37fF
C212 a_9009_1004.n7 VNB 0.59fF
C213 a_9009_1004.n8 VNB 0.65fF
C214 a_9009_1004.n9 VNB 0.04fF
C215 a_9009_1004.n10 VNB 0.33fF
C216 a_9009_1004.n11 VNB 0.06fF
C217 a_2141_1004.n0 VNB 0.04fF
C218 a_2141_1004.n1 VNB 0.55fF
C219 a_2141_1004.n2 VNB 0.65fF
C220 a_2141_1004.n3 VNB 0.33fF
C221 a_2141_1004.n4 VNB 0.36fF
C222 a_2141_1004.n5 VNB 0.67fF
C223 a_2141_1004.n6 VNB 0.62fF
C224 a_2141_1004.n7 VNB 0.04fF
C225 a_2141_1004.n8 VNB 0.29fF
C226 a_2141_1004.n9 VNB 0.06fF
C227 a_16318_73.n0 VNB 0.13fF
C228 a_16318_73.n1 VNB 0.13fF
C229 a_16318_73.n2 VNB 0.14fF
C230 a_5552_182.n0 VNB 0.07fF
C231 a_5552_182.n1 VNB 0.09fF
C232 a_5552_182.n2 VNB 0.13fF
C233 a_5552_182.n3 VNB 0.11fF
C234 a_5552_182.n4 VNB 0.02fF
C235 a_5552_182.n5 VNB 0.03fF
C236 a_5552_182.n6 VNB 0.06fF
C237 a_5552_182.n7 VNB 0.03fF
C238 a_5552_182.n8 VNB 0.12fF
C239 a_5552_182.n9 VNB 0.06fF
C240 a_5552_182.n10 VNB 0.01fF
C241 a_5552_182.t0 VNB 0.33fF
C242 a_5271_75.n0 VNB 0.20fF
C243 a_5271_75.n1 VNB 0.04fF
C244 a_5271_75.n2 VNB 0.01fF
C245 a_5271_75.n3 VNB 0.08fF
C246 a_5271_75.n4 VNB 0.06fF
C247 a_5271_75.n5 VNB 0.07fF
C248 a_372_182.n0 VNB 0.07fF
C249 a_372_182.n1 VNB 0.09fF
C250 a_372_182.n2 VNB 0.13fF
C251 a_372_182.n3 VNB 0.11fF
C252 a_372_182.n4 VNB 0.02fF
C253 a_372_182.n5 VNB 0.03fF
C254 a_372_182.n6 VNB 0.06fF
C255 a_372_182.n7 VNB 0.03fF
C256 a_372_182.n8 VNB 0.12fF
C257 a_372_182.n9 VNB 0.06fF
C258 a_372_182.n10 VNB 0.01fF
C259 a_372_182.t0 VNB 0.33fF
C260 a_91_75.n0 VNB 0.19fF
C261 a_91_75.n1 VNB 0.04fF
C262 a_91_75.n2 VNB 0.01fF
C263 a_91_75.n3 VNB 0.08fF
C264 a_91_75.n4 VNB 0.06fF
C265 a_91_75.n5 VNB 0.06fF
C266 a_3643_75.n0 VNB 0.09fF
C267 a_3643_75.n1 VNB 0.10fF
C268 a_3643_75.n2 VNB 0.05fF
C269 a_3643_75.n3 VNB 0.03fF
C270 a_3643_75.n4 VNB 0.04fF
C271 a_3643_75.n5 VNB 0.11fF
C272 a_3643_75.n6 VNB 0.04fF
C273 a_15932_181.n0 VNB 0.04fF
C274 a_15932_181.n1 VNB 0.42fF
C275 a_15932_181.n2 VNB 0.51fF
C276 a_15932_181.n3 VNB 0.48fF
C277 a_15932_181.n4 VNB 0.06fF
C278 a_15932_181.n5 VNB 0.03fF
C279 a_15932_181.n6 VNB 0.08fF
C280 a_15932_181.n7 VNB 0.41fF
C281 a_15932_181.n8 VNB 0.04fF
C282 a_15932_181.n9 VNB 0.05fF
C283 a_15932_181.n10 VNB 0.03fF
C284 a_15932_181.n11 VNB 0.10fF
C285 a_15932_181.n12 VNB 1.08fF
C286 a_15932_181.n13 VNB 0.03fF
C287 a_15932_181.n14 VNB 0.09fF
C288 a_15932_181.n15 VNB 0.05fF
C289 a_599_943.n0 VNB 0.04fF
C290 a_599_943.n1 VNB 0.59fF
C291 a_599_943.n2 VNB 0.59fF
C292 a_599_943.n3 VNB 0.69fF
C293 a_599_943.n4 VNB 0.22fF
C294 a_599_943.n5 VNB 0.35fF
C295 a_599_943.n6 VNB 0.43fF
C296 a_599_943.n7 VNB 0.42fF
C297 a_599_943.n8 VNB 0.43fF
C298 a_599_943.t12 VNB 0.57fF
C299 a_599_943.n9 VNB 0.42fF
C300 a_599_943.n10 VNB 1.37fF
C301 a_599_943.n11 VNB 0.49fF
C302 a_599_943.n12 VNB 0.04fF
C303 a_599_943.n13 VNB 0.31fF
C304 a_599_943.n14 VNB 0.06fF
C305 a_13041_75.n0 VNB 0.20fF
C306 a_13041_75.n1 VNB 0.04fF
C307 a_13041_75.n2 VNB 0.01fF
C308 a_13041_75.n3 VNB 0.03fF
C309 a_13041_75.n4 VNB 0.05fF
C310 a_13041_75.n5 VNB 0.09fF
C311 a_13041_75.n6 VNB 0.07fF
C312 a_14284_182.n0 VNB 0.02fF
C313 a_14284_182.n1 VNB 0.09fF
C314 a_14284_182.n2 VNB 0.13fF
C315 a_14284_182.n3 VNB 0.11fF
C316 a_14284_182.t1 VNB 0.30fF
C317 a_14284_182.n4 VNB 0.09fF
C318 a_14284_182.n5 VNB 0.06fF
C319 a_14284_182.n6 VNB 0.01fF
C320 a_14284_182.n7 VNB 0.03fF
C321 a_14284_182.n8 VNB 0.11fF
C322 a_14284_182.n9 VNB 0.02fF
C323 a_14284_182.n10 VNB 0.05fF
C324 a_14284_182.n11 VNB 0.03fF
C325 a_10637_1004.n0 VNB 0.07fF
C326 a_10637_1004.n1 VNB 0.91fF
C327 a_10637_1004.n2 VNB 0.91fF
C328 a_10637_1004.n3 VNB 1.07fF
C329 a_10637_1004.n4 VNB 0.34fF
C330 a_10637_1004.n5 VNB 0.49fF
C331 a_10637_1004.n6 VNB 0.54fF
C332 a_10637_1004.n7 VNB 1.00fF
C333 a_10637_1004.n8 VNB 0.54fF
C334 a_10637_1004.n9 VNB 0.80fF
C335 a_10637_1004.n10 VNB 4.00fF
C336 a_10637_1004.n11 VNB 0.76fF
C337 a_10637_1004.n12 VNB 0.06fF
C338 a_10637_1004.n13 VNB 0.53fF
C339 a_10637_1004.n14 VNB 0.09fF
C340 a_15757_1005.n0 VNB 0.36fF
C341 a_15757_1005.n1 VNB 0.32fF
C342 a_15757_1005.n2 VNB 0.23fF
C343 a_15757_1005.n3 VNB 0.62fF
C344 a_15757_1005.n4 VNB 0.28fF
C345 a_15757_1005.n5 VNB 0.40fF
C346 a_16421_1005.n0 VNB 0.28fF
C347 a_16421_1005.n1 VNB 0.29fF
C348 a_16421_1005.n2 VNB 0.20fF
C349 a_16421_1005.n3 VNB 0.56fF
C350 a_16421_1005.n4 VNB 0.25fF
C351 a_16421_1005.n5 VNB 0.35fF
C352 a_4151_943.n0 VNB 1.21fF
C353 a_4151_943.n1 VNB 0.90fF
C354 a_4151_943.n2 VNB 1.06fF
C355 a_4151_943.n3 VNB 1.32fF
C356 a_4151_943.t6 VNB 1.00fF
C357 a_4151_943.n4 VNB 0.79fF
C358 a_4151_943.n5 VNB 4.66fF
C359 a_4151_943.n6 VNB 0.96fF
C360 a_4151_943.t12 VNB 1.12fF
C361 a_4151_943.n7 VNB 0.83fF
C362 a_4151_943.n8 VNB 19.51fF
C363 a_4151_943.n9 VNB 0.09fF
C364 a_4151_943.n10 VNB 0.12fF
C365 a_4151_943.n11 VNB 0.08fF
C366 a_4151_943.n12 VNB 0.57fF
C367 a_4151_943.n13 VNB 0.96fF
C368 a_4151_943.n14 VNB 0.80fF
C369 a_4151_943.n15 VNB 1.44fF
C370 a_277_1004.n0 VNB 0.79fF
C371 a_277_1004.n1 VNB 0.79fF
C372 a_277_1004.n2 VNB 0.93fF
C373 a_277_1004.n3 VNB 0.29fF
C374 a_277_1004.n4 VNB 0.42fF
C375 a_277_1004.n5 VNB 0.47fF
C376 a_277_1004.n6 VNB 0.87fF
C377 a_277_1004.n7 VNB 0.47fF
C378 a_277_1004.n8 VNB 0.70fF
C379 a_277_1004.n9 VNB 3.48fF
C380 a_277_1004.n10 VNB 0.67fF
C381 a_277_1004.n11 VNB 0.12fF
C382 a_277_1004.n12 VNB 0.45fF
C383 a_277_1004.n13 VNB 0.07fF
C384 a_147_159.n0 VNB 0.37fF
C385 a_147_159.t20 VNB 0.73fF
C386 a_147_159.n1 VNB 0.48fF
C387 a_147_159.n2 VNB 0.42fF
C388 a_147_159.n3 VNB 0.50fF
C389 a_147_159.n4 VNB 0.40fF
C390 a_147_159.n5 VNB 0.69fF
C391 a_147_159.n6 VNB 0.69fF
C392 a_147_159.n7 VNB 0.81fF
C393 a_147_159.n8 VNB 0.25fF
C394 a_147_159.n9 VNB 0.33fF
C395 a_147_159.n10 VNB 0.05fF
C396 a_147_159.n11 VNB 0.07fF
C397 a_147_159.n12 VNB 0.45fF
C398 a_147_159.n13 VNB 0.60fF
C399 a_147_159.n14 VNB 0.71fF
C400 a_147_159.n15 VNB 0.37fF
C401 a_147_159.t21 VNB 0.73fF
C402 a_147_159.n16 VNB 0.48fF
C403 a_147_159.n17 VNB 0.37fF
C404 a_147_159.n18 VNB 0.71fF
C405 a_147_159.n19 VNB 2.70fF
C406 a_147_159.n20 VNB 1.10fF
C407 a_147_159.n21 VNB 0.05fF
C408 a_147_159.n22 VNB 0.07fF
C409 a_147_159.n23 VNB 0.04fF
C410 a_147_159.n24 VNB 0.44fF
C411 a_147_159.n25 VNB 0.57fF
C412 a_147_159.n26 VNB 0.69fF
C413 a_147_159.n27 VNB 0.81fF
C414 a_147_159.n28 VNB 0.25fF
C415 a_147_159.n29 VNB 0.33fF
C416 a_147_159.n30 VNB 0.69fF
C417 a_5457_1004.n0 VNB 0.07fF
C418 a_5457_1004.n1 VNB 0.88fF
C419 a_5457_1004.n2 VNB 0.88fF
C420 a_5457_1004.n3 VNB 1.04fF
C421 a_5457_1004.n4 VNB 0.33fF
C422 a_5457_1004.n5 VNB 0.47fF
C423 a_5457_1004.n6 VNB 0.52fF
C424 a_5457_1004.n7 VNB 0.98fF
C425 a_5457_1004.n8 VNB 0.52fF
C426 a_5457_1004.n9 VNB 0.78fF
C427 a_5457_1004.n10 VNB 3.88fF
C428 a_5457_1004.n11 VNB 0.73fF
C429 a_5457_1004.n12 VNB 0.06fF
C430 a_5457_1004.n13 VNB 0.52fF
C431 a_5457_1004.n14 VNB 0.09fF
C432 a_5779_943.n0 VNB 0.74fF
C433 a_5779_943.n1 VNB 0.74fF
C434 a_5779_943.n2 VNB 0.87fF
C435 a_5779_943.n3 VNB 0.27fF
C436 a_5779_943.n4 VNB 0.44fF
C437 a_5779_943.n5 VNB 0.54fF
C438 a_5779_943.n6 VNB 0.53fF
C439 a_5779_943.n7 VNB 0.54fF
C440 a_5779_943.t11 VNB 0.71fF
C441 a_5779_943.n8 VNB 0.53fF
C442 a_5779_943.n9 VNB 1.72fF
C443 a_5779_943.n10 VNB 0.63fF
C444 a_5779_943.n11 VNB 0.11fF
C445 a_5779_943.n12 VNB 0.38fF
C446 a_5779_943.n13 VNB 0.06fF
C447 a_6514_182.n0 VNB 0.07fF
C448 a_6514_182.n1 VNB 0.13fF
C449 a_6514_182.n2 VNB 0.07fF
C450 a_6514_182.n3 VNB 0.02fF
C451 a_6514_182.n4 VNB 0.03fF
C452 a_6514_182.n5 VNB 0.06fF
C453 a_6514_182.n6 VNB 0.05fF
C454 a_6514_182.n7 VNB 0.06fF
C455 a_6514_182.n8 VNB 0.07fF
C456 a_6514_182.n9 VNB 0.07fF
C457 a_6514_182.n10 VNB 0.03fF
C458 a_6514_182.n11 VNB 0.01fF
C459 a_6514_182.n12 VNB 0.12fF
C460 a_6514_182.t0 VNB 0.28fF
C461 a_6233_75.n0 VNB 0.20fF
C462 a_6233_75.n1 VNB 0.04fF
C463 a_6233_75.n2 VNB 0.01fF
C464 a_6233_75.n3 VNB 0.08fF
C465 a_6233_75.n4 VNB 0.06fF
C466 a_6233_75.n5 VNB 0.07fF
C467 a_9806_73.n0 VNB 0.05fF
C468 a_9806_73.n1 VNB 0.02fF
C469 a_9806_73.n2 VNB 0.12fF
C470 a_9806_73.n3 VNB 0.04fF
C471 a_9806_73.n4 VNB 0.17fF
C472 a_5327_159.n0 VNB 0.07fF
C473 a_5327_159.n1 VNB 0.94fF
C474 a_5327_159.n2 VNB 0.94fF
C475 a_5327_159.n3 VNB 1.11fF
C476 a_5327_159.n4 VNB 0.35fF
C477 a_5327_159.n5 VNB 0.45fF
C478 a_5327_159.n6 VNB 0.51fF
C479 a_5327_159.t7 VNB 1.00fF
C480 a_5327_159.n7 VNB 0.73fF
C481 a_5327_159.n8 VNB 0.51fF
C482 a_5327_159.t9 VNB 1.00fF
C483 a_5327_159.n9 VNB 0.66fF
C484 a_5327_159.n10 VNB 0.50fF
C485 a_5327_159.n11 VNB 0.97fF
C486 a_5327_159.n12 VNB 3.69fF
C487 a_5327_159.n13 VNB 2.91fF
C488 a_5327_159.n14 VNB 0.78fF
C489 a_5327_159.n15 VNB 0.06fF
C490 a_5327_159.n16 VNB 0.60fF
C491 a_5327_159.n17 VNB 0.09fF
C492 a_9331_943.n0 VNB 0.08fF
C493 a_9331_943.n1 VNB 0.78fF
C494 a_9331_943.n2 VNB 0.92fF
C495 a_9331_943.n3 VNB 0.47fF
C496 a_9331_943.n4 VNB 0.38fF
C497 a_9331_943.n5 VNB 0.43fF
C498 a_9331_943.n6 VNB 1.07fF
C499 a_9331_943.n7 VNB 0.79fF
C500 a_9331_943.n8 VNB 0.67fF
C501 a_9331_943.n9 VNB 0.51fF
C502 a_9331_943.n10 VNB 0.69fF
C503 a_9331_943.n11 VNB 3.13fF
C504 a_9331_943.n12 VNB 0.78fF
C505 a_9331_943.n13 VNB 0.92fF
C506 a_9331_943.n14 VNB 0.47fF
C507 a_9331_943.n15 VNB 0.06fF
C508 a_9331_943.n16 VNB 0.08fF
C509 a_9331_943.n17 VNB 0.05fF
C510 a_9331_943.n18 VNB 0.41fF
C511 a_9331_943.n19 VNB 0.61fF
C512 a_9331_943.n20 VNB 0.42fF
C513 a_9331_943.n21 VNB 0.57fF
C514 a_9331_943.n22 VNB 0.56fF
C515 a_9331_943.n23 VNB 0.42fF
C516 a_9331_943.n24 VNB 0.79fF
C517 a_9331_943.n25 VNB 0.79fF
C518 a_9331_943.n26 VNB 0.93fF
C519 a_9331_943.n27 VNB 0.29fF
C520 a_9331_943.n28 VNB 0.47fF
C521 a_9331_943.n29 VNB 0.06fF
C522 a_9331_943.n30 VNB 0.08fF
C523 a_9331_943.n31 VNB 0.05fF
C524 a_9331_943.n32 VNB 0.41fF
C525 a_9331_943.n33 VNB 0.65fF
C526 a_9331_943.n34 VNB 0.91fF
C527 a_9331_943.n35 VNB 0.57fF
C528 a_9331_943.t22 VNB 0.76fF
C529 a_9331_943.n36 VNB 0.53fF
C530 a_9331_943.n37 VNB 1.17fF
C531 a_9331_943.n38 VNB 0.57fF
C532 a_9331_943.t25 VNB 0.76fF
C533 a_9331_943.n39 VNB 0.55fF
C534 a_9331_943.n40 VNB 1.50fF
C535 a_9331_943.n41 VNB 0.61fF
C536 a_9331_943.n42 VNB 0.04fF
C537 a_9331_943.n43 VNB 0.41fF
C538 a_9331_943.n44 VNB 0.07fF
C539 a_14511_943.n0 VNB 0.59fF
C540 a_14511_943.n1 VNB 0.32fF
C541 a_14511_943.n2 VNB 0.36fF
C542 a_14511_943.t12 VNB 0.64fF
C543 a_14511_943.n3 VNB 1.08fF
C544 a_14511_943.n4 VNB 0.76fF
C545 a_14511_943.t11 VNB 0.61fF
C546 a_14511_943.n5 VNB 0.34fF
C547 a_14511_943.n6 VNB 0.40fF
C548 a_14511_943.t5 VNB 0.61fF
C549 a_14511_943.n7 VNB 0.42fF
C550 a_14511_943.n8 VNB 1.27fF
C551 a_14511_943.n9 VNB 0.05fF
C552 a_14511_943.n10 VNB 0.06fF
C553 a_14511_943.n11 VNB 0.04fF
C554 a_14511_943.n12 VNB 0.35fF
C555 a_14511_943.n13 VNB 0.47fF
C556 a_14511_943.n14 VNB 0.32fF
C557 a_14511_943.n15 VNB 0.70fF
C558 VPB.n0 VNB 0.03fF
C559 VPB.n1 VNB 0.04fF
C560 VPB.n2 VNB 0.02fF
C561 VPB.n3 VNB 0.19fF
C562 VPB.n5 VNB 0.02fF
C563 VPB.n6 VNB 0.02fF
C564 VPB.n7 VNB 0.02fF
C565 VPB.n8 VNB 0.02fF
C566 VPB.n10 VNB 0.02fF
C567 VPB.n11 VNB 0.02fF
C568 VPB.n12 VNB 0.02fF
C569 VPB.n14 VNB 0.10fF
C570 VPB.n15 VNB 0.10fF
C571 VPB.n16 VNB 0.02fF
C572 VPB.n17 VNB 0.02fF
C573 VPB.n18 VNB 0.02fF
C574 VPB.n19 VNB 0.04fF
C575 VPB.n20 VNB 0.02fF
C576 VPB.n21 VNB 0.29fF
C577 VPB.n22 VNB 0.04fF
C578 VPB.n24 VNB 0.02fF
C579 VPB.n25 VNB 0.02fF
C580 VPB.n26 VNB 0.02fF
C581 VPB.n27 VNB 0.02fF
C582 VPB.n29 VNB 0.02fF
C583 VPB.n30 VNB 0.02fF
C584 VPB.n31 VNB 0.02fF
C585 VPB.n33 VNB 0.28fF
C586 VPB.n35 VNB 0.03fF
C587 VPB.n36 VNB 0.02fF
C588 VPB.n37 VNB 0.03fF
C589 VPB.n38 VNB 0.03fF
C590 VPB.n39 VNB 0.28fF
C591 VPB.n40 VNB 0.01fF
C592 VPB.n41 VNB 0.02fF
C593 VPB.n42 VNB 0.28fF
C594 VPB.n43 VNB 0.02fF
C595 VPB.n44 VNB 0.02fF
C596 VPB.n45 VNB 0.05fF
C597 VPB.n46 VNB 0.21fF
C598 VPB.n47 VNB 0.02fF
C599 VPB.n48 VNB 0.01fF
C600 VPB.n49 VNB 0.14fF
C601 VPB.n50 VNB 0.16fF
C602 VPB.n51 VNB 0.02fF
C603 VPB.n52 VNB 0.02fF
C604 VPB.n53 VNB 0.14fF
C605 VPB.n54 VNB 0.16fF
C606 VPB.n55 VNB 0.02fF
C607 VPB.n56 VNB 0.02fF
C608 VPB.n57 VNB 0.02fF
C609 VPB.n58 VNB 0.14fF
C610 VPB.n59 VNB 0.15fF
C611 VPB.n60 VNB 0.02fF
C612 VPB.n61 VNB 0.02fF
C613 VPB.n62 VNB 0.14fF
C614 VPB.n63 VNB 0.15fF
C615 VPB.n64 VNB 0.02fF
C616 VPB.n65 VNB 0.02fF
C617 VPB.n66 VNB 0.02fF
C618 VPB.n67 VNB 0.14fF
C619 VPB.n68 VNB 0.16fF
C620 VPB.n69 VNB 0.02fF
C621 VPB.n70 VNB 0.02fF
C622 VPB.n71 VNB 0.14fF
C623 VPB.n72 VNB 0.16fF
C624 VPB.n73 VNB 0.02fF
C625 VPB.n74 VNB 0.02fF
C626 VPB.n75 VNB 0.21fF
C627 VPB.n76 VNB 0.02fF
C628 VPB.n77 VNB 0.01fF
C629 VPB.n78 VNB 0.06fF
C630 VPB.n79 VNB 0.28fF
C631 VPB.n80 VNB 0.02fF
C632 VPB.n81 VNB 0.02fF
C633 VPB.n82 VNB 0.02fF
C634 VPB.n83 VNB 0.02fF
C635 VPB.n84 VNB 0.02fF
C636 VPB.n85 VNB 0.04fF
C637 VPB.n86 VNB 0.02fF
C638 VPB.n87 VNB 0.29fF
C639 VPB.n88 VNB 0.04fF
C640 VPB.n90 VNB 0.02fF
C641 VPB.n91 VNB 0.02fF
C642 VPB.n92 VNB 0.02fF
C643 VPB.n93 VNB 0.02fF
C644 VPB.n95 VNB 0.02fF
C645 VPB.n96 VNB 0.02fF
C646 VPB.n97 VNB 0.02fF
C647 VPB.n99 VNB 0.28fF
C648 VPB.n101 VNB 0.03fF
C649 VPB.n102 VNB 0.02fF
C650 VPB.n103 VNB 0.10fF
C651 VPB.n104 VNB 0.10fF
C652 VPB.n105 VNB 0.02fF
C653 VPB.n106 VNB 0.02fF
C654 VPB.n107 VNB 0.02fF
C655 VPB.n108 VNB 0.04fF
C656 VPB.n109 VNB 0.02fF
C657 VPB.n110 VNB 0.24fF
C658 VPB.n111 VNB 0.04fF
C659 VPB.n113 VNB 0.02fF
C660 VPB.n114 VNB 0.02fF
C661 VPB.n115 VNB 0.02fF
C662 VPB.n116 VNB 0.02fF
C663 VPB.n118 VNB 0.02fF
C664 VPB.n119 VNB 0.02fF
C665 VPB.n120 VNB 0.02fF
C666 VPB.n122 VNB 0.28fF
C667 VPB.n124 VNB 0.03fF
C668 VPB.n125 VNB 0.02fF
C669 VPB.n126 VNB 0.03fF
C670 VPB.n127 VNB 0.03fF
C671 VPB.n128 VNB 0.28fF
C672 VPB.n129 VNB 0.01fF
C673 VPB.n130 VNB 0.02fF
C674 VPB.n131 VNB 0.28fF
C675 VPB.n132 VNB 0.02fF
C676 VPB.n133 VNB 0.02fF
C677 VPB.n134 VNB 0.05fF
C678 VPB.n135 VNB 0.21fF
C679 VPB.n136 VNB 0.02fF
C680 VPB.n137 VNB 0.01fF
C681 VPB.n138 VNB 0.14fF
C682 VPB.n139 VNB 0.16fF
C683 VPB.n140 VNB 0.02fF
C684 VPB.n141 VNB 0.02fF
C685 VPB.n142 VNB 0.14fF
C686 VPB.n143 VNB 0.16fF
C687 VPB.n144 VNB 0.02fF
C688 VPB.n145 VNB 0.02fF
C689 VPB.n146 VNB 0.02fF
C690 VPB.n147 VNB 0.14fF
C691 VPB.n148 VNB 0.15fF
C692 VPB.n149 VNB 0.02fF
C693 VPB.n150 VNB 0.02fF
C694 VPB.n151 VNB 0.14fF
C695 VPB.n152 VNB 0.15fF
C696 VPB.n153 VNB 0.02fF
C697 VPB.n154 VNB 0.02fF
C698 VPB.n155 VNB 0.02fF
C699 VPB.n156 VNB 0.14fF
C700 VPB.n157 VNB 0.16fF
C701 VPB.n158 VNB 0.02fF
C702 VPB.n159 VNB 0.02fF
C703 VPB.n160 VNB 0.14fF
C704 VPB.n161 VNB 0.16fF
C705 VPB.n162 VNB 0.02fF
C706 VPB.n163 VNB 0.02fF
C707 VPB.n164 VNB 0.21fF
C708 VPB.n165 VNB 0.02fF
C709 VPB.n166 VNB 0.01fF
C710 VPB.n167 VNB 0.06fF
C711 VPB.n168 VNB 0.28fF
C712 VPB.n169 VNB 0.02fF
C713 VPB.n170 VNB 0.02fF
C714 VPB.n171 VNB 0.02fF
C715 VPB.n172 VNB 0.02fF
C716 VPB.n173 VNB 0.02fF
C717 VPB.n174 VNB 0.14fF
C718 VPB.n175 VNB 0.03fF
C719 VPB.n176 VNB 0.02fF
C720 VPB.n177 VNB 0.05fF
C721 VPB.n178 VNB 0.01fF
C722 VPB.n179 VNB 0.02fF
C723 VPB.n180 VNB 0.02fF
C724 VPB.n183 VNB 0.02fF
C725 VPB.n184 VNB 0.02fF
C726 VPB.n185 VNB 0.02fF
C727 VPB.n188 VNB 0.46fF
C728 VPB.n190 VNB 0.04fF
C729 VPB.n191 VNB 0.04fF
C730 VPB.n192 VNB 0.28fF
C731 VPB.n193 VNB 0.03fF
C732 VPB.n194 VNB 0.04fF
C733 VPB.n195 VNB 0.28fF
C734 VPB.n196 VNB 0.02fF
C735 VPB.n197 VNB 0.02fF
C736 VPB.n198 VNB 0.28fF
C737 VPB.n199 VNB 0.02fF
C738 VPB.n200 VNB 0.02fF
C739 VPB.n201 VNB 0.28fF
C740 VPB.n202 VNB 0.02fF
C741 VPB.n203 VNB 0.02fF
C742 VPB.n204 VNB 0.00fF
C743 VPB.n205 VNB 0.10fF
C744 VPB.n206 VNB 0.02fF
C745 VPB.n207 VNB 0.28fF
C746 VPB.n208 VNB 0.02fF
C747 VPB.n209 VNB 0.02fF
C748 VPB.n210 VNB 0.02fF
C749 VPB.n211 VNB 0.28fF
C750 VPB.n212 VNB 0.02fF
C751 VPB.n213 VNB 0.02fF
C752 VPB.n214 VNB 0.02fF
C753 VPB.n215 VNB 0.28fF
C754 VPB.n216 VNB 0.02fF
C755 VPB.n217 VNB 0.02fF
C756 VPB.n218 VNB 0.02fF
C757 VPB.n219 VNB 0.28fF
C758 VPB.n220 VNB 0.01fF
C759 VPB.n221 VNB 0.02fF
C760 VPB.n222 VNB 0.04fF
C761 VPB.n223 VNB 0.02fF
C762 VPB.n224 VNB 0.02fF
C763 VPB.n225 VNB 0.02fF
C764 VPB.n226 VNB 0.04fF
C765 VPB.n227 VNB 0.02fF
C766 VPB.n228 VNB 0.20fF
C767 VPB.n229 VNB 0.04fF
C768 VPB.n231 VNB 0.02fF
C769 VPB.n232 VNB 0.02fF
C770 VPB.n233 VNB 0.02fF
C771 VPB.n234 VNB 0.02fF
C772 VPB.n236 VNB 0.02fF
C773 VPB.n237 VNB 0.02fF
C774 VPB.n238 VNB 0.02fF
C775 VPB.n240 VNB 0.28fF
C776 VPB.n242 VNB 0.03fF
C777 VPB.n243 VNB 0.02fF
C778 VPB.n244 VNB 0.03fF
C779 VPB.n245 VNB 0.03fF
C780 VPB.n246 VNB 0.28fF
C781 VPB.n247 VNB 0.01fF
C782 VPB.n248 VNB 0.02fF
C783 VPB.n249 VNB 0.04fF
C784 VPB.n250 VNB 0.28fF
C785 VPB.n251 VNB 0.02fF
C786 VPB.n252 VNB 0.02fF
C787 VPB.n253 VNB 0.02fF
C788 VPB.n254 VNB 0.28fF
C789 VPB.n255 VNB 0.02fF
C790 VPB.n256 VNB 0.02fF
C791 VPB.n257 VNB 0.02fF
C792 VPB.n258 VNB 0.28fF
C793 VPB.n259 VNB 0.02fF
C794 VPB.n260 VNB 0.02fF
C795 VPB.n261 VNB 0.02fF
C796 VPB.n262 VNB 0.28fF
C797 VPB.n263 VNB 0.02fF
C798 VPB.n264 VNB 0.02fF
C799 VPB.n265 VNB 0.02fF
C800 VPB.n266 VNB 0.28fF
C801 VPB.n267 VNB 0.02fF
C802 VPB.n268 VNB 0.02fF
C803 VPB.n269 VNB 0.02fF
C804 VPB.n270 VNB 0.28fF
C805 VPB.n271 VNB 0.02fF
C806 VPB.n272 VNB 0.02fF
C807 VPB.n273 VNB 0.02fF
C808 VPB.n274 VNB 0.28fF
C809 VPB.n275 VNB 0.01fF
C810 VPB.n276 VNB 0.02fF
C811 VPB.n277 VNB 0.04fF
C812 VPB.n278 VNB 0.02fF
C813 VPB.n279 VNB 0.02fF
C814 VPB.n280 VNB 0.02fF
C815 VPB.n281 VNB 0.04fF
C816 VPB.n282 VNB 0.02fF
C817 VPB.n283 VNB 0.20fF
C818 VPB.n284 VNB 0.04fF
C819 VPB.n286 VNB 0.02fF
C820 VPB.n287 VNB 0.02fF
C821 VPB.n288 VNB 0.02fF
C822 VPB.n289 VNB 0.02fF
C823 VPB.n291 VNB 0.02fF
C824 VPB.n292 VNB 0.02fF
C825 VPB.n293 VNB 0.02fF
C826 VPB.n295 VNB 0.28fF
C827 VPB.n297 VNB 0.03fF
C828 VPB.n298 VNB 0.02fF
C829 VPB.n299 VNB 0.03fF
C830 VPB.n300 VNB 0.03fF
C831 VPB.n301 VNB 0.28fF
C832 VPB.n302 VNB 0.01fF
C833 VPB.n303 VNB 0.02fF
C834 VPB.n304 VNB 0.04fF
C835 VPB.n305 VNB 0.06fF
C836 VPB.n306 VNB 0.23fF
C837 VPB.n307 VNB 0.02fF
C838 VPB.n308 VNB 0.01fF
C839 VPB.n309 VNB 0.02fF
C840 VPB.n310 VNB 0.14fF
C841 VPB.n311 VNB 0.16fF
C842 VPB.n312 VNB 0.02fF
C843 VPB.n313 VNB 0.02fF
C844 VPB.n314 VNB 0.02fF
C845 VPB.n315 VNB 0.10fF
C846 VPB.n316 VNB 0.02fF
C847 VPB.n317 VNB 0.14fF
C848 VPB.n318 VNB 0.15fF
C849 VPB.n319 VNB 0.02fF
C850 VPB.n320 VNB 0.02fF
C851 VPB.n321 VNB 0.02fF
C852 VPB.n322 VNB 0.14fF
C853 VPB.n323 VNB 0.15fF
C854 VPB.n324 VNB 0.02fF
C855 VPB.n325 VNB 0.02fF
C856 VPB.n326 VNB 0.02fF
C857 VPB.n327 VNB 0.14fF
C858 VPB.n328 VNB 0.16fF
C859 VPB.n329 VNB 0.02fF
C860 VPB.n330 VNB 0.02fF
C861 VPB.n331 VNB 0.02fF
C862 VPB.n332 VNB 0.06fF
C863 VPB.n333 VNB 0.24fF
C864 VPB.n334 VNB 0.02fF
C865 VPB.n335 VNB 0.01fF
C866 VPB.n336 VNB 0.02fF
C867 VPB.n337 VNB 0.28fF
C868 VPB.n338 VNB 0.01fF
C869 VPB.n339 VNB 0.02fF
C870 VPB.n340 VNB 0.04fF
C871 VPB.n341 VNB 0.02fF
C872 VPB.n342 VNB 0.02fF
C873 VPB.n343 VNB 0.02fF
C874 VPB.n344 VNB 0.04fF
C875 VPB.n345 VNB 0.02fF
C876 VPB.n346 VNB 0.20fF
C877 VPB.n347 VNB 0.04fF
C878 VPB.n349 VNB 0.02fF
C879 VPB.n350 VNB 0.02fF
C880 VPB.n351 VNB 0.02fF
C881 VPB.n352 VNB 0.02fF
C882 VPB.n354 VNB 0.02fF
C883 VPB.n355 VNB 0.02fF
C884 VPB.n356 VNB 0.02fF
C885 VPB.n358 VNB 0.28fF
C886 VPB.n360 VNB 0.03fF
C887 VPB.n361 VNB 0.02fF
C888 VPB.n362 VNB 0.03fF
C889 VPB.n363 VNB 0.03fF
C890 VPB.n364 VNB 0.28fF
C891 VPB.n365 VNB 0.01fF
C892 VPB.n366 VNB 0.02fF
C893 VPB.n367 VNB 0.04fF
C894 VPB.n368 VNB 0.05fF
C895 VPB.n369 VNB 0.23fF
C896 VPB.n370 VNB 0.02fF
C897 VPB.n371 VNB 0.01fF
C898 VPB.n372 VNB 0.02fF
C899 VPB.n373 VNB 0.14fF
C900 VPB.n374 VNB 0.16fF
C901 VPB.n375 VNB 0.02fF
C902 VPB.n376 VNB 0.02fF
C903 VPB.n377 VNB 0.02fF
C904 VPB.n378 VNB 0.10fF
C905 VPB.n379 VNB 0.02fF
C906 VPB.n380 VNB 0.14fF
C907 VPB.n381 VNB 0.15fF
C908 VPB.n382 VNB 0.02fF
C909 VPB.n383 VNB 0.02fF
C910 VPB.n384 VNB 0.02fF
C911 VPB.n385 VNB 0.14fF
C912 VPB.n386 VNB 0.15fF
C913 VPB.n387 VNB 0.02fF
C914 VPB.n388 VNB 0.02fF
C915 VPB.n389 VNB 0.02fF
C916 VPB.n390 VNB 0.14fF
C917 VPB.n391 VNB 0.16fF
C918 VPB.n392 VNB 0.02fF
C919 VPB.n393 VNB 0.02fF
C920 VPB.n394 VNB 0.02fF
C921 VPB.n395 VNB 0.06fF
C922 VPB.n396 VNB 0.24fF
C923 VPB.n397 VNB 0.02fF
C924 VPB.n398 VNB 0.01fF
C925 VPB.n399 VNB 0.02fF
C926 VPB.n400 VNB 0.28fF
C927 VPB.n401 VNB 0.01fF
C928 VPB.n402 VNB 0.02fF
C929 VPB.n403 VNB 0.04fF
C930 VPB.n404 VNB 0.02fF
C931 VPB.n405 VNB 0.02fF
C932 VPB.n406 VNB 0.02fF
C933 VPB.n407 VNB 0.04fF
C934 VPB.n408 VNB 0.02fF
C935 VPB.n409 VNB 0.24fF
C936 VPB.n410 VNB 0.04fF
C937 VPB.n412 VNB 0.02fF
C938 VPB.n413 VNB 0.02fF
C939 VPB.n414 VNB 0.02fF
C940 VPB.n415 VNB 0.02fF
C941 VPB.n417 VNB 0.02fF
C942 VPB.n418 VNB 0.02fF
C943 VPB.n419 VNB 0.02fF
C944 VPB.n421 VNB 0.28fF
C945 VPB.n423 VNB 0.03fF
C946 VPB.n424 VNB 0.02fF
C947 VPB.n425 VNB 0.03fF
C948 VPB.n426 VNB 0.03fF
C949 VPB.n427 VNB 0.28fF
C950 VPB.n428 VNB 0.01fF
C951 VPB.n429 VNB 0.02fF
C952 VPB.n430 VNB 0.04fF
C953 VPB.n431 VNB 0.28fF
C954 VPB.n432 VNB 0.02fF
C955 VPB.n433 VNB 0.02fF
C956 VPB.n434 VNB 0.02fF
C957 VPB.n435 VNB 0.05fF
C958 VPB.n436 VNB 0.21fF
C959 VPB.n437 VNB 0.02fF
C960 VPB.n438 VNB 0.01fF
C961 VPB.n439 VNB 0.02fF
C962 VPB.n440 VNB 0.14fF
C963 VPB.n441 VNB 0.16fF
C964 VPB.n442 VNB 0.02fF
C965 VPB.n443 VNB 0.02fF
C966 VPB.n444 VNB 0.02fF
C967 VPB.n445 VNB 0.10fF
C968 VPB.n446 VNB 0.02fF
C969 VPB.n447 VNB 0.14fF
C970 VPB.n448 VNB 0.16fF
C971 VPB.n449 VNB 0.02fF
C972 VPB.n450 VNB 0.02fF
C973 VPB.n451 VNB 0.02fF
C974 VPB.n452 VNB 0.14fF
C975 VPB.n453 VNB 0.15fF
C976 VPB.n454 VNB 0.02fF
C977 VPB.n455 VNB 0.02fF
C978 VPB.n456 VNB 0.02fF
C979 VPB.n457 VNB 0.14fF
C980 VPB.n458 VNB 0.15fF
C981 VPB.n459 VNB 0.02fF
C982 VPB.n460 VNB 0.02fF
C983 VPB.n461 VNB 0.02fF
C984 VPB.n462 VNB 0.10fF
C985 VPB.n463 VNB 0.02fF
C986 VPB.n464 VNB 0.14fF
C987 VPB.n465 VNB 0.16fF
C988 VPB.n466 VNB 0.02fF
C989 VPB.n467 VNB 0.02fF
C990 VPB.n468 VNB 0.02fF
C991 VPB.n469 VNB 0.14fF
C992 VPB.n470 VNB 0.16fF
C993 VPB.n471 VNB 0.02fF
C994 VPB.n472 VNB 0.02fF
C995 VPB.n473 VNB 0.02fF
C996 VPB.n474 VNB 0.06fF
C997 VPB.n475 VNB 0.21fF
C998 VPB.n476 VNB 0.02fF
C999 VPB.n477 VNB 0.01fF
C1000 VPB.n478 VNB 0.02fF
C1001 VPB.n479 VNB 0.28fF
C1002 VPB.n480 VNB 0.02fF
C1003 VPB.n481 VNB 0.02fF
C1004 VPB.n482 VNB 0.02fF
C1005 VPB.n483 VNB 0.28fF
C1006 VPB.n484 VNB 0.01fF
C1007 VPB.n485 VNB 0.02fF
C1008 VPB.n486 VNB 0.04fF
C1009 VPB.n487 VNB 0.02fF
C1010 VPB.n488 VNB 0.02fF
C1011 VPB.n489 VNB 0.02fF
C1012 VPB.n490 VNB 0.04fF
C1013 VPB.n491 VNB 0.02fF
C1014 VPB.n492 VNB 0.29fF
C1015 VPB.n493 VNB 0.04fF
C1016 VPB.n495 VNB 0.02fF
C1017 VPB.n496 VNB 0.02fF
C1018 VPB.n497 VNB 0.02fF
C1019 VPB.n498 VNB 0.02fF
C1020 VPB.n500 VNB 0.02fF
C1021 VPB.n501 VNB 0.02fF
C1022 VPB.n502 VNB 0.02fF
C1023 VPB.n504 VNB 0.28fF
C1024 VPB.n506 VNB 0.03fF
C1025 VPB.n507 VNB 0.02fF
C1026 VPB.n508 VNB 0.03fF
C1027 VPB.n509 VNB 0.03fF
C1028 VPB.n510 VNB 0.28fF
C1029 VPB.n511 VNB 0.01fF
C1030 VPB.n512 VNB 0.02fF
C1031 VPB.n513 VNB 0.04fF
C1032 VPB.n514 VNB 0.28fF
C1033 VPB.n515 VNB 0.02fF
C1034 VPB.n516 VNB 0.02fF
C1035 VPB.n517 VNB 0.02fF
C1036 VPB.n518 VNB 0.05fF
C1037 VPB.n519 VNB 0.21fF
C1038 VPB.n520 VNB 0.02fF
C1039 VPB.n521 VNB 0.01fF
C1040 VPB.n522 VNB 0.02fF
C1041 VPB.n523 VNB 0.14fF
C1042 VPB.n524 VNB 0.16fF
C1043 VPB.n525 VNB 0.02fF
C1044 VPB.n526 VNB 0.02fF
C1045 VPB.n527 VNB 0.02fF
C1046 VPB.n528 VNB 0.10fF
C1047 VPB.n529 VNB 0.02fF
C1048 VPB.n530 VNB 0.14fF
C1049 VPB.n531 VNB 0.16fF
C1050 VPB.n532 VNB 0.02fF
C1051 VPB.n533 VNB 0.02fF
C1052 VPB.n534 VNB 0.02fF
C1053 VPB.n535 VNB 0.14fF
C1054 VPB.n536 VNB 0.15fF
C1055 VPB.n537 VNB 0.02fF
C1056 VPB.n538 VNB 0.02fF
C1057 VPB.n539 VNB 0.02fF
C1058 VPB.n540 VNB 0.14fF
C1059 VPB.n541 VNB 0.15fF
C1060 VPB.n542 VNB 0.02fF
C1061 VPB.n543 VNB 0.02fF
C1062 VPB.n544 VNB 0.02fF
C1063 VPB.n545 VNB 0.10fF
C1064 VPB.n546 VNB 0.02fF
C1065 VPB.n547 VNB 0.14fF
C1066 VPB.n548 VNB 0.16fF
C1067 VPB.n549 VNB 0.02fF
C1068 VPB.n550 VNB 0.02fF
C1069 VPB.n551 VNB 0.02fF
C1070 VPB.n552 VNB 0.14fF
C1071 VPB.n553 VNB 0.16fF
C1072 VPB.n554 VNB 0.02fF
C1073 VPB.n555 VNB 0.02fF
C1074 VPB.n556 VNB 0.02fF
C1075 VPB.n557 VNB 0.06fF
C1076 VPB.n558 VNB 0.21fF
C1077 VPB.n559 VNB 0.02fF
C1078 VPB.n560 VNB 0.01fF
C1079 VPB.n561 VNB 0.02fF
C1080 VPB.n562 VNB 0.28fF
C1081 VPB.n563 VNB 0.02fF
C1082 VPB.n564 VNB 0.02fF
C1083 VPB.n565 VNB 0.02fF
C1084 VPB.n566 VNB 0.28fF
C1085 VPB.n567 VNB 0.01fF
C1086 VPB.n568 VNB 0.02fF
C1087 VPB.n569 VNB 0.04fF
C1088 VPB.n570 VNB 0.02fF
C1089 VPB.n571 VNB 0.02fF
C1090 VPB.n572 VNB 0.02fF
C1091 VPB.n573 VNB 0.04fF
C1092 VPB.n574 VNB 0.02fF
C1093 VPB.n575 VNB 0.24fF
C1094 VPB.n576 VNB 0.04fF
C1095 VPB.n578 VNB 0.02fF
C1096 VPB.n579 VNB 0.02fF
C1097 VPB.n580 VNB 0.02fF
C1098 VPB.n581 VNB 0.02fF
C1099 VPB.n583 VNB 0.02fF
C1100 VPB.n584 VNB 0.02fF
C1101 VPB.n585 VNB 0.02fF
C1102 VPB.n587 VNB 0.28fF
C1103 VPB.n589 VNB 0.03fF
C1104 VPB.n590 VNB 0.02fF
C1105 VPB.n591 VNB 0.03fF
C1106 VPB.n592 VNB 0.03fF
C1107 VPB.n593 VNB 0.28fF
C1108 VPB.n594 VNB 0.01fF
C1109 VPB.n595 VNB 0.02fF
C1110 VPB.n596 VNB 0.04fF
C1111 VPB.n597 VNB 0.05fF
C1112 VPB.n598 VNB 0.23fF
C1113 VPB.n599 VNB 0.02fF
C1114 VPB.n600 VNB 0.01fF
C1115 VPB.n601 VNB 0.02fF
C1116 VPB.n602 VNB 0.14fF
C1117 VPB.n603 VNB 0.16fF
C1118 VPB.n604 VNB 0.02fF
C1119 VPB.n605 VNB 0.02fF
C1120 VPB.n606 VNB 0.02fF
C1121 VPB.n607 VNB 0.10fF
C1122 VPB.n608 VNB 0.02fF
C1123 VPB.n609 VNB 0.14fF
C1124 VPB.n610 VNB 0.15fF
C1125 VPB.n611 VNB 0.02fF
C1126 VPB.n612 VNB 0.02fF
C1127 VPB.n613 VNB 0.02fF
C1128 VPB.n614 VNB 0.14fF
C1129 VPB.n615 VNB 0.15fF
C1130 VPB.n616 VNB 0.02fF
C1131 VPB.n617 VNB 0.02fF
C1132 VPB.n618 VNB 0.02fF
C1133 VPB.n619 VNB 0.14fF
C1134 VPB.n620 VNB 0.16fF
C1135 VPB.n621 VNB 0.02fF
C1136 VPB.n622 VNB 0.02fF
C1137 VPB.n623 VNB 0.02fF
C1138 VPB.n624 VNB 0.06fF
C1139 VPB.n625 VNB 0.24fF
C1140 VPB.n626 VNB 0.02fF
C1141 VPB.n627 VNB 0.01fF
C1142 VPB.n628 VNB 0.02fF
C1143 VPB.n629 VNB 0.28fF
C1144 VPB.n630 VNB 0.01fF
C1145 VPB.n631 VNB 0.02fF
C1146 VPB.n632 VNB 0.04fF
C1147 VPB.n633 VNB 0.02fF
C1148 VPB.n634 VNB 0.02fF
C1149 VPB.n635 VNB 0.02fF
C1150 VPB.n636 VNB 0.04fF
C1151 VPB.n637 VNB 0.02fF
C1152 VPB.n638 VNB 0.24fF
C1153 VPB.n639 VNB 0.04fF
C1154 VPB.n641 VNB 0.02fF
C1155 VPB.n642 VNB 0.02fF
C1156 VPB.n643 VNB 0.02fF
C1157 VPB.n644 VNB 0.02fF
C1158 VPB.n646 VNB 0.02fF
C1159 VPB.n647 VNB 0.02fF
C1160 VPB.n648 VNB 0.02fF
C1161 VPB.n650 VNB 0.28fF
C1162 VPB.n652 VNB 0.03fF
C1163 VPB.n653 VNB 0.02fF
C1164 VPB.n654 VNB 0.03fF
C1165 VPB.n655 VNB 0.03fF
C1166 VPB.n656 VNB 0.28fF
C1167 VPB.n657 VNB 0.01fF
C1168 VPB.n658 VNB 0.02fF
C1169 VPB.n659 VNB 0.04fF
C1170 VPB.n660 VNB 0.28fF
C1171 VPB.n661 VNB 0.02fF
C1172 VPB.n662 VNB 0.02fF
C1173 VPB.n663 VNB 0.02fF
C1174 VPB.n664 VNB 0.05fF
C1175 VPB.n665 VNB 0.21fF
C1176 VPB.n666 VNB 0.02fF
C1177 VPB.n667 VNB 0.01fF
C1178 VPB.n668 VNB 0.02fF
C1179 VPB.n669 VNB 0.14fF
C1180 VPB.n670 VNB 0.16fF
C1181 VPB.n671 VNB 0.02fF
C1182 VPB.n672 VNB 0.02fF
C1183 VPB.n673 VNB 0.02fF
C1184 VPB.n674 VNB 0.10fF
C1185 VPB.n675 VNB 0.02fF
C1186 VPB.n676 VNB 0.14fF
C1187 VPB.n677 VNB 0.16fF
C1188 VPB.n678 VNB 0.02fF
C1189 VPB.n679 VNB 0.02fF
C1190 VPB.n680 VNB 0.02fF
C1191 VPB.n681 VNB 0.14fF
C1192 VPB.n682 VNB 0.15fF
C1193 VPB.n683 VNB 0.02fF
C1194 VPB.n684 VNB 0.02fF
C1195 VPB.n685 VNB 0.02fF
C1196 VPB.n686 VNB 0.14fF
C1197 VPB.n687 VNB 0.15fF
C1198 VPB.n688 VNB 0.02fF
C1199 VPB.n689 VNB 0.02fF
C1200 VPB.n690 VNB 0.02fF
C1201 VPB.n691 VNB 0.10fF
C1202 VPB.n692 VNB 0.02fF
C1203 VPB.n693 VNB 0.14fF
C1204 VPB.n694 VNB 0.16fF
C1205 VPB.n695 VNB 0.02fF
C1206 VPB.n696 VNB 0.02fF
C1207 VPB.n697 VNB 0.02fF
C1208 VPB.n698 VNB 0.14fF
C1209 VPB.n699 VNB 0.16fF
C1210 VPB.n700 VNB 0.02fF
C1211 VPB.n701 VNB 0.02fF
C1212 VPB.n702 VNB 0.02fF
C1213 VPB.n703 VNB 0.06fF
C1214 VPB.n704 VNB 0.21fF
C1215 VPB.n705 VNB 0.02fF
C1216 VPB.n706 VNB 0.01fF
C1217 VPB.n707 VNB 0.02fF
C1218 VPB.n708 VNB 0.28fF
C1219 VPB.n709 VNB 0.02fF
C1220 VPB.n710 VNB 0.02fF
C1221 VPB.n711 VNB 0.02fF
C1222 VPB.n712 VNB 0.28fF
C1223 VPB.n713 VNB 0.01fF
C1224 VPB.n714 VNB 0.02fF
C1225 VPB.n715 VNB 0.04fF
C1226 VPB.n716 VNB 0.02fF
C1227 VPB.n717 VNB 0.02fF
C1228 VPB.n718 VNB 0.02fF
C1229 VPB.n719 VNB 0.04fF
C1230 VPB.n720 VNB 0.02fF
C1231 VPB.n721 VNB 0.29fF
C1232 VPB.n722 VNB 0.04fF
C1233 VPB.n724 VNB 0.02fF
C1234 VPB.n725 VNB 0.02fF
C1235 VPB.n726 VNB 0.02fF
C1236 VPB.n727 VNB 0.02fF
C1237 VPB.n729 VNB 0.02fF
C1238 VPB.n730 VNB 0.02fF
C1239 VPB.n731 VNB 0.02fF
C1240 VPB.n733 VNB 0.28fF
C1241 VPB.n735 VNB 0.03fF
C1242 VPB.n736 VNB 0.02fF
C1243 VPB.n737 VNB 0.03fF
C1244 VPB.n738 VNB 0.03fF
C1245 VPB.n739 VNB 0.28fF
C1246 VPB.n740 VNB 0.01fF
C1247 VPB.n741 VNB 0.02fF
C1248 VPB.n742 VNB 0.04fF
C1249 VPB.n743 VNB 0.28fF
C1250 VPB.n744 VNB 0.02fF
C1251 VPB.n745 VNB 0.02fF
C1252 VPB.n746 VNB 0.02fF
C1253 VPB.n747 VNB 0.05fF
C1254 VPB.n748 VNB 0.21fF
C1255 VPB.n749 VNB 0.02fF
C1256 VPB.n750 VNB 0.01fF
C1257 VPB.n751 VNB 0.02fF
C1258 VPB.n752 VNB 0.14fF
C1259 VPB.n753 VNB 0.16fF
C1260 VPB.n754 VNB 0.02fF
C1261 VPB.n755 VNB 0.02fF
C1262 VPB.n756 VNB 0.02fF
C1263 VPB.n757 VNB 0.10fF
C1264 VPB.n758 VNB 0.02fF
C1265 VPB.n759 VNB 0.14fF
C1266 VPB.n760 VNB 0.16fF
C1267 VPB.n761 VNB 0.02fF
C1268 VPB.n762 VNB 0.02fF
C1269 VPB.n763 VNB 0.02fF
C1270 VPB.n764 VNB 0.14fF
C1271 VPB.n765 VNB 0.15fF
C1272 VPB.n766 VNB 0.02fF
C1273 VPB.n767 VNB 0.02fF
C1274 VPB.n768 VNB 0.02fF
C1275 VPB.n769 VNB 0.14fF
C1276 VPB.n770 VNB 0.15fF
C1277 VPB.n771 VNB 0.02fF
C1278 VPB.n772 VNB 0.02fF
C1279 VPB.n773 VNB 0.02fF
C1280 VPB.n774 VNB 0.10fF
C1281 VPB.n775 VNB 0.02fF
C1282 VPB.n776 VNB 0.14fF
C1283 VPB.n777 VNB 0.16fF
C1284 VPB.n778 VNB 0.02fF
C1285 VPB.n779 VNB 0.02fF
C1286 VPB.n780 VNB 0.02fF
C1287 VPB.n781 VNB 0.14fF
C1288 VPB.n782 VNB 0.16fF
C1289 VPB.n783 VNB 0.02fF
C1290 VPB.n784 VNB 0.02fF
C1291 VPB.n785 VNB 0.02fF
C1292 VPB.n786 VNB 0.06fF
C1293 VPB.n787 VNB 0.21fF
C1294 VPB.n788 VNB 0.02fF
C1295 VPB.n789 VNB 0.01fF
C1296 VPB.n790 VNB 0.02fF
C1297 VPB.n791 VNB 0.28fF
C1298 VPB.n792 VNB 0.02fF
C1299 VPB.n793 VNB 0.02fF
C1300 VPB.n794 VNB 0.02fF
C1301 VPB.n795 VNB 0.28fF
C1302 VPB.n796 VNB 0.01fF
C1303 VPB.n797 VNB 0.02fF
C1304 VPB.n798 VNB 0.04fF
C1305 VPB.n799 VNB 0.02fF
C1306 VPB.n800 VNB 0.02fF
C1307 VPB.n801 VNB 0.02fF
C1308 VPB.n802 VNB 0.04fF
C1309 VPB.n803 VNB 0.02fF
C1310 VPB.n804 VNB 0.24fF
C1311 VPB.n805 VNB 0.04fF
C1312 VPB.n807 VNB 0.02fF
C1313 VPB.n808 VNB 0.02fF
C1314 VPB.n809 VNB 0.02fF
C1315 VPB.n810 VNB 0.02fF
C1316 VPB.n812 VNB 0.02fF
C1317 VPB.n813 VNB 0.02fF
C1318 VPB.n814 VNB 0.02fF
C1319 VPB.n816 VNB 0.28fF
C1320 VPB.n818 VNB 0.03fF
C1321 VPB.n819 VNB 0.02fF
C1322 VPB.n820 VNB 0.03fF
C1323 VPB.n821 VNB 0.03fF
C1324 VPB.n822 VNB 0.28fF
C1325 VPB.n823 VNB 0.01fF
C1326 VPB.n824 VNB 0.02fF
C1327 VPB.n825 VNB 0.04fF
C1328 VPB.n826 VNB 0.05fF
C1329 VPB.n827 VNB 0.23fF
C1330 VPB.n828 VNB 0.02fF
C1331 VPB.n829 VNB 0.01fF
C1332 VPB.n830 VNB 0.02fF
C1333 VPB.n831 VNB 0.14fF
C1334 VPB.n832 VNB 0.16fF
C1335 VPB.n833 VNB 0.02fF
C1336 VPB.n834 VNB 0.02fF
C1337 VPB.n835 VNB 0.02fF
C1338 VPB.n836 VNB 0.10fF
C1339 VPB.n837 VNB 0.02fF
C1340 VPB.n838 VNB 0.14fF
C1341 VPB.n839 VNB 0.15fF
C1342 VPB.n840 VNB 0.02fF
C1343 VPB.n841 VNB 0.02fF
C1344 VPB.n842 VNB 0.02fF
C1345 VPB.n843 VNB 0.14fF
C1346 VPB.n844 VNB 0.15fF
C1347 VPB.n845 VNB 0.02fF
C1348 VPB.n846 VNB 0.02fF
C1349 VPB.n847 VNB 0.02fF
C1350 VPB.n848 VNB 0.14fF
C1351 VPB.n849 VNB 0.16fF
C1352 VPB.n850 VNB 0.02fF
C1353 VPB.n851 VNB 0.02fF
C1354 VPB.n852 VNB 0.02fF
C1355 VPB.n853 VNB 0.06fF
C1356 VPB.n854 VNB 0.24fF
C1357 VPB.n855 VNB 0.02fF
C1358 VPB.n856 VNB 0.01fF
C1359 VPB.n857 VNB 0.02fF
C1360 VPB.n858 VNB 0.28fF
C1361 VPB.n859 VNB 0.01fF
C1362 VPB.n860 VNB 0.02fF
C1363 VPB.n861 VNB 0.04fF
C1364 VPB.n862 VNB 0.04fF
C1365 VPB.n863 VNB 0.02fF
C1366 VPB.n864 VNB 0.02fF
C1367 VPB.n865 VNB 0.02fF
C1368 VPB.n866 VNB 0.02fF
C1369 VPB.n867 VNB 0.02fF
C1370 VPB.n868 VNB 0.02fF
C1371 VPB.n869 VNB 0.02fF
C1372 VPB.n870 VNB 0.02fF
C1373 VPB.n871 VNB 0.02fF
C1374 VPB.n872 VNB 0.02fF
C1375 VPB.n873 VNB 0.02fF
C1376 VPB.n874 VNB 0.28fF
C1377 VPB.n875 VNB 0.01fF
C1378 VPB.n876 VNB 0.02fF
C1379 VPB.n877 VNB 0.03fF
C1380 VPB.n878 VNB 0.03fF
C1381 VPB.n879 VNB 0.28fF
C1382 VPB.n880 VNB 0.01fF
C1383 VPB.n881 VNB 0.02fF
C1384 VPB.n882 VNB 0.03fF
C1385 VPB.n883 VNB 0.28fF
C1386 VPB.n884 VNB 0.02fF
C1387 VPB.n885 VNB 0.02fF
C1388 VPB.n886 VNB 0.02fF
C1389 VPB.n887 VNB 0.05fF
C1390 VPB.n888 VNB 0.21fF
C1391 VPB.n889 VNB 0.02fF
C1392 VPB.n890 VNB 0.01fF
C1393 VPB.n891 VNB 0.02fF
C1394 VPB.n892 VNB 0.14fF
C1395 VPB.n893 VNB 0.16fF
C1396 VPB.n894 VNB 0.02fF
C1397 VPB.n895 VNB 0.02fF
C1398 VPB.n896 VNB 0.02fF
C1399 VPB.n897 VNB 0.10fF
C1400 VPB.n898 VNB 0.02fF
C1401 VPB.n899 VNB 0.14fF
C1402 VPB.n900 VNB 0.16fF
C1403 VPB.n901 VNB 0.02fF
C1404 VPB.n902 VNB 0.02fF
C1405 VPB.n903 VNB 0.02fF
C1406 VPB.n904 VNB 0.14fF
C1407 VPB.n905 VNB 0.15fF
C1408 VPB.n906 VNB 0.02fF
C1409 VPB.n907 VNB 0.02fF
C1410 VPB.n908 VNB 0.02fF
C1411 VPB.n909 VNB 0.14fF
C1412 VPB.n910 VNB 0.15fF
C1413 VPB.n911 VNB 0.02fF
C1414 VPB.n912 VNB 0.02fF
C1415 VPB.n913 VNB 0.02fF
C1416 VPB.n914 VNB 0.10fF
C1417 VPB.n915 VNB 0.02fF
C1418 VPB.n916 VNB 0.14fF
C1419 VPB.n917 VNB 0.16fF
C1420 VPB.n918 VNB 0.02fF
C1421 VPB.n919 VNB 0.02fF
C1422 VPB.n920 VNB 0.02fF
C1423 VPB.n921 VNB 0.14fF
C1424 VPB.n922 VNB 0.16fF
C1425 VPB.n923 VNB 0.02fF
C1426 VPB.n924 VNB 0.02fF
C1427 VPB.n925 VNB 0.02fF
C1428 VPB.n926 VNB 0.06fF
C1429 VPB.n927 VNB 0.21fF
C1430 VPB.n928 VNB 0.02fF
C1431 VPB.n929 VNB 0.01fF
C1432 VPB.n930 VNB 0.02fF
C1433 VPB.n931 VNB 0.28fF
C1434 VPB.n932 VNB 0.02fF
C1435 VPB.n933 VNB 0.02fF
C1436 VPB.n934 VNB 0.02fF
C1437 VPB.n935 VNB 0.28fF
C1438 VPB.n936 VNB 0.01fF
C1439 VPB.n937 VNB 0.02fF
C1440 VPB.n938 VNB 0.04fF
C1441 VPB.n939 VNB 0.02fF
C1442 VPB.n940 VNB 0.02fF
C1443 VPB.n941 VNB 0.02fF
C1444 VPB.n942 VNB 0.04fF
C1445 VPB.n943 VNB 0.02fF
C1446 VPB.n944 VNB 0.24fF
C1447 VPB.n945 VNB 0.04fF
C1448 VPB.n947 VNB 0.02fF
C1449 VPB.n948 VNB 0.02fF
C1450 VPB.n949 VNB 0.02fF
C1451 VPB.n950 VNB 0.02fF
C1452 VPB.n952 VNB 0.02fF
C1453 VPB.n953 VNB 0.02fF
C1454 VPB.n954 VNB 0.02fF
C1455 VPB.n956 VNB 0.28fF
C1456 VPB.n958 VNB 0.03fF
C1457 VPB.n959 VNB 0.02fF
C1458 VPB.n960 VNB 0.03fF
C1459 VPB.n961 VNB 0.03fF
C1460 VPB.n962 VNB 0.28fF
C1461 VPB.n963 VNB 0.01fF
C1462 VPB.n964 VNB 0.02fF
C1463 VPB.n965 VNB 0.04fF
C1464 VPB.n966 VNB 0.05fF
C1465 VPB.n967 VNB 0.23fF
C1466 VPB.n968 VNB 0.02fF
C1467 VPB.n969 VNB 0.01fF
C1468 VPB.n970 VNB 0.02fF
C1469 VPB.n971 VNB 0.14fF
C1470 VPB.n972 VNB 0.16fF
C1471 VPB.n973 VNB 0.02fF
C1472 VPB.n974 VNB 0.02fF
C1473 VPB.n975 VNB 0.02fF
C1474 VPB.n976 VNB 0.10fF
C1475 VPB.n977 VNB 0.02fF
C1476 VPB.n978 VNB 0.14fF
C1477 VPB.n979 VNB 0.15fF
C1478 VPB.n980 VNB 0.02fF
C1479 VPB.n981 VNB 0.02fF
C1480 VPB.n982 VNB 0.02fF
C1481 VPB.n983 VNB 0.14fF
C1482 VPB.n984 VNB 0.15fF
C1483 VPB.n985 VNB 0.02fF
C1484 VPB.n986 VNB 0.02fF
C1485 VPB.n987 VNB 0.02fF
C1486 VPB.n988 VNB 0.14fF
C1487 VPB.n989 VNB 0.16fF
C1488 VPB.n990 VNB 0.02fF
C1489 VPB.n991 VNB 0.02fF
C1490 VPB.n992 VNB 0.02fF
C1491 VPB.n993 VNB 0.06fF
C1492 VPB.n994 VNB 0.24fF
C1493 VPB.n995 VNB 0.02fF
C1494 VPB.n996 VNB 0.01fF
C1495 VPB.n997 VNB 0.02fF
C1496 VPB.n998 VNB 0.28fF
C1497 VPB.n999 VNB 0.01fF
C1498 VPB.n1000 VNB 0.02fF
C1499 VPB.n1001 VNB 0.04fF
C1500 VPB.n1002 VNB 0.02fF
C1501 VPB.n1003 VNB 0.02fF
C1502 VPB.n1004 VNB 0.02fF
C1503 VPB.n1005 VNB 0.04fF
C1504 VPB.n1006 VNB 0.02fF
C1505 VPB.n1007 VNB 0.24fF
C1506 VPB.n1008 VNB 0.04fF
C1507 VPB.n1010 VNB 0.02fF
C1508 VPB.n1011 VNB 0.02fF
C1509 VPB.n1012 VNB 0.02fF
C1510 VPB.n1013 VNB 0.02fF
C1511 VPB.n1015 VNB 0.02fF
C1512 VPB.n1016 VNB 0.02fF
C1513 VPB.n1017 VNB 0.02fF
C1514 VPB.n1019 VNB 0.28fF
C1515 VPB.n1021 VNB 0.03fF
C1516 VPB.n1022 VNB 0.02fF
C1517 VPB.n1023 VNB 0.03fF
C1518 VPB.n1024 VNB 0.03fF
C1519 VPB.n1025 VNB 0.28fF
C1520 VPB.n1026 VNB 0.01fF
C1521 VPB.n1027 VNB 0.02fF
C1522 VPB.n1028 VNB 0.04fF
C1523 VPB.n1029 VNB 0.28fF
C1524 VPB.n1030 VNB 0.02fF
C1525 VPB.n1031 VNB 0.02fF
C1526 VPB.n1032 VNB 0.02fF
C1527 VPB.n1033 VNB 0.05fF
C1528 VPB.n1034 VNB 0.21fF
C1529 VPB.n1035 VNB 0.02fF
C1530 VPB.n1036 VNB 0.01fF
C1531 VPB.n1037 VNB 0.02fF
C1532 VPB.n1038 VNB 0.14fF
C1533 VPB.n1039 VNB 0.16fF
C1534 VPB.n1040 VNB 0.02fF
C1535 VPB.n1041 VNB 0.02fF
C1536 VPB.n1042 VNB 0.02fF
C1537 VPB.n1043 VNB 0.10fF
C1538 VPB.n1044 VNB 0.02fF
C1539 VPB.n1045 VNB 0.14fF
C1540 VPB.n1046 VNB 0.16fF
C1541 VPB.n1047 VNB 0.02fF
C1542 VPB.n1048 VNB 0.02fF
C1543 VPB.n1049 VNB 0.02fF
C1544 VPB.n1050 VNB 0.14fF
C1545 VPB.n1051 VNB 0.15fF
C1546 VPB.n1052 VNB 0.02fF
C1547 VPB.n1053 VNB 0.02fF
C1548 VPB.n1054 VNB 0.02fF
C1549 VPB.n1055 VNB 0.14fF
C1550 VPB.n1056 VNB 0.15fF
C1551 VPB.n1057 VNB 0.02fF
C1552 VPB.n1058 VNB 0.02fF
C1553 VPB.n1059 VNB 0.02fF
C1554 VPB.n1060 VNB 0.10fF
C1555 VPB.n1061 VNB 0.02fF
C1556 VPB.n1062 VNB 0.14fF
C1557 VPB.n1063 VNB 0.16fF
C1558 VPB.n1064 VNB 0.02fF
C1559 VPB.n1065 VNB 0.02fF
C1560 VPB.n1066 VNB 0.02fF
C1561 VPB.n1067 VNB 0.14fF
C1562 VPB.n1068 VNB 0.16fF
C1563 VPB.n1069 VNB 0.02fF
C1564 VPB.n1070 VNB 0.02fF
C1565 VPB.n1071 VNB 0.02fF
C1566 VPB.n1072 VNB 0.06fF
C1567 VPB.n1073 VNB 0.21fF
C1568 VPB.n1074 VNB 0.02fF
C1569 VPB.n1075 VNB 0.01fF
C1570 VPB.n1076 VNB 0.02fF
C1571 VPB.n1077 VNB 0.28fF
C1572 VPB.n1078 VNB 0.02fF
C1573 VPB.n1079 VNB 0.02fF
C1574 VPB.n1080 VNB 0.02fF
C1575 VPB.n1081 VNB 0.28fF
C1576 VPB.n1082 VNB 0.01fF
C1577 VPB.n1083 VNB 0.02fF
C1578 VPB.n1084 VNB 0.04fF
C1579 VPB.n1085 VNB 0.02fF
C1580 VPB.n1086 VNB 0.02fF
C1581 VPB.n1087 VNB 0.02fF
C1582 VPB.n1088 VNB 0.04fF
C1583 VPB.n1089 VNB 0.02fF
C1584 VPB.n1090 VNB 0.29fF
C1585 VPB.n1091 VNB 0.04fF
C1586 VPB.n1093 VNB 0.02fF
C1587 VPB.n1094 VNB 0.02fF
C1588 VPB.n1095 VNB 0.02fF
C1589 VPB.n1096 VNB 0.02fF
C1590 VPB.n1098 VNB 0.02fF
C1591 VPB.n1099 VNB 0.02fF
C1592 VPB.n1100 VNB 0.02fF
C1593 VPB.n1102 VNB 0.28fF
C1594 VPB.n1104 VNB 0.03fF
C1595 VPB.n1105 VNB 0.02fF
C1596 VPB.n1106 VNB 0.03fF
C1597 VPB.n1107 VNB 0.03fF
C1598 VPB.n1108 VNB 0.28fF
C1599 VPB.n1109 VNB 0.01fF
C1600 VPB.n1110 VNB 0.02fF
C1601 VPB.n1111 VNB 0.04fF
C1602 VPB.n1112 VNB 0.28fF
C1603 VPB.n1113 VNB 0.02fF
C1604 VPB.n1114 VNB 0.02fF
C1605 VPB.n1115 VNB 0.02fF
C1606 VPB.n1116 VNB 0.05fF
C1607 VPB.n1117 VNB 0.21fF
C1608 VPB.n1118 VNB 0.02fF
C1609 VPB.n1119 VNB 0.01fF
C1610 VPB.n1120 VNB 0.02fF
C1611 VPB.n1121 VNB 0.14fF
C1612 VPB.n1122 VNB 0.16fF
C1613 VPB.n1123 VNB 0.02fF
C1614 VPB.n1124 VNB 0.02fF
C1615 VPB.n1125 VNB 0.02fF
C1616 VPB.n1126 VNB 0.10fF
C1617 VPB.n1127 VNB 0.02fF
C1618 VPB.n1128 VNB 0.14fF
C1619 VPB.n1129 VNB 0.16fF
C1620 VPB.n1130 VNB 0.02fF
C1621 VPB.n1131 VNB 0.02fF
C1622 VPB.n1132 VNB 0.02fF
C1623 VPB.n1133 VNB 0.14fF
C1624 VPB.n1134 VNB 0.15fF
C1625 VPB.n1135 VNB 0.02fF
C1626 VPB.n1136 VNB 0.02fF
C1627 VPB.n1137 VNB 0.02fF
C1628 VPB.n1138 VNB 0.14fF
C1629 VPB.n1139 VNB 0.15fF
C1630 VPB.n1140 VNB 0.02fF
C1631 VPB.n1141 VNB 0.02fF
C1632 VPB.n1142 VNB 0.02fF
C1633 VPB.n1143 VNB 0.10fF
C1634 VPB.n1144 VNB 0.02fF
C1635 VPB.n1145 VNB 0.14fF
C1636 VPB.n1146 VNB 0.16fF
C1637 VPB.n1147 VNB 0.02fF
C1638 VPB.n1148 VNB 0.02fF
C1639 VPB.n1149 VNB 0.02fF
C1640 VPB.n1150 VNB 0.14fF
C1641 VPB.n1151 VNB 0.16fF
C1642 VPB.n1152 VNB 0.02fF
C1643 VPB.n1153 VNB 0.02fF
C1644 VPB.n1154 VNB 0.02fF
C1645 VPB.n1155 VNB 0.06fF
C1646 VPB.n1156 VNB 0.21fF
C1647 VPB.n1157 VNB 0.02fF
C1648 VPB.n1158 VNB 0.01fF
C1649 VPB.n1159 VNB 0.02fF
C1650 VPB.n1160 VNB 0.28fF
C1651 VPB.n1161 VNB 0.02fF
C1652 VPB.n1162 VNB 0.02fF
C1653 VPB.n1163 VNB 0.02fF
C1654 VPB.n1164 VNB 0.28fF
C1655 VPB.n1165 VNB 0.01fF
C1656 VPB.n1166 VNB 0.02fF
C1657 VPB.n1167 VNB 0.04fF
C1658 VPB.n1168 VNB 0.02fF
C1659 VPB.n1169 VNB 0.02fF
C1660 VPB.n1170 VNB 0.02fF
C1661 VPB.n1171 VNB 0.04fF
C1662 VPB.n1172 VNB 0.02fF
C1663 VPB.n1173 VNB 0.24fF
C1664 VPB.n1174 VNB 0.04fF
C1665 VPB.n1176 VNB 0.02fF
C1666 VPB.n1177 VNB 0.02fF
C1667 VPB.n1178 VNB 0.02fF
C1668 VPB.n1179 VNB 0.02fF
C1669 VPB.n1181 VNB 0.02fF
C1670 VPB.n1182 VNB 0.02fF
C1671 VPB.n1183 VNB 0.02fF
C1672 VPB.n1185 VNB 0.28fF
C1673 VPB.n1187 VNB 0.03fF
C1674 VPB.n1188 VNB 0.02fF
C1675 VPB.n1189 VNB 0.03fF
C1676 VPB.n1190 VNB 0.03fF
C1677 VPB.n1191 VNB 0.28fF
C1678 VPB.n1192 VNB 0.01fF
C1679 VPB.n1193 VNB 0.02fF
C1680 VPB.n1194 VNB 0.04fF
C1681 VPB.n1195 VNB 0.05fF
C1682 VPB.n1196 VNB 0.23fF
C1683 VPB.n1197 VNB 0.02fF
C1684 VPB.n1198 VNB 0.01fF
C1685 VPB.n1199 VNB 0.02fF
C1686 VPB.n1200 VNB 0.14fF
C1687 VPB.n1201 VNB 0.16fF
C1688 VPB.n1202 VNB 0.02fF
C1689 VPB.n1203 VNB 0.02fF
C1690 VPB.n1204 VNB 0.02fF
C1691 VPB.n1205 VNB 0.10fF
C1692 VPB.n1206 VNB 0.02fF
C1693 VPB.n1207 VNB 0.14fF
C1694 VPB.n1208 VNB 0.15fF
C1695 VPB.n1209 VNB 0.02fF
C1696 VPB.n1210 VNB 0.02fF
C1697 VPB.n1211 VNB 0.02fF
C1698 VPB.n1212 VNB 0.14fF
C1699 VPB.n1213 VNB 0.15fF
C1700 VPB.n1214 VNB 0.02fF
C1701 VPB.n1215 VNB 0.02fF
C1702 VPB.n1216 VNB 0.02fF
C1703 VPB.n1217 VNB 0.14fF
C1704 VPB.n1218 VNB 0.16fF
C1705 VPB.n1219 VNB 0.02fF
C1706 VPB.n1220 VNB 0.02fF
C1707 VPB.n1221 VNB 0.02fF
C1708 VPB.n1222 VNB 0.06fF
C1709 VPB.n1223 VNB 0.24fF
C1710 VPB.n1224 VNB 0.02fF
C1711 VPB.n1225 VNB 0.01fF
C1712 VPB.n1226 VNB 0.02fF
C1713 VPB.n1227 VNB 0.28fF
C1714 VPB.n1228 VNB 0.01fF
C1715 VPB.n1229 VNB 0.02fF
C1716 VPB.n1230 VNB 0.04fF
C1717 VPB.n1231 VNB 0.02fF
C1718 VPB.n1232 VNB 0.02fF
C1719 VPB.n1233 VNB 0.02fF
C1720 VPB.n1234 VNB 0.04fF
C1721 VPB.n1235 VNB 0.02fF
C1722 VPB.n1236 VNB 0.24fF
C1723 VPB.n1237 VNB 0.04fF
C1724 VPB.n1239 VNB 0.02fF
C1725 VPB.n1240 VNB 0.02fF
C1726 VPB.n1241 VNB 0.02fF
C1727 VPB.n1242 VNB 0.02fF
C1728 VPB.n1244 VNB 0.02fF
C1729 VPB.n1245 VNB 0.02fF
C1730 VPB.n1246 VNB 0.02fF
C1731 VPB.n1248 VNB 0.28fF
C1732 VPB.n1250 VNB 0.03fF
C1733 VPB.n1251 VNB 0.02fF
C1734 VPB.n1252 VNB 0.03fF
C1735 VPB.n1253 VNB 0.03fF
C1736 VPB.n1254 VNB 0.28fF
C1737 VPB.n1255 VNB 0.01fF
C1738 VPB.n1256 VNB 0.02fF
C1739 VPB.n1257 VNB 0.04fF
C1740 VPB.n1258 VNB 0.28fF
C1741 VPB.n1259 VNB 0.02fF
C1742 VPB.n1260 VNB 0.02fF
C1743 VPB.n1261 VNB 0.02fF
C1744 VPB.n1262 VNB 0.05fF
C1745 VPB.n1263 VNB 0.21fF
C1746 VPB.n1264 VNB 0.02fF
C1747 VPB.n1265 VNB 0.01fF
C1748 VPB.n1266 VNB 0.02fF
C1749 VPB.n1267 VNB 0.14fF
C1750 VPB.n1268 VNB 0.16fF
C1751 VPB.n1269 VNB 0.02fF
C1752 VPB.n1270 VNB 0.02fF
C1753 VPB.n1271 VNB 0.02fF
C1754 VPB.n1272 VNB 0.10fF
C1755 VPB.n1273 VNB 0.02fF
C1756 VPB.n1274 VNB 0.14fF
C1757 VPB.n1275 VNB 0.16fF
C1758 VPB.n1276 VNB 0.02fF
C1759 VPB.n1277 VNB 0.02fF
C1760 VPB.n1278 VNB 0.02fF
C1761 VPB.n1279 VNB 0.14fF
C1762 VPB.n1280 VNB 0.15fF
C1763 VPB.n1281 VNB 0.02fF
C1764 VPB.n1282 VNB 0.02fF
C1765 VPB.n1283 VNB 0.02fF
C1766 VPB.n1284 VNB 0.14fF
C1767 VPB.n1285 VNB 0.15fF
C1768 VPB.n1286 VNB 0.02fF
C1769 VPB.n1287 VNB 0.02fF
C1770 VPB.n1288 VNB 0.02fF
C1771 VPB.n1289 VNB 0.10fF
C1772 VPB.n1290 VNB 0.02fF
C1773 VPB.n1291 VNB 0.14fF
C1774 VPB.n1292 VNB 0.16fF
C1775 VPB.n1293 VNB 0.02fF
C1776 VPB.n1294 VNB 0.02fF
C1777 VPB.n1295 VNB 0.02fF
C1778 VPB.n1296 VNB 0.14fF
C1779 VPB.n1297 VNB 0.16fF
C1780 VPB.n1298 VNB 0.02fF
C1781 VPB.n1299 VNB 0.02fF
C1782 VPB.n1300 VNB 0.02fF
C1783 VPB.n1301 VNB 0.06fF
C1784 VPB.n1302 VNB 0.21fF
C1785 VPB.n1303 VNB 0.02fF
C1786 VPB.n1304 VNB 0.01fF
C1787 VPB.n1305 VNB 0.02fF
C1788 VPB.n1306 VNB 0.28fF
C1789 VPB.n1307 VNB 0.02fF
C1790 VPB.n1308 VNB 0.02fF
C1791 VPB.n1309 VNB 0.02fF
C1792 VPB.n1310 VNB 0.28fF
C1793 VPB.n1311 VNB 0.01fF
C1794 VPB.n1312 VNB 0.02fF
C1795 VPB.n1313 VNB 0.04fF
C1796 VPB.n1314 VNB 0.02fF
C1797 VPB.n1315 VNB 0.02fF
C1798 VPB.n1316 VNB 0.02fF
C1799 VPB.n1317 VNB 0.04fF
C1800 VPB.n1318 VNB 0.02fF
C1801 VPB.n1319 VNB 0.29fF
C1802 VPB.n1320 VNB 0.04fF
C1803 VPB.n1322 VNB 0.02fF
C1804 VPB.n1323 VNB 0.02fF
C1805 VPB.n1324 VNB 0.02fF
C1806 VPB.n1325 VNB 0.02fF
C1807 VPB.n1327 VNB 0.02fF
C1808 VPB.n1328 VNB 0.02fF
C1809 VPB.n1329 VNB 0.02fF
C1810 VPB.n1331 VNB 0.28fF
C1811 VPB.n1333 VNB 0.03fF
C1812 VPB.n1334 VNB 0.02fF
C1813 VPB.n1335 VNB 0.03fF
C1814 VPB.n1336 VNB 0.03fF
C1815 VPB.n1337 VNB 0.28fF
C1816 VPB.n1338 VNB 0.01fF
C1817 VPB.n1339 VNB 0.02fF
C1818 VPB.n1340 VNB 0.04fF
C1819 VPB.n1341 VNB 0.28fF
C1820 VPB.n1342 VNB 0.02fF
C1821 VPB.n1343 VNB 0.02fF
C1822 VPB.n1344 VNB 0.02fF
C1823 VPB.n1345 VNB 0.05fF
C1824 VPB.n1346 VNB 0.21fF
C1825 VPB.n1347 VNB 0.02fF
C1826 VPB.n1348 VNB 0.01fF
C1827 VPB.n1349 VNB 0.02fF
C1828 VPB.n1350 VNB 0.14fF
C1829 VPB.n1351 VNB 0.16fF
C1830 VPB.n1352 VNB 0.02fF
C1831 VPB.n1353 VNB 0.02fF
C1832 VPB.n1354 VNB 0.02fF
C1833 VPB.n1355 VNB 0.10fF
C1834 VPB.n1356 VNB 0.02fF
C1835 VPB.n1357 VNB 0.14fF
C1836 VPB.n1358 VNB 0.16fF
C1837 VPB.n1359 VNB 0.02fF
C1838 VPB.n1360 VNB 0.02fF
C1839 VPB.n1361 VNB 0.02fF
C1840 VPB.n1362 VNB 0.14fF
C1841 VPB.n1363 VNB 0.15fF
C1842 VPB.n1364 VNB 0.02fF
C1843 VPB.n1365 VNB 0.02fF
C1844 VPB.n1366 VNB 0.02fF
C1845 VPB.n1367 VNB 0.14fF
C1846 VPB.n1368 VNB 0.15fF
C1847 VPB.n1369 VNB 0.02fF
C1848 VPB.n1370 VNB 0.02fF
C1849 VPB.n1371 VNB 0.02fF
C1850 VPB.n1372 VNB 0.10fF
C1851 VPB.n1373 VNB 0.02fF
C1852 VPB.n1374 VNB 0.14fF
C1853 VPB.n1375 VNB 0.16fF
C1854 VPB.n1376 VNB 0.02fF
C1855 VPB.n1377 VNB 0.02fF
C1856 VPB.n1378 VNB 0.02fF
C1857 VPB.n1379 VNB 0.14fF
C1858 VPB.n1380 VNB 0.16fF
C1859 VPB.n1381 VNB 0.02fF
C1860 VPB.n1382 VNB 0.02fF
C1861 VPB.n1383 VNB 0.02fF
C1862 VPB.n1384 VNB 0.06fF
C1863 VPB.n1385 VNB 0.21fF
C1864 VPB.n1386 VNB 0.02fF
C1865 VPB.n1387 VNB 0.01fF
C1866 VPB.n1388 VNB 0.02fF
C1867 VPB.n1389 VNB 0.28fF
C1868 VPB.n1390 VNB 0.02fF
C1869 VPB.n1391 VNB 0.02fF
C1870 VPB.n1392 VNB 0.02fF
C1871 VPB.n1393 VNB 0.28fF
C1872 VPB.n1394 VNB 0.01fF
C1873 VPB.n1395 VNB 0.02fF
C1874 VPB.n1396 VNB 0.04fF
C1875 VPB.n1397 VNB 0.02fF
C1876 VPB.n1398 VNB 0.02fF
C1877 VPB.n1399 VNB 0.02fF
C1878 VPB.n1400 VNB 0.04fF
C1879 VPB.n1401 VNB 0.02fF
C1880 VPB.n1402 VNB 0.24fF
C1881 VPB.n1403 VNB 0.04fF
C1882 VPB.n1405 VNB 0.02fF
C1883 VPB.n1406 VNB 0.02fF
C1884 VPB.n1407 VNB 0.02fF
C1885 VPB.n1408 VNB 0.02fF
C1886 VPB.n1410 VNB 0.02fF
C1887 VPB.n1411 VNB 0.02fF
C1888 VPB.n1412 VNB 0.02fF
C1889 VPB.n1414 VNB 0.28fF
C1890 VPB.n1416 VNB 0.03fF
C1891 VPB.n1417 VNB 0.02fF
C1892 VPB.n1418 VNB 0.03fF
C1893 VPB.n1419 VNB 0.03fF
C1894 VPB.n1420 VNB 0.28fF
C1895 VPB.n1421 VNB 0.01fF
C1896 VPB.n1422 VNB 0.02fF
C1897 VPB.n1423 VNB 0.04fF
C1898 VPB.n1424 VNB 0.05fF
C1899 VPB.n1425 VNB 0.23fF
C1900 VPB.n1426 VNB 0.02fF
C1901 VPB.n1427 VNB 0.01fF
C1902 VPB.n1428 VNB 0.02fF
C1903 VPB.n1429 VNB 0.14fF
C1904 VPB.n1430 VNB 0.16fF
C1905 VPB.n1431 VNB 0.02fF
C1906 VPB.n1432 VNB 0.02fF
C1907 VPB.n1433 VNB 0.02fF
C1908 VPB.n1434 VNB 0.10fF
C1909 VPB.n1435 VNB 0.02fF
C1910 VPB.n1436 VNB 0.14fF
C1911 VPB.n1437 VNB 0.15fF
C1912 VPB.n1438 VNB 0.02fF
C1913 VPB.n1439 VNB 0.02fF
C1914 VPB.n1440 VNB 0.02fF
C1915 VPB.n1441 VNB 0.14fF
C1916 VPB.n1442 VNB 0.15fF
C1917 VPB.n1443 VNB 0.02fF
C1918 VPB.n1444 VNB 0.02fF
C1919 VPB.n1445 VNB 0.02fF
C1920 VPB.n1446 VNB 0.14fF
C1921 VPB.n1447 VNB 0.16fF
C1922 VPB.n1448 VNB 0.02fF
C1923 VPB.n1449 VNB 0.02fF
C1924 VPB.n1450 VNB 0.02fF
C1925 VPB.n1451 VNB 0.06fF
C1926 VPB.n1452 VNB 0.24fF
C1927 VPB.n1453 VNB 0.02fF
C1928 VPB.n1454 VNB 0.01fF
C1929 VPB.n1455 VNB 0.02fF
C1930 VPB.n1456 VNB 0.28fF
C1931 VPB.n1457 VNB 0.01fF
C1932 VPB.n1458 VNB 0.02fF
C1933 VPB.n1459 VNB 0.04fF
C1934 VPB.n1460 VNB 0.02fF
C1935 VPB.n1461 VNB 0.02fF
C1936 VPB.n1462 VNB 0.02fF
C1937 VPB.n1463 VNB 0.04fF
C1938 VPB.n1464 VNB 0.02fF
C1939 VPB.n1465 VNB 0.24fF
C1940 VPB.n1466 VNB 0.04fF
C1941 VPB.n1468 VNB 0.02fF
C1942 VPB.n1469 VNB 0.02fF
C1943 VPB.n1470 VNB 0.02fF
C1944 VPB.n1471 VNB 0.02fF
C1945 VPB.n1473 VNB 0.02fF
C1946 VPB.n1474 VNB 0.02fF
C1947 VPB.n1475 VNB 0.02fF
C1948 VPB.n1477 VNB 0.28fF
C1949 VPB.n1479 VNB 0.03fF
C1950 VPB.n1480 VNB 0.02fF
C1951 VPB.n1481 VNB 0.03fF
C1952 VPB.n1482 VNB 0.03fF
C1953 VPB.n1483 VNB 0.28fF
C1954 VPB.n1484 VNB 0.01fF
C1955 VPB.n1485 VNB 0.02fF
C1956 VPB.n1486 VNB 0.04fF
C1957 VPB.n1487 VNB 0.28fF
C1958 VPB.n1488 VNB 0.02fF
C1959 VPB.n1489 VNB 0.02fF
C1960 VPB.n1490 VNB 0.02fF
C1961 VPB.n1491 VNB 0.05fF
C1962 VPB.n1492 VNB 0.21fF
C1963 VPB.n1493 VNB 0.02fF
C1964 VPB.n1494 VNB 0.01fF
C1965 VPB.n1495 VNB 0.02fF
C1966 VPB.n1496 VNB 0.14fF
C1967 VPB.n1497 VNB 0.16fF
C1968 VPB.n1498 VNB 0.02fF
C1969 VPB.n1499 VNB 0.02fF
C1970 VPB.n1500 VNB 0.02fF
C1971 VPB.n1501 VNB 0.10fF
C1972 VPB.n1502 VNB 0.02fF
C1973 VPB.n1503 VNB 0.14fF
C1974 VPB.n1504 VNB 0.16fF
C1975 VPB.n1505 VNB 0.02fF
C1976 VPB.n1506 VNB 0.02fF
C1977 VPB.n1507 VNB 0.02fF
C1978 VPB.n1508 VNB 0.14fF
C1979 VPB.n1509 VNB 0.15fF
C1980 VPB.n1510 VNB 0.02fF
C1981 VPB.n1511 VNB 0.02fF
C1982 VPB.n1512 VNB 0.02fF
C1983 VPB.n1513 VNB 0.14fF
C1984 VPB.n1514 VNB 0.15fF
C1985 VPB.n1515 VNB 0.02fF
C1986 VPB.n1516 VNB 0.02fF
C1987 VPB.n1517 VNB 0.02fF
C1988 VPB.n1518 VNB 0.10fF
C1989 VPB.n1519 VNB 0.02fF
C1990 VPB.n1520 VNB 0.14fF
C1991 VPB.n1521 VNB 0.16fF
C1992 VPB.n1522 VNB 0.02fF
C1993 VPB.n1523 VNB 0.02fF
C1994 VPB.n1524 VNB 0.02fF
C1995 VPB.n1525 VNB 0.14fF
C1996 VPB.n1526 VNB 0.16fF
C1997 VPB.n1527 VNB 0.02fF
C1998 VPB.n1528 VNB 0.02fF
C1999 VPB.n1529 VNB 0.02fF
C2000 VPB.n1530 VNB 0.06fF
C2001 VPB.n1531 VNB 0.21fF
C2002 VPB.n1532 VNB 0.02fF
C2003 VPB.n1533 VNB 0.01fF
C2004 VPB.n1534 VNB 0.02fF
C2005 VPB.n1535 VNB 0.28fF
C2006 VPB.n1536 VNB 0.02fF
C2007 VPB.n1537 VNB 0.02fF
C2008 VPB.n1538 VNB 0.02fF
C2009 VPB.n1539 VNB 0.28fF
C2010 VPB.n1540 VNB 0.01fF
C2011 VPB.n1541 VNB 0.02fF
C2012 VPB.n1542 VNB 0.04fF
C2013 VPB.n1543 VNB 0.04fF
C2014 VPB.n1544 VNB 0.02fF
C2015 VPB.n1545 VNB 0.02fF
C2016 VPB.n1546 VNB 0.02fF
C2017 VPB.n1547 VNB 0.02fF
C2018 VPB.n1548 VNB 0.02fF
C2019 VPB.n1549 VNB 0.02fF
C2020 VPB.n1550 VNB 0.02fF
C2021 VPB.n1551 VNB 0.02fF
C2022 VPB.n1552 VNB 0.02fF
C2023 VPB.n1553 VNB 0.02fF
C2024 VPB.n1554 VNB 0.03fF
C2025 VPB.n1555 VNB 0.04fF
C2026 VPB.n1556 VNB 0.02fF
C2027 VPB.n1557 VNB 0.02fF
C2028 VPB.n1558 VNB 0.02fF
C2029 VPB.n1559 VNB 0.04fF
C2030 VPB.n1560 VNB 0.04fF
C2031 VPB.n1562 VNB 0.43fF
C2032 a_10507_159.n0 VNB 0.05fF
C2033 a_10507_159.n1 VNB 0.72fF
C2034 a_10507_159.n2 VNB 0.72fF
C2035 a_10507_159.n3 VNB 0.84fF
C2036 a_10507_159.n4 VNB 0.26fF
C2037 a_10507_159.n5 VNB 0.34fF
C2038 a_10507_159.n6 VNB 0.38fF
C2039 a_10507_159.t22 VNB 0.76fF
C2040 a_10507_159.n7 VNB 0.50fF
C2041 a_10507_159.n8 VNB 0.43fF
C2042 a_10507_159.n9 VNB 0.52fF
C2043 a_10507_159.n10 VNB 0.41fF
C2044 a_10507_159.n11 VNB 0.72fF
C2045 a_10507_159.n12 VNB 0.72fF
C2046 a_10507_159.n13 VNB 0.84fF
C2047 a_10507_159.n14 VNB 0.26fF
C2048 a_10507_159.n15 VNB 0.34fF
C2049 a_10507_159.n16 VNB 0.59fF
C2050 a_10507_159.n17 VNB 0.63fF
C2051 a_10507_159.n18 VNB 0.74fF
C2052 a_10507_159.n19 VNB 0.38fF
C2053 a_10507_159.t25 VNB 0.76fF
C2054 a_10507_159.n20 VNB 0.50fF
C2055 a_10507_159.n21 VNB 0.38fF
C2056 a_10507_159.n22 VNB 0.74fF
C2057 a_10507_159.n23 VNB 2.80fF
C2058 a_10507_159.n24 VNB 1.14fF
C2059 a_10507_159.n25 VNB 0.59fF
C2060 a_10507_159.n26 VNB 0.05fF
C2061 a_10507_159.n27 VNB 0.46fF
C2062 a_10507_159.n28 VNB 0.07fF
.ends
