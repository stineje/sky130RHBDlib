* SPICE3 file created from TIEHI.ext - technology: sky130A

.subckt TIEHI Y VDD GND
M1000 a_121_411# a_121_411# GND GND nshort w=3u l=0.15u
+  ad=0p pd=0u as=1.1408p ps=8.1u
M1001 Y a_121_411# VDD VDD pshort w=2u l=0.15u M=2
+  ad=0.58p pd=4.58u as=1.1p ps=9.1u
C0 a_121_411# Y 0.23fF
C1 VDD Y 0.76fF
C2 a_121_411# VDD 0.12fF
R0 VDD.n52 VDD.n51 13.653
R1 VDD.n51 VDD.n50 13.653
R2 VDD.n4 VDD.n2 12.915
R3 VDD.n4 VDD.n3 12.66
R4 VDD.n12 VDD.n11 12.343
R5 VDD.n10 VDD.n9 12.343
R6 VDD.n7 VDD.n6 12.343
R7 VDD.n35 VDD.n34 7.5
R8 VDD.n38 VDD.n37 7.5
R9 VDD.n40 VDD.n39 7.5
R10 VDD.n43 VDD.n42 7.5
R11 VDD.n49 VDD.n48 7.5
R12 VDD.n20 VDD.n16 7.5
R13 VDD.n2 VDD.n1 7.5
R14 VDD.n6 VDD.n5 7.5
R15 VDD.n9 VDD.n8 7.5
R16 VDD.n19 VDD.n18 7.5
R17 VDD.n14 VDD.n0 7.5
R18 VDD.n48 VDD.n47 6.772
R19 VDD.n36 VDD.n33 6.772
R20 VDD.n41 VDD.n38 6.772
R21 VDD.n45 VDD.n43 6.772
R22 VDD.n45 VDD.n44 6.772
R23 VDD.n41 VDD.n40 6.772
R24 VDD.n36 VDD.n35 6.772
R25 VDD.n47 VDD.n32 6.772
R26 VDD.n16 VDD.n15 6.458
R27 VDD.n28 VDD.n24 1.967
R28 VDD.n58 VDD.n57 1.967
R29 VDD.n14 VDD.n7 1.329
R30 VDD.n14 VDD.n10 1.329
R31 VDD.n14 VDD.n12 1.329
R32 VDD.n14 VDD.n13 1.329
R33 VDD.n15 VDD.n14 0.696
R34 VDD.n14 VDD.n4 0.696
R35 VDD.n46 VDD.n45 0.365
R36 VDD.n46 VDD.n41 0.365
R37 VDD.n46 VDD.n36 0.365
R38 VDD.n47 VDD.n46 0.365
R39 VDD.n53 VDD 0.207
R40 VDD.n63 VDD.n29 0.157
R41 VDD.n63 VDD.n59 0.157
R42 VDD.n59 VDD.n53 0.145
R43 Y.n1 Y.n0 192.895
R44 Y.n0 Y.t0 14.282
R45 Y.n0 Y.t1 14.282
R46 Y.n1 Y 0.046
C3 Y.t0 GND 0.14fF
C4 Y.t1 GND 0.14fF
C5 Y.n0 GND 0.74fF
C6 Y.n1 GND 0.11fF
C7 VDD.n0 GND 0.10fF
C8 VDD.n1 GND 0.02fF
C9 VDD.n2 GND 0.02fF
C10 VDD.n3 GND 0.04fF
C11 VDD.n4 GND 0.01fF
C12 VDD.n5 GND 0.02fF
C13 VDD.n6 GND 0.02fF
C14 VDD.n8 GND 0.02fF
C15 VDD.n9 GND 0.02fF
C16 VDD.n11 GND 0.02fF
C17 VDD.n14 GND 0.39fF
C18 VDD.n16 GND 0.03fF
C19 VDD.n18 GND 0.02fF
C20 VDD.n19 GND 0.02fF
C21 VDD.n20 GND 0.03fF
C22 VDD.n24 GND 0.05fF
C23 VDD.n28 GND 0.01fF
C24 VDD.n29 GND 0.06fF
C25 VDD.n32 GND 0.02fF
C26 VDD.n33 GND 0.02fF
C27 VDD.n34 GND 0.02fF
C28 VDD.n35 GND 0.02fF
C29 VDD.n37 GND 0.02fF
C30 VDD.n38 GND 0.02fF
C31 VDD.n39 GND 0.02fF
C32 VDD.n40 GND 0.02fF
C33 VDD.n42 GND 0.03fF
C34 VDD.n43 GND 0.02fF
C35 VDD.n44 GND 0.10fF
C36 VDD.n46 GND 0.39fF
C37 VDD.n48 GND 0.03fF
C38 VDD.n49 GND 0.03fF
C39 VDD.n50 GND 0.23fF
C40 VDD.n51 GND 0.02fF
C41 VDD.n52 GND 0.03fF
C42 VDD.n53 GND 0.02fF
C43 VDD.n57 GND 0.05fF
C44 VDD.n58 GND 0.01fF
C45 VDD.n59 GND 0.02fF
C46 VDD.n63 GND 0.02fF
.ends
