* SPICE3 file created from TMRDFFQNX1.ext - technology: sky130A

.subckt TMRDFFQNX1 QN D CLK VDD GND
X0 VDD CLK a_277_1004 VDD pshort w=2 l=0.15 M=2
X1 a_3177_1004 a_3303_383 a_3072_73 GND nshort w=3 l=0.15
X2 a_13757_1005 a_7595_383 QN VDD pshort w=2 l=0.15 M=2
X3 a_3177_1004 a_3303_383 VDD VDD pshort w=2 l=0.15 M=2
X4 a_4439_159 CLK a_6698_73 GND nshort w=3 l=0.15
X5 a_6137_1004 a_4439_159 a_6032_73 GND nshort w=3 l=0.15
X6 GND a_147_159 a_91_75 GND nshort w=3 l=0.15
X7 VDD CLK a_147_159 VDD pshort w=2 l=0.15 M=2
X8 a_8956_182 CLK a_8675_75 GND nshort w=3 l=0.15
X9 a_11887_383 a_8731_159 VDD VDD pshort w=2 l=0.15 M=2
X10 VDD a_11887_383 a_11761_1004 VDD pshort w=2 l=0.15 M=2
X11 QN a_7595_383 a_14320_73 GND nshort w=3 l=0.15
X12 GND a_8861_1004 a_11656_73 GND nshort w=3 l=0.15
X13 VDD CLK a_4439_159 VDD pshort w=2 l=0.15 M=2
X14 a_9183_943 D VDD VDD pshort w=2 l=0.15 M=2
X15 GND a_10429_1004 a_10990_73 GND nshort w=3 l=0.15
X16 GND a_4439_159 a_4383_75 GND nshort w=3 l=0.15
X17 a_3303_383 a_3177_1004 VDD VDD pshort w=2 l=0.15 M=2
X18 VDD a_599_943 a_277_1004 VDD pshort w=2 l=0.15 M=2
X19 VDD a_277_1004 a_599_943 VDD pshort w=2 l=0.15 M=2
X20 a_8731_159 a_10429_1004 VDD VDD pshort w=2 l=0.15 M=2
X21 a_4569_1004 a_4891_943 VDD VDD pshort w=2 l=0.15 M=2
X22 a_13757_1005 a_3303_383 QN VDD pshort w=2 l=0.15 M=2
X23 VDD a_147_159 a_3303_383 VDD pshort w=2 l=0.15 M=2
X24 VDD a_9183_943 a_10429_1004 VDD pshort w=2 l=0.15 M=2
X25 a_7595_383 a_7469_1004 VDD VDD pshort w=2 l=0.15 M=2
X26 VDD a_4569_1004 a_7469_1004 VDD pshort w=2 l=0.15 M=2
X27 a_1845_1004 a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X28 a_8861_1004 a_9183_943 VDD VDD pshort w=2 l=0.15 M=2
X29 VDD a_4439_159 a_4569_1004 VDD pshort w=2 l=0.15 M=2
X30 a_7595_383 a_4439_159 a_8030_73 GND nshort w=3 l=0.15
X31 GND a_4569_1004 a_5366_73 GND nshort w=3 l=0.15
X32 GND a_599_943 a_1740_73 GND nshort w=3 l=0.15
X33 a_6137_1004 a_4439_159 VDD VDD pshort w=2 l=0.15 M=2
X34 a_372_182 CLK a_91_75 GND nshort w=3 l=0.15
X35 a_9183_943 a_8861_1004 VDD VDD pshort w=2 l=0.15 M=2
X36 GND a_11887_383 a_13654_73 GND nshort w=3 l=0.15
X37 a_13093_1005 a_3303_383 a_13757_1005 VDD pshort w=2 l=0.15 M=2
X38 VDD a_7595_383 a_13093_1005 VDD pshort w=2 l=0.15 M=2
X39 GND a_11887_383 a_12988_73 GND nshort w=3 l=0.15
X40 VDD D a_599_943 VDD pshort w=2 l=0.15 M=2
X41 a_8731_159 CLK VDD VDD pshort w=2 l=0.15 M=2
X42 a_13757_1005 a_11887_383 a_13093_1005 VDD pshort w=2 l=0.15 M=2
X43 VDD a_8731_159 a_10429_1004 VDD pshort w=2 l=0.15 M=2
X44 a_147_159 CLK a_2406_73 GND nshort w=3 l=0.15
X45 a_4439_159 a_6137_1004 VDD VDD pshort w=2 l=0.15 M=2
X46 a_277_1004 a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X47 a_4664_182 CLK a_4383_75 GND nshort w=3 l=0.15
X48 VDD a_7595_383 a_7469_1004 VDD pshort w=2 l=0.15 M=2
X49 VDD CLK a_4569_1004 VDD pshort w=2 l=0.15 M=2
X50 a_9183_943 D a_9658_73 GND nshort w=3 l=0.15
X51 VDD a_599_943 a_1845_1004 VDD pshort w=2 l=0.15 M=2
X52 GND a_4569_1004 a_7364_73 GND nshort w=3 l=0.15
X53 GND a_3177_1004 a_3738_73 GND nshort w=3 l=0.15
X54 a_11761_1004 a_8861_1004 VDD VDD pshort w=2 l=0.15 M=2
X55 GND a_9183_943 a_10324_73 GND nshort w=3 l=0.15
X56 VDD a_11887_383 a_13093_1005 VDD pshort w=2 l=0.15 M=2
X57 a_4891_943 D VDD VDD pshort w=2 l=0.15 M=2
X58 a_8861_1004 a_9183_943 a_8956_182 GND nshort w=3 l=0.15
X59 a_11761_1004 a_11887_383 a_11656_73 GND nshort w=3 l=0.15
X60 GND a_277_1004 a_1074_73 GND nshort w=3 l=0.15
X61 VDD a_277_1004 a_3177_1004 VDD pshort w=2 l=0.15 M=2
X62 a_8731_159 CLK a_10990_73 GND nshort w=3 l=0.15
X63 VDD a_11761_1004 a_11887_383 VDD pshort w=2 l=0.15 M=2
X64 a_4891_943 a_4569_1004 VDD VDD pshort w=2 l=0.15 M=2
X65 a_1845_1004 a_147_159 a_1740_73 GND nshort w=3 l=0.15
X66 a_7595_383 a_4439_159 VDD VDD pshort w=2 l=0.15 M=2
X67 GND a_11761_1004 a_12322_73 GND nshort w=3 l=0.15
X68 a_8861_1004 a_8731_159 VDD VDD pshort w=2 l=0.15 M=2
X69 a_4891_943 D a_5366_73 GND nshort w=3 l=0.15
X70 a_147_159 a_1845_1004 VDD VDD pshort w=2 l=0.15 M=2
X71 VDD CLK a_8861_1004 VDD pshort w=2 l=0.15 M=2
X72 QN a_3303_383 a_13654_73 GND nshort w=3 l=0.15
X73 VDD a_4891_943 a_6137_1004 VDD pshort w=2 l=0.15 M=2
X74 GND a_6137_1004 a_6698_73 GND nshort w=3 l=0.15
X75 GND a_277_1004 a_3072_73 GND nshort w=3 l=0.15
X76 QN a_7595_383 a_12988_73 GND nshort w=3 l=0.15
X77 GND a_4891_943 a_6032_73 GND nshort w=3 l=0.15
X78 GND a_3303_383 a_14320_73 GND nshort w=3 l=0.15
X79 a_3303_383 a_147_159 a_3738_73 GND nshort w=3 l=0.15
X80 a_7469_1004 a_7595_383 a_7364_73 GND nshort w=3 l=0.15
X81 a_10429_1004 a_8731_159 a_10324_73 GND nshort w=3 l=0.15
X82 GND a_8731_159 a_8675_75 GND nshort w=3 l=0.15
X83 GND a_7469_1004 a_8030_73 GND nshort w=3 l=0.15
X84 a_599_943 D a_1074_73 GND nshort w=3 l=0.15
X85 a_11887_383 a_8731_159 a_12322_73 GND nshort w=3 l=0.15
X86 GND a_1845_1004 a_2406_73 GND nshort w=3 l=0.15
X87 a_277_1004 a_599_943 a_372_182 GND nshort w=3 l=0.15
X88 GND a_8861_1004 a_9658_73 GND nshort w=3 l=0.15
X89 a_4569_1004 a_4891_943 a_4664_182 GND nshort w=3 l=0.15
C0 VDD a_4439_159 3.02fF
C1 VDD a_4569_1004 2.49fF
C2 VDD a_8731_159 3.06fF
C3 a_147_159 CLK 4.49fF
C4 a_3303_383 D 7.42fF
C5 a_7595_383 D 2.68fF
C6 a_4439_159 CLK 4.81fF
C7 VDD a_8861_1004 2.49fF
C8 CLK a_8731_159 3.25fF
C9 VDD a_277_1004 2.32fF
C10 a_4439_159 a_4569_1004 3.00fF
C11 VDD a_11887_383 2.40fF
C12 VDD a_3303_383 2.61fF
C13 VDD a_7595_383 2.62fF
C14 VDD CLK 5.18fF
C15 a_147_159 a_277_1004 3.00fF
C16 a_3303_383 a_7595_383 2.76fF
C17 VDD a_147_159 3.05fF
C18 a_8861_1004 a_8731_159 3.00fF
C19 VDD GND 35.35fF
C20 a_7595_383 GND 2.22fF **FLOATING
C21 a_3303_383 GND 3.23fF **FLOATING
.ends
