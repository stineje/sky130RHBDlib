magic
tech sky130A
magscale 1 2
timestamp 1670369075
<< error_s >>
rect 198 296 214 312
rect 392 296 408 312
rect 586 296 602 312
rect 274 266 304 296
rect 468 266 498 296
rect 662 266 692 296
rect 198 250 214 266
rect 258 250 274 266
rect 393 252 408 266
rect 392 251 408 252
rect 452 252 467 266
rect 587 252 602 266
rect 452 251 468 252
rect 586 251 602 252
rect 646 252 661 266
rect 646 251 662 252
rect 391 250 392 251
rect 468 250 469 251
rect 585 250 586 251
rect 662 250 663 251
rect 198 165 214 181
rect 258 165 274 181
rect 392 165 408 181
rect 452 165 468 181
rect 586 165 602 181
rect 646 165 662 181
rect 168 135 198 165
rect 274 135 304 165
rect 362 135 392 165
rect 468 135 498 165
rect 556 135 586 165
rect 662 135 692 165
<< nwell >>
rect 87 786 953 1550
<< pwell >>
rect 34 34 632 544
rect 34 -34 928 34
<< pdiffc >>
rect 141 1331 175 1365
rect 229 1331 263 1365
rect 317 1331 351 1365
rect 493 1331 527 1365
rect 613 1331 647 1365
rect 789 1331 823 1365
rect 141 1059 175 1093
rect 317 1059 351 1093
rect 405 1059 439 1093
<< psubdiff >>
rect 34 482 928 544
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 928 17
rect 34 -34 928 -17
<< nsubdiff >>
rect 34 1497 928 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 928 1497
rect 34 822 928 884
<< psubdiffcont >>
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
<< poly >>
rect 619 944 659 974
rect 168 375 198 413
rect 362 382 392 383
rect 556 382 586 413
<< locali >>
rect 34 1497 928 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 928 1497
rect 34 1446 928 1463
rect 141 1365 175 1405
rect 141 1313 175 1331
rect 229 1365 263 1446
rect 229 1313 263 1331
rect 317 1365 527 1399
rect 317 1313 351 1331
rect 493 1313 527 1331
rect 613 1365 823 1399
rect 613 1297 647 1331
rect 789 1297 823 1331
rect 141 1093 175 1111
rect 317 1093 351 1111
rect 141 1025 351 1059
rect 405 1093 439 1111
rect 613 1059 647 1111
rect 405 1025 647 1059
rect 701 1059 735 1111
rect 701 1025 757 1059
rect 205 433 239 942
rect 353 908 361 942
rect 353 441 387 908
rect 353 433 357 441
rect 575 419 609 908
rect 723 348 757 1025
rect 219 314 757 348
rect 219 233 253 314
rect 413 233 447 314
rect 607 234 641 314
rect 122 34 156 73
rect 219 34 253 89
rect 316 34 350 73
rect 413 34 447 89
rect 510 34 544 73
rect 607 34 641 89
rect 704 34 738 89
rect 34 17 928 34
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 928 17
rect 34 -34 928 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
<< metal1 >>
rect 34 1497 928 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 928 1497
rect 34 1446 928 1463
rect 34 17 928 34
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 928 17
rect 34 -34 928 -17
use diff_ring_side  diff_ring_side_0
timestamp 1652319726
transform 1 0 962 0 1 0
box -87 -34 87 1550
use diff_ring_side  diff_ring_side_1
timestamp 1652319726
transform 1 0 0 0 1 0
box -87 -34 87 1550
use nmos_top_trim1  nmos_top_trim1_1
timestamp 1651256895
transform -1 0 360 0 1 73
box 0 0 248 309
use nmos_top_trim2  nmos_top_trim2_0
timestamp 1651256905
transform -1 0 554 0 1 73
box 0 0 248 309
use nmos_top_trim2  nmos_top_trim2_1
timestamp 1651256905
transform -1 0 748 0 1 73
box 0 0 248 309
use pmos2_1  pmos2_1_0
timestamp 1647326732
transform 1 0 43 0 1 1404
box 52 -460 352 37
use pmos2_1  pmos2_1_1
timestamp 1647326732
transform 1 0 219 0 1 1404
box 52 -460 352 37
use pmos2_1  pmos2_1_2
timestamp 1647326732
transform 1 0 515 0 1 1404
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 192 -1 0 942
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 223 -1 0 417
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 -1 369 1 0 415
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 378 -1 0 942
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_4
timestamp 1648060378
transform 0 -1 591 1 0 415
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_5
timestamp 1648060378
transform 0 1 593 -1 0 942
box -32 -28 34 26
<< end >>
