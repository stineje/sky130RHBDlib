// File: nmos_bottom.spi.NMOS_BOTTOM.pxi
// Created: Tue Oct 15 15:58:05 2024
// 
simulator lang=spectre
cc_1 ( noxref_1 noxref_2 ) capacitor c=0.0420464f //x=0.43 //y=0.5 //x2=0 //y2=0
cc_2 ( noxref_1 noxref_3 ) capacitor c=0.0170906f //x=0.43 //y=0.5 //x2=0.62 \
 //y2=0.925
cc_3 ( noxref_2 noxref_3 ) capacitor c=0.106466f //x=0 //y=0 //x2=0.62 \
 //y2=0.925
