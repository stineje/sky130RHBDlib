magic
tech sky130A
magscale 1 2
timestamp 1670369097
<< error_s >>
rect -98 296 -82 312
rect 96 296 112 312
rect 290 296 306 312
rect 851 297 867 313
rect -22 266 8 296
rect 172 266 202 296
rect 366 266 396 296
rect 927 267 957 297
rect -98 250 -82 266
rect -38 250 -22 266
rect 97 252 112 266
rect 96 251 112 252
rect 156 252 171 266
rect 291 252 306 266
rect 156 251 172 252
rect 290 251 306 252
rect 350 252 365 266
rect 350 251 366 252
rect 851 251 867 267
rect 911 251 927 267
rect 95 250 96 251
rect 172 250 173 251
rect 289 250 290 251
rect 366 250 367 251
rect -98 165 -82 181
rect -38 165 -22 181
rect 96 165 112 181
rect 156 165 172 181
rect 290 165 306 181
rect 350 165 366 181
rect 851 166 867 182
rect 911 166 927 182
rect -128 135 -98 165
rect -22 135 8 165
rect 66 135 96 165
rect 172 135 202 165
rect 260 135 290 165
rect 366 135 396 165
rect 821 136 851 166
rect 927 136 957 166
<< metal1 >>
rect 491 649 761 683
use invx1_pcell  invx1_pcell_0
timestamp 1652329846
transform 1 0 666 0 1 0
box -87 -34 531 1550
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 444 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 814 0 1 666
box -53 -33 29 33
use nor3x1_pcell  nor3x1_pcell_0
timestamp 1670369075
transform 1 0 -296 0 1 0
box -87 -34 1049 1550
<< end >>
