// File: AND3X1.spi.AND3X1.pxi
// Created: Tue Oct 15 15:44:31 2024
// 
simulator lang=spectre
x_PM_AND3X1\%GND ( GND N_GND_c_4_p N_GND_c_31_p N_GND_c_1_p N_GND_c_5_p \
 N_GND_c_6_p N_GND_c_73_p N_GND_c_7_p N_GND_c_22_p N_GND_c_2_p N_GND_c_3_p \
 N_GND_M0_noxref_d N_GND_M3_noxref_s )  PM_AND3X1\%GND
x_PM_AND3X1\%VDD ( VDD N_VDD_c_92_p N_VDD_c_89_n N_VDD_c_97_p N_VDD_c_98_p \
 N_VDD_c_104_p N_VDD_c_108_p N_VDD_c_115_p N_VDD_c_90_n N_VDD_c_91_n \
 N_VDD_M4_noxref_s N_VDD_M5_noxref_d N_VDD_M7_noxref_d N_VDD_M9_noxref_d \
 N_VDD_M10_noxref_s N_VDD_M11_noxref_d )  PM_AND3X1\%VDD
x_PM_AND3X1\%noxref_3 ( N_noxref_3_c_172_n N_noxref_3_c_178_n \
 N_noxref_3_c_202_n N_noxref_3_c_206_n N_noxref_3_c_208_n N_noxref_3_c_212_n \
 N_noxref_3_c_179_n N_noxref_3_c_285_p N_noxref_3_c_216_n N_noxref_3_c_181_n \
 N_noxref_3_c_257_p N_noxref_3_c_263_p N_noxref_3_M3_noxref_g \
 N_noxref_3_M10_noxref_g N_noxref_3_M11_noxref_g N_noxref_3_c_186_n \
 N_noxref_3_c_301_p N_noxref_3_c_302_p N_noxref_3_c_188_n N_noxref_3_c_226_n \
 N_noxref_3_c_227_n N_noxref_3_c_189_n N_noxref_3_c_293_p N_noxref_3_c_190_n \
 N_noxref_3_c_192_n N_noxref_3_c_193_n N_noxref_3_M2_noxref_d \
 N_noxref_3_M4_noxref_d N_noxref_3_M6_noxref_d N_noxref_3_M8_noxref_d )  \
 PM_AND3X1\%noxref_3
x_PM_AND3X1\%A ( A A A A A A A N_A_c_313_n N_A_M0_noxref_g N_A_M4_noxref_g \
 N_A_M5_noxref_g N_A_c_314_n N_A_c_316_n N_A_c_317_n N_A_c_318_n N_A_c_319_n \
 N_A_c_320_n N_A_c_321_n N_A_c_323_n N_A_c_336_n N_A_c_331_n )  PM_AND3X1\%A
x_PM_AND3X1\%B ( B B B B B B B N_B_c_368_n N_B_M1_noxref_g N_B_M6_noxref_g \
 N_B_M7_noxref_g N_B_c_390_n N_B_c_393_n N_B_c_426_p N_B_c_433_p N_B_c_395_n \
 N_B_c_396_n N_B_c_397_n N_B_c_398_n N_B_c_381_n N_B_c_382_n )  PM_AND3X1\%B
x_PM_AND3X1\%noxref_6 ( N_noxref_6_c_457_n N_noxref_6_c_438_n \
 N_noxref_6_c_442_n N_noxref_6_c_446_n N_noxref_6_c_469_n \
 N_noxref_6_M0_noxref_s )  PM_AND3X1\%noxref_6
x_PM_AND3X1\%C ( C C C C C C C N_C_c_483_n N_C_M2_noxref_g N_C_M8_noxref_g \
 N_C_M9_noxref_g N_C_c_497_n N_C_c_498_n N_C_c_499_n N_C_c_500_n N_C_c_501_n \
 N_C_c_503_n N_C_c_504_n N_C_c_506_n N_C_c_507_n N_C_c_509_n )  PM_AND3X1\%C
x_PM_AND3X1\%noxref_8 ( N_noxref_8_c_537_n N_noxref_8_c_540_n \
 N_noxref_8_c_544_n N_noxref_8_c_547_n N_noxref_8_c_558_n \
 N_noxref_8_M1_noxref_d N_noxref_8_M2_noxref_s )  PM_AND3X1\%noxref_8
x_PM_AND3X1\%Y ( Y Y Y Y Y Y Y N_Y_c_592_n N_Y_c_616_n N_Y_c_602_n N_Y_c_605_n \
 N_Y_M3_noxref_d N_Y_M10_noxref_d )  PM_AND3X1\%Y
cc_1 ( N_GND_c_1_p N_VDD_c_89_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_90_n ) capacitor c=0.00855708f //x=4.81 //y=0 \
 //x2=4.81 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_91_n ) capacitor c=0.00989031f //x=6.41 //y=0 \
 //x2=6.29 //y2=7.4
cc_4 ( N_GND_c_4_p N_noxref_3_c_172_n ) capacitor c=0.0116268f //x=6.29 //y=0 \
 //x2=5.435 //y2=3.33
cc_5 ( N_GND_c_5_p N_noxref_3_c_172_n ) capacitor c=0.0016229f //x=4.64 //y=0 \
 //x2=5.435 //y2=3.33
cc_6 ( N_GND_c_6_p N_noxref_3_c_172_n ) capacitor c=0.00110325f //x=5.355 \
 //y=0 //x2=5.435 //y2=3.33
cc_7 ( N_GND_c_7_p N_noxref_3_c_172_n ) capacitor c=2.76195e-19 //x=5.84 \
 //y=0.535 //x2=5.435 //y2=3.33
cc_8 ( N_GND_c_2_p N_noxref_3_c_172_n ) capacitor c=0.00820844f //x=4.81 //y=0 \
 //x2=5.435 //y2=3.33
cc_9 ( N_GND_M3_noxref_s N_noxref_3_c_172_n ) capacitor c=0.00164577f \
 //x=5.305 //y=0.37 //x2=5.435 //y2=3.33
cc_10 ( N_GND_c_4_p N_noxref_3_c_178_n ) capacitor c=0.00177092f //x=6.29 \
 //y=0 //x2=4.185 //y2=3.33
cc_11 ( N_GND_c_2_p N_noxref_3_c_179_n ) capacitor c=0.0458509f //x=4.81 //y=0 \
 //x2=3.985 //y2=1.665
cc_12 ( N_GND_M3_noxref_s N_noxref_3_c_179_n ) capacitor c=3.19788e-19 \
 //x=5.305 //y=0.37 //x2=3.985 //y2=1.665
cc_13 ( N_GND_c_4_p N_noxref_3_c_181_n ) capacitor c=0.00184963f //x=6.29 \
 //y=0 //x2=5.55 //y2=2.085
cc_14 ( N_GND_c_7_p N_noxref_3_c_181_n ) capacitor c=7.87839e-19 //x=5.84 \
 //y=0.535 //x2=5.55 //y2=2.085
cc_15 ( N_GND_c_2_p N_noxref_3_c_181_n ) capacitor c=0.029021f //x=4.81 //y=0 \
 //x2=5.55 //y2=2.085
cc_16 ( N_GND_c_3_p N_noxref_3_c_181_n ) capacitor c=0.00118981f //x=6.41 \
 //y=0 //x2=5.55 //y2=2.085
cc_17 ( N_GND_M3_noxref_s N_noxref_3_c_181_n ) capacitor c=0.0108503f \
 //x=5.305 //y=0.37 //x2=5.55 //y2=2.085
cc_18 ( N_GND_c_7_p N_noxref_3_c_186_n ) capacitor c=0.0121757f //x=5.84 \
 //y=0.535 //x2=5.66 //y2=0.91
cc_19 ( N_GND_M3_noxref_s N_noxref_3_c_186_n ) capacitor c=0.0318107f \
 //x=5.305 //y=0.37 //x2=5.66 //y2=0.91
cc_20 ( N_GND_c_2_p N_noxref_3_c_188_n ) capacitor c=0.00561485f //x=4.81 \
 //y=0 //x2=5.66 //y2=1.92
cc_21 ( N_GND_M3_noxref_s N_noxref_3_c_189_n ) capacitor c=0.00483274f \
 //x=5.305 //y=0.37 //x2=6.035 //y2=0.755
cc_22 ( N_GND_c_22_p N_noxref_3_c_190_n ) capacitor c=0.0118602f //x=6.325 \
 //y=0.535 //x2=6.19 //y2=0.91
cc_23 ( N_GND_M3_noxref_s N_noxref_3_c_190_n ) capacitor c=0.0143355f \
 //x=5.305 //y=0.37 //x2=6.19 //y2=0.91
cc_24 ( N_GND_M3_noxref_s N_noxref_3_c_192_n ) capacitor c=0.0074042f \
 //x=5.305 //y=0.37 //x2=6.19 //y2=1.255
cc_25 ( N_GND_c_7_p N_noxref_3_c_193_n ) capacitor c=2.1838e-19 //x=5.84 \
 //y=0.535 //x2=5.55 //y2=2.085
cc_26 ( N_GND_c_2_p N_noxref_3_c_193_n ) capacitor c=0.0108179f //x=4.81 //y=0 \
 //x2=5.55 //y2=2.085
cc_27 ( N_GND_M3_noxref_s N_noxref_3_c_193_n ) capacitor c=0.00655738f \
 //x=5.305 //y=0.37 //x2=5.55 //y2=2.085
cc_28 ( N_GND_c_2_p N_noxref_3_M2_noxref_d ) capacitor c=0.00591582f //x=4.81 \
 //y=0 //x2=3.395 //y2=0.915
cc_29 ( N_GND_M3_noxref_s N_noxref_3_M2_noxref_d ) capacitor c=2.07235e-19 \
 //x=5.305 //y=0.37 //x2=3.395 //y2=0.915
cc_30 ( N_GND_c_1_p N_A_c_313_n ) capacitor c=0.0180363f //x=0.74 //y=0 \
 //x2=1.11 //y2=2.08
cc_31 ( N_GND_c_31_p N_A_c_314_n ) capacitor c=0.00132755f //x=0.99 //y=0 \
 //x2=0.81 //y2=0.875
cc_32 ( N_GND_M0_noxref_d N_A_c_314_n ) capacitor c=0.00211996f //x=0.885 \
 //y=0.875 //x2=0.81 //y2=0.875
cc_33 ( N_GND_M0_noxref_d N_A_c_316_n ) capacitor c=0.00255985f //x=0.885 \
 //y=0.875 //x2=0.81 //y2=1.22
cc_34 ( N_GND_c_1_p N_A_c_317_n ) capacitor c=0.00295461f //x=0.74 //y=0 \
 //x2=0.81 //y2=1.53
cc_35 ( N_GND_c_1_p N_A_c_318_n ) capacitor c=0.0134214f //x=0.74 //y=0 \
 //x2=0.81 //y2=1.915
cc_36 ( N_GND_M0_noxref_d N_A_c_319_n ) capacitor c=0.0131341f //x=0.885 \
 //y=0.875 //x2=1.185 //y2=0.72
cc_37 ( N_GND_M0_noxref_d N_A_c_320_n ) capacitor c=0.00193146f //x=0.885 \
 //y=0.875 //x2=1.185 //y2=1.375
cc_38 ( N_GND_c_5_p N_A_c_321_n ) capacitor c=0.00129018f //x=4.64 //y=0 \
 //x2=1.34 //y2=0.875
cc_39 ( N_GND_M0_noxref_d N_A_c_321_n ) capacitor c=0.00257848f //x=0.885 \
 //y=0.875 //x2=1.34 //y2=0.875
cc_40 ( N_GND_M0_noxref_d N_A_c_323_n ) capacitor c=0.00255985f //x=0.885 \
 //y=0.875 //x2=1.34 //y2=1.22
cc_41 ( N_GND_c_1_p N_B_c_368_n ) capacitor c=7.64246e-19 //x=0.74 //y=0 \
 //x2=2.22 //y2=2.08
cc_42 ( N_GND_c_4_p N_noxref_6_c_438_n ) capacitor c=0.00710541f //x=6.29 \
 //y=0 //x2=1.475 //y2=1.59
cc_43 ( N_GND_c_31_p N_noxref_6_c_438_n ) capacitor c=0.00110021f //x=0.99 \
 //y=0 //x2=1.475 //y2=1.59
cc_44 ( N_GND_c_5_p N_noxref_6_c_438_n ) capacitor c=0.00179185f //x=4.64 \
 //y=0 //x2=1.475 //y2=1.59
cc_45 ( N_GND_M0_noxref_d N_noxref_6_c_438_n ) capacitor c=0.00900091f \
 //x=0.885 //y=0.875 //x2=1.475 //y2=1.59
cc_46 ( N_GND_c_4_p N_noxref_6_c_442_n ) capacitor c=0.00709506f //x=6.29 \
 //y=0 //x2=1.56 //y2=0.625
cc_47 ( N_GND_c_5_p N_noxref_6_c_442_n ) capacitor c=0.0140218f //x=4.64 //y=0 \
 //x2=1.56 //y2=0.625
cc_48 ( N_GND_c_3_p N_noxref_6_c_442_n ) capacitor c=0.00138062f //x=6.41 \
 //y=0 //x2=1.56 //y2=0.625
cc_49 ( N_GND_M0_noxref_d N_noxref_6_c_442_n ) capacitor c=0.033954f //x=0.885 \
 //y=0.875 //x2=1.56 //y2=0.625
cc_50 ( N_GND_c_4_p N_noxref_6_c_446_n ) capacitor c=0.0192401f //x=6.29 //y=0 \
 //x2=2.445 //y2=0.54
cc_51 ( N_GND_c_5_p N_noxref_6_c_446_n ) capacitor c=0.0356078f //x=4.64 //y=0 \
 //x2=2.445 //y2=0.54
cc_52 ( N_GND_c_3_p N_noxref_6_c_446_n ) capacitor c=0.00264707f //x=6.41 \
 //y=0 //x2=2.445 //y2=0.54
cc_53 ( N_GND_c_4_p N_noxref_6_M0_noxref_s ) capacitor c=0.0139221f //x=6.29 \
 //y=0 //x2=0.455 //y2=0.375
cc_54 ( N_GND_c_31_p N_noxref_6_M0_noxref_s ) capacitor c=0.0140218f //x=0.99 \
 //y=0 //x2=0.455 //y2=0.375
cc_55 ( N_GND_c_1_p N_noxref_6_M0_noxref_s ) capacitor c=0.0712607f //x=0.74 \
 //y=0 //x2=0.455 //y2=0.375
cc_56 ( N_GND_c_5_p N_noxref_6_M0_noxref_s ) capacitor c=0.0131422f //x=4.64 \
 //y=0 //x2=0.455 //y2=0.375
cc_57 ( N_GND_c_2_p N_noxref_6_M0_noxref_s ) capacitor c=3.31601e-19 //x=4.81 \
 //y=0 //x2=0.455 //y2=0.375
cc_58 ( N_GND_c_3_p N_noxref_6_M0_noxref_s ) capacitor c=0.00272322f //x=6.41 \
 //y=0 //x2=0.455 //y2=0.375
cc_59 ( N_GND_M0_noxref_d N_noxref_6_M0_noxref_s ) capacitor c=0.033718f \
 //x=0.885 //y=0.875 //x2=0.455 //y2=0.375
cc_60 ( N_GND_c_2_p N_C_c_483_n ) capacitor c=9.53263e-19 //x=4.81 //y=0 \
 //x2=3.33 //y2=2.08
cc_61 ( N_GND_c_4_p N_noxref_8_c_537_n ) capacitor c=0.00789826f //x=6.29 \
 //y=0 //x2=3.015 //y2=0.995
cc_62 ( N_GND_c_5_p N_noxref_8_c_537_n ) capacitor c=0.00829979f //x=4.64 \
 //y=0 //x2=3.015 //y2=0.995
cc_63 ( N_GND_c_3_p N_noxref_8_c_537_n ) capacitor c=3.53825e-19 //x=6.41 \
 //y=0 //x2=3.015 //y2=0.995
cc_64 ( N_GND_c_4_p N_noxref_8_c_540_n ) capacitor c=0.00709506f //x=6.29 \
 //y=0 //x2=3.1 //y2=0.625
cc_65 ( N_GND_c_5_p N_noxref_8_c_540_n ) capacitor c=0.0140218f //x=4.64 //y=0 \
 //x2=3.1 //y2=0.625
cc_66 ( N_GND_c_3_p N_noxref_8_c_540_n ) capacitor c=0.00138062f //x=6.41 \
 //y=0 //x2=3.1 //y2=0.625
cc_67 ( N_GND_M0_noxref_d N_noxref_8_c_540_n ) capacitor c=6.21394e-19 \
 //x=0.885 //y=0.875 //x2=3.1 //y2=0.625
cc_68 ( N_GND_c_4_p N_noxref_8_c_544_n ) capacitor c=0.018306f //x=6.29 //y=0 \
 //x2=3.985 //y2=0.54
cc_69 ( N_GND_c_5_p N_noxref_8_c_544_n ) capacitor c=0.0362762f //x=4.64 //y=0 \
 //x2=3.985 //y2=0.54
cc_70 ( N_GND_c_3_p N_noxref_8_c_544_n ) capacitor c=0.00282763f //x=6.41 \
 //y=0 //x2=3.985 //y2=0.54
cc_71 ( N_GND_c_4_p N_noxref_8_c_547_n ) capacitor c=0.00286759f //x=6.29 \
 //y=0 //x2=4.07 //y2=0.625
cc_72 ( N_GND_c_5_p N_noxref_8_c_547_n ) capacitor c=0.0142605f //x=4.64 //y=0 \
 //x2=4.07 //y2=0.625
cc_73 ( N_GND_c_73_p N_noxref_8_c_547_n ) capacitor c=9.29926e-19 //x=5.44 \
 //y=0.45 //x2=4.07 //y2=0.625
cc_74 ( N_GND_c_2_p N_noxref_8_c_547_n ) capacitor c=0.0404137f //x=4.81 //y=0 \
 //x2=4.07 //y2=0.625
cc_75 ( N_GND_c_3_p N_noxref_8_c_547_n ) capacitor c=0.0013725f //x=6.41 //y=0 \
 //x2=4.07 //y2=0.625
cc_76 ( N_GND_M0_noxref_d N_noxref_8_M1_noxref_d ) capacitor c=0.00162435f \
 //x=0.885 //y=0.875 //x2=1.86 //y2=0.91
cc_77 ( N_GND_c_1_p N_noxref_8_M2_noxref_s ) capacitor c=8.16352e-19 //x=0.74 \
 //y=0 //x2=2.965 //y2=0.375
cc_78 ( N_GND_c_2_p N_noxref_8_M2_noxref_s ) capacitor c=0.00183149f //x=4.81 \
 //y=0 //x2=2.965 //y2=0.375
cc_79 ( N_GND_M3_noxref_s N_noxref_8_M2_noxref_s ) capacitor c=9.29926e-19 \
 //x=5.305 //y=0.37 //x2=2.965 //y2=0.375
cc_80 ( N_GND_c_2_p Y ) capacitor c=8.10282e-19 //x=4.81 //y=0 //x2=6.29 \
 //y2=2.22
cc_81 ( N_GND_c_4_p N_Y_c_592_n ) capacitor c=0.00180637f //x=6.29 //y=0 \
 //x2=6.205 //y2=2.08
cc_82 ( N_GND_c_3_p N_Y_c_592_n ) capacitor c=0.0301661f //x=6.41 //y=0 \
 //x2=6.205 //y2=2.08
cc_83 ( N_GND_M3_noxref_s N_Y_c_592_n ) capacitor c=0.00999304f //x=5.305 \
 //y=0.37 //x2=6.205 //y2=2.08
cc_84 ( N_GND_c_4_p N_Y_M3_noxref_d ) capacitor c=0.00194883f //x=6.29 //y=0 \
 //x2=5.735 //y2=0.91
cc_85 ( N_GND_c_7_p N_Y_M3_noxref_d ) capacitor c=0.0146043f //x=5.84 \
 //y=0.535 //x2=5.735 //y2=0.91
cc_86 ( N_GND_c_2_p N_Y_M3_noxref_d ) capacitor c=0.00924905f //x=4.81 //y=0 \
 //x2=5.735 //y2=0.91
cc_87 ( N_GND_c_3_p N_Y_M3_noxref_d ) capacitor c=0.00973758f //x=6.41 //y=0 \
 //x2=5.735 //y2=0.91
cc_88 ( N_GND_M3_noxref_s N_Y_M3_noxref_d ) capacitor c=0.076995f //x=5.305 \
 //y=0.37 //x2=5.735 //y2=0.91
cc_89 ( N_VDD_c_92_p N_noxref_3_c_172_n ) capacitor c=0.00920603f //x=6.29 \
 //y=7.4 //x2=5.435 //y2=3.33
cc_90 ( N_VDD_c_90_n N_noxref_3_c_172_n ) capacitor c=0.0069465f //x=4.81 \
 //y=7.4 //x2=5.435 //y2=3.33
cc_91 ( N_VDD_M10_noxref_s N_noxref_3_c_172_n ) capacitor c=0.00106085f \
 //x=5.35 //y=5.02 //x2=5.435 //y2=3.33
cc_92 ( N_VDD_c_92_p N_noxref_3_c_178_n ) capacitor c=0.00163378f //x=6.29 \
 //y=7.4 //x2=4.185 //y2=3.33
cc_93 ( N_VDD_c_92_p N_noxref_3_c_202_n ) capacitor c=0.0059154f //x=6.29 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_94 ( N_VDD_c_97_p N_noxref_3_c_202_n ) capacitor c=4.18223e-19 //x=1.885 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_95 ( N_VDD_c_98_p N_noxref_3_c_202_n ) capacitor c=4.18223e-19 //x=2.765 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_96 ( N_VDD_M5_noxref_d N_noxref_3_c_202_n ) capacitor c=0.0119114f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_97 ( N_VDD_c_89_n N_noxref_3_c_206_n ) capacitor c=0.00880189f //x=0.74 \
 //y=7.4 //x2=1.615 //y2=5.155
cc_98 ( N_VDD_M4_noxref_s N_noxref_3_c_206_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_99 ( N_VDD_c_92_p N_noxref_3_c_208_n ) capacitor c=0.00593264f //x=6.29 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_100 ( N_VDD_c_98_p N_noxref_3_c_208_n ) capacitor c=4.18223e-19 //x=2.765 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_101 ( N_VDD_c_104_p N_noxref_3_c_208_n ) capacitor c=4.18223e-19 //x=3.645 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_102 ( N_VDD_M7_noxref_d N_noxref_3_c_208_n ) capacitor c=0.0119114f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_103 ( N_VDD_c_92_p N_noxref_3_c_212_n ) capacitor c=0.00592985f //x=6.29 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_104 ( N_VDD_c_104_p N_noxref_3_c_212_n ) capacitor c=6.98646e-19 //x=3.645 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_105 ( N_VDD_c_108_p N_noxref_3_c_212_n ) capacitor c=0.00179956f //x=4.64 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_106 ( N_VDD_M9_noxref_d N_noxref_3_c_212_n ) capacitor c=0.0119114f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_107 ( N_VDD_c_90_n N_noxref_3_c_216_n ) capacitor c=0.0456169f //x=4.81 \
 //y=7.4 //x2=4.07 //y2=3.33
cc_108 ( N_VDD_c_92_p N_noxref_3_c_181_n ) capacitor c=0.00160122f //x=6.29 \
 //y=7.4 //x2=5.55 //y2=2.085
cc_109 ( N_VDD_c_90_n N_noxref_3_c_181_n ) capacitor c=0.0272885f //x=4.81 \
 //y=7.4 //x2=5.55 //y2=2.085
cc_110 ( N_VDD_c_91_n N_noxref_3_c_181_n ) capacitor c=0.00144809f //x=6.29 \
 //y=7.4 //x2=5.55 //y2=2.085
cc_111 ( N_VDD_M10_noxref_s N_noxref_3_c_181_n ) capacitor c=0.00971593f \
 //x=5.35 //y=5.02 //x2=5.55 //y2=2.085
cc_112 ( N_VDD_c_115_p N_noxref_3_M10_noxref_g ) capacitor c=0.00748034f \
 //x=6.28 //y=7.4 //x2=5.705 //y2=6.02
cc_113 ( N_VDD_c_90_n N_noxref_3_M10_noxref_g ) capacitor c=0.00935943f \
 //x=4.81 //y=7.4 //x2=5.705 //y2=6.02
cc_114 ( N_VDD_M10_noxref_s N_noxref_3_M10_noxref_g ) capacitor c=0.0528676f \
 //x=5.35 //y=5.02 //x2=5.705 //y2=6.02
cc_115 ( N_VDD_c_115_p N_noxref_3_M11_noxref_g ) capacitor c=0.00697478f \
 //x=6.28 //y=7.4 //x2=6.145 //y2=6.02
cc_116 ( N_VDD_M11_noxref_d N_noxref_3_M11_noxref_g ) capacitor c=0.0528676f \
 //x=6.22 //y=5.02 //x2=6.145 //y2=6.02
cc_117 ( N_VDD_c_91_n N_noxref_3_c_226_n ) capacitor c=0.0287802f //x=6.29 \
 //y=7.4 //x2=6.07 //y2=4.79
cc_118 ( N_VDD_c_90_n N_noxref_3_c_227_n ) capacitor c=0.011132f //x=4.81 \
 //y=7.4 //x2=5.78 //y2=4.79
cc_119 ( N_VDD_M10_noxref_s N_noxref_3_c_227_n ) capacitor c=0.00527247f \
 //x=5.35 //y=5.02 //x2=5.78 //y2=4.79
cc_120 ( N_VDD_c_92_p N_noxref_3_M4_noxref_d ) capacitor c=0.00706456f \
 //x=6.29 //y=7.4 //x2=1.385 //y2=5.02
cc_121 ( N_VDD_c_97_p N_noxref_3_M4_noxref_d ) capacitor c=0.0138437f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_122 ( N_VDD_c_91_n N_noxref_3_M4_noxref_d ) capacitor c=0.00135292f \
 //x=6.29 //y=7.4 //x2=1.385 //y2=5.02
cc_123 ( N_VDD_M5_noxref_d N_noxref_3_M4_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_124 ( N_VDD_c_92_p N_noxref_3_M6_noxref_d ) capacitor c=0.00706456f \
 //x=6.29 //y=7.4 //x2=2.265 //y2=5.02
cc_125 ( N_VDD_c_98_p N_noxref_3_M6_noxref_d ) capacitor c=0.0138437f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_126 ( N_VDD_c_90_n N_noxref_3_M6_noxref_d ) capacitor c=4.9285e-19 //x=4.81 \
 //y=7.4 //x2=2.265 //y2=5.02
cc_127 ( N_VDD_c_91_n N_noxref_3_M6_noxref_d ) capacitor c=0.00135292f \
 //x=6.29 //y=7.4 //x2=2.265 //y2=5.02
cc_128 ( N_VDD_M4_noxref_s N_noxref_3_M6_noxref_d ) capacitor c=0.00130656f \
 //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_129 ( N_VDD_M5_noxref_d N_noxref_3_M6_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_130 ( N_VDD_M7_noxref_d N_noxref_3_M6_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_131 ( N_VDD_c_92_p N_noxref_3_M8_noxref_d ) capacitor c=0.00706456f \
 //x=6.29 //y=7.4 //x2=3.145 //y2=5.02
cc_132 ( N_VDD_c_104_p N_noxref_3_M8_noxref_d ) capacitor c=0.0137718f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_133 ( N_VDD_c_90_n N_noxref_3_M8_noxref_d ) capacitor c=0.00939849f \
 //x=4.81 //y=7.4 //x2=3.145 //y2=5.02
cc_134 ( N_VDD_c_91_n N_noxref_3_M8_noxref_d ) capacitor c=0.00135292f \
 //x=6.29 //y=7.4 //x2=3.145 //y2=5.02
cc_135 ( N_VDD_M7_noxref_d N_noxref_3_M8_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_136 ( N_VDD_M9_noxref_d N_noxref_3_M8_noxref_d ) capacitor c=0.0664752f \
 //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_137 ( N_VDD_M10_noxref_s N_noxref_3_M8_noxref_d ) capacitor c=5.22106e-19 \
 //x=5.35 //y=5.02 //x2=3.145 //y2=5.02
cc_138 ( N_VDD_c_92_p N_A_c_313_n ) capacitor c=0.00112336f //x=6.29 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_139 ( N_VDD_c_89_n N_A_c_313_n ) capacitor c=0.0168497f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_140 ( N_VDD_M4_noxref_s N_A_c_313_n ) capacitor c=0.0130213f //x=0.955 \
 //y=5.02 //x2=1.11 //y2=2.08
cc_141 ( N_VDD_c_97_p N_A_M4_noxref_g ) capacitor c=0.00749687f //x=1.885 \
 //y=7.4 //x2=1.31 //y2=6.02
cc_142 ( N_VDD_M4_noxref_s N_A_M4_noxref_g ) capacitor c=0.0477201f //x=0.955 \
 //y=5.02 //x2=1.31 //y2=6.02
cc_143 ( N_VDD_c_97_p N_A_M5_noxref_g ) capacitor c=0.00675175f //x=1.885 \
 //y=7.4 //x2=1.75 //y2=6.02
cc_144 ( N_VDD_M5_noxref_d N_A_M5_noxref_g ) capacitor c=0.015318f //x=1.825 \
 //y=5.02 //x2=1.75 //y2=6.02
cc_145 ( N_VDD_c_89_n N_A_c_331_n ) capacitor c=0.0076931f //x=0.74 //y=7.4 \
 //x2=1.385 //y2=4.79
cc_146 ( N_VDD_M4_noxref_s N_A_c_331_n ) capacitor c=0.00442959f //x=0.955 \
 //y=5.02 //x2=1.385 //y2=4.79
cc_147 ( N_VDD_c_92_p N_B_c_368_n ) capacitor c=2.41299e-19 //x=6.29 //y=7.4 \
 //x2=2.22 //y2=2.08
cc_148 ( N_VDD_c_89_n N_B_c_368_n ) capacitor c=7.34553e-19 //x=0.74 //y=7.4 \
 //x2=2.22 //y2=2.08
cc_149 ( N_VDD_c_98_p N_B_M6_noxref_g ) capacitor c=0.00676195f //x=2.765 \
 //y=7.4 //x2=2.19 //y2=6.02
cc_150 ( N_VDD_M5_noxref_d N_B_M6_noxref_g ) capacitor c=0.015318f //x=1.825 \
 //y=5.02 //x2=2.19 //y2=6.02
cc_151 ( N_VDD_c_98_p N_B_M7_noxref_g ) capacitor c=0.00675175f //x=2.765 \
 //y=7.4 //x2=2.63 //y2=6.02
cc_152 ( N_VDD_M7_noxref_d N_B_M7_noxref_g ) capacitor c=0.015318f //x=2.705 \
 //y=5.02 //x2=2.63 //y2=6.02
cc_153 ( N_VDD_c_90_n N_C_c_483_n ) capacitor c=8.81482e-19 //x=4.81 //y=7.4 \
 //x2=3.33 //y2=2.08
cc_154 ( N_VDD_c_104_p N_C_M8_noxref_g ) capacitor c=0.00675175f //x=3.645 \
 //y=7.4 //x2=3.07 //y2=6.02
cc_155 ( N_VDD_M7_noxref_d N_C_M8_noxref_g ) capacitor c=0.015318f //x=2.705 \
 //y=5.02 //x2=3.07 //y2=6.02
cc_156 ( N_VDD_c_104_p N_C_M9_noxref_g ) capacitor c=0.00675379f //x=3.645 \
 //y=7.4 //x2=3.51 //y2=6.02
cc_157 ( N_VDD_M9_noxref_d N_C_M9_noxref_g ) capacitor c=0.0394719f //x=3.585 \
 //y=5.02 //x2=3.51 //y2=6.02
cc_158 ( N_VDD_c_90_n Y ) capacitor c=4.80934e-19 //x=4.81 //y=7.4 //x2=6.29 \
 //y2=2.22
cc_159 ( N_VDD_c_91_n Y ) capacitor c=0.0232778f //x=6.29 //y=7.4 //x2=6.29 \
 //y2=2.22
cc_160 ( N_VDD_c_92_p N_Y_c_602_n ) capacitor c=0.00190861f //x=6.29 //y=7.4 \
 //x2=6.205 //y2=4.58
cc_161 ( N_VDD_c_115_p N_Y_c_602_n ) capacitor c=8.8179e-19 //x=6.28 //y=7.4 \
 //x2=6.205 //y2=4.58
cc_162 ( N_VDD_M11_noxref_d N_Y_c_602_n ) capacitor c=0.00641434f //x=6.22 \
 //y=5.02 //x2=6.205 //y2=4.58
cc_163 ( N_VDD_c_90_n N_Y_c_605_n ) capacitor c=0.017572f //x=4.81 //y=7.4 \
 //x2=6.01 //y2=4.58
cc_164 ( N_VDD_c_92_p N_Y_M10_noxref_d ) capacitor c=0.00708604f //x=6.29 \
 //y=7.4 //x2=5.78 //y2=5.02
cc_165 ( N_VDD_c_115_p N_Y_M10_noxref_d ) capacitor c=0.0139004f //x=6.28 \
 //y=7.4 //x2=5.78 //y2=5.02
cc_166 ( N_VDD_c_91_n N_Y_M10_noxref_d ) capacitor c=0.0219131f //x=6.29 \
 //y=7.4 //x2=5.78 //y2=5.02
cc_167 ( N_VDD_M10_noxref_s N_Y_M10_noxref_d ) capacitor c=0.0843065f //x=5.35 \
 //y=5.02 //x2=5.78 //y2=5.02
cc_168 ( N_VDD_M11_noxref_d N_Y_M10_noxref_d ) capacitor c=0.0832641f //x=6.22 \
 //y=5.02 //x2=5.78 //y2=5.02
cc_169 ( N_noxref_3_c_206_n N_A_M4_noxref_g ) capacitor c=0.0213876f //x=1.615 \
 //y=5.155 //x2=1.31 //y2=6.02
cc_170 ( N_noxref_3_c_202_n N_A_M5_noxref_g ) capacitor c=0.0204065f //x=2.325 \
 //y=5.155 //x2=1.75 //y2=6.02
cc_171 ( N_noxref_3_M4_noxref_d N_A_M5_noxref_g ) capacitor c=0.0180032f \
 //x=1.385 //y=5.02 //x2=1.75 //y2=6.02
cc_172 ( N_noxref_3_c_206_n N_A_c_336_n ) capacitor c=0.00437952f //x=1.615 \
 //y=5.155 //x2=1.675 //y2=4.79
cc_173 ( N_noxref_3_c_202_n N_B_c_368_n ) capacitor c=0.0149929f //x=2.325 \
 //y=5.155 //x2=2.22 //y2=2.08
cc_174 ( N_noxref_3_c_216_n N_B_c_368_n ) capacitor c=0.00326759f //x=4.07 \
 //y=3.33 //x2=2.22 //y2=2.08
cc_175 ( N_noxref_3_c_202_n N_B_M6_noxref_g ) capacitor c=0.0170029f //x=2.325 \
 //y=5.155 //x2=2.19 //y2=6.02
cc_176 ( N_noxref_3_M6_noxref_d N_B_M6_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.19 //y2=6.02
cc_177 ( N_noxref_3_c_208_n N_B_M7_noxref_g ) capacitor c=0.0209317f //x=3.205 \
 //y=5.155 //x2=2.63 //y2=6.02
cc_178 ( N_noxref_3_M6_noxref_d N_B_M7_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.63 //y2=6.02
cc_179 ( N_noxref_3_c_257_p N_B_c_381_n ) capacitor c=0.004361f //x=2.41 \
 //y=5.155 //x2=2.555 //y2=4.79
cc_180 ( N_noxref_3_c_202_n N_B_c_382_n ) capacitor c=0.0032428f //x=2.325 \
 //y=5.155 //x2=2.22 //y2=4.7
cc_181 ( N_noxref_3_M2_noxref_d N_noxref_6_M0_noxref_s ) capacitor \
 c=0.00309936f //x=3.395 //y=0.915 //x2=0.455 //y2=0.375
cc_182 ( N_noxref_3_c_178_n N_C_c_483_n ) capacitor c=0.00717888f //x=4.185 \
 //y=3.33 //x2=3.33 //y2=2.08
cc_183 ( N_noxref_3_c_216_n N_C_c_483_n ) capacitor c=0.0910677f //x=4.07 \
 //y=3.33 //x2=3.33 //y2=2.08
cc_184 ( N_noxref_3_c_181_n N_C_c_483_n ) capacitor c=0.00126776f //x=5.55 \
 //y=2.085 //x2=3.33 //y2=2.08
cc_185 ( N_noxref_3_c_263_p N_C_c_483_n ) capacitor c=0.0176831f //x=3.29 \
 //y=5.155 //x2=3.33 //y2=2.08
cc_186 ( N_noxref_3_c_208_n N_C_M8_noxref_g ) capacitor c=0.0209317f //x=3.205 \
 //y=5.155 //x2=3.07 //y2=6.02
cc_187 ( N_noxref_3_M8_noxref_d N_C_M8_noxref_g ) capacitor c=0.0180032f \
 //x=3.145 //y=5.02 //x2=3.07 //y2=6.02
cc_188 ( N_noxref_3_c_212_n N_C_M9_noxref_g ) capacitor c=0.0230698f //x=3.985 \
 //y=5.155 //x2=3.51 //y2=6.02
cc_189 ( N_noxref_3_M8_noxref_d N_C_M9_noxref_g ) capacitor c=0.0194246f \
 //x=3.145 //y=5.02 //x2=3.51 //y2=6.02
cc_190 ( N_noxref_3_M2_noxref_d N_C_c_497_n ) capacitor c=0.00217566f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=0.915
cc_191 ( N_noxref_3_M2_noxref_d N_C_c_498_n ) capacitor c=0.0034598f //x=3.395 \
 //y=0.915 //x2=3.32 //y2=1.26
cc_192 ( N_noxref_3_M2_noxref_d N_C_c_499_n ) capacitor c=0.00544291f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=1.57
cc_193 ( N_noxref_3_M2_noxref_d N_C_c_500_n ) capacitor c=0.00241102f \
 //x=3.395 //y=0.915 //x2=3.695 //y2=0.76
cc_194 ( N_noxref_3_c_179_n N_C_c_501_n ) capacitor c=0.00359704f //x=3.985 \
 //y=1.665 //x2=3.695 //y2=1.415
cc_195 ( N_noxref_3_M2_noxref_d N_C_c_501_n ) capacitor c=0.0140297f //x=3.395 \
 //y=0.915 //x2=3.695 //y2=1.415
cc_196 ( N_noxref_3_M2_noxref_d N_C_c_503_n ) capacitor c=0.00219619f \
 //x=3.395 //y=0.915 //x2=3.85 //y2=0.915
cc_197 ( N_noxref_3_c_179_n N_C_c_504_n ) capacitor c=0.00457401f //x=3.985 \
 //y=1.665 //x2=3.85 //y2=1.26
cc_198 ( N_noxref_3_M2_noxref_d N_C_c_504_n ) capacitor c=0.00603828f \
 //x=3.395 //y=0.915 //x2=3.85 //y2=1.26
cc_199 ( N_noxref_3_c_216_n N_C_c_506_n ) capacitor c=0.00877984f //x=4.07 \
 //y=3.33 //x2=3.33 //y2=2.08
cc_200 ( N_noxref_3_c_216_n N_C_c_507_n ) capacitor c=0.00283672f //x=4.07 \
 //y=3.33 //x2=3.33 //y2=1.915
cc_201 ( N_noxref_3_M2_noxref_d N_C_c_507_n ) capacitor c=0.00661782f \
 //x=3.395 //y=0.915 //x2=3.33 //y2=1.915
cc_202 ( N_noxref_3_c_212_n N_C_c_509_n ) capacitor c=0.00201851f //x=3.985 \
 //y=5.155 //x2=3.33 //y2=4.7
cc_203 ( N_noxref_3_c_216_n N_C_c_509_n ) capacitor c=0.013844f //x=4.07 \
 //y=3.33 //x2=3.33 //y2=4.7
cc_204 ( N_noxref_3_c_263_p N_C_c_509_n ) capacitor c=0.00475314f //x=3.29 \
 //y=5.155 //x2=3.33 //y2=4.7
cc_205 ( N_noxref_3_c_179_n N_noxref_8_c_544_n ) capacitor c=0.00469128f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_206 ( N_noxref_3_M2_noxref_d N_noxref_8_c_544_n ) capacitor c=0.0118457f \
 //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_207 ( N_noxref_3_c_285_p N_noxref_8_c_558_n ) capacitor c=0.0200405f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_208 ( N_noxref_3_M2_noxref_d N_noxref_8_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_209 ( N_noxref_3_c_179_n N_noxref_8_M2_noxref_s ) capacitor c=0.020752f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_210 ( N_noxref_3_M2_noxref_d N_noxref_8_M2_noxref_s ) capacitor \
 c=0.0426368f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
cc_211 ( N_noxref_3_c_172_n Y ) capacitor c=0.00582634f //x=5.435 //y=3.33 \
 //x2=6.29 //y2=2.22
cc_212 ( N_noxref_3_c_216_n Y ) capacitor c=0.00126776f //x=4.07 //y=3.33 \
 //x2=6.29 //y2=2.22
cc_213 ( N_noxref_3_c_181_n Y ) capacitor c=0.0711303f //x=5.55 //y=2.085 \
 //x2=6.29 //y2=2.22
cc_214 ( N_noxref_3_c_193_n Y ) capacitor c=8.49451e-19 //x=5.55 //y=2.085 \
 //x2=6.29 //y2=2.22
cc_215 ( N_noxref_3_c_293_p N_Y_c_592_n ) capacitor c=0.0023507f //x=6.035 \
 //y=1.41 //x2=6.205 //y2=2.08
cc_216 ( N_noxref_3_c_193_n N_Y_c_616_n ) capacitor c=0.0167852f //x=5.55 \
 //y=2.085 //x2=6.005 //y2=2.08
cc_217 ( N_noxref_3_c_226_n N_Y_c_602_n ) capacitor c=0.0101013f //x=6.07 \
 //y=4.79 //x2=6.205 //y2=4.58
cc_218 ( N_noxref_3_c_181_n N_Y_c_605_n ) capacitor c=0.0250789f //x=5.55 \
 //y=2.085 //x2=6.01 //y2=4.58
cc_219 ( N_noxref_3_c_227_n N_Y_c_605_n ) capacitor c=0.00962086f //x=5.78 \
 //y=4.79 //x2=6.01 //y2=4.58
cc_220 ( N_noxref_3_c_216_n N_Y_M3_noxref_d ) capacitor c=3.36976e-19 //x=4.07 \
 //y=3.33 //x2=5.735 //y2=0.91
cc_221 ( N_noxref_3_c_181_n N_Y_M3_noxref_d ) capacitor c=0.0175773f //x=5.55 \
 //y=2.085 //x2=5.735 //y2=0.91
cc_222 ( N_noxref_3_c_186_n N_Y_M3_noxref_d ) capacitor c=0.00218556f //x=5.66 \
 //y=0.91 //x2=5.735 //y2=0.91
cc_223 ( N_noxref_3_c_301_p N_Y_M3_noxref_d ) capacitor c=0.00347355f //x=5.66 \
 //y=1.255 //x2=5.735 //y2=0.91
cc_224 ( N_noxref_3_c_302_p N_Y_M3_noxref_d ) capacitor c=0.00742431f //x=5.66 \
 //y=1.565 //x2=5.735 //y2=0.91
cc_225 ( N_noxref_3_c_188_n N_Y_M3_noxref_d ) capacitor c=0.00957707f //x=5.66 \
 //y=1.92 //x2=5.735 //y2=0.91
cc_226 ( N_noxref_3_c_189_n N_Y_M3_noxref_d ) capacitor c=0.00220879f \
 //x=6.035 //y=0.755 //x2=5.735 //y2=0.91
cc_227 ( N_noxref_3_c_293_p N_Y_M3_noxref_d ) capacitor c=0.0138447f //x=6.035 \
 //y=1.41 //x2=5.735 //y2=0.91
cc_228 ( N_noxref_3_c_190_n N_Y_M3_noxref_d ) capacitor c=0.00218624f //x=6.19 \
 //y=0.91 //x2=5.735 //y2=0.91
cc_229 ( N_noxref_3_c_192_n N_Y_M3_noxref_d ) capacitor c=0.00601286f //x=6.19 \
 //y=1.255 //x2=5.735 //y2=0.91
cc_230 ( N_noxref_3_c_216_n N_Y_M10_noxref_d ) capacitor c=6.5427e-19 //x=4.07 \
 //y=3.33 //x2=5.78 //y2=5.02
cc_231 ( N_noxref_3_M10_noxref_g N_Y_M10_noxref_d ) capacitor c=0.0219309f \
 //x=5.705 //y=6.02 //x2=5.78 //y2=5.02
cc_232 ( N_noxref_3_M11_noxref_g N_Y_M10_noxref_d ) capacitor c=0.021902f \
 //x=6.145 //y=6.02 //x2=5.78 //y2=5.02
cc_233 ( N_noxref_3_c_226_n N_Y_M10_noxref_d ) capacitor c=0.0148755f //x=6.07 \
 //y=4.79 //x2=5.78 //y2=5.02
cc_234 ( N_noxref_3_c_227_n N_Y_M10_noxref_d ) capacitor c=0.00307344f \
 //x=5.78 //y=4.79 //x2=5.78 //y2=5.02
cc_235 ( N_A_c_313_n N_B_c_368_n ) capacitor c=0.0585104f //x=1.11 //y=2.08 \
 //x2=2.22 //y2=2.08
cc_236 ( N_A_c_318_n N_B_c_368_n ) capacitor c=0.00238338f //x=0.81 //y=1.915 \
 //x2=2.22 //y2=2.08
cc_237 ( N_A_c_336_n N_B_c_368_n ) capacitor c=0.00147352f //x=1.675 //y=4.79 \
 //x2=2.22 //y2=2.08
cc_238 ( N_A_c_331_n N_B_c_368_n ) capacitor c=0.00142741f //x=1.385 //y=4.79 \
 //x2=2.22 //y2=2.08
cc_239 ( N_A_M4_noxref_g N_B_M6_noxref_g ) capacitor c=0.0105869f //x=1.31 \
 //y=6.02 //x2=2.19 //y2=6.02
cc_240 ( N_A_M5_noxref_g N_B_M6_noxref_g ) capacitor c=0.10632f //x=1.75 \
 //y=6.02 //x2=2.19 //y2=6.02
cc_241 ( N_A_M5_noxref_g N_B_M7_noxref_g ) capacitor c=0.0101598f //x=1.75 \
 //y=6.02 //x2=2.63 //y2=6.02
cc_242 ( N_A_c_314_n N_B_c_390_n ) capacitor c=5.72482e-19 //x=0.81 //y=0.875 \
 //x2=1.785 //y2=0.91
cc_243 ( N_A_c_316_n N_B_c_390_n ) capacitor c=0.00149976f //x=0.81 //y=1.22 \
 //x2=1.785 //y2=0.91
cc_244 ( N_A_c_321_n N_B_c_390_n ) capacitor c=0.0160123f //x=1.34 //y=0.875 \
 //x2=1.785 //y2=0.91
cc_245 ( N_A_c_317_n N_B_c_393_n ) capacitor c=0.00111227f //x=0.81 //y=1.53 \
 //x2=1.785 //y2=1.22
cc_246 ( N_A_c_323_n N_B_c_393_n ) capacitor c=0.0124075f //x=1.34 //y=1.22 \
 //x2=1.785 //y2=1.22
cc_247 ( N_A_c_321_n N_B_c_395_n ) capacitor c=0.00103227f //x=1.34 //y=0.875 \
 //x2=2.31 //y2=0.91
cc_248 ( N_A_c_323_n N_B_c_396_n ) capacitor c=0.0010154f //x=1.34 //y=1.22 \
 //x2=2.31 //y2=1.22
cc_249 ( N_A_c_323_n N_B_c_397_n ) capacitor c=9.23422e-19 //x=1.34 //y=1.22 \
 //x2=2.31 //y2=1.45
cc_250 ( N_A_c_313_n N_B_c_398_n ) capacitor c=0.00231304f //x=1.11 //y=2.08 \
 //x2=2.31 //y2=1.915
cc_251 ( N_A_c_318_n N_B_c_398_n ) capacitor c=0.00964411f //x=0.81 //y=1.915 \
 //x2=2.31 //y2=1.915
cc_252 ( N_A_c_313_n N_B_c_382_n ) capacitor c=0.00183762f //x=1.11 //y=2.08 \
 //x2=2.22 //y2=4.7
cc_253 ( N_A_c_336_n N_B_c_382_n ) capacitor c=0.0168581f //x=1.675 //y=4.79 \
 //x2=2.22 //y2=4.7
cc_254 ( N_A_c_331_n N_B_c_382_n ) capacitor c=0.00484466f //x=1.385 //y=4.79 \
 //x2=2.22 //y2=4.7
cc_255 ( N_A_c_318_n N_noxref_6_c_457_n ) capacitor c=0.0034165f //x=0.81 \
 //y=1.915 //x2=0.59 //y2=1.505
cc_256 ( N_A_c_313_n N_noxref_6_c_438_n ) capacitor c=0.0122915f //x=1.11 \
 //y=2.08 //x2=1.475 //y2=1.59
cc_257 ( N_A_c_317_n N_noxref_6_c_438_n ) capacitor c=0.00703864f //x=0.81 \
 //y=1.53 //x2=1.475 //y2=1.59
cc_258 ( N_A_c_318_n N_noxref_6_c_438_n ) capacitor c=0.0259045f //x=0.81 \
 //y=1.915 //x2=1.475 //y2=1.59
cc_259 ( N_A_c_320_n N_noxref_6_c_438_n ) capacitor c=0.00708583f //x=1.185 \
 //y=1.375 //x2=1.475 //y2=1.59
cc_260 ( N_A_c_323_n N_noxref_6_c_438_n ) capacitor c=0.00698822f //x=1.34 \
 //y=1.22 //x2=1.475 //y2=1.59
cc_261 ( N_A_c_314_n N_noxref_6_M0_noxref_s ) capacitor c=0.0327271f //x=0.81 \
 //y=0.875 //x2=0.455 //y2=0.375
cc_262 ( N_A_c_317_n N_noxref_6_M0_noxref_s ) capacitor c=7.99997e-19 //x=0.81 \
 //y=1.53 //x2=0.455 //y2=0.375
cc_263 ( N_A_c_318_n N_noxref_6_M0_noxref_s ) capacitor c=0.00122123f //x=0.81 \
 //y=1.915 //x2=0.455 //y2=0.375
cc_264 ( N_A_c_321_n N_noxref_6_M0_noxref_s ) capacitor c=0.0121427f //x=1.34 \
 //y=0.875 //x2=0.455 //y2=0.375
cc_265 ( N_A_c_313_n N_C_c_483_n ) capacitor c=0.00155228f //x=1.11 //y=2.08 \
 //x2=3.33 //y2=2.08
cc_266 ( N_B_c_390_n N_noxref_6_c_446_n ) capacitor c=0.0167228f //x=1.785 \
 //y=0.91 //x2=2.445 //y2=0.54
cc_267 ( N_B_c_395_n N_noxref_6_c_446_n ) capacitor c=0.00534519f //x=2.31 \
 //y=0.91 //x2=2.445 //y2=0.54
cc_268 ( N_B_c_368_n N_noxref_6_c_469_n ) capacitor c=0.0124072f //x=2.22 \
 //y=2.08 //x2=2.445 //y2=1.59
cc_269 ( N_B_c_393_n N_noxref_6_c_469_n ) capacitor c=0.0153476f //x=1.785 \
 //y=1.22 //x2=2.445 //y2=1.59
cc_270 ( N_B_c_398_n N_noxref_6_c_469_n ) capacitor c=0.023396f //x=2.31 \
 //y=1.915 //x2=2.445 //y2=1.59
cc_271 ( N_B_c_390_n N_noxref_6_M0_noxref_s ) capacitor c=0.00798959f \
 //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_272 ( N_B_c_397_n N_noxref_6_M0_noxref_s ) capacitor c=0.00212176f //x=2.31 \
 //y=1.45 //x2=0.455 //y2=0.375
cc_273 ( N_B_c_398_n N_noxref_6_M0_noxref_s ) capacitor c=0.00298115f //x=2.31 \
 //y=1.915 //x2=0.455 //y2=0.375
cc_274 ( N_B_c_368_n N_C_c_483_n ) capacitor c=0.05827f //x=2.22 //y=2.08 \
 //x2=3.33 //y2=2.08
cc_275 ( N_B_c_398_n N_C_c_483_n ) capacitor c=0.0023343f //x=2.31 //y=1.915 \
 //x2=3.33 //y2=2.08
cc_276 ( N_B_c_382_n N_C_c_483_n ) capacitor c=0.00142741f //x=2.22 //y=4.7 \
 //x2=3.33 //y2=2.08
cc_277 ( N_B_M6_noxref_g N_C_M8_noxref_g ) capacitor c=0.0101598f //x=2.19 \
 //y=6.02 //x2=3.07 //y2=6.02
cc_278 ( N_B_M7_noxref_g N_C_M8_noxref_g ) capacitor c=0.0602553f //x=2.63 \
 //y=6.02 //x2=3.07 //y2=6.02
cc_279 ( N_B_M7_noxref_g N_C_M9_noxref_g ) capacitor c=0.0101598f //x=2.63 \
 //y=6.02 //x2=3.51 //y2=6.02
cc_280 ( N_B_c_395_n N_C_c_497_n ) capacitor c=0.00456962f //x=2.31 //y=0.91 \
 //x2=3.32 //y2=0.915
cc_281 ( N_B_c_396_n N_C_c_498_n ) capacitor c=0.00438372f //x=2.31 //y=1.22 \
 //x2=3.32 //y2=1.26
cc_282 ( N_B_c_397_n N_C_c_499_n ) capacitor c=0.00438372f //x=2.31 //y=1.45 \
 //x2=3.32 //y2=1.57
cc_283 ( N_B_c_368_n N_C_c_506_n ) capacitor c=0.00228632f //x=2.22 //y=2.08 \
 //x2=3.33 //y2=2.08
cc_284 ( N_B_c_398_n N_C_c_506_n ) capacitor c=0.00933826f //x=2.31 //y=1.915 \
 //x2=3.33 //y2=2.08
cc_285 ( N_B_c_398_n N_C_c_507_n ) capacitor c=0.00438372f //x=2.31 //y=1.915 \
 //x2=3.33 //y2=1.915
cc_286 ( N_B_c_368_n N_C_c_509_n ) capacitor c=0.00219458f //x=2.22 //y=2.08 \
 //x2=3.33 //y2=4.7
cc_287 ( N_B_c_381_n N_C_c_509_n ) capacitor c=0.0611812f //x=2.555 //y=4.79 \
 //x2=3.33 //y2=4.7
cc_288 ( N_B_c_382_n N_C_c_509_n ) capacitor c=0.00487508f //x=2.22 //y=4.7 \
 //x2=3.33 //y2=4.7
cc_289 ( N_B_c_426_p N_noxref_8_c_537_n ) capacitor c=2.14837e-19 //x=2.155 \
 //y=0.755 //x2=3.015 //y2=0.995
cc_290 ( N_B_c_395_n N_noxref_8_c_537_n ) capacitor c=0.00123426f //x=2.31 \
 //y=0.91 //x2=3.015 //y2=0.995
cc_291 ( N_B_c_396_n N_noxref_8_c_537_n ) capacitor c=0.0129288f //x=2.31 \
 //y=1.22 //x2=3.015 //y2=0.995
cc_292 ( N_B_c_397_n N_noxref_8_c_537_n ) capacitor c=0.00142359f //x=2.31 \
 //y=1.45 //x2=3.015 //y2=0.995
cc_293 ( N_B_c_390_n N_noxref_8_M1_noxref_d ) capacitor c=0.00223875f \
 //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_294 ( N_B_c_393_n N_noxref_8_M1_noxref_d ) capacitor c=0.00262485f \
 //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_295 ( N_B_c_426_p N_noxref_8_M1_noxref_d ) capacitor c=0.00220746f \
 //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_296 ( N_B_c_433_p N_noxref_8_M1_noxref_d ) capacitor c=0.00194798f \
 //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_297 ( N_B_c_395_n N_noxref_8_M1_noxref_d ) capacitor c=0.00198465f //x=2.31 \
 //y=0.91 //x2=1.86 //y2=0.91
cc_298 ( N_B_c_396_n N_noxref_8_M1_noxref_d ) capacitor c=0.00128384f //x=2.31 \
 //y=1.22 //x2=1.86 //y2=0.91
cc_299 ( N_B_c_395_n N_noxref_8_M2_noxref_s ) capacitor c=7.21316e-19 //x=2.31 \
 //y=0.91 //x2=2.965 //y2=0.375
cc_300 ( N_B_c_396_n N_noxref_8_M2_noxref_s ) capacitor c=0.00348171f //x=2.31 \
 //y=1.22 //x2=2.965 //y2=0.375
cc_301 ( N_noxref_6_c_446_n N_noxref_8_c_537_n ) capacitor c=0.0136048f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_302 ( N_noxref_6_c_469_n N_noxref_8_c_537_n ) capacitor c=0.0102337f \
 //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_303 ( N_noxref_6_M0_noxref_s N_noxref_8_c_537_n ) capacitor c=0.023368f \
 //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_304 ( N_noxref_6_M0_noxref_s N_noxref_8_c_540_n ) capacitor c=0.0180035f \
 //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_305 ( N_noxref_6_c_446_n N_noxref_8_M1_noxref_d ) capacitor c=0.0129526f \
 //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_306 ( N_noxref_6_c_469_n N_noxref_8_M1_noxref_d ) capacitor c=0.0091401f \
 //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_307 ( N_noxref_6_M0_noxref_s N_noxref_8_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_308 ( N_noxref_6_M0_noxref_s N_noxref_8_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_309 ( N_C_c_483_n N_noxref_8_c_544_n ) capacitor c=0.00210069f //x=3.33 \
 //y=2.08 //x2=3.985 //y2=0.54
cc_310 ( N_C_c_497_n N_noxref_8_c_544_n ) capacitor c=0.0192822f //x=3.32 \
 //y=0.915 //x2=3.985 //y2=0.54
cc_311 ( N_C_c_503_n N_noxref_8_c_544_n ) capacitor c=0.00656458f //x=3.85 \
 //y=0.915 //x2=3.985 //y2=0.54
cc_312 ( N_C_c_506_n N_noxref_8_c_544_n ) capacitor c=2.20712e-19 //x=3.33 \
 //y=2.08 //x2=3.985 //y2=0.54
cc_313 ( N_C_c_498_n N_noxref_8_c_558_n ) capacitor c=0.00538829f //x=3.32 \
 //y=1.26 //x2=3.1 //y2=0.995
cc_314 ( N_C_c_497_n N_noxref_8_M2_noxref_s ) capacitor c=0.00538829f //x=3.32 \
 //y=0.915 //x2=2.965 //y2=0.375
cc_315 ( N_C_c_499_n N_noxref_8_M2_noxref_s ) capacitor c=0.00538829f //x=3.32 \
 //y=1.57 //x2=2.965 //y2=0.375
cc_316 ( N_C_c_503_n N_noxref_8_M2_noxref_s ) capacitor c=0.0143002f //x=3.85 \
 //y=0.915 //x2=2.965 //y2=0.375
cc_317 ( N_C_c_504_n N_noxref_8_M2_noxref_s ) capacitor c=0.00290153f //x=3.85 \
 //y=1.26 //x2=2.965 //y2=0.375
