* SPICE3 file created from HA.ext - technology: sky130A

.subckt HA SUM COUT A B VPB VNB
M1000 SUM B a_1666_74.t0 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.14u as=0p ps=0u
M1001 VNB A a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=3.9597p pd=29.01u as=0p ps=0u
M1002 SUM a_1295_182.t3 a_2351_1004.t3 pshort w=2u l=0.15u
+  ad=1.16p pd=9.16u as=0p ps=0u
M1003 a_1917_943.t1 B VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VNB a_1917_943.t3 a_2332_74.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t9 A a_217_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_851_182.t2 a_217_1004.t5 VPB.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_1685_1004.t1 a_1917_943.t4 SUM pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t5 B a_217_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 SUM a_1917_943.t5 a_1685_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t10 A a_1685_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 SUM a_1295_182.t4 a_2332_74.t1 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t12 a_217_1004.t6 a_851_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPB.t7 A a_1295_182.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_2351_1004.t1 B VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_217_1004.t3 A VPB.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VNB A a_1666_74.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_2351_1004.t2 a_1295_182.t5 SUM pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_217_1004.t1 B VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1685_1004.t2 A VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPB.t2 B a_2351_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPB.t0 B a_1917_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1295_182.t1 A VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 A B 2.16fF
C1 A SUM 0.07fF
C2 SUM B 1.08fF
C3 A VPB 0.67fF
C4 B VPB 0.65fF
C5 SUM VPB 0.53fF
R0 a_1917_943.n2 a_1917_943.t5 477.179
R1 a_1917_943.n4 a_1917_943.t3 420.747
R2 a_1917_943.n2 a_1917_943.t4 406.485
R3 a_1917_943.n3 a_1917_943.n2 211.151
R4 a_1917_943.n6 a_1917_943.n4 188.704
R5 a_1917_943.n3 a_1917_943.n1 114.038
R6 a_1917_943.n4 a_1917_943.n3 53.105
R7 a_1917_943.n6 a_1917_943.n5 30
R8 a_1917_943.n7 a_1917_943.n0 24.383
R9 a_1917_943.n7 a_1917_943.n6 23.684
R10 a_1917_943.n1 a_1917_943.t0 14.282
R11 a_1917_943.n1 a_1917_943.t1 14.282
R12 a_2332_74.n10 a_2332_74.n9 93.333
R13 a_2332_74.n2 a_2332_74.n1 41.622
R14 a_2332_74.n13 a_2332_74.n12 26.667
R15 a_2332_74.n6 a_2332_74.n5 24.977
R16 a_2332_74.t0 a_2332_74.n2 21.209
R17 a_2332_74.t0 a_2332_74.n3 11.595
R18 a_2332_74.t1 a_2332_74.n8 8.137
R19 a_2332_74.t0 a_2332_74.n0 6.109
R20 a_2332_74.t1 a_2332_74.n7 4.864
R21 a_2332_74.t0 a_2332_74.n4 3.871
R22 a_2332_74.t0 a_2332_74.n13 2.535
R23 a_2332_74.n13 a_2332_74.t1 1.145
R24 a_2332_74.n7 a_2332_74.n6 1.13
R25 a_2332_74.t1 a_2332_74.n11 0.804
R26 a_2332_74.n11 a_2332_74.n10 0.136
R27 VNB VNB.n339 300.778
R28 VNB.n185 VNB.n184 199.897
R29 VNB.n85 VNB.n84 199.897
R30 VNB.n237 VNB.n236 199.897
R31 VNB.n295 VNB.n294 199.897
R32 VNB.n18 VNB.n17 199.897
R33 VNB.n266 VNB.n265 158.304
R34 VNB.n108 VNB.n106 154.509
R35 VNB.n194 VNB.n192 154.509
R36 VNB.n304 VNB.n302 154.509
R37 VNB.n246 VNB.n244 154.509
R38 VNB.n46 VNB.n44 154.509
R39 VNB.n120 VNB.n119 121.366
R40 VNB.n58 VNB.n57 121.366
R41 VNB.n255 VNB.n254 105.536
R42 VNB.n95 VNB.n91 85.201
R43 VNB.n155 VNB.n147 76.136
R44 VNB.n155 VNB.n154 76
R45 VNB.n326 VNB.n325 76
R46 VNB.n314 VNB.n313 76
R47 VNB.n306 VNB.n305 76
R48 VNB.n284 VNB.n283 76
R49 VNB.n280 VNB.n279 76
R50 VNB.n270 VNB.n269 76
R51 VNB.n258 VNB.n257 76
R52 VNB.n248 VNB.n247 76
R53 VNB.n226 VNB.n225 76
R54 VNB.n222 VNB.n219 76
R55 VNB.n208 VNB.n207 76
R56 VNB.n204 VNB.n203 76
R57 VNB.n200 VNB.n199 76
R58 VNB.n196 VNB.n195 76
R59 VNB.n174 VNB.n173 76
R60 VNB.n170 VNB.n169 76
R61 VNB.n162 VNB.n161 76
R62 VNB.n124 VNB.n74 64.194
R63 VNB.n62 VNB.n7 63.835
R64 VNB.n34 VNB.n33 49.896
R65 VNB.n274 VNB.t2 39.412
R66 VNB.n121 VNB.n120 36.937
R67 VNB.n59 VNB.n58 36.937
R68 VNB.n97 VNB.n96 36.678
R69 VNB.n252 VNB.n251 35.01
R70 VNB.n309 VNB.n308 35.01
R71 VNB.t5 VNB.n26 32.601
R72 VNB.n74 VNB.n73 28.421
R73 VNB.n7 VNB.n6 28.421
R74 VNB.n127 VNB.n126 27.855
R75 VNB.n267 VNB.n264 27.855
R76 VNB.n65 VNB.n64 27.855
R77 VNB.n74 VNB.n72 25.263
R78 VNB.n7 VNB.n5 25.263
R79 VNB.n72 VNB.n71 24.383
R80 VNB.n5 VNB.n4 24.383
R81 VNB.n147 VNB.n144 20.452
R82 VNB.n327 VNB.n326 20.452
R83 VNB.n151 VNB.n150 20.094
R84 VNB.n158 VNB.n157 20.094
R85 VNB.n166 VNB.n165 20.094
R86 VNB.n253 VNB.n252 20.094
R87 VNB.n263 VNB.n262 20.094
R88 VNB.n276 VNB.n275 20.094
R89 VNB.n310 VNB.n309 20.094
R90 VNB.n32 VNB.n31 20.094
R91 VNB.n39 VNB.n29 20.094
R92 VNB.n252 VNB.n250 19.017
R93 VNB.n309 VNB.n307 19.017
R94 VNB.n156 VNB.t0 18.552
R95 VNB.n160 VNB.n159 18.269
R96 VNB.n28 VNB.t5 17.353
R97 VNB.n274 VNB.n273 17.185
R98 VNB.n128 VNB.n127 16.721
R99 VNB.n268 VNB.n267 16.721
R100 VNB.n66 VNB.n65 16.721
R101 VNB.n154 VNB.n153 13.653
R102 VNB.n153 VNB.n152 13.653
R103 VNB.n161 VNB.n160 13.653
R104 VNB.n169 VNB.n168 13.653
R105 VNB.n168 VNB.n167 13.653
R106 VNB.n173 VNB.n172 13.653
R107 VNB.n172 VNB.n171 13.653
R108 VNB.n195 VNB.n194 13.653
R109 VNB.n194 VNB.n193 13.653
R110 VNB.n199 VNB.n198 13.653
R111 VNB.n198 VNB.n197 13.653
R112 VNB.n203 VNB.n202 13.653
R113 VNB.n202 VNB.n201 13.653
R114 VNB.n207 VNB.n206 13.653
R115 VNB.n206 VNB.n205 13.653
R116 VNB.n94 VNB.n93 13.653
R117 VNB.n93 VNB.n92 13.653
R118 VNB.n98 VNB.n97 13.653
R119 VNB.n101 VNB.n100 13.653
R120 VNB.n100 VNB.n99 13.653
R121 VNB.n104 VNB.n103 13.653
R122 VNB.n103 VNB.n102 13.653
R123 VNB.n109 VNB.n108 13.653
R124 VNB.n108 VNB.n107 13.653
R125 VNB.n112 VNB.n111 13.653
R126 VNB.n111 VNB.n110 13.653
R127 VNB.n115 VNB.n114 13.653
R128 VNB.n114 VNB.n113 13.653
R129 VNB.n118 VNB.n117 13.653
R130 VNB.n117 VNB.n116 13.653
R131 VNB.n123 VNB.n122 13.653
R132 VNB.n122 VNB.n121 13.653
R133 VNB.n129 VNB.n128 13.653
R134 VNB.n222 VNB.n221 13.653
R135 VNB.n221 VNB.n220 13.653
R136 VNB.n225 VNB.n224 13.653
R137 VNB.n224 VNB.n223 13.653
R138 VNB.n247 VNB.n246 13.653
R139 VNB.n246 VNB.n245 13.653
R140 VNB.n257 VNB.n256 13.653
R141 VNB.n256 VNB.n255 13.653
R142 VNB.n269 VNB.n268 13.653
R143 VNB.n279 VNB.n278 13.653
R144 VNB.n278 VNB.n277 13.653
R145 VNB.n283 VNB.n282 13.653
R146 VNB.n282 VNB.n281 13.653
R147 VNB.n305 VNB.n304 13.653
R148 VNB.n304 VNB.n303 13.653
R149 VNB.n313 VNB.n312 13.653
R150 VNB.n312 VNB.n311 13.653
R151 VNB.n35 VNB.n34 13.653
R152 VNB.n38 VNB.n37 13.653
R153 VNB.n37 VNB.n36 13.653
R154 VNB.n42 VNB.n41 13.653
R155 VNB.n41 VNB.n40 13.653
R156 VNB.n47 VNB.n46 13.653
R157 VNB.n46 VNB.n45 13.653
R158 VNB.n50 VNB.n49 13.653
R159 VNB.n49 VNB.n48 13.653
R160 VNB.n53 VNB.n52 13.653
R161 VNB.n52 VNB.n51 13.653
R162 VNB.n56 VNB.n55 13.653
R163 VNB.n55 VNB.n54 13.653
R164 VNB.n61 VNB.n60 13.653
R165 VNB.n60 VNB.n59 13.653
R166 VNB.n67 VNB.n66 13.653
R167 VNB.n70 VNB.n69 13.653
R168 VNB.n69 VNB.n68 13.653
R169 VNB.n326 VNB.n0 13.653
R170 VNB VNB.n0 13.653
R171 VNB.n147 VNB.n146 13.653
R172 VNB.n146 VNB.n145 13.653
R173 VNB.n165 VNB.n164 13.608
R174 VNB.n334 VNB.n331 13.577
R175 VNB.n132 VNB.n130 13.276
R176 VNB.n144 VNB.n132 13.276
R177 VNB.n177 VNB.n175 13.276
R178 VNB.n190 VNB.n177 13.276
R179 VNB.n77 VNB.n75 13.276
R180 VNB.n90 VNB.n77 13.276
R181 VNB.n229 VNB.n227 13.276
R182 VNB.n242 VNB.n229 13.276
R183 VNB.n287 VNB.n285 13.276
R184 VNB.n300 VNB.n287 13.276
R185 VNB.n10 VNB.n8 13.276
R186 VNB.n23 VNB.n10 13.276
R187 VNB.n195 VNB.n191 13.276
R188 VNB.n101 VNB.n98 13.276
R189 VNB.n104 VNB.n101 13.276
R190 VNB.n105 VNB.n104 13.276
R191 VNB.n109 VNB.n105 13.276
R192 VNB.n112 VNB.n109 13.276
R193 VNB.n115 VNB.n112 13.276
R194 VNB.n118 VNB.n115 13.276
R195 VNB.n123 VNB.n118 13.276
R196 VNB.n222 VNB.n129 13.276
R197 VNB.n225 VNB.n222 13.276
R198 VNB.n247 VNB.n243 13.276
R199 VNB.n305 VNB.n301 13.276
R200 VNB.n38 VNB.n35 13.276
R201 VNB.n43 VNB.n42 13.276
R202 VNB.n47 VNB.n43 13.276
R203 VNB.n50 VNB.n47 13.276
R204 VNB.n53 VNB.n50 13.276
R205 VNB.n56 VNB.n53 13.276
R206 VNB.n61 VNB.n56 13.276
R207 VNB.n70 VNB.n67 13.276
R208 VNB.n326 VNB.n70 13.276
R209 VNB.n3 VNB.n1 13.276
R210 VNB.n327 VNB.n3 13.276
R211 VNB.n29 VNB.n28 12.837
R212 VNB.n150 VNB.n149 10.853
R213 VNB.n95 VNB.n94 10.764
R214 VNB.n124 VNB.n123 10.764
R215 VNB.n62 VNB.n61 10.764
R216 VNB.n149 VNB.n148 10.417
R217 VNB.n42 VNB.n39 9.329
R218 VNB.n164 VNB.n163 7.858
R219 VNB.n28 VNB.n27 7.566
R220 VNB.n250 VNB.n249 7.5
R221 VNB.n261 VNB.n260 7.5
R222 VNB.n336 VNB.n335 7.5
R223 VNB.n183 VNB.n182 7.5
R224 VNB.n179 VNB.n178 7.5
R225 VNB.n177 VNB.n176 7.5
R226 VNB.n190 VNB.n189 7.5
R227 VNB.n83 VNB.n82 7.5
R228 VNB.n79 VNB.n78 7.5
R229 VNB.n77 VNB.n76 7.5
R230 VNB.n90 VNB.n89 7.5
R231 VNB.n235 VNB.n234 7.5
R232 VNB.n231 VNB.n230 7.5
R233 VNB.n229 VNB.n228 7.5
R234 VNB.n242 VNB.n241 7.5
R235 VNB.n293 VNB.n292 7.5
R236 VNB.n289 VNB.n288 7.5
R237 VNB.n287 VNB.n286 7.5
R238 VNB.n300 VNB.n299 7.5
R239 VNB.n16 VNB.n15 7.5
R240 VNB.n12 VNB.n11 7.5
R241 VNB.n10 VNB.n9 7.5
R242 VNB.n23 VNB.n22 7.5
R243 VNB.n328 VNB.n327 7.5
R244 VNB.n3 VNB.n2 7.5
R245 VNB.n333 VNB.n332 7.5
R246 VNB.n138 VNB.n137 7.5
R247 VNB.n134 VNB.n133 7.5
R248 VNB.n132 VNB.n131 7.5
R249 VNB.n144 VNB.n143 7.5
R250 VNB.n191 VNB.n190 7.176
R251 VNB.n105 VNB.n90 7.176
R252 VNB.n243 VNB.n242 7.176
R253 VNB.n301 VNB.n300 7.176
R254 VNB.n43 VNB.n23 7.176
R255 VNB.n338 VNB.n336 7.011
R256 VNB.n186 VNB.n183 7.011
R257 VNB.n181 VNB.n179 7.011
R258 VNB.n86 VNB.n83 7.011
R259 VNB.n81 VNB.n79 7.011
R260 VNB.n238 VNB.n235 7.011
R261 VNB.n233 VNB.n231 7.011
R262 VNB.n296 VNB.n293 7.011
R263 VNB.n291 VNB.n289 7.011
R264 VNB.n19 VNB.n16 7.011
R265 VNB.n14 VNB.n12 7.011
R266 VNB.n140 VNB.n138 7.011
R267 VNB.n136 VNB.n134 7.011
R268 VNB.n189 VNB.n188 7.01
R269 VNB.n181 VNB.n180 7.01
R270 VNB.n186 VNB.n185 7.01
R271 VNB.n89 VNB.n88 7.01
R272 VNB.n81 VNB.n80 7.01
R273 VNB.n86 VNB.n85 7.01
R274 VNB.n241 VNB.n240 7.01
R275 VNB.n233 VNB.n232 7.01
R276 VNB.n238 VNB.n237 7.01
R277 VNB.n299 VNB.n298 7.01
R278 VNB.n291 VNB.n290 7.01
R279 VNB.n296 VNB.n295 7.01
R280 VNB.n22 VNB.n21 7.01
R281 VNB.n14 VNB.n13 7.01
R282 VNB.n19 VNB.n18 7.01
R283 VNB.n143 VNB.n142 7.01
R284 VNB.n136 VNB.n135 7.01
R285 VNB.n140 VNB.n139 7.01
R286 VNB.n338 VNB.n337 7.01
R287 VNB.n334 VNB.n333 6.788
R288 VNB.n329 VNB.n328 6.788
R289 VNB.n275 VNB.n274 6.139
R290 VNB.n272 VNB.n271 4.551
R291 VNB.n25 VNB.n24 4.551
R292 VNB.n169 VNB.n166 4.305
R293 VNB.n257 VNB.n253 4.305
R294 VNB.n313 VNB.n310 4.305
R295 VNB.n154 VNB.n151 3.947
R296 VNB.n279 VNB.n276 3.947
R297 VNB.n39 VNB.n38 3.947
R298 VNB.n98 VNB.n95 2.511
R299 VNB.n129 VNB.n124 2.511
R300 VNB.n67 VNB.n62 2.511
R301 VNB.t2 VNB.n272 2.238
R302 VNB.t5 VNB.n25 2.238
R303 VNB.n127 VNB.n125 1.99
R304 VNB.n267 VNB.n266 1.99
R305 VNB.n65 VNB.n63 1.99
R306 VNB.n260 VNB.n259 1.935
R307 VNB.n339 VNB.n330 0.921
R308 VNB.n339 VNB.n334 0.476
R309 VNB.n339 VNB.n329 0.475
R310 VNB.n157 VNB.n156 0.358
R311 VNB.n262 VNB.n261 0.358
R312 VNB.n31 VNB.n30 0.358
R313 VNB.n196 VNB.n174 0.272
R314 VNB.n213 VNB.n212 0.272
R315 VNB.n248 VNB.n226 0.272
R316 VNB.n306 VNB.n284 0.272
R317 VNB.n318 VNB.n317 0.272
R318 VNB.n187 VNB.n181 0.246
R319 VNB.n188 VNB.n187 0.246
R320 VNB.n187 VNB.n186 0.246
R321 VNB.n87 VNB.n81 0.246
R322 VNB.n88 VNB.n87 0.246
R323 VNB.n87 VNB.n86 0.246
R324 VNB.n239 VNB.n233 0.246
R325 VNB.n240 VNB.n239 0.246
R326 VNB.n239 VNB.n238 0.246
R327 VNB.n297 VNB.n291 0.246
R328 VNB.n298 VNB.n297 0.246
R329 VNB.n297 VNB.n296 0.246
R330 VNB.n20 VNB.n14 0.246
R331 VNB.n21 VNB.n20 0.246
R332 VNB.n20 VNB.n19 0.246
R333 VNB.n141 VNB.n136 0.246
R334 VNB.n142 VNB.n141 0.246
R335 VNB.n141 VNB.n140 0.246
R336 VNB.n339 VNB.n338 0.246
R337 VNB.n325 VNB 0.198
R338 VNB.n161 VNB.n158 0.179
R339 VNB.n269 VNB.n263 0.179
R340 VNB.n35 VNB.n32 0.179
R341 VNB.n162 VNB.n155 0.136
R342 VNB.n170 VNB.n162 0.136
R343 VNB.n174 VNB.n170 0.136
R344 VNB.n200 VNB.n196 0.136
R345 VNB.n204 VNB.n200 0.136
R346 VNB.n208 VNB.n204 0.136
R347 VNB.n209 VNB.n208 0.136
R348 VNB.n210 VNB.n209 0.136
R349 VNB.n211 VNB.n210 0.136
R350 VNB.n212 VNB.n211 0.136
R351 VNB.n214 VNB.n213 0.136
R352 VNB.n215 VNB.n214 0.136
R353 VNB.n216 VNB.n215 0.136
R354 VNB.n217 VNB.n216 0.136
R355 VNB.n218 VNB.n217 0.136
R356 VNB.n219 VNB.n218 0.136
R357 VNB.n258 VNB.n248 0.136
R358 VNB.n270 VNB.n258 0.136
R359 VNB.n280 VNB.n270 0.136
R360 VNB.n284 VNB.n280 0.136
R361 VNB.n314 VNB.n306 0.136
R362 VNB.n315 VNB.n314 0.136
R363 VNB.n316 VNB.n315 0.136
R364 VNB.n317 VNB.n316 0.136
R365 VNB.n319 VNB.n318 0.136
R366 VNB.n320 VNB.n319 0.136
R367 VNB.n321 VNB.n320 0.136
R368 VNB.n322 VNB.n321 0.136
R369 VNB.n323 VNB.n322 0.136
R370 VNB.n324 VNB.n323 0.136
R371 VNB.n325 VNB.n324 0.136
R372 VNB.n219 VNB 0.068
R373 VNB.n226 VNB 0.068
R374 a_1295_182.n1 a_1295_182.t3 477.179
R375 a_1295_182.n1 a_1295_182.t5 406.485
R376 a_1295_182.n2 a_1295_182.t4 225.731
R377 a_1295_182.n3 a_1295_182.n0 220.249
R378 a_1295_182.n2 a_1295_182.n1 161.6
R379 a_1295_182.n3 a_1295_182.n2 156.579
R380 a_1295_182.n5 a_1295_182.n3 142.121
R381 a_1295_182.n5 a_1295_182.n4 15.218
R382 a_1295_182.n0 a_1295_182.t0 14.282
R383 a_1295_182.n0 a_1295_182.t1 14.282
R384 a_1295_182.n6 a_1295_182.n5 12.014
R385 a_2351_1004.t2 a_2351_1004.n0 101.663
R386 a_2351_1004.n0 a_2351_1004.t0 101.661
R387 a_2351_1004.n0 a_2351_1004.t3 14.294
R388 a_2351_1004.n0 a_2351_1004.t1 14.282
R389 VPB VPB.n337 126.832
R390 VPB.n50 VPB.n48 94.117
R391 VPB.n310 VPB.n308 94.117
R392 VPB.n263 VPB.n261 94.117
R393 VPB.n118 VPB.n116 94.117
R394 VPB.n206 VPB.n204 94.117
R395 VPB.n167 VPB.n161 76.136
R396 VPB.n167 VPB.n166 76
R397 VPB.n171 VPB.n170 76
R398 VPB.n177 VPB.n176 76
R399 VPB.n181 VPB.n180 76
R400 VPB.n208 VPB.n207 76
R401 VPB.n212 VPB.n211 76
R402 VPB.n216 VPB.n215 76
R403 VPB.n220 VPB.n219 76
R404 VPB.n234 VPB.n231 76
R405 VPB.n238 VPB.n237 76
R406 VPB.n265 VPB.n264 76
R407 VPB.n271 VPB.n270 76
R408 VPB.n275 VPB.n274 76
R409 VPB.n281 VPB.n280 76
R410 VPB.n285 VPB.n284 76
R411 VPB.n312 VPB.n311 76
R412 VPB.n318 VPB.n317 76
R413 VPB.n330 VPB.n329 76
R414 VPB.n164 VPB.n163 68.979
R415 VPB.n278 VPB.n277 68.979
R416 VPB.n40 VPB.n39 68.979
R417 VPB.n133 VPB.n77 65.944
R418 VPB.n104 VPB.n99 65.944
R419 VPB.n174 VPB.n173 64.528
R420 VPB.n268 VPB.n267 64.528
R421 VPB.n315 VPB.n314 64.528
R422 VPB.n21 VPB.n20 61.764
R423 VPB.n292 VPB.n291 61.764
R424 VPB.n245 VPB.n244 61.764
R425 VPB.n84 VPB.n83 61.764
R426 VPB.n188 VPB.n187 61.764
R427 VPB.n73 VPB.t8 55.106
R428 VPB.n43 VPB.t13 55.106
R429 VPB.n313 VPB.t12 55.106
R430 VPB.n276 VPB.t6 55.106
R431 VPB.n266 VPB.t7 55.106
R432 VPB.n172 VPB.t1 55.106
R433 VPB.n162 VPB.t0 55.106
R434 VPB.n55 VPB.t5 55.106
R435 VPB.n57 VPB.n56 48.952
R436 VPB.n106 VPB.n105 44.502
R437 VPB.n135 VPB.n134 44.502
R438 VPB.n70 VPB.n69 44.502
R439 VPB.n64 VPB.n14 40.824
R440 VPB.n334 VPB.n330 20.452
R441 VPB.n161 VPB.n158 20.452
R442 VPB.n61 VPB.n60 17.801
R443 VPB.n14 VPB.t4 14.282
R444 VPB.n14 VPB.t9 14.282
R445 VPB.n77 VPB.t11 14.282
R446 VPB.n77 VPB.t10 14.282
R447 VPB.n99 VPB.t3 14.282
R448 VPB.n99 VPB.t2 14.282
R449 VPB.n161 VPB.n160 13.653
R450 VPB.n160 VPB.n159 13.653
R451 VPB.n166 VPB.n165 13.653
R452 VPB.n165 VPB.n164 13.653
R453 VPB.n170 VPB.n169 13.653
R454 VPB.n169 VPB.n168 13.653
R455 VPB.n176 VPB.n175 13.653
R456 VPB.n175 VPB.n174 13.653
R457 VPB.n180 VPB.n179 13.653
R458 VPB.n179 VPB.n178 13.653
R459 VPB.n207 VPB.n206 13.653
R460 VPB.n206 VPB.n205 13.653
R461 VPB.n211 VPB.n210 13.653
R462 VPB.n210 VPB.n209 13.653
R463 VPB.n215 VPB.n214 13.653
R464 VPB.n214 VPB.n213 13.653
R465 VPB.n219 VPB.n218 13.653
R466 VPB.n218 VPB.n217 13.653
R467 VPB.n103 VPB.n102 13.653
R468 VPB.n102 VPB.n101 13.653
R469 VPB.n108 VPB.n107 13.653
R470 VPB.n107 VPB.n106 13.653
R471 VPB.n111 VPB.n110 13.653
R472 VPB.n110 VPB.n109 13.653
R473 VPB.n114 VPB.n113 13.653
R474 VPB.n113 VPB.n112 13.653
R475 VPB.n119 VPB.n118 13.653
R476 VPB.n118 VPB.n117 13.653
R477 VPB.n122 VPB.n121 13.653
R478 VPB.n121 VPB.n120 13.653
R479 VPB.n125 VPB.n124 13.653
R480 VPB.n124 VPB.n123 13.653
R481 VPB.n128 VPB.n127 13.653
R482 VPB.n127 VPB.n126 13.653
R483 VPB.n132 VPB.n131 13.653
R484 VPB.n131 VPB.n130 13.653
R485 VPB.n137 VPB.n136 13.653
R486 VPB.n136 VPB.n135 13.653
R487 VPB.n234 VPB.n233 13.653
R488 VPB.n233 VPB.n232 13.653
R489 VPB.n237 VPB.n236 13.653
R490 VPB.n236 VPB.n235 13.653
R491 VPB.n264 VPB.n263 13.653
R492 VPB.n263 VPB.n262 13.653
R493 VPB.n270 VPB.n269 13.653
R494 VPB.n269 VPB.n268 13.653
R495 VPB.n274 VPB.n273 13.653
R496 VPB.n273 VPB.n272 13.653
R497 VPB.n280 VPB.n279 13.653
R498 VPB.n279 VPB.n278 13.653
R499 VPB.n284 VPB.n283 13.653
R500 VPB.n283 VPB.n282 13.653
R501 VPB.n311 VPB.n310 13.653
R502 VPB.n310 VPB.n309 13.653
R503 VPB.n317 VPB.n316 13.653
R504 VPB.n316 VPB.n315 13.653
R505 VPB.n38 VPB.n37 13.653
R506 VPB.n37 VPB.n36 13.653
R507 VPB.n42 VPB.n41 13.653
R508 VPB.n41 VPB.n40 13.653
R509 VPB.n46 VPB.n45 13.653
R510 VPB.n45 VPB.n44 13.653
R511 VPB.n51 VPB.n50 13.653
R512 VPB.n50 VPB.n49 13.653
R513 VPB.n54 VPB.n53 13.653
R514 VPB.n53 VPB.n52 13.653
R515 VPB.n59 VPB.n58 13.653
R516 VPB.n58 VPB.n57 13.653
R517 VPB.n63 VPB.n62 13.653
R518 VPB.n62 VPB.n61 13.653
R519 VPB.n68 VPB.n67 13.653
R520 VPB.n67 VPB.n66 13.653
R521 VPB.n72 VPB.n71 13.653
R522 VPB.n71 VPB.n70 13.653
R523 VPB.n76 VPB.n75 13.653
R524 VPB.n75 VPB.n74 13.653
R525 VPB.n330 VPB.n0 13.653
R526 VPB VPB.n0 13.653
R527 VPB.n101 VPB.n100 13.35
R528 VPB.n130 VPB.n129 13.35
R529 VPB.n66 VPB.n65 13.35
R530 VPB.n334 VPB.n333 13.276
R531 VPB.n333 VPB.n331 13.276
R532 VPB.n35 VPB.n17 13.276
R533 VPB.n17 VPB.n15 13.276
R534 VPB.n306 VPB.n288 13.276
R535 VPB.n288 VPB.n286 13.276
R536 VPB.n259 VPB.n241 13.276
R537 VPB.n241 VPB.n239 13.276
R538 VPB.n98 VPB.n80 13.276
R539 VPB.n80 VPB.n78 13.276
R540 VPB.n202 VPB.n184 13.276
R541 VPB.n184 VPB.n182 13.276
R542 VPB.n207 VPB.n203 13.276
R543 VPB.n111 VPB.n108 13.276
R544 VPB.n114 VPB.n111 13.276
R545 VPB.n115 VPB.n114 13.276
R546 VPB.n119 VPB.n115 13.276
R547 VPB.n122 VPB.n119 13.276
R548 VPB.n125 VPB.n122 13.276
R549 VPB.n128 VPB.n125 13.276
R550 VPB.n132 VPB.n128 13.276
R551 VPB.n234 VPB.n137 13.276
R552 VPB.n237 VPB.n234 13.276
R553 VPB.n264 VPB.n260 13.276
R554 VPB.n311 VPB.n307 13.276
R555 VPB.n42 VPB.n38 13.276
R556 VPB.n47 VPB.n46 13.276
R557 VPB.n51 VPB.n47 13.276
R558 VPB.n54 VPB.n51 13.276
R559 VPB.n63 VPB.n59 13.276
R560 VPB.n72 VPB.n68 13.276
R561 VPB.n330 VPB.n76 13.276
R562 VPB.n158 VPB.n140 13.276
R563 VPB.n140 VPB.n138 13.276
R564 VPB.n145 VPB.n143 12.796
R565 VPB.n145 VPB.n144 12.564
R566 VPB.n153 VPB.n152 12.198
R567 VPB.n153 VPB.n150 12.198
R568 VPB.n148 VPB.n147 12.198
R569 VPB.n59 VPB.n55 11.841
R570 VPB.n73 VPB.n72 11.482
R571 VPB.n46 VPB.n43 10.944
R572 VPB.n104 VPB.n103 8.97
R573 VPB.n133 VPB.n132 8.97
R574 VPB.n158 VPB.n157 7.5
R575 VPB.n143 VPB.n142 7.5
R576 VPB.n147 VPB.n146 7.5
R577 VPB.n152 VPB.n151 7.5
R578 VPB.n140 VPB.n139 7.5
R579 VPB.n155 VPB.n141 7.5
R580 VPB.n184 VPB.n183 7.5
R581 VPB.n197 VPB.n196 7.5
R582 VPB.n191 VPB.n190 7.5
R583 VPB.n193 VPB.n192 7.5
R584 VPB.n186 VPB.n185 7.5
R585 VPB.n202 VPB.n201 7.5
R586 VPB.n80 VPB.n79 7.5
R587 VPB.n93 VPB.n92 7.5
R588 VPB.n87 VPB.n86 7.5
R589 VPB.n89 VPB.n88 7.5
R590 VPB.n82 VPB.n81 7.5
R591 VPB.n98 VPB.n97 7.5
R592 VPB.n241 VPB.n240 7.5
R593 VPB.n254 VPB.n253 7.5
R594 VPB.n248 VPB.n247 7.5
R595 VPB.n250 VPB.n249 7.5
R596 VPB.n243 VPB.n242 7.5
R597 VPB.n259 VPB.n258 7.5
R598 VPB.n288 VPB.n287 7.5
R599 VPB.n301 VPB.n300 7.5
R600 VPB.n295 VPB.n294 7.5
R601 VPB.n297 VPB.n296 7.5
R602 VPB.n290 VPB.n289 7.5
R603 VPB.n306 VPB.n305 7.5
R604 VPB.n17 VPB.n16 7.5
R605 VPB.n30 VPB.n29 7.5
R606 VPB.n24 VPB.n23 7.5
R607 VPB.n26 VPB.n25 7.5
R608 VPB.n19 VPB.n18 7.5
R609 VPB.n35 VPB.n34 7.5
R610 VPB.n333 VPB.n332 7.5
R611 VPB.n12 VPB.n11 7.5
R612 VPB.n6 VPB.n5 7.5
R613 VPB.n8 VPB.n7 7.5
R614 VPB.n2 VPB.n1 7.5
R615 VPB.n335 VPB.n334 7.5
R616 VPB.n47 VPB.n35 7.176
R617 VPB.n307 VPB.n306 7.176
R618 VPB.n260 VPB.n259 7.176
R619 VPB.n115 VPB.n98 7.176
R620 VPB.n203 VPB.n202 7.176
R621 VPB.n68 VPB.n64 6.817
R622 VPB.n198 VPB.n195 6.729
R623 VPB.n194 VPB.n191 6.729
R624 VPB.n189 VPB.n186 6.729
R625 VPB.n94 VPB.n91 6.729
R626 VPB.n90 VPB.n87 6.729
R627 VPB.n85 VPB.n82 6.729
R628 VPB.n255 VPB.n252 6.729
R629 VPB.n251 VPB.n248 6.729
R630 VPB.n246 VPB.n243 6.729
R631 VPB.n302 VPB.n299 6.729
R632 VPB.n298 VPB.n295 6.729
R633 VPB.n293 VPB.n290 6.729
R634 VPB.n31 VPB.n28 6.729
R635 VPB.n27 VPB.n24 6.729
R636 VPB.n22 VPB.n19 6.729
R637 VPB.n13 VPB.n10 6.729
R638 VPB.n9 VPB.n6 6.729
R639 VPB.n4 VPB.n2 6.729
R640 VPB.n189 VPB.n188 6.728
R641 VPB.n194 VPB.n193 6.728
R642 VPB.n198 VPB.n197 6.728
R643 VPB.n201 VPB.n200 6.728
R644 VPB.n85 VPB.n84 6.728
R645 VPB.n90 VPB.n89 6.728
R646 VPB.n94 VPB.n93 6.728
R647 VPB.n97 VPB.n96 6.728
R648 VPB.n246 VPB.n245 6.728
R649 VPB.n251 VPB.n250 6.728
R650 VPB.n255 VPB.n254 6.728
R651 VPB.n258 VPB.n257 6.728
R652 VPB.n293 VPB.n292 6.728
R653 VPB.n298 VPB.n297 6.728
R654 VPB.n302 VPB.n301 6.728
R655 VPB.n305 VPB.n304 6.728
R656 VPB.n22 VPB.n21 6.728
R657 VPB.n27 VPB.n26 6.728
R658 VPB.n31 VPB.n30 6.728
R659 VPB.n34 VPB.n33 6.728
R660 VPB.n4 VPB.n3 6.728
R661 VPB.n9 VPB.n8 6.728
R662 VPB.n13 VPB.n12 6.728
R663 VPB.n336 VPB.n335 6.728
R664 VPB.n64 VPB.n63 6.458
R665 VPB.n157 VPB.n156 6.398
R666 VPB.n108 VPB.n104 4.305
R667 VPB.n137 VPB.n133 4.305
R668 VPB.n176 VPB.n172 2.691
R669 VPB.n270 VPB.n266 2.691
R670 VPB.n317 VPB.n313 2.691
R671 VPB.n166 VPB.n162 2.332
R672 VPB.n280 VPB.n276 2.332
R673 VPB.n43 VPB.n42 2.332
R674 VPB.n76 VPB.n73 1.794
R675 VPB.n55 VPB.n54 1.435
R676 VPB.n155 VPB.n148 1.402
R677 VPB.n155 VPB.n149 1.402
R678 VPB.n155 VPB.n153 1.402
R679 VPB.n155 VPB.n154 1.402
R680 VPB.n156 VPB.n155 0.735
R681 VPB.n155 VPB.n145 0.735
R682 VPB.n199 VPB.n198 0.387
R683 VPB.n199 VPB.n194 0.387
R684 VPB.n199 VPB.n189 0.387
R685 VPB.n200 VPB.n199 0.387
R686 VPB.n95 VPB.n94 0.387
R687 VPB.n95 VPB.n90 0.387
R688 VPB.n95 VPB.n85 0.387
R689 VPB.n96 VPB.n95 0.387
R690 VPB.n256 VPB.n255 0.387
R691 VPB.n256 VPB.n251 0.387
R692 VPB.n256 VPB.n246 0.387
R693 VPB.n257 VPB.n256 0.387
R694 VPB.n303 VPB.n302 0.387
R695 VPB.n303 VPB.n298 0.387
R696 VPB.n303 VPB.n293 0.387
R697 VPB.n304 VPB.n303 0.387
R698 VPB.n32 VPB.n31 0.387
R699 VPB.n32 VPB.n27 0.387
R700 VPB.n32 VPB.n22 0.387
R701 VPB.n33 VPB.n32 0.387
R702 VPB.n337 VPB.n13 0.387
R703 VPB.n337 VPB.n9 0.387
R704 VPB.n337 VPB.n4 0.387
R705 VPB.n337 VPB.n336 0.387
R706 VPB.n208 VPB.n181 0.272
R707 VPB.n225 VPB.n224 0.272
R708 VPB.n265 VPB.n238 0.272
R709 VPB.n312 VPB.n285 0.272
R710 VPB.n322 VPB.n321 0.272
R711 VPB.n329 VPB 0.198
R712 VPB.n171 VPB.n167 0.136
R713 VPB.n177 VPB.n171 0.136
R714 VPB.n181 VPB.n177 0.136
R715 VPB.n212 VPB.n208 0.136
R716 VPB.n216 VPB.n212 0.136
R717 VPB.n220 VPB.n216 0.136
R718 VPB.n221 VPB.n220 0.136
R719 VPB.n222 VPB.n221 0.136
R720 VPB.n223 VPB.n222 0.136
R721 VPB.n224 VPB.n223 0.136
R722 VPB.n226 VPB.n225 0.136
R723 VPB.n227 VPB.n226 0.136
R724 VPB.n228 VPB.n227 0.136
R725 VPB.n229 VPB.n228 0.136
R726 VPB.n230 VPB.n229 0.136
R727 VPB.n231 VPB.n230 0.136
R728 VPB.n271 VPB.n265 0.136
R729 VPB.n275 VPB.n271 0.136
R730 VPB.n281 VPB.n275 0.136
R731 VPB.n285 VPB.n281 0.136
R732 VPB.n318 VPB.n312 0.136
R733 VPB.n319 VPB.n318 0.136
R734 VPB.n320 VPB.n319 0.136
R735 VPB.n321 VPB.n320 0.136
R736 VPB.n323 VPB.n322 0.136
R737 VPB.n324 VPB.n323 0.136
R738 VPB.n325 VPB.n324 0.136
R739 VPB.n326 VPB.n325 0.136
R740 VPB.n327 VPB.n326 0.136
R741 VPB.n328 VPB.n327 0.136
R742 VPB.n329 VPB.n328 0.136
R743 VPB.n231 VPB 0.068
R744 VPB.n238 VPB 0.068
R745 a_217_1004.n4 a_217_1004.t6 512.525
R746 a_217_1004.n4 a_217_1004.t5 371.139
R747 a_217_1004.n5 a_217_1004.t7 220.263
R748 a_217_1004.n8 a_217_1004.n6 194.086
R749 a_217_1004.n6 a_217_1004.n3 162.547
R750 a_217_1004.n5 a_217_1004.n4 158.3
R751 a_217_1004.n6 a_217_1004.n5 153.043
R752 a_217_1004.n3 a_217_1004.n2 76.002
R753 a_217_1004.n8 a_217_1004.n7 30
R754 a_217_1004.n9 a_217_1004.n0 24.383
R755 a_217_1004.n9 a_217_1004.n8 23.684
R756 a_217_1004.n1 a_217_1004.t2 14.282
R757 a_217_1004.n1 a_217_1004.t1 14.282
R758 a_217_1004.n2 a_217_1004.t4 14.282
R759 a_217_1004.n2 a_217_1004.t3 14.282
R760 a_217_1004.n3 a_217_1004.n1 12.85
R761 a_851_182.n2 a_851_182.n0 362.371
R762 a_851_182.n2 a_851_182.n1 15.218
R763 a_851_182.n0 a_851_182.t1 14.282
R764 a_851_182.n0 a_851_182.t2 14.282
R765 a_851_182.n3 a_851_182.n2 12.014
R766 a_1685_1004.t1 a_1685_1004.n0 101.663
R767 a_1685_1004.n0 a_1685_1004.t3 101.661
R768 a_1685_1004.n0 a_1685_1004.t0 14.294
R769 a_1685_1004.n0 a_1685_1004.t2 14.282
R770 a_112_73.t0 a_112_73.n1 34.62
R771 a_112_73.t0 a_112_73.n0 8.137
R772 a_112_73.t0 a_112_73.n2 4.69
R773 a_1666_74.t0 a_1666_74.n1 34.62
R774 a_1666_74.t0 a_1666_74.n0 8.137
R775 a_1666_74.t0 a_1666_74.n2 4.69
C6 VPB VNB 13.92fF
C7 a_1666_74.n0 VNB 0.05fF
C8 a_1666_74.n1 VNB 0.12fF
C9 a_1666_74.n2 VNB 0.04fF
C10 a_112_73.n0 VNB 0.05fF
C11 a_112_73.n1 VNB 0.12fF
C12 a_112_73.n2 VNB 0.04fF
C13 a_1685_1004.n0 VNB 0.52fF
C14 a_851_182.n0 VNB 1.15fF
C15 a_851_182.n1 VNB 0.10fF
C16 a_851_182.n2 VNB 0.54fF
C17 a_851_182.n3 VNB 0.05fF
C18 a_217_1004.n0 VNB 0.04fF
C19 a_217_1004.n1 VNB 0.49fF
C20 a_217_1004.n2 VNB 0.58fF
C21 a_217_1004.n3 VNB 0.30fF
C22 a_217_1004.n4 VNB 0.33fF
C23 a_217_1004.t7 VNB 0.48fF
C24 a_217_1004.n5 VNB 0.53fF
C25 a_217_1004.n6 VNB 0.53fF
C26 a_217_1004.n7 VNB 0.03fF
C27 a_217_1004.n8 VNB 0.26fF
C28 a_217_1004.n9 VNB 0.05fF
C29 VPB.n0 VNB 0.03fF
C30 VPB.n1 VNB 0.04fF
C31 VPB.n2 VNB 0.02fF
C32 VPB.n3 VNB 0.14fF
C33 VPB.n5 VNB 0.02fF
C34 VPB.n6 VNB 0.02fF
C35 VPB.n7 VNB 0.02fF
C36 VPB.n8 VNB 0.02fF
C37 VPB.n10 VNB 0.02fF
C38 VPB.n11 VNB 0.02fF
C39 VPB.n12 VNB 0.02fF
C40 VPB.n14 VNB 0.10fF
C41 VPB.n15 VNB 0.02fF
C42 VPB.n16 VNB 0.02fF
C43 VPB.n17 VNB 0.02fF
C44 VPB.n18 VNB 0.04fF
C45 VPB.n19 VNB 0.02fF
C46 VPB.n20 VNB 0.17fF
C47 VPB.n21 VNB 0.04fF
C48 VPB.n23 VNB 0.02fF
C49 VPB.n24 VNB 0.02fF
C50 VPB.n25 VNB 0.02fF
C51 VPB.n26 VNB 0.02fF
C52 VPB.n28 VNB 0.02fF
C53 VPB.n29 VNB 0.02fF
C54 VPB.n30 VNB 0.02fF
C55 VPB.n32 VNB 0.27fF
C56 VPB.n34 VNB 0.03fF
C57 VPB.n35 VNB 0.02fF
C58 VPB.n36 VNB 0.16fF
C59 VPB.n37 VNB 0.02fF
C60 VPB.n38 VNB 0.02fF
C61 VPB.n39 VNB 0.14fF
C62 VPB.n40 VNB 0.19fF
C63 VPB.n41 VNB 0.02fF
C64 VPB.n42 VNB 0.01fF
C65 VPB.n43 VNB 0.06fF
C66 VPB.n44 VNB 0.27fF
C67 VPB.n45 VNB 0.01fF
C68 VPB.n46 VNB 0.02fF
C69 VPB.n47 VNB 0.03fF
C70 VPB.n48 VNB 0.03fF
C71 VPB.n49 VNB 0.27fF
C72 VPB.n50 VNB 0.01fF
C73 VPB.n51 VNB 0.02fF
C74 VPB.n52 VNB 0.23fF
C75 VPB.n53 VNB 0.02fF
C76 VPB.n54 VNB 0.01fF
C77 VPB.n55 VNB 0.05fF
C78 VPB.n56 VNB 0.14fF
C79 VPB.n57 VNB 0.16fF
C80 VPB.n58 VNB 0.02fF
C81 VPB.n59 VNB 0.02fF
C82 VPB.n60 VNB 0.14fF
C83 VPB.n61 VNB 0.15fF
C84 VPB.n62 VNB 0.02fF
C85 VPB.n63 VNB 0.02fF
C86 VPB.n64 VNB 0.02fF
C87 VPB.n65 VNB 0.14fF
C88 VPB.n66 VNB 0.15fF
C89 VPB.n67 VNB 0.02fF
C90 VPB.n68 VNB 0.02fF
C91 VPB.n69 VNB 0.14fF
C92 VPB.n70 VNB 0.16fF
C93 VPB.n71 VNB 0.02fF
C94 VPB.n72 VNB 0.02fF
C95 VPB.n73 VNB 0.06fF
C96 VPB.n74 VNB 0.24fF
C97 VPB.n75 VNB 0.02fF
C98 VPB.n76 VNB 0.01fF
C99 VPB.n77 VNB 0.10fF
C100 VPB.n78 VNB 0.02fF
C101 VPB.n79 VNB 0.02fF
C102 VPB.n80 VNB 0.02fF
C103 VPB.n81 VNB 0.04fF
C104 VPB.n82 VNB 0.02fF
C105 VPB.n83 VNB 0.19fF
C106 VPB.n84 VNB 0.04fF
C107 VPB.n86 VNB 0.02fF
C108 VPB.n87 VNB 0.02fF
C109 VPB.n88 VNB 0.02fF
C110 VPB.n89 VNB 0.02fF
C111 VPB.n91 VNB 0.02fF
C112 VPB.n92 VNB 0.02fF
C113 VPB.n93 VNB 0.02fF
C114 VPB.n95 VNB 0.27fF
C115 VPB.n97 VNB 0.03fF
C116 VPB.n98 VNB 0.02fF
C117 VPB.n99 VNB 0.10fF
C118 VPB.n100 VNB 0.14fF
C119 VPB.n101 VNB 0.15fF
C120 VPB.n102 VNB 0.02fF
C121 VPB.n103 VNB 0.02fF
C122 VPB.n104 VNB 0.03fF
C123 VPB.n105 VNB 0.14fF
C124 VPB.n106 VNB 0.16fF
C125 VPB.n107 VNB 0.02fF
C126 VPB.n108 VNB 0.02fF
C127 VPB.n109 VNB 0.24fF
C128 VPB.n110 VNB 0.02fF
C129 VPB.n111 VNB 0.02fF
C130 VPB.n112 VNB 0.27fF
C131 VPB.n113 VNB 0.01fF
C132 VPB.n114 VNB 0.02fF
C133 VPB.n115 VNB 0.03fF
C134 VPB.n116 VNB 0.03fF
C135 VPB.n117 VNB 0.27fF
C136 VPB.n118 VNB 0.01fF
C137 VPB.n119 VNB 0.02fF
C138 VPB.n120 VNB 0.27fF
C139 VPB.n121 VNB 0.02fF
C140 VPB.n122 VNB 0.02fF
C141 VPB.n123 VNB 0.27fF
C142 VPB.n124 VNB 0.02fF
C143 VPB.n125 VNB 0.02fF
C144 VPB.n126 VNB 0.27fF
C145 VPB.n127 VNB 0.02fF
C146 VPB.n128 VNB 0.02fF
C147 VPB.n129 VNB 0.14fF
C148 VPB.n130 VNB 0.15fF
C149 VPB.n131 VNB 0.02fF
C150 VPB.n132 VNB 0.02fF
C151 VPB.n133 VNB 0.03fF
C152 VPB.n134 VNB 0.14fF
C153 VPB.n135 VNB 0.16fF
C154 VPB.n136 VNB 0.02fF
C155 VPB.n137 VNB 0.02fF
C156 VPB.n138 VNB 0.02fF
C157 VPB.n139 VNB 0.02fF
C158 VPB.n140 VNB 0.02fF
C159 VPB.n141 VNB 0.11fF
C160 VPB.n142 VNB 0.03fF
C161 VPB.n143 VNB 0.02fF
C162 VPB.n144 VNB 0.05fF
C163 VPB.n145 VNB 0.01fF
C164 VPB.n146 VNB 0.02fF
C165 VPB.n147 VNB 0.02fF
C166 VPB.n150 VNB 0.02fF
C167 VPB.n151 VNB 0.02fF
C168 VPB.n152 VNB 0.02fF
C169 VPB.n155 VNB 0.46fF
C170 VPB.n157 VNB 0.04fF
C171 VPB.n158 VNB 0.04fF
C172 VPB.n159 VNB 0.27fF
C173 VPB.n160 VNB 0.03fF
C174 VPB.n161 VNB 0.03fF
C175 VPB.n162 VNB 0.06fF
C176 VPB.n163 VNB 0.14fF
C177 VPB.n164 VNB 0.19fF
C178 VPB.n165 VNB 0.02fF
C179 VPB.n166 VNB 0.01fF
C180 VPB.n167 VNB 0.07fF
C181 VPB.n168 VNB 0.16fF
C182 VPB.n169 VNB 0.02fF
C183 VPB.n170 VNB 0.02fF
C184 VPB.n171 VNB 0.02fF
C185 VPB.n172 VNB 0.06fF
C186 VPB.n173 VNB 0.14fF
C187 VPB.n174 VNB 0.19fF
C188 VPB.n175 VNB 0.02fF
C189 VPB.n176 VNB 0.01fF
C190 VPB.n177 VNB 0.02fF
C191 VPB.n178 VNB 0.27fF
C192 VPB.n179 VNB 0.01fF
C193 VPB.n180 VNB 0.02fF
C194 VPB.n181 VNB 0.04fF
C195 VPB.n182 VNB 0.02fF
C196 VPB.n183 VNB 0.02fF
C197 VPB.n184 VNB 0.02fF
C198 VPB.n185 VNB 0.04fF
C199 VPB.n186 VNB 0.02fF
C200 VPB.n187 VNB 0.17fF
C201 VPB.n188 VNB 0.04fF
C202 VPB.n190 VNB 0.02fF
C203 VPB.n191 VNB 0.02fF
C204 VPB.n192 VNB 0.02fF
C205 VPB.n193 VNB 0.02fF
C206 VPB.n195 VNB 0.02fF
C207 VPB.n196 VNB 0.02fF
C208 VPB.n197 VNB 0.02fF
C209 VPB.n199 VNB 0.27fF
C210 VPB.n201 VNB 0.03fF
C211 VPB.n202 VNB 0.02fF
C212 VPB.n203 VNB 0.03fF
C213 VPB.n204 VNB 0.03fF
C214 VPB.n205 VNB 0.27fF
C215 VPB.n206 VNB 0.01fF
C216 VPB.n207 VNB 0.02fF
C217 VPB.n208 VNB 0.04fF
C218 VPB.n209 VNB 0.27fF
C219 VPB.n210 VNB 0.02fF
C220 VPB.n211 VNB 0.02fF
C221 VPB.n212 VNB 0.02fF
C222 VPB.n213 VNB 0.27fF
C223 VPB.n214 VNB 0.02fF
C224 VPB.n215 VNB 0.02fF
C225 VPB.n216 VNB 0.02fF
C226 VPB.n217 VNB 0.27fF
C227 VPB.n218 VNB 0.02fF
C228 VPB.n219 VNB 0.02fF
C229 VPB.n220 VNB 0.02fF
C230 VPB.n221 VNB 0.02fF
C231 VPB.n222 VNB 0.02fF
C232 VPB.n223 VNB 0.02fF
C233 VPB.n224 VNB 0.04fF
C234 VPB.n225 VNB 0.04fF
C235 VPB.n226 VNB 0.02fF
C236 VPB.n227 VNB 0.02fF
C237 VPB.n228 VNB 0.02fF
C238 VPB.n229 VNB 0.02fF
C239 VPB.n230 VNB 0.02fF
C240 VPB.n231 VNB 0.02fF
C241 VPB.n232 VNB 0.24fF
C242 VPB.n233 VNB 0.02fF
C243 VPB.n234 VNB 0.02fF
C244 VPB.n235 VNB 0.27fF
C245 VPB.n236 VNB 0.01fF
C246 VPB.n237 VNB 0.02fF
C247 VPB.n238 VNB 0.03fF
C248 VPB.n239 VNB 0.02fF
C249 VPB.n240 VNB 0.02fF
C250 VPB.n241 VNB 0.02fF
C251 VPB.n242 VNB 0.04fF
C252 VPB.n243 VNB 0.02fF
C253 VPB.n244 VNB 0.16fF
C254 VPB.n245 VNB 0.04fF
C255 VPB.n247 VNB 0.02fF
C256 VPB.n248 VNB 0.02fF
C257 VPB.n249 VNB 0.02fF
C258 VPB.n250 VNB 0.02fF
C259 VPB.n252 VNB 0.02fF
C260 VPB.n253 VNB 0.02fF
C261 VPB.n254 VNB 0.02fF
C262 VPB.n256 VNB 0.27fF
C263 VPB.n258 VNB 0.03fF
C264 VPB.n259 VNB 0.02fF
C265 VPB.n260 VNB 0.03fF
C266 VPB.n261 VNB 0.03fF
C267 VPB.n262 VNB 0.27fF
C268 VPB.n263 VNB 0.01fF
C269 VPB.n264 VNB 0.02fF
C270 VPB.n265 VNB 0.04fF
C271 VPB.n266 VNB 0.06fF
C272 VPB.n267 VNB 0.14fF
C273 VPB.n268 VNB 0.19fF
C274 VPB.n269 VNB 0.02fF
C275 VPB.n270 VNB 0.01fF
C276 VPB.n271 VNB 0.02fF
C277 VPB.n272 VNB 0.16fF
C278 VPB.n273 VNB 0.02fF
C279 VPB.n274 VNB 0.02fF
C280 VPB.n275 VNB 0.02fF
C281 VPB.n276 VNB 0.06fF
C282 VPB.n277 VNB 0.14fF
C283 VPB.n278 VNB 0.19fF
C284 VPB.n279 VNB 0.02fF
C285 VPB.n280 VNB 0.01fF
C286 VPB.n281 VNB 0.02fF
C287 VPB.n282 VNB 0.27fF
C288 VPB.n283 VNB 0.01fF
C289 VPB.n284 VNB 0.02fF
C290 VPB.n285 VNB 0.04fF
C291 VPB.n286 VNB 0.02fF
C292 VPB.n287 VNB 0.02fF
C293 VPB.n288 VNB 0.02fF
C294 VPB.n289 VNB 0.04fF
C295 VPB.n290 VNB 0.02fF
C296 VPB.n291 VNB 0.13fF
C297 VPB.n292 VNB 0.04fF
C298 VPB.n294 VNB 0.02fF
C299 VPB.n295 VNB 0.02fF
C300 VPB.n296 VNB 0.02fF
C301 VPB.n297 VNB 0.02fF
C302 VPB.n299 VNB 0.02fF
C303 VPB.n300 VNB 0.02fF
C304 VPB.n301 VNB 0.02fF
C305 VPB.n303 VNB 0.27fF
C306 VPB.n305 VNB 0.03fF
C307 VPB.n306 VNB 0.02fF
C308 VPB.n307 VNB 0.03fF
C309 VPB.n308 VNB 0.03fF
C310 VPB.n309 VNB 0.27fF
C311 VPB.n310 VNB 0.01fF
C312 VPB.n311 VNB 0.02fF
C313 VPB.n312 VNB 0.04fF
C314 VPB.n313 VNB 0.06fF
C315 VPB.n314 VNB 0.14fF
C316 VPB.n315 VNB 0.19fF
C317 VPB.n316 VNB 0.02fF
C318 VPB.n317 VNB 0.01fF
C319 VPB.n318 VNB 0.02fF
C320 VPB.n319 VNB 0.02fF
C321 VPB.n320 VNB 0.02fF
C322 VPB.n321 VNB 0.04fF
C323 VPB.n322 VNB 0.04fF
C324 VPB.n323 VNB 0.02fF
C325 VPB.n324 VNB 0.02fF
C326 VPB.n325 VNB 0.02fF
C327 VPB.n326 VNB 0.02fF
C328 VPB.n327 VNB 0.02fF
C329 VPB.n328 VNB 0.02fF
C330 VPB.n329 VNB 0.03fF
C331 VPB.n330 VNB 0.03fF
C332 VPB.n331 VNB 0.02fF
C333 VPB.n332 VNB 0.02fF
C334 VPB.n333 VNB 0.02fF
C335 VPB.n334 VNB 0.04fF
C336 VPB.n335 VNB 0.04fF
C337 VPB.n337 VNB 0.43fF
C338 a_2351_1004.n0 VNB 0.52fF
C339 a_1295_182.n0 VNB 1.05fF
C340 a_1295_182.n1 VNB 0.59fF
C341 a_1295_182.n2 VNB 1.20fF
C342 a_1295_182.n3 VNB 1.28fF
C343 a_1295_182.n4 VNB 0.11fF
C344 a_1295_182.n5 VNB 0.25fF
C345 a_1295_182.n6 VNB 0.06fF
C346 a_2332_74.n0 VNB 0.02fF
C347 a_2332_74.n1 VNB 0.10fF
C348 a_2332_74.n2 VNB 0.07fF
C349 a_2332_74.n3 VNB 0.05fF
C350 a_2332_74.n4 VNB 0.00fF
C351 a_2332_74.n5 VNB 0.04fF
C352 a_2332_74.n6 VNB 0.05fF
C353 a_2332_74.n7 VNB 0.02fF
C354 a_2332_74.n8 VNB 0.05fF
C355 a_2332_74.n9 VNB 0.02fF
C356 a_2332_74.n10 VNB 0.08fF
C357 a_2332_74.n11 VNB 0.17fF
C358 a_2332_74.n12 VNB 0.09fF
C359 a_2332_74.n13 VNB 0.00fF
C360 a_1917_943.n0 VNB 0.07fF
C361 a_1917_943.n1 VNB 1.14fF
C362 a_1917_943.n2 VNB 1.24fF
C363 a_1917_943.n3 VNB 1.37fF
C364 a_1917_943.n4 VNB 1.55fF
C365 a_1917_943.n5 VNB 0.06fF
C366 a_1917_943.n6 VNB 0.46fF
C367 a_1917_943.n7 VNB 0.09fF
.ends
