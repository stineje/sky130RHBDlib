magic
tech sky130A
magscale 1 2
timestamp 1645210163
use sky130_fd_pr__hvdfl1sd2__example_55959141808143  sky130_fd_pr__hvdfl1sd2__example_55959141808143_0
timestamp 1645210163
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_0
timestamp 1645210163
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808102  sky130_fd_pr__hvdfl1sd__example_55959141808102_1
timestamp 1645210163
transform 1 0 256 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 284 267 284 267 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 7298952
string GDS_START 7297380
<< end >>
