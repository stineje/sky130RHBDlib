// File: nor2x1_pcell.spi.NOR2X1_PCELL.pxi
// Created: Tue Oct 15 15:59:23 2024
// 
simulator lang=spectre
x_PM_NOR2X1_PCELL\%noxref_1 ( N_noxref_1_c_3_p N_noxref_1_c_4_p \
 N_noxref_1_c_11_p N_noxref_1_c_16_p N_noxref_1_c_20_p N_noxref_1_c_1_p \
 N_noxref_1_c_2_p N_noxref_1_M0_noxref_s )  PM_NOR2X1_PCELL\%noxref_1
x_PM_NOR2X1_PCELL\%noxref_2 ( N_noxref_2_c_64_p N_noxref_2_c_43_p \
 N_noxref_2_c_38_n N_noxref_2_c_39_n N_noxref_2_M2_noxref_d )  \
 PM_NOR2X1_PCELL\%noxref_2
x_PM_NOR2X1_PCELL\%noxref_3 ( N_noxref_3_c_74_n N_noxref_3_c_86_n \
 N_noxref_3_M0_noxref_g N_noxref_3_M2_noxref_g N_noxref_3_M3_noxref_g \
 N_noxref_3_c_77_n N_noxref_3_c_104_p N_noxref_3_c_105_p N_noxref_3_c_79_n \
 N_noxref_3_c_81_n N_noxref_3_c_127_p N_noxref_3_c_95_p N_noxref_3_c_82_n \
 N_noxref_3_c_84_n N_noxref_3_c_93_n )  PM_NOR2X1_PCELL\%noxref_3
x_PM_NOR2X1_PCELL\%noxref_4 ( N_noxref_4_c_151_n N_noxref_4_c_139_n \
 N_noxref_4_M1_noxref_g N_noxref_4_M4_noxref_g N_noxref_4_M5_noxref_g \
 N_noxref_4_c_141_n N_noxref_4_c_161_n N_noxref_4_c_164_n N_noxref_4_c_181_p \
 N_noxref_4_c_143_n N_noxref_4_c_144_n N_noxref_4_c_145_n N_noxref_4_c_168_n \
 N_noxref_4_c_169_n N_noxref_4_c_171_n N_noxref_4_c_172_n )  \
 PM_NOR2X1_PCELL\%noxref_4
x_PM_NOR2X1_PCELL\%noxref_5 ( N_noxref_5_c_205_n N_noxref_5_c_228_n \
 N_noxref_5_c_221_n N_noxref_5_c_222_n N_noxref_5_c_209_n N_noxref_5_c_213_n \
 N_noxref_5_M0_noxref_d N_noxref_5_M1_noxref_d N_noxref_5_M4_noxref_d )  \
 PM_NOR2X1_PCELL\%noxref_5
x_PM_NOR2X1_PCELL\%noxref_6 ( N_noxref_6_c_270_n N_noxref_6_c_273_n \
 N_noxref_6_c_274_n N_noxref_6_c_275_n N_noxref_6_M2_noxref_s \
 N_noxref_6_M3_noxref_d N_noxref_6_M5_noxref_d )  PM_NOR2X1_PCELL\%noxref_6
cc_1 ( N_noxref_1_c_1_p N_noxref_2_c_38_n ) capacitor c=0.00989031f //x=0.695 \
 //y=0 //x2=0.74 //y2=7.4
cc_2 ( N_noxref_1_c_2_p N_noxref_2_c_39_n ) capacitor c=0.00989031f //x=2.635 \
 //y=0 //x2=2.59 //y2=7.4
cc_3 ( N_noxref_1_c_3_p N_noxref_3_c_74_n ) capacitor c=6.7762e-19 //x=2.59 \
 //y=0 //x2=1.11 //y2=2.08
cc_4 ( N_noxref_1_c_4_p N_noxref_3_c_74_n ) capacitor c=0.00136072f //x=1.095 \
 //y=0.53 //x2=1.11 //y2=2.08
cc_5 ( N_noxref_1_c_1_p N_noxref_3_c_74_n ) capacitor c=0.0176887f //x=0.695 \
 //y=0 //x2=1.11 //y2=2.08
cc_6 ( N_noxref_1_c_4_p N_noxref_3_c_77_n ) capacitor c=0.0122371f //x=1.095 \
 //y=0.53 //x2=0.915 //y2=0.905
cc_7 ( N_noxref_1_M0_noxref_s N_noxref_3_c_77_n ) capacitor c=0.0318086f \
 //x=0.56 //y=0.365 //x2=0.915 //y2=0.905
cc_8 ( N_noxref_1_c_4_p N_noxref_3_c_79_n ) capacitor c=2.1838e-19 //x=1.095 \
 //y=0.53 //x2=0.915 //y2=1.915
cc_9 ( N_noxref_1_c_1_p N_noxref_3_c_79_n ) capacitor c=0.0196165f //x=0.695 \
 //y=0 //x2=0.915 //y2=1.915
cc_10 ( N_noxref_1_M0_noxref_s N_noxref_3_c_81_n ) capacitor c=0.00474433f \
 //x=0.56 //y=0.365 //x2=1.29 //y2=0.75
cc_11 ( N_noxref_1_c_11_p N_noxref_3_c_82_n ) capacitor c=0.0113089f //x=1.58 \
 //y=0.53 //x2=1.445 //y2=0.905
cc_12 ( N_noxref_1_M0_noxref_s N_noxref_3_c_82_n ) capacitor c=0.00514143f \
 //x=0.56 //y=0.365 //x2=1.445 //y2=0.905
cc_13 ( N_noxref_1_M0_noxref_s N_noxref_3_c_84_n ) capacitor c=8.33128e-19 \
 //x=0.56 //y=0.365 //x2=1.445 //y2=1.25
cc_14 ( N_noxref_1_c_1_p N_noxref_4_c_139_n ) capacitor c=9.2064e-19 //x=0.695 \
 //y=0 //x2=1.85 //y2=2.08
cc_15 ( N_noxref_1_c_2_p N_noxref_4_c_139_n ) capacitor c=9.53263e-19 \
 //x=2.635 //y=0 //x2=1.85 //y2=2.08
cc_16 ( N_noxref_1_c_16_p N_noxref_4_c_141_n ) capacitor c=0.0109802f \
 //x=2.065 //y=0.53 //x2=1.885 //y2=0.905
cc_17 ( N_noxref_1_M0_noxref_s N_noxref_4_c_141_n ) capacitor c=0.00590563f \
 //x=0.56 //y=0.365 //x2=1.885 //y2=0.905
cc_18 ( N_noxref_1_M0_noxref_s N_noxref_4_c_143_n ) capacitor c=0.00466751f \
 //x=0.56 //y=0.365 //x2=2.26 //y2=0.75
cc_19 ( N_noxref_1_M0_noxref_s N_noxref_4_c_144_n ) capacitor c=0.00316186f \
 //x=0.56 //y=0.365 //x2=2.26 //y2=1.405
cc_20 ( N_noxref_1_c_20_p N_noxref_4_c_145_n ) capacitor c=0.0112321f //x=2.55 \
 //y=0.53 //x2=2.415 //y2=0.905
cc_21 ( N_noxref_1_M0_noxref_s N_noxref_4_c_145_n ) capacitor c=0.0142835f \
 //x=0.56 //y=0.365 //x2=2.415 //y2=0.905
cc_22 ( N_noxref_1_c_3_p N_noxref_5_c_205_n ) capacitor c=0.00359057f //x=2.59 \
 //y=0 //x2=2.065 //y2=1.655
cc_23 ( N_noxref_1_c_11_p N_noxref_5_c_205_n ) capacitor c=0.00381844f \
 //x=1.58 //y=0.53 //x2=2.065 //y2=1.655
cc_24 ( N_noxref_1_c_16_p N_noxref_5_c_205_n ) capacitor c=0.00323369f \
 //x=2.065 //y=0.53 //x2=2.065 //y2=1.655
cc_25 ( N_noxref_1_M0_noxref_s N_noxref_5_c_205_n ) capacitor c=0.0173679f \
 //x=0.56 //y=0.365 //x2=2.065 //y2=1.655
cc_26 ( N_noxref_1_c_3_p N_noxref_5_c_209_n ) capacitor c=0.00295442f //x=2.59 \
 //y=0 //x2=2.505 //y2=1.655
cc_27 ( N_noxref_1_c_20_p N_noxref_5_c_209_n ) capacitor c=0.0047981f //x=2.55 \
 //y=0.53 //x2=2.505 //y2=1.655
cc_28 ( N_noxref_1_c_2_p N_noxref_5_c_209_n ) capacitor c=0.0471746f //x=2.635 \
 //y=0 //x2=2.505 //y2=1.655
cc_29 ( N_noxref_1_M0_noxref_s N_noxref_5_c_209_n ) capacitor c=0.016186f \
 //x=0.56 //y=0.365 //x2=2.505 //y2=1.655
cc_30 ( N_noxref_1_c_1_p N_noxref_5_c_213_n ) capacitor c=0.00101801f \
 //x=0.695 //y=0 //x2=2.59 //y2=5.125
cc_31 ( N_noxref_1_c_3_p N_noxref_5_M0_noxref_d ) capacitor c=0.00175924f \
 //x=2.59 //y=0 //x2=0.99 //y2=0.905
cc_32 ( N_noxref_1_c_1_p N_noxref_5_M0_noxref_d ) capacitor c=0.00416273f \
 //x=0.695 //y=0 //x2=0.99 //y2=0.905
cc_33 ( N_noxref_1_c_2_p N_noxref_5_M0_noxref_d ) capacitor c=4.88559e-19 \
 //x=2.635 //y=0 //x2=0.99 //y2=0.905
cc_34 ( N_noxref_1_M0_noxref_s N_noxref_5_M0_noxref_d ) capacitor c=0.0770866f \
 //x=0.56 //y=0.365 //x2=0.99 //y2=0.905
cc_35 ( N_noxref_1_c_3_p N_noxref_5_M1_noxref_d ) capacitor c=0.00195394f \
 //x=2.59 //y=0 //x2=1.96 //y2=0.905
cc_36 ( N_noxref_1_c_2_p N_noxref_5_M1_noxref_d ) capacitor c=0.00634044f \
 //x=2.635 //y=0 //x2=1.96 //y2=0.905
cc_37 ( N_noxref_1_M0_noxref_s N_noxref_5_M1_noxref_d ) capacitor c=0.0610175f \
 //x=0.56 //y=0.365 //x2=1.96 //y2=0.905
cc_38 ( N_noxref_2_c_38_n N_noxref_3_c_74_n ) capacitor c=0.0104719f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_39 ( N_noxref_2_c_38_n N_noxref_3_c_86_n ) capacitor c=0.008636f //x=0.74 \
 //y=7.4 //x2=0.955 //y2=4.705
cc_40 ( N_noxref_2_M2_noxref_d N_noxref_3_c_86_n ) capacitor c=2.85008e-19 \
 //x=1.085 //y=5.025 //x2=0.955 //y2=4.705
cc_41 ( N_noxref_2_c_43_p N_noxref_3_M2_noxref_g ) capacitor c=0.0067918f \
 //x=1.145 //y=7.4 //x2=1.01 //y2=6.025
cc_42 ( N_noxref_2_c_38_n N_noxref_3_M2_noxref_g ) capacitor c=0.0237757f \
 //x=0.74 //y=7.4 //x2=1.01 //y2=6.025
cc_43 ( N_noxref_2_M2_noxref_d N_noxref_3_M2_noxref_g ) capacitor c=0.0156786f \
 //x=1.085 //y=5.025 //x2=1.01 //y2=6.025
cc_44 ( N_noxref_2_c_39_n N_noxref_3_M3_noxref_g ) capacitor c=0.00678153f \
 //x=2.59 //y=7.4 //x2=1.45 //y2=6.025
cc_45 ( N_noxref_2_M2_noxref_d N_noxref_3_M3_noxref_g ) capacitor c=0.0183011f \
 //x=1.085 //y=5.025 //x2=1.45 //y2=6.025
cc_46 ( N_noxref_2_c_38_n N_noxref_3_c_93_n ) capacitor c=0.00890932f //x=0.74 \
 //y=7.4 //x2=0.955 //y2=4.705
cc_47 ( N_noxref_2_c_38_n N_noxref_4_c_139_n ) capacitor c=7.02327e-19 \
 //x=0.74 //y=7.4 //x2=1.85 //y2=2.08
cc_48 ( N_noxref_2_c_39_n N_noxref_4_c_139_n ) capacitor c=6.16704e-19 \
 //x=2.59 //y=7.4 //x2=1.85 //y2=2.08
cc_49 ( N_noxref_2_c_39_n N_noxref_4_M4_noxref_g ) capacitor c=0.00513565f \
 //x=2.59 //y=7.4 //x2=1.89 //y2=6.025
cc_50 ( N_noxref_2_c_39_n N_noxref_4_M5_noxref_g ) capacitor c=0.0322288f \
 //x=2.59 //y=7.4 //x2=2.33 //y2=6.025
cc_51 ( N_noxref_2_c_39_n N_noxref_5_c_221_n ) capacitor c=9.65117e-19 \
 //x=2.59 //y=7.4 //x2=2.505 //y2=5.21
cc_52 ( N_noxref_2_c_38_n N_noxref_5_c_222_n ) capacitor c=8.9933e-19 //x=0.74 \
 //y=7.4 //x2=2.195 //y2=5.21
cc_53 ( N_noxref_2_c_38_n N_noxref_5_c_213_n ) capacitor c=0.00163766f \
 //x=0.74 //y=7.4 //x2=2.59 //y2=5.125
cc_54 ( N_noxref_2_c_39_n N_noxref_5_c_213_n ) capacitor c=0.0469841f //x=2.59 \
 //y=7.4 //x2=2.59 //y2=5.125
cc_55 ( N_noxref_2_c_39_n N_noxref_5_M4_noxref_d ) capacitor c=0.00991513f \
 //x=2.59 //y=7.4 //x2=1.965 //y2=5.025
cc_56 ( N_noxref_2_M2_noxref_d N_noxref_5_M4_noxref_d ) capacitor \
 c=0.00561178f //x=1.085 //y=5.025 //x2=1.965 //y2=5.025
cc_57 ( N_noxref_2_c_43_p N_noxref_6_c_270_n ) capacitor c=5.81484e-19 \
 //x=1.145 //y=7.4 //x2=1.585 //y2=5.21
cc_58 ( N_noxref_2_c_39_n N_noxref_6_c_270_n ) capacitor c=0.0034744f //x=2.59 \
 //y=7.4 //x2=1.585 //y2=5.21
cc_59 ( N_noxref_2_M2_noxref_d N_noxref_6_c_270_n ) capacitor c=0.0132432f \
 //x=1.085 //y=5.025 //x2=1.585 //y2=5.21
cc_60 ( N_noxref_2_c_38_n N_noxref_6_c_273_n ) capacitor c=0.0679103f //x=0.74 \
 //y=7.4 //x2=0.875 //y2=5.21
cc_61 ( N_noxref_2_c_39_n N_noxref_6_c_274_n ) capacitor c=0.00356149f \
 //x=2.59 //y=7.4 //x2=2.465 //y2=6.91
cc_62 ( N_noxref_2_c_64_p N_noxref_6_c_275_n ) capacitor c=0.0370274f //x=2.59 \
 //y=7.4 //x2=1.755 //y2=6.91
cc_63 ( N_noxref_2_c_39_n N_noxref_6_c_275_n ) capacitor c=0.059856f //x=2.59 \
 //y=7.4 //x2=1.755 //y2=6.91
cc_64 ( N_noxref_2_c_64_p N_noxref_6_M2_noxref_s ) capacitor c=0.00726388f \
 //x=2.59 //y=7.4 //x2=0.655 //y2=5.025
cc_65 ( N_noxref_2_c_43_p N_noxref_6_M2_noxref_s ) capacitor c=0.0141117f \
 //x=1.145 //y=7.4 //x2=0.655 //y2=5.025
cc_66 ( N_noxref_2_c_39_n N_noxref_6_M2_noxref_s ) capacitor c=0.00138926f \
 //x=2.59 //y=7.4 //x2=0.655 //y2=5.025
cc_67 ( N_noxref_2_M2_noxref_d N_noxref_6_M2_noxref_s ) capacitor c=0.0667021f \
 //x=1.085 //y=5.025 //x2=0.655 //y2=5.025
cc_68 ( N_noxref_2_c_38_n N_noxref_6_M3_noxref_d ) capacitor c=8.88629e-19 \
 //x=0.74 //y=7.4 //x2=1.525 //y2=5.025
cc_69 ( N_noxref_2_M2_noxref_d N_noxref_6_M3_noxref_d ) capacitor c=0.0659925f \
 //x=1.085 //y=5.025 //x2=1.525 //y2=5.025
cc_70 ( N_noxref_2_c_39_n N_noxref_6_M5_noxref_d ) capacitor c=0.0528345f \
 //x=2.59 //y=7.4 //x2=2.405 //y2=5.025
cc_71 ( N_noxref_2_M2_noxref_d N_noxref_6_M5_noxref_d ) capacitor \
 c=0.00107819f //x=1.085 //y=5.025 //x2=2.405 //y2=5.025
cc_72 ( N_noxref_3_c_86_n N_noxref_4_c_151_n ) capacitor c=0.0482889f \
 //x=0.955 //y=4.705 //x2=1.85 //y2=4.54
cc_73 ( N_noxref_3_c_95_p N_noxref_4_c_151_n ) capacitor c=0.00146509f \
 //x=1.375 //y=4.795 //x2=1.85 //y2=4.54
cc_74 ( N_noxref_3_c_93_n N_noxref_4_c_151_n ) capacitor c=0.00112871f \
 //x=0.955 //y=4.705 //x2=1.85 //y2=4.54
cc_75 ( N_noxref_3_c_74_n N_noxref_4_c_139_n ) capacitor c=0.0455438f //x=1.11 \
 //y=2.08 //x2=1.85 //y2=2.08
cc_76 ( N_noxref_3_c_79_n N_noxref_4_c_139_n ) capacitor c=0.00308814f \
 //x=0.915 //y=1.915 //x2=1.85 //y2=2.08
cc_77 ( N_noxref_3_M2_noxref_g N_noxref_4_M4_noxref_g ) capacitor c=0.0100243f \
 //x=1.01 //y=6.025 //x2=1.89 //y2=6.025
cc_78 ( N_noxref_3_M3_noxref_g N_noxref_4_M4_noxref_g ) capacitor c=0.107798f \
 //x=1.45 //y=6.025 //x2=1.89 //y2=6.025
cc_79 ( N_noxref_3_M3_noxref_g N_noxref_4_M5_noxref_g ) capacitor c=0.0094155f \
 //x=1.45 //y=6.025 //x2=2.33 //y2=6.025
cc_80 ( N_noxref_3_c_77_n N_noxref_4_c_141_n ) capacitor c=0.00125788f \
 //x=0.915 //y=0.905 //x2=1.885 //y2=0.905
cc_81 ( N_noxref_3_c_82_n N_noxref_4_c_141_n ) capacitor c=0.0126654f \
 //x=1.445 //y=0.905 //x2=1.885 //y2=0.905
cc_82 ( N_noxref_3_c_104_p N_noxref_4_c_161_n ) capacitor c=0.00148539f \
 //x=0.915 //y=1.25 //x2=1.885 //y2=1.255
cc_83 ( N_noxref_3_c_105_p N_noxref_4_c_161_n ) capacitor c=0.00105591f \
 //x=0.915 //y=1.56 //x2=1.885 //y2=1.255
cc_84 ( N_noxref_3_c_84_n N_noxref_4_c_161_n ) capacitor c=0.0126654f \
 //x=1.445 //y=1.25 //x2=1.885 //y2=1.255
cc_85 ( N_noxref_3_c_105_p N_noxref_4_c_164_n ) capacitor c=0.00109549f \
 //x=0.915 //y=1.56 //x2=1.885 //y2=1.56
cc_86 ( N_noxref_3_c_84_n N_noxref_4_c_164_n ) capacitor c=0.00886999f \
 //x=1.445 //y=1.25 //x2=1.885 //y2=1.56
cc_87 ( N_noxref_3_c_84_n N_noxref_4_c_144_n ) capacitor c=0.00123863f \
 //x=1.445 //y=1.25 //x2=2.26 //y2=1.405
cc_88 ( N_noxref_3_c_82_n N_noxref_4_c_145_n ) capacitor c=0.00132934f \
 //x=1.445 //y=0.905 //x2=2.415 //y2=0.905
cc_89 ( N_noxref_3_c_84_n N_noxref_4_c_168_n ) capacitor c=0.00150734f \
 //x=1.445 //y=1.25 //x2=2.415 //y2=1.255
cc_90 ( N_noxref_3_c_74_n N_noxref_4_c_169_n ) capacitor c=0.00307062f \
 //x=1.11 //y=2.08 //x2=1.85 //y2=2.08
cc_91 ( N_noxref_3_c_79_n N_noxref_4_c_169_n ) capacitor c=0.0179092f \
 //x=0.915 //y=1.915 //x2=1.85 //y2=2.08
cc_92 ( N_noxref_3_c_79_n N_noxref_4_c_171_n ) capacitor c=0.00577193f \
 //x=0.915 //y=1.915 //x2=1.85 //y2=1.915
cc_93 ( N_noxref_3_c_86_n N_noxref_4_c_172_n ) capacitor c=0.00336963f \
 //x=0.955 //y=4.705 //x2=1.885 //y2=4.705
cc_94 ( N_noxref_3_c_95_p N_noxref_4_c_172_n ) capacitor c=0.020271f //x=1.375 \
 //y=4.795 //x2=1.885 //y2=4.705
cc_95 ( N_noxref_3_c_93_n N_noxref_4_c_172_n ) capacitor c=0.00546725f \
 //x=0.955 //y=4.705 //x2=1.885 //y2=4.705
cc_96 ( N_noxref_3_c_84_n N_noxref_5_c_205_n ) capacitor c=0.00431513f \
 //x=1.445 //y=1.25 //x2=2.065 //y2=1.655
cc_97 ( N_noxref_3_c_74_n N_noxref_5_c_228_n ) capacitor c=0.0112169f //x=1.11 \
 //y=2.08 //x2=1.265 //y2=1.655
cc_98 ( N_noxref_3_c_79_n N_noxref_5_c_228_n ) capacitor c=0.00589082f \
 //x=0.915 //y=1.915 //x2=1.265 //y2=1.655
cc_99 ( N_noxref_3_c_74_n N_noxref_5_c_213_n ) capacitor c=0.00380766f \
 //x=1.11 //y=2.08 //x2=2.59 //y2=5.125
cc_100 ( N_noxref_3_c_77_n N_noxref_5_M0_noxref_d ) capacitor c=0.0013184f \
 //x=0.915 //y=0.905 //x2=0.99 //y2=0.905
cc_101 ( N_noxref_3_c_104_p N_noxref_5_M0_noxref_d ) capacitor c=0.0034598f \
 //x=0.915 //y=1.25 //x2=0.99 //y2=0.905
cc_102 ( N_noxref_3_c_105_p N_noxref_5_M0_noxref_d ) capacitor c=0.00300148f \
 //x=0.915 //y=1.56 //x2=0.99 //y2=0.905
cc_103 ( N_noxref_3_c_79_n N_noxref_5_M0_noxref_d ) capacitor c=0.00273686f \
 //x=0.915 //y=1.915 //x2=0.99 //y2=0.905
cc_104 ( N_noxref_3_c_81_n N_noxref_5_M0_noxref_d ) capacitor c=0.00241102f \
 //x=1.29 //y=0.75 //x2=0.99 //y2=0.905
cc_105 ( N_noxref_3_c_127_p N_noxref_5_M0_noxref_d ) capacitor c=0.0123304f \
 //x=1.29 //y=1.405 //x2=0.99 //y2=0.905
cc_106 ( N_noxref_3_c_82_n N_noxref_5_M0_noxref_d ) capacitor c=0.00219619f \
 //x=1.445 //y=0.905 //x2=0.99 //y2=0.905
cc_107 ( N_noxref_3_c_84_n N_noxref_5_M0_noxref_d ) capacitor c=0.00603828f \
 //x=1.445 //y=1.25 //x2=0.99 //y2=0.905
cc_108 ( N_noxref_3_c_86_n N_noxref_6_c_270_n ) capacitor c=0.00630079f \
 //x=0.955 //y=4.705 //x2=1.585 //y2=5.21
cc_109 ( N_noxref_3_M2_noxref_g N_noxref_6_c_270_n ) capacitor c=0.0182669f \
 //x=1.01 //y=6.025 //x2=1.585 //y2=5.21
cc_110 ( N_noxref_3_M3_noxref_g N_noxref_6_c_270_n ) capacitor c=0.0204082f \
 //x=1.45 //y=6.025 //x2=1.585 //y2=5.21
cc_111 ( N_noxref_3_c_95_p N_noxref_6_c_270_n ) capacitor c=0.00365818f \
 //x=1.375 //y=4.795 //x2=1.585 //y2=5.21
cc_112 ( N_noxref_3_c_93_n N_noxref_6_c_270_n ) capacitor c=0.0017421f \
 //x=0.955 //y=4.705 //x2=1.585 //y2=5.21
cc_113 ( N_noxref_3_c_86_n N_noxref_6_c_273_n ) capacitor c=0.0118415f \
 //x=0.955 //y=4.705 //x2=0.875 //y2=5.21
cc_114 ( N_noxref_3_c_93_n N_noxref_6_c_273_n ) capacitor c=0.00613395f \
 //x=0.955 //y=4.705 //x2=0.875 //y2=5.21
cc_115 ( N_noxref_3_M2_noxref_g N_noxref_6_M2_noxref_s ) capacitor \
 c=0.0473218f //x=1.01 //y=6.025 //x2=0.655 //y2=5.025
cc_116 ( N_noxref_3_M3_noxref_g N_noxref_6_M3_noxref_d ) capacitor \
 c=0.0170604f //x=1.45 //y=6.025 //x2=1.525 //y2=5.025
cc_117 ( N_noxref_4_c_139_n N_noxref_5_c_205_n ) capacitor c=0.0162392f \
 //x=1.85 //y=2.08 //x2=2.065 //y2=1.655
cc_118 ( N_noxref_4_c_164_n N_noxref_5_c_205_n ) capacitor c=0.00218915f \
 //x=1.885 //y=1.56 //x2=2.065 //y2=1.655
cc_119 ( N_noxref_4_c_169_n N_noxref_5_c_205_n ) capacitor c=0.00633758f \
 //x=1.85 //y=2.08 //x2=2.065 //y2=1.655
cc_120 ( N_noxref_4_c_171_n N_noxref_5_c_205_n ) capacitor c=0.0189958f \
 //x=1.85 //y=1.915 //x2=2.065 //y2=1.655
cc_121 ( N_noxref_4_M5_noxref_g N_noxref_5_c_221_n ) capacitor c=0.0217751f \
 //x=2.33 //y=6.025 //x2=2.505 //y2=5.21
cc_122 ( N_noxref_4_M4_noxref_g N_noxref_5_c_222_n ) capacitor c=0.0132788f \
 //x=1.89 //y=6.025 //x2=2.195 //y2=5.21
cc_123 ( N_noxref_4_c_181_p N_noxref_5_c_222_n ) capacitor c=0.00417892f \
 //x=2.255 //y=4.795 //x2=2.195 //y2=5.21
cc_124 ( N_noxref_4_c_144_n N_noxref_5_c_209_n ) capacitor c=0.00801563f \
 //x=2.26 //y=1.405 //x2=2.505 //y2=1.655
cc_125 ( N_noxref_4_c_151_n N_noxref_5_c_213_n ) capacitor c=0.0102183f \
 //x=1.85 //y=4.54 //x2=2.59 //y2=5.125
cc_126 ( N_noxref_4_c_139_n N_noxref_5_c_213_n ) capacitor c=0.0842481f \
 //x=1.85 //y=2.08 //x2=2.59 //y2=5.125
cc_127 ( N_noxref_4_c_181_p N_noxref_5_c_213_n ) capacitor c=0.0144455f \
 //x=2.255 //y=4.795 //x2=2.59 //y2=5.125
cc_128 ( N_noxref_4_c_169_n N_noxref_5_c_213_n ) capacitor c=0.00877984f \
 //x=1.85 //y=2.08 //x2=2.59 //y2=5.125
cc_129 ( N_noxref_4_c_171_n N_noxref_5_c_213_n ) capacitor c=0.00306024f \
 //x=1.85 //y=1.915 //x2=2.59 //y2=5.125
cc_130 ( N_noxref_4_c_172_n N_noxref_5_c_213_n ) capacitor c=0.00537091f \
 //x=1.885 //y=4.705 //x2=2.59 //y2=5.125
cc_131 ( N_noxref_4_c_164_n N_noxref_5_M0_noxref_d ) capacitor c=0.00148728f \
 //x=1.885 //y=1.56 //x2=0.99 //y2=0.905
cc_132 ( N_noxref_4_c_141_n N_noxref_5_M1_noxref_d ) capacitor c=0.00226395f \
 //x=1.885 //y=0.905 //x2=1.96 //y2=0.905
cc_133 ( N_noxref_4_c_161_n N_noxref_5_M1_noxref_d ) capacitor c=0.0035101f \
 //x=1.885 //y=1.255 //x2=1.96 //y2=0.905
cc_134 ( N_noxref_4_c_164_n N_noxref_5_M1_noxref_d ) capacitor c=0.00546704f \
 //x=1.885 //y=1.56 //x2=1.96 //y2=0.905
cc_135 ( N_noxref_4_c_143_n N_noxref_5_M1_noxref_d ) capacitor c=0.00241102f \
 //x=2.26 //y=0.75 //x2=1.96 //y2=0.905
cc_136 ( N_noxref_4_c_144_n N_noxref_5_M1_noxref_d ) capacitor c=0.0158021f \
 //x=2.26 //y=1.405 //x2=1.96 //y2=0.905
cc_137 ( N_noxref_4_c_145_n N_noxref_5_M1_noxref_d ) capacitor c=0.00132831f \
 //x=2.415 //y=0.905 //x2=1.96 //y2=0.905
cc_138 ( N_noxref_4_c_168_n N_noxref_5_M1_noxref_d ) capacitor c=0.0035101f \
 //x=2.415 //y=1.255 //x2=1.96 //y2=0.905
cc_139 ( N_noxref_4_c_171_n N_noxref_5_M1_noxref_d ) capacitor c=3.4952e-19 \
 //x=1.85 //y=1.915 //x2=1.96 //y2=0.905
cc_140 ( N_noxref_4_M5_noxref_g N_noxref_5_M4_noxref_d ) capacitor \
 c=0.0136385f //x=2.33 //y=6.025 //x2=1.965 //y2=5.025
cc_141 ( N_noxref_4_M4_noxref_g N_noxref_6_c_270_n ) capacitor c=0.0170604f \
 //x=1.89 //y=6.025 //x2=1.585 //y2=5.21
cc_142 ( N_noxref_4_c_172_n N_noxref_6_c_270_n ) capacitor c=2.3112e-19 \
 //x=1.885 //y=4.705 //x2=1.585 //y2=5.21
cc_143 ( N_noxref_4_c_151_n N_noxref_6_c_274_n ) capacitor c=0.00109004f \
 //x=1.85 //y=4.54 //x2=2.465 //y2=6.91
cc_144 ( N_noxref_4_M4_noxref_g N_noxref_6_c_274_n ) capacitor c=0.0148484f \
 //x=1.89 //y=6.025 //x2=2.465 //y2=6.91
cc_145 ( N_noxref_4_M5_noxref_g N_noxref_6_c_274_n ) capacitor c=0.0163196f \
 //x=2.33 //y=6.025 //x2=2.465 //y2=6.91
cc_146 ( N_noxref_4_M5_noxref_g N_noxref_6_M5_noxref_d ) capacitor \
 c=0.0351101f //x=2.33 //y=6.025 //x2=2.405 //y2=5.025
cc_147 ( N_noxref_5_c_222_n N_noxref_6_c_270_n ) capacitor c=0.0348754f \
 //x=2.195 //y=5.21 //x2=1.585 //y2=5.21
cc_148 ( N_noxref_5_c_221_n N_noxref_6_c_274_n ) capacitor c=0.00194034f \
 //x=2.505 //y=5.21 //x2=2.465 //y2=6.91
cc_149 ( N_noxref_5_M4_noxref_d N_noxref_6_c_274_n ) capacitor c=0.0118172f \
 //x=1.965 //y=5.025 //x2=2.465 //y2=6.91
cc_150 ( N_noxref_5_M4_noxref_d N_noxref_6_M2_noxref_s ) capacitor \
 c=0.00107541f //x=1.965 //y=5.025 //x2=0.655 //y2=5.025
cc_151 ( N_noxref_5_M4_noxref_d N_noxref_6_M3_noxref_d ) capacitor \
 c=0.0348754f //x=1.965 //y=5.025 //x2=1.525 //y2=5.025
cc_152 ( N_noxref_5_c_221_n N_noxref_6_M5_noxref_d ) capacitor c=0.0164221f \
 //x=2.505 //y=5.21 //x2=2.405 //y2=5.025
cc_153 ( N_noxref_5_M4_noxref_d N_noxref_6_M5_noxref_d ) capacitor \
 c=0.0458293f //x=1.965 //y=5.025 //x2=2.405 //y2=5.025
