magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 8 67 1103 203
rect 29 -17 63 67
rect 285 21 1103 67
<< locali >>
rect 85 199 155 339
rect 189 199 247 265
rect 559 357 623 475
rect 559 290 601 357
rect 775 325 825 493
rect 943 325 993 493
rect 535 199 601 290
rect 647 289 734 323
rect 775 291 1087 325
rect 647 199 681 289
rect 1041 181 1087 291
rect 783 145 1087 181
rect 783 51 833 145
rect 935 51 1001 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 407 69 491
rect 103 441 169 527
rect 225 459 489 493
rect 225 407 259 459
rect 17 373 259 407
rect 302 391 421 425
rect 17 165 51 373
rect 198 305 319 339
rect 281 265 319 305
rect 281 199 339 265
rect 281 165 319 199
rect 17 90 80 165
rect 131 17 165 165
rect 215 131 319 165
rect 387 165 421 391
rect 455 199 489 459
rect 680 359 730 527
rect 859 359 909 527
rect 1027 359 1077 527
rect 715 215 1007 249
rect 715 165 749 215
rect 387 131 749 165
rect 215 90 249 131
rect 303 17 369 96
rect 419 61 453 131
rect 493 17 559 97
rect 593 61 627 131
rect 671 17 747 97
rect 867 17 901 111
rect 1035 17 1069 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 647 199 681 289 6 A
port 1 nsew signal input
rlabel locali s 647 289 734 323 6 A
port 1 nsew signal input
rlabel locali s 535 199 601 290 6 B
port 2 nsew signal input
rlabel locali s 559 290 601 357 6 B
port 2 nsew signal input
rlabel locali s 559 357 623 475 6 B
port 2 nsew signal input
rlabel locali s 85 199 155 339 6 C_N
port 3 nsew signal input
rlabel locali s 189 199 247 265 6 D_N
port 4 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 285 21 1103 67 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 29 -17 63 67 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 8 67 1103 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 935 51 1001 145 6 X
port 9 nsew signal output
rlabel locali s 783 51 833 145 6 X
port 9 nsew signal output
rlabel locali s 783 145 1087 181 6 X
port 9 nsew signal output
rlabel locali s 1041 181 1087 291 6 X
port 9 nsew signal output
rlabel locali s 775 291 1087 325 6 X
port 9 nsew signal output
rlabel locali s 943 325 993 493 6 X
port 9 nsew signal output
rlabel locali s 775 325 825 493 6 X
port 9 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1104 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 8888
string GDS_START 130
<< end >>
