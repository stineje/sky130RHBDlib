// File: TMRDFFQNX1.spi.TMRDFFQNX1.pxi
// Created: Tue Oct 15 15:51:34 2024
// 
simulator lang=spectre
x_PM_TMRDFFQNX1\%GND ( GND N_GND_c_23_p N_GND_c_113_p N_GND_c_1_p N_GND_c_24_p \
 N_GND_c_25_p N_GND_c_74_p N_GND_c_33_p N_GND_c_40_p N_GND_c_50_p N_GND_c_57_p \
 N_GND_c_77_p N_GND_c_84_p N_GND_c_91_p N_GND_c_98_p N_GND_c_206_p \
 N_GND_c_213_p N_GND_c_162_p N_GND_c_169_p N_GND_c_130_p N_GND_c_137_p \
 N_GND_c_146_p N_GND_c_153_p N_GND_c_172_p N_GND_c_179_p N_GND_c_186_p \
 N_GND_c_193_p N_GND_c_350_p N_GND_c_357_p N_GND_c_306_p N_GND_c_313_p \
 N_GND_c_265_p N_GND_c_272_p N_GND_c_281_p N_GND_c_288_p N_GND_c_316_p \
 N_GND_c_323_p N_GND_c_330_p N_GND_c_337_p N_GND_c_372_p N_GND_c_379_p \
 N_GND_c_382_p N_GND_c_388_p N_GND_c_469_p N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p \
 N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p N_GND_c_8_p N_GND_c_9_p N_GND_c_10_p \
 N_GND_c_11_p N_GND_c_12_p N_GND_c_13_p N_GND_c_14_p N_GND_c_15_p N_GND_c_16_p \
 N_GND_c_17_p N_GND_c_18_p N_GND_c_19_p N_GND_c_20_p N_GND_c_21_p N_GND_c_22_p \
 N_GND_M0_noxref_d N_GND_M3_noxref_d N_GND_M5_noxref_d N_GND_M7_noxref_d \
 N_GND_M9_noxref_d N_GND_M11_noxref_d N_GND_M13_noxref_d N_GND_M16_noxref_d \
 N_GND_M18_noxref_d N_GND_M20_noxref_d N_GND_M22_noxref_d N_GND_M24_noxref_d \
 N_GND_M26_noxref_d N_GND_M29_noxref_d N_GND_M31_noxref_d N_GND_M33_noxref_d \
 N_GND_M35_noxref_d N_GND_M37_noxref_d N_GND_M39_noxref_d N_GND_M41_noxref_d \
 N_GND_M43_noxref_d )  PM_TMRDFFQNX1\%GND
x_PM_TMRDFFQNX1\%VDD ( VDD N_VDD_c_960_p N_VDD_c_937_n N_VDD_c_1027_p \
 N_VDD_c_1028_p N_VDD_c_975_p N_VDD_c_1038_p N_VDD_c_1447_p N_VDD_c_961_p \
 N_VDD_c_962_p N_VDD_c_1449_p N_VDD_c_1450_p N_VDD_c_973_p N_VDD_c_997_p \
 N_VDD_c_1452_p N_VDD_c_1453_p N_VDD_c_1008_p N_VDD_c_1121_p N_VDD_c_1465_p \
 N_VDD_c_1466_p N_VDD_c_1045_p N_VDD_c_1074_p N_VDD_c_1491_p N_VDD_c_1492_p \
 N_VDD_c_1085_p N_VDD_c_1142_p N_VDD_c_1494_p N_VDD_c_1495_p N_VDD_c_1228_p \
 N_VDD_c_1229_p N_VDD_c_1176_p N_VDD_c_1239_p N_VDD_c_1474_p N_VDD_c_1162_p \
 N_VDD_c_1163_p N_VDD_c_1476_p N_VDD_c_1477_p N_VDD_c_1174_p N_VDD_c_1198_p \
 N_VDD_c_1479_p N_VDD_c_1480_p N_VDD_c_1209_p N_VDD_c_1318_p N_VDD_c_1504_p \
 N_VDD_c_1505_p N_VDD_c_1246_p N_VDD_c_1275_p N_VDD_c_1507_p N_VDD_c_1508_p \
 N_VDD_c_1286_p N_VDD_c_1339_p N_VDD_c_1510_p N_VDD_c_1511_p N_VDD_c_1512_p \
 N_VDD_c_1572_p N_VDD_c_1394_p N_VDD_c_1524_p N_VDD_c_1525_p N_VDD_c_1380_p \
 N_VDD_c_1373_p N_VDD_c_1527_p N_VDD_c_1528_p N_VDD_c_1392_p N_VDD_c_1416_p \
 N_VDD_c_1530_p N_VDD_c_1531_p N_VDD_c_1427_p N_VDD_c_1576_p N_VDD_c_1673_p \
 N_VDD_c_1674_p N_VDD_c_1600_p N_VDD_c_1638_p N_VDD_c_1628_p N_VDD_c_1629_p \
 N_VDD_c_1630_p N_VDD_c_1710_p N_VDD_c_1739_p N_VDD_c_1734_p N_VDD_c_1817_p \
 N_VDD_c_1838_p N_VDD_c_1772_p N_VDD_c_938_n N_VDD_c_939_n N_VDD_c_940_n \
 N_VDD_c_941_n N_VDD_c_942_n N_VDD_c_943_n N_VDD_c_944_n N_VDD_c_945_n \
 N_VDD_c_946_n N_VDD_c_947_n N_VDD_c_948_n N_VDD_c_949_n N_VDD_c_950_n \
 N_VDD_c_951_n N_VDD_c_952_n N_VDD_c_953_n N_VDD_c_954_n N_VDD_c_955_n \
 N_VDD_c_956_n N_VDD_c_957_n N_VDD_c_958_n N_VDD_M45_noxref_s \
 N_VDD_M46_noxref_d N_VDD_M48_noxref_d N_VDD_M50_noxref_d N_VDD_M51_noxref_s \
 N_VDD_M52_noxref_d N_VDD_M54_noxref_d N_VDD_M55_noxref_s N_VDD_M56_noxref_d \
 N_VDD_M58_noxref_d N_VDD_M59_noxref_s N_VDD_M60_noxref_d N_VDD_M62_noxref_d \
 N_VDD_M63_noxref_s N_VDD_M64_noxref_d N_VDD_M66_noxref_d N_VDD_M67_noxref_s \
 N_VDD_M68_noxref_d N_VDD_M70_noxref_d N_VDD_M71_noxref_s N_VDD_M72_noxref_d \
 N_VDD_M74_noxref_d N_VDD_M76_noxref_d N_VDD_M77_noxref_s N_VDD_M78_noxref_d \
 N_VDD_M80_noxref_d N_VDD_M81_noxref_s N_VDD_M82_noxref_d N_VDD_M84_noxref_d \
 N_VDD_M85_noxref_s N_VDD_M86_noxref_d N_VDD_M88_noxref_d N_VDD_M89_noxref_s \
 N_VDD_M90_noxref_d N_VDD_M92_noxref_d N_VDD_M93_noxref_s N_VDD_M94_noxref_d \
 N_VDD_M96_noxref_d N_VDD_M97_noxref_s N_VDD_M98_noxref_d N_VDD_M100_noxref_d \
 N_VDD_M102_noxref_d N_VDD_M103_noxref_s N_VDD_M104_noxref_d \
 N_VDD_M106_noxref_d N_VDD_M107_noxref_s N_VDD_M108_noxref_d \
 N_VDD_M110_noxref_d N_VDD_M111_noxref_s N_VDD_M112_noxref_d \
 N_VDD_M114_noxref_d N_VDD_M115_noxref_s N_VDD_M116_noxref_d \
 N_VDD_M118_noxref_d N_VDD_M119_noxref_s N_VDD_M120_noxref_d \
 N_VDD_M122_noxref_d N_VDD_M123_noxref_s N_VDD_M124_noxref_d \
 N_VDD_M126_noxref_d )  PM_TMRDFFQNX1\%VDD
x_PM_TMRDFFQNX1\%noxref_3 ( N_noxref_3_c_1935_n N_noxref_3_c_1939_n \
 N_noxref_3_c_1940_n N_noxref_3_c_2007_p N_noxref_3_c_1941_n \
 N_noxref_3_c_1959_n N_noxref_3_c_1963_n N_noxref_3_c_1965_n \
 N_noxref_3_c_1942_n N_noxref_3_c_2079_p N_noxref_3_c_1943_n \
 N_noxref_3_c_1944_n N_noxref_3_c_2099_p N_noxref_3_M2_noxref_g \
 N_noxref_3_M5_noxref_g N_noxref_3_M49_noxref_g N_noxref_3_M50_noxref_g \
 N_noxref_3_M55_noxref_g N_noxref_3_M56_noxref_g N_noxref_3_c_2034_p \
 N_noxref_3_c_2035_p N_noxref_3_c_2036_p N_noxref_3_c_2037_p \
 N_noxref_3_c_2014_p N_noxref_3_c_2039_p N_noxref_3_c_2015_p \
 N_noxref_3_c_1945_n N_noxref_3_c_1947_n N_noxref_3_c_1948_n \
 N_noxref_3_c_1949_n N_noxref_3_c_1950_n N_noxref_3_c_1951_n \
 N_noxref_3_c_1952_n N_noxref_3_c_1954_n N_noxref_3_c_2021_p \
 N_noxref_3_c_2022_p N_noxref_3_c_2013_p N_noxref_3_c_1982_n \
 N_noxref_3_M4_noxref_d N_noxref_3_M51_noxref_d N_noxref_3_M53_noxref_d )  \
 PM_TMRDFFQNX1\%noxref_3
x_PM_TMRDFFQNX1\%noxref_4 ( N_noxref_4_c_2167_n N_noxref_4_c_2215_n \
 N_noxref_4_c_2184_n N_noxref_4_c_2188_n N_noxref_4_c_2190_n \
 N_noxref_4_c_2168_n N_noxref_4_c_2266_p N_noxref_4_c_2169_n \
 N_noxref_4_c_2170_n N_noxref_4_c_2251_p N_noxref_4_M7_noxref_g \
 N_noxref_4_M59_noxref_g N_noxref_4_M60_noxref_g N_noxref_4_c_2171_n \
 N_noxref_4_c_2173_n N_noxref_4_c_2174_n N_noxref_4_c_2175_n \
 N_noxref_4_c_2176_n N_noxref_4_c_2177_n N_noxref_4_c_2178_n \
 N_noxref_4_c_2180_n N_noxref_4_c_2203_n N_noxref_4_M6_noxref_d \
 N_noxref_4_M55_noxref_d N_noxref_4_M57_noxref_d )  PM_TMRDFFQNX1\%noxref_4
x_PM_TMRDFFQNX1\%noxref_5 ( N_noxref_5_c_2388_n N_noxref_5_c_2389_n \
 N_noxref_5_c_2317_n N_noxref_5_c_2396_n N_noxref_5_c_2342_n \
 N_noxref_5_c_2346_n N_noxref_5_c_2348_n N_noxref_5_c_2352_n \
 N_noxref_5_c_2318_n N_noxref_5_c_2402_n N_noxref_5_c_2356_n \
 N_noxref_5_c_2319_n N_noxref_5_c_2320_n N_noxref_5_c_2497_p \
 N_noxref_5_c_2414_n N_noxref_5_M3_noxref_g N_noxref_5_M9_noxref_g \
 N_noxref_5_M51_noxref_g N_noxref_5_M52_noxref_g N_noxref_5_M63_noxref_g \
 N_noxref_5_M64_noxref_g N_noxref_5_c_2321_n N_noxref_5_c_2323_n \
 N_noxref_5_c_2324_n N_noxref_5_c_2325_n N_noxref_5_c_2326_n \
 N_noxref_5_c_2327_n N_noxref_5_c_2328_n N_noxref_5_c_2330_n \
 N_noxref_5_c_2331_n N_noxref_5_c_2333_n N_noxref_5_c_2334_n \
 N_noxref_5_c_2335_n N_noxref_5_c_2336_n N_noxref_5_c_2337_n \
 N_noxref_5_c_2338_n N_noxref_5_c_2340_n N_noxref_5_c_2371_n \
 N_noxref_5_c_2372_n N_noxref_5_M2_noxref_d N_noxref_5_M45_noxref_d \
 N_noxref_5_M47_noxref_d N_noxref_5_M49_noxref_d )  PM_TMRDFFQNX1\%noxref_5
x_PM_TMRDFFQNX1\%noxref_6 ( N_noxref_6_c_2619_p N_noxref_6_c_2612_n \
 N_noxref_6_c_2581_n N_noxref_6_c_2585_n N_noxref_6_c_2587_n \
 N_noxref_6_c_2565_n N_noxref_6_c_2649_p N_noxref_6_c_2566_n \
 N_noxref_6_c_2567_n N_noxref_6_c_2685_p N_noxref_6_M11_noxref_g \
 N_noxref_6_M67_noxref_g N_noxref_6_M68_noxref_g N_noxref_6_c_2568_n \
 N_noxref_6_c_2570_n N_noxref_6_c_2571_n N_noxref_6_c_2572_n \
 N_noxref_6_c_2573_n N_noxref_6_c_2574_n N_noxref_6_c_2575_n \
 N_noxref_6_c_2577_n N_noxref_6_c_2600_n N_noxref_6_M10_noxref_d \
 N_noxref_6_M63_noxref_d N_noxref_6_M65_noxref_d )  PM_TMRDFFQNX1\%noxref_6
x_PM_TMRDFFQNX1\%noxref_7 ( N_noxref_7_c_2715_n N_noxref_7_c_2716_n \
 N_noxref_7_c_2744_n N_noxref_7_c_2801_n N_noxref_7_c_2745_n \
 N_noxref_7_c_2747_n N_noxref_7_c_2717_n N_noxref_7_c_2803_n \
 N_noxref_7_c_2718_n N_noxref_7_c_2753_n N_noxref_7_c_2757_n \
 N_noxref_7_c_2759_n N_noxref_7_c_2720_n N_noxref_7_c_2919_p \
 N_noxref_7_c_2721_n N_noxref_7_c_2888_n N_noxref_7_c_2722_n \
 N_noxref_7_c_2981_p N_noxref_7_M0_noxref_g N_noxref_7_M6_noxref_g \
 N_noxref_7_M12_noxref_g N_noxref_7_M45_noxref_g N_noxref_7_M46_noxref_g \
 N_noxref_7_M57_noxref_g N_noxref_7_M58_noxref_g N_noxref_7_M69_noxref_g \
 N_noxref_7_M70_noxref_g N_noxref_7_c_2724_n N_noxref_7_c_2726_n \
 N_noxref_7_c_2727_n N_noxref_7_c_2728_n N_noxref_7_c_2729_n \
 N_noxref_7_c_2730_n N_noxref_7_c_2731_n N_noxref_7_c_2733_n \
 N_noxref_7_c_2882_n N_noxref_7_c_2781_n N_noxref_7_c_2812_n \
 N_noxref_7_c_2815_n N_noxref_7_c_2817_n N_noxref_7_c_2849_n \
 N_noxref_7_c_2851_n N_noxref_7_c_2852_n N_noxref_7_c_2820_n \
 N_noxref_7_c_2821_n N_noxref_7_c_2897_n N_noxref_7_c_2900_n \
 N_noxref_7_c_2902_n N_noxref_7_c_2946_p N_noxref_7_c_3020_p \
 N_noxref_7_c_3007_p N_noxref_7_c_2905_n N_noxref_7_c_2906_n \
 N_noxref_7_c_2822_n N_noxref_7_c_2858_n N_noxref_7_c_2824_n \
 N_noxref_7_c_2907_n N_noxref_7_c_3014_p N_noxref_7_c_2909_n \
 N_noxref_7_M8_noxref_d N_noxref_7_M59_noxref_d N_noxref_7_M61_noxref_d )  \
 PM_TMRDFFQNX1\%noxref_7
x_PM_TMRDFFQNX1\%noxref_8 ( N_noxref_8_c_3129_p N_noxref_8_c_3144_p \
 N_noxref_8_c_3121_p N_noxref_8_c_3134_p N_noxref_8_c_3068_n \
 N_noxref_8_c_3086_n N_noxref_8_c_3090_n N_noxref_8_c_3092_n \
 N_noxref_8_c_3069_n N_noxref_8_c_3209_p N_noxref_8_c_3070_n \
 N_noxref_8_c_3071_n N_noxref_8_c_3229_p N_noxref_8_M15_noxref_g \
 N_noxref_8_M18_noxref_g N_noxref_8_M75_noxref_g N_noxref_8_M76_noxref_g \
 N_noxref_8_M81_noxref_g N_noxref_8_M82_noxref_g N_noxref_8_c_3160_p \
 N_noxref_8_c_3161_p N_noxref_8_c_3162_p N_noxref_8_c_3163_p \
 N_noxref_8_c_3141_p N_noxref_8_c_3165_p N_noxref_8_c_3142_p \
 N_noxref_8_c_3072_n N_noxref_8_c_3074_n N_noxref_8_c_3075_n \
 N_noxref_8_c_3076_n N_noxref_8_c_3077_n N_noxref_8_c_3078_n \
 N_noxref_8_c_3079_n N_noxref_8_c_3081_n N_noxref_8_c_3147_p \
 N_noxref_8_c_3148_p N_noxref_8_c_3140_p N_noxref_8_c_3109_n \
 N_noxref_8_M17_noxref_d N_noxref_8_M77_noxref_d N_noxref_8_M79_noxref_d )  \
 PM_TMRDFFQNX1\%noxref_8
x_PM_TMRDFFQNX1\%noxref_9 ( N_noxref_9_c_3355_p N_noxref_9_c_3347_n \
 N_noxref_9_c_3316_n N_noxref_9_c_3320_n N_noxref_9_c_3322_n \
 N_noxref_9_c_3300_n N_noxref_9_c_3398_p N_noxref_9_c_3301_n \
 N_noxref_9_c_3302_n N_noxref_9_c_3383_p N_noxref_9_M20_noxref_g \
 N_noxref_9_M85_noxref_g N_noxref_9_M86_noxref_g N_noxref_9_c_3303_n \
 N_noxref_9_c_3305_n N_noxref_9_c_3306_n N_noxref_9_c_3307_n \
 N_noxref_9_c_3308_n N_noxref_9_c_3309_n N_noxref_9_c_3310_n \
 N_noxref_9_c_3312_n N_noxref_9_c_3335_n N_noxref_9_M19_noxref_d \
 N_noxref_9_M81_noxref_d N_noxref_9_M83_noxref_d )  PM_TMRDFFQNX1\%noxref_9
x_PM_TMRDFFQNX1\%noxref_10 ( N_noxref_10_c_3523_n N_noxref_10_c_3524_n \
 N_noxref_10_c_3526_n N_noxref_10_c_3531_n N_noxref_10_c_3477_n \
 N_noxref_10_c_3481_n N_noxref_10_c_3483_n N_noxref_10_c_3487_n \
 N_noxref_10_c_3453_n N_noxref_10_c_3594_p N_noxref_10_c_3491_n \
 N_noxref_10_c_3454_n N_noxref_10_c_3455_n N_noxref_10_c_3633_p \
 N_noxref_10_c_3548_n N_noxref_10_M16_noxref_g N_noxref_10_M22_noxref_g \
 N_noxref_10_M77_noxref_g N_noxref_10_M78_noxref_g N_noxref_10_M89_noxref_g \
 N_noxref_10_M90_noxref_g N_noxref_10_c_3456_n N_noxref_10_c_3458_n \
 N_noxref_10_c_3459_n N_noxref_10_c_3460_n N_noxref_10_c_3461_n \
 N_noxref_10_c_3462_n N_noxref_10_c_3463_n N_noxref_10_c_3465_n \
 N_noxref_10_c_3466_n N_noxref_10_c_3468_n N_noxref_10_c_3469_n \
 N_noxref_10_c_3470_n N_noxref_10_c_3471_n N_noxref_10_c_3472_n \
 N_noxref_10_c_3473_n N_noxref_10_c_3475_n N_noxref_10_c_3506_n \
 N_noxref_10_c_3507_n N_noxref_10_M15_noxref_d N_noxref_10_M71_noxref_d \
 N_noxref_10_M73_noxref_d N_noxref_10_M75_noxref_d )  PM_TMRDFFQNX1\%noxref_10
x_PM_TMRDFFQNX1\%noxref_11 ( N_noxref_11_c_3765_p N_noxref_11_c_3758_n \
 N_noxref_11_c_3727_n N_noxref_11_c_3731_n N_noxref_11_c_3733_n \
 N_noxref_11_c_3711_n N_noxref_11_c_3804_p N_noxref_11_c_3712_n \
 N_noxref_11_c_3713_n N_noxref_11_c_3828_p N_noxref_11_M24_noxref_g \
 N_noxref_11_M93_noxref_g N_noxref_11_M94_noxref_g N_noxref_11_c_3714_n \
 N_noxref_11_c_3716_n N_noxref_11_c_3717_n N_noxref_11_c_3718_n \
 N_noxref_11_c_3719_n N_noxref_11_c_3720_n N_noxref_11_c_3721_n \
 N_noxref_11_c_3723_n N_noxref_11_c_3746_n N_noxref_11_M23_noxref_d \
 N_noxref_11_M89_noxref_d N_noxref_11_M91_noxref_d )  PM_TMRDFFQNX1\%noxref_11
x_PM_TMRDFFQNX1\%noxref_12 ( N_noxref_12_c_3882_n N_noxref_12_c_3884_n \
 N_noxref_12_c_3885_n N_noxref_12_c_3944_n N_noxref_12_c_3886_n \
 N_noxref_12_c_3888_n N_noxref_12_c_3862_n N_noxref_12_c_3946_n \
 N_noxref_12_c_3863_n N_noxref_12_c_3894_n N_noxref_12_c_3898_n \
 N_noxref_12_c_3900_n N_noxref_12_c_3865_n N_noxref_12_c_4059_p \
 N_noxref_12_c_3866_n N_noxref_12_c_4030_n N_noxref_12_c_3867_n \
 N_noxref_12_c_4121_p N_noxref_12_M13_noxref_g N_noxref_12_M19_noxref_g \
 N_noxref_12_M25_noxref_g N_noxref_12_M71_noxref_g N_noxref_12_M72_noxref_g \
 N_noxref_12_M83_noxref_g N_noxref_12_M84_noxref_g N_noxref_12_M95_noxref_g \
 N_noxref_12_M96_noxref_g N_noxref_12_c_3869_n N_noxref_12_c_3871_n \
 N_noxref_12_c_3872_n N_noxref_12_c_3873_n N_noxref_12_c_3874_n \
 N_noxref_12_c_3875_n N_noxref_12_c_3876_n N_noxref_12_c_3878_n \
 N_noxref_12_c_4024_n N_noxref_12_c_3922_n N_noxref_12_c_3955_n \
 N_noxref_12_c_3958_n N_noxref_12_c_3960_n N_noxref_12_c_3992_n \
 N_noxref_12_c_3994_n N_noxref_12_c_3995_n N_noxref_12_c_3963_n \
 N_noxref_12_c_3964_n N_noxref_12_c_4039_n N_noxref_12_c_4042_n \
 N_noxref_12_c_4044_n N_noxref_12_c_4083_p N_noxref_12_c_4162_p \
 N_noxref_12_c_4139_p N_noxref_12_c_4047_n N_noxref_12_c_4048_n \
 N_noxref_12_c_3965_n N_noxref_12_c_4001_n N_noxref_12_c_3967_n \
 N_noxref_12_c_4049_n N_noxref_12_c_4156_p N_noxref_12_c_4051_n \
 N_noxref_12_M21_noxref_d N_noxref_12_M85_noxref_d N_noxref_12_M87_noxref_d )  \
 PM_TMRDFFQNX1\%noxref_12
x_PM_TMRDFFQNX1\%D ( N_D_c_4217_n N_D_c_4236_n N_D_c_4238_n N_D_c_4251_n D D D \
 D N_D_c_4289_n N_D_c_4253_n N_D_c_4381_n N_D_c_4255_n N_D_c_4465_p \
 N_D_c_4257_n N_D_M4_noxref_g N_D_M17_noxref_g N_D_M30_noxref_g \
 N_D_M53_noxref_g N_D_M54_noxref_g N_D_M79_noxref_g N_D_M80_noxref_g \
 N_D_M105_noxref_g N_D_M106_noxref_g N_D_c_4299_n N_D_c_4300_n N_D_c_4301_n \
 N_D_c_4302_n N_D_c_4304_n N_D_c_4305_n N_D_c_4307_n N_D_c_4308_n N_D_c_4391_n \
 N_D_c_4392_n N_D_c_4393_n N_D_c_4394_n N_D_c_4396_n N_D_c_4397_n N_D_c_4399_n \
 N_D_c_4400_n N_D_c_4480_p N_D_c_4481_p N_D_c_4482_p N_D_c_4474_p N_D_c_4483_p \
 N_D_c_4469_p N_D_c_4485_p N_D_c_4470_p N_D_c_4310_n N_D_c_4311_n N_D_c_4313_n \
 N_D_c_4402_n N_D_c_4403_n N_D_c_4405_n N_D_c_4475_p N_D_c_4476_p N_D_c_4467_p \
 )  PM_TMRDFFQNX1\%D
x_PM_TMRDFFQNX1\%noxref_14 ( N_noxref_14_c_4694_n N_noxref_14_c_4696_n \
 N_noxref_14_c_4724_p N_noxref_14_c_4697_n N_noxref_14_c_4641_n \
 N_noxref_14_c_4659_n N_noxref_14_c_4663_n N_noxref_14_c_4665_n \
 N_noxref_14_c_4642_n N_noxref_14_c_4835_p N_noxref_14_c_4643_n \
 N_noxref_14_c_4644_n N_noxref_14_c_4713_n N_noxref_14_M28_noxref_g \
 N_noxref_14_M31_noxref_g N_noxref_14_M101_noxref_g N_noxref_14_M102_noxref_g \
 N_noxref_14_M107_noxref_g N_noxref_14_M108_noxref_g N_noxref_14_c_4749_p \
 N_noxref_14_c_4750_p N_noxref_14_c_4751_p N_noxref_14_c_4792_p \
 N_noxref_14_c_4770_p N_noxref_14_c_4794_p N_noxref_14_c_4771_p \
 N_noxref_14_c_4645_n N_noxref_14_c_4647_n N_noxref_14_c_4648_n \
 N_noxref_14_c_4649_n N_noxref_14_c_4650_n N_noxref_14_c_4651_n \
 N_noxref_14_c_4652_n N_noxref_14_c_4654_n N_noxref_14_c_4744_p \
 N_noxref_14_c_4754_p N_noxref_14_c_4739_p N_noxref_14_c_4682_n \
 N_noxref_14_M30_noxref_d N_noxref_14_M103_noxref_d N_noxref_14_M105_noxref_d ) \
 PM_TMRDFFQNX1\%noxref_14
x_PM_TMRDFFQNX1\%noxref_15 ( N_noxref_15_c_4936_p N_noxref_15_c_4921_n \
 N_noxref_15_c_4890_n N_noxref_15_c_4894_n N_noxref_15_c_4896_n \
 N_noxref_15_c_4874_n N_noxref_15_c_5000_p N_noxref_15_c_4875_n \
 N_noxref_15_c_4876_n N_noxref_15_c_4985_p N_noxref_15_M33_noxref_g \
 N_noxref_15_M111_noxref_g N_noxref_15_M112_noxref_g N_noxref_15_c_4877_n \
 N_noxref_15_c_4879_n N_noxref_15_c_4880_n N_noxref_15_c_4881_n \
 N_noxref_15_c_4882_n N_noxref_15_c_4883_n N_noxref_15_c_4884_n \
 N_noxref_15_c_4886_n N_noxref_15_c_4909_n N_noxref_15_M32_noxref_d \
 N_noxref_15_M107_noxref_d N_noxref_15_M109_noxref_d )  PM_TMRDFFQNX1\%noxref_15
x_PM_TMRDFFQNX1\%CLK ( N_CLK_c_5034_n N_CLK_c_5052_n N_CLK_c_5053_n \
 N_CLK_c_5060_n N_CLK_c_5061_n N_CLK_c_5079_n N_CLK_c_5092_n N_CLK_c_5111_n \
 N_CLK_c_5112_n N_CLK_c_5130_n CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK \
 CLK CLK CLK CLK CLK CLK CLK N_CLK_c_5025_n N_CLK_c_5203_n N_CLK_c_5026_n \
 N_CLK_c_5028_n N_CLK_c_5363_n N_CLK_c_5029_n N_CLK_c_5031_n N_CLK_c_5543_n \
 N_CLK_c_5032_n N_CLK_M1_noxref_g N_CLK_M8_noxref_g N_CLK_M14_noxref_g \
 N_CLK_M21_noxref_g N_CLK_M27_noxref_g N_CLK_M34_noxref_g N_CLK_M47_noxref_g \
 N_CLK_M48_noxref_g N_CLK_M61_noxref_g N_CLK_M62_noxref_g N_CLK_M73_noxref_g \
 N_CLK_M74_noxref_g N_CLK_M87_noxref_g N_CLK_M88_noxref_g N_CLK_M99_noxref_g \
 N_CLK_M100_noxref_g N_CLK_M113_noxref_g N_CLK_M114_noxref_g N_CLK_c_5300_n \
 N_CLK_c_5303_n N_CLK_c_5698_p N_CLK_c_5705_p N_CLK_c_5187_n N_CLK_c_5188_n \
 N_CLK_c_5189_n N_CLK_c_5190_n N_CLK_c_5193_n N_CLK_c_5212_n N_CLK_c_5215_n \
 N_CLK_c_5217_n N_CLK_c_5313_n N_CLK_c_5315_n N_CLK_c_5316_n N_CLK_c_5220_n \
 N_CLK_c_5221_n N_CLK_c_5461_n N_CLK_c_5464_n N_CLK_c_5727_p N_CLK_c_5734_p \
 N_CLK_c_5347_n N_CLK_c_5348_n N_CLK_c_5349_n N_CLK_c_5350_n N_CLK_c_5353_n \
 N_CLK_c_5372_n N_CLK_c_5375_n N_CLK_c_5377_n N_CLK_c_5474_n N_CLK_c_5476_n \
 N_CLK_c_5477_n N_CLK_c_5380_n N_CLK_c_5381_n N_CLK_c_5627_p N_CLK_c_5629_p \
 N_CLK_c_5756_p N_CLK_c_5763_p N_CLK_c_5529_n N_CLK_c_5530_n N_CLK_c_5531_n \
 N_CLK_c_5532_n N_CLK_c_5535_n N_CLK_c_5552_n N_CLK_c_5555_n N_CLK_c_5557_n \
 N_CLK_c_5596_p N_CLK_c_5647_p N_CLK_c_5614_p N_CLK_c_5560_n N_CLK_c_5561_n \
 N_CLK_c_5194_n N_CLK_c_5222_n N_CLK_c_5326_n N_CLK_c_5224_n N_CLK_c_5354_n \
 N_CLK_c_5382_n N_CLK_c_5486_n N_CLK_c_5384_n N_CLK_c_5536_n N_CLK_c_5562_n \
 N_CLK_c_5621_p N_CLK_c_5564_n )  PM_TMRDFFQNX1\%CLK
x_PM_TMRDFFQNX1\%noxref_17 ( N_noxref_17_c_5873_n N_noxref_17_c_5874_n \
 N_noxref_17_c_5847_n N_noxref_17_c_5848_n N_noxref_17_c_5801_n \
 N_noxref_17_c_5805_n N_noxref_17_c_5807_n N_noxref_17_c_5811_n \
 N_noxref_17_c_5777_n N_noxref_17_c_5990_p N_noxref_17_c_5815_n \
 N_noxref_17_c_5778_n N_noxref_17_c_5779_n N_noxref_17_c_5934_n \
 N_noxref_17_c_5898_n N_noxref_17_M29_noxref_g N_noxref_17_M35_noxref_g \
 N_noxref_17_M103_noxref_g N_noxref_17_M104_noxref_g N_noxref_17_M115_noxref_g \
 N_noxref_17_M116_noxref_g N_noxref_17_c_5780_n N_noxref_17_c_5782_n \
 N_noxref_17_c_5783_n N_noxref_17_c_5784_n N_noxref_17_c_5785_n \
 N_noxref_17_c_5786_n N_noxref_17_c_5787_n N_noxref_17_c_5789_n \
 N_noxref_17_c_5790_n N_noxref_17_c_5792_n N_noxref_17_c_5793_n \
 N_noxref_17_c_5794_n N_noxref_17_c_5795_n N_noxref_17_c_5796_n \
 N_noxref_17_c_5797_n N_noxref_17_c_5799_n N_noxref_17_c_5830_n \
 N_noxref_17_c_5831_n N_noxref_17_M28_noxref_d N_noxref_17_M97_noxref_d \
 N_noxref_17_M99_noxref_d N_noxref_17_M101_noxref_d )  PM_TMRDFFQNX1\%noxref_17
x_PM_TMRDFFQNX1\%noxref_18 ( N_noxref_18_c_6048_n N_noxref_18_c_6054_n \
 N_noxref_18_c_6057_n N_noxref_18_c_6061_n N_noxref_18_c_6063_n \
 N_noxref_18_c_6032_n N_noxref_18_c_6167_p N_noxref_18_c_6033_n \
 N_noxref_18_c_6034_n N_noxref_18_c_6153_p N_noxref_18_M37_noxref_g \
 N_noxref_18_M119_noxref_g N_noxref_18_M120_noxref_g N_noxref_18_c_6035_n \
 N_noxref_18_c_6037_n N_noxref_18_c_6038_n N_noxref_18_c_6039_n \
 N_noxref_18_c_6040_n N_noxref_18_c_6041_n N_noxref_18_c_6042_n \
 N_noxref_18_c_6044_n N_noxref_18_c_6076_n N_noxref_18_M36_noxref_d \
 N_noxref_18_M115_noxref_d N_noxref_18_M117_noxref_d )  PM_TMRDFFQNX1\%noxref_18
x_PM_TMRDFFQNX1\%noxref_19 ( N_noxref_19_c_6210_n N_noxref_19_c_6212_n \
 N_noxref_19_c_6213_n N_noxref_19_c_6284_n N_noxref_19_c_6215_n \
 N_noxref_19_c_6222_n N_noxref_19_c_6190_n N_noxref_19_c_6286_n \
 N_noxref_19_c_6191_n N_noxref_19_c_6230_n N_noxref_19_c_6234_n \
 N_noxref_19_c_6236_n N_noxref_19_c_6193_n N_noxref_19_c_6504_p \
 N_noxref_19_c_6194_n N_noxref_19_c_6440_n N_noxref_19_c_6195_n \
 N_noxref_19_c_6381_n N_noxref_19_M26_noxref_g N_noxref_19_M32_noxref_g \
 N_noxref_19_M38_noxref_g N_noxref_19_M97_noxref_g N_noxref_19_M98_noxref_g \
 N_noxref_19_M109_noxref_g N_noxref_19_M110_noxref_g N_noxref_19_M121_noxref_g \
 N_noxref_19_M122_noxref_g N_noxref_19_c_6197_n N_noxref_19_c_6199_n \
 N_noxref_19_c_6200_n N_noxref_19_c_6201_n N_noxref_19_c_6202_n \
 N_noxref_19_c_6203_n N_noxref_19_c_6204_n N_noxref_19_c_6206_n \
 N_noxref_19_c_6395_n N_noxref_19_c_6258_n N_noxref_19_c_6295_n \
 N_noxref_19_c_6298_n N_noxref_19_c_6300_n N_noxref_19_c_6332_n \
 N_noxref_19_c_6334_n N_noxref_19_c_6335_n N_noxref_19_c_6303_n \
 N_noxref_19_c_6304_n N_noxref_19_c_6449_n N_noxref_19_c_6452_n \
 N_noxref_19_c_6454_n N_noxref_19_c_6465_p N_noxref_19_c_6494_p \
 N_noxref_19_c_6478_p N_noxref_19_c_6457_n N_noxref_19_c_6458_n \
 N_noxref_19_c_6305_n N_noxref_19_c_6341_n N_noxref_19_c_6307_n \
 N_noxref_19_c_6459_n N_noxref_19_c_6485_p N_noxref_19_c_6461_n \
 N_noxref_19_M34_noxref_d N_noxref_19_M111_noxref_d N_noxref_19_M113_noxref_d ) \
 PM_TMRDFFQNX1\%noxref_19
x_PM_TMRDFFQNX1\%noxref_20 ( N_noxref_20_c_6592_n N_noxref_20_c_6653_n \
 N_noxref_20_c_6593_n N_noxref_20_c_6595_n N_noxref_20_c_6597_n \
 N_noxref_20_c_6602_n N_noxref_20_c_6655_n N_noxref_20_c_6560_n \
 N_noxref_20_c_6608_n N_noxref_20_c_6612_n N_noxref_20_c_6614_n \
 N_noxref_20_c_6562_n N_noxref_20_c_6762_p N_noxref_20_c_6563_n \
 N_noxref_20_c_6564_n N_noxref_20_c_6567_n N_noxref_20_c_6743_n \
 N_noxref_20_M36_noxref_g N_noxref_20_M39_noxref_g N_noxref_20_M41_noxref_g \
 N_noxref_20_M117_noxref_g N_noxref_20_M118_noxref_g N_noxref_20_M123_noxref_g \
 N_noxref_20_M124_noxref_g N_noxref_20_M127_noxref_g N_noxref_20_M128_noxref_g \
 N_noxref_20_c_6663_n N_noxref_20_c_6666_n N_noxref_20_c_6668_n \
 N_noxref_20_c_6703_n N_noxref_20_c_6705_n N_noxref_20_c_6706_n \
 N_noxref_20_c_6671_n N_noxref_20_c_6672_n N_noxref_20_c_6569_n \
 N_noxref_20_c_6571_n N_noxref_20_c_6572_n N_noxref_20_c_6573_n \
 N_noxref_20_c_6574_n N_noxref_20_c_6575_n N_noxref_20_c_6775_p \
 N_noxref_20_c_6639_n N_noxref_20_c_6576_n N_noxref_20_c_6578_n \
 N_noxref_20_c_6579_n N_noxref_20_c_6581_n N_noxref_20_c_6844_p \
 N_noxref_20_c_6582_n N_noxref_20_c_6583_n N_noxref_20_c_6584_n \
 N_noxref_20_c_6585_n N_noxref_20_c_6587_n N_noxref_20_c_6673_n \
 N_noxref_20_c_6712_n N_noxref_20_c_6675_n N_noxref_20_c_6588_n \
 N_noxref_20_c_6641_n N_noxref_20_M38_noxref_d N_noxref_20_M119_noxref_d \
 N_noxref_20_M121_noxref_d )  PM_TMRDFFQNX1\%noxref_20
x_PM_TMRDFFQNX1\%noxref_21 ( N_noxref_21_c_6904_n N_noxref_21_c_6909_n \
 N_noxref_21_c_6911_n N_noxref_21_c_6935_n N_noxref_21_c_6938_n \
 N_noxref_21_c_6956_n N_noxref_21_c_7001_n N_noxref_21_c_6939_n \
 N_noxref_21_c_6959_n N_noxref_21_c_6963_n N_noxref_21_c_6965_n \
 N_noxref_21_c_6941_n N_noxref_21_c_7334_p N_noxref_21_c_6942_n \
 N_noxref_21_c_6970_n N_noxref_21_c_6944_n N_noxref_21_c_6946_n \
 N_noxref_21_c_7080_n N_noxref_21_c_7243_p N_noxref_21_M23_noxref_g \
 N_noxref_21_M40_noxref_g N_noxref_21_M44_noxref_g N_noxref_21_M91_noxref_g \
 N_noxref_21_M92_noxref_g N_noxref_21_M125_noxref_g N_noxref_21_M126_noxref_g \
 N_noxref_21_M133_noxref_g N_noxref_21_M134_noxref_g N_noxref_21_c_7009_n \
 N_noxref_21_c_7012_n N_noxref_21_c_7014_n N_noxref_21_c_7046_n \
 N_noxref_21_c_7048_n N_noxref_21_c_7049_n N_noxref_21_c_7017_n \
 N_noxref_21_c_7018_n N_noxref_21_c_7186_n N_noxref_21_c_7189_n \
 N_noxref_21_c_7191_n N_noxref_21_c_6986_n N_noxref_21_c_7274_p \
 N_noxref_21_c_7275_p N_noxref_21_c_7195_n N_noxref_21_c_7196_n \
 N_noxref_21_c_7239_p N_noxref_21_c_7250_p N_noxref_21_c_7241_p \
 N_noxref_21_c_7291_p N_noxref_21_c_7282_p N_noxref_21_c_7252_p \
 N_noxref_21_c_7249_p N_noxref_21_c_7253_p N_noxref_21_c_7019_n \
 N_noxref_21_c_7055_n N_noxref_21_c_7021_n N_noxref_21_c_6948_n \
 N_noxref_21_c_7394_p N_noxref_21_c_6987_n N_noxref_21_c_7226_p \
 N_noxref_21_c_7293_p N_noxref_21_c_7233_p N_noxref_21_M25_noxref_d \
 N_noxref_21_M93_noxref_d N_noxref_21_M95_noxref_d )  PM_TMRDFFQNX1\%noxref_21
x_PM_TMRDFFQNX1\%noxref_22 ( N_noxref_22_c_7406_n N_noxref_22_c_7412_n \
 N_noxref_22_c_7417_n N_noxref_22_c_7421_n N_noxref_22_c_7423_n \
 N_noxref_22_c_7426_n N_noxref_22_c_7452_n N_noxref_22_c_7428_n \
 N_noxref_22_c_7471_p N_noxref_22_M123_noxref_d N_noxref_22_M125_noxref_d \
 N_noxref_22_M127_noxref_s N_noxref_22_M128_noxref_d N_noxref_22_M130_noxref_d \
 )  PM_TMRDFFQNX1\%noxref_22
x_PM_TMRDFFQNX1\%noxref_23 ( N_noxref_23_c_7497_n N_noxref_23_c_7578_n \
 N_noxref_23_c_7498_n N_noxref_23_c_7641_n N_noxref_23_c_7513_n \
 N_noxref_23_c_7514_n N_noxref_23_c_7579_n N_noxref_23_c_7515_n \
 N_noxref_23_c_7540_n N_noxref_23_c_7544_n N_noxref_23_c_7546_n \
 N_noxref_23_c_7517_n N_noxref_23_c_7713_n N_noxref_23_c_7518_n \
 N_noxref_23_c_7519_n N_noxref_23_c_7521_n N_noxref_23_c_7657_n \
 N_noxref_23_M10_noxref_g N_noxref_23_M42_noxref_g N_noxref_23_M43_noxref_g \
 N_noxref_23_M65_noxref_g N_noxref_23_M66_noxref_g N_noxref_23_M129_noxref_g \
 N_noxref_23_M130_noxref_g N_noxref_23_M131_noxref_g N_noxref_23_M132_noxref_g \
 N_noxref_23_c_7587_n N_noxref_23_c_7590_n N_noxref_23_c_7592_n \
 N_noxref_23_c_7624_n N_noxref_23_c_7626_n N_noxref_23_c_7627_n \
 N_noxref_23_c_7595_n N_noxref_23_c_7596_n N_noxref_23_c_7789_n \
 N_noxref_23_c_7792_n N_noxref_23_c_7863_p N_noxref_23_c_7794_n \
 N_noxref_23_c_7891_p N_noxref_23_c_7892_p N_noxref_23_c_7565_n \
 N_noxref_23_c_7798_n N_noxref_23_c_7799_n N_noxref_23_c_7800_n \
 N_noxref_23_c_7522_n N_noxref_23_c_7523_n N_noxref_23_c_7525_n \
 N_noxref_23_c_7828_n N_noxref_23_c_7526_n N_noxref_23_c_7527_n \
 N_noxref_23_c_7528_n N_noxref_23_c_7830_n N_noxref_23_c_7566_n \
 N_noxref_23_c_7529_n N_noxref_23_c_7531_n N_noxref_23_c_7597_n \
 N_noxref_23_c_7633_n N_noxref_23_c_7599_n N_noxref_23_c_7532_n \
 N_noxref_23_M12_noxref_d N_noxref_23_M67_noxref_d N_noxref_23_M69_noxref_d )  \
 PM_TMRDFFQNX1\%noxref_23
x_PM_TMRDFFQNX1\%noxref_24 ( N_noxref_24_c_7956_n N_noxref_24_c_7960_n \
 N_noxref_24_c_7971_n N_noxref_24_c_7962_n N_noxref_24_c_7963_n \
 N_noxref_24_c_7964_n N_noxref_24_c_7983_n N_noxref_24_c_7966_n \
 N_noxref_24_c_7984_n N_noxref_24_M127_noxref_d N_noxref_24_M129_noxref_d \
 N_noxref_24_M131_noxref_s N_noxref_24_M132_noxref_d N_noxref_24_M134_noxref_d \
 )  PM_TMRDFFQNX1\%noxref_24
x_PM_TMRDFFQNX1\%QN ( N_QN_c_8045_n N_QN_c_8052_n N_QN_c_8053_n N_QN_c_8059_n \
 QN QN QN QN QN QN QN QN N_QN_c_8112_n N_QN_c_8074_n N_QN_c_8075_n \
 N_QN_c_8061_n N_QN_c_8119_n N_QN_c_8120_n N_QN_M40_noxref_d N_QN_M42_noxref_d \
 N_QN_M44_noxref_d N_QN_M131_noxref_d N_QN_M133_noxref_d )  PM_TMRDFFQNX1\%QN
x_PM_TMRDFFQNX1\%noxref_26 ( N_noxref_26_c_8231_n N_noxref_26_c_8214_n \
 N_noxref_26_c_8218_n N_noxref_26_c_8221_n N_noxref_26_c_8239_n \
 N_noxref_26_M0_noxref_s )  PM_TMRDFFQNX1\%noxref_26
x_PM_TMRDFFQNX1\%noxref_27 ( N_noxref_27_c_8261_n N_noxref_27_c_8263_n \
 N_noxref_27_c_8266_n N_noxref_27_c_8269_n N_noxref_27_c_8280_n \
 N_noxref_27_M1_noxref_d N_noxref_27_M2_noxref_s )  PM_TMRDFFQNX1\%noxref_27
x_PM_TMRDFFQNX1\%noxref_28 ( N_noxref_28_c_8333_n N_noxref_28_c_8314_n \
 N_noxref_28_c_8318_n N_noxref_28_c_8321_n N_noxref_28_c_8322_n \
 N_noxref_28_c_8325_n N_noxref_28_M3_noxref_s )  PM_TMRDFFQNX1\%noxref_28
x_PM_TMRDFFQNX1\%noxref_29 ( N_noxref_29_c_8387_n N_noxref_29_c_8368_n \
 N_noxref_29_c_8372_n N_noxref_29_c_8375_n N_noxref_29_c_8376_n \
 N_noxref_29_c_8379_n N_noxref_29_M5_noxref_s )  PM_TMRDFFQNX1\%noxref_29
x_PM_TMRDFFQNX1\%noxref_30 ( N_noxref_30_c_8439_n N_noxref_30_c_8420_n \
 N_noxref_30_c_8424_n N_noxref_30_c_8427_n N_noxref_30_c_8428_n \
 N_noxref_30_c_8431_n N_noxref_30_M7_noxref_s )  PM_TMRDFFQNX1\%noxref_30
x_PM_TMRDFFQNX1\%noxref_31 ( N_noxref_31_c_8491_n N_noxref_31_c_8472_n \
 N_noxref_31_c_8476_n N_noxref_31_c_8479_n N_noxref_31_c_8480_n \
 N_noxref_31_c_8483_n N_noxref_31_M9_noxref_s )  PM_TMRDFFQNX1\%noxref_31
x_PM_TMRDFFQNX1\%noxref_32 ( N_noxref_32_c_8543_n N_noxref_32_c_8524_n \
 N_noxref_32_c_8528_n N_noxref_32_c_8531_n N_noxref_32_c_8532_n \
 N_noxref_32_c_8535_n N_noxref_32_M11_noxref_s )  PM_TMRDFFQNX1\%noxref_32
x_PM_TMRDFFQNX1\%noxref_33 ( N_noxref_33_c_8593_n N_noxref_33_c_8576_n \
 N_noxref_33_c_8580_n N_noxref_33_c_8583_n N_noxref_33_c_8605_n \
 N_noxref_33_M13_noxref_s )  PM_TMRDFFQNX1\%noxref_33
x_PM_TMRDFFQNX1\%noxref_34 ( N_noxref_34_c_8626_n N_noxref_34_c_8628_n \
 N_noxref_34_c_8631_n N_noxref_34_c_8634_n N_noxref_34_c_8644_n \
 N_noxref_34_M14_noxref_d N_noxref_34_M15_noxref_s )  PM_TMRDFFQNX1\%noxref_34
x_PM_TMRDFFQNX1\%noxref_35 ( N_noxref_35_c_8698_n N_noxref_35_c_8679_n \
 N_noxref_35_c_8683_n N_noxref_35_c_8686_n N_noxref_35_c_8687_n \
 N_noxref_35_c_8690_n N_noxref_35_M16_noxref_s )  PM_TMRDFFQNX1\%noxref_35
x_PM_TMRDFFQNX1\%noxref_36 ( N_noxref_36_c_8752_n N_noxref_36_c_8733_n \
 N_noxref_36_c_8737_n N_noxref_36_c_8740_n N_noxref_36_c_8741_n \
 N_noxref_36_c_8744_n N_noxref_36_M18_noxref_s )  PM_TMRDFFQNX1\%noxref_36
x_PM_TMRDFFQNX1\%noxref_37 ( N_noxref_37_c_8804_n N_noxref_37_c_8785_n \
 N_noxref_37_c_8789_n N_noxref_37_c_8792_n N_noxref_37_c_8793_n \
 N_noxref_37_c_8796_n N_noxref_37_M20_noxref_s )  PM_TMRDFFQNX1\%noxref_37
x_PM_TMRDFFQNX1\%noxref_38 ( N_noxref_38_c_8856_n N_noxref_38_c_8837_n \
 N_noxref_38_c_8841_n N_noxref_38_c_8844_n N_noxref_38_c_8845_n \
 N_noxref_38_c_8848_n N_noxref_38_M22_noxref_s )  PM_TMRDFFQNX1\%noxref_38
x_PM_TMRDFFQNX1\%noxref_39 ( N_noxref_39_c_8910_n N_noxref_39_c_8891_n \
 N_noxref_39_c_8895_n N_noxref_39_c_8898_n N_noxref_39_c_8899_n \
 N_noxref_39_c_8902_n N_noxref_39_M24_noxref_s )  PM_TMRDFFQNX1\%noxref_39
x_PM_TMRDFFQNX1\%noxref_40 ( N_noxref_40_c_8970_n N_noxref_40_c_8945_n \
 N_noxref_40_c_8949_n N_noxref_40_c_8952_n N_noxref_40_c_8963_n \
 N_noxref_40_M26_noxref_s )  PM_TMRDFFQNX1\%noxref_40
x_PM_TMRDFFQNX1\%noxref_41 ( N_noxref_41_c_8995_n N_noxref_41_c_8997_n \
 N_noxref_41_c_9000_n N_noxref_41_c_9003_n N_noxref_41_c_9013_n \
 N_noxref_41_M27_noxref_d N_noxref_41_M28_noxref_s )  PM_TMRDFFQNX1\%noxref_41
x_PM_TMRDFFQNX1\%noxref_42 ( N_noxref_42_c_9076_n N_noxref_42_c_9048_n \
 N_noxref_42_c_9052_n N_noxref_42_c_9055_n N_noxref_42_c_9056_n \
 N_noxref_42_c_9059_n N_noxref_42_M29_noxref_s )  PM_TMRDFFQNX1\%noxref_42
x_PM_TMRDFFQNX1\%noxref_43 ( N_noxref_43_c_9119_n N_noxref_43_c_9100_n \
 N_noxref_43_c_9104_n N_noxref_43_c_9107_n N_noxref_43_c_9108_n \
 N_noxref_43_c_9111_n N_noxref_43_M31_noxref_s )  PM_TMRDFFQNX1\%noxref_43
x_PM_TMRDFFQNX1\%noxref_44 ( N_noxref_44_c_9171_n N_noxref_44_c_9152_n \
 N_noxref_44_c_9156_n N_noxref_44_c_9159_n N_noxref_44_c_9160_n \
 N_noxref_44_c_9163_n N_noxref_44_M33_noxref_s )  PM_TMRDFFQNX1\%noxref_44
x_PM_TMRDFFQNX1\%noxref_45 ( N_noxref_45_c_9223_n N_noxref_45_c_9204_n \
 N_noxref_45_c_9208_n N_noxref_45_c_9211_n N_noxref_45_c_9212_n \
 N_noxref_45_c_9215_n N_noxref_45_M35_noxref_s )  PM_TMRDFFQNX1\%noxref_45
x_PM_TMRDFFQNX1\%noxref_46 ( N_noxref_46_c_9275_n N_noxref_46_c_9256_n \
 N_noxref_46_c_9260_n N_noxref_46_c_9263_n N_noxref_46_c_9264_n \
 N_noxref_46_c_9267_n N_noxref_46_M37_noxref_s )  PM_TMRDFFQNX1\%noxref_46
x_PM_TMRDFFQNX1\%noxref_47 ( N_noxref_47_c_9327_n N_noxref_47_c_9308_n \
 N_noxref_47_c_9312_n N_noxref_47_c_9315_n N_noxref_47_c_9316_n \
 N_noxref_47_c_9319_n N_noxref_47_M39_noxref_s )  PM_TMRDFFQNX1\%noxref_47
x_PM_TMRDFFQNX1\%noxref_48 ( N_noxref_48_c_9384_n N_noxref_48_c_9366_n \
 N_noxref_48_c_9369_n N_noxref_48_c_9372_n N_noxref_48_c_9373_n \
 N_noxref_48_c_9376_n N_noxref_48_M41_noxref_s )  PM_TMRDFFQNX1\%noxref_48
x_PM_TMRDFFQNX1\%noxref_49 ( N_noxref_49_c_9449_n N_noxref_49_c_9422_n \
 N_noxref_49_c_9425_n N_noxref_49_c_9428_n N_noxref_49_c_9429_n \
 N_noxref_49_c_9431_n N_noxref_49_M43_noxref_s )  PM_TMRDFFQNX1\%noxref_49
cc_1 ( N_GND_c_1_p N_VDD_c_937_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_938_n ) capacitor c=0.00989031f //x=73.63 //y=0 \
 //x2=73.63 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_939_n ) capacitor c=0.00500587f //x=4.81 //y=0 \
 //x2=4.81 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_940_n ) capacitor c=0.0057235f //x=8.14 //y=0 \
 //x2=8.14 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_941_n ) capacitor c=0.0057235f //x=11.47 //y=0 \
 //x2=11.47 //y2=7.4
cc_6 ( N_GND_c_6_p N_VDD_c_942_n ) capacitor c=0.0057235f //x=14.8 //y=0 \
 //x2=14.8 //y2=7.4
cc_7 ( N_GND_c_7_p N_VDD_c_943_n ) capacitor c=0.0057235f //x=18.13 //y=0 \
 //x2=18.13 //y2=7.4
cc_8 ( N_GND_c_8_p N_VDD_c_944_n ) capacitor c=0.00989031f //x=21.46 //y=0 \
 //x2=21.46 //y2=7.4
cc_9 ( N_GND_c_9_p N_VDD_c_945_n ) capacitor c=0.0057235f //x=26.27 //y=0 \
 //x2=26.27 //y2=7.4
cc_10 ( N_GND_c_10_p N_VDD_c_946_n ) capacitor c=0.0057235f //x=29.6 //y=0 \
 //x2=29.6 //y2=7.4
cc_11 ( N_GND_c_11_p N_VDD_c_947_n ) capacitor c=0.0057235f //x=32.93 //y=0 \
 //x2=32.93 //y2=7.4
cc_12 ( N_GND_c_12_p N_VDD_c_948_n ) capacitor c=0.0057235f //x=36.26 //y=0 \
 //x2=36.26 //y2=7.4
cc_13 ( N_GND_c_13_p N_VDD_c_949_n ) capacitor c=0.0057235f //x=39.59 //y=0 \
 //x2=39.59 //y2=7.4
cc_14 ( N_GND_c_14_p N_VDD_c_950_n ) capacitor c=0.00989031f //x=42.92 //y=0 \
 //x2=42.92 //y2=7.4
cc_15 ( N_GND_c_15_p N_VDD_c_951_n ) capacitor c=0.0057235f //x=47.73 //y=0 \
 //x2=47.73 //y2=7.4
cc_16 ( N_GND_c_16_p N_VDD_c_952_n ) capacitor c=0.00474727f //x=51.06 //y=0 \
 //x2=51.06 //y2=7.4
cc_17 ( N_GND_c_17_p N_VDD_c_953_n ) capacitor c=0.00474727f //x=54.39 //y=0 \
 //x2=54.39 //y2=7.4
cc_18 ( N_GND_c_18_p N_VDD_c_954_n ) capacitor c=0.00474727f //x=57.72 //y=0 \
 //x2=57.72 //y2=7.4
cc_19 ( N_GND_c_19_p N_VDD_c_955_n ) capacitor c=0.00474727f //x=61.05 //y=0 \
 //x2=61.05 //y2=7.4
cc_20 ( N_GND_c_20_p N_VDD_c_956_n ) capacitor c=0.00802221f //x=64.38 //y=0 \
 //x2=64.38 //y2=7.4
cc_21 ( N_GND_c_21_p N_VDD_c_957_n ) capacitor c=0.00482014f //x=67.71 //y=0 \
 //x2=67.71 //y2=7.4
cc_22 ( N_GND_c_22_p N_VDD_c_958_n ) capacitor c=0.00553669f //x=71.04 //y=0 \
 //x2=71.04 //y2=7.4
cc_23 ( N_GND_c_23_p N_noxref_3_c_1935_n ) capacitor c=0.0232424f //x=73.63 \
 //y=0 //x2=7.285 //y2=3.33
cc_24 ( N_GND_c_24_p N_noxref_3_c_1935_n ) capacitor c=0.00174514f //x=4.64 \
 //y=0 //x2=7.285 //y2=3.33
cc_25 ( N_GND_c_25_p N_noxref_3_c_1935_n ) capacitor c=0.00192599f //x=5.905 \
 //y=0 //x2=7.285 //y2=3.33
cc_26 ( N_GND_c_3_p N_noxref_3_c_1935_n ) capacitor c=0.00820844f //x=4.81 \
 //y=0 //x2=7.285 //y2=3.33
cc_27 ( N_GND_c_23_p N_noxref_3_c_1939_n ) capacitor c=0.00172266f //x=73.63 \
 //y=0 //x2=3.445 //y2=3.33
cc_28 ( N_GND_c_4_p N_noxref_3_c_1940_n ) capacitor c=0.00505527f //x=8.14 \
 //y=0 //x2=9.135 //y2=3.33
cc_29 ( N_GND_c_3_p N_noxref_3_c_1941_n ) capacitor c=0.00123372f //x=4.81 \
 //y=0 //x2=3.33 //y2=2.08
cc_30 ( N_GND_c_4_p N_noxref_3_c_1942_n ) capacitor c=0.0435122f //x=8.14 \
 //y=0 //x2=7.315 //y2=1.655
cc_31 ( N_GND_c_3_p N_noxref_3_c_1943_n ) capacitor c=9.64732e-19 //x=4.81 \
 //y=0 //x2=7.4 //y2=3.33
cc_32 ( N_GND_c_4_p N_noxref_3_c_1944_n ) capacitor c=0.0152765f //x=8.14 \
 //y=0 //x2=9.25 //y2=2.08
cc_33 ( N_GND_c_33_p N_noxref_3_c_1945_n ) capacitor c=0.00135046f //x=9.235 \
 //y=0 //x2=9.055 //y2=0.865
cc_34 ( N_GND_M5_noxref_d N_noxref_3_c_1945_n ) capacitor c=0.00220047f \
 //x=9.13 //y=0.865 //x2=9.055 //y2=0.865
cc_35 ( N_GND_M5_noxref_d N_noxref_3_c_1947_n ) capacitor c=0.00255985f \
 //x=9.13 //y=0.865 //x2=9.055 //y2=1.21
cc_36 ( N_GND_c_4_p N_noxref_3_c_1948_n ) capacitor c=0.0018059f //x=8.14 \
 //y=0 //x2=9.055 //y2=1.52
cc_37 ( N_GND_c_4_p N_noxref_3_c_1949_n ) capacitor c=0.0114883f //x=8.14 \
 //y=0 //x2=9.055 //y2=1.915
cc_38 ( N_GND_M5_noxref_d N_noxref_3_c_1950_n ) capacitor c=0.0131326f \
 //x=9.13 //y=0.865 //x2=9.43 //y2=0.71
cc_39 ( N_GND_M5_noxref_d N_noxref_3_c_1951_n ) capacitor c=0.00193127f \
 //x=9.13 //y=0.865 //x2=9.43 //y2=1.365
cc_40 ( N_GND_c_40_p N_noxref_3_c_1952_n ) capacitor c=0.00130622f //x=11.3 \
 //y=0 //x2=9.585 //y2=0.865
cc_41 ( N_GND_M5_noxref_d N_noxref_3_c_1952_n ) capacitor c=0.00257848f \
 //x=9.13 //y=0.865 //x2=9.585 //y2=0.865
cc_42 ( N_GND_M5_noxref_d N_noxref_3_c_1954_n ) capacitor c=0.00255985f \
 //x=9.13 //y=0.865 //x2=9.585 //y2=1.21
cc_43 ( N_GND_c_3_p N_noxref_3_M4_noxref_d ) capacitor c=8.58106e-19 //x=4.81 \
 //y=0 //x2=6.77 //y2=0.905
cc_44 ( N_GND_c_4_p N_noxref_3_M4_noxref_d ) capacitor c=0.00616547f //x=8.14 \
 //y=0 //x2=6.77 //y2=0.905
cc_45 ( N_GND_M3_noxref_d N_noxref_3_M4_noxref_d ) capacitor c=0.00143464f \
 //x=5.8 //y=0.865 //x2=6.77 //y2=0.905
cc_46 ( N_GND_c_5_p N_noxref_4_c_2167_n ) capacitor c=0.00505527f //x=11.47 \
 //y=0 //x2=12.465 //y2=3.33
cc_47 ( N_GND_c_5_p N_noxref_4_c_2168_n ) capacitor c=0.0436694f //x=11.47 \
 //y=0 //x2=10.645 //y2=1.655
cc_48 ( N_GND_c_4_p N_noxref_4_c_2169_n ) capacitor c=9.64732e-19 //x=8.14 \
 //y=0 //x2=10.73 //y2=3.33
cc_49 ( N_GND_c_5_p N_noxref_4_c_2170_n ) capacitor c=0.0153491f //x=11.47 \
 //y=0 //x2=12.58 //y2=2.08
cc_50 ( N_GND_c_50_p N_noxref_4_c_2171_n ) capacitor c=0.00135046f //x=12.565 \
 //y=0 //x2=12.385 //y2=0.865
cc_51 ( N_GND_M7_noxref_d N_noxref_4_c_2171_n ) capacitor c=0.00220047f \
 //x=12.46 //y=0.865 //x2=12.385 //y2=0.865
cc_52 ( N_GND_M7_noxref_d N_noxref_4_c_2173_n ) capacitor c=0.00255985f \
 //x=12.46 //y=0.865 //x2=12.385 //y2=1.21
cc_53 ( N_GND_c_5_p N_noxref_4_c_2174_n ) capacitor c=0.0018059f //x=11.47 \
 //y=0 //x2=12.385 //y2=1.52
cc_54 ( N_GND_c_5_p N_noxref_4_c_2175_n ) capacitor c=0.0114883f //x=11.47 \
 //y=0 //x2=12.385 //y2=1.915
cc_55 ( N_GND_M7_noxref_d N_noxref_4_c_2176_n ) capacitor c=0.0131326f \
 //x=12.46 //y=0.865 //x2=12.76 //y2=0.71
cc_56 ( N_GND_M7_noxref_d N_noxref_4_c_2177_n ) capacitor c=0.00193127f \
 //x=12.46 //y=0.865 //x2=12.76 //y2=1.365
cc_57 ( N_GND_c_57_p N_noxref_4_c_2178_n ) capacitor c=0.00130622f //x=14.63 \
 //y=0 //x2=12.915 //y2=0.865
cc_58 ( N_GND_M7_noxref_d N_noxref_4_c_2178_n ) capacitor c=0.00257848f \
 //x=12.46 //y=0.865 //x2=12.915 //y2=0.865
cc_59 ( N_GND_M7_noxref_d N_noxref_4_c_2180_n ) capacitor c=0.00255985f \
 //x=12.46 //y=0.865 //x2=12.915 //y2=1.21
cc_60 ( N_GND_c_4_p N_noxref_4_M6_noxref_d ) capacitor c=8.58106e-19 //x=8.14 \
 //y=0 //x2=10.1 //y2=0.905
cc_61 ( N_GND_c_5_p N_noxref_4_M6_noxref_d ) capacitor c=0.00616547f //x=11.47 \
 //y=0 //x2=10.1 //y2=0.905
cc_62 ( N_GND_M5_noxref_d N_noxref_4_M6_noxref_d ) capacitor c=0.00143464f \
 //x=9.13 //y=0.865 //x2=10.1 //y2=0.905
cc_63 ( N_GND_c_6_p N_noxref_5_c_2317_n ) capacitor c=0.0034979f //x=14.8 \
 //y=0 //x2=15.795 //y2=3.7
cc_64 ( N_GND_c_3_p N_noxref_5_c_2318_n ) capacitor c=0.0456054f //x=4.81 \
 //y=0 //x2=3.985 //y2=1.665
cc_65 ( N_GND_c_3_p N_noxref_5_c_2319_n ) capacitor c=0.0175874f //x=4.81 \
 //y=0 //x2=5.92 //y2=2.08
cc_66 ( N_GND_c_6_p N_noxref_5_c_2320_n ) capacitor c=0.0153491f //x=14.8 \
 //y=0 //x2=15.91 //y2=2.08
cc_67 ( N_GND_c_25_p N_noxref_5_c_2321_n ) capacitor c=0.00135046f //x=5.905 \
 //y=0 //x2=5.725 //y2=0.865
cc_68 ( N_GND_M3_noxref_d N_noxref_5_c_2321_n ) capacitor c=0.00220047f \
 //x=5.8 //y=0.865 //x2=5.725 //y2=0.865
cc_69 ( N_GND_M3_noxref_d N_noxref_5_c_2323_n ) capacitor c=0.00255985f \
 //x=5.8 //y=0.865 //x2=5.725 //y2=1.21
cc_70 ( N_GND_c_3_p N_noxref_5_c_2324_n ) capacitor c=0.00189421f //x=4.81 \
 //y=0 //x2=5.725 //y2=1.52
cc_71 ( N_GND_c_3_p N_noxref_5_c_2325_n ) capacitor c=0.0114883f //x=4.81 \
 //y=0 //x2=5.725 //y2=1.915
cc_72 ( N_GND_M3_noxref_d N_noxref_5_c_2326_n ) capacitor c=0.0131326f //x=5.8 \
 //y=0.865 //x2=6.1 //y2=0.71
cc_73 ( N_GND_M3_noxref_d N_noxref_5_c_2327_n ) capacitor c=0.00193127f \
 //x=5.8 //y=0.865 //x2=6.1 //y2=1.365
cc_74 ( N_GND_c_74_p N_noxref_5_c_2328_n ) capacitor c=0.00130622f //x=7.97 \
 //y=0 //x2=6.255 //y2=0.865
cc_75 ( N_GND_M3_noxref_d N_noxref_5_c_2328_n ) capacitor c=0.00257848f \
 //x=5.8 //y=0.865 //x2=6.255 //y2=0.865
cc_76 ( N_GND_M3_noxref_d N_noxref_5_c_2330_n ) capacitor c=0.00255985f \
 //x=5.8 //y=0.865 //x2=6.255 //y2=1.21
cc_77 ( N_GND_c_77_p N_noxref_5_c_2331_n ) capacitor c=0.00135046f //x=15.895 \
 //y=0 //x2=15.715 //y2=0.865
cc_78 ( N_GND_M9_noxref_d N_noxref_5_c_2331_n ) capacitor c=0.00220047f \
 //x=15.79 //y=0.865 //x2=15.715 //y2=0.865
cc_79 ( N_GND_M9_noxref_d N_noxref_5_c_2333_n ) capacitor c=0.00255985f \
 //x=15.79 //y=0.865 //x2=15.715 //y2=1.21
cc_80 ( N_GND_c_6_p N_noxref_5_c_2334_n ) capacitor c=0.0018059f //x=14.8 \
 //y=0 //x2=15.715 //y2=1.52
cc_81 ( N_GND_c_6_p N_noxref_5_c_2335_n ) capacitor c=0.0114883f //x=14.8 \
 //y=0 //x2=15.715 //y2=1.915
cc_82 ( N_GND_M9_noxref_d N_noxref_5_c_2336_n ) capacitor c=0.0131326f \
 //x=15.79 //y=0.865 //x2=16.09 //y2=0.71
cc_83 ( N_GND_M9_noxref_d N_noxref_5_c_2337_n ) capacitor c=0.00193127f \
 //x=15.79 //y=0.865 //x2=16.09 //y2=1.365
cc_84 ( N_GND_c_84_p N_noxref_5_c_2338_n ) capacitor c=0.00130622f //x=17.96 \
 //y=0 //x2=16.245 //y2=0.865
cc_85 ( N_GND_M9_noxref_d N_noxref_5_c_2338_n ) capacitor c=0.00257848f \
 //x=15.79 //y=0.865 //x2=16.245 //y2=0.865
cc_86 ( N_GND_M9_noxref_d N_noxref_5_c_2340_n ) capacitor c=0.00255985f \
 //x=15.79 //y=0.865 //x2=16.245 //y2=1.21
cc_87 ( N_GND_c_3_p N_noxref_5_M2_noxref_d ) capacitor c=0.00591582f //x=4.81 \
 //y=0 //x2=3.395 //y2=0.915
cc_88 ( N_GND_c_7_p N_noxref_6_c_2565_n ) capacitor c=0.0436694f //x=18.13 \
 //y=0 //x2=17.305 //y2=1.655
cc_89 ( N_GND_c_6_p N_noxref_6_c_2566_n ) capacitor c=9.64732e-19 //x=14.8 \
 //y=0 //x2=17.39 //y2=3.7
cc_90 ( N_GND_c_7_p N_noxref_6_c_2567_n ) capacitor c=0.0153491f //x=18.13 \
 //y=0 //x2=19.24 //y2=2.08
cc_91 ( N_GND_c_91_p N_noxref_6_c_2568_n ) capacitor c=0.00135046f //x=19.225 \
 //y=0 //x2=19.045 //y2=0.865
cc_92 ( N_GND_M11_noxref_d N_noxref_6_c_2568_n ) capacitor c=0.00220047f \
 //x=19.12 //y=0.865 //x2=19.045 //y2=0.865
cc_93 ( N_GND_M11_noxref_d N_noxref_6_c_2570_n ) capacitor c=0.00255985f \
 //x=19.12 //y=0.865 //x2=19.045 //y2=1.21
cc_94 ( N_GND_c_7_p N_noxref_6_c_2571_n ) capacitor c=0.0018059f //x=18.13 \
 //y=0 //x2=19.045 //y2=1.52
cc_95 ( N_GND_c_7_p N_noxref_6_c_2572_n ) capacitor c=0.0114883f //x=18.13 \
 //y=0 //x2=19.045 //y2=1.915
cc_96 ( N_GND_M11_noxref_d N_noxref_6_c_2573_n ) capacitor c=0.0131326f \
 //x=19.12 //y=0.865 //x2=19.42 //y2=0.71
cc_97 ( N_GND_M11_noxref_d N_noxref_6_c_2574_n ) capacitor c=0.00193127f \
 //x=19.12 //y=0.865 //x2=19.42 //y2=1.365
cc_98 ( N_GND_c_98_p N_noxref_6_c_2575_n ) capacitor c=0.00130622f //x=21.29 \
 //y=0 //x2=19.575 //y2=0.865
cc_99 ( N_GND_M11_noxref_d N_noxref_6_c_2575_n ) capacitor c=0.00257848f \
 //x=19.12 //y=0.865 //x2=19.575 //y2=0.865
cc_100 ( N_GND_M11_noxref_d N_noxref_6_c_2577_n ) capacitor c=0.00255985f \
 //x=19.12 //y=0.865 //x2=19.575 //y2=1.21
cc_101 ( N_GND_c_6_p N_noxref_6_M10_noxref_d ) capacitor c=8.58106e-19 \
 //x=14.8 //y=0 //x2=16.76 //y2=0.905
cc_102 ( N_GND_c_7_p N_noxref_6_M10_noxref_d ) capacitor c=0.00616547f \
 //x=18.13 //y=0 //x2=16.76 //y2=0.905
cc_103 ( N_GND_M9_noxref_d N_noxref_6_M10_noxref_d ) capacitor c=0.00143464f \
 //x=15.79 //y=0.865 //x2=16.76 //y2=0.905
cc_104 ( N_GND_c_23_p N_noxref_7_c_2715_n ) capacitor c=0.0122686f //x=73.63 \
 //y=0 //x2=9.875 //y2=4.07
cc_105 ( N_GND_c_23_p N_noxref_7_c_2716_n ) capacitor c=0.0015877f //x=73.63 \
 //y=0 //x2=1.225 //y2=4.07
cc_106 ( N_GND_c_1_p N_noxref_7_c_2717_n ) capacitor c=0.0180363f //x=0.74 \
 //y=0 //x2=1.11 //y2=2.08
cc_107 ( N_GND_c_4_p N_noxref_7_c_2718_n ) capacitor c=8.24484e-19 //x=8.14 \
 //y=0 //x2=9.99 //y2=2.08
cc_108 ( N_GND_c_5_p N_noxref_7_c_2718_n ) capacitor c=7.09207e-19 //x=11.47 \
 //y=0 //x2=9.99 //y2=2.08
cc_109 ( N_GND_c_6_p N_noxref_7_c_2720_n ) capacitor c=0.0436694f //x=14.8 \
 //y=0 //x2=13.975 //y2=1.655
cc_110 ( N_GND_c_5_p N_noxref_7_c_2721_n ) capacitor c=9.64732e-19 //x=11.47 \
 //y=0 //x2=14.06 //y2=4.07
cc_111 ( N_GND_c_7_p N_noxref_7_c_2722_n ) capacitor c=7.51486e-19 //x=18.13 \
 //y=0 //x2=19.98 //y2=2.08
cc_112 ( N_GND_c_8_p N_noxref_7_c_2722_n ) capacitor c=7.09207e-19 //x=21.46 \
 //y=0 //x2=19.98 //y2=2.08
cc_113 ( N_GND_c_113_p N_noxref_7_c_2724_n ) capacitor c=0.00132755f //x=0.99 \
 //y=0 //x2=0.81 //y2=0.875
cc_114 ( N_GND_M0_noxref_d N_noxref_7_c_2724_n ) capacitor c=0.00211996f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=0.875
cc_115 ( N_GND_M0_noxref_d N_noxref_7_c_2726_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=1.22
cc_116 ( N_GND_c_1_p N_noxref_7_c_2727_n ) capacitor c=0.00295461f //x=0.74 \
 //y=0 //x2=0.81 //y2=1.53
cc_117 ( N_GND_c_1_p N_noxref_7_c_2728_n ) capacitor c=0.0134214f //x=0.74 \
 //y=0 //x2=0.81 //y2=1.915
cc_118 ( N_GND_M0_noxref_d N_noxref_7_c_2729_n ) capacitor c=0.0131341f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=0.72
cc_119 ( N_GND_M0_noxref_d N_noxref_7_c_2730_n ) capacitor c=0.00193146f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=1.375
cc_120 ( N_GND_c_24_p N_noxref_7_c_2731_n ) capacitor c=0.00129018f //x=4.64 \
 //y=0 //x2=1.34 //y2=0.875
cc_121 ( N_GND_M0_noxref_d N_noxref_7_c_2731_n ) capacitor c=0.00257848f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=0.875
cc_122 ( N_GND_M0_noxref_d N_noxref_7_c_2733_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=1.22
cc_123 ( N_GND_c_5_p N_noxref_7_M8_noxref_d ) capacitor c=8.58106e-19 \
 //x=11.47 //y=0 //x2=13.43 //y2=0.905
cc_124 ( N_GND_c_6_p N_noxref_7_M8_noxref_d ) capacitor c=0.00616547f //x=14.8 \
 //y=0 //x2=13.43 //y2=0.905
cc_125 ( N_GND_M7_noxref_d N_noxref_7_M8_noxref_d ) capacitor c=0.00143464f \
 //x=12.46 //y=0.865 //x2=13.43 //y2=0.905
cc_126 ( N_GND_c_9_p N_noxref_8_c_3068_n ) capacitor c=7.82389e-19 //x=26.27 \
 //y=0 //x2=24.79 //y2=2.08
cc_127 ( N_GND_c_10_p N_noxref_8_c_3069_n ) capacitor c=0.0435122f //x=29.6 \
 //y=0 //x2=28.775 //y2=1.655
cc_128 ( N_GND_c_9_p N_noxref_8_c_3070_n ) capacitor c=9.64732e-19 //x=26.27 \
 //y=0 //x2=28.86 //y2=3.33
cc_129 ( N_GND_c_10_p N_noxref_8_c_3071_n ) capacitor c=0.0152765f //x=29.6 \
 //y=0 //x2=30.71 //y2=2.08
cc_130 ( N_GND_c_130_p N_noxref_8_c_3072_n ) capacitor c=0.00135046f \
 //x=30.695 //y=0 //x2=30.515 //y2=0.865
cc_131 ( N_GND_M18_noxref_d N_noxref_8_c_3072_n ) capacitor c=0.00220047f \
 //x=30.59 //y=0.865 //x2=30.515 //y2=0.865
cc_132 ( N_GND_M18_noxref_d N_noxref_8_c_3074_n ) capacitor c=0.00255985f \
 //x=30.59 //y=0.865 //x2=30.515 //y2=1.21
cc_133 ( N_GND_c_10_p N_noxref_8_c_3075_n ) capacitor c=0.0018059f //x=29.6 \
 //y=0 //x2=30.515 //y2=1.52
cc_134 ( N_GND_c_10_p N_noxref_8_c_3076_n ) capacitor c=0.0114883f //x=29.6 \
 //y=0 //x2=30.515 //y2=1.915
cc_135 ( N_GND_M18_noxref_d N_noxref_8_c_3077_n ) capacitor c=0.0131326f \
 //x=30.59 //y=0.865 //x2=30.89 //y2=0.71
cc_136 ( N_GND_M18_noxref_d N_noxref_8_c_3078_n ) capacitor c=0.00193127f \
 //x=30.59 //y=0.865 //x2=30.89 //y2=1.365
cc_137 ( N_GND_c_137_p N_noxref_8_c_3079_n ) capacitor c=0.00130622f //x=32.76 \
 //y=0 //x2=31.045 //y2=0.865
cc_138 ( N_GND_M18_noxref_d N_noxref_8_c_3079_n ) capacitor c=0.00257848f \
 //x=30.59 //y=0.865 //x2=31.045 //y2=0.865
cc_139 ( N_GND_M18_noxref_d N_noxref_8_c_3081_n ) capacitor c=0.00255985f \
 //x=30.59 //y=0.865 //x2=31.045 //y2=1.21
cc_140 ( N_GND_c_9_p N_noxref_8_M17_noxref_d ) capacitor c=8.58106e-19 \
 //x=26.27 //y=0 //x2=28.23 //y2=0.905
cc_141 ( N_GND_c_10_p N_noxref_8_M17_noxref_d ) capacitor c=0.00616547f \
 //x=29.6 //y=0 //x2=28.23 //y2=0.905
cc_142 ( N_GND_M16_noxref_d N_noxref_8_M17_noxref_d ) capacitor c=0.00143464f \
 //x=27.26 //y=0.865 //x2=28.23 //y2=0.905
cc_143 ( N_GND_c_11_p N_noxref_9_c_3300_n ) capacitor c=0.0436694f //x=32.93 \
 //y=0 //x2=32.105 //y2=1.655
cc_144 ( N_GND_c_10_p N_noxref_9_c_3301_n ) capacitor c=9.64732e-19 //x=29.6 \
 //y=0 //x2=32.19 //y2=3.33
cc_145 ( N_GND_c_11_p N_noxref_9_c_3302_n ) capacitor c=0.0153491f //x=32.93 \
 //y=0 //x2=34.04 //y2=2.08
cc_146 ( N_GND_c_146_p N_noxref_9_c_3303_n ) capacitor c=0.00135046f \
 //x=34.025 //y=0 //x2=33.845 //y2=0.865
cc_147 ( N_GND_M20_noxref_d N_noxref_9_c_3303_n ) capacitor c=0.00220047f \
 //x=33.92 //y=0.865 //x2=33.845 //y2=0.865
cc_148 ( N_GND_M20_noxref_d N_noxref_9_c_3305_n ) capacitor c=0.00255985f \
 //x=33.92 //y=0.865 //x2=33.845 //y2=1.21
cc_149 ( N_GND_c_11_p N_noxref_9_c_3306_n ) capacitor c=0.0018059f //x=32.93 \
 //y=0 //x2=33.845 //y2=1.52
cc_150 ( N_GND_c_11_p N_noxref_9_c_3307_n ) capacitor c=0.0114883f //x=32.93 \
 //y=0 //x2=33.845 //y2=1.915
cc_151 ( N_GND_M20_noxref_d N_noxref_9_c_3308_n ) capacitor c=0.0131326f \
 //x=33.92 //y=0.865 //x2=34.22 //y2=0.71
cc_152 ( N_GND_M20_noxref_d N_noxref_9_c_3309_n ) capacitor c=0.00193127f \
 //x=33.92 //y=0.865 //x2=34.22 //y2=1.365
cc_153 ( N_GND_c_153_p N_noxref_9_c_3310_n ) capacitor c=0.00130622f //x=36.09 \
 //y=0 //x2=34.375 //y2=0.865
cc_154 ( N_GND_M20_noxref_d N_noxref_9_c_3310_n ) capacitor c=0.00257848f \
 //x=33.92 //y=0.865 //x2=34.375 //y2=0.865
cc_155 ( N_GND_M20_noxref_d N_noxref_9_c_3312_n ) capacitor c=0.00255985f \
 //x=33.92 //y=0.865 //x2=34.375 //y2=1.21
cc_156 ( N_GND_c_10_p N_noxref_9_M19_noxref_d ) capacitor c=8.58106e-19 \
 //x=29.6 //y=0 //x2=31.56 //y2=0.905
cc_157 ( N_GND_c_11_p N_noxref_9_M19_noxref_d ) capacitor c=0.00616547f \
 //x=32.93 //y=0 //x2=31.56 //y2=0.905
cc_158 ( N_GND_M18_noxref_d N_noxref_9_M19_noxref_d ) capacitor c=0.00143464f \
 //x=30.59 //y=0.865 //x2=31.56 //y2=0.905
cc_159 ( N_GND_c_9_p N_noxref_10_c_3453_n ) capacitor c=0.0432803f //x=26.27 \
 //y=0 //x2=25.445 //y2=1.665
cc_160 ( N_GND_c_9_p N_noxref_10_c_3454_n ) capacitor c=0.0152578f //x=26.27 \
 //y=0 //x2=27.38 //y2=2.08
cc_161 ( N_GND_c_12_p N_noxref_10_c_3455_n ) capacitor c=0.0151426f //x=36.26 \
 //y=0 //x2=37.37 //y2=2.08
cc_162 ( N_GND_c_162_p N_noxref_10_c_3456_n ) capacitor c=0.00135046f \
 //x=27.365 //y=0 //x2=27.185 //y2=0.865
cc_163 ( N_GND_M16_noxref_d N_noxref_10_c_3456_n ) capacitor c=0.00220047f \
 //x=27.26 //y=0.865 //x2=27.185 //y2=0.865
cc_164 ( N_GND_M16_noxref_d N_noxref_10_c_3458_n ) capacitor c=0.00255985f \
 //x=27.26 //y=0.865 //x2=27.185 //y2=1.21
cc_165 ( N_GND_c_9_p N_noxref_10_c_3459_n ) capacitor c=0.00189421f //x=26.27 \
 //y=0 //x2=27.185 //y2=1.52
cc_166 ( N_GND_c_9_p N_noxref_10_c_3460_n ) capacitor c=0.0114883f //x=26.27 \
 //y=0 //x2=27.185 //y2=1.915
cc_167 ( N_GND_M16_noxref_d N_noxref_10_c_3461_n ) capacitor c=0.0131326f \
 //x=27.26 //y=0.865 //x2=27.56 //y2=0.71
cc_168 ( N_GND_M16_noxref_d N_noxref_10_c_3462_n ) capacitor c=0.00193127f \
 //x=27.26 //y=0.865 //x2=27.56 //y2=1.365
cc_169 ( N_GND_c_169_p N_noxref_10_c_3463_n ) capacitor c=0.00130622f \
 //x=29.43 //y=0 //x2=27.715 //y2=0.865
cc_170 ( N_GND_M16_noxref_d N_noxref_10_c_3463_n ) capacitor c=0.00257848f \
 //x=27.26 //y=0.865 //x2=27.715 //y2=0.865
cc_171 ( N_GND_M16_noxref_d N_noxref_10_c_3465_n ) capacitor c=0.00255985f \
 //x=27.26 //y=0.865 //x2=27.715 //y2=1.21
cc_172 ( N_GND_c_172_p N_noxref_10_c_3466_n ) capacitor c=0.00135046f \
 //x=37.355 //y=0 //x2=37.175 //y2=0.865
cc_173 ( N_GND_M22_noxref_d N_noxref_10_c_3466_n ) capacitor c=0.00220047f \
 //x=37.25 //y=0.865 //x2=37.175 //y2=0.865
cc_174 ( N_GND_M22_noxref_d N_noxref_10_c_3468_n ) capacitor c=0.00255985f \
 //x=37.25 //y=0.865 //x2=37.175 //y2=1.21
cc_175 ( N_GND_c_12_p N_noxref_10_c_3469_n ) capacitor c=0.0018059f //x=36.26 \
 //y=0 //x2=37.175 //y2=1.52
cc_176 ( N_GND_c_12_p N_noxref_10_c_3470_n ) capacitor c=0.0106743f //x=36.26 \
 //y=0 //x2=37.175 //y2=1.915
cc_177 ( N_GND_M22_noxref_d N_noxref_10_c_3471_n ) capacitor c=0.0131326f \
 //x=37.25 //y=0.865 //x2=37.55 //y2=0.71
cc_178 ( N_GND_M22_noxref_d N_noxref_10_c_3472_n ) capacitor c=0.00193127f \
 //x=37.25 //y=0.865 //x2=37.55 //y2=1.365
cc_179 ( N_GND_c_179_p N_noxref_10_c_3473_n ) capacitor c=0.00130622f \
 //x=39.42 //y=0 //x2=37.705 //y2=0.865
cc_180 ( N_GND_M22_noxref_d N_noxref_10_c_3473_n ) capacitor c=0.00257848f \
 //x=37.25 //y=0.865 //x2=37.705 //y2=0.865
cc_181 ( N_GND_M22_noxref_d N_noxref_10_c_3475_n ) capacitor c=0.00255985f \
 //x=37.25 //y=0.865 //x2=37.705 //y2=1.21
cc_182 ( N_GND_c_9_p N_noxref_10_M15_noxref_d ) capacitor c=0.00591582f \
 //x=26.27 //y=0 //x2=24.855 //y2=0.915
cc_183 ( N_GND_c_13_p N_noxref_11_c_3711_n ) capacitor c=0.0408098f //x=39.59 \
 //y=0 //x2=38.765 //y2=1.655
cc_184 ( N_GND_c_12_p N_noxref_11_c_3712_n ) capacitor c=9.64732e-19 //x=36.26 \
 //y=0 //x2=38.85 //y2=3.7
cc_185 ( N_GND_c_13_p N_noxref_11_c_3713_n ) capacitor c=0.0130105f //x=39.59 \
 //y=0 //x2=40.7 //y2=2.08
cc_186 ( N_GND_c_186_p N_noxref_11_c_3714_n ) capacitor c=0.00135046f \
 //x=40.685 //y=0 //x2=40.505 //y2=0.865
cc_187 ( N_GND_M24_noxref_d N_noxref_11_c_3714_n ) capacitor c=0.00220047f \
 //x=40.58 //y=0.865 //x2=40.505 //y2=0.865
cc_188 ( N_GND_M24_noxref_d N_noxref_11_c_3716_n ) capacitor c=0.00255985f \
 //x=40.58 //y=0.865 //x2=40.505 //y2=1.21
cc_189 ( N_GND_c_13_p N_noxref_11_c_3717_n ) capacitor c=0.0018059f //x=39.59 \
 //y=0 //x2=40.505 //y2=1.52
cc_190 ( N_GND_c_13_p N_noxref_11_c_3718_n ) capacitor c=0.00992619f //x=39.59 \
 //y=0 //x2=40.505 //y2=1.915
cc_191 ( N_GND_M24_noxref_d N_noxref_11_c_3719_n ) capacitor c=0.0131326f \
 //x=40.58 //y=0.865 //x2=40.88 //y2=0.71
cc_192 ( N_GND_M24_noxref_d N_noxref_11_c_3720_n ) capacitor c=0.00193127f \
 //x=40.58 //y=0.865 //x2=40.88 //y2=1.365
cc_193 ( N_GND_c_193_p N_noxref_11_c_3721_n ) capacitor c=0.00130622f \
 //x=42.75 //y=0 //x2=41.035 //y2=0.865
cc_194 ( N_GND_M24_noxref_d N_noxref_11_c_3721_n ) capacitor c=0.00257848f \
 //x=40.58 //y=0.865 //x2=41.035 //y2=0.865
cc_195 ( N_GND_M24_noxref_d N_noxref_11_c_3723_n ) capacitor c=0.00255985f \
 //x=40.58 //y=0.865 //x2=41.035 //y2=1.21
cc_196 ( N_GND_c_12_p N_noxref_11_M23_noxref_d ) capacitor c=8.58106e-19 \
 //x=36.26 //y=0 //x2=38.22 //y2=0.905
cc_197 ( N_GND_c_13_p N_noxref_11_M23_noxref_d ) capacitor c=0.00616547f \
 //x=39.59 //y=0 //x2=38.22 //y2=0.905
cc_198 ( N_GND_M22_noxref_d N_noxref_11_M23_noxref_d ) capacitor c=0.00143464f \
 //x=37.25 //y=0.865 //x2=38.22 //y2=0.905
cc_199 ( N_GND_c_8_p N_noxref_12_c_3862_n ) capacitor c=0.0153336f //x=21.46 \
 //y=0 //x2=22.57 //y2=2.08
cc_200 ( N_GND_c_10_p N_noxref_12_c_3863_n ) capacitor c=8.24484e-19 //x=29.6 \
 //y=0 //x2=31.45 //y2=2.08
cc_201 ( N_GND_c_11_p N_noxref_12_c_3863_n ) capacitor c=7.09207e-19 //x=32.93 \
 //y=0 //x2=31.45 //y2=2.08
cc_202 ( N_GND_c_12_p N_noxref_12_c_3865_n ) capacitor c=0.0432816f //x=36.26 \
 //y=0 //x2=35.435 //y2=1.655
cc_203 ( N_GND_c_11_p N_noxref_12_c_3866_n ) capacitor c=9.64732e-19 //x=32.93 \
 //y=0 //x2=35.52 //y2=4.07
cc_204 ( N_GND_c_13_p N_noxref_12_c_3867_n ) capacitor c=6.07681e-19 //x=39.59 \
 //y=0 //x2=41.44 //y2=2.08
cc_205 ( N_GND_c_14_p N_noxref_12_c_3867_n ) capacitor c=6.28327e-19 //x=42.92 \
 //y=0 //x2=41.44 //y2=2.08
cc_206 ( N_GND_c_206_p N_noxref_12_c_3869_n ) capacitor c=0.00132755f \
 //x=22.45 //y=0 //x2=22.27 //y2=0.875
cc_207 ( N_GND_M13_noxref_d N_noxref_12_c_3869_n ) capacitor c=0.00211996f \
 //x=22.345 //y=0.875 //x2=22.27 //y2=0.875
cc_208 ( N_GND_M13_noxref_d N_noxref_12_c_3871_n ) capacitor c=0.00255985f \
 //x=22.345 //y=0.875 //x2=22.27 //y2=1.22
cc_209 ( N_GND_c_8_p N_noxref_12_c_3872_n ) capacitor c=0.00195164f //x=21.46 \
 //y=0 //x2=22.27 //y2=1.53
cc_210 ( N_GND_c_8_p N_noxref_12_c_3873_n ) capacitor c=0.0126573f //x=21.46 \
 //y=0 //x2=22.27 //y2=1.915
cc_211 ( N_GND_M13_noxref_d N_noxref_12_c_3874_n ) capacitor c=0.0131341f \
 //x=22.345 //y=0.875 //x2=22.645 //y2=0.72
cc_212 ( N_GND_M13_noxref_d N_noxref_12_c_3875_n ) capacitor c=0.00193146f \
 //x=22.345 //y=0.875 //x2=22.645 //y2=1.375
cc_213 ( N_GND_c_213_p N_noxref_12_c_3876_n ) capacitor c=0.00129018f //x=26.1 \
 //y=0 //x2=22.8 //y2=0.875
cc_214 ( N_GND_M13_noxref_d N_noxref_12_c_3876_n ) capacitor c=0.00257848f \
 //x=22.345 //y=0.875 //x2=22.8 //y2=0.875
cc_215 ( N_GND_M13_noxref_d N_noxref_12_c_3878_n ) capacitor c=0.00255985f \
 //x=22.345 //y=0.875 //x2=22.8 //y2=1.22
cc_216 ( N_GND_c_11_p N_noxref_12_M21_noxref_d ) capacitor c=8.58106e-19 \
 //x=32.93 //y=0 //x2=34.89 //y2=0.905
cc_217 ( N_GND_c_12_p N_noxref_12_M21_noxref_d ) capacitor c=0.00616547f \
 //x=36.26 //y=0 //x2=34.89 //y2=0.905
cc_218 ( N_GND_M20_noxref_d N_noxref_12_M21_noxref_d ) capacitor c=0.00143464f \
 //x=33.92 //y=0.865 //x2=34.89 //y2=0.905
cc_219 ( N_GND_c_23_p N_D_c_4217_n ) capacitor c=0.175795f //x=73.63 //y=0 \
 //x2=28.005 //y2=2.59
cc_220 ( N_GND_c_74_p N_D_c_4217_n ) capacitor c=0.00251335f //x=7.97 //y=0 \
 //x2=28.005 //y2=2.59
cc_221 ( N_GND_c_33_p N_D_c_4217_n ) capacitor c=0.00280978f //x=9.235 //y=0 \
 //x2=28.005 //y2=2.59
cc_222 ( N_GND_c_40_p N_D_c_4217_n ) capacitor c=0.00326905f //x=11.3 //y=0 \
 //x2=28.005 //y2=2.59
cc_223 ( N_GND_c_50_p N_D_c_4217_n ) capacitor c=0.00280978f //x=12.565 //y=0 \
 //x2=28.005 //y2=2.59
cc_224 ( N_GND_c_57_p N_D_c_4217_n ) capacitor c=0.00326905f //x=14.63 //y=0 \
 //x2=28.005 //y2=2.59
cc_225 ( N_GND_c_77_p N_D_c_4217_n ) capacitor c=0.00280978f //x=15.895 //y=0 \
 //x2=28.005 //y2=2.59
cc_226 ( N_GND_c_84_p N_D_c_4217_n ) capacitor c=0.00326905f //x=17.96 //y=0 \
 //x2=28.005 //y2=2.59
cc_227 ( N_GND_c_91_p N_D_c_4217_n ) capacitor c=0.00280978f //x=19.225 //y=0 \
 //x2=28.005 //y2=2.59
cc_228 ( N_GND_c_98_p N_D_c_4217_n ) capacitor c=0.00326905f //x=21.29 //y=0 \
 //x2=28.005 //y2=2.59
cc_229 ( N_GND_c_206_p N_D_c_4217_n ) capacitor c=0.00221947f //x=22.45 //y=0 \
 //x2=28.005 //y2=2.59
cc_230 ( N_GND_c_213_p N_D_c_4217_n ) capacitor c=0.00344363f //x=26.1 //y=0 \
 //x2=28.005 //y2=2.59
cc_231 ( N_GND_c_162_p N_D_c_4217_n ) capacitor c=0.00280978f //x=27.365 //y=0 \
 //x2=28.005 //y2=2.59
cc_232 ( N_GND_c_4_p N_D_c_4217_n ) capacitor c=0.0360747f //x=8.14 //y=0 \
 //x2=28.005 //y2=2.59
cc_233 ( N_GND_c_5_p N_D_c_4217_n ) capacitor c=0.0360747f //x=11.47 //y=0 \
 //x2=28.005 //y2=2.59
cc_234 ( N_GND_c_6_p N_D_c_4217_n ) capacitor c=0.0377057f //x=14.8 //y=0 \
 //x2=28.005 //y2=2.59
cc_235 ( N_GND_c_7_p N_D_c_4217_n ) capacitor c=0.0338055f //x=18.13 //y=0 \
 //x2=28.005 //y2=2.59
cc_236 ( N_GND_c_8_p N_D_c_4217_n ) capacitor c=0.0338055f //x=21.46 //y=0 \
 //x2=28.005 //y2=2.59
cc_237 ( N_GND_c_9_p N_D_c_4217_n ) capacitor c=0.0338055f //x=26.27 //y=0 \
 //x2=28.005 //y2=2.59
cc_238 ( N_GND_c_23_p N_D_c_4236_n ) capacitor c=0.00219267f //x=73.63 //y=0 \
 //x2=6.775 //y2=2.59
cc_239 ( N_GND_c_74_p N_D_c_4236_n ) capacitor c=2.30913e-19 //x=7.97 //y=0 \
 //x2=6.775 //y2=2.59
cc_240 ( N_GND_c_23_p N_D_c_4238_n ) capacitor c=0.125054f //x=73.63 //y=0 \
 //x2=49.465 //y2=2.59
cc_241 ( N_GND_c_169_p N_D_c_4238_n ) capacitor c=0.00251335f //x=29.43 //y=0 \
 //x2=49.465 //y2=2.59
cc_242 ( N_GND_c_130_p N_D_c_4238_n ) capacitor c=0.00280978f //x=30.695 //y=0 \
 //x2=49.465 //y2=2.59
cc_243 ( N_GND_c_137_p N_D_c_4238_n ) capacitor c=0.00326905f //x=32.76 //y=0 \
 //x2=49.465 //y2=2.59
cc_244 ( N_GND_c_146_p N_D_c_4238_n ) capacitor c=0.00280978f //x=34.025 //y=0 \
 //x2=49.465 //y2=2.59
cc_245 ( N_GND_c_153_p N_D_c_4238_n ) capacitor c=0.00326905f //x=36.09 //y=0 \
 //x2=49.465 //y2=2.59
cc_246 ( N_GND_c_172_p N_D_c_4238_n ) capacitor c=0.00280978f //x=37.355 //y=0 \
 //x2=49.465 //y2=2.59
cc_247 ( N_GND_c_10_p N_D_c_4238_n ) capacitor c=0.0338055f //x=29.6 //y=0 \
 //x2=49.465 //y2=2.59
cc_248 ( N_GND_c_11_p N_D_c_4238_n ) capacitor c=0.0338055f //x=32.93 //y=0 \
 //x2=49.465 //y2=2.59
cc_249 ( N_GND_c_12_p N_D_c_4238_n ) capacitor c=0.0338055f //x=36.26 //y=0 \
 //x2=49.465 //y2=2.59
cc_250 ( N_GND_c_13_p N_D_c_4238_n ) capacitor c=0.0215583f //x=39.59 //y=0 \
 //x2=49.465 //y2=2.59
cc_251 ( N_GND_c_14_p N_D_c_4238_n ) capacitor c=0.0215583f //x=42.92 //y=0 \
 //x2=49.465 //y2=2.59
cc_252 ( N_GND_c_15_p N_D_c_4238_n ) capacitor c=0.0215583f //x=47.73 //y=0 \
 //x2=49.465 //y2=2.59
cc_253 ( N_GND_c_23_p N_D_c_4251_n ) capacitor c=0.00193173f //x=73.63 //y=0 \
 //x2=28.235 //y2=2.59
cc_254 ( N_GND_c_169_p N_D_c_4251_n ) capacitor c=2.30913e-19 //x=29.43 //y=0 \
 //x2=28.235 //y2=2.59
cc_255 ( N_GND_c_3_p N_D_c_4253_n ) capacitor c=0.00100253f //x=4.81 //y=0 \
 //x2=6.66 //y2=2.08
cc_256 ( N_GND_c_4_p N_D_c_4253_n ) capacitor c=7.51387e-19 //x=8.14 //y=0 \
 //x2=6.66 //y2=2.08
cc_257 ( N_GND_c_9_p N_D_c_4255_n ) capacitor c=7.72952e-19 //x=26.27 //y=0 \
 //x2=28.12 //y2=2.08
cc_258 ( N_GND_c_10_p N_D_c_4255_n ) capacitor c=7.51387e-19 //x=29.6 //y=0 \
 //x2=28.12 //y2=2.08
cc_259 ( N_GND_c_15_p N_D_c_4257_n ) capacitor c=5.63192e-19 //x=47.73 //y=0 \
 //x2=49.58 //y2=2.08
cc_260 ( N_GND_c_16_p N_D_c_4257_n ) capacitor c=9.37396e-19 //x=51.06 //y=0 \
 //x2=49.58 //y2=2.08
cc_261 ( N_GND_c_15_p N_noxref_14_c_4641_n ) capacitor c=6.05804e-19 //x=47.73 \
 //y=0 //x2=46.25 //y2=2.08
cc_262 ( N_GND_c_16_p N_noxref_14_c_4642_n ) capacitor c=0.0430593f //x=51.06 \
 //y=0 //x2=50.235 //y2=1.655
cc_263 ( N_GND_c_15_p N_noxref_14_c_4643_n ) capacitor c=9.64732e-19 //x=47.73 \
 //y=0 //x2=50.32 //y2=3.33
cc_264 ( N_GND_c_16_p N_noxref_14_c_4644_n ) capacitor c=0.0154158f //x=51.06 \
 //y=0 //x2=52.17 //y2=2.08
cc_265 ( N_GND_c_265_p N_noxref_14_c_4645_n ) capacitor c=0.00135046f \
 //x=52.155 //y=0 //x2=51.975 //y2=0.865
cc_266 ( N_GND_M31_noxref_d N_noxref_14_c_4645_n ) capacitor c=0.00220047f \
 //x=52.05 //y=0.865 //x2=51.975 //y2=0.865
cc_267 ( N_GND_M31_noxref_d N_noxref_14_c_4647_n ) capacitor c=0.00255985f \
 //x=52.05 //y=0.865 //x2=51.975 //y2=1.21
cc_268 ( N_GND_c_16_p N_noxref_14_c_4648_n ) capacitor c=0.0018059f //x=51.06 \
 //y=0 //x2=51.975 //y2=1.52
cc_269 ( N_GND_c_16_p N_noxref_14_c_4649_n ) capacitor c=0.0101006f //x=51.06 \
 //y=0 //x2=51.975 //y2=1.915
cc_270 ( N_GND_M31_noxref_d N_noxref_14_c_4650_n ) capacitor c=0.0131326f \
 //x=52.05 //y=0.865 //x2=52.35 //y2=0.71
cc_271 ( N_GND_M31_noxref_d N_noxref_14_c_4651_n ) capacitor c=0.00193127f \
 //x=52.05 //y=0.865 //x2=52.35 //y2=1.365
cc_272 ( N_GND_c_272_p N_noxref_14_c_4652_n ) capacitor c=0.00130622f \
 //x=54.22 //y=0 //x2=52.505 //y2=0.865
cc_273 ( N_GND_M31_noxref_d N_noxref_14_c_4652_n ) capacitor c=0.00257848f \
 //x=52.05 //y=0.865 //x2=52.505 //y2=0.865
cc_274 ( N_GND_M31_noxref_d N_noxref_14_c_4654_n ) capacitor c=0.00255985f \
 //x=52.05 //y=0.865 //x2=52.505 //y2=1.21
cc_275 ( N_GND_c_15_p N_noxref_14_M30_noxref_d ) capacitor c=8.58106e-19 \
 //x=47.73 //y=0 //x2=49.69 //y2=0.905
cc_276 ( N_GND_c_16_p N_noxref_14_M30_noxref_d ) capacitor c=0.00616547f \
 //x=51.06 //y=0 //x2=49.69 //y2=0.905
cc_277 ( N_GND_M29_noxref_d N_noxref_14_M30_noxref_d ) capacitor c=0.00143464f \
 //x=48.72 //y=0.865 //x2=49.69 //y2=0.905
cc_278 ( N_GND_c_17_p N_noxref_15_c_4874_n ) capacitor c=0.0436694f //x=54.39 \
 //y=0 //x2=53.565 //y2=1.655
cc_279 ( N_GND_c_16_p N_noxref_15_c_4875_n ) capacitor c=9.64732e-19 //x=51.06 \
 //y=0 //x2=53.65 //y2=3.33
cc_280 ( N_GND_c_17_p N_noxref_15_c_4876_n ) capacitor c=0.0156954f //x=54.39 \
 //y=0 //x2=55.5 //y2=2.08
cc_281 ( N_GND_c_281_p N_noxref_15_c_4877_n ) capacitor c=0.00135046f \
 //x=55.485 //y=0 //x2=55.305 //y2=0.865
cc_282 ( N_GND_M33_noxref_d N_noxref_15_c_4877_n ) capacitor c=0.00220047f \
 //x=55.38 //y=0.865 //x2=55.305 //y2=0.865
cc_283 ( N_GND_M33_noxref_d N_noxref_15_c_4879_n ) capacitor c=0.00255985f \
 //x=55.38 //y=0.865 //x2=55.305 //y2=1.21
cc_284 ( N_GND_c_17_p N_noxref_15_c_4880_n ) capacitor c=0.0018059f //x=54.39 \
 //y=0 //x2=55.305 //y2=1.52
cc_285 ( N_GND_c_17_p N_noxref_15_c_4881_n ) capacitor c=0.0101006f //x=54.39 \
 //y=0 //x2=55.305 //y2=1.915
cc_286 ( N_GND_M33_noxref_d N_noxref_15_c_4882_n ) capacitor c=0.0131326f \
 //x=55.38 //y=0.865 //x2=55.68 //y2=0.71
cc_287 ( N_GND_M33_noxref_d N_noxref_15_c_4883_n ) capacitor c=0.00193127f \
 //x=55.38 //y=0.865 //x2=55.68 //y2=1.365
cc_288 ( N_GND_c_288_p N_noxref_15_c_4884_n ) capacitor c=0.00130622f \
 //x=57.55 //y=0 //x2=55.835 //y2=0.865
cc_289 ( N_GND_M33_noxref_d N_noxref_15_c_4884_n ) capacitor c=0.00257848f \
 //x=55.38 //y=0.865 //x2=55.835 //y2=0.865
cc_290 ( N_GND_M33_noxref_d N_noxref_15_c_4886_n ) capacitor c=0.00255985f \
 //x=55.38 //y=0.865 //x2=55.835 //y2=1.21
cc_291 ( N_GND_c_16_p N_noxref_15_M32_noxref_d ) capacitor c=8.58106e-19 \
 //x=51.06 //y=0 //x2=53.02 //y2=0.905
cc_292 ( N_GND_c_17_p N_noxref_15_M32_noxref_d ) capacitor c=0.00616547f \
 //x=54.39 //y=0 //x2=53.02 //y2=0.905
cc_293 ( N_GND_M31_noxref_d N_noxref_15_M32_noxref_d ) capacitor c=0.00143464f \
 //x=52.05 //y=0.865 //x2=53.02 //y2=0.905
cc_294 ( N_GND_c_1_p N_CLK_c_5025_n ) capacitor c=7.64246e-19 //x=0.74 //y=0 \
 //x2=2.22 //y2=2.08
cc_295 ( N_GND_c_5_p N_CLK_c_5026_n ) capacitor c=7.51486e-19 //x=11.47 //y=0 \
 //x2=13.32 //y2=2.08
cc_296 ( N_GND_c_6_p N_CLK_c_5026_n ) capacitor c=7.09207e-19 //x=14.8 //y=0 \
 //x2=13.32 //y2=2.08
cc_297 ( N_GND_c_8_p N_CLK_c_5028_n ) capacitor c=6.4925e-19 //x=21.46 //y=0 \
 //x2=23.68 //y2=2.08
cc_298 ( N_GND_c_11_p N_CLK_c_5029_n ) capacitor c=7.51486e-19 //x=32.93 //y=0 \
 //x2=34.78 //y2=2.08
cc_299 ( N_GND_c_12_p N_CLK_c_5029_n ) capacitor c=8.18953e-19 //x=36.26 //y=0 \
 //x2=34.78 //y2=2.08
cc_300 ( N_GND_c_14_p N_CLK_c_5031_n ) capacitor c=4.85592e-19 //x=42.92 //y=0 \
 //x2=45.14 //y2=2.08
cc_301 ( N_GND_c_17_p N_CLK_c_5032_n ) capacitor c=7.1088e-19 //x=54.39 //y=0 \
 //x2=56.24 //y2=2.08
cc_302 ( N_GND_c_18_p N_CLK_c_5032_n ) capacitor c=7.76678e-19 //x=57.72 //y=0 \
 //x2=56.24 //y2=2.08
cc_303 ( N_GND_c_15_p N_noxref_17_c_5777_n ) capacitor c=0.040668f //x=47.73 \
 //y=0 //x2=46.905 //y2=1.665
cc_304 ( N_GND_c_15_p N_noxref_17_c_5778_n ) capacitor c=0.0130128f //x=47.73 \
 //y=0 //x2=48.84 //y2=2.08
cc_305 ( N_GND_c_18_p N_noxref_17_c_5779_n ) capacitor c=0.0156954f //x=57.72 \
 //y=0 //x2=58.83 //y2=2.08
cc_306 ( N_GND_c_306_p N_noxref_17_c_5780_n ) capacitor c=0.00135046f \
 //x=48.825 //y=0 //x2=48.645 //y2=0.865
cc_307 ( N_GND_M29_noxref_d N_noxref_17_c_5780_n ) capacitor c=0.00220047f \
 //x=48.72 //y=0.865 //x2=48.645 //y2=0.865
cc_308 ( N_GND_M29_noxref_d N_noxref_17_c_5782_n ) capacitor c=0.00255985f \
 //x=48.72 //y=0.865 //x2=48.645 //y2=1.21
cc_309 ( N_GND_c_15_p N_noxref_17_c_5783_n ) capacitor c=0.00189421f //x=47.73 \
 //y=0 //x2=48.645 //y2=1.52
cc_310 ( N_GND_c_15_p N_noxref_17_c_5784_n ) capacitor c=0.0101006f //x=47.73 \
 //y=0 //x2=48.645 //y2=1.915
cc_311 ( N_GND_M29_noxref_d N_noxref_17_c_5785_n ) capacitor c=0.0131326f \
 //x=48.72 //y=0.865 //x2=49.02 //y2=0.71
cc_312 ( N_GND_M29_noxref_d N_noxref_17_c_5786_n ) capacitor c=0.00193127f \
 //x=48.72 //y=0.865 //x2=49.02 //y2=1.365
cc_313 ( N_GND_c_313_p N_noxref_17_c_5787_n ) capacitor c=0.00130622f \
 //x=50.89 //y=0 //x2=49.175 //y2=0.865
cc_314 ( N_GND_M29_noxref_d N_noxref_17_c_5787_n ) capacitor c=0.00257848f \
 //x=48.72 //y=0.865 //x2=49.175 //y2=0.865
cc_315 ( N_GND_M29_noxref_d N_noxref_17_c_5789_n ) capacitor c=0.00255985f \
 //x=48.72 //y=0.865 //x2=49.175 //y2=1.21
cc_316 ( N_GND_c_316_p N_noxref_17_c_5790_n ) capacitor c=0.00135046f \
 //x=58.815 //y=0 //x2=58.635 //y2=0.865
cc_317 ( N_GND_M35_noxref_d N_noxref_17_c_5790_n ) capacitor c=0.00220047f \
 //x=58.71 //y=0.865 //x2=58.635 //y2=0.865
cc_318 ( N_GND_M35_noxref_d N_noxref_17_c_5792_n ) capacitor c=0.00255985f \
 //x=58.71 //y=0.865 //x2=58.635 //y2=1.21
cc_319 ( N_GND_c_18_p N_noxref_17_c_5793_n ) capacitor c=0.0018059f //x=57.72 \
 //y=0 //x2=58.635 //y2=1.52
cc_320 ( N_GND_c_18_p N_noxref_17_c_5794_n ) capacitor c=0.0101006f //x=57.72 \
 //y=0 //x2=58.635 //y2=1.915
cc_321 ( N_GND_M35_noxref_d N_noxref_17_c_5795_n ) capacitor c=0.0131326f \
 //x=58.71 //y=0.865 //x2=59.01 //y2=0.71
cc_322 ( N_GND_M35_noxref_d N_noxref_17_c_5796_n ) capacitor c=0.00193127f \
 //x=58.71 //y=0.865 //x2=59.01 //y2=1.365
cc_323 ( N_GND_c_323_p N_noxref_17_c_5797_n ) capacitor c=0.00130622f \
 //x=60.88 //y=0 //x2=59.165 //y2=0.865
cc_324 ( N_GND_M35_noxref_d N_noxref_17_c_5797_n ) capacitor c=0.00257848f \
 //x=58.71 //y=0.865 //x2=59.165 //y2=0.865
cc_325 ( N_GND_M35_noxref_d N_noxref_17_c_5799_n ) capacitor c=0.00255985f \
 //x=58.71 //y=0.865 //x2=59.165 //y2=1.21
cc_326 ( N_GND_c_15_p N_noxref_17_M28_noxref_d ) capacitor c=0.00591582f \
 //x=47.73 //y=0 //x2=46.315 //y2=0.915
cc_327 ( N_GND_c_19_p N_noxref_18_c_6032_n ) capacitor c=0.0436694f //x=61.05 \
 //y=0 //x2=60.225 //y2=1.655
cc_328 ( N_GND_c_18_p N_noxref_18_c_6033_n ) capacitor c=9.64732e-19 //x=57.72 \
 //y=0 //x2=60.31 //y2=4.44
cc_329 ( N_GND_c_19_p N_noxref_18_c_6034_n ) capacitor c=0.0156954f //x=61.05 \
 //y=0 //x2=62.16 //y2=2.08
cc_330 ( N_GND_c_330_p N_noxref_18_c_6035_n ) capacitor c=0.00135046f \
 //x=62.145 //y=0 //x2=61.965 //y2=0.865
cc_331 ( N_GND_M37_noxref_d N_noxref_18_c_6035_n ) capacitor c=0.00220047f \
 //x=62.04 //y=0.865 //x2=61.965 //y2=0.865
cc_332 ( N_GND_M37_noxref_d N_noxref_18_c_6037_n ) capacitor c=0.00255985f \
 //x=62.04 //y=0.865 //x2=61.965 //y2=1.21
cc_333 ( N_GND_c_19_p N_noxref_18_c_6038_n ) capacitor c=0.0018059f //x=61.05 \
 //y=0 //x2=61.965 //y2=1.52
cc_334 ( N_GND_c_19_p N_noxref_18_c_6039_n ) capacitor c=0.0101006f //x=61.05 \
 //y=0 //x2=61.965 //y2=1.915
cc_335 ( N_GND_M37_noxref_d N_noxref_18_c_6040_n ) capacitor c=0.0131326f \
 //x=62.04 //y=0.865 //x2=62.34 //y2=0.71
cc_336 ( N_GND_M37_noxref_d N_noxref_18_c_6041_n ) capacitor c=0.00193127f \
 //x=62.04 //y=0.865 //x2=62.34 //y2=1.365
cc_337 ( N_GND_c_337_p N_noxref_18_c_6042_n ) capacitor c=0.00130622f \
 //x=64.21 //y=0 //x2=62.495 //y2=0.865
cc_338 ( N_GND_M37_noxref_d N_noxref_18_c_6042_n ) capacitor c=0.00257848f \
 //x=62.04 //y=0.865 //x2=62.495 //y2=0.865
cc_339 ( N_GND_M37_noxref_d N_noxref_18_c_6044_n ) capacitor c=0.00255985f \
 //x=62.04 //y=0.865 //x2=62.495 //y2=1.21
cc_340 ( N_GND_c_18_p N_noxref_18_M36_noxref_d ) capacitor c=8.58106e-19 \
 //x=57.72 //y=0 //x2=59.68 //y2=0.905
cc_341 ( N_GND_c_19_p N_noxref_18_M36_noxref_d ) capacitor c=0.00616547f \
 //x=61.05 //y=0 //x2=59.68 //y2=0.905
cc_342 ( N_GND_M35_noxref_d N_noxref_18_M36_noxref_d ) capacitor c=0.00143464f \
 //x=58.71 //y=0.865 //x2=59.68 //y2=0.905
cc_343 ( N_GND_c_14_p N_noxref_19_c_6190_n ) capacitor c=0.0130099f //x=42.92 \
 //y=0 //x2=44.03 //y2=2.08
cc_344 ( N_GND_c_16_p N_noxref_19_c_6191_n ) capacitor c=9.9063e-19 //x=51.06 \
 //y=0 //x2=52.91 //y2=2.08
cc_345 ( N_GND_c_17_p N_noxref_19_c_6191_n ) capacitor c=7.76678e-19 //x=54.39 \
 //y=0 //x2=52.91 //y2=2.08
cc_346 ( N_GND_c_18_p N_noxref_19_c_6193_n ) capacitor c=0.0436694f //x=57.72 \
 //y=0 //x2=56.895 //y2=1.655
cc_347 ( N_GND_c_17_p N_noxref_19_c_6194_n ) capacitor c=9.64732e-19 //x=54.39 \
 //y=0 //x2=56.98 //y2=4.07
cc_348 ( N_GND_c_19_p N_noxref_19_c_6195_n ) capacitor c=7.1088e-19 //x=61.05 \
 //y=0 //x2=62.9 //y2=2.08
cc_349 ( N_GND_c_20_p N_noxref_19_c_6195_n ) capacitor c=8.13269e-19 //x=64.38 \
 //y=0 //x2=62.9 //y2=2.08
cc_350 ( N_GND_c_350_p N_noxref_19_c_6197_n ) capacitor c=0.00132755f \
 //x=43.91 //y=0 //x2=43.73 //y2=0.875
cc_351 ( N_GND_M26_noxref_d N_noxref_19_c_6197_n ) capacitor c=0.00211996f \
 //x=43.805 //y=0.875 //x2=43.73 //y2=0.875
cc_352 ( N_GND_M26_noxref_d N_noxref_19_c_6199_n ) capacitor c=0.00255985f \
 //x=43.805 //y=0.875 //x2=43.73 //y2=1.22
cc_353 ( N_GND_c_14_p N_noxref_19_c_6200_n ) capacitor c=0.00195164f //x=42.92 \
 //y=0 //x2=43.73 //y2=1.53
cc_354 ( N_GND_c_14_p N_noxref_19_c_6201_n ) capacitor c=0.0110952f //x=42.92 \
 //y=0 //x2=43.73 //y2=1.915
cc_355 ( N_GND_M26_noxref_d N_noxref_19_c_6202_n ) capacitor c=0.0131341f \
 //x=43.805 //y=0.875 //x2=44.105 //y2=0.72
cc_356 ( N_GND_M26_noxref_d N_noxref_19_c_6203_n ) capacitor c=0.00193146f \
 //x=43.805 //y=0.875 //x2=44.105 //y2=1.375
cc_357 ( N_GND_c_357_p N_noxref_19_c_6204_n ) capacitor c=0.00129018f \
 //x=47.56 //y=0 //x2=44.26 //y2=0.875
cc_358 ( N_GND_M26_noxref_d N_noxref_19_c_6204_n ) capacitor c=0.00257848f \
 //x=43.805 //y=0.875 //x2=44.26 //y2=0.875
cc_359 ( N_GND_M26_noxref_d N_noxref_19_c_6206_n ) capacitor c=0.00255985f \
 //x=43.805 //y=0.875 //x2=44.26 //y2=1.22
cc_360 ( N_GND_c_17_p N_noxref_19_M34_noxref_d ) capacitor c=8.58106e-19 \
 //x=54.39 //y=0 //x2=56.35 //y2=0.905
cc_361 ( N_GND_c_18_p N_noxref_19_M34_noxref_d ) capacitor c=0.00616547f \
 //x=57.72 //y=0 //x2=56.35 //y2=0.905
cc_362 ( N_GND_M33_noxref_d N_noxref_19_M34_noxref_d ) capacitor c=0.00143464f \
 //x=55.38 //y=0.865 //x2=56.35 //y2=0.905
cc_363 ( N_GND_c_18_p N_noxref_20_c_6560_n ) capacitor c=7.1088e-19 //x=57.72 \
 //y=0 //x2=59.57 //y2=2.08
cc_364 ( N_GND_c_19_p N_noxref_20_c_6560_n ) capacitor c=7.76678e-19 //x=61.05 \
 //y=0 //x2=59.57 //y2=2.08
cc_365 ( N_GND_c_20_p N_noxref_20_c_6562_n ) capacitor c=0.043499f //x=64.38 \
 //y=0 //x2=63.555 //y2=1.655
cc_366 ( N_GND_c_19_p N_noxref_20_c_6563_n ) capacitor c=9.64732e-19 //x=61.05 \
 //y=0 //x2=63.64 //y2=3.7
cc_367 ( N_GND_c_23_p N_noxref_20_c_6564_n ) capacitor c=2.87616e-19 //x=73.63 \
 //y=0 //x2=65.12 //y2=2.08
cc_368 ( N_GND_c_20_p N_noxref_20_c_6564_n ) capacitor c=0.0269204f //x=64.38 \
 //y=0 //x2=65.12 //y2=2.08
cc_369 ( N_GND_c_21_p N_noxref_20_c_6564_n ) capacitor c=4.75835e-19 //x=67.71 \
 //y=0 //x2=65.12 //y2=2.08
cc_370 ( N_GND_c_21_p N_noxref_20_c_6567_n ) capacitor c=0.0177157f //x=67.71 \
 //y=0 //x2=68.82 //y2=2.08
cc_371 ( N_GND_c_22_p N_noxref_20_c_6567_n ) capacitor c=7.87427e-19 //x=71.04 \
 //y=0 //x2=68.82 //y2=2.08
cc_372 ( N_GND_c_372_p N_noxref_20_c_6569_n ) capacitor c=0.0013864f \
 //x=65.475 //y=0 //x2=65.295 //y2=0.865
cc_373 ( N_GND_M39_noxref_d N_noxref_20_c_6569_n ) capacitor c=0.00220047f \
 //x=65.37 //y=0.865 //x2=65.295 //y2=0.865
cc_374 ( N_GND_M39_noxref_d N_noxref_20_c_6571_n ) capacitor c=0.00255985f \
 //x=65.37 //y=0.865 //x2=65.295 //y2=1.21
cc_375 ( N_GND_c_20_p N_noxref_20_c_6572_n ) capacitor c=0.0018059f //x=64.38 \
 //y=0 //x2=65.295 //y2=1.52
cc_376 ( N_GND_c_20_p N_noxref_20_c_6573_n ) capacitor c=0.00369987f //x=64.38 \
 //y=0 //x2=65.295 //y2=1.915
cc_377 ( N_GND_M39_noxref_d N_noxref_20_c_6574_n ) capacitor c=0.0131326f \
 //x=65.37 //y=0.865 //x2=65.67 //y2=0.71
cc_378 ( N_GND_M39_noxref_d N_noxref_20_c_6575_n ) capacitor c=0.00193127f \
 //x=65.37 //y=0.865 //x2=65.67 //y2=1.365
cc_379 ( N_GND_c_379_p N_noxref_20_c_6576_n ) capacitor c=0.00130622f \
 //x=67.54 //y=0 //x2=65.825 //y2=0.865
cc_380 ( N_GND_M39_noxref_d N_noxref_20_c_6576_n ) capacitor c=0.00257848f \
 //x=65.37 //y=0.865 //x2=65.825 //y2=0.865
cc_381 ( N_GND_M39_noxref_d N_noxref_20_c_6578_n ) capacitor c=0.00255985f \
 //x=65.37 //y=0.865 //x2=65.825 //y2=1.21
cc_382 ( N_GND_c_382_p N_noxref_20_c_6579_n ) capacitor c=0.00135046f \
 //x=68.805 //y=0 //x2=68.625 //y2=0.865
cc_383 ( N_GND_M41_noxref_d N_noxref_20_c_6579_n ) capacitor c=0.00220047f \
 //x=68.7 //y=0.865 //x2=68.625 //y2=0.865
cc_384 ( N_GND_M41_noxref_d N_noxref_20_c_6581_n ) capacitor c=0.00272336f \
 //x=68.7 //y=0.865 //x2=68.625 //y2=1.21
cc_385 ( N_GND_c_21_p N_noxref_20_c_6582_n ) capacitor c=0.00976978f //x=67.71 \
 //y=0 //x2=68.625 //y2=1.915
cc_386 ( N_GND_M41_noxref_d N_noxref_20_c_6583_n ) capacitor c=0.0131326f \
 //x=68.7 //y=0.865 //x2=69 //y2=0.71
cc_387 ( N_GND_M41_noxref_d N_noxref_20_c_6584_n ) capacitor c=0.00167494f \
 //x=68.7 //y=0.865 //x2=69 //y2=1.365
cc_388 ( N_GND_c_388_p N_noxref_20_c_6585_n ) capacitor c=0.00130622f \
 //x=70.87 //y=0 //x2=69.155 //y2=0.865
cc_389 ( N_GND_M41_noxref_d N_noxref_20_c_6585_n ) capacitor c=0.00257848f \
 //x=68.7 //y=0.865 //x2=69.155 //y2=0.865
cc_390 ( N_GND_M41_noxref_d N_noxref_20_c_6587_n ) capacitor c=0.00272336f \
 //x=68.7 //y=0.865 //x2=69.155 //y2=1.21
cc_391 ( N_GND_c_20_p N_noxref_20_c_6588_n ) capacitor c=0.00888771f //x=64.38 \
 //y=0 //x2=65.12 //y2=2.08
cc_392 ( N_GND_c_19_p N_noxref_20_M38_noxref_d ) capacitor c=8.58106e-19 \
 //x=61.05 //y=0 //x2=63.01 //y2=0.905
cc_393 ( N_GND_c_20_p N_noxref_20_M38_noxref_d ) capacitor c=0.00616146f \
 //x=64.38 //y=0 //x2=63.01 //y2=0.905
cc_394 ( N_GND_M37_noxref_d N_noxref_20_M38_noxref_d ) capacitor c=0.00143464f \
 //x=62.04 //y=0.865 //x2=63.01 //y2=0.905
cc_395 ( N_GND_c_23_p N_noxref_21_c_6904_n ) capacitor c=0.036509f //x=73.63 \
 //y=0 //x2=42.065 //y2=2.22
cc_396 ( N_GND_c_179_p N_noxref_21_c_6904_n ) capacitor c=0.00311072f \
 //x=39.42 //y=0 //x2=42.065 //y2=2.22
cc_397 ( N_GND_c_186_p N_noxref_21_c_6904_n ) capacitor c=0.00347653f \
 //x=40.685 //y=0 //x2=42.065 //y2=2.22
cc_398 ( N_GND_c_193_p N_noxref_21_c_6904_n ) capacitor c=0.0010086f //x=42.75 \
 //y=0 //x2=42.065 //y2=2.22
cc_399 ( N_GND_c_13_p N_noxref_21_c_6904_n ) capacitor c=0.0379964f //x=39.59 \
 //y=0 //x2=42.065 //y2=2.22
cc_400 ( N_GND_c_23_p N_noxref_21_c_6909_n ) capacitor c=0.00214183f //x=73.63 \
 //y=0 //x2=38.225 //y2=2.22
cc_401 ( N_GND_c_179_p N_noxref_21_c_6909_n ) capacitor c=3.68204e-19 \
 //x=39.42 //y=0 //x2=38.225 //y2=2.22
cc_402 ( N_GND_c_23_p N_noxref_21_c_6911_n ) capacitor c=0.227735f //x=73.63 \
 //y=0 //x2=66.115 //y2=2.22
cc_403 ( N_GND_c_193_p N_noxref_21_c_6911_n ) capacitor c=0.00286739f \
 //x=42.75 //y=0 //x2=66.115 //y2=2.22
cc_404 ( N_GND_c_350_p N_noxref_21_c_6911_n ) capacitor c=0.00274252f \
 //x=43.91 //y=0 //x2=66.115 //y2=2.22
cc_405 ( N_GND_c_357_p N_noxref_21_c_6911_n ) capacitor c=0.00450506f \
 //x=47.56 //y=0 //x2=66.115 //y2=2.22
cc_406 ( N_GND_c_306_p N_noxref_21_c_6911_n ) capacitor c=0.00347653f \
 //x=48.825 //y=0 //x2=66.115 //y2=2.22
cc_407 ( N_GND_c_313_p N_noxref_21_c_6911_n ) capacitor c=0.00411932f \
 //x=50.89 //y=0 //x2=66.115 //y2=2.22
cc_408 ( N_GND_c_265_p N_noxref_21_c_6911_n ) capacitor c=0.00347653f \
 //x=52.155 //y=0 //x2=66.115 //y2=2.22
cc_409 ( N_GND_c_272_p N_noxref_21_c_6911_n ) capacitor c=0.00411932f \
 //x=54.22 //y=0 //x2=66.115 //y2=2.22
cc_410 ( N_GND_c_281_p N_noxref_21_c_6911_n ) capacitor c=0.00347653f \
 //x=55.485 //y=0 //x2=66.115 //y2=2.22
cc_411 ( N_GND_c_288_p N_noxref_21_c_6911_n ) capacitor c=0.00411932f \
 //x=57.55 //y=0 //x2=66.115 //y2=2.22
cc_412 ( N_GND_c_316_p N_noxref_21_c_6911_n ) capacitor c=0.00347653f \
 //x=58.815 //y=0 //x2=66.115 //y2=2.22
cc_413 ( N_GND_c_323_p N_noxref_21_c_6911_n ) capacitor c=0.00411932f \
 //x=60.88 //y=0 //x2=66.115 //y2=2.22
cc_414 ( N_GND_c_330_p N_noxref_21_c_6911_n ) capacitor c=0.00347653f \
 //x=62.145 //y=0 //x2=66.115 //y2=2.22
cc_415 ( N_GND_c_337_p N_noxref_21_c_6911_n ) capacitor c=0.00411932f \
 //x=64.21 //y=0 //x2=66.115 //y2=2.22
cc_416 ( N_GND_c_372_p N_noxref_21_c_6911_n ) capacitor c=0.00291512f \
 //x=65.475 //y=0 //x2=66.115 //y2=2.22
cc_417 ( N_GND_c_379_p N_noxref_21_c_6911_n ) capacitor c=3.68204e-19 \
 //x=67.54 //y=0 //x2=66.115 //y2=2.22
cc_418 ( N_GND_c_14_p N_noxref_21_c_6911_n ) capacitor c=0.0379964f //x=42.92 \
 //y=0 //x2=66.115 //y2=2.22
cc_419 ( N_GND_c_15_p N_noxref_21_c_6911_n ) capacitor c=0.0379964f //x=47.73 \
 //y=0 //x2=66.115 //y2=2.22
cc_420 ( N_GND_c_16_p N_noxref_21_c_6911_n ) capacitor c=0.0401775f //x=51.06 \
 //y=0 //x2=66.115 //y2=2.22
cc_421 ( N_GND_c_17_p N_noxref_21_c_6911_n ) capacitor c=0.0401775f //x=54.39 \
 //y=0 //x2=66.115 //y2=2.22
cc_422 ( N_GND_c_18_p N_noxref_21_c_6911_n ) capacitor c=0.0401775f //x=57.72 \
 //y=0 //x2=66.115 //y2=2.22
cc_423 ( N_GND_c_19_p N_noxref_21_c_6911_n ) capacitor c=0.0401775f //x=61.05 \
 //y=0 //x2=66.115 //y2=2.22
cc_424 ( N_GND_c_20_p N_noxref_21_c_6911_n ) capacitor c=0.0389307f //x=64.38 \
 //y=0 //x2=66.115 //y2=2.22
cc_425 ( N_GND_c_21_p N_noxref_21_c_6911_n ) capacitor c=0.00415531f //x=67.71 \
 //y=0 //x2=66.115 //y2=2.22
cc_426 ( N_GND_c_23_p N_noxref_21_c_6935_n ) capacitor c=0.00232052f //x=73.63 \
 //y=0 //x2=42.295 //y2=2.22
cc_427 ( N_GND_c_193_p N_noxref_21_c_6935_n ) capacitor c=2.19784e-19 \
 //x=42.75 //y=0 //x2=42.295 //y2=2.22
cc_428 ( N_GND_c_14_p N_noxref_21_c_6935_n ) capacitor c=0.00209945f //x=42.92 \
 //y=0 //x2=42.295 //y2=2.22
cc_429 ( N_GND_c_22_p N_noxref_21_c_6938_n ) capacitor c=0.00281233f //x=71.04 \
 //y=0 //x2=72.775 //y2=4.07
cc_430 ( N_GND_c_12_p N_noxref_21_c_6939_n ) capacitor c=7.74776e-19 //x=36.26 \
 //y=0 //x2=38.11 //y2=2.08
cc_431 ( N_GND_c_13_p N_noxref_21_c_6939_n ) capacitor c=5.93203e-19 //x=39.59 \
 //y=0 //x2=38.11 //y2=2.08
cc_432 ( N_GND_c_14_p N_noxref_21_c_6941_n ) capacitor c=0.0402988f //x=42.92 \
 //y=0 //x2=42.095 //y2=1.655
cc_433 ( N_GND_c_13_p N_noxref_21_c_6942_n ) capacitor c=9.64732e-19 //x=39.59 \
 //y=0 //x2=42.18 //y2=2.22
cc_434 ( N_GND_c_14_p N_noxref_21_c_6942_n ) capacitor c=5.56859e-19 //x=42.92 \
 //y=0 //x2=42.18 //y2=2.22
cc_435 ( N_GND_c_20_p N_noxref_21_c_6944_n ) capacitor c=9.60509e-19 //x=64.38 \
 //y=0 //x2=66.23 //y2=2.08
cc_436 ( N_GND_c_21_p N_noxref_21_c_6944_n ) capacitor c=0.0111266f //x=67.71 \
 //y=0 //x2=66.23 //y2=2.08
cc_437 ( N_GND_c_2_p N_noxref_21_c_6946_n ) capacitor c=0.00128267f //x=73.63 \
 //y=0 //x2=72.89 //y2=2.08
cc_438 ( N_GND_c_22_p N_noxref_21_c_6946_n ) capacitor c=8.50308e-19 //x=71.04 \
 //y=0 //x2=72.89 //y2=2.08
cc_439 ( N_GND_c_21_p N_noxref_21_c_6948_n ) capacitor c=2.63786e-19 //x=67.71 \
 //y=0 //x2=66.23 //y2=2.08
cc_440 ( N_GND_c_13_p N_noxref_21_M25_noxref_d ) capacitor c=8.58106e-19 \
 //x=39.59 //y=0 //x2=41.55 //y2=0.905
cc_441 ( N_GND_c_14_p N_noxref_21_M25_noxref_d ) capacitor c=0.00616547f \
 //x=42.92 //y=0 //x2=41.55 //y2=0.905
cc_442 ( N_GND_M24_noxref_d N_noxref_21_M25_noxref_d ) capacitor c=0.00143464f \
 //x=40.58 //y=0.865 //x2=41.55 //y2=0.905
cc_443 ( N_GND_c_7_p N_noxref_23_c_7497_n ) capacitor c=0.00750857f //x=18.13 \
 //y=0 //x2=20.605 //y2=2.96
cc_444 ( N_GND_c_23_p N_noxref_23_c_7498_n ) capacitor c=0.112259f //x=73.63 \
 //y=0 //x2=70.185 //y2=2.96
cc_445 ( N_GND_c_8_p N_noxref_23_c_7498_n ) capacitor c=0.00750857f //x=21.46 \
 //y=0 //x2=70.185 //y2=2.96
cc_446 ( N_GND_c_9_p N_noxref_23_c_7498_n ) capacitor c=0.00750857f //x=26.27 \
 //y=0 //x2=70.185 //y2=2.96
cc_447 ( N_GND_c_10_p N_noxref_23_c_7498_n ) capacitor c=0.00750857f //x=29.6 \
 //y=0 //x2=70.185 //y2=2.96
cc_448 ( N_GND_c_11_p N_noxref_23_c_7498_n ) capacitor c=0.00750857f //x=32.93 \
 //y=0 //x2=70.185 //y2=2.96
cc_449 ( N_GND_c_12_p N_noxref_23_c_7498_n ) capacitor c=0.00750857f //x=36.26 \
 //y=0 //x2=70.185 //y2=2.96
cc_450 ( N_GND_c_13_p N_noxref_23_c_7498_n ) capacitor c=0.00750857f //x=39.59 \
 //y=0 //x2=70.185 //y2=2.96
cc_451 ( N_GND_c_14_p N_noxref_23_c_7498_n ) capacitor c=0.00750857f //x=42.92 \
 //y=0 //x2=70.185 //y2=2.96
cc_452 ( N_GND_c_15_p N_noxref_23_c_7498_n ) capacitor c=0.00750857f //x=47.73 \
 //y=0 //x2=70.185 //y2=2.96
cc_453 ( N_GND_c_16_p N_noxref_23_c_7498_n ) capacitor c=0.00949826f //x=51.06 \
 //y=0 //x2=70.185 //y2=2.96
cc_454 ( N_GND_c_17_p N_noxref_23_c_7498_n ) capacitor c=0.00949826f //x=54.39 \
 //y=0 //x2=70.185 //y2=2.96
cc_455 ( N_GND_c_18_p N_noxref_23_c_7498_n ) capacitor c=0.00949826f //x=57.72 \
 //y=0 //x2=70.185 //y2=2.96
cc_456 ( N_GND_c_19_p N_noxref_23_c_7498_n ) capacitor c=0.00949826f //x=61.05 \
 //y=0 //x2=70.185 //y2=2.96
cc_457 ( N_GND_c_20_p N_noxref_23_c_7498_n ) capacitor c=0.00949826f //x=64.38 \
 //y=0 //x2=70.185 //y2=2.96
cc_458 ( N_GND_c_21_p N_noxref_23_c_7498_n ) capacitor c=0.0128764f //x=67.71 \
 //y=0 //x2=70.185 //y2=2.96
cc_459 ( N_GND_c_22_p N_noxref_23_c_7513_n ) capacitor c=0.0396043f //x=71.04 \
 //y=0 //x2=71.665 //y2=2.08
cc_460 ( N_GND_c_22_p N_noxref_23_c_7514_n ) capacitor c=0.00128384f //x=71.04 \
 //y=0 //x2=70.415 //y2=2.08
cc_461 ( N_GND_c_6_p N_noxref_23_c_7515_n ) capacitor c=7.51486e-19 //x=14.8 \
 //y=0 //x2=16.65 //y2=2.08
cc_462 ( N_GND_c_7_p N_noxref_23_c_7515_n ) capacitor c=7.09207e-19 //x=18.13 \
 //y=0 //x2=16.65 //y2=2.08
cc_463 ( N_GND_c_8_p N_noxref_23_c_7517_n ) capacitor c=0.0436242f //x=21.46 \
 //y=0 //x2=20.635 //y2=1.655
cc_464 ( N_GND_c_7_p N_noxref_23_c_7518_n ) capacitor c=9.64732e-19 //x=18.13 \
 //y=0 //x2=20.72 //y2=2.96
cc_465 ( N_GND_c_21_p N_noxref_23_c_7519_n ) capacitor c=6.95291e-19 //x=67.71 \
 //y=0 //x2=70.3 //y2=2.08
cc_466 ( N_GND_c_22_p N_noxref_23_c_7519_n ) capacitor c=0.0266762f //x=71.04 \
 //y=0 //x2=70.3 //y2=2.08
cc_467 ( N_GND_c_22_p N_noxref_23_c_7521_n ) capacitor c=0.0266762f //x=71.04 \
 //y=0 //x2=71.78 //y2=2.08
cc_468 ( N_GND_c_22_p N_noxref_23_c_7522_n ) capacitor c=0.0103285f //x=71.04 \
 //y=0 //x2=70.125 //y2=1.915
cc_469 ( N_GND_c_469_p N_noxref_23_c_7523_n ) capacitor c=0.0013864f \
 //x=72.135 //y=0 //x2=71.955 //y2=0.865
cc_470 ( N_GND_M43_noxref_d N_noxref_23_c_7523_n ) capacitor c=0.00220047f \
 //x=72.03 //y=0.865 //x2=71.955 //y2=0.865
cc_471 ( N_GND_M43_noxref_d N_noxref_23_c_7525_n ) capacitor c=0.00272336f \
 //x=72.03 //y=0.865 //x2=71.955 //y2=1.21
cc_472 ( N_GND_c_22_p N_noxref_23_c_7526_n ) capacitor c=0.00369763f //x=71.04 \
 //y=0 //x2=71.955 //y2=1.915
cc_473 ( N_GND_M43_noxref_d N_noxref_23_c_7527_n ) capacitor c=0.0131326f \
 //x=72.03 //y=0.865 //x2=72.33 //y2=0.71
cc_474 ( N_GND_M43_noxref_d N_noxref_23_c_7528_n ) capacitor c=0.00167494f \
 //x=72.03 //y=0.865 //x2=72.33 //y2=1.365
cc_475 ( N_GND_c_2_p N_noxref_23_c_7529_n ) capacitor c=0.00130622f //x=73.63 \
 //y=0 //x2=72.485 //y2=0.865
cc_476 ( N_GND_M43_noxref_d N_noxref_23_c_7529_n ) capacitor c=0.00257848f \
 //x=72.03 //y=0.865 //x2=72.485 //y2=0.865
cc_477 ( N_GND_M43_noxref_d N_noxref_23_c_7531_n ) capacitor c=0.00272336f \
 //x=72.03 //y=0.865 //x2=72.485 //y2=1.21
cc_478 ( N_GND_c_22_p N_noxref_23_c_7532_n ) capacitor c=0.00662863f //x=71.04 \
 //y=0 //x2=71.78 //y2=2.08
cc_479 ( N_GND_c_7_p N_noxref_23_M12_noxref_d ) capacitor c=8.58106e-19 \
 //x=18.13 //y=0 //x2=20.09 //y2=0.905
cc_480 ( N_GND_c_8_p N_noxref_23_M12_noxref_d ) capacitor c=0.00616547f \
 //x=21.46 //y=0 //x2=20.09 //y2=0.905
cc_481 ( N_GND_M11_noxref_d N_noxref_23_M12_noxref_d ) capacitor c=0.00143464f \
 //x=19.12 //y=0.865 //x2=20.09 //y2=0.905
cc_482 ( N_GND_c_23_p N_QN_c_8045_n ) capacitor c=0.0695894f //x=73.63 //y=0 \
 //x2=69.745 //y2=1.18
cc_483 ( N_GND_c_379_p N_QN_c_8045_n ) capacitor c=0.0081414f //x=67.54 //y=0 \
 //x2=69.745 //y2=1.18
cc_484 ( N_GND_c_382_p N_QN_c_8045_n ) capacitor c=0.0101988f //x=68.805 //y=0 \
 //x2=69.745 //y2=1.18
cc_485 ( N_GND_c_388_p N_QN_c_8045_n ) capacitor c=0.00469062f //x=70.87 //y=0 \
 //x2=69.745 //y2=1.18
cc_486 ( N_GND_c_2_p N_QN_c_8045_n ) capacitor c=0.00132022f //x=73.63 //y=0 \
 //x2=69.745 //y2=1.18
cc_487 ( N_GND_c_21_p N_QN_c_8045_n ) capacitor c=0.0412927f //x=67.71 //y=0 \
 //x2=69.745 //y2=1.18
cc_488 ( N_GND_M41_noxref_d N_QN_c_8045_n ) capacitor c=0.00960943f //x=68.7 \
 //y=0.865 //x2=69.745 //y2=1.18
cc_489 ( N_GND_c_23_p N_QN_c_8052_n ) capacitor c=0.00715563f //x=73.63 //y=0 \
 //x2=66.645 //y2=1.18
cc_490 ( N_GND_c_23_p N_QN_c_8053_n ) capacitor c=0.0769193f //x=73.63 //y=0 \
 //x2=73.075 //y2=1.18
cc_491 ( N_GND_c_388_p N_QN_c_8053_n ) capacitor c=0.00788597f //x=70.87 //y=0 \
 //x2=73.075 //y2=1.18
cc_492 ( N_GND_c_469_p N_QN_c_8053_n ) capacitor c=0.00974891f //x=72.135 \
 //y=0 //x2=73.075 //y2=1.18
cc_493 ( N_GND_c_2_p N_QN_c_8053_n ) capacitor c=0.0057803f //x=73.63 //y=0 \
 //x2=73.075 //y2=1.18
cc_494 ( N_GND_c_22_p N_QN_c_8053_n ) capacitor c=0.0384312f //x=71.04 //y=0 \
 //x2=73.075 //y2=1.18
cc_495 ( N_GND_M43_noxref_d N_QN_c_8053_n ) capacitor c=0.00960943f //x=72.03 \
 //y=0.865 //x2=73.075 //y2=1.18
cc_496 ( N_GND_c_23_p N_QN_c_8059_n ) capacitor c=0.00664346f //x=73.63 //y=0 \
 //x2=69.975 //y2=1.18
cc_497 ( N_GND_c_22_p QN ) capacitor c=0.00109945f //x=71.04 //y=0 //x2=73.63 \
 //y2=2.22
cc_498 ( N_GND_c_2_p N_QN_c_8061_n ) capacitor c=0.04686f //x=73.63 //y=0 \
 //x2=73.545 //y2=1.645
cc_499 ( N_GND_c_23_p N_QN_M40_noxref_d ) capacitor c=2.00936e-19 //x=73.63 \
 //y=0 //x2=66.34 //y2=0.905
cc_500 ( N_GND_c_21_p N_QN_M40_noxref_d ) capacitor c=0.00141366f //x=67.71 \
 //y=0 //x2=66.34 //y2=0.905
cc_501 ( N_GND_M39_noxref_d N_QN_M40_noxref_d ) capacitor c=0.00128667f \
 //x=65.37 //y=0.865 //x2=66.34 //y2=0.905
cc_502 ( N_GND_c_23_p N_QN_M42_noxref_d ) capacitor c=2.00936e-19 //x=73.63 \
 //y=0 //x2=69.67 //y2=0.905
cc_503 ( N_GND_c_22_p N_QN_M42_noxref_d ) capacitor c=0.0014176f //x=71.04 \
 //y=0 //x2=69.67 //y2=0.905
cc_504 ( N_GND_M41_noxref_d N_QN_M42_noxref_d ) capacitor c=0.0012247f \
 //x=68.7 //y=0.865 //x2=69.67 //y2=0.905
cc_505 ( N_GND_c_23_p N_QN_M44_noxref_d ) capacitor c=2.00936e-19 //x=73.63 \
 //y=0 //x2=73 //y2=0.905
cc_506 ( N_GND_c_2_p N_QN_M44_noxref_d ) capacitor c=0.00524992f //x=73.63 \
 //y=0 //x2=73 //y2=0.905
cc_507 ( N_GND_c_22_p N_QN_M44_noxref_d ) capacitor c=8.62423e-19 //x=71.04 \
 //y=0 //x2=73 //y2=0.905
cc_508 ( N_GND_M43_noxref_d N_QN_M44_noxref_d ) capacitor c=0.0012247f \
 //x=72.03 //y=0.865 //x2=73 //y2=0.905
cc_509 ( N_GND_c_23_p N_noxref_26_c_8214_n ) capacitor c=0.00618812f //x=73.63 \
 //y=0 //x2=1.475 //y2=1.59
cc_510 ( N_GND_c_113_p N_noxref_26_c_8214_n ) capacitor c=0.00110021f //x=0.99 \
 //y=0 //x2=1.475 //y2=1.59
cc_511 ( N_GND_c_24_p N_noxref_26_c_8214_n ) capacitor c=0.00179185f //x=4.64 \
 //y=0 //x2=1.475 //y2=1.59
cc_512 ( N_GND_M0_noxref_d N_noxref_26_c_8214_n ) capacitor c=0.00894788f \
 //x=0.885 //y=0.875 //x2=1.475 //y2=1.59
cc_513 ( N_GND_c_23_p N_noxref_26_c_8218_n ) capacitor c=0.00575184f //x=73.63 \
 //y=0 //x2=1.56 //y2=0.625
cc_514 ( N_GND_c_24_p N_noxref_26_c_8218_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=1.56 //y2=0.625
cc_515 ( N_GND_M0_noxref_d N_noxref_26_c_8218_n ) capacitor c=0.033954f \
 //x=0.885 //y=0.875 //x2=1.56 //y2=0.625
cc_516 ( N_GND_c_23_p N_noxref_26_c_8221_n ) capacitor c=0.0139021f //x=73.63 \
 //y=0 //x2=2.445 //y2=0.54
cc_517 ( N_GND_c_24_p N_noxref_26_c_8221_n ) capacitor c=0.0356078f //x=4.64 \
 //y=0 //x2=2.445 //y2=0.54
cc_518 ( N_GND_c_2_p N_noxref_26_c_8221_n ) capacitor c=0.00178035f //x=73.63 \
 //y=0 //x2=2.445 //y2=0.54
cc_519 ( N_GND_c_23_p N_noxref_26_M0_noxref_s ) capacitor c=0.0125336f \
 //x=73.63 //y=0 //x2=0.455 //y2=0.375
cc_520 ( N_GND_c_113_p N_noxref_26_M0_noxref_s ) capacitor c=0.0140218f \
 //x=0.99 //y=0 //x2=0.455 //y2=0.375
cc_521 ( N_GND_c_1_p N_noxref_26_M0_noxref_s ) capacitor c=0.0712607f //x=0.74 \
 //y=0 //x2=0.455 //y2=0.375
cc_522 ( N_GND_c_24_p N_noxref_26_M0_noxref_s ) capacitor c=0.0131422f \
 //x=4.64 //y=0 //x2=0.455 //y2=0.375
cc_523 ( N_GND_c_3_p N_noxref_26_M0_noxref_s ) capacitor c=3.31601e-19 \
 //x=4.81 //y=0 //x2=0.455 //y2=0.375
cc_524 ( N_GND_M0_noxref_d N_noxref_26_M0_noxref_s ) capacitor c=0.033718f \
 //x=0.885 //y=0.875 //x2=0.455 //y2=0.375
cc_525 ( N_GND_c_23_p N_noxref_27_c_8261_n ) capacitor c=0.00402784f //x=73.63 \
 //y=0 //x2=3.015 //y2=0.995
cc_526 ( N_GND_c_24_p N_noxref_27_c_8261_n ) capacitor c=0.00829979f //x=4.64 \
 //y=0 //x2=3.015 //y2=0.995
cc_527 ( N_GND_c_23_p N_noxref_27_c_8263_n ) capacitor c=0.00575184f //x=73.63 \
 //y=0 //x2=3.1 //y2=0.625
cc_528 ( N_GND_c_24_p N_noxref_27_c_8263_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=3.1 //y2=0.625
cc_529 ( N_GND_M0_noxref_d N_noxref_27_c_8263_n ) capacitor c=6.21394e-19 \
 //x=0.885 //y=0.875 //x2=3.1 //y2=0.625
cc_530 ( N_GND_c_23_p N_noxref_27_c_8266_n ) capacitor c=0.0118365f //x=73.63 \
 //y=0 //x2=3.985 //y2=0.54
cc_531 ( N_GND_c_24_p N_noxref_27_c_8266_n ) capacitor c=0.0365413f //x=4.64 \
 //y=0 //x2=3.985 //y2=0.54
cc_532 ( N_GND_c_2_p N_noxref_27_c_8266_n ) capacitor c=0.00190179f //x=73.63 \
 //y=0 //x2=3.985 //y2=0.54
cc_533 ( N_GND_c_23_p N_noxref_27_c_8269_n ) capacitor c=0.00287549f //x=73.63 \
 //y=0 //x2=4.07 //y2=0.625
cc_534 ( N_GND_c_24_p N_noxref_27_c_8269_n ) capacitor c=0.0142658f //x=4.64 \
 //y=0 //x2=4.07 //y2=0.625
cc_535 ( N_GND_c_3_p N_noxref_27_c_8269_n ) capacitor c=0.0404137f //x=4.81 \
 //y=0 //x2=4.07 //y2=0.625
cc_536 ( N_GND_M0_noxref_d N_noxref_27_M1_noxref_d ) capacitor c=0.00162435f \
 //x=0.885 //y=0.875 //x2=1.86 //y2=0.91
cc_537 ( N_GND_c_1_p N_noxref_27_M2_noxref_s ) capacitor c=8.16352e-19 \
 //x=0.74 //y=0 //x2=2.965 //y2=0.375
cc_538 ( N_GND_c_3_p N_noxref_27_M2_noxref_s ) capacitor c=0.00183576f \
 //x=4.81 //y=0 //x2=2.965 //y2=0.375
cc_539 ( N_GND_c_23_p N_noxref_28_c_8314_n ) capacitor c=0.00552526f //x=73.63 \
 //y=0 //x2=6.39 //y2=1.58
cc_540 ( N_GND_c_25_p N_noxref_28_c_8314_n ) capacitor c=0.00113001f //x=5.905 \
 //y=0 //x2=6.39 //y2=1.58
cc_541 ( N_GND_c_74_p N_noxref_28_c_8314_n ) capacitor c=0.0018242f //x=7.97 \
 //y=0 //x2=6.39 //y2=1.58
cc_542 ( N_GND_M3_noxref_d N_noxref_28_c_8314_n ) capacitor c=0.00897209f \
 //x=5.8 //y=0.865 //x2=6.39 //y2=1.58
cc_543 ( N_GND_c_23_p N_noxref_28_c_8318_n ) capacitor c=0.00287501f //x=73.63 \
 //y=0 //x2=6.475 //y2=0.615
cc_544 ( N_GND_c_74_p N_noxref_28_c_8318_n ) capacitor c=0.014584f //x=7.97 \
 //y=0 //x2=6.475 //y2=0.615
cc_545 ( N_GND_M3_noxref_d N_noxref_28_c_8318_n ) capacitor c=0.033812f \
 //x=5.8 //y=0.865 //x2=6.475 //y2=0.615
cc_546 ( N_GND_c_3_p N_noxref_28_c_8321_n ) capacitor c=2.91423e-19 //x=4.81 \
 //y=0 //x2=6.475 //y2=1.495
cc_547 ( N_GND_c_23_p N_noxref_28_c_8322_n ) capacitor c=0.0111758f //x=73.63 \
 //y=0 //x2=7.36 //y2=0.53
cc_548 ( N_GND_c_74_p N_noxref_28_c_8322_n ) capacitor c=0.0374722f //x=7.97 \
 //y=0 //x2=7.36 //y2=0.53
cc_549 ( N_GND_c_2_p N_noxref_28_c_8322_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=7.36 //y2=0.53
cc_550 ( N_GND_c_23_p N_noxref_28_c_8325_n ) capacitor c=0.00271457f //x=73.63 \
 //y=0 //x2=7.445 //y2=0.615
cc_551 ( N_GND_c_74_p N_noxref_28_c_8325_n ) capacitor c=0.0147189f //x=7.97 \
 //y=0 //x2=7.445 //y2=0.615
cc_552 ( N_GND_c_4_p N_noxref_28_c_8325_n ) capacitor c=0.0431718f //x=8.14 \
 //y=0 //x2=7.445 //y2=0.615
cc_553 ( N_GND_c_23_p N_noxref_28_M3_noxref_s ) capacitor c=0.00293348f \
 //x=73.63 //y=0 //x2=5.37 //y2=0.365
cc_554 ( N_GND_c_25_p N_noxref_28_M3_noxref_s ) capacitor c=0.0149357f \
 //x=5.905 //y=0 //x2=5.37 //y2=0.365
cc_555 ( N_GND_c_3_p N_noxref_28_M3_noxref_s ) capacitor c=0.0583534f //x=4.81 \
 //y=0 //x2=5.37 //y2=0.365
cc_556 ( N_GND_c_4_p N_noxref_28_M3_noxref_s ) capacitor c=0.00198043f \
 //x=8.14 //y=0 //x2=5.37 //y2=0.365
cc_557 ( N_GND_M3_noxref_d N_noxref_28_M3_noxref_s ) capacitor c=0.0334197f \
 //x=5.8 //y=0.865 //x2=5.37 //y2=0.365
cc_558 ( N_GND_c_23_p N_noxref_29_c_8368_n ) capacitor c=0.00530453f //x=73.63 \
 //y=0 //x2=9.72 //y2=1.58
cc_559 ( N_GND_c_33_p N_noxref_29_c_8368_n ) capacitor c=0.00112921f //x=9.235 \
 //y=0 //x2=9.72 //y2=1.58
cc_560 ( N_GND_c_40_p N_noxref_29_c_8368_n ) capacitor c=0.00182339f //x=11.3 \
 //y=0 //x2=9.72 //y2=1.58
cc_561 ( N_GND_M5_noxref_d N_noxref_29_c_8368_n ) capacitor c=0.00879185f \
 //x=9.13 //y=0.865 //x2=9.72 //y2=1.58
cc_562 ( N_GND_c_23_p N_noxref_29_c_8372_n ) capacitor c=0.00271584f //x=73.63 \
 //y=0 //x2=9.805 //y2=0.615
cc_563 ( N_GND_c_40_p N_noxref_29_c_8372_n ) capacitor c=0.014783f //x=11.3 \
 //y=0 //x2=9.805 //y2=0.615
cc_564 ( N_GND_M5_noxref_d N_noxref_29_c_8372_n ) capacitor c=0.033812f \
 //x=9.13 //y=0.865 //x2=9.805 //y2=0.615
cc_565 ( N_GND_c_4_p N_noxref_29_c_8375_n ) capacitor c=2.91423e-19 //x=8.14 \
 //y=0 //x2=9.805 //y2=1.495
cc_566 ( N_GND_c_23_p N_noxref_29_c_8376_n ) capacitor c=0.0111861f //x=73.63 \
 //y=0 //x2=10.69 //y2=0.53
cc_567 ( N_GND_c_40_p N_noxref_29_c_8376_n ) capacitor c=0.0374741f //x=11.3 \
 //y=0 //x2=10.69 //y2=0.53
cc_568 ( N_GND_c_2_p N_noxref_29_c_8376_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=10.69 //y2=0.53
cc_569 ( N_GND_c_23_p N_noxref_29_c_8379_n ) capacitor c=0.00271457f //x=73.63 \
 //y=0 //x2=10.775 //y2=0.615
cc_570 ( N_GND_c_40_p N_noxref_29_c_8379_n ) capacitor c=0.0147189f //x=11.3 \
 //y=0 //x2=10.775 //y2=0.615
cc_571 ( N_GND_c_5_p N_noxref_29_c_8379_n ) capacitor c=0.0431718f //x=11.47 \
 //y=0 //x2=10.775 //y2=0.615
cc_572 ( N_GND_c_23_p N_noxref_29_M5_noxref_s ) capacitor c=0.00271584f \
 //x=73.63 //y=0 //x2=8.7 //y2=0.365
cc_573 ( N_GND_c_33_p N_noxref_29_M5_noxref_s ) capacitor c=0.014783f \
 //x=9.235 //y=0 //x2=8.7 //y2=0.365
cc_574 ( N_GND_c_4_p N_noxref_29_M5_noxref_s ) capacitor c=0.058339f //x=8.14 \
 //y=0 //x2=8.7 //y2=0.365
cc_575 ( N_GND_c_5_p N_noxref_29_M5_noxref_s ) capacitor c=0.00198043f \
 //x=11.47 //y=0 //x2=8.7 //y2=0.365
cc_576 ( N_GND_M5_noxref_d N_noxref_29_M5_noxref_s ) capacitor c=0.0334197f \
 //x=9.13 //y=0.865 //x2=8.7 //y2=0.365
cc_577 ( N_GND_c_23_p N_noxref_30_c_8420_n ) capacitor c=0.00530453f //x=73.63 \
 //y=0 //x2=13.05 //y2=1.58
cc_578 ( N_GND_c_50_p N_noxref_30_c_8420_n ) capacitor c=0.00112921f \
 //x=12.565 //y=0 //x2=13.05 //y2=1.58
cc_579 ( N_GND_c_57_p N_noxref_30_c_8420_n ) capacitor c=0.00182339f //x=14.63 \
 //y=0 //x2=13.05 //y2=1.58
cc_580 ( N_GND_M7_noxref_d N_noxref_30_c_8420_n ) capacitor c=0.00879185f \
 //x=12.46 //y=0.865 //x2=13.05 //y2=1.58
cc_581 ( N_GND_c_23_p N_noxref_30_c_8424_n ) capacitor c=0.00271584f //x=73.63 \
 //y=0 //x2=13.135 //y2=0.615
cc_582 ( N_GND_c_57_p N_noxref_30_c_8424_n ) capacitor c=0.014783f //x=14.63 \
 //y=0 //x2=13.135 //y2=0.615
cc_583 ( N_GND_M7_noxref_d N_noxref_30_c_8424_n ) capacitor c=0.033812f \
 //x=12.46 //y=0.865 //x2=13.135 //y2=0.615
cc_584 ( N_GND_c_5_p N_noxref_30_c_8427_n ) capacitor c=2.91423e-19 //x=11.47 \
 //y=0 //x2=13.135 //y2=1.495
cc_585 ( N_GND_c_23_p N_noxref_30_c_8428_n ) capacitor c=0.0111861f //x=73.63 \
 //y=0 //x2=14.02 //y2=0.53
cc_586 ( N_GND_c_57_p N_noxref_30_c_8428_n ) capacitor c=0.0374741f //x=14.63 \
 //y=0 //x2=14.02 //y2=0.53
cc_587 ( N_GND_c_2_p N_noxref_30_c_8428_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=14.02 //y2=0.53
cc_588 ( N_GND_c_23_p N_noxref_30_c_8431_n ) capacitor c=0.00271457f //x=73.63 \
 //y=0 //x2=14.105 //y2=0.615
cc_589 ( N_GND_c_57_p N_noxref_30_c_8431_n ) capacitor c=0.0147189f //x=14.63 \
 //y=0 //x2=14.105 //y2=0.615
cc_590 ( N_GND_c_6_p N_noxref_30_c_8431_n ) capacitor c=0.0431718f //x=14.8 \
 //y=0 //x2=14.105 //y2=0.615
cc_591 ( N_GND_c_23_p N_noxref_30_M7_noxref_s ) capacitor c=0.00271584f \
 //x=73.63 //y=0 //x2=12.03 //y2=0.365
cc_592 ( N_GND_c_50_p N_noxref_30_M7_noxref_s ) capacitor c=0.014783f \
 //x=12.565 //y=0 //x2=12.03 //y2=0.365
cc_593 ( N_GND_c_5_p N_noxref_30_M7_noxref_s ) capacitor c=0.058339f //x=11.47 \
 //y=0 //x2=12.03 //y2=0.365
cc_594 ( N_GND_c_6_p N_noxref_30_M7_noxref_s ) capacitor c=0.00198043f \
 //x=14.8 //y=0 //x2=12.03 //y2=0.365
cc_595 ( N_GND_M7_noxref_d N_noxref_30_M7_noxref_s ) capacitor c=0.0334197f \
 //x=12.46 //y=0.865 //x2=12.03 //y2=0.365
cc_596 ( N_GND_c_23_p N_noxref_31_c_8472_n ) capacitor c=0.00530453f //x=73.63 \
 //y=0 //x2=16.38 //y2=1.58
cc_597 ( N_GND_c_77_p N_noxref_31_c_8472_n ) capacitor c=0.00112921f \
 //x=15.895 //y=0 //x2=16.38 //y2=1.58
cc_598 ( N_GND_c_84_p N_noxref_31_c_8472_n ) capacitor c=0.00182339f //x=17.96 \
 //y=0 //x2=16.38 //y2=1.58
cc_599 ( N_GND_M9_noxref_d N_noxref_31_c_8472_n ) capacitor c=0.00879185f \
 //x=15.79 //y=0.865 //x2=16.38 //y2=1.58
cc_600 ( N_GND_c_23_p N_noxref_31_c_8476_n ) capacitor c=0.00271584f //x=73.63 \
 //y=0 //x2=16.465 //y2=0.615
cc_601 ( N_GND_c_84_p N_noxref_31_c_8476_n ) capacitor c=0.014783f //x=17.96 \
 //y=0 //x2=16.465 //y2=0.615
cc_602 ( N_GND_M9_noxref_d N_noxref_31_c_8476_n ) capacitor c=0.033812f \
 //x=15.79 //y=0.865 //x2=16.465 //y2=0.615
cc_603 ( N_GND_c_6_p N_noxref_31_c_8479_n ) capacitor c=2.91423e-19 //x=14.8 \
 //y=0 //x2=16.465 //y2=1.495
cc_604 ( N_GND_c_23_p N_noxref_31_c_8480_n ) capacitor c=0.0111861f //x=73.63 \
 //y=0 //x2=17.35 //y2=0.53
cc_605 ( N_GND_c_84_p N_noxref_31_c_8480_n ) capacitor c=0.0374741f //x=17.96 \
 //y=0 //x2=17.35 //y2=0.53
cc_606 ( N_GND_c_2_p N_noxref_31_c_8480_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=17.35 //y2=0.53
cc_607 ( N_GND_c_23_p N_noxref_31_c_8483_n ) capacitor c=0.00271457f //x=73.63 \
 //y=0 //x2=17.435 //y2=0.615
cc_608 ( N_GND_c_84_p N_noxref_31_c_8483_n ) capacitor c=0.0147189f //x=17.96 \
 //y=0 //x2=17.435 //y2=0.615
cc_609 ( N_GND_c_7_p N_noxref_31_c_8483_n ) capacitor c=0.0431718f //x=18.13 \
 //y=0 //x2=17.435 //y2=0.615
cc_610 ( N_GND_c_23_p N_noxref_31_M9_noxref_s ) capacitor c=0.00271584f \
 //x=73.63 //y=0 //x2=15.36 //y2=0.365
cc_611 ( N_GND_c_77_p N_noxref_31_M9_noxref_s ) capacitor c=0.014783f \
 //x=15.895 //y=0 //x2=15.36 //y2=0.365
cc_612 ( N_GND_c_6_p N_noxref_31_M9_noxref_s ) capacitor c=0.058339f //x=14.8 \
 //y=0 //x2=15.36 //y2=0.365
cc_613 ( N_GND_c_7_p N_noxref_31_M9_noxref_s ) capacitor c=0.00198043f \
 //x=18.13 //y=0 //x2=15.36 //y2=0.365
cc_614 ( N_GND_M9_noxref_d N_noxref_31_M9_noxref_s ) capacitor c=0.0334197f \
 //x=15.79 //y=0.865 //x2=15.36 //y2=0.365
cc_615 ( N_GND_c_23_p N_noxref_32_c_8524_n ) capacitor c=0.00530453f //x=73.63 \
 //y=0 //x2=19.71 //y2=1.58
cc_616 ( N_GND_c_91_p N_noxref_32_c_8524_n ) capacitor c=0.00112921f \
 //x=19.225 //y=0 //x2=19.71 //y2=1.58
cc_617 ( N_GND_c_98_p N_noxref_32_c_8524_n ) capacitor c=0.00182339f //x=21.29 \
 //y=0 //x2=19.71 //y2=1.58
cc_618 ( N_GND_M11_noxref_d N_noxref_32_c_8524_n ) capacitor c=0.00879185f \
 //x=19.12 //y=0.865 //x2=19.71 //y2=1.58
cc_619 ( N_GND_c_23_p N_noxref_32_c_8528_n ) capacitor c=0.00271584f //x=73.63 \
 //y=0 //x2=19.795 //y2=0.615
cc_620 ( N_GND_c_98_p N_noxref_32_c_8528_n ) capacitor c=0.014783f //x=21.29 \
 //y=0 //x2=19.795 //y2=0.615
cc_621 ( N_GND_M11_noxref_d N_noxref_32_c_8528_n ) capacitor c=0.033812f \
 //x=19.12 //y=0.865 //x2=19.795 //y2=0.615
cc_622 ( N_GND_c_7_p N_noxref_32_c_8531_n ) capacitor c=2.91423e-19 //x=18.13 \
 //y=0 //x2=19.795 //y2=1.495
cc_623 ( N_GND_c_23_p N_noxref_32_c_8532_n ) capacitor c=0.0111861f //x=73.63 \
 //y=0 //x2=20.68 //y2=0.53
cc_624 ( N_GND_c_98_p N_noxref_32_c_8532_n ) capacitor c=0.0374741f //x=21.29 \
 //y=0 //x2=20.68 //y2=0.53
cc_625 ( N_GND_c_2_p N_noxref_32_c_8532_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=20.68 //y2=0.53
cc_626 ( N_GND_c_23_p N_noxref_32_c_8535_n ) capacitor c=0.00271457f //x=73.63 \
 //y=0 //x2=20.765 //y2=0.615
cc_627 ( N_GND_c_98_p N_noxref_32_c_8535_n ) capacitor c=0.0147189f //x=21.29 \
 //y=0 //x2=20.765 //y2=0.615
cc_628 ( N_GND_c_8_p N_noxref_32_c_8535_n ) capacitor c=0.0431718f //x=21.46 \
 //y=0 //x2=20.765 //y2=0.615
cc_629 ( N_GND_c_23_p N_noxref_32_M11_noxref_s ) capacitor c=0.00271584f \
 //x=73.63 //y=0 //x2=18.69 //y2=0.365
cc_630 ( N_GND_c_91_p N_noxref_32_M11_noxref_s ) capacitor c=0.014783f \
 //x=19.225 //y=0 //x2=18.69 //y2=0.365
cc_631 ( N_GND_c_7_p N_noxref_32_M11_noxref_s ) capacitor c=0.058339f \
 //x=18.13 //y=0 //x2=18.69 //y2=0.365
cc_632 ( N_GND_c_8_p N_noxref_32_M11_noxref_s ) capacitor c=0.00198098f \
 //x=21.46 //y=0 //x2=18.69 //y2=0.365
cc_633 ( N_GND_M11_noxref_d N_noxref_32_M11_noxref_s ) capacitor c=0.0334197f \
 //x=19.12 //y=0.865 //x2=18.69 //y2=0.365
cc_634 ( N_GND_c_23_p N_noxref_33_c_8576_n ) capacitor c=0.00529827f //x=73.63 \
 //y=0 //x2=22.935 //y2=1.59
cc_635 ( N_GND_c_206_p N_noxref_33_c_8576_n ) capacitor c=0.00111496f \
 //x=22.45 //y=0 //x2=22.935 //y2=1.59
cc_636 ( N_GND_c_213_p N_noxref_33_c_8576_n ) capacitor c=0.0018066f //x=26.1 \
 //y=0 //x2=22.935 //y2=1.59
cc_637 ( N_GND_M13_noxref_d N_noxref_33_c_8576_n ) capacitor c=0.00869643f \
 //x=22.345 //y=0.875 //x2=22.935 //y2=1.59
cc_638 ( N_GND_c_23_p N_noxref_33_c_8580_n ) capacitor c=0.00266608f //x=73.63 \
 //y=0 //x2=23.02 //y2=0.625
cc_639 ( N_GND_c_213_p N_noxref_33_c_8580_n ) capacitor c=0.0141814f //x=26.1 \
 //y=0 //x2=23.02 //y2=0.625
cc_640 ( N_GND_M13_noxref_d N_noxref_33_c_8580_n ) capacitor c=0.033954f \
 //x=22.345 //y=0.875 //x2=23.02 //y2=0.625
cc_641 ( N_GND_c_23_p N_noxref_33_c_8583_n ) capacitor c=0.0109327f //x=73.63 \
 //y=0 //x2=23.905 //y2=0.54
cc_642 ( N_GND_c_213_p N_noxref_33_c_8583_n ) capacitor c=0.0361235f //x=26.1 \
 //y=0 //x2=23.905 //y2=0.54
cc_643 ( N_GND_c_2_p N_noxref_33_c_8583_n ) capacitor c=0.00178035f //x=73.63 \
 //y=0 //x2=23.905 //y2=0.54
cc_644 ( N_GND_c_23_p N_noxref_33_M13_noxref_s ) capacitor c=0.00532331f \
 //x=73.63 //y=0 //x2=21.915 //y2=0.375
cc_645 ( N_GND_c_206_p N_noxref_33_M13_noxref_s ) capacitor c=0.0141814f \
 //x=22.45 //y=0 //x2=21.915 //y2=0.375
cc_646 ( N_GND_c_213_p N_noxref_33_M13_noxref_s ) capacitor c=0.0132355f \
 //x=26.1 //y=0 //x2=21.915 //y2=0.375
cc_647 ( N_GND_c_8_p N_noxref_33_M13_noxref_s ) capacitor c=0.0696963f \
 //x=21.46 //y=0 //x2=21.915 //y2=0.375
cc_648 ( N_GND_c_9_p N_noxref_33_M13_noxref_s ) capacitor c=3.31601e-19 \
 //x=26.27 //y=0 //x2=21.915 //y2=0.375
cc_649 ( N_GND_M13_noxref_d N_noxref_33_M13_noxref_s ) capacitor c=0.033718f \
 //x=22.345 //y=0.875 //x2=21.915 //y2=0.375
cc_650 ( N_GND_c_23_p N_noxref_34_c_8626_n ) capacitor c=0.00364762f //x=73.63 \
 //y=0 //x2=24.475 //y2=0.995
cc_651 ( N_GND_c_213_p N_noxref_34_c_8626_n ) capacitor c=0.00940048f //x=26.1 \
 //y=0 //x2=24.475 //y2=0.995
cc_652 ( N_GND_c_23_p N_noxref_34_c_8628_n ) capacitor c=0.00266608f //x=73.63 \
 //y=0 //x2=24.56 //y2=0.625
cc_653 ( N_GND_c_213_p N_noxref_34_c_8628_n ) capacitor c=0.0141814f //x=26.1 \
 //y=0 //x2=24.56 //y2=0.625
cc_654 ( N_GND_M13_noxref_d N_noxref_34_c_8628_n ) capacitor c=6.21394e-19 \
 //x=22.345 //y=0.875 //x2=24.56 //y2=0.625
cc_655 ( N_GND_c_23_p N_noxref_34_c_8631_n ) capacitor c=0.0110123f //x=73.63 \
 //y=0 //x2=25.445 //y2=0.54
cc_656 ( N_GND_c_213_p N_noxref_34_c_8631_n ) capacitor c=0.0364631f //x=26.1 \
 //y=0 //x2=25.445 //y2=0.54
cc_657 ( N_GND_c_2_p N_noxref_34_c_8631_n ) capacitor c=0.00190179f //x=73.63 \
 //y=0 //x2=25.445 //y2=0.54
cc_658 ( N_GND_c_23_p N_noxref_34_c_8634_n ) capacitor c=0.00266421f //x=73.63 \
 //y=0 //x2=25.53 //y2=0.625
cc_659 ( N_GND_c_213_p N_noxref_34_c_8634_n ) capacitor c=0.0141195f //x=26.1 \
 //y=0 //x2=25.53 //y2=0.625
cc_660 ( N_GND_c_9_p N_noxref_34_c_8634_n ) capacitor c=0.0404137f //x=26.27 \
 //y=0 //x2=25.53 //y2=0.625
cc_661 ( N_GND_M13_noxref_d N_noxref_34_M14_noxref_d ) capacitor c=0.00162435f \
 //x=22.345 //y=0.875 //x2=23.32 //y2=0.91
cc_662 ( N_GND_c_8_p N_noxref_34_M15_noxref_s ) capacitor c=8.16352e-19 \
 //x=21.46 //y=0 //x2=24.425 //y2=0.375
cc_663 ( N_GND_c_9_p N_noxref_34_M15_noxref_s ) capacitor c=0.00183576f \
 //x=26.27 //y=0 //x2=24.425 //y2=0.375
cc_664 ( N_GND_c_23_p N_noxref_35_c_8679_n ) capacitor c=0.00530453f //x=73.63 \
 //y=0 //x2=27.85 //y2=1.58
cc_665 ( N_GND_c_162_p N_noxref_35_c_8679_n ) capacitor c=0.00112921f \
 //x=27.365 //y=0 //x2=27.85 //y2=1.58
cc_666 ( N_GND_c_169_p N_noxref_35_c_8679_n ) capacitor c=0.00182339f \
 //x=29.43 //y=0 //x2=27.85 //y2=1.58
cc_667 ( N_GND_M16_noxref_d N_noxref_35_c_8679_n ) capacitor c=0.00879185f \
 //x=27.26 //y=0.865 //x2=27.85 //y2=1.58
cc_668 ( N_GND_c_23_p N_noxref_35_c_8683_n ) capacitor c=0.00271498f //x=73.63 \
 //y=0 //x2=27.935 //y2=0.615
cc_669 ( N_GND_c_169_p N_noxref_35_c_8683_n ) capacitor c=0.0147824f //x=29.43 \
 //y=0 //x2=27.935 //y2=0.615
cc_670 ( N_GND_M16_noxref_d N_noxref_35_c_8683_n ) capacitor c=0.033812f \
 //x=27.26 //y=0.865 //x2=27.935 //y2=0.615
cc_671 ( N_GND_c_9_p N_noxref_35_c_8686_n ) capacitor c=2.91423e-19 //x=26.27 \
 //y=0 //x2=27.935 //y2=1.495
cc_672 ( N_GND_c_23_p N_noxref_35_c_8687_n ) capacitor c=0.0111758f //x=73.63 \
 //y=0 //x2=28.82 //y2=0.53
cc_673 ( N_GND_c_169_p N_noxref_35_c_8687_n ) capacitor c=0.0374722f //x=29.43 \
 //y=0 //x2=28.82 //y2=0.53
cc_674 ( N_GND_c_2_p N_noxref_35_c_8687_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=28.82 //y2=0.53
cc_675 ( N_GND_c_23_p N_noxref_35_c_8690_n ) capacitor c=0.00271457f //x=73.63 \
 //y=0 //x2=28.905 //y2=0.615
cc_676 ( N_GND_c_169_p N_noxref_35_c_8690_n ) capacitor c=0.0147189f //x=29.43 \
 //y=0 //x2=28.905 //y2=0.615
cc_677 ( N_GND_c_10_p N_noxref_35_c_8690_n ) capacitor c=0.0431718f //x=29.6 \
 //y=0 //x2=28.905 //y2=0.615
cc_678 ( N_GND_c_23_p N_noxref_35_M16_noxref_s ) capacitor c=0.00271584f \
 //x=73.63 //y=0 //x2=26.83 //y2=0.365
cc_679 ( N_GND_c_162_p N_noxref_35_M16_noxref_s ) capacitor c=0.014783f \
 //x=27.365 //y=0 //x2=26.83 //y2=0.365
cc_680 ( N_GND_c_9_p N_noxref_35_M16_noxref_s ) capacitor c=0.0583534f \
 //x=26.27 //y=0 //x2=26.83 //y2=0.365
cc_681 ( N_GND_c_10_p N_noxref_35_M16_noxref_s ) capacitor c=0.00198043f \
 //x=29.6 //y=0 //x2=26.83 //y2=0.365
cc_682 ( N_GND_M16_noxref_d N_noxref_35_M16_noxref_s ) capacitor c=0.0334197f \
 //x=27.26 //y=0.865 //x2=26.83 //y2=0.365
cc_683 ( N_GND_c_23_p N_noxref_36_c_8733_n ) capacitor c=0.00530453f //x=73.63 \
 //y=0 //x2=31.18 //y2=1.58
cc_684 ( N_GND_c_130_p N_noxref_36_c_8733_n ) capacitor c=0.00112921f \
 //x=30.695 //y=0 //x2=31.18 //y2=1.58
cc_685 ( N_GND_c_137_p N_noxref_36_c_8733_n ) capacitor c=0.00182339f \
 //x=32.76 //y=0 //x2=31.18 //y2=1.58
cc_686 ( N_GND_M18_noxref_d N_noxref_36_c_8733_n ) capacitor c=0.00879185f \
 //x=30.59 //y=0.865 //x2=31.18 //y2=1.58
cc_687 ( N_GND_c_23_p N_noxref_36_c_8737_n ) capacitor c=0.00271584f //x=73.63 \
 //y=0 //x2=31.265 //y2=0.615
cc_688 ( N_GND_c_137_p N_noxref_36_c_8737_n ) capacitor c=0.014783f //x=32.76 \
 //y=0 //x2=31.265 //y2=0.615
cc_689 ( N_GND_M18_noxref_d N_noxref_36_c_8737_n ) capacitor c=0.033812f \
 //x=30.59 //y=0.865 //x2=31.265 //y2=0.615
cc_690 ( N_GND_c_10_p N_noxref_36_c_8740_n ) capacitor c=2.91423e-19 //x=29.6 \
 //y=0 //x2=31.265 //y2=1.495
cc_691 ( N_GND_c_23_p N_noxref_36_c_8741_n ) capacitor c=0.0111861f //x=73.63 \
 //y=0 //x2=32.15 //y2=0.53
cc_692 ( N_GND_c_137_p N_noxref_36_c_8741_n ) capacitor c=0.0374741f //x=32.76 \
 //y=0 //x2=32.15 //y2=0.53
cc_693 ( N_GND_c_2_p N_noxref_36_c_8741_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=32.15 //y2=0.53
cc_694 ( N_GND_c_23_p N_noxref_36_c_8744_n ) capacitor c=0.00271457f //x=73.63 \
 //y=0 //x2=32.235 //y2=0.615
cc_695 ( N_GND_c_137_p N_noxref_36_c_8744_n ) capacitor c=0.0147189f //x=32.76 \
 //y=0 //x2=32.235 //y2=0.615
cc_696 ( N_GND_c_11_p N_noxref_36_c_8744_n ) capacitor c=0.0431718f //x=32.93 \
 //y=0 //x2=32.235 //y2=0.615
cc_697 ( N_GND_c_23_p N_noxref_36_M18_noxref_s ) capacitor c=0.00271584f \
 //x=73.63 //y=0 //x2=30.16 //y2=0.365
cc_698 ( N_GND_c_130_p N_noxref_36_M18_noxref_s ) capacitor c=0.014783f \
 //x=30.695 //y=0 //x2=30.16 //y2=0.365
cc_699 ( N_GND_c_10_p N_noxref_36_M18_noxref_s ) capacitor c=0.058339f \
 //x=29.6 //y=0 //x2=30.16 //y2=0.365
cc_700 ( N_GND_c_11_p N_noxref_36_M18_noxref_s ) capacitor c=0.00198043f \
 //x=32.93 //y=0 //x2=30.16 //y2=0.365
cc_701 ( N_GND_M18_noxref_d N_noxref_36_M18_noxref_s ) capacitor c=0.0334197f \
 //x=30.59 //y=0.865 //x2=30.16 //y2=0.365
cc_702 ( N_GND_c_23_p N_noxref_37_c_8785_n ) capacitor c=0.00530453f //x=73.63 \
 //y=0 //x2=34.51 //y2=1.58
cc_703 ( N_GND_c_146_p N_noxref_37_c_8785_n ) capacitor c=0.00112921f \
 //x=34.025 //y=0 //x2=34.51 //y2=1.58
cc_704 ( N_GND_c_153_p N_noxref_37_c_8785_n ) capacitor c=0.00182339f \
 //x=36.09 //y=0 //x2=34.51 //y2=1.58
cc_705 ( N_GND_M20_noxref_d N_noxref_37_c_8785_n ) capacitor c=0.00879185f \
 //x=33.92 //y=0.865 //x2=34.51 //y2=1.58
cc_706 ( N_GND_c_23_p N_noxref_37_c_8789_n ) capacitor c=0.00271584f //x=73.63 \
 //y=0 //x2=34.595 //y2=0.615
cc_707 ( N_GND_c_153_p N_noxref_37_c_8789_n ) capacitor c=0.014783f //x=36.09 \
 //y=0 //x2=34.595 //y2=0.615
cc_708 ( N_GND_M20_noxref_d N_noxref_37_c_8789_n ) capacitor c=0.033812f \
 //x=33.92 //y=0.865 //x2=34.595 //y2=0.615
cc_709 ( N_GND_c_11_p N_noxref_37_c_8792_n ) capacitor c=2.91423e-19 //x=32.93 \
 //y=0 //x2=34.595 //y2=1.495
cc_710 ( N_GND_c_23_p N_noxref_37_c_8793_n ) capacitor c=0.0111861f //x=73.63 \
 //y=0 //x2=35.48 //y2=0.53
cc_711 ( N_GND_c_153_p N_noxref_37_c_8793_n ) capacitor c=0.0374741f //x=36.09 \
 //y=0 //x2=35.48 //y2=0.53
cc_712 ( N_GND_c_2_p N_noxref_37_c_8793_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=35.48 //y2=0.53
cc_713 ( N_GND_c_23_p N_noxref_37_c_8796_n ) capacitor c=0.00271457f //x=73.63 \
 //y=0 //x2=35.565 //y2=0.615
cc_714 ( N_GND_c_153_p N_noxref_37_c_8796_n ) capacitor c=0.0147189f //x=36.09 \
 //y=0 //x2=35.565 //y2=0.615
cc_715 ( N_GND_c_12_p N_noxref_37_c_8796_n ) capacitor c=0.0431718f //x=36.26 \
 //y=0 //x2=35.565 //y2=0.615
cc_716 ( N_GND_c_23_p N_noxref_37_M20_noxref_s ) capacitor c=0.00271584f \
 //x=73.63 //y=0 //x2=33.49 //y2=0.365
cc_717 ( N_GND_c_146_p N_noxref_37_M20_noxref_s ) capacitor c=0.014783f \
 //x=34.025 //y=0 //x2=33.49 //y2=0.365
cc_718 ( N_GND_c_11_p N_noxref_37_M20_noxref_s ) capacitor c=0.058339f \
 //x=32.93 //y=0 //x2=33.49 //y2=0.365
cc_719 ( N_GND_c_12_p N_noxref_37_M20_noxref_s ) capacitor c=0.00198043f \
 //x=36.26 //y=0 //x2=33.49 //y2=0.365
cc_720 ( N_GND_M20_noxref_d N_noxref_37_M20_noxref_s ) capacitor c=0.0334197f \
 //x=33.92 //y=0.865 //x2=33.49 //y2=0.365
cc_721 ( N_GND_c_23_p N_noxref_38_c_8837_n ) capacitor c=0.00530453f //x=73.63 \
 //y=0 //x2=37.84 //y2=1.58
cc_722 ( N_GND_c_172_p N_noxref_38_c_8837_n ) capacitor c=0.00112921f \
 //x=37.355 //y=0 //x2=37.84 //y2=1.58
cc_723 ( N_GND_c_179_p N_noxref_38_c_8837_n ) capacitor c=0.00182339f \
 //x=39.42 //y=0 //x2=37.84 //y2=1.58
cc_724 ( N_GND_M22_noxref_d N_noxref_38_c_8837_n ) capacitor c=0.00879185f \
 //x=37.25 //y=0.865 //x2=37.84 //y2=1.58
cc_725 ( N_GND_c_23_p N_noxref_38_c_8841_n ) capacitor c=0.00268165f //x=73.63 \
 //y=0 //x2=37.925 //y2=0.615
cc_726 ( N_GND_c_179_p N_noxref_38_c_8841_n ) capacitor c=0.014447f //x=39.42 \
 //y=0 //x2=37.925 //y2=0.615
cc_727 ( N_GND_M22_noxref_d N_noxref_38_c_8841_n ) capacitor c=0.033812f \
 //x=37.25 //y=0.865 //x2=37.925 //y2=0.615
cc_728 ( N_GND_c_12_p N_noxref_38_c_8844_n ) capacitor c=2.91423e-19 //x=36.26 \
 //y=0 //x2=37.925 //y2=1.495
cc_729 ( N_GND_c_23_p N_noxref_38_c_8845_n ) capacitor c=0.0106805f //x=73.63 \
 //y=0 //x2=38.81 //y2=0.53
cc_730 ( N_GND_c_179_p N_noxref_38_c_8845_n ) capacitor c=0.0374231f //x=39.42 \
 //y=0 //x2=38.81 //y2=0.53
cc_731 ( N_GND_c_2_p N_noxref_38_c_8845_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=38.81 //y2=0.53
cc_732 ( N_GND_c_23_p N_noxref_38_c_8848_n ) capacitor c=0.00258845f //x=73.63 \
 //y=0 //x2=38.895 //y2=0.615
cc_733 ( N_GND_c_179_p N_noxref_38_c_8848_n ) capacitor c=0.0146256f //x=39.42 \
 //y=0 //x2=38.895 //y2=0.615
cc_734 ( N_GND_c_13_p N_noxref_38_c_8848_n ) capacitor c=0.0431718f //x=39.59 \
 //y=0 //x2=38.895 //y2=0.615
cc_735 ( N_GND_c_23_p N_noxref_38_M22_noxref_s ) capacitor c=0.00271584f \
 //x=73.63 //y=0 //x2=36.82 //y2=0.365
cc_736 ( N_GND_c_172_p N_noxref_38_M22_noxref_s ) capacitor c=0.014783f \
 //x=37.355 //y=0 //x2=36.82 //y2=0.365
cc_737 ( N_GND_c_12_p N_noxref_38_M22_noxref_s ) capacitor c=0.058339f \
 //x=36.26 //y=0 //x2=36.82 //y2=0.365
cc_738 ( N_GND_c_13_p N_noxref_38_M22_noxref_s ) capacitor c=0.00198043f \
 //x=39.59 //y=0 //x2=36.82 //y2=0.365
cc_739 ( N_GND_M22_noxref_d N_noxref_38_M22_noxref_s ) capacitor c=0.0334197f \
 //x=37.25 //y=0.865 //x2=36.82 //y2=0.365
cc_740 ( N_GND_c_23_p N_noxref_39_c_8891_n ) capacitor c=0.00517234f //x=73.63 \
 //y=0 //x2=41.17 //y2=1.58
cc_741 ( N_GND_c_186_p N_noxref_39_c_8891_n ) capacitor c=0.00112872f \
 //x=40.685 //y=0 //x2=41.17 //y2=1.58
cc_742 ( N_GND_c_193_p N_noxref_39_c_8891_n ) capacitor c=0.0018229f //x=42.75 \
 //y=0 //x2=41.17 //y2=1.58
cc_743 ( N_GND_M24_noxref_d N_noxref_39_c_8891_n ) capacitor c=0.008625f \
 //x=40.58 //y=0.865 //x2=41.17 //y2=1.58
cc_744 ( N_GND_c_23_p N_noxref_39_c_8895_n ) capacitor c=0.00259029f //x=73.63 \
 //y=0 //x2=41.255 //y2=0.615
cc_745 ( N_GND_c_193_p N_noxref_39_c_8895_n ) capacitor c=0.0146901f //x=42.75 \
 //y=0 //x2=41.255 //y2=0.615
cc_746 ( N_GND_M24_noxref_d N_noxref_39_c_8895_n ) capacitor c=0.033812f \
 //x=40.58 //y=0.865 //x2=41.255 //y2=0.615
cc_747 ( N_GND_c_13_p N_noxref_39_c_8898_n ) capacitor c=2.91423e-19 //x=39.59 \
 //y=0 //x2=41.255 //y2=1.495
cc_748 ( N_GND_c_23_p N_noxref_39_c_8899_n ) capacitor c=0.0106879f //x=73.63 \
 //y=0 //x2=42.14 //y2=0.53
cc_749 ( N_GND_c_193_p N_noxref_39_c_8899_n ) capacitor c=0.0374232f //x=42.75 \
 //y=0 //x2=42.14 //y2=0.53
cc_750 ( N_GND_c_2_p N_noxref_39_c_8899_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=42.14 //y2=0.53
cc_751 ( N_GND_c_23_p N_noxref_39_c_8902_n ) capacitor c=0.00257855f //x=73.63 \
 //y=0 //x2=42.225 //y2=0.615
cc_752 ( N_GND_c_193_p N_noxref_39_c_8902_n ) capacitor c=0.0146181f //x=42.75 \
 //y=0 //x2=42.225 //y2=0.615
cc_753 ( N_GND_c_14_p N_noxref_39_c_8902_n ) capacitor c=0.0431718f //x=42.92 \
 //y=0 //x2=42.225 //y2=0.615
cc_754 ( N_GND_c_23_p N_noxref_39_M24_noxref_s ) capacitor c=0.00259029f \
 //x=73.63 //y=0 //x2=40.15 //y2=0.365
cc_755 ( N_GND_c_186_p N_noxref_39_M24_noxref_s ) capacitor c=0.0146901f \
 //x=40.685 //y=0 //x2=40.15 //y2=0.365
cc_756 ( N_GND_c_13_p N_noxref_39_M24_noxref_s ) capacitor c=0.058339f \
 //x=39.59 //y=0 //x2=40.15 //y2=0.365
cc_757 ( N_GND_c_14_p N_noxref_39_M24_noxref_s ) capacitor c=0.00198098f \
 //x=42.92 //y=0 //x2=40.15 //y2=0.365
cc_758 ( N_GND_M24_noxref_d N_noxref_39_M24_noxref_s ) capacitor c=0.0334197f \
 //x=40.58 //y=0.865 //x2=40.15 //y2=0.365
cc_759 ( N_GND_c_23_p N_noxref_40_c_8945_n ) capacitor c=0.00517576f //x=73.63 \
 //y=0 //x2=44.395 //y2=1.59
cc_760 ( N_GND_c_350_p N_noxref_40_c_8945_n ) capacitor c=0.00111448f \
 //x=43.91 //y=0 //x2=44.395 //y2=1.59
cc_761 ( N_GND_c_357_p N_noxref_40_c_8945_n ) capacitor c=0.00180612f \
 //x=47.56 //y=0 //x2=44.395 //y2=1.59
cc_762 ( N_GND_M26_noxref_d N_noxref_40_c_8945_n ) capacitor c=0.00853078f \
 //x=43.805 //y=0.875 //x2=44.395 //y2=1.59
cc_763 ( N_GND_c_23_p N_noxref_40_c_8949_n ) capacitor c=0.00254475f //x=73.63 \
 //y=0 //x2=44.48 //y2=0.625
cc_764 ( N_GND_c_357_p N_noxref_40_c_8949_n ) capacitor c=0.0140928f //x=47.56 \
 //y=0 //x2=44.48 //y2=0.625
cc_765 ( N_GND_M26_noxref_d N_noxref_40_c_8949_n ) capacitor c=0.033954f \
 //x=43.805 //y=0.875 //x2=44.48 //y2=0.625
cc_766 ( N_GND_c_23_p N_noxref_40_c_8952_n ) capacitor c=0.0104506f //x=73.63 \
 //y=0 //x2=45.365 //y2=0.54
cc_767 ( N_GND_c_357_p N_noxref_40_c_8952_n ) capacitor c=0.0360726f //x=47.56 \
 //y=0 //x2=45.365 //y2=0.54
cc_768 ( N_GND_c_2_p N_noxref_40_c_8952_n ) capacitor c=0.00178035f //x=73.63 \
 //y=0 //x2=45.365 //y2=0.54
cc_769 ( N_GND_c_23_p N_noxref_40_M26_noxref_s ) capacitor c=0.00507657f \
 //x=73.63 //y=0 //x2=43.375 //y2=0.375
cc_770 ( N_GND_c_350_p N_noxref_40_M26_noxref_s ) capacitor c=0.0140928f \
 //x=43.91 //y=0 //x2=43.375 //y2=0.375
cc_771 ( N_GND_c_357_p N_noxref_40_M26_noxref_s ) capacitor c=0.0136651f \
 //x=47.56 //y=0 //x2=43.375 //y2=0.375
cc_772 ( N_GND_c_14_p N_noxref_40_M26_noxref_s ) capacitor c=0.0696963f \
 //x=42.92 //y=0 //x2=43.375 //y2=0.375
cc_773 ( N_GND_c_15_p N_noxref_40_M26_noxref_s ) capacitor c=3.31601e-19 \
 //x=47.73 //y=0 //x2=43.375 //y2=0.375
cc_774 ( N_GND_M26_noxref_d N_noxref_40_M26_noxref_s ) capacitor c=0.033718f \
 //x=43.805 //y=0.875 //x2=43.375 //y2=0.375
cc_775 ( N_GND_c_23_p N_noxref_41_c_8995_n ) capacitor c=0.00352952f //x=73.63 \
 //y=0 //x2=45.935 //y2=0.995
cc_776 ( N_GND_c_357_p N_noxref_41_c_8995_n ) capacitor c=0.00934524f \
 //x=47.56 //y=0 //x2=45.935 //y2=0.995
cc_777 ( N_GND_c_23_p N_noxref_41_c_8997_n ) capacitor c=0.00254475f //x=73.63 \
 //y=0 //x2=46.02 //y2=0.625
cc_778 ( N_GND_c_357_p N_noxref_41_c_8997_n ) capacitor c=0.0140928f //x=47.56 \
 //y=0 //x2=46.02 //y2=0.625
cc_779 ( N_GND_M26_noxref_d N_noxref_41_c_8997_n ) capacitor c=6.21394e-19 \
 //x=43.805 //y=0.875 //x2=46.02 //y2=0.625
cc_780 ( N_GND_c_23_p N_noxref_41_c_9000_n ) capacitor c=0.0105317f //x=73.63 \
 //y=0 //x2=46.905 //y2=0.54
cc_781 ( N_GND_c_357_p N_noxref_41_c_9000_n ) capacitor c=0.036415f //x=47.56 \
 //y=0 //x2=46.905 //y2=0.54
cc_782 ( N_GND_c_2_p N_noxref_41_c_9000_n ) capacitor c=0.00190179f //x=73.63 \
 //y=0 //x2=46.905 //y2=0.54
cc_783 ( N_GND_c_23_p N_noxref_41_c_9003_n ) capacitor c=0.00254232f //x=73.63 \
 //y=0 //x2=46.99 //y2=0.625
cc_784 ( N_GND_c_357_p N_noxref_41_c_9003_n ) capacitor c=0.0140304f //x=47.56 \
 //y=0 //x2=46.99 //y2=0.625
cc_785 ( N_GND_c_15_p N_noxref_41_c_9003_n ) capacitor c=0.0404137f //x=47.73 \
 //y=0 //x2=46.99 //y2=0.625
cc_786 ( N_GND_M26_noxref_d N_noxref_41_M27_noxref_d ) capacitor c=0.00162435f \
 //x=43.805 //y=0.875 //x2=44.78 //y2=0.91
cc_787 ( N_GND_c_14_p N_noxref_41_M28_noxref_s ) capacitor c=8.16352e-19 \
 //x=42.92 //y=0 //x2=45.885 //y2=0.375
cc_788 ( N_GND_c_15_p N_noxref_41_M28_noxref_s ) capacitor c=0.00183576f \
 //x=47.73 //y=0 //x2=45.885 //y2=0.375
cc_789 ( N_GND_c_23_p N_noxref_42_c_9048_n ) capacitor c=0.00517234f //x=73.63 \
 //y=0 //x2=49.31 //y2=1.58
cc_790 ( N_GND_c_306_p N_noxref_42_c_9048_n ) capacitor c=0.00112872f \
 //x=48.825 //y=0 //x2=49.31 //y2=1.58
cc_791 ( N_GND_c_313_p N_noxref_42_c_9048_n ) capacitor c=0.0018229f //x=50.89 \
 //y=0 //x2=49.31 //y2=1.58
cc_792 ( N_GND_M29_noxref_d N_noxref_42_c_9048_n ) capacitor c=0.008625f \
 //x=48.72 //y=0.865 //x2=49.31 //y2=1.58
cc_793 ( N_GND_c_23_p N_noxref_42_c_9052_n ) capacitor c=0.00259029f //x=73.63 \
 //y=0 //x2=49.395 //y2=0.615
cc_794 ( N_GND_c_313_p N_noxref_42_c_9052_n ) capacitor c=0.0146901f //x=50.89 \
 //y=0 //x2=49.395 //y2=0.615
cc_795 ( N_GND_M29_noxref_d N_noxref_42_c_9052_n ) capacitor c=0.033812f \
 //x=48.72 //y=0.865 //x2=49.395 //y2=0.615
cc_796 ( N_GND_c_15_p N_noxref_42_c_9055_n ) capacitor c=2.91423e-19 //x=47.73 \
 //y=0 //x2=49.395 //y2=1.495
cc_797 ( N_GND_c_23_p N_noxref_42_c_9056_n ) capacitor c=0.0106919f //x=73.63 \
 //y=0 //x2=50.28 //y2=0.53
cc_798 ( N_GND_c_313_p N_noxref_42_c_9056_n ) capacitor c=0.0374253f //x=50.89 \
 //y=0 //x2=50.28 //y2=0.53
cc_799 ( N_GND_c_2_p N_noxref_42_c_9056_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=50.28 //y2=0.53
cc_800 ( N_GND_c_23_p N_noxref_42_c_9059_n ) capacitor c=0.00258845f //x=73.63 \
 //y=0 //x2=50.365 //y2=0.615
cc_801 ( N_GND_c_313_p N_noxref_42_c_9059_n ) capacitor c=0.0146256f //x=50.89 \
 //y=0 //x2=50.365 //y2=0.615
cc_802 ( N_GND_c_16_p N_noxref_42_c_9059_n ) capacitor c=0.0431718f //x=51.06 \
 //y=0 //x2=50.365 //y2=0.615
cc_803 ( N_GND_c_23_p N_noxref_42_M29_noxref_s ) capacitor c=0.00259029f \
 //x=73.63 //y=0 //x2=48.29 //y2=0.365
cc_804 ( N_GND_c_306_p N_noxref_42_M29_noxref_s ) capacitor c=0.0146901f \
 //x=48.825 //y=0 //x2=48.29 //y2=0.365
cc_805 ( N_GND_c_15_p N_noxref_42_M29_noxref_s ) capacitor c=0.0583534f \
 //x=47.73 //y=0 //x2=48.29 //y2=0.365
cc_806 ( N_GND_c_16_p N_noxref_42_M29_noxref_s ) capacitor c=0.00198043f \
 //x=51.06 //y=0 //x2=48.29 //y2=0.365
cc_807 ( N_GND_M29_noxref_d N_noxref_42_M29_noxref_s ) capacitor c=0.0334197f \
 //x=48.72 //y=0.865 //x2=48.29 //y2=0.365
cc_808 ( N_GND_c_23_p N_noxref_43_c_9100_n ) capacitor c=0.00517234f //x=73.63 \
 //y=0 //x2=52.64 //y2=1.58
cc_809 ( N_GND_c_265_p N_noxref_43_c_9100_n ) capacitor c=0.00112872f \
 //x=52.155 //y=0 //x2=52.64 //y2=1.58
cc_810 ( N_GND_c_272_p N_noxref_43_c_9100_n ) capacitor c=0.0018229f //x=54.22 \
 //y=0 //x2=52.64 //y2=1.58
cc_811 ( N_GND_M31_noxref_d N_noxref_43_c_9100_n ) capacitor c=0.008625f \
 //x=52.05 //y=0.865 //x2=52.64 //y2=1.58
cc_812 ( N_GND_c_23_p N_noxref_43_c_9104_n ) capacitor c=0.00259029f //x=73.63 \
 //y=0 //x2=52.725 //y2=0.615
cc_813 ( N_GND_c_272_p N_noxref_43_c_9104_n ) capacitor c=0.0146901f //x=54.22 \
 //y=0 //x2=52.725 //y2=0.615
cc_814 ( N_GND_M31_noxref_d N_noxref_43_c_9104_n ) capacitor c=0.033812f \
 //x=52.05 //y=0.865 //x2=52.725 //y2=0.615
cc_815 ( N_GND_c_16_p N_noxref_43_c_9107_n ) capacitor c=2.91423e-19 //x=51.06 \
 //y=0 //x2=52.725 //y2=1.495
cc_816 ( N_GND_c_23_p N_noxref_43_c_9108_n ) capacitor c=0.0106919f //x=73.63 \
 //y=0 //x2=53.61 //y2=0.53
cc_817 ( N_GND_c_272_p N_noxref_43_c_9108_n ) capacitor c=0.0374253f //x=54.22 \
 //y=0 //x2=53.61 //y2=0.53
cc_818 ( N_GND_c_2_p N_noxref_43_c_9108_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=53.61 //y2=0.53
cc_819 ( N_GND_c_23_p N_noxref_43_c_9111_n ) capacitor c=0.00258845f //x=73.63 \
 //y=0 //x2=53.695 //y2=0.615
cc_820 ( N_GND_c_272_p N_noxref_43_c_9111_n ) capacitor c=0.0146256f //x=54.22 \
 //y=0 //x2=53.695 //y2=0.615
cc_821 ( N_GND_c_17_p N_noxref_43_c_9111_n ) capacitor c=0.0431718f //x=54.39 \
 //y=0 //x2=53.695 //y2=0.615
cc_822 ( N_GND_c_23_p N_noxref_43_M31_noxref_s ) capacitor c=0.00259029f \
 //x=73.63 //y=0 //x2=51.62 //y2=0.365
cc_823 ( N_GND_c_265_p N_noxref_43_M31_noxref_s ) capacitor c=0.0146901f \
 //x=52.155 //y=0 //x2=51.62 //y2=0.365
cc_824 ( N_GND_c_16_p N_noxref_43_M31_noxref_s ) capacitor c=0.058339f \
 //x=51.06 //y=0 //x2=51.62 //y2=0.365
cc_825 ( N_GND_c_17_p N_noxref_43_M31_noxref_s ) capacitor c=0.00198043f \
 //x=54.39 //y=0 //x2=51.62 //y2=0.365
cc_826 ( N_GND_M31_noxref_d N_noxref_43_M31_noxref_s ) capacitor c=0.0334197f \
 //x=52.05 //y=0.865 //x2=51.62 //y2=0.365
cc_827 ( N_GND_c_23_p N_noxref_44_c_9152_n ) capacitor c=0.00517234f //x=73.63 \
 //y=0 //x2=55.97 //y2=1.58
cc_828 ( N_GND_c_281_p N_noxref_44_c_9152_n ) capacitor c=0.00112872f \
 //x=55.485 //y=0 //x2=55.97 //y2=1.58
cc_829 ( N_GND_c_288_p N_noxref_44_c_9152_n ) capacitor c=0.0018229f //x=57.55 \
 //y=0 //x2=55.97 //y2=1.58
cc_830 ( N_GND_M33_noxref_d N_noxref_44_c_9152_n ) capacitor c=0.008625f \
 //x=55.38 //y=0.865 //x2=55.97 //y2=1.58
cc_831 ( N_GND_c_23_p N_noxref_44_c_9156_n ) capacitor c=0.00259029f //x=73.63 \
 //y=0 //x2=56.055 //y2=0.615
cc_832 ( N_GND_c_288_p N_noxref_44_c_9156_n ) capacitor c=0.0146901f //x=57.55 \
 //y=0 //x2=56.055 //y2=0.615
cc_833 ( N_GND_M33_noxref_d N_noxref_44_c_9156_n ) capacitor c=0.033812f \
 //x=55.38 //y=0.865 //x2=56.055 //y2=0.615
cc_834 ( N_GND_c_17_p N_noxref_44_c_9159_n ) capacitor c=2.91423e-19 //x=54.39 \
 //y=0 //x2=56.055 //y2=1.495
cc_835 ( N_GND_c_23_p N_noxref_44_c_9160_n ) capacitor c=0.0106919f //x=73.63 \
 //y=0 //x2=56.94 //y2=0.53
cc_836 ( N_GND_c_288_p N_noxref_44_c_9160_n ) capacitor c=0.0374253f //x=57.55 \
 //y=0 //x2=56.94 //y2=0.53
cc_837 ( N_GND_c_2_p N_noxref_44_c_9160_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=56.94 //y2=0.53
cc_838 ( N_GND_c_23_p N_noxref_44_c_9163_n ) capacitor c=0.00258845f //x=73.63 \
 //y=0 //x2=57.025 //y2=0.615
cc_839 ( N_GND_c_288_p N_noxref_44_c_9163_n ) capacitor c=0.0146256f //x=57.55 \
 //y=0 //x2=57.025 //y2=0.615
cc_840 ( N_GND_c_18_p N_noxref_44_c_9163_n ) capacitor c=0.0431718f //x=57.72 \
 //y=0 //x2=57.025 //y2=0.615
cc_841 ( N_GND_c_23_p N_noxref_44_M33_noxref_s ) capacitor c=0.00259029f \
 //x=73.63 //y=0 //x2=54.95 //y2=0.365
cc_842 ( N_GND_c_281_p N_noxref_44_M33_noxref_s ) capacitor c=0.0146901f \
 //x=55.485 //y=0 //x2=54.95 //y2=0.365
cc_843 ( N_GND_c_17_p N_noxref_44_M33_noxref_s ) capacitor c=0.058339f \
 //x=54.39 //y=0 //x2=54.95 //y2=0.365
cc_844 ( N_GND_c_18_p N_noxref_44_M33_noxref_s ) capacitor c=0.00198043f \
 //x=57.72 //y=0 //x2=54.95 //y2=0.365
cc_845 ( N_GND_M33_noxref_d N_noxref_44_M33_noxref_s ) capacitor c=0.0334197f \
 //x=55.38 //y=0.865 //x2=54.95 //y2=0.365
cc_846 ( N_GND_c_23_p N_noxref_45_c_9204_n ) capacitor c=0.00517234f //x=73.63 \
 //y=0 //x2=59.3 //y2=1.58
cc_847 ( N_GND_c_316_p N_noxref_45_c_9204_n ) capacitor c=0.00112872f \
 //x=58.815 //y=0 //x2=59.3 //y2=1.58
cc_848 ( N_GND_c_323_p N_noxref_45_c_9204_n ) capacitor c=0.0018229f //x=60.88 \
 //y=0 //x2=59.3 //y2=1.58
cc_849 ( N_GND_M35_noxref_d N_noxref_45_c_9204_n ) capacitor c=0.008625f \
 //x=58.71 //y=0.865 //x2=59.3 //y2=1.58
cc_850 ( N_GND_c_23_p N_noxref_45_c_9208_n ) capacitor c=0.00259029f //x=73.63 \
 //y=0 //x2=59.385 //y2=0.615
cc_851 ( N_GND_c_323_p N_noxref_45_c_9208_n ) capacitor c=0.0143795f //x=60.88 \
 //y=0 //x2=59.385 //y2=0.615
cc_852 ( N_GND_M35_noxref_d N_noxref_45_c_9208_n ) capacitor c=0.033812f \
 //x=58.71 //y=0.865 //x2=59.385 //y2=0.615
cc_853 ( N_GND_c_18_p N_noxref_45_c_9211_n ) capacitor c=2.91423e-19 //x=57.72 \
 //y=0 //x2=59.385 //y2=1.495
cc_854 ( N_GND_c_23_p N_noxref_45_c_9212_n ) capacitor c=0.0106919f //x=73.63 \
 //y=0 //x2=60.27 //y2=0.53
cc_855 ( N_GND_c_323_p N_noxref_45_c_9212_n ) capacitor c=0.0374253f //x=60.88 \
 //y=0 //x2=60.27 //y2=0.53
cc_856 ( N_GND_c_2_p N_noxref_45_c_9212_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=60.27 //y2=0.53
cc_857 ( N_GND_c_23_p N_noxref_45_c_9215_n ) capacitor c=0.00258845f //x=73.63 \
 //y=0 //x2=60.355 //y2=0.615
cc_858 ( N_GND_c_323_p N_noxref_45_c_9215_n ) capacitor c=0.0146256f //x=60.88 \
 //y=0 //x2=60.355 //y2=0.615
cc_859 ( N_GND_c_19_p N_noxref_45_c_9215_n ) capacitor c=0.0431718f //x=61.05 \
 //y=0 //x2=60.355 //y2=0.615
cc_860 ( N_GND_c_23_p N_noxref_45_M35_noxref_s ) capacitor c=0.00259029f \
 //x=73.63 //y=0 //x2=58.28 //y2=0.365
cc_861 ( N_GND_c_316_p N_noxref_45_M35_noxref_s ) capacitor c=0.0146901f \
 //x=58.815 //y=0 //x2=58.28 //y2=0.365
cc_862 ( N_GND_c_18_p N_noxref_45_M35_noxref_s ) capacitor c=0.058339f \
 //x=57.72 //y=0 //x2=58.28 //y2=0.365
cc_863 ( N_GND_c_19_p N_noxref_45_M35_noxref_s ) capacitor c=0.00198043f \
 //x=61.05 //y=0 //x2=58.28 //y2=0.365
cc_864 ( N_GND_M35_noxref_d N_noxref_45_M35_noxref_s ) capacitor c=0.0334197f \
 //x=58.71 //y=0.865 //x2=58.28 //y2=0.365
cc_865 ( N_GND_c_23_p N_noxref_46_c_9256_n ) capacitor c=0.00517234f //x=73.63 \
 //y=0 //x2=62.63 //y2=1.58
cc_866 ( N_GND_c_330_p N_noxref_46_c_9256_n ) capacitor c=0.00112872f \
 //x=62.145 //y=0 //x2=62.63 //y2=1.58
cc_867 ( N_GND_c_337_p N_noxref_46_c_9256_n ) capacitor c=0.0018229f //x=64.21 \
 //y=0 //x2=62.63 //y2=1.58
cc_868 ( N_GND_M37_noxref_d N_noxref_46_c_9256_n ) capacitor c=0.008625f \
 //x=62.04 //y=0.865 //x2=62.63 //y2=1.58
cc_869 ( N_GND_c_23_p N_noxref_46_c_9260_n ) capacitor c=0.00259029f //x=73.63 \
 //y=0 //x2=62.715 //y2=0.615
cc_870 ( N_GND_c_337_p N_noxref_46_c_9260_n ) capacitor c=0.0146901f //x=64.21 \
 //y=0 //x2=62.715 //y2=0.615
cc_871 ( N_GND_M37_noxref_d N_noxref_46_c_9260_n ) capacitor c=0.033812f \
 //x=62.04 //y=0.865 //x2=62.715 //y2=0.615
cc_872 ( N_GND_c_19_p N_noxref_46_c_9263_n ) capacitor c=2.91423e-19 //x=61.05 \
 //y=0 //x2=62.715 //y2=1.495
cc_873 ( N_GND_c_23_p N_noxref_46_c_9264_n ) capacitor c=0.0106919f //x=73.63 \
 //y=0 //x2=63.6 //y2=0.53
cc_874 ( N_GND_c_337_p N_noxref_46_c_9264_n ) capacitor c=0.0374253f //x=64.21 \
 //y=0 //x2=63.6 //y2=0.53
cc_875 ( N_GND_c_2_p N_noxref_46_c_9264_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=63.6 //y2=0.53
cc_876 ( N_GND_c_23_p N_noxref_46_c_9267_n ) capacitor c=0.00258845f //x=73.63 \
 //y=0 //x2=63.685 //y2=0.615
cc_877 ( N_GND_c_337_p N_noxref_46_c_9267_n ) capacitor c=0.0146256f //x=64.21 \
 //y=0 //x2=63.685 //y2=0.615
cc_878 ( N_GND_c_20_p N_noxref_46_c_9267_n ) capacitor c=0.0427915f //x=64.38 \
 //y=0 //x2=63.685 //y2=0.615
cc_879 ( N_GND_c_23_p N_noxref_46_M37_noxref_s ) capacitor c=0.00259029f \
 //x=73.63 //y=0 //x2=61.61 //y2=0.365
cc_880 ( N_GND_c_330_p N_noxref_46_M37_noxref_s ) capacitor c=0.0146901f \
 //x=62.145 //y=0 //x2=61.61 //y2=0.365
cc_881 ( N_GND_c_19_p N_noxref_46_M37_noxref_s ) capacitor c=0.058339f \
 //x=61.05 //y=0 //x2=61.61 //y2=0.365
cc_882 ( N_GND_c_20_p N_noxref_46_M37_noxref_s ) capacitor c=0.00198098f \
 //x=64.38 //y=0 //x2=61.61 //y2=0.365
cc_883 ( N_GND_M37_noxref_d N_noxref_46_M37_noxref_s ) capacitor c=0.0334197f \
 //x=62.04 //y=0.865 //x2=61.61 //y2=0.365
cc_884 ( N_GND_c_23_p N_noxref_47_c_9308_n ) capacitor c=0.00521624f //x=73.63 \
 //y=0 //x2=65.96 //y2=1.58
cc_885 ( N_GND_c_372_p N_noxref_47_c_9308_n ) capacitor c=0.00112872f \
 //x=65.475 //y=0 //x2=65.96 //y2=1.58
cc_886 ( N_GND_c_379_p N_noxref_47_c_9308_n ) capacitor c=0.0018229f //x=67.54 \
 //y=0 //x2=65.96 //y2=1.58
cc_887 ( N_GND_M39_noxref_d N_noxref_47_c_9308_n ) capacitor c=0.00892401f \
 //x=65.37 //y=0.865 //x2=65.96 //y2=1.58
cc_888 ( N_GND_c_23_p N_noxref_47_c_9312_n ) capacitor c=0.00258934f //x=73.63 \
 //y=0 //x2=66.045 //y2=0.615
cc_889 ( N_GND_c_379_p N_noxref_47_c_9312_n ) capacitor c=0.0146894f //x=67.54 \
 //y=0 //x2=66.045 //y2=0.615
cc_890 ( N_GND_M39_noxref_d N_noxref_47_c_9312_n ) capacitor c=0.0336822f \
 //x=65.37 //y=0.865 //x2=66.045 //y2=0.615
cc_891 ( N_GND_c_20_p N_noxref_47_c_9315_n ) capacitor c=2.91423e-19 //x=64.38 \
 //y=0 //x2=66.045 //y2=1.495
cc_892 ( N_GND_c_23_p N_noxref_47_c_9316_n ) capacitor c=0.00942854f //x=73.63 \
 //y=0 //x2=66.93 //y2=0.53
cc_893 ( N_GND_c_379_p N_noxref_47_c_9316_n ) capacitor c=0.0374756f //x=67.54 \
 //y=0 //x2=66.93 //y2=0.53
cc_894 ( N_GND_c_2_p N_noxref_47_c_9316_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=66.93 //y2=0.53
cc_895 ( N_GND_c_23_p N_noxref_47_c_9319_n ) capacitor c=0.00212661f //x=73.63 \
 //y=0 //x2=67.015 //y2=0.615
cc_896 ( N_GND_c_379_p N_noxref_47_c_9319_n ) capacitor c=0.0143168f //x=67.54 \
 //y=0 //x2=67.015 //y2=0.615
cc_897 ( N_GND_c_21_p N_noxref_47_c_9319_n ) capacitor c=0.0554337f //x=67.71 \
 //y=0 //x2=67.015 //y2=0.615
cc_898 ( N_GND_c_23_p N_noxref_47_M39_noxref_s ) capacitor c=0.00259029f \
 //x=73.63 //y=0 //x2=64.94 //y2=0.365
cc_899 ( N_GND_c_372_p N_noxref_47_M39_noxref_s ) capacitor c=0.0146901f \
 //x=65.475 //y=0 //x2=64.94 //y2=0.365
cc_900 ( N_GND_c_20_p N_noxref_47_M39_noxref_s ) capacitor c=0.0587986f \
 //x=64.38 //y=0 //x2=64.94 //y2=0.365
cc_901 ( N_GND_c_21_p N_noxref_47_M39_noxref_s ) capacitor c=0.00181744f \
 //x=67.71 //y=0 //x2=64.94 //y2=0.365
cc_902 ( N_GND_M39_noxref_d N_noxref_47_M39_noxref_s ) capacitor c=0.0333456f \
 //x=65.37 //y=0.865 //x2=64.94 //y2=0.365
cc_903 ( N_GND_c_382_p N_noxref_48_c_9366_n ) capacitor c=8.01905e-19 \
 //x=68.805 //y=0 //x2=69.29 //y2=1.58
cc_904 ( N_GND_c_388_p N_noxref_48_c_9366_n ) capacitor c=0.00161527f \
 //x=70.87 //y=0 //x2=69.29 //y2=1.58
cc_905 ( N_GND_M41_noxref_d N_noxref_48_c_9366_n ) capacitor c=0.0073276f \
 //x=68.7 //y=0.865 //x2=69.29 //y2=1.58
cc_906 ( N_GND_c_23_p N_noxref_48_c_9369_n ) capacitor c=0.00212661f //x=73.63 \
 //y=0 //x2=69.375 //y2=0.615
cc_907 ( N_GND_c_388_p N_noxref_48_c_9369_n ) capacitor c=0.0143168f //x=70.87 \
 //y=0 //x2=69.375 //y2=0.615
cc_908 ( N_GND_M41_noxref_d N_noxref_48_c_9369_n ) capacitor c=0.0336587f \
 //x=68.7 //y=0.865 //x2=69.375 //y2=0.615
cc_909 ( N_GND_c_21_p N_noxref_48_c_9372_n ) capacitor c=2.91423e-19 //x=67.71 \
 //y=0 //x2=69.375 //y2=1.495
cc_910 ( N_GND_c_23_p N_noxref_48_c_9373_n ) capacitor c=0.00884129f //x=73.63 \
 //y=0 //x2=70.26 //y2=0.53
cc_911 ( N_GND_c_388_p N_noxref_48_c_9373_n ) capacitor c=0.0373651f //x=70.87 \
 //y=0 //x2=70.26 //y2=0.53
cc_912 ( N_GND_c_2_p N_noxref_48_c_9373_n ) capacitor c=0.00199232f //x=73.63 \
 //y=0 //x2=70.26 //y2=0.53
cc_913 ( N_GND_c_23_p N_noxref_48_c_9376_n ) capacitor c=0.00212661f //x=73.63 \
 //y=0 //x2=70.345 //y2=0.615
cc_914 ( N_GND_c_388_p N_noxref_48_c_9376_n ) capacitor c=0.0143168f //x=70.87 \
 //y=0 //x2=70.345 //y2=0.615
cc_915 ( N_GND_c_22_p N_noxref_48_c_9376_n ) capacitor c=0.0548042f //x=71.04 \
 //y=0 //x2=70.345 //y2=0.615
cc_916 ( N_GND_c_23_p N_noxref_48_M41_noxref_s ) capacitor c=0.00212661f \
 //x=73.63 //y=0 //x2=68.27 //y2=0.365
cc_917 ( N_GND_c_382_p N_noxref_48_M41_noxref_s ) capacitor c=0.0143168f \
 //x=68.805 //y=0 //x2=68.27 //y2=0.365
cc_918 ( N_GND_c_21_p N_noxref_48_M41_noxref_s ) capacitor c=0.0561194f \
 //x=67.71 //y=0 //x2=68.27 //y2=0.365
cc_919 ( N_GND_c_22_p N_noxref_48_M41_noxref_s ) capacitor c=0.0022128f \
 //x=71.04 //y=0 //x2=68.27 //y2=0.365
cc_920 ( N_GND_M41_noxref_d N_noxref_48_M41_noxref_s ) capacitor c=0.0332904f \
 //x=68.7 //y=0.865 //x2=68.27 //y2=0.365
cc_921 ( N_GND_c_469_p N_noxref_49_c_9422_n ) capacitor c=8.01912e-19 \
 //x=72.135 //y=0 //x2=72.62 //y2=1.58
cc_922 ( N_GND_c_2_p N_noxref_49_c_9422_n ) capacitor c=0.00161527f //x=73.63 \
 //y=0 //x2=72.62 //y2=1.58
cc_923 ( N_GND_M43_noxref_d N_noxref_49_c_9422_n ) capacitor c=0.0073482f \
 //x=72.03 //y=0.865 //x2=72.62 //y2=1.58
cc_924 ( N_GND_c_23_p N_noxref_49_c_9425_n ) capacitor c=0.00212661f //x=73.63 \
 //y=0 //x2=72.705 //y2=0.615
cc_925 ( N_GND_c_2_p N_noxref_49_c_9425_n ) capacitor c=0.0143168f //x=73.63 \
 //y=0 //x2=72.705 //y2=0.615
cc_926 ( N_GND_M43_noxref_d N_noxref_49_c_9425_n ) capacitor c=0.0336587f \
 //x=72.03 //y=0.865 //x2=72.705 //y2=0.615
cc_927 ( N_GND_c_22_p N_noxref_49_c_9428_n ) capacitor c=2.91423e-19 //x=71.04 \
 //y=0 //x2=72.705 //y2=1.495
cc_928 ( N_GND_c_23_p N_noxref_49_c_9429_n ) capacitor c=0.0127012f //x=73.63 \
 //y=0 //x2=73.59 //y2=0.53
cc_929 ( N_GND_c_2_p N_noxref_49_c_9429_n ) capacitor c=0.0391711f //x=73.63 \
 //y=0 //x2=73.59 //y2=0.53
cc_930 ( N_GND_c_23_p N_noxref_49_c_9431_n ) capacitor c=0.00719686f //x=73.63 \
 //y=0 //x2=73.675 //y2=0.615
cc_931 ( N_GND_c_2_p N_noxref_49_c_9431_n ) capacitor c=0.0581858f //x=73.63 \
 //y=0 //x2=73.675 //y2=0.615
cc_932 ( N_GND_c_23_p N_noxref_49_M43_noxref_s ) capacitor c=0.00212661f \
 //x=73.63 //y=0 //x2=71.6 //y2=0.365
cc_933 ( N_GND_c_469_p N_noxref_49_M43_noxref_s ) capacitor c=0.0143168f \
 //x=72.135 //y=0 //x2=71.6 //y2=0.365
cc_934 ( N_GND_c_2_p N_noxref_49_M43_noxref_s ) capacitor c=0.00202267f \
 //x=73.63 //y=0 //x2=71.6 //y2=0.365
cc_935 ( N_GND_c_22_p N_noxref_49_M43_noxref_s ) capacitor c=0.0555228f \
 //x=71.04 //y=0 //x2=71.6 //y2=0.365
cc_936 ( N_GND_M43_noxref_d N_noxref_49_M43_noxref_s ) capacitor c=0.0332904f \
 //x=72.03 //y=0.865 //x2=71.6 //y2=0.365
cc_937 ( N_VDD_c_939_n N_noxref_3_c_1941_n ) capacitor c=6.58823e-19 //x=4.81 \
 //y=7.4 //x2=3.33 //y2=2.08
cc_938 ( N_VDD_c_960_p N_noxref_3_c_1959_n ) capacitor c=0.00453663f //x=73.63 \
 //y=7.4 //x2=6.835 //y2=5.2
cc_939 ( N_VDD_c_961_p N_noxref_3_c_1959_n ) capacitor c=4.48391e-19 //x=6.395 \
 //y=7.4 //x2=6.835 //y2=5.2
cc_940 ( N_VDD_c_962_p N_noxref_3_c_1959_n ) capacitor c=4.48391e-19 //x=7.275 \
 //y=7.4 //x2=6.835 //y2=5.2
cc_941 ( N_VDD_M52_noxref_d N_noxref_3_c_1959_n ) capacitor c=0.0124542f \
 //x=6.335 //y=5.02 //x2=6.835 //y2=5.2
cc_942 ( N_VDD_c_939_n N_noxref_3_c_1963_n ) capacitor c=0.00985474f //x=4.81 \
 //y=7.4 //x2=6.125 //y2=5.2
cc_943 ( N_VDD_M51_noxref_s N_noxref_3_c_1963_n ) capacitor c=0.087833f \
 //x=5.465 //y=5.02 //x2=6.125 //y2=5.2
cc_944 ( N_VDD_c_960_p N_noxref_3_c_1965_n ) capacitor c=0.00301575f //x=73.63 \
 //y=7.4 //x2=7.315 //y2=5.2
cc_945 ( N_VDD_c_962_p N_noxref_3_c_1965_n ) capacitor c=7.72068e-19 //x=7.275 \
 //y=7.4 //x2=7.315 //y2=5.2
cc_946 ( N_VDD_M54_noxref_d N_noxref_3_c_1965_n ) capacitor c=0.0158515f \
 //x=7.215 //y=5.02 //x2=7.315 //y2=5.2
cc_947 ( N_VDD_M55_noxref_s N_noxref_3_c_1965_n ) capacitor c=2.44532e-19 \
 //x=8.795 //y=5.02 //x2=7.315 //y2=5.2
cc_948 ( N_VDD_c_939_n N_noxref_3_c_1943_n ) capacitor c=0.00151618f //x=4.81 \
 //y=7.4 //x2=7.4 //y2=3.33
cc_949 ( N_VDD_c_940_n N_noxref_3_c_1943_n ) capacitor c=0.0429414f //x=8.14 \
 //y=7.4 //x2=7.4 //y2=3.33
cc_950 ( N_VDD_c_960_p N_noxref_3_c_1944_n ) capacitor c=0.00125279f //x=73.63 \
 //y=7.4 //x2=9.25 //y2=2.08
cc_951 ( N_VDD_c_973_p N_noxref_3_c_1944_n ) capacitor c=2.87256e-19 //x=9.725 \
 //y=7.4 //x2=9.25 //y2=2.08
cc_952 ( N_VDD_c_940_n N_noxref_3_c_1944_n ) capacitor c=0.0134208f //x=8.14 \
 //y=7.4 //x2=9.25 //y2=2.08
cc_953 ( N_VDD_c_975_p N_noxref_3_M49_noxref_g ) capacitor c=0.00675175f \
 //x=3.645 //y=7.4 //x2=3.07 //y2=6.02
cc_954 ( N_VDD_M48_noxref_d N_noxref_3_M49_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=3.07 //y2=6.02
cc_955 ( N_VDD_c_975_p N_noxref_3_M50_noxref_g ) capacitor c=0.00675379f \
 //x=3.645 //y=7.4 //x2=3.51 //y2=6.02
cc_956 ( N_VDD_M50_noxref_d N_noxref_3_M50_noxref_g ) capacitor c=0.0394719f \
 //x=3.585 //y=5.02 //x2=3.51 //y2=6.02
cc_957 ( N_VDD_c_973_p N_noxref_3_M55_noxref_g ) capacitor c=0.00726866f \
 //x=9.725 //y=7.4 //x2=9.15 //y2=6.02
cc_958 ( N_VDD_M55_noxref_s N_noxref_3_M55_noxref_g ) capacitor c=0.054195f \
 //x=8.795 //y=5.02 //x2=9.15 //y2=6.02
cc_959 ( N_VDD_c_973_p N_noxref_3_M56_noxref_g ) capacitor c=0.00672952f \
 //x=9.725 //y=7.4 //x2=9.59 //y2=6.02
cc_960 ( N_VDD_M56_noxref_d N_noxref_3_M56_noxref_g ) capacitor c=0.015318f \
 //x=9.665 //y=5.02 //x2=9.59 //y2=6.02
cc_961 ( N_VDD_c_940_n N_noxref_3_c_1982_n ) capacitor c=0.0150435f //x=8.14 \
 //y=7.4 //x2=9.25 //y2=4.7
cc_962 ( N_VDD_c_960_p N_noxref_3_M51_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=5.895 //y2=5.02
cc_963 ( N_VDD_c_961_p N_noxref_3_M51_noxref_d ) capacitor c=0.0140317f \
 //x=6.395 //y=7.4 //x2=5.895 //y2=5.02
cc_964 ( N_VDD_c_940_n N_noxref_3_M51_noxref_d ) capacitor c=6.94454e-19 \
 //x=8.14 //y=7.4 //x2=5.895 //y2=5.02
cc_965 ( N_VDD_M52_noxref_d N_noxref_3_M51_noxref_d ) capacitor c=0.0664752f \
 //x=6.335 //y=5.02 //x2=5.895 //y2=5.02
cc_966 ( N_VDD_c_960_p N_noxref_3_M53_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=6.775 //y2=5.02
cc_967 ( N_VDD_c_962_p N_noxref_3_M53_noxref_d ) capacitor c=0.0140317f \
 //x=7.275 //y=7.4 //x2=6.775 //y2=5.02
cc_968 ( N_VDD_c_940_n N_noxref_3_M53_noxref_d ) capacitor c=0.0120541f \
 //x=8.14 //y=7.4 //x2=6.775 //y2=5.02
cc_969 ( N_VDD_M51_noxref_s N_noxref_3_M53_noxref_d ) capacitor c=0.00111971f \
 //x=5.465 //y=5.02 //x2=6.775 //y2=5.02
cc_970 ( N_VDD_M52_noxref_d N_noxref_3_M53_noxref_d ) capacitor c=0.0664752f \
 //x=6.335 //y=5.02 //x2=6.775 //y2=5.02
cc_971 ( N_VDD_M54_noxref_d N_noxref_3_M53_noxref_d ) capacitor c=0.0664752f \
 //x=7.215 //y=5.02 //x2=6.775 //y2=5.02
cc_972 ( N_VDD_M55_noxref_s N_noxref_3_M53_noxref_d ) capacitor c=4.54516e-19 \
 //x=8.795 //y=5.02 //x2=6.775 //y2=5.02
cc_973 ( N_VDD_c_960_p N_noxref_4_c_2184_n ) capacitor c=0.00453663f //x=73.63 \
 //y=7.4 //x2=10.165 //y2=5.2
cc_974 ( N_VDD_c_973_p N_noxref_4_c_2184_n ) capacitor c=4.48391e-19 //x=9.725 \
 //y=7.4 //x2=10.165 //y2=5.2
cc_975 ( N_VDD_c_997_p N_noxref_4_c_2184_n ) capacitor c=4.48391e-19 \
 //x=10.605 //y=7.4 //x2=10.165 //y2=5.2
cc_976 ( N_VDD_M56_noxref_d N_noxref_4_c_2184_n ) capacitor c=0.0124542f \
 //x=9.665 //y=5.02 //x2=10.165 //y2=5.2
cc_977 ( N_VDD_c_940_n N_noxref_4_c_2188_n ) capacitor c=0.00985474f //x=8.14 \
 //y=7.4 //x2=9.455 //y2=5.2
cc_978 ( N_VDD_M55_noxref_s N_noxref_4_c_2188_n ) capacitor c=0.087833f \
 //x=8.795 //y=5.02 //x2=9.455 //y2=5.2
cc_979 ( N_VDD_c_960_p N_noxref_4_c_2190_n ) capacitor c=0.00301575f //x=73.63 \
 //y=7.4 //x2=10.645 //y2=5.2
cc_980 ( N_VDD_c_997_p N_noxref_4_c_2190_n ) capacitor c=7.72068e-19 \
 //x=10.605 //y=7.4 //x2=10.645 //y2=5.2
cc_981 ( N_VDD_M58_noxref_d N_noxref_4_c_2190_n ) capacitor c=0.0158515f \
 //x=10.545 //y=5.02 //x2=10.645 //y2=5.2
cc_982 ( N_VDD_M59_noxref_s N_noxref_4_c_2190_n ) capacitor c=2.44532e-19 \
 //x=12.125 //y=5.02 //x2=10.645 //y2=5.2
cc_983 ( N_VDD_c_940_n N_noxref_4_c_2169_n ) capacitor c=0.00151618f //x=8.14 \
 //y=7.4 //x2=10.73 //y2=3.33
cc_984 ( N_VDD_c_941_n N_noxref_4_c_2169_n ) capacitor c=0.0427674f //x=11.47 \
 //y=7.4 //x2=10.73 //y2=3.33
cc_985 ( N_VDD_c_960_p N_noxref_4_c_2170_n ) capacitor c=0.00125279f //x=73.63 \
 //y=7.4 //x2=12.58 //y2=2.08
cc_986 ( N_VDD_c_1008_p N_noxref_4_c_2170_n ) capacitor c=2.87256e-19 \
 //x=13.055 //y=7.4 //x2=12.58 //y2=2.08
cc_987 ( N_VDD_c_941_n N_noxref_4_c_2170_n ) capacitor c=0.0133228f //x=11.47 \
 //y=7.4 //x2=12.58 //y2=2.08
cc_988 ( N_VDD_c_1008_p N_noxref_4_M59_noxref_g ) capacitor c=0.00726866f \
 //x=13.055 //y=7.4 //x2=12.48 //y2=6.02
cc_989 ( N_VDD_M59_noxref_s N_noxref_4_M59_noxref_g ) capacitor c=0.054195f \
 //x=12.125 //y=5.02 //x2=12.48 //y2=6.02
cc_990 ( N_VDD_c_1008_p N_noxref_4_M60_noxref_g ) capacitor c=0.00672952f \
 //x=13.055 //y=7.4 //x2=12.92 //y2=6.02
cc_991 ( N_VDD_M60_noxref_d N_noxref_4_M60_noxref_g ) capacitor c=0.015318f \
 //x=12.995 //y=5.02 //x2=12.92 //y2=6.02
cc_992 ( N_VDD_c_941_n N_noxref_4_c_2203_n ) capacitor c=0.0149273f //x=11.47 \
 //y=7.4 //x2=12.58 //y2=4.7
cc_993 ( N_VDD_c_960_p N_noxref_4_M55_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=9.225 //y2=5.02
cc_994 ( N_VDD_c_973_p N_noxref_4_M55_noxref_d ) capacitor c=0.0140317f \
 //x=9.725 //y=7.4 //x2=9.225 //y2=5.02
cc_995 ( N_VDD_c_941_n N_noxref_4_M55_noxref_d ) capacitor c=6.94454e-19 \
 //x=11.47 //y=7.4 //x2=9.225 //y2=5.02
cc_996 ( N_VDD_M56_noxref_d N_noxref_4_M55_noxref_d ) capacitor c=0.0664752f \
 //x=9.665 //y=5.02 //x2=9.225 //y2=5.02
cc_997 ( N_VDD_c_960_p N_noxref_4_M57_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=10.105 //y2=5.02
cc_998 ( N_VDD_c_997_p N_noxref_4_M57_noxref_d ) capacitor c=0.0140317f \
 //x=10.605 //y=7.4 //x2=10.105 //y2=5.02
cc_999 ( N_VDD_c_941_n N_noxref_4_M57_noxref_d ) capacitor c=0.0120541f \
 //x=11.47 //y=7.4 //x2=10.105 //y2=5.02
cc_1000 ( N_VDD_M55_noxref_s N_noxref_4_M57_noxref_d ) capacitor c=0.00111971f \
 //x=8.795 //y=5.02 //x2=10.105 //y2=5.02
cc_1001 ( N_VDD_M56_noxref_d N_noxref_4_M57_noxref_d ) capacitor c=0.0664752f \
 //x=9.665 //y=5.02 //x2=10.105 //y2=5.02
cc_1002 ( N_VDD_M58_noxref_d N_noxref_4_M57_noxref_d ) capacitor c=0.0664752f \
 //x=10.545 //y=5.02 //x2=10.105 //y2=5.02
cc_1003 ( N_VDD_M59_noxref_s N_noxref_4_M57_noxref_d ) capacitor c=4.54516e-19 \
 //x=12.125 //y=5.02 //x2=10.105 //y2=5.02
cc_1004 ( N_VDD_c_960_p N_noxref_5_c_2342_n ) capacitor c=0.00449316f \
 //x=73.63 //y=7.4 //x2=2.325 //y2=5.155
cc_1005 ( N_VDD_c_1027_p N_noxref_5_c_2342_n ) capacitor c=4.32228e-19 \
 //x=1.885 //y=7.4 //x2=2.325 //y2=5.155
cc_1006 ( N_VDD_c_1028_p N_noxref_5_c_2342_n ) capacitor c=4.31906e-19 \
 //x=2.765 //y=7.4 //x2=2.325 //y2=5.155
cc_1007 ( N_VDD_M46_noxref_d N_noxref_5_c_2342_n ) capacitor c=0.0115147f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_1008 ( N_VDD_c_937_n N_noxref_5_c_2346_n ) capacitor c=0.00880189f //x=0.74 \
 //y=7.4 //x2=1.615 //y2=5.155
cc_1009 ( N_VDD_M45_noxref_s N_noxref_5_c_2346_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_1010 ( N_VDD_c_960_p N_noxref_5_c_2348_n ) capacitor c=0.0044221f //x=73.63 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_1011 ( N_VDD_c_1028_p N_noxref_5_c_2348_n ) capacitor c=4.31931e-19 \
 //x=2.765 //y=7.4 //x2=3.205 //y2=5.155
cc_1012 ( N_VDD_c_975_p N_noxref_5_c_2348_n ) capacitor c=4.31931e-19 \
 //x=3.645 //y=7.4 //x2=3.205 //y2=5.155
cc_1013 ( N_VDD_M48_noxref_d N_noxref_5_c_2348_n ) capacitor c=0.0112985f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_1014 ( N_VDD_c_960_p N_noxref_5_c_2352_n ) capacitor c=0.00434174f \
 //x=73.63 //y=7.4 //x2=3.985 //y2=5.155
cc_1015 ( N_VDD_c_975_p N_noxref_5_c_2352_n ) capacitor c=7.46626e-19 \
 //x=3.645 //y=7.4 //x2=3.985 //y2=5.155
cc_1016 ( N_VDD_c_1038_p N_noxref_5_c_2352_n ) capacitor c=0.00198565f \
 //x=4.64 //y=7.4 //x2=3.985 //y2=5.155
cc_1017 ( N_VDD_M50_noxref_d N_noxref_5_c_2352_n ) capacitor c=0.0112985f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_1018 ( N_VDD_c_939_n N_noxref_5_c_2356_n ) capacitor c=0.0426341f //x=4.81 \
 //y=7.4 //x2=4.07 //y2=3.7
cc_1019 ( N_VDD_c_960_p N_noxref_5_c_2319_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=5.92 //y2=2.08
cc_1020 ( N_VDD_c_961_p N_noxref_5_c_2319_n ) capacitor c=2.87256e-19 \
 //x=6.395 //y=7.4 //x2=5.92 //y2=2.08
cc_1021 ( N_VDD_c_939_n N_noxref_5_c_2319_n ) capacitor c=0.0134665f //x=4.81 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_1022 ( N_VDD_c_960_p N_noxref_5_c_2320_n ) capacitor c=0.00125292f \
 //x=73.63 //y=7.4 //x2=15.91 //y2=2.08
cc_1023 ( N_VDD_c_1045_p N_noxref_5_c_2320_n ) capacitor c=2.87264e-19 \
 //x=16.385 //y=7.4 //x2=15.91 //y2=2.08
cc_1024 ( N_VDD_c_942_n N_noxref_5_c_2320_n ) capacitor c=0.0135534f //x=14.8 \
 //y=7.4 //x2=15.91 //y2=2.08
cc_1025 ( N_VDD_c_961_p N_noxref_5_M51_noxref_g ) capacitor c=0.00726866f \
 //x=6.395 //y=7.4 //x2=5.82 //y2=6.02
cc_1026 ( N_VDD_M51_noxref_s N_noxref_5_M51_noxref_g ) capacitor c=0.054195f \
 //x=5.465 //y=5.02 //x2=5.82 //y2=6.02
cc_1027 ( N_VDD_c_961_p N_noxref_5_M52_noxref_g ) capacitor c=0.00672952f \
 //x=6.395 //y=7.4 //x2=6.26 //y2=6.02
cc_1028 ( N_VDD_M52_noxref_d N_noxref_5_M52_noxref_g ) capacitor c=0.015318f \
 //x=6.335 //y=5.02 //x2=6.26 //y2=6.02
cc_1029 ( N_VDD_c_1045_p N_noxref_5_M63_noxref_g ) capacitor c=0.00726866f \
 //x=16.385 //y=7.4 //x2=15.81 //y2=6.02
cc_1030 ( N_VDD_M63_noxref_s N_noxref_5_M63_noxref_g ) capacitor c=0.054195f \
 //x=15.455 //y=5.02 //x2=15.81 //y2=6.02
cc_1031 ( N_VDD_c_1045_p N_noxref_5_M64_noxref_g ) capacitor c=0.00672952f \
 //x=16.385 //y=7.4 //x2=16.25 //y2=6.02
cc_1032 ( N_VDD_M64_noxref_d N_noxref_5_M64_noxref_g ) capacitor c=0.015318f \
 //x=16.325 //y=5.02 //x2=16.25 //y2=6.02
cc_1033 ( N_VDD_c_939_n N_noxref_5_c_2371_n ) capacitor c=0.015293f //x=4.81 \
 //y=7.4 //x2=5.92 //y2=4.7
cc_1034 ( N_VDD_c_942_n N_noxref_5_c_2372_n ) capacitor c=0.0149273f //x=14.8 \
 //y=7.4 //x2=15.91 //y2=4.7
cc_1035 ( N_VDD_c_960_p N_noxref_5_M45_noxref_d ) capacitor c=0.00285091f \
 //x=73.63 //y=7.4 //x2=1.385 //y2=5.02
cc_1036 ( N_VDD_c_1027_p N_noxref_5_M45_noxref_d ) capacitor c=0.0141016f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_1037 ( N_VDD_M46_noxref_d N_noxref_5_M45_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_1038 ( N_VDD_c_960_p N_noxref_5_M47_noxref_d ) capacitor c=0.00275186f \
 //x=73.63 //y=7.4 //x2=2.265 //y2=5.02
cc_1039 ( N_VDD_c_1028_p N_noxref_5_M47_noxref_d ) capacitor c=0.0140346f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_1040 ( N_VDD_c_939_n N_noxref_5_M47_noxref_d ) capacitor c=4.9285e-19 \
 //x=4.81 //y=7.4 //x2=2.265 //y2=5.02
cc_1041 ( N_VDD_M45_noxref_s N_noxref_5_M47_noxref_d ) capacitor c=0.00130656f \
 //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_1042 ( N_VDD_M46_noxref_d N_noxref_5_M47_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_1043 ( N_VDD_M48_noxref_d N_noxref_5_M47_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_1044 ( N_VDD_c_960_p N_noxref_5_M49_noxref_d ) capacitor c=0.00275235f \
 //x=73.63 //y=7.4 //x2=3.145 //y2=5.02
cc_1045 ( N_VDD_c_975_p N_noxref_5_M49_noxref_d ) capacitor c=0.0137384f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_1046 ( N_VDD_c_939_n N_noxref_5_M49_noxref_d ) capacitor c=0.00939849f \
 //x=4.81 //y=7.4 //x2=3.145 //y2=5.02
cc_1047 ( N_VDD_M48_noxref_d N_noxref_5_M49_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_1048 ( N_VDD_M50_noxref_d N_noxref_5_M49_noxref_d ) capacitor c=0.0664752f \
 //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_1049 ( N_VDD_M51_noxref_s N_noxref_5_M49_noxref_d ) capacitor c=4.52683e-19 \
 //x=5.465 //y=5.02 //x2=3.145 //y2=5.02
cc_1050 ( N_VDD_c_960_p N_noxref_6_c_2581_n ) capacitor c=0.00453752f \
 //x=73.63 //y=7.4 //x2=16.825 //y2=5.2
cc_1051 ( N_VDD_c_1045_p N_noxref_6_c_2581_n ) capacitor c=4.48395e-19 \
 //x=16.385 //y=7.4 //x2=16.825 //y2=5.2
cc_1052 ( N_VDD_c_1074_p N_noxref_6_c_2581_n ) capacitor c=4.48393e-19 \
 //x=17.265 //y=7.4 //x2=16.825 //y2=5.2
cc_1053 ( N_VDD_M64_noxref_d N_noxref_6_c_2581_n ) capacitor c=0.0124581f \
 //x=16.325 //y=5.02 //x2=16.825 //y2=5.2
cc_1054 ( N_VDD_c_942_n N_noxref_6_c_2585_n ) capacitor c=0.00985474f //x=14.8 \
 //y=7.4 //x2=16.115 //y2=5.2
cc_1055 ( N_VDD_M63_noxref_s N_noxref_6_c_2585_n ) capacitor c=0.087833f \
 //x=15.455 //y=5.02 //x2=16.115 //y2=5.2
cc_1056 ( N_VDD_c_960_p N_noxref_6_c_2587_n ) capacitor c=0.00301575f \
 //x=73.63 //y=7.4 //x2=17.305 //y2=5.2
cc_1057 ( N_VDD_c_1074_p N_noxref_6_c_2587_n ) capacitor c=7.72068e-19 \
 //x=17.265 //y=7.4 //x2=17.305 //y2=5.2
cc_1058 ( N_VDD_M66_noxref_d N_noxref_6_c_2587_n ) capacitor c=0.0158515f \
 //x=17.205 //y=5.02 //x2=17.305 //y2=5.2
cc_1059 ( N_VDD_M67_noxref_s N_noxref_6_c_2587_n ) capacitor c=2.44532e-19 \
 //x=18.785 //y=5.02 //x2=17.305 //y2=5.2
cc_1060 ( N_VDD_c_942_n N_noxref_6_c_2566_n ) capacitor c=0.00151618f //x=14.8 \
 //y=7.4 //x2=17.39 //y2=3.7
cc_1061 ( N_VDD_c_943_n N_noxref_6_c_2566_n ) capacitor c=0.0429414f //x=18.13 \
 //y=7.4 //x2=17.39 //y2=3.7
cc_1062 ( N_VDD_c_960_p N_noxref_6_c_2567_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=19.24 //y2=2.08
cc_1063 ( N_VDD_c_1085_p N_noxref_6_c_2567_n ) capacitor c=2.87256e-19 \
 //x=19.715 //y=7.4 //x2=19.24 //y2=2.08
cc_1064 ( N_VDD_c_943_n N_noxref_6_c_2567_n ) capacitor c=0.0134208f //x=18.13 \
 //y=7.4 //x2=19.24 //y2=2.08
cc_1065 ( N_VDD_c_1085_p N_noxref_6_M67_noxref_g ) capacitor c=0.00726866f \
 //x=19.715 //y=7.4 //x2=19.14 //y2=6.02
cc_1066 ( N_VDD_M67_noxref_s N_noxref_6_M67_noxref_g ) capacitor c=0.054195f \
 //x=18.785 //y=5.02 //x2=19.14 //y2=6.02
cc_1067 ( N_VDD_c_1085_p N_noxref_6_M68_noxref_g ) capacitor c=0.00672952f \
 //x=19.715 //y=7.4 //x2=19.58 //y2=6.02
cc_1068 ( N_VDD_M68_noxref_d N_noxref_6_M68_noxref_g ) capacitor c=0.015318f \
 //x=19.655 //y=5.02 //x2=19.58 //y2=6.02
cc_1069 ( N_VDD_c_943_n N_noxref_6_c_2600_n ) capacitor c=0.0150435f //x=18.13 \
 //y=7.4 //x2=19.24 //y2=4.7
cc_1070 ( N_VDD_c_960_p N_noxref_6_M63_noxref_d ) capacitor c=0.00275364f \
 //x=73.63 //y=7.4 //x2=15.885 //y2=5.02
cc_1071 ( N_VDD_c_1045_p N_noxref_6_M63_noxref_d ) capacitor c=0.0140327f \
 //x=16.385 //y=7.4 //x2=15.885 //y2=5.02
cc_1072 ( N_VDD_c_943_n N_noxref_6_M63_noxref_d ) capacitor c=6.94454e-19 \
 //x=18.13 //y=7.4 //x2=15.885 //y2=5.02
cc_1073 ( N_VDD_M64_noxref_d N_noxref_6_M63_noxref_d ) capacitor c=0.0664752f \
 //x=16.325 //y=5.02 //x2=15.885 //y2=5.02
cc_1074 ( N_VDD_c_960_p N_noxref_6_M65_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=16.765 //y2=5.02
cc_1075 ( N_VDD_c_1074_p N_noxref_6_M65_noxref_d ) capacitor c=0.0140317f \
 //x=17.265 //y=7.4 //x2=16.765 //y2=5.02
cc_1076 ( N_VDD_c_943_n N_noxref_6_M65_noxref_d ) capacitor c=0.0120541f \
 //x=18.13 //y=7.4 //x2=16.765 //y2=5.02
cc_1077 ( N_VDD_M63_noxref_s N_noxref_6_M65_noxref_d ) capacitor c=0.00111971f \
 //x=15.455 //y=5.02 //x2=16.765 //y2=5.02
cc_1078 ( N_VDD_M64_noxref_d N_noxref_6_M65_noxref_d ) capacitor c=0.0664752f \
 //x=16.325 //y=5.02 //x2=16.765 //y2=5.02
cc_1079 ( N_VDD_M66_noxref_d N_noxref_6_M65_noxref_d ) capacitor c=0.0664752f \
 //x=17.205 //y=5.02 //x2=16.765 //y2=5.02
cc_1080 ( N_VDD_M67_noxref_s N_noxref_6_M65_noxref_d ) capacitor c=4.54516e-19 \
 //x=18.785 //y=5.02 //x2=16.765 //y2=5.02
cc_1081 ( N_VDD_c_960_p N_noxref_7_c_2715_n ) capacitor c=0.035625f //x=73.63 \
 //y=7.4 //x2=9.875 //y2=4.07
cc_1082 ( N_VDD_c_1027_p N_noxref_7_c_2715_n ) capacitor c=0.00113322f \
 //x=1.885 //y=7.4 //x2=9.875 //y2=4.07
cc_1083 ( N_VDD_c_939_n N_noxref_7_c_2715_n ) capacitor c=0.0140578f //x=4.81 \
 //y=7.4 //x2=9.875 //y2=4.07
cc_1084 ( N_VDD_c_940_n N_noxref_7_c_2715_n ) capacitor c=0.0140578f //x=8.14 \
 //y=7.4 //x2=9.875 //y2=4.07
cc_1085 ( N_VDD_c_960_p N_noxref_7_c_2716_n ) capacitor c=0.00189266f \
 //x=73.63 //y=7.4 //x2=1.225 //y2=4.07
cc_1086 ( N_VDD_c_937_n N_noxref_7_c_2716_n ) capacitor c=0.0017219f //x=0.74 \
 //y=7.4 //x2=1.225 //y2=4.07
cc_1087 ( N_VDD_M45_noxref_s N_noxref_7_c_2716_n ) capacitor c=0.00128242f \
 //x=0.955 //y=5.02 //x2=1.225 //y2=4.07
cc_1088 ( N_VDD_c_941_n N_noxref_7_c_2744_n ) capacitor c=0.0140578f //x=11.47 \
 //y=7.4 //x2=13.945 //y2=4.07
cc_1089 ( N_VDD_c_942_n N_noxref_7_c_2745_n ) capacitor c=0.0142127f //x=14.8 \
 //y=7.4 //x2=19.865 //y2=4.07
cc_1090 ( N_VDD_c_943_n N_noxref_7_c_2745_n ) capacitor c=0.0140578f //x=18.13 \
 //y=7.4 //x2=19.865 //y2=4.07
cc_1091 ( N_VDD_c_942_n N_noxref_7_c_2747_n ) capacitor c=0.00104972f //x=14.8 \
 //y=7.4 //x2=14.175 //y2=4.07
cc_1092 ( N_VDD_c_960_p N_noxref_7_c_2717_n ) capacitor c=9.2251e-19 //x=73.63 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_1093 ( N_VDD_c_937_n N_noxref_7_c_2717_n ) capacitor c=0.0159723f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_1094 ( N_VDD_M45_noxref_s N_noxref_7_c_2717_n ) capacitor c=0.0122951f \
 //x=0.955 //y=5.02 //x2=1.11 //y2=2.08
cc_1095 ( N_VDD_c_940_n N_noxref_7_c_2718_n ) capacitor c=4.57806e-19 //x=8.14 \
 //y=7.4 //x2=9.99 //y2=2.08
cc_1096 ( N_VDD_c_941_n N_noxref_7_c_2718_n ) capacitor c=3.69525e-19 \
 //x=11.47 //y=7.4 //x2=9.99 //y2=2.08
cc_1097 ( N_VDD_c_960_p N_noxref_7_c_2753_n ) capacitor c=0.00453473f \
 //x=73.63 //y=7.4 //x2=13.495 //y2=5.2
cc_1098 ( N_VDD_c_1008_p N_noxref_7_c_2753_n ) capacitor c=4.48391e-19 \
 //x=13.055 //y=7.4 //x2=13.495 //y2=5.2
cc_1099 ( N_VDD_c_1121_p N_noxref_7_c_2753_n ) capacitor c=4.48377e-19 \
 //x=13.935 //y=7.4 //x2=13.495 //y2=5.2
cc_1100 ( N_VDD_M60_noxref_d N_noxref_7_c_2753_n ) capacitor c=0.0124506f \
 //x=12.995 //y=5.02 //x2=13.495 //y2=5.2
cc_1101 ( N_VDD_c_941_n N_noxref_7_c_2757_n ) capacitor c=0.00985474f \
 //x=11.47 //y=7.4 //x2=12.785 //y2=5.2
cc_1102 ( N_VDD_M59_noxref_s N_noxref_7_c_2757_n ) capacitor c=0.087833f \
 //x=12.125 //y=5.02 //x2=12.785 //y2=5.2
cc_1103 ( N_VDD_c_960_p N_noxref_7_c_2759_n ) capacitor c=0.00301658f \
 //x=73.63 //y=7.4 //x2=13.975 //y2=5.2
cc_1104 ( N_VDD_c_1121_p N_noxref_7_c_2759_n ) capacitor c=7.72084e-19 \
 //x=13.935 //y=7.4 //x2=13.975 //y2=5.2
cc_1105 ( N_VDD_M62_noxref_d N_noxref_7_c_2759_n ) capacitor c=0.0158564f \
 //x=13.875 //y=5.02 //x2=13.975 //y2=5.2
cc_1106 ( N_VDD_M63_noxref_s N_noxref_7_c_2759_n ) capacitor c=2.44532e-19 \
 //x=15.455 //y=5.02 //x2=13.975 //y2=5.2
cc_1107 ( N_VDD_c_941_n N_noxref_7_c_2721_n ) capacitor c=0.00151618f \
 //x=11.47 //y=7.4 //x2=14.06 //y2=4.07
cc_1108 ( N_VDD_c_942_n N_noxref_7_c_2721_n ) capacitor c=0.0432014f //x=14.8 \
 //y=7.4 //x2=14.06 //y2=4.07
cc_1109 ( N_VDD_c_943_n N_noxref_7_c_2722_n ) capacitor c=4.57806e-19 \
 //x=18.13 //y=7.4 //x2=19.98 //y2=2.08
cc_1110 ( N_VDD_c_944_n N_noxref_7_c_2722_n ) capacitor c=4.17938e-19 \
 //x=21.46 //y=7.4 //x2=19.98 //y2=2.08
cc_1111 ( N_VDD_c_1027_p N_noxref_7_M45_noxref_g ) capacitor c=0.00749687f \
 //x=1.885 //y=7.4 //x2=1.31 //y2=6.02
cc_1112 ( N_VDD_M45_noxref_s N_noxref_7_M45_noxref_g ) capacitor c=0.0477201f \
 //x=0.955 //y=5.02 //x2=1.31 //y2=6.02
cc_1113 ( N_VDD_c_1027_p N_noxref_7_M46_noxref_g ) capacitor c=0.00675175f \
 //x=1.885 //y=7.4 //x2=1.75 //y2=6.02
cc_1114 ( N_VDD_M46_noxref_d N_noxref_7_M46_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=1.75 //y2=6.02
cc_1115 ( N_VDD_c_997_p N_noxref_7_M57_noxref_g ) capacitor c=0.00673971f \
 //x=10.605 //y=7.4 //x2=10.03 //y2=6.02
cc_1116 ( N_VDD_M56_noxref_d N_noxref_7_M57_noxref_g ) capacitor c=0.015318f \
 //x=9.665 //y=5.02 //x2=10.03 //y2=6.02
cc_1117 ( N_VDD_c_997_p N_noxref_7_M58_noxref_g ) capacitor c=0.00672952f \
 //x=10.605 //y=7.4 //x2=10.47 //y2=6.02
cc_1118 ( N_VDD_c_941_n N_noxref_7_M58_noxref_g ) capacitor c=0.00864163f \
 //x=11.47 //y=7.4 //x2=10.47 //y2=6.02
cc_1119 ( N_VDD_M58_noxref_d N_noxref_7_M58_noxref_g ) capacitor c=0.0430452f \
 //x=10.545 //y=5.02 //x2=10.47 //y2=6.02
cc_1120 ( N_VDD_c_1142_p N_noxref_7_M69_noxref_g ) capacitor c=0.00673971f \
 //x=20.595 //y=7.4 //x2=20.02 //y2=6.02
cc_1121 ( N_VDD_M68_noxref_d N_noxref_7_M69_noxref_g ) capacitor c=0.015318f \
 //x=19.655 //y=5.02 //x2=20.02 //y2=6.02
cc_1122 ( N_VDD_c_1142_p N_noxref_7_M70_noxref_g ) capacitor c=0.00672952f \
 //x=20.595 //y=7.4 //x2=20.46 //y2=6.02
cc_1123 ( N_VDD_c_944_n N_noxref_7_M70_noxref_g ) capacitor c=0.00928743f \
 //x=21.46 //y=7.4 //x2=20.46 //y2=6.02
cc_1124 ( N_VDD_M70_noxref_d N_noxref_7_M70_noxref_g ) capacitor c=0.0430452f \
 //x=20.535 //y=5.02 //x2=20.46 //y2=6.02
cc_1125 ( N_VDD_c_937_n N_noxref_7_c_2781_n ) capacitor c=0.00757682f //x=0.74 \
 //y=7.4 //x2=1.385 //y2=4.79
cc_1126 ( N_VDD_M45_noxref_s N_noxref_7_c_2781_n ) capacitor c=0.00445117f \
 //x=0.955 //y=5.02 //x2=1.385 //y2=4.79
cc_1127 ( N_VDD_c_960_p N_noxref_7_M59_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=12.555 //y2=5.02
cc_1128 ( N_VDD_c_1008_p N_noxref_7_M59_noxref_d ) capacitor c=0.0140317f \
 //x=13.055 //y=7.4 //x2=12.555 //y2=5.02
cc_1129 ( N_VDD_c_942_n N_noxref_7_M59_noxref_d ) capacitor c=6.94454e-19 \
 //x=14.8 //y=7.4 //x2=12.555 //y2=5.02
cc_1130 ( N_VDD_M60_noxref_d N_noxref_7_M59_noxref_d ) capacitor c=0.0664752f \
 //x=12.995 //y=5.02 //x2=12.555 //y2=5.02
cc_1131 ( N_VDD_c_960_p N_noxref_7_M61_noxref_d ) capacitor c=0.00275364f \
 //x=73.63 //y=7.4 //x2=13.435 //y2=5.02
cc_1132 ( N_VDD_c_1121_p N_noxref_7_M61_noxref_d ) capacitor c=0.0140327f \
 //x=13.935 //y=7.4 //x2=13.435 //y2=5.02
cc_1133 ( N_VDD_c_942_n N_noxref_7_M61_noxref_d ) capacitor c=0.0120541f \
 //x=14.8 //y=7.4 //x2=13.435 //y2=5.02
cc_1134 ( N_VDD_M59_noxref_s N_noxref_7_M61_noxref_d ) capacitor c=0.00111971f \
 //x=12.125 //y=5.02 //x2=13.435 //y2=5.02
cc_1135 ( N_VDD_M60_noxref_d N_noxref_7_M61_noxref_d ) capacitor c=0.0664752f \
 //x=12.995 //y=5.02 //x2=13.435 //y2=5.02
cc_1136 ( N_VDD_M62_noxref_d N_noxref_7_M61_noxref_d ) capacitor c=0.0664752f \
 //x=13.875 //y=5.02 //x2=13.435 //y2=5.02
cc_1137 ( N_VDD_M63_noxref_s N_noxref_7_M61_noxref_d ) capacitor c=4.54516e-19 \
 //x=15.455 //y=5.02 //x2=13.435 //y2=5.02
cc_1138 ( N_VDD_c_945_n N_noxref_8_c_3068_n ) capacitor c=6.58823e-19 \
 //x=26.27 //y=7.4 //x2=24.79 //y2=2.08
cc_1139 ( N_VDD_c_960_p N_noxref_8_c_3086_n ) capacitor c=0.00453663f \
 //x=73.63 //y=7.4 //x2=28.295 //y2=5.2
cc_1140 ( N_VDD_c_1162_p N_noxref_8_c_3086_n ) capacitor c=4.48391e-19 \
 //x=27.855 //y=7.4 //x2=28.295 //y2=5.2
cc_1141 ( N_VDD_c_1163_p N_noxref_8_c_3086_n ) capacitor c=4.48391e-19 \
 //x=28.735 //y=7.4 //x2=28.295 //y2=5.2
cc_1142 ( N_VDD_M78_noxref_d N_noxref_8_c_3086_n ) capacitor c=0.0124542f \
 //x=27.795 //y=5.02 //x2=28.295 //y2=5.2
cc_1143 ( N_VDD_c_945_n N_noxref_8_c_3090_n ) capacitor c=0.00985474f \
 //x=26.27 //y=7.4 //x2=27.585 //y2=5.2
cc_1144 ( N_VDD_M77_noxref_s N_noxref_8_c_3090_n ) capacitor c=0.087833f \
 //x=26.925 //y=5.02 //x2=27.585 //y2=5.2
cc_1145 ( N_VDD_c_960_p N_noxref_8_c_3092_n ) capacitor c=0.00301575f \
 //x=73.63 //y=7.4 //x2=28.775 //y2=5.2
cc_1146 ( N_VDD_c_1163_p N_noxref_8_c_3092_n ) capacitor c=7.72068e-19 \
 //x=28.735 //y=7.4 //x2=28.775 //y2=5.2
cc_1147 ( N_VDD_M80_noxref_d N_noxref_8_c_3092_n ) capacitor c=0.0158515f \
 //x=28.675 //y=5.02 //x2=28.775 //y2=5.2
cc_1148 ( N_VDD_M81_noxref_s N_noxref_8_c_3092_n ) capacitor c=2.44532e-19 \
 //x=30.255 //y=5.02 //x2=28.775 //y2=5.2
cc_1149 ( N_VDD_c_945_n N_noxref_8_c_3070_n ) capacitor c=0.00151618f \
 //x=26.27 //y=7.4 //x2=28.86 //y2=3.33
cc_1150 ( N_VDD_c_946_n N_noxref_8_c_3070_n ) capacitor c=0.0429414f //x=29.6 \
 //y=7.4 //x2=28.86 //y2=3.33
cc_1151 ( N_VDD_c_960_p N_noxref_8_c_3071_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=30.71 //y2=2.08
cc_1152 ( N_VDD_c_1174_p N_noxref_8_c_3071_n ) capacitor c=2.87256e-19 \
 //x=31.185 //y=7.4 //x2=30.71 //y2=2.08
cc_1153 ( N_VDD_c_946_n N_noxref_8_c_3071_n ) capacitor c=0.0134208f //x=29.6 \
 //y=7.4 //x2=30.71 //y2=2.08
cc_1154 ( N_VDD_c_1176_p N_noxref_8_M75_noxref_g ) capacitor c=0.00675175f \
 //x=25.105 //y=7.4 //x2=24.53 //y2=6.02
cc_1155 ( N_VDD_M74_noxref_d N_noxref_8_M75_noxref_g ) capacitor c=0.015318f \
 //x=24.165 //y=5.02 //x2=24.53 //y2=6.02
cc_1156 ( N_VDD_c_1176_p N_noxref_8_M76_noxref_g ) capacitor c=0.00675379f \
 //x=25.105 //y=7.4 //x2=24.97 //y2=6.02
cc_1157 ( N_VDD_M76_noxref_d N_noxref_8_M76_noxref_g ) capacitor c=0.0394719f \
 //x=25.045 //y=5.02 //x2=24.97 //y2=6.02
cc_1158 ( N_VDD_c_1174_p N_noxref_8_M81_noxref_g ) capacitor c=0.00726866f \
 //x=31.185 //y=7.4 //x2=30.61 //y2=6.02
cc_1159 ( N_VDD_M81_noxref_s N_noxref_8_M81_noxref_g ) capacitor c=0.054195f \
 //x=30.255 //y=5.02 //x2=30.61 //y2=6.02
cc_1160 ( N_VDD_c_1174_p N_noxref_8_M82_noxref_g ) capacitor c=0.00672952f \
 //x=31.185 //y=7.4 //x2=31.05 //y2=6.02
cc_1161 ( N_VDD_M82_noxref_d N_noxref_8_M82_noxref_g ) capacitor c=0.015318f \
 //x=31.125 //y=5.02 //x2=31.05 //y2=6.02
cc_1162 ( N_VDD_c_946_n N_noxref_8_c_3109_n ) capacitor c=0.0150435f //x=29.6 \
 //y=7.4 //x2=30.71 //y2=4.7
cc_1163 ( N_VDD_c_960_p N_noxref_8_M77_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=27.355 //y2=5.02
cc_1164 ( N_VDD_c_1162_p N_noxref_8_M77_noxref_d ) capacitor c=0.0140317f \
 //x=27.855 //y=7.4 //x2=27.355 //y2=5.02
cc_1165 ( N_VDD_c_946_n N_noxref_8_M77_noxref_d ) capacitor c=6.94454e-19 \
 //x=29.6 //y=7.4 //x2=27.355 //y2=5.02
cc_1166 ( N_VDD_M78_noxref_d N_noxref_8_M77_noxref_d ) capacitor c=0.0664752f \
 //x=27.795 //y=5.02 //x2=27.355 //y2=5.02
cc_1167 ( N_VDD_c_960_p N_noxref_8_M79_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=28.235 //y2=5.02
cc_1168 ( N_VDD_c_1163_p N_noxref_8_M79_noxref_d ) capacitor c=0.0140317f \
 //x=28.735 //y=7.4 //x2=28.235 //y2=5.02
cc_1169 ( N_VDD_c_946_n N_noxref_8_M79_noxref_d ) capacitor c=0.0120541f \
 //x=29.6 //y=7.4 //x2=28.235 //y2=5.02
cc_1170 ( N_VDD_M77_noxref_s N_noxref_8_M79_noxref_d ) capacitor c=0.00111971f \
 //x=26.925 //y=5.02 //x2=28.235 //y2=5.02
cc_1171 ( N_VDD_M78_noxref_d N_noxref_8_M79_noxref_d ) capacitor c=0.0664752f \
 //x=27.795 //y=5.02 //x2=28.235 //y2=5.02
cc_1172 ( N_VDD_M80_noxref_d N_noxref_8_M79_noxref_d ) capacitor c=0.0664752f \
 //x=28.675 //y=5.02 //x2=28.235 //y2=5.02
cc_1173 ( N_VDD_M81_noxref_s N_noxref_8_M79_noxref_d ) capacitor c=4.54516e-19 \
 //x=30.255 //y=5.02 //x2=28.235 //y2=5.02
cc_1174 ( N_VDD_c_960_p N_noxref_9_c_3316_n ) capacitor c=0.00453663f \
 //x=73.63 //y=7.4 //x2=31.625 //y2=5.2
cc_1175 ( N_VDD_c_1174_p N_noxref_9_c_3316_n ) capacitor c=4.48391e-19 \
 //x=31.185 //y=7.4 //x2=31.625 //y2=5.2
cc_1176 ( N_VDD_c_1198_p N_noxref_9_c_3316_n ) capacitor c=4.48391e-19 \
 //x=32.065 //y=7.4 //x2=31.625 //y2=5.2
cc_1177 ( N_VDD_M82_noxref_d N_noxref_9_c_3316_n ) capacitor c=0.0124542f \
 //x=31.125 //y=5.02 //x2=31.625 //y2=5.2
cc_1178 ( N_VDD_c_946_n N_noxref_9_c_3320_n ) capacitor c=0.00985474f //x=29.6 \
 //y=7.4 //x2=30.915 //y2=5.2
cc_1179 ( N_VDD_M81_noxref_s N_noxref_9_c_3320_n ) capacitor c=0.087833f \
 //x=30.255 //y=5.02 //x2=30.915 //y2=5.2
cc_1180 ( N_VDD_c_960_p N_noxref_9_c_3322_n ) capacitor c=0.00301575f \
 //x=73.63 //y=7.4 //x2=32.105 //y2=5.2
cc_1181 ( N_VDD_c_1198_p N_noxref_9_c_3322_n ) capacitor c=7.72068e-19 \
 //x=32.065 //y=7.4 //x2=32.105 //y2=5.2
cc_1182 ( N_VDD_M84_noxref_d N_noxref_9_c_3322_n ) capacitor c=0.0158515f \
 //x=32.005 //y=5.02 //x2=32.105 //y2=5.2
cc_1183 ( N_VDD_M85_noxref_s N_noxref_9_c_3322_n ) capacitor c=2.44532e-19 \
 //x=33.585 //y=5.02 //x2=32.105 //y2=5.2
cc_1184 ( N_VDD_c_946_n N_noxref_9_c_3301_n ) capacitor c=0.00151618f //x=29.6 \
 //y=7.4 //x2=32.19 //y2=3.33
cc_1185 ( N_VDD_c_947_n N_noxref_9_c_3301_n ) capacitor c=0.0427674f //x=32.93 \
 //y=7.4 //x2=32.19 //y2=3.33
cc_1186 ( N_VDD_c_960_p N_noxref_9_c_3302_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=34.04 //y2=2.08
cc_1187 ( N_VDD_c_1209_p N_noxref_9_c_3302_n ) capacitor c=2.87256e-19 \
 //x=34.515 //y=7.4 //x2=34.04 //y2=2.08
cc_1188 ( N_VDD_c_947_n N_noxref_9_c_3302_n ) capacitor c=0.0133228f //x=32.93 \
 //y=7.4 //x2=34.04 //y2=2.08
cc_1189 ( N_VDD_c_1209_p N_noxref_9_M85_noxref_g ) capacitor c=0.00726866f \
 //x=34.515 //y=7.4 //x2=33.94 //y2=6.02
cc_1190 ( N_VDD_M85_noxref_s N_noxref_9_M85_noxref_g ) capacitor c=0.054195f \
 //x=33.585 //y=5.02 //x2=33.94 //y2=6.02
cc_1191 ( N_VDD_c_1209_p N_noxref_9_M86_noxref_g ) capacitor c=0.00672952f \
 //x=34.515 //y=7.4 //x2=34.38 //y2=6.02
cc_1192 ( N_VDD_M86_noxref_d N_noxref_9_M86_noxref_g ) capacitor c=0.015318f \
 //x=34.455 //y=5.02 //x2=34.38 //y2=6.02
cc_1193 ( N_VDD_c_947_n N_noxref_9_c_3335_n ) capacitor c=0.0149273f //x=32.93 \
 //y=7.4 //x2=34.04 //y2=4.7
cc_1194 ( N_VDD_c_960_p N_noxref_9_M81_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=30.685 //y2=5.02
cc_1195 ( N_VDD_c_1174_p N_noxref_9_M81_noxref_d ) capacitor c=0.0140317f \
 //x=31.185 //y=7.4 //x2=30.685 //y2=5.02
cc_1196 ( N_VDD_c_947_n N_noxref_9_M81_noxref_d ) capacitor c=6.94454e-19 \
 //x=32.93 //y=7.4 //x2=30.685 //y2=5.02
cc_1197 ( N_VDD_M82_noxref_d N_noxref_9_M81_noxref_d ) capacitor c=0.0664752f \
 //x=31.125 //y=5.02 //x2=30.685 //y2=5.02
cc_1198 ( N_VDD_c_960_p N_noxref_9_M83_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=31.565 //y2=5.02
cc_1199 ( N_VDD_c_1198_p N_noxref_9_M83_noxref_d ) capacitor c=0.0140317f \
 //x=32.065 //y=7.4 //x2=31.565 //y2=5.02
cc_1200 ( N_VDD_c_947_n N_noxref_9_M83_noxref_d ) capacitor c=0.0120541f \
 //x=32.93 //y=7.4 //x2=31.565 //y2=5.02
cc_1201 ( N_VDD_M81_noxref_s N_noxref_9_M83_noxref_d ) capacitor c=0.00111971f \
 //x=30.255 //y=5.02 //x2=31.565 //y2=5.02
cc_1202 ( N_VDD_M82_noxref_d N_noxref_9_M83_noxref_d ) capacitor c=0.0664752f \
 //x=31.125 //y=5.02 //x2=31.565 //y2=5.02
cc_1203 ( N_VDD_M84_noxref_d N_noxref_9_M83_noxref_d ) capacitor c=0.0664752f \
 //x=32.005 //y=5.02 //x2=31.565 //y2=5.02
cc_1204 ( N_VDD_M85_noxref_s N_noxref_9_M83_noxref_d ) capacitor c=4.54516e-19 \
 //x=33.585 //y=5.02 //x2=31.565 //y2=5.02
cc_1205 ( N_VDD_c_960_p N_noxref_10_c_3477_n ) capacitor c=0.00444751f \
 //x=73.63 //y=7.4 //x2=23.785 //y2=5.155
cc_1206 ( N_VDD_c_1228_p N_noxref_10_c_3477_n ) capacitor c=4.31931e-19 \
 //x=23.345 //y=7.4 //x2=23.785 //y2=5.155
cc_1207 ( N_VDD_c_1229_p N_noxref_10_c_3477_n ) capacitor c=4.31906e-19 \
 //x=24.225 //y=7.4 //x2=23.785 //y2=5.155
cc_1208 ( N_VDD_M72_noxref_d N_noxref_10_c_3477_n ) capacitor c=0.0112985f \
 //x=23.285 //y=5.02 //x2=23.785 //y2=5.155
cc_1209 ( N_VDD_c_944_n N_noxref_10_c_3481_n ) capacitor c=0.00863585f \
 //x=21.46 //y=7.4 //x2=23.075 //y2=5.155
cc_1210 ( N_VDD_M71_noxref_s N_noxref_10_c_3481_n ) capacitor c=0.0831083f \
 //x=22.415 //y=5.02 //x2=23.075 //y2=5.155
cc_1211 ( N_VDD_c_960_p N_noxref_10_c_3483_n ) capacitor c=0.0044221f \
 //x=73.63 //y=7.4 //x2=24.665 //y2=5.155
cc_1212 ( N_VDD_c_1229_p N_noxref_10_c_3483_n ) capacitor c=4.31931e-19 \
 //x=24.225 //y=7.4 //x2=24.665 //y2=5.155
cc_1213 ( N_VDD_c_1176_p N_noxref_10_c_3483_n ) capacitor c=4.31931e-19 \
 //x=25.105 //y=7.4 //x2=24.665 //y2=5.155
cc_1214 ( N_VDD_M74_noxref_d N_noxref_10_c_3483_n ) capacitor c=0.0112985f \
 //x=24.165 //y=5.02 //x2=24.665 //y2=5.155
cc_1215 ( N_VDD_c_960_p N_noxref_10_c_3487_n ) capacitor c=0.00434174f \
 //x=73.63 //y=7.4 //x2=25.445 //y2=5.155
cc_1216 ( N_VDD_c_1176_p N_noxref_10_c_3487_n ) capacitor c=7.46626e-19 \
 //x=25.105 //y=7.4 //x2=25.445 //y2=5.155
cc_1217 ( N_VDD_c_1239_p N_noxref_10_c_3487_n ) capacitor c=0.00198565f \
 //x=26.1 //y=7.4 //x2=25.445 //y2=5.155
cc_1218 ( N_VDD_M76_noxref_d N_noxref_10_c_3487_n ) capacitor c=0.0112985f \
 //x=25.045 //y=5.02 //x2=25.445 //y2=5.155
cc_1219 ( N_VDD_c_945_n N_noxref_10_c_3491_n ) capacitor c=0.0426341f \
 //x=26.27 //y=7.4 //x2=25.53 //y2=3.7
cc_1220 ( N_VDD_c_960_p N_noxref_10_c_3454_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=27.38 //y2=2.08
cc_1221 ( N_VDD_c_1162_p N_noxref_10_c_3454_n ) capacitor c=2.87256e-19 \
 //x=27.855 //y=7.4 //x2=27.38 //y2=2.08
cc_1222 ( N_VDD_c_945_n N_noxref_10_c_3454_n ) capacitor c=0.0134665f \
 //x=26.27 //y=7.4 //x2=27.38 //y2=2.08
cc_1223 ( N_VDD_c_960_p N_noxref_10_c_3455_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=37.37 //y2=2.08
cc_1224 ( N_VDD_c_1246_p N_noxref_10_c_3455_n ) capacitor c=2.87256e-19 \
 //x=37.845 //y=7.4 //x2=37.37 //y2=2.08
cc_1225 ( N_VDD_c_948_n N_noxref_10_c_3455_n ) capacitor c=0.0133642f \
 //x=36.26 //y=7.4 //x2=37.37 //y2=2.08
cc_1226 ( N_VDD_c_1162_p N_noxref_10_M77_noxref_g ) capacitor c=0.00726866f \
 //x=27.855 //y=7.4 //x2=27.28 //y2=6.02
cc_1227 ( N_VDD_M77_noxref_s N_noxref_10_M77_noxref_g ) capacitor c=0.054195f \
 //x=26.925 //y=5.02 //x2=27.28 //y2=6.02
cc_1228 ( N_VDD_c_1162_p N_noxref_10_M78_noxref_g ) capacitor c=0.00672952f \
 //x=27.855 //y=7.4 //x2=27.72 //y2=6.02
cc_1229 ( N_VDD_M78_noxref_d N_noxref_10_M78_noxref_g ) capacitor c=0.015318f \
 //x=27.795 //y=5.02 //x2=27.72 //y2=6.02
cc_1230 ( N_VDD_c_1246_p N_noxref_10_M89_noxref_g ) capacitor c=0.00726866f \
 //x=37.845 //y=7.4 //x2=37.27 //y2=6.02
cc_1231 ( N_VDD_M89_noxref_s N_noxref_10_M89_noxref_g ) capacitor c=0.054195f \
 //x=36.915 //y=5.02 //x2=37.27 //y2=6.02
cc_1232 ( N_VDD_c_1246_p N_noxref_10_M90_noxref_g ) capacitor c=0.00672952f \
 //x=37.845 //y=7.4 //x2=37.71 //y2=6.02
cc_1233 ( N_VDD_M90_noxref_d N_noxref_10_M90_noxref_g ) capacitor c=0.015318f \
 //x=37.785 //y=5.02 //x2=37.71 //y2=6.02
cc_1234 ( N_VDD_c_945_n N_noxref_10_c_3506_n ) capacitor c=0.015293f //x=26.27 \
 //y=7.4 //x2=27.38 //y2=4.7
cc_1235 ( N_VDD_c_948_n N_noxref_10_c_3507_n ) capacitor c=0.0149273f \
 //x=36.26 //y=7.4 //x2=37.37 //y2=4.7
cc_1236 ( N_VDD_c_960_p N_noxref_10_M71_noxref_d ) capacitor c=0.00275235f \
 //x=73.63 //y=7.4 //x2=22.845 //y2=5.02
cc_1237 ( N_VDD_c_1228_p N_noxref_10_M71_noxref_d ) capacitor c=0.014035f \
 //x=23.345 //y=7.4 //x2=22.845 //y2=5.02
cc_1238 ( N_VDD_M72_noxref_d N_noxref_10_M71_noxref_d ) capacitor c=0.0664752f \
 //x=23.285 //y=5.02 //x2=22.845 //y2=5.02
cc_1239 ( N_VDD_c_960_p N_noxref_10_M73_noxref_d ) capacitor c=0.00275186f \
 //x=73.63 //y=7.4 //x2=23.725 //y2=5.02
cc_1240 ( N_VDD_c_1229_p N_noxref_10_M73_noxref_d ) capacitor c=0.0140346f \
 //x=24.225 //y=7.4 //x2=23.725 //y2=5.02
cc_1241 ( N_VDD_c_945_n N_noxref_10_M73_noxref_d ) capacitor c=4.9285e-19 \
 //x=26.27 //y=7.4 //x2=23.725 //y2=5.02
cc_1242 ( N_VDD_M71_noxref_s N_noxref_10_M73_noxref_d ) capacitor \
 c=0.00130656f //x=22.415 //y=5.02 //x2=23.725 //y2=5.02
cc_1243 ( N_VDD_M72_noxref_d N_noxref_10_M73_noxref_d ) capacitor c=0.0664752f \
 //x=23.285 //y=5.02 //x2=23.725 //y2=5.02
cc_1244 ( N_VDD_M74_noxref_d N_noxref_10_M73_noxref_d ) capacitor c=0.0664752f \
 //x=24.165 //y=5.02 //x2=23.725 //y2=5.02
cc_1245 ( N_VDD_c_960_p N_noxref_10_M75_noxref_d ) capacitor c=0.00275235f \
 //x=73.63 //y=7.4 //x2=24.605 //y2=5.02
cc_1246 ( N_VDD_c_1176_p N_noxref_10_M75_noxref_d ) capacitor c=0.0137384f \
 //x=25.105 //y=7.4 //x2=24.605 //y2=5.02
cc_1247 ( N_VDD_c_945_n N_noxref_10_M75_noxref_d ) capacitor c=0.00939849f \
 //x=26.27 //y=7.4 //x2=24.605 //y2=5.02
cc_1248 ( N_VDD_M74_noxref_d N_noxref_10_M75_noxref_d ) capacitor c=0.0664752f \
 //x=24.165 //y=5.02 //x2=24.605 //y2=5.02
cc_1249 ( N_VDD_M76_noxref_d N_noxref_10_M75_noxref_d ) capacitor c=0.0664752f \
 //x=25.045 //y=5.02 //x2=24.605 //y2=5.02
cc_1250 ( N_VDD_M77_noxref_s N_noxref_10_M75_noxref_d ) capacitor \
 c=4.52683e-19 //x=26.925 //y=5.02 //x2=24.605 //y2=5.02
cc_1251 ( N_VDD_c_960_p N_noxref_11_c_3727_n ) capacitor c=0.00453663f \
 //x=73.63 //y=7.4 //x2=38.285 //y2=5.2
cc_1252 ( N_VDD_c_1246_p N_noxref_11_c_3727_n ) capacitor c=4.48391e-19 \
 //x=37.845 //y=7.4 //x2=38.285 //y2=5.2
cc_1253 ( N_VDD_c_1275_p N_noxref_11_c_3727_n ) capacitor c=4.48391e-19 \
 //x=38.725 //y=7.4 //x2=38.285 //y2=5.2
cc_1254 ( N_VDD_M90_noxref_d N_noxref_11_c_3727_n ) capacitor c=0.0124542f \
 //x=37.785 //y=5.02 //x2=38.285 //y2=5.2
cc_1255 ( N_VDD_c_948_n N_noxref_11_c_3731_n ) capacitor c=0.00985474f \
 //x=36.26 //y=7.4 //x2=37.575 //y2=5.2
cc_1256 ( N_VDD_M89_noxref_s N_noxref_11_c_3731_n ) capacitor c=0.087833f \
 //x=36.915 //y=5.02 //x2=37.575 //y2=5.2
cc_1257 ( N_VDD_c_960_p N_noxref_11_c_3733_n ) capacitor c=0.00301575f \
 //x=73.63 //y=7.4 //x2=38.765 //y2=5.2
cc_1258 ( N_VDD_c_1275_p N_noxref_11_c_3733_n ) capacitor c=7.72068e-19 \
 //x=38.725 //y=7.4 //x2=38.765 //y2=5.2
cc_1259 ( N_VDD_M92_noxref_d N_noxref_11_c_3733_n ) capacitor c=0.0158515f \
 //x=38.665 //y=5.02 //x2=38.765 //y2=5.2
cc_1260 ( N_VDD_M93_noxref_s N_noxref_11_c_3733_n ) capacitor c=2.44532e-19 \
 //x=40.245 //y=5.02 //x2=38.765 //y2=5.2
cc_1261 ( N_VDD_c_948_n N_noxref_11_c_3712_n ) capacitor c=0.00151618f \
 //x=36.26 //y=7.4 //x2=38.85 //y2=3.7
cc_1262 ( N_VDD_c_949_n N_noxref_11_c_3712_n ) capacitor c=0.0429414f \
 //x=39.59 //y=7.4 //x2=38.85 //y2=3.7
cc_1263 ( N_VDD_c_960_p N_noxref_11_c_3713_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=40.7 //y2=2.08
cc_1264 ( N_VDD_c_1286_p N_noxref_11_c_3713_n ) capacitor c=2.87256e-19 \
 //x=41.175 //y=7.4 //x2=40.7 //y2=2.08
cc_1265 ( N_VDD_c_949_n N_noxref_11_c_3713_n ) capacitor c=0.0134208f \
 //x=39.59 //y=7.4 //x2=40.7 //y2=2.08
cc_1266 ( N_VDD_c_1286_p N_noxref_11_M93_noxref_g ) capacitor c=0.00726866f \
 //x=41.175 //y=7.4 //x2=40.6 //y2=6.02
cc_1267 ( N_VDD_M93_noxref_s N_noxref_11_M93_noxref_g ) capacitor c=0.054195f \
 //x=40.245 //y=5.02 //x2=40.6 //y2=6.02
cc_1268 ( N_VDD_c_1286_p N_noxref_11_M94_noxref_g ) capacitor c=0.00672952f \
 //x=41.175 //y=7.4 //x2=41.04 //y2=6.02
cc_1269 ( N_VDD_M94_noxref_d N_noxref_11_M94_noxref_g ) capacitor c=0.015318f \
 //x=41.115 //y=5.02 //x2=41.04 //y2=6.02
cc_1270 ( N_VDD_c_949_n N_noxref_11_c_3746_n ) capacitor c=0.0150435f \
 //x=39.59 //y=7.4 //x2=40.7 //y2=4.7
cc_1271 ( N_VDD_c_960_p N_noxref_11_M89_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=37.345 //y2=5.02
cc_1272 ( N_VDD_c_1246_p N_noxref_11_M89_noxref_d ) capacitor c=0.0140317f \
 //x=37.845 //y=7.4 //x2=37.345 //y2=5.02
cc_1273 ( N_VDD_c_949_n N_noxref_11_M89_noxref_d ) capacitor c=6.94454e-19 \
 //x=39.59 //y=7.4 //x2=37.345 //y2=5.02
cc_1274 ( N_VDD_M90_noxref_d N_noxref_11_M89_noxref_d ) capacitor c=0.0664752f \
 //x=37.785 //y=5.02 //x2=37.345 //y2=5.02
cc_1275 ( N_VDD_c_960_p N_noxref_11_M91_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=38.225 //y2=5.02
cc_1276 ( N_VDD_c_1275_p N_noxref_11_M91_noxref_d ) capacitor c=0.0140317f \
 //x=38.725 //y=7.4 //x2=38.225 //y2=5.02
cc_1277 ( N_VDD_c_949_n N_noxref_11_M91_noxref_d ) capacitor c=0.0120541f \
 //x=39.59 //y=7.4 //x2=38.225 //y2=5.02
cc_1278 ( N_VDD_M89_noxref_s N_noxref_11_M91_noxref_d ) capacitor \
 c=0.00111971f //x=36.915 //y=5.02 //x2=38.225 //y2=5.02
cc_1279 ( N_VDD_M90_noxref_d N_noxref_11_M91_noxref_d ) capacitor c=0.0664752f \
 //x=37.785 //y=5.02 //x2=38.225 //y2=5.02
cc_1280 ( N_VDD_M92_noxref_d N_noxref_11_M91_noxref_d ) capacitor c=0.0664752f \
 //x=38.665 //y=5.02 //x2=38.225 //y2=5.02
cc_1281 ( N_VDD_M93_noxref_s N_noxref_11_M91_noxref_d ) capacitor \
 c=4.54516e-19 //x=40.245 //y=5.02 //x2=38.225 //y2=5.02
cc_1282 ( N_VDD_c_945_n N_noxref_12_c_3882_n ) capacitor c=0.0140578f \
 //x=26.27 //y=7.4 //x2=31.335 //y2=4.07
cc_1283 ( N_VDD_c_946_n N_noxref_12_c_3882_n ) capacitor c=0.0140578f //x=29.6 \
 //y=7.4 //x2=31.335 //y2=4.07
cc_1284 ( N_VDD_c_944_n N_noxref_12_c_3884_n ) capacitor c=0.00116746f \
 //x=21.46 //y=7.4 //x2=22.685 //y2=4.07
cc_1285 ( N_VDD_c_947_n N_noxref_12_c_3885_n ) capacitor c=0.0140578f \
 //x=32.93 //y=7.4 //x2=35.405 //y2=4.07
cc_1286 ( N_VDD_c_948_n N_noxref_12_c_3886_n ) capacitor c=0.0140578f \
 //x=36.26 //y=7.4 //x2=41.325 //y2=4.07
cc_1287 ( N_VDD_c_949_n N_noxref_12_c_3886_n ) capacitor c=0.0140578f \
 //x=39.59 //y=7.4 //x2=41.325 //y2=4.07
cc_1288 ( N_VDD_c_948_n N_noxref_12_c_3888_n ) capacitor c=0.00104972f \
 //x=36.26 //y=7.4 //x2=35.635 //y2=4.07
cc_1289 ( N_VDD_c_960_p N_noxref_12_c_3862_n ) capacitor c=9.10347e-19 \
 //x=73.63 //y=7.4 //x2=22.57 //y2=2.08
cc_1290 ( N_VDD_c_944_n N_noxref_12_c_3862_n ) capacitor c=0.0137129f \
 //x=21.46 //y=7.4 //x2=22.57 //y2=2.08
cc_1291 ( N_VDD_M71_noxref_s N_noxref_12_c_3862_n ) capacitor c=0.0120327f \
 //x=22.415 //y=5.02 //x2=22.57 //y2=2.08
cc_1292 ( N_VDD_c_946_n N_noxref_12_c_3863_n ) capacitor c=4.57806e-19 \
 //x=29.6 //y=7.4 //x2=31.45 //y2=2.08
cc_1293 ( N_VDD_c_947_n N_noxref_12_c_3863_n ) capacitor c=3.69525e-19 \
 //x=32.93 //y=7.4 //x2=31.45 //y2=2.08
cc_1294 ( N_VDD_c_960_p N_noxref_12_c_3894_n ) capacitor c=0.00453473f \
 //x=73.63 //y=7.4 //x2=34.955 //y2=5.2
cc_1295 ( N_VDD_c_1209_p N_noxref_12_c_3894_n ) capacitor c=4.48391e-19 \
 //x=34.515 //y=7.4 //x2=34.955 //y2=5.2
cc_1296 ( N_VDD_c_1318_p N_noxref_12_c_3894_n ) capacitor c=4.48377e-19 \
 //x=35.395 //y=7.4 //x2=34.955 //y2=5.2
cc_1297 ( N_VDD_M86_noxref_d N_noxref_12_c_3894_n ) capacitor c=0.0124506f \
 //x=34.455 //y=5.02 //x2=34.955 //y2=5.2
cc_1298 ( N_VDD_c_947_n N_noxref_12_c_3898_n ) capacitor c=0.00985474f \
 //x=32.93 //y=7.4 //x2=34.245 //y2=5.2
cc_1299 ( N_VDD_M85_noxref_s N_noxref_12_c_3898_n ) capacitor c=0.087833f \
 //x=33.585 //y=5.02 //x2=34.245 //y2=5.2
cc_1300 ( N_VDD_c_960_p N_noxref_12_c_3900_n ) capacitor c=0.00301575f \
 //x=73.63 //y=7.4 //x2=35.435 //y2=5.2
cc_1301 ( N_VDD_c_1318_p N_noxref_12_c_3900_n ) capacitor c=7.72068e-19 \
 //x=35.395 //y=7.4 //x2=35.435 //y2=5.2
cc_1302 ( N_VDD_M88_noxref_d N_noxref_12_c_3900_n ) capacitor c=0.0158515f \
 //x=35.335 //y=5.02 //x2=35.435 //y2=5.2
cc_1303 ( N_VDD_M89_noxref_s N_noxref_12_c_3900_n ) capacitor c=2.44532e-19 \
 //x=36.915 //y=5.02 //x2=35.435 //y2=5.2
cc_1304 ( N_VDD_c_947_n N_noxref_12_c_3866_n ) capacitor c=0.00151618f \
 //x=32.93 //y=7.4 //x2=35.52 //y2=4.07
cc_1305 ( N_VDD_c_948_n N_noxref_12_c_3866_n ) capacitor c=0.043035f //x=36.26 \
 //y=7.4 //x2=35.52 //y2=4.07
cc_1306 ( N_VDD_c_949_n N_noxref_12_c_3867_n ) capacitor c=4.57806e-19 \
 //x=39.59 //y=7.4 //x2=41.44 //y2=2.08
cc_1307 ( N_VDD_c_950_n N_noxref_12_c_3867_n ) capacitor c=4.17938e-19 \
 //x=42.92 //y=7.4 //x2=41.44 //y2=2.08
cc_1308 ( N_VDD_c_1228_p N_noxref_12_M71_noxref_g ) capacitor c=0.00749687f \
 //x=23.345 //y=7.4 //x2=22.77 //y2=6.02
cc_1309 ( N_VDD_M71_noxref_s N_noxref_12_M71_noxref_g ) capacitor c=0.0477201f \
 //x=22.415 //y=5.02 //x2=22.77 //y2=6.02
cc_1310 ( N_VDD_c_1228_p N_noxref_12_M72_noxref_g ) capacitor c=0.00675175f \
 //x=23.345 //y=7.4 //x2=23.21 //y2=6.02
cc_1311 ( N_VDD_M72_noxref_d N_noxref_12_M72_noxref_g ) capacitor c=0.015318f \
 //x=23.285 //y=5.02 //x2=23.21 //y2=6.02
cc_1312 ( N_VDD_c_1198_p N_noxref_12_M83_noxref_g ) capacitor c=0.00673971f \
 //x=32.065 //y=7.4 //x2=31.49 //y2=6.02
cc_1313 ( N_VDD_M82_noxref_d N_noxref_12_M83_noxref_g ) capacitor c=0.015318f \
 //x=31.125 //y=5.02 //x2=31.49 //y2=6.02
cc_1314 ( N_VDD_c_1198_p N_noxref_12_M84_noxref_g ) capacitor c=0.00672952f \
 //x=32.065 //y=7.4 //x2=31.93 //y2=6.02
cc_1315 ( N_VDD_c_947_n N_noxref_12_M84_noxref_g ) capacitor c=0.00864163f \
 //x=32.93 //y=7.4 //x2=31.93 //y2=6.02
cc_1316 ( N_VDD_M84_noxref_d N_noxref_12_M84_noxref_g ) capacitor c=0.0430452f \
 //x=32.005 //y=5.02 //x2=31.93 //y2=6.02
cc_1317 ( N_VDD_c_1339_p N_noxref_12_M95_noxref_g ) capacitor c=0.00673971f \
 //x=42.055 //y=7.4 //x2=41.48 //y2=6.02
cc_1318 ( N_VDD_M94_noxref_d N_noxref_12_M95_noxref_g ) capacitor c=0.015318f \
 //x=41.115 //y=5.02 //x2=41.48 //y2=6.02
cc_1319 ( N_VDD_c_1339_p N_noxref_12_M96_noxref_g ) capacitor c=0.00672952f \
 //x=42.055 //y=7.4 //x2=41.92 //y2=6.02
cc_1320 ( N_VDD_c_950_n N_noxref_12_M96_noxref_g ) capacitor c=0.00928743f \
 //x=42.92 //y=7.4 //x2=41.92 //y2=6.02
cc_1321 ( N_VDD_M96_noxref_d N_noxref_12_M96_noxref_g ) capacitor c=0.0430452f \
 //x=41.995 //y=5.02 //x2=41.92 //y2=6.02
cc_1322 ( N_VDD_c_944_n N_noxref_12_c_3922_n ) capacitor c=0.00757682f \
 //x=21.46 //y=7.4 //x2=22.845 //y2=4.79
cc_1323 ( N_VDD_M71_noxref_s N_noxref_12_c_3922_n ) capacitor c=0.00444914f \
 //x=22.415 //y=5.02 //x2=22.845 //y2=4.79
cc_1324 ( N_VDD_c_960_p N_noxref_12_M85_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=34.015 //y2=5.02
cc_1325 ( N_VDD_c_1209_p N_noxref_12_M85_noxref_d ) capacitor c=0.0140317f \
 //x=34.515 //y=7.4 //x2=34.015 //y2=5.02
cc_1326 ( N_VDD_c_948_n N_noxref_12_M85_noxref_d ) capacitor c=6.94454e-19 \
 //x=36.26 //y=7.4 //x2=34.015 //y2=5.02
cc_1327 ( N_VDD_M86_noxref_d N_noxref_12_M85_noxref_d ) capacitor c=0.0664752f \
 //x=34.455 //y=5.02 //x2=34.015 //y2=5.02
cc_1328 ( N_VDD_c_960_p N_noxref_12_M87_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=34.895 //y2=5.02
cc_1329 ( N_VDD_c_1318_p N_noxref_12_M87_noxref_d ) capacitor c=0.0140317f \
 //x=35.395 //y=7.4 //x2=34.895 //y2=5.02
cc_1330 ( N_VDD_c_948_n N_noxref_12_M87_noxref_d ) capacitor c=0.0120541f \
 //x=36.26 //y=7.4 //x2=34.895 //y2=5.02
cc_1331 ( N_VDD_M85_noxref_s N_noxref_12_M87_noxref_d ) capacitor \
 c=0.00111971f //x=33.585 //y=5.02 //x2=34.895 //y2=5.02
cc_1332 ( N_VDD_M86_noxref_d N_noxref_12_M87_noxref_d ) capacitor c=0.0664752f \
 //x=34.455 //y=5.02 //x2=34.895 //y2=5.02
cc_1333 ( N_VDD_M88_noxref_d N_noxref_12_M87_noxref_d ) capacitor c=0.0664752f \
 //x=35.335 //y=5.02 //x2=34.895 //y2=5.02
cc_1334 ( N_VDD_M89_noxref_s N_noxref_12_M87_noxref_d ) capacitor \
 c=4.54516e-19 //x=36.915 //y=5.02 //x2=34.895 //y2=5.02
cc_1335 ( N_VDD_c_939_n N_D_c_4253_n ) capacitor c=4.47073e-19 //x=4.81 \
 //y=7.4 //x2=6.66 //y2=2.08
cc_1336 ( N_VDD_c_940_n N_D_c_4253_n ) capacitor c=3.37458e-19 //x=8.14 \
 //y=7.4 //x2=6.66 //y2=2.08
cc_1337 ( N_VDD_c_945_n N_D_c_4255_n ) capacitor c=4.47073e-19 //x=26.27 \
 //y=7.4 //x2=28.12 //y2=2.08
cc_1338 ( N_VDD_c_946_n N_D_c_4255_n ) capacitor c=3.37458e-19 //x=29.6 \
 //y=7.4 //x2=28.12 //y2=2.08
cc_1339 ( N_VDD_c_951_n N_D_c_4257_n ) capacitor c=4.47073e-19 //x=47.73 \
 //y=7.4 //x2=49.58 //y2=2.08
cc_1340 ( N_VDD_c_952_n N_D_c_4257_n ) capacitor c=3.37458e-19 //x=51.06 \
 //y=7.4 //x2=49.58 //y2=2.08
cc_1341 ( N_VDD_c_962_p N_D_M53_noxref_g ) capacitor c=0.00673971f //x=7.275 \
 //y=7.4 //x2=6.7 //y2=6.02
cc_1342 ( N_VDD_M52_noxref_d N_D_M53_noxref_g ) capacitor c=0.015318f \
 //x=6.335 //y=5.02 //x2=6.7 //y2=6.02
cc_1343 ( N_VDD_c_962_p N_D_M54_noxref_g ) capacitor c=0.00672952f //x=7.275 \
 //y=7.4 //x2=7.14 //y2=6.02
cc_1344 ( N_VDD_c_940_n N_D_M54_noxref_g ) capacitor c=0.00864163f //x=8.14 \
 //y=7.4 //x2=7.14 //y2=6.02
cc_1345 ( N_VDD_M54_noxref_d N_D_M54_noxref_g ) capacitor c=0.0430452f \
 //x=7.215 //y=5.02 //x2=7.14 //y2=6.02
cc_1346 ( N_VDD_c_1163_p N_D_M79_noxref_g ) capacitor c=0.00673971f //x=28.735 \
 //y=7.4 //x2=28.16 //y2=6.02
cc_1347 ( N_VDD_M78_noxref_d N_D_M79_noxref_g ) capacitor c=0.015318f \
 //x=27.795 //y=5.02 //x2=28.16 //y2=6.02
cc_1348 ( N_VDD_c_1163_p N_D_M80_noxref_g ) capacitor c=0.00672952f //x=28.735 \
 //y=7.4 //x2=28.6 //y2=6.02
cc_1349 ( N_VDD_c_946_n N_D_M80_noxref_g ) capacitor c=0.00864163f //x=29.6 \
 //y=7.4 //x2=28.6 //y2=6.02
cc_1350 ( N_VDD_M80_noxref_d N_D_M80_noxref_g ) capacitor c=0.0430452f \
 //x=28.675 //y=5.02 //x2=28.6 //y2=6.02
cc_1351 ( N_VDD_c_1373_p N_D_M105_noxref_g ) capacitor c=0.00673971f \
 //x=50.195 //y=7.4 //x2=49.62 //y2=6.02
cc_1352 ( N_VDD_M104_noxref_d N_D_M105_noxref_g ) capacitor c=0.015318f \
 //x=49.255 //y=5.02 //x2=49.62 //y2=6.02
cc_1353 ( N_VDD_c_1373_p N_D_M106_noxref_g ) capacitor c=0.00672952f \
 //x=50.195 //y=7.4 //x2=50.06 //y2=6.02
cc_1354 ( N_VDD_c_952_n N_D_M106_noxref_g ) capacitor c=0.00864163f //x=51.06 \
 //y=7.4 //x2=50.06 //y2=6.02
cc_1355 ( N_VDD_M106_noxref_d N_D_M106_noxref_g ) capacitor c=0.0430452f \
 //x=50.135 //y=5.02 //x2=50.06 //y2=6.02
cc_1356 ( N_VDD_c_951_n N_noxref_14_c_4641_n ) capacitor c=6.58823e-19 \
 //x=47.73 //y=7.4 //x2=46.25 //y2=2.08
cc_1357 ( N_VDD_c_960_p N_noxref_14_c_4659_n ) capacitor c=0.00453663f \
 //x=73.63 //y=7.4 //x2=49.755 //y2=5.2
cc_1358 ( N_VDD_c_1380_p N_noxref_14_c_4659_n ) capacitor c=4.48391e-19 \
 //x=49.315 //y=7.4 //x2=49.755 //y2=5.2
cc_1359 ( N_VDD_c_1373_p N_noxref_14_c_4659_n ) capacitor c=4.48391e-19 \
 //x=50.195 //y=7.4 //x2=49.755 //y2=5.2
cc_1360 ( N_VDD_M104_noxref_d N_noxref_14_c_4659_n ) capacitor c=0.0124542f \
 //x=49.255 //y=5.02 //x2=49.755 //y2=5.2
cc_1361 ( N_VDD_c_951_n N_noxref_14_c_4663_n ) capacitor c=0.00985474f \
 //x=47.73 //y=7.4 //x2=49.045 //y2=5.2
cc_1362 ( N_VDD_M103_noxref_s N_noxref_14_c_4663_n ) capacitor c=0.087833f \
 //x=48.385 //y=5.02 //x2=49.045 //y2=5.2
cc_1363 ( N_VDD_c_960_p N_noxref_14_c_4665_n ) capacitor c=0.00301575f \
 //x=73.63 //y=7.4 //x2=50.235 //y2=5.2
cc_1364 ( N_VDD_c_1373_p N_noxref_14_c_4665_n ) capacitor c=7.72068e-19 \
 //x=50.195 //y=7.4 //x2=50.235 //y2=5.2
cc_1365 ( N_VDD_M106_noxref_d N_noxref_14_c_4665_n ) capacitor c=0.0158515f \
 //x=50.135 //y=5.02 //x2=50.235 //y2=5.2
cc_1366 ( N_VDD_M107_noxref_s N_noxref_14_c_4665_n ) capacitor c=2.44532e-19 \
 //x=51.715 //y=5.02 //x2=50.235 //y2=5.2
cc_1367 ( N_VDD_c_951_n N_noxref_14_c_4643_n ) capacitor c=0.00151618f \
 //x=47.73 //y=7.4 //x2=50.32 //y2=3.33
cc_1368 ( N_VDD_c_952_n N_noxref_14_c_4643_n ) capacitor c=0.0429414f \
 //x=51.06 //y=7.4 //x2=50.32 //y2=3.33
cc_1369 ( N_VDD_c_960_p N_noxref_14_c_4644_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=52.17 //y2=2.08
cc_1370 ( N_VDD_c_1392_p N_noxref_14_c_4644_n ) capacitor c=2.87256e-19 \
 //x=52.645 //y=7.4 //x2=52.17 //y2=2.08
cc_1371 ( N_VDD_c_952_n N_noxref_14_c_4644_n ) capacitor c=0.0134208f \
 //x=51.06 //y=7.4 //x2=52.17 //y2=2.08
cc_1372 ( N_VDD_c_1394_p N_noxref_14_M101_noxref_g ) capacitor c=0.00675175f \
 //x=46.565 //y=7.4 //x2=45.99 //y2=6.02
cc_1373 ( N_VDD_M100_noxref_d N_noxref_14_M101_noxref_g ) capacitor \
 c=0.015318f //x=45.625 //y=5.02 //x2=45.99 //y2=6.02
cc_1374 ( N_VDD_c_1394_p N_noxref_14_M102_noxref_g ) capacitor c=0.00675379f \
 //x=46.565 //y=7.4 //x2=46.43 //y2=6.02
cc_1375 ( N_VDD_M102_noxref_d N_noxref_14_M102_noxref_g ) capacitor \
 c=0.0394719f //x=46.505 //y=5.02 //x2=46.43 //y2=6.02
cc_1376 ( N_VDD_c_1392_p N_noxref_14_M107_noxref_g ) capacitor c=0.00726866f \
 //x=52.645 //y=7.4 //x2=52.07 //y2=6.02
cc_1377 ( N_VDD_M107_noxref_s N_noxref_14_M107_noxref_g ) capacitor \
 c=0.054195f //x=51.715 //y=5.02 //x2=52.07 //y2=6.02
cc_1378 ( N_VDD_c_1392_p N_noxref_14_M108_noxref_g ) capacitor c=0.00672952f \
 //x=52.645 //y=7.4 //x2=52.51 //y2=6.02
cc_1379 ( N_VDD_M108_noxref_d N_noxref_14_M108_noxref_g ) capacitor \
 c=0.015318f //x=52.585 //y=5.02 //x2=52.51 //y2=6.02
cc_1380 ( N_VDD_c_952_n N_noxref_14_c_4682_n ) capacitor c=0.0150435f \
 //x=51.06 //y=7.4 //x2=52.17 //y2=4.7
cc_1381 ( N_VDD_c_960_p N_noxref_14_M103_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=48.815 //y2=5.02
cc_1382 ( N_VDD_c_1380_p N_noxref_14_M103_noxref_d ) capacitor c=0.0140317f \
 //x=49.315 //y=7.4 //x2=48.815 //y2=5.02
cc_1383 ( N_VDD_c_952_n N_noxref_14_M103_noxref_d ) capacitor c=6.94454e-19 \
 //x=51.06 //y=7.4 //x2=48.815 //y2=5.02
cc_1384 ( N_VDD_M104_noxref_d N_noxref_14_M103_noxref_d ) capacitor \
 c=0.0664752f //x=49.255 //y=5.02 //x2=48.815 //y2=5.02
cc_1385 ( N_VDD_c_960_p N_noxref_14_M105_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=49.695 //y2=5.02
cc_1386 ( N_VDD_c_1373_p N_noxref_14_M105_noxref_d ) capacitor c=0.0140317f \
 //x=50.195 //y=7.4 //x2=49.695 //y2=5.02
cc_1387 ( N_VDD_c_952_n N_noxref_14_M105_noxref_d ) capacitor c=0.0120541f \
 //x=51.06 //y=7.4 //x2=49.695 //y2=5.02
cc_1388 ( N_VDD_M103_noxref_s N_noxref_14_M105_noxref_d ) capacitor \
 c=0.00111971f //x=48.385 //y=5.02 //x2=49.695 //y2=5.02
cc_1389 ( N_VDD_M104_noxref_d N_noxref_14_M105_noxref_d ) capacitor \
 c=0.0664752f //x=49.255 //y=5.02 //x2=49.695 //y2=5.02
cc_1390 ( N_VDD_M106_noxref_d N_noxref_14_M105_noxref_d ) capacitor \
 c=0.0664752f //x=50.135 //y=5.02 //x2=49.695 //y2=5.02
cc_1391 ( N_VDD_M107_noxref_s N_noxref_14_M105_noxref_d ) capacitor \
 c=4.54516e-19 //x=51.715 //y=5.02 //x2=49.695 //y2=5.02
cc_1392 ( N_VDD_c_960_p N_noxref_15_c_4890_n ) capacitor c=0.00453663f \
 //x=73.63 //y=7.4 //x2=53.085 //y2=5.2
cc_1393 ( N_VDD_c_1392_p N_noxref_15_c_4890_n ) capacitor c=4.48391e-19 \
 //x=52.645 //y=7.4 //x2=53.085 //y2=5.2
cc_1394 ( N_VDD_c_1416_p N_noxref_15_c_4890_n ) capacitor c=4.48391e-19 \
 //x=53.525 //y=7.4 //x2=53.085 //y2=5.2
cc_1395 ( N_VDD_M108_noxref_d N_noxref_15_c_4890_n ) capacitor c=0.0124542f \
 //x=52.585 //y=5.02 //x2=53.085 //y2=5.2
cc_1396 ( N_VDD_c_952_n N_noxref_15_c_4894_n ) capacitor c=0.00985474f \
 //x=51.06 //y=7.4 //x2=52.375 //y2=5.2
cc_1397 ( N_VDD_M107_noxref_s N_noxref_15_c_4894_n ) capacitor c=0.087833f \
 //x=51.715 //y=5.02 //x2=52.375 //y2=5.2
cc_1398 ( N_VDD_c_960_p N_noxref_15_c_4896_n ) capacitor c=0.00301575f \
 //x=73.63 //y=7.4 //x2=53.565 //y2=5.2
cc_1399 ( N_VDD_c_1416_p N_noxref_15_c_4896_n ) capacitor c=7.72068e-19 \
 //x=53.525 //y=7.4 //x2=53.565 //y2=5.2
cc_1400 ( N_VDD_M110_noxref_d N_noxref_15_c_4896_n ) capacitor c=0.0158515f \
 //x=53.465 //y=5.02 //x2=53.565 //y2=5.2
cc_1401 ( N_VDD_M111_noxref_s N_noxref_15_c_4896_n ) capacitor c=2.44532e-19 \
 //x=55.045 //y=5.02 //x2=53.565 //y2=5.2
cc_1402 ( N_VDD_c_952_n N_noxref_15_c_4875_n ) capacitor c=0.00151618f \
 //x=51.06 //y=7.4 //x2=53.65 //y2=3.33
cc_1403 ( N_VDD_c_953_n N_noxref_15_c_4875_n ) capacitor c=0.0427674f \
 //x=54.39 //y=7.4 //x2=53.65 //y2=3.33
cc_1404 ( N_VDD_c_960_p N_noxref_15_c_4876_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=55.5 //y2=2.08
cc_1405 ( N_VDD_c_1427_p N_noxref_15_c_4876_n ) capacitor c=2.87256e-19 \
 //x=55.975 //y=7.4 //x2=55.5 //y2=2.08
cc_1406 ( N_VDD_c_953_n N_noxref_15_c_4876_n ) capacitor c=0.0133228f \
 //x=54.39 //y=7.4 //x2=55.5 //y2=2.08
cc_1407 ( N_VDD_c_1427_p N_noxref_15_M111_noxref_g ) capacitor c=0.00726866f \
 //x=55.975 //y=7.4 //x2=55.4 //y2=6.02
cc_1408 ( N_VDD_M111_noxref_s N_noxref_15_M111_noxref_g ) capacitor \
 c=0.054195f //x=55.045 //y=5.02 //x2=55.4 //y2=6.02
cc_1409 ( N_VDD_c_1427_p N_noxref_15_M112_noxref_g ) capacitor c=0.00672952f \
 //x=55.975 //y=7.4 //x2=55.84 //y2=6.02
cc_1410 ( N_VDD_M112_noxref_d N_noxref_15_M112_noxref_g ) capacitor \
 c=0.015318f //x=55.915 //y=5.02 //x2=55.84 //y2=6.02
cc_1411 ( N_VDD_c_953_n N_noxref_15_c_4909_n ) capacitor c=0.0149273f \
 //x=54.39 //y=7.4 //x2=55.5 //y2=4.7
cc_1412 ( N_VDD_c_960_p N_noxref_15_M107_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=52.145 //y2=5.02
cc_1413 ( N_VDD_c_1392_p N_noxref_15_M107_noxref_d ) capacitor c=0.0140317f \
 //x=52.645 //y=7.4 //x2=52.145 //y2=5.02
cc_1414 ( N_VDD_c_953_n N_noxref_15_M107_noxref_d ) capacitor c=6.94454e-19 \
 //x=54.39 //y=7.4 //x2=52.145 //y2=5.02
cc_1415 ( N_VDD_M108_noxref_d N_noxref_15_M107_noxref_d ) capacitor \
 c=0.0664752f //x=52.585 //y=5.02 //x2=52.145 //y2=5.02
cc_1416 ( N_VDD_c_960_p N_noxref_15_M109_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=53.025 //y2=5.02
cc_1417 ( N_VDD_c_1416_p N_noxref_15_M109_noxref_d ) capacitor c=0.0140317f \
 //x=53.525 //y=7.4 //x2=53.025 //y2=5.02
cc_1418 ( N_VDD_c_953_n N_noxref_15_M109_noxref_d ) capacitor c=0.0120541f \
 //x=54.39 //y=7.4 //x2=53.025 //y2=5.02
cc_1419 ( N_VDD_M107_noxref_s N_noxref_15_M109_noxref_d ) capacitor \
 c=0.00111971f //x=51.715 //y=5.02 //x2=53.025 //y2=5.02
cc_1420 ( N_VDD_M108_noxref_d N_noxref_15_M109_noxref_d ) capacitor \
 c=0.0664752f //x=52.585 //y=5.02 //x2=53.025 //y2=5.02
cc_1421 ( N_VDD_M110_noxref_d N_noxref_15_M109_noxref_d ) capacitor \
 c=0.0664752f //x=53.465 //y=5.02 //x2=53.025 //y2=5.02
cc_1422 ( N_VDD_M111_noxref_s N_noxref_15_M109_noxref_d ) capacitor \
 c=4.54516e-19 //x=55.045 //y=5.02 //x2=53.025 //y2=5.02
cc_1423 ( N_VDD_c_960_p N_CLK_c_5034_n ) capacitor c=0.0809378f //x=73.63 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1424 ( N_VDD_c_1038_p N_CLK_c_5034_n ) capacitor c=0.00258496f //x=4.64 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1425 ( N_VDD_c_1447_p N_CLK_c_5034_n ) capacitor c=0.00209689f //x=5.515 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1426 ( N_VDD_c_961_p N_CLK_c_5034_n ) capacitor c=7.81728e-19 //x=6.395 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1427 ( N_VDD_c_1449_p N_CLK_c_5034_n ) capacitor c=0.00205475f //x=7.97 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1428 ( N_VDD_c_1450_p N_CLK_c_5034_n ) capacitor c=0.00209689f //x=8.845 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1429 ( N_VDD_c_973_p N_CLK_c_5034_n ) capacitor c=7.81728e-19 //x=9.725 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1430 ( N_VDD_c_1452_p N_CLK_c_5034_n ) capacitor c=0.00205475f //x=11.3 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1431 ( N_VDD_c_1453_p N_CLK_c_5034_n ) capacitor c=0.00209689f //x=12.175 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1432 ( N_VDD_c_1008_p N_CLK_c_5034_n ) capacitor c=7.81728e-19 //x=13.055 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1433 ( N_VDD_c_939_n N_CLK_c_5034_n ) capacitor c=0.0389825f //x=4.81 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1434 ( N_VDD_c_940_n N_CLK_c_5034_n ) capacitor c=0.0389825f //x=8.14 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1435 ( N_VDD_c_941_n N_CLK_c_5034_n ) capacitor c=0.0389825f //x=11.47 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_1436 ( N_VDD_M51_noxref_s N_CLK_c_5034_n ) capacitor c=0.00541054f \
 //x=5.465 //y=5.02 //x2=13.205 //y2=4.44
cc_1437 ( N_VDD_M54_noxref_d N_CLK_c_5034_n ) capacitor c=6.7165e-19 //x=7.215 \
 //y=5.02 //x2=13.205 //y2=4.44
cc_1438 ( N_VDD_M55_noxref_s N_CLK_c_5034_n ) capacitor c=0.00541054f \
 //x=8.795 //y=5.02 //x2=13.205 //y2=4.44
cc_1439 ( N_VDD_M58_noxref_d N_CLK_c_5034_n ) capacitor c=6.7165e-19 \
 //x=10.545 //y=5.02 //x2=13.205 //y2=4.44
cc_1440 ( N_VDD_M59_noxref_s N_CLK_c_5034_n ) capacitor c=0.00541054f \
 //x=12.125 //y=5.02 //x2=13.205 //y2=4.44
cc_1441 ( N_VDD_c_960_p N_CLK_c_5052_n ) capacitor c=0.00146064f //x=73.63 \
 //y=7.4 //x2=2.335 //y2=4.44
cc_1442 ( N_VDD_c_960_p N_CLK_c_5053_n ) capacitor c=0.023948f //x=73.63 \
 //y=7.4 //x2=16.745 //y2=4.442
cc_1443 ( N_VDD_c_1465_p N_CLK_c_5053_n ) capacitor c=0.0020391f //x=14.63 \
 //y=7.4 //x2=16.745 //y2=4.442
cc_1444 ( N_VDD_c_1466_p N_CLK_c_5053_n ) capacitor c=0.002081f //x=15.505 \
 //y=7.4 //x2=16.745 //y2=4.442
cc_1445 ( N_VDD_c_1045_p N_CLK_c_5053_n ) capacitor c=7.79455e-19 //x=16.385 \
 //y=7.4 //x2=16.745 //y2=4.442
cc_1446 ( N_VDD_c_942_n N_CLK_c_5053_n ) capacitor c=0.037674f //x=14.8 \
 //y=7.4 //x2=16.745 //y2=4.442
cc_1447 ( N_VDD_M62_noxref_d N_CLK_c_5053_n ) capacitor c=6.65538e-19 \
 //x=13.875 //y=5.02 //x2=16.745 //y2=4.442
cc_1448 ( N_VDD_M63_noxref_s N_CLK_c_5053_n ) capacitor c=0.00527639f \
 //x=15.455 //y=5.02 //x2=16.745 //y2=4.442
cc_1449 ( N_VDD_c_960_p N_CLK_c_5060_n ) capacitor c=0.00149167f //x=73.63 \
 //y=7.4 //x2=13.465 //y2=4.442
cc_1450 ( N_VDD_c_960_p N_CLK_c_5061_n ) capacitor c=0.0809378f //x=73.63 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1451 ( N_VDD_c_1239_p N_CLK_c_5061_n ) capacitor c=0.00258496f //x=26.1 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1452 ( N_VDD_c_1474_p N_CLK_c_5061_n ) capacitor c=0.00209689f //x=26.975 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1453 ( N_VDD_c_1162_p N_CLK_c_5061_n ) capacitor c=7.81728e-19 //x=27.855 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1454 ( N_VDD_c_1476_p N_CLK_c_5061_n ) capacitor c=0.00205475f //x=29.43 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1455 ( N_VDD_c_1477_p N_CLK_c_5061_n ) capacitor c=0.00209689f //x=30.305 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1456 ( N_VDD_c_1174_p N_CLK_c_5061_n ) capacitor c=7.81728e-19 //x=31.185 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1457 ( N_VDD_c_1479_p N_CLK_c_5061_n ) capacitor c=0.00205475f //x=32.76 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1458 ( N_VDD_c_1480_p N_CLK_c_5061_n ) capacitor c=0.00209689f //x=33.635 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1459 ( N_VDD_c_1209_p N_CLK_c_5061_n ) capacitor c=7.81728e-19 //x=34.515 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1460 ( N_VDD_c_945_n N_CLK_c_5061_n ) capacitor c=0.0389825f //x=26.27 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1461 ( N_VDD_c_946_n N_CLK_c_5061_n ) capacitor c=0.0389825f //x=29.6 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1462 ( N_VDD_c_947_n N_CLK_c_5061_n ) capacitor c=0.0389825f //x=32.93 \
 //y=7.4 //x2=34.665 //y2=4.44
cc_1463 ( N_VDD_M77_noxref_s N_CLK_c_5061_n ) capacitor c=0.00541054f \
 //x=26.925 //y=5.02 //x2=34.665 //y2=4.44
cc_1464 ( N_VDD_M80_noxref_d N_CLK_c_5061_n ) capacitor c=6.7165e-19 \
 //x=28.675 //y=5.02 //x2=34.665 //y2=4.44
cc_1465 ( N_VDD_M81_noxref_s N_CLK_c_5061_n ) capacitor c=0.00541054f \
 //x=30.255 //y=5.02 //x2=34.665 //y2=4.44
cc_1466 ( N_VDD_M84_noxref_d N_CLK_c_5061_n ) capacitor c=6.7165e-19 \
 //x=32.005 //y=5.02 //x2=34.665 //y2=4.44
cc_1467 ( N_VDD_M85_noxref_s N_CLK_c_5061_n ) capacitor c=0.00541054f \
 //x=33.585 //y=5.02 //x2=34.665 //y2=4.44
cc_1468 ( N_VDD_c_960_p N_CLK_c_5079_n ) capacitor c=0.0526102f //x=73.63 \
 //y=7.4 //x2=23.795 //y2=4.44
cc_1469 ( N_VDD_c_1491_p N_CLK_c_5079_n ) capacitor c=0.00205475f //x=17.96 \
 //y=7.4 //x2=23.795 //y2=4.44
cc_1470 ( N_VDD_c_1492_p N_CLK_c_5079_n ) capacitor c=0.00209689f //x=18.835 \
 //y=7.4 //x2=23.795 //y2=4.44
cc_1471 ( N_VDD_c_1085_p N_CLK_c_5079_n ) capacitor c=7.81728e-19 //x=19.715 \
 //y=7.4 //x2=23.795 //y2=4.44
cc_1472 ( N_VDD_c_1494_p N_CLK_c_5079_n ) capacitor c=0.00205475f //x=21.29 \
 //y=7.4 //x2=23.795 //y2=4.44
cc_1473 ( N_VDD_c_1495_p N_CLK_c_5079_n ) capacitor c=0.00328994f //x=22.465 \
 //y=7.4 //x2=23.795 //y2=4.44
cc_1474 ( N_VDD_c_1228_p N_CLK_c_5079_n ) capacitor c=0.00135925f //x=23.345 \
 //y=7.4 //x2=23.795 //y2=4.44
cc_1475 ( N_VDD_c_943_n N_CLK_c_5079_n ) capacitor c=0.0389825f //x=18.13 \
 //y=7.4 //x2=23.795 //y2=4.44
cc_1476 ( N_VDD_c_944_n N_CLK_c_5079_n ) capacitor c=0.0404757f //x=21.46 \
 //y=7.4 //x2=23.795 //y2=4.44
cc_1477 ( N_VDD_M66_noxref_d N_CLK_c_5079_n ) capacitor c=6.7165e-19 \
 //x=17.205 //y=5.02 //x2=23.795 //y2=4.44
cc_1478 ( N_VDD_M67_noxref_s N_CLK_c_5079_n ) capacitor c=0.00541054f \
 //x=18.785 //y=5.02 //x2=23.795 //y2=4.44
cc_1479 ( N_VDD_M70_noxref_d N_CLK_c_5079_n ) capacitor c=6.7165e-19 \
 //x=20.535 //y=5.02 //x2=23.795 //y2=4.44
cc_1480 ( N_VDD_M71_noxref_s N_CLK_c_5079_n ) capacitor c=0.00179496f \
 //x=22.415 //y=5.02 //x2=23.795 //y2=4.44
cc_1481 ( N_VDD_c_960_p N_CLK_c_5092_n ) capacitor c=0.0758142f //x=73.63 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1482 ( N_VDD_c_1504_p N_CLK_c_5092_n ) capacitor c=0.00205475f //x=36.09 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1483 ( N_VDD_c_1505_p N_CLK_c_5092_n ) capacitor c=0.00209689f //x=36.965 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1484 ( N_VDD_c_1246_p N_CLK_c_5092_n ) capacitor c=7.81728e-19 //x=37.845 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1485 ( N_VDD_c_1507_p N_CLK_c_5092_n ) capacitor c=0.00205475f //x=39.42 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1486 ( N_VDD_c_1508_p N_CLK_c_5092_n ) capacitor c=0.00209689f //x=40.295 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1487 ( N_VDD_c_1286_p N_CLK_c_5092_n ) capacitor c=7.81728e-19 //x=41.175 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1488 ( N_VDD_c_1510_p N_CLK_c_5092_n ) capacitor c=0.00205475f //x=42.75 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1489 ( N_VDD_c_1511_p N_CLK_c_5092_n ) capacitor c=0.00328994f //x=43.925 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1490 ( N_VDD_c_1512_p N_CLK_c_5092_n ) capacitor c=0.00135925f //x=44.805 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1491 ( N_VDD_c_948_n N_CLK_c_5092_n ) capacitor c=0.0389825f //x=36.26 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1492 ( N_VDD_c_949_n N_CLK_c_5092_n ) capacitor c=0.0389825f //x=39.59 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1493 ( N_VDD_c_950_n N_CLK_c_5092_n ) capacitor c=0.0404757f //x=42.92 \
 //y=7.4 //x2=45.025 //y2=4.44
cc_1494 ( N_VDD_M88_noxref_d N_CLK_c_5092_n ) capacitor c=6.7165e-19 \
 //x=35.335 //y=5.02 //x2=45.025 //y2=4.44
cc_1495 ( N_VDD_M89_noxref_s N_CLK_c_5092_n ) capacitor c=0.00541054f \
 //x=36.915 //y=5.02 //x2=45.025 //y2=4.44
cc_1496 ( N_VDD_M92_noxref_d N_CLK_c_5092_n ) capacitor c=6.7165e-19 \
 //x=38.665 //y=5.02 //x2=45.025 //y2=4.44
cc_1497 ( N_VDD_M93_noxref_s N_CLK_c_5092_n ) capacitor c=0.00541054f \
 //x=40.245 //y=5.02 //x2=45.025 //y2=4.44
cc_1498 ( N_VDD_M96_noxref_d N_CLK_c_5092_n ) capacitor c=6.7165e-19 \
 //x=41.995 //y=5.02 //x2=45.025 //y2=4.44
cc_1499 ( N_VDD_M97_noxref_s N_CLK_c_5092_n ) capacitor c=0.00179496f \
 //x=43.875 //y=5.02 //x2=45.025 //y2=4.44
cc_1500 ( N_VDD_c_960_p N_CLK_c_5111_n ) capacitor c=0.00123805f //x=73.63 \
 //y=7.4 //x2=34.895 //y2=4.44
cc_1501 ( N_VDD_c_960_p N_CLK_c_5112_n ) capacitor c=0.0824294f //x=73.63 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1502 ( N_VDD_c_1524_p N_CLK_c_5112_n ) capacitor c=0.00258496f //x=47.56 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1503 ( N_VDD_c_1525_p N_CLK_c_5112_n ) capacitor c=0.00209689f //x=48.435 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1504 ( N_VDD_c_1380_p N_CLK_c_5112_n ) capacitor c=7.81728e-19 //x=49.315 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1505 ( N_VDD_c_1527_p N_CLK_c_5112_n ) capacitor c=0.00205475f //x=50.89 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1506 ( N_VDD_c_1528_p N_CLK_c_5112_n ) capacitor c=0.00209689f //x=51.765 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1507 ( N_VDD_c_1392_p N_CLK_c_5112_n ) capacitor c=7.81728e-19 //x=52.645 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1508 ( N_VDD_c_1530_p N_CLK_c_5112_n ) capacitor c=0.00205475f //x=54.22 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1509 ( N_VDD_c_1531_p N_CLK_c_5112_n ) capacitor c=0.00209689f //x=55.095 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1510 ( N_VDD_c_1427_p N_CLK_c_5112_n ) capacitor c=7.81728e-19 //x=55.975 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1511 ( N_VDD_c_951_n N_CLK_c_5112_n ) capacitor c=0.0389825f //x=47.73 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1512 ( N_VDD_c_952_n N_CLK_c_5112_n ) capacitor c=0.0389825f //x=51.06 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1513 ( N_VDD_c_953_n N_CLK_c_5112_n ) capacitor c=0.0389825f //x=54.39 \
 //y=7.4 //x2=56.125 //y2=4.44
cc_1514 ( N_VDD_M103_noxref_s N_CLK_c_5112_n ) capacitor c=0.00541054f \
 //x=48.385 //y=5.02 //x2=56.125 //y2=4.44
cc_1515 ( N_VDD_M106_noxref_d N_CLK_c_5112_n ) capacitor c=6.7165e-19 \
 //x=50.135 //y=5.02 //x2=56.125 //y2=4.44
cc_1516 ( N_VDD_M107_noxref_s N_CLK_c_5112_n ) capacitor c=0.00541054f \
 //x=51.715 //y=5.02 //x2=56.125 //y2=4.44
cc_1517 ( N_VDD_M110_noxref_d N_CLK_c_5112_n ) capacitor c=6.7165e-19 \
 //x=53.465 //y=5.02 //x2=56.125 //y2=4.44
cc_1518 ( N_VDD_M111_noxref_s N_CLK_c_5112_n ) capacitor c=0.00541054f \
 //x=55.045 //y=5.02 //x2=56.125 //y2=4.44
cc_1519 ( N_VDD_c_960_p N_CLK_c_5130_n ) capacitor c=0.00120845f //x=73.63 \
 //y=7.4 //x2=45.255 //y2=4.44
cc_1520 ( N_VDD_c_960_p N_CLK_c_5025_n ) capacitor c=2.03287e-19 //x=73.63 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_1521 ( N_VDD_c_937_n N_CLK_c_5025_n ) capacitor c=9.53425e-19 //x=0.74 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_1522 ( N_VDD_c_941_n N_CLK_c_5026_n ) capacitor c=5.27482e-19 //x=11.47 \
 //y=7.4 //x2=13.32 //y2=2.08
cc_1523 ( N_VDD_c_942_n N_CLK_c_5026_n ) capacitor c=4.23917e-19 //x=14.8 \
 //y=7.4 //x2=13.32 //y2=2.08
cc_1524 ( N_VDD_c_960_p N_CLK_c_5028_n ) capacitor c=2.03287e-19 //x=73.63 \
 //y=7.4 //x2=23.68 //y2=2.08
cc_1525 ( N_VDD_c_944_n N_CLK_c_5028_n ) capacitor c=7.21466e-19 //x=21.46 \
 //y=7.4 //x2=23.68 //y2=2.08
cc_1526 ( N_VDD_c_947_n N_CLK_c_5029_n ) capacitor c=5.27482e-19 //x=32.93 \
 //y=7.4 //x2=34.78 //y2=2.08
cc_1527 ( N_VDD_c_948_n N_CLK_c_5029_n ) capacitor c=3.91923e-19 //x=36.26 \
 //y=7.4 //x2=34.78 //y2=2.08
cc_1528 ( N_VDD_c_960_p N_CLK_c_5031_n ) capacitor c=2.03287e-19 //x=73.63 \
 //y=7.4 //x2=45.14 //y2=2.08
cc_1529 ( N_VDD_c_950_n N_CLK_c_5031_n ) capacitor c=7.21466e-19 //x=42.92 \
 //y=7.4 //x2=45.14 //y2=2.08
cc_1530 ( N_VDD_c_953_n N_CLK_c_5032_n ) capacitor c=5.27482e-19 //x=54.39 \
 //y=7.4 //x2=56.24 //y2=2.08
cc_1531 ( N_VDD_c_954_n N_CLK_c_5032_n ) capacitor c=7.54518e-19 //x=57.72 \
 //y=7.4 //x2=56.24 //y2=2.08
cc_1532 ( N_VDD_c_1028_p N_CLK_M47_noxref_g ) capacitor c=0.00676195f \
 //x=2.765 //y=7.4 //x2=2.19 //y2=6.02
cc_1533 ( N_VDD_M46_noxref_d N_CLK_M47_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=2.19 //y2=6.02
cc_1534 ( N_VDD_c_1028_p N_CLK_M48_noxref_g ) capacitor c=0.00675175f \
 //x=2.765 //y=7.4 //x2=2.63 //y2=6.02
cc_1535 ( N_VDD_M48_noxref_d N_CLK_M48_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=2.63 //y2=6.02
cc_1536 ( N_VDD_c_1121_p N_CLK_M61_noxref_g ) capacitor c=0.00673971f \
 //x=13.935 //y=7.4 //x2=13.36 //y2=6.02
cc_1537 ( N_VDD_M60_noxref_d N_CLK_M61_noxref_g ) capacitor c=0.015318f \
 //x=12.995 //y=5.02 //x2=13.36 //y2=6.02
cc_1538 ( N_VDD_c_1121_p N_CLK_M62_noxref_g ) capacitor c=0.00672952f \
 //x=13.935 //y=7.4 //x2=13.8 //y2=6.02
cc_1539 ( N_VDD_c_942_n N_CLK_M62_noxref_g ) capacitor c=0.00864163f //x=14.8 \
 //y=7.4 //x2=13.8 //y2=6.02
cc_1540 ( N_VDD_M62_noxref_d N_CLK_M62_noxref_g ) capacitor c=0.0430452f \
 //x=13.875 //y=5.02 //x2=13.8 //y2=6.02
cc_1541 ( N_VDD_c_1229_p N_CLK_M73_noxref_g ) capacitor c=0.00676195f \
 //x=24.225 //y=7.4 //x2=23.65 //y2=6.02
cc_1542 ( N_VDD_M72_noxref_d N_CLK_M73_noxref_g ) capacitor c=0.015318f \
 //x=23.285 //y=5.02 //x2=23.65 //y2=6.02
cc_1543 ( N_VDD_c_1229_p N_CLK_M74_noxref_g ) capacitor c=0.00675175f \
 //x=24.225 //y=7.4 //x2=24.09 //y2=6.02
cc_1544 ( N_VDD_M74_noxref_d N_CLK_M74_noxref_g ) capacitor c=0.015318f \
 //x=24.165 //y=5.02 //x2=24.09 //y2=6.02
cc_1545 ( N_VDD_c_1318_p N_CLK_M87_noxref_g ) capacitor c=0.00673971f \
 //x=35.395 //y=7.4 //x2=34.82 //y2=6.02
cc_1546 ( N_VDD_M86_noxref_d N_CLK_M87_noxref_g ) capacitor c=0.015318f \
 //x=34.455 //y=5.02 //x2=34.82 //y2=6.02
cc_1547 ( N_VDD_c_1318_p N_CLK_M88_noxref_g ) capacitor c=0.00672952f \
 //x=35.395 //y=7.4 //x2=35.26 //y2=6.02
cc_1548 ( N_VDD_c_948_n N_CLK_M88_noxref_g ) capacitor c=0.00864163f //x=36.26 \
 //y=7.4 //x2=35.26 //y2=6.02
cc_1549 ( N_VDD_M88_noxref_d N_CLK_M88_noxref_g ) capacitor c=0.0430452f \
 //x=35.335 //y=5.02 //x2=35.26 //y2=6.02
cc_1550 ( N_VDD_c_1572_p N_CLK_M99_noxref_g ) capacitor c=0.00676195f \
 //x=45.685 //y=7.4 //x2=45.11 //y2=6.02
cc_1551 ( N_VDD_M98_noxref_d N_CLK_M99_noxref_g ) capacitor c=0.015318f \
 //x=44.745 //y=5.02 //x2=45.11 //y2=6.02
cc_1552 ( N_VDD_c_1572_p N_CLK_M100_noxref_g ) capacitor c=0.00675175f \
 //x=45.685 //y=7.4 //x2=45.55 //y2=6.02
cc_1553 ( N_VDD_M100_noxref_d N_CLK_M100_noxref_g ) capacitor c=0.015318f \
 //x=45.625 //y=5.02 //x2=45.55 //y2=6.02
cc_1554 ( N_VDD_c_1576_p N_CLK_M113_noxref_g ) capacitor c=0.00673971f \
 //x=56.855 //y=7.4 //x2=56.28 //y2=6.02
cc_1555 ( N_VDD_M112_noxref_d N_CLK_M113_noxref_g ) capacitor c=0.015318f \
 //x=55.915 //y=5.02 //x2=56.28 //y2=6.02
cc_1556 ( N_VDD_c_1576_p N_CLK_M114_noxref_g ) capacitor c=0.00672952f \
 //x=56.855 //y=7.4 //x2=56.72 //y2=6.02
cc_1557 ( N_VDD_c_954_n N_CLK_M114_noxref_g ) capacitor c=0.00864163f \
 //x=57.72 //y=7.4 //x2=56.72 //y2=6.02
cc_1558 ( N_VDD_M114_noxref_d N_CLK_M114_noxref_g ) capacitor c=0.0430452f \
 //x=56.795 //y=5.02 //x2=56.72 //y2=6.02
cc_1559 ( N_VDD_c_960_p N_noxref_17_c_5801_n ) capacitor c=0.00444751f \
 //x=73.63 //y=7.4 //x2=45.245 //y2=5.155
cc_1560 ( N_VDD_c_1512_p N_noxref_17_c_5801_n ) capacitor c=4.31931e-19 \
 //x=44.805 //y=7.4 //x2=45.245 //y2=5.155
cc_1561 ( N_VDD_c_1572_p N_noxref_17_c_5801_n ) capacitor c=4.31906e-19 \
 //x=45.685 //y=7.4 //x2=45.245 //y2=5.155
cc_1562 ( N_VDD_M98_noxref_d N_noxref_17_c_5801_n ) capacitor c=0.0112985f \
 //x=44.745 //y=5.02 //x2=45.245 //y2=5.155
cc_1563 ( N_VDD_c_950_n N_noxref_17_c_5805_n ) capacitor c=0.00863585f \
 //x=42.92 //y=7.4 //x2=44.535 //y2=5.155
cc_1564 ( N_VDD_M97_noxref_s N_noxref_17_c_5805_n ) capacitor c=0.0831083f \
 //x=43.875 //y=5.02 //x2=44.535 //y2=5.155
cc_1565 ( N_VDD_c_960_p N_noxref_17_c_5807_n ) capacitor c=0.0044221f \
 //x=73.63 //y=7.4 //x2=46.125 //y2=5.155
cc_1566 ( N_VDD_c_1572_p N_noxref_17_c_5807_n ) capacitor c=4.31931e-19 \
 //x=45.685 //y=7.4 //x2=46.125 //y2=5.155
cc_1567 ( N_VDD_c_1394_p N_noxref_17_c_5807_n ) capacitor c=4.31931e-19 \
 //x=46.565 //y=7.4 //x2=46.125 //y2=5.155
cc_1568 ( N_VDD_M100_noxref_d N_noxref_17_c_5807_n ) capacitor c=0.0112985f \
 //x=45.625 //y=5.02 //x2=46.125 //y2=5.155
cc_1569 ( N_VDD_c_960_p N_noxref_17_c_5811_n ) capacitor c=0.00434174f \
 //x=73.63 //y=7.4 //x2=46.905 //y2=5.155
cc_1570 ( N_VDD_c_1394_p N_noxref_17_c_5811_n ) capacitor c=7.46626e-19 \
 //x=46.565 //y=7.4 //x2=46.905 //y2=5.155
cc_1571 ( N_VDD_c_1524_p N_noxref_17_c_5811_n ) capacitor c=0.00198565f \
 //x=47.56 //y=7.4 //x2=46.905 //y2=5.155
cc_1572 ( N_VDD_M102_noxref_d N_noxref_17_c_5811_n ) capacitor c=0.0112985f \
 //x=46.505 //y=5.02 //x2=46.905 //y2=5.155
cc_1573 ( N_VDD_c_951_n N_noxref_17_c_5815_n ) capacitor c=0.0426341f \
 //x=47.73 //y=7.4 //x2=46.99 //y2=3.7
cc_1574 ( N_VDD_c_960_p N_noxref_17_c_5778_n ) capacitor c=0.00125279f \
 //x=73.63 //y=7.4 //x2=48.84 //y2=2.08
cc_1575 ( N_VDD_c_1380_p N_noxref_17_c_5778_n ) capacitor c=2.87256e-19 \
 //x=49.315 //y=7.4 //x2=48.84 //y2=2.08
cc_1576 ( N_VDD_c_951_n N_noxref_17_c_5778_n ) capacitor c=0.0134665f \
 //x=47.73 //y=7.4 //x2=48.84 //y2=2.08
cc_1577 ( N_VDD_c_960_p N_noxref_17_c_5779_n ) capacitor c=0.00126216f \
 //x=73.63 //y=7.4 //x2=58.83 //y2=2.08
cc_1578 ( N_VDD_c_1600_p N_noxref_17_c_5779_n ) capacitor c=2.87813e-19 \
 //x=59.305 //y=7.4 //x2=58.83 //y2=2.08
cc_1579 ( N_VDD_c_954_n N_noxref_17_c_5779_n ) capacitor c=0.015485f //x=57.72 \
 //y=7.4 //x2=58.83 //y2=2.08
cc_1580 ( N_VDD_c_1380_p N_noxref_17_M103_noxref_g ) capacitor c=0.00726866f \
 //x=49.315 //y=7.4 //x2=48.74 //y2=6.02
cc_1581 ( N_VDD_M103_noxref_s N_noxref_17_M103_noxref_g ) capacitor \
 c=0.054195f //x=48.385 //y=5.02 //x2=48.74 //y2=6.02
cc_1582 ( N_VDD_c_1380_p N_noxref_17_M104_noxref_g ) capacitor c=0.00672952f \
 //x=49.315 //y=7.4 //x2=49.18 //y2=6.02
cc_1583 ( N_VDD_M104_noxref_d N_noxref_17_M104_noxref_g ) capacitor \
 c=0.015318f //x=49.255 //y=5.02 //x2=49.18 //y2=6.02
cc_1584 ( N_VDD_c_1600_p N_noxref_17_M115_noxref_g ) capacitor c=0.00726866f \
 //x=59.305 //y=7.4 //x2=58.73 //y2=6.02
cc_1585 ( N_VDD_M115_noxref_s N_noxref_17_M115_noxref_g ) capacitor \
 c=0.054195f //x=58.375 //y=5.02 //x2=58.73 //y2=6.02
cc_1586 ( N_VDD_c_1600_p N_noxref_17_M116_noxref_g ) capacitor c=0.00672952f \
 //x=59.305 //y=7.4 //x2=59.17 //y2=6.02
cc_1587 ( N_VDD_M116_noxref_d N_noxref_17_M116_noxref_g ) capacitor \
 c=0.015318f //x=59.245 //y=5.02 //x2=59.17 //y2=6.02
cc_1588 ( N_VDD_c_951_n N_noxref_17_c_5830_n ) capacitor c=0.015293f //x=47.73 \
 //y=7.4 //x2=48.84 //y2=4.7
cc_1589 ( N_VDD_c_954_n N_noxref_17_c_5831_n ) capacitor c=0.0149273f \
 //x=57.72 //y=7.4 //x2=58.83 //y2=4.7
cc_1590 ( N_VDD_c_960_p N_noxref_17_M97_noxref_d ) capacitor c=0.00275235f \
 //x=73.63 //y=7.4 //x2=44.305 //y2=5.02
cc_1591 ( N_VDD_c_1512_p N_noxref_17_M97_noxref_d ) capacitor c=0.014035f \
 //x=44.805 //y=7.4 //x2=44.305 //y2=5.02
cc_1592 ( N_VDD_M98_noxref_d N_noxref_17_M97_noxref_d ) capacitor c=0.0664752f \
 //x=44.745 //y=5.02 //x2=44.305 //y2=5.02
cc_1593 ( N_VDD_c_960_p N_noxref_17_M99_noxref_d ) capacitor c=0.00275186f \
 //x=73.63 //y=7.4 //x2=45.185 //y2=5.02
cc_1594 ( N_VDD_c_1572_p N_noxref_17_M99_noxref_d ) capacitor c=0.0140346f \
 //x=45.685 //y=7.4 //x2=45.185 //y2=5.02
cc_1595 ( N_VDD_c_951_n N_noxref_17_M99_noxref_d ) capacitor c=4.9285e-19 \
 //x=47.73 //y=7.4 //x2=45.185 //y2=5.02
cc_1596 ( N_VDD_M97_noxref_s N_noxref_17_M99_noxref_d ) capacitor \
 c=0.00130656f //x=43.875 //y=5.02 //x2=45.185 //y2=5.02
cc_1597 ( N_VDD_M98_noxref_d N_noxref_17_M99_noxref_d ) capacitor c=0.0664752f \
 //x=44.745 //y=5.02 //x2=45.185 //y2=5.02
cc_1598 ( N_VDD_M100_noxref_d N_noxref_17_M99_noxref_d ) capacitor \
 c=0.0664752f //x=45.625 //y=5.02 //x2=45.185 //y2=5.02
cc_1599 ( N_VDD_c_960_p N_noxref_17_M101_noxref_d ) capacitor c=0.00275235f \
 //x=73.63 //y=7.4 //x2=46.065 //y2=5.02
cc_1600 ( N_VDD_c_1394_p N_noxref_17_M101_noxref_d ) capacitor c=0.0137384f \
 //x=46.565 //y=7.4 //x2=46.065 //y2=5.02
cc_1601 ( N_VDD_c_951_n N_noxref_17_M101_noxref_d ) capacitor c=0.00939849f \
 //x=47.73 //y=7.4 //x2=46.065 //y2=5.02
cc_1602 ( N_VDD_M100_noxref_d N_noxref_17_M101_noxref_d ) capacitor \
 c=0.0664752f //x=45.625 //y=5.02 //x2=46.065 //y2=5.02
cc_1603 ( N_VDD_M102_noxref_d N_noxref_17_M101_noxref_d ) capacitor \
 c=0.0664752f //x=46.505 //y=5.02 //x2=46.065 //y2=5.02
cc_1604 ( N_VDD_M103_noxref_s N_noxref_17_M101_noxref_d ) capacitor \
 c=4.52683e-19 //x=48.385 //y=5.02 //x2=46.065 //y2=5.02
cc_1605 ( N_VDD_c_960_p N_noxref_18_c_6048_n ) capacitor c=0.0143704f \
 //x=73.63 //y=7.4 //x2=62.045 //y2=4.44
cc_1606 ( N_VDD_c_1628_p N_noxref_18_c_6048_n ) capacitor c=0.00196877f \
 //x=60.88 //y=7.4 //x2=62.045 //y2=4.44
cc_1607 ( N_VDD_c_1629_p N_noxref_18_c_6048_n ) capacitor c=0.00209689f \
 //x=61.755 //y=7.4 //x2=62.045 //y2=4.44
cc_1608 ( N_VDD_c_1630_p N_noxref_18_c_6048_n ) capacitor c=9.71854e-19 \
 //x=62.635 //y=7.4 //x2=62.045 //y2=4.44
cc_1609 ( N_VDD_c_955_n N_noxref_18_c_6048_n ) capacitor c=0.0397717f \
 //x=61.05 //y=7.4 //x2=62.045 //y2=4.44
cc_1610 ( N_VDD_M119_noxref_s N_noxref_18_c_6048_n ) capacitor c=0.00541054f \
 //x=61.705 //y=5.02 //x2=62.045 //y2=4.44
cc_1611 ( N_VDD_c_960_p N_noxref_18_c_6054_n ) capacitor c=0.00215478f \
 //x=73.63 //y=7.4 //x2=60.425 //y2=4.44
cc_1612 ( N_VDD_c_955_n N_noxref_18_c_6054_n ) capacitor c=0.00102529f \
 //x=61.05 //y=7.4 //x2=60.425 //y2=4.44
cc_1613 ( N_VDD_M118_noxref_d N_noxref_18_c_6054_n ) capacitor c=6.90267e-19 \
 //x=60.125 //y=5.02 //x2=60.425 //y2=4.44
cc_1614 ( N_VDD_c_960_p N_noxref_18_c_6057_n ) capacitor c=0.00460134f \
 //x=73.63 //y=7.4 //x2=59.745 //y2=5.2
cc_1615 ( N_VDD_c_1600_p N_noxref_18_c_6057_n ) capacitor c=4.48705e-19 \
 //x=59.305 //y=7.4 //x2=59.745 //y2=5.2
cc_1616 ( N_VDD_c_1638_p N_noxref_18_c_6057_n ) capacitor c=4.48705e-19 \
 //x=60.185 //y=7.4 //x2=59.745 //y2=5.2
cc_1617 ( N_VDD_M116_noxref_d N_noxref_18_c_6057_n ) capacitor c=0.0126924f \
 //x=59.245 //y=5.02 //x2=59.745 //y2=5.2
cc_1618 ( N_VDD_c_954_n N_noxref_18_c_6061_n ) capacitor c=0.00985474f \
 //x=57.72 //y=7.4 //x2=59.035 //y2=5.2
cc_1619 ( N_VDD_M115_noxref_s N_noxref_18_c_6061_n ) capacitor c=0.087833f \
 //x=58.375 //y=5.02 //x2=59.035 //y2=5.2
cc_1620 ( N_VDD_c_960_p N_noxref_18_c_6063_n ) capacitor c=0.00304119f \
 //x=73.63 //y=7.4 //x2=60.225 //y2=5.2
cc_1621 ( N_VDD_c_1638_p N_noxref_18_c_6063_n ) capacitor c=7.73167e-19 \
 //x=60.185 //y=7.4 //x2=60.225 //y2=5.2
cc_1622 ( N_VDD_M118_noxref_d N_noxref_18_c_6063_n ) capacitor c=0.0151251f \
 //x=60.125 //y=5.02 //x2=60.225 //y2=5.2
cc_1623 ( N_VDD_M119_noxref_s N_noxref_18_c_6063_n ) capacitor c=2.44532e-19 \
 //x=61.705 //y=5.02 //x2=60.225 //y2=5.2
cc_1624 ( N_VDD_c_954_n N_noxref_18_c_6033_n ) capacitor c=0.00151618f \
 //x=57.72 //y=7.4 //x2=60.31 //y2=4.44
cc_1625 ( N_VDD_c_955_n N_noxref_18_c_6033_n ) capacitor c=0.042956f //x=61.05 \
 //y=7.4 //x2=60.31 //y2=4.44
cc_1626 ( N_VDD_c_960_p N_noxref_18_c_6034_n ) capacitor c=0.00125199f \
 //x=73.63 //y=7.4 //x2=62.16 //y2=2.08
cc_1627 ( N_VDD_c_1630_p N_noxref_18_c_6034_n ) capacitor c=2.87208e-19 \
 //x=62.635 //y=7.4 //x2=62.16 //y2=2.08
cc_1628 ( N_VDD_c_955_n N_noxref_18_c_6034_n ) capacitor c=0.0131445f \
 //x=61.05 //y=7.4 //x2=62.16 //y2=2.08
cc_1629 ( N_VDD_c_1630_p N_noxref_18_M119_noxref_g ) capacitor c=0.00726866f \
 //x=62.635 //y=7.4 //x2=62.06 //y2=6.02
cc_1630 ( N_VDD_M119_noxref_s N_noxref_18_M119_noxref_g ) capacitor \
 c=0.054195f //x=61.705 //y=5.02 //x2=62.06 //y2=6.02
cc_1631 ( N_VDD_c_1630_p N_noxref_18_M120_noxref_g ) capacitor c=0.00672952f \
 //x=62.635 //y=7.4 //x2=62.5 //y2=6.02
cc_1632 ( N_VDD_M120_noxref_d N_noxref_18_M120_noxref_g ) capacitor \
 c=0.015318f //x=62.575 //y=5.02 //x2=62.5 //y2=6.02
cc_1633 ( N_VDD_c_955_n N_noxref_18_c_6076_n ) capacitor c=0.0149273f \
 //x=61.05 //y=7.4 //x2=62.16 //y2=4.7
cc_1634 ( N_VDD_c_960_p N_noxref_18_M115_noxref_d ) capacitor c=0.00285083f \
 //x=73.63 //y=7.4 //x2=58.805 //y2=5.02
cc_1635 ( N_VDD_c_1600_p N_noxref_18_M115_noxref_d ) capacitor c=0.0140984f \
 //x=59.305 //y=7.4 //x2=58.805 //y2=5.02
cc_1636 ( N_VDD_c_955_n N_noxref_18_M115_noxref_d ) capacitor c=6.94454e-19 \
 //x=61.05 //y=7.4 //x2=58.805 //y2=5.02
cc_1637 ( N_VDD_M116_noxref_d N_noxref_18_M115_noxref_d ) capacitor \
 c=0.0664752f //x=59.245 //y=5.02 //x2=58.805 //y2=5.02
cc_1638 ( N_VDD_c_960_p N_noxref_18_M117_noxref_d ) capacitor c=0.00285083f \
 //x=73.63 //y=7.4 //x2=59.685 //y2=5.02
cc_1639 ( N_VDD_c_1638_p N_noxref_18_M117_noxref_d ) capacitor c=0.0140984f \
 //x=60.185 //y=7.4 //x2=59.685 //y2=5.02
cc_1640 ( N_VDD_c_955_n N_noxref_18_M117_noxref_d ) capacitor c=0.0120541f \
 //x=61.05 //y=7.4 //x2=59.685 //y2=5.02
cc_1641 ( N_VDD_M115_noxref_s N_noxref_18_M117_noxref_d ) capacitor \
 c=0.00111971f //x=58.375 //y=5.02 //x2=59.685 //y2=5.02
cc_1642 ( N_VDD_M116_noxref_d N_noxref_18_M117_noxref_d ) capacitor \
 c=0.0664752f //x=59.245 //y=5.02 //x2=59.685 //y2=5.02
cc_1643 ( N_VDD_M118_noxref_d N_noxref_18_M117_noxref_d ) capacitor \
 c=0.0664752f //x=60.125 //y=5.02 //x2=59.685 //y2=5.02
cc_1644 ( N_VDD_M119_noxref_s N_noxref_18_M117_noxref_d ) capacitor \
 c=4.54516e-19 //x=61.705 //y=5.02 //x2=59.685 //y2=5.02
cc_1645 ( N_VDD_c_951_n N_noxref_19_c_6210_n ) capacitor c=0.0140578f \
 //x=47.73 //y=7.4 //x2=52.795 //y2=4.07
cc_1646 ( N_VDD_c_952_n N_noxref_19_c_6210_n ) capacitor c=0.0140578f \
 //x=51.06 //y=7.4 //x2=52.795 //y2=4.07
cc_1647 ( N_VDD_c_950_n N_noxref_19_c_6212_n ) capacitor c=0.00116746f \
 //x=42.92 //y=7.4 //x2=44.145 //y2=4.07
cc_1648 ( N_VDD_c_960_p N_noxref_19_c_6213_n ) capacitor c=0.0158405f \
 //x=73.63 //y=7.4 //x2=56.865 //y2=4.07
cc_1649 ( N_VDD_c_953_n N_noxref_19_c_6213_n ) capacitor c=0.0140578f \
 //x=54.39 //y=7.4 //x2=56.865 //y2=4.07
cc_1650 ( N_VDD_c_960_p N_noxref_19_c_6215_n ) capacitor c=0.0332843f \
 //x=73.63 //y=7.4 //x2=62.785 //y2=4.07
cc_1651 ( N_VDD_c_1673_p N_noxref_19_c_6215_n ) capacitor c=0.00161566f \
 //x=57.55 //y=7.4 //x2=62.785 //y2=4.07
cc_1652 ( N_VDD_c_1674_p N_noxref_19_c_6215_n ) capacitor c=0.00172186f \
 //x=58.425 //y=7.4 //x2=62.785 //y2=4.07
cc_1653 ( N_VDD_c_1600_p N_noxref_19_c_6215_n ) capacitor c=6.61469e-19 \
 //x=59.305 //y=7.4 //x2=62.785 //y2=4.07
cc_1654 ( N_VDD_c_954_n N_noxref_19_c_6215_n ) capacitor c=0.0269494f \
 //x=57.72 //y=7.4 //x2=62.785 //y2=4.07
cc_1655 ( N_VDD_c_955_n N_noxref_19_c_6215_n ) capacitor c=0.0140578f \
 //x=61.05 //y=7.4 //x2=62.785 //y2=4.07
cc_1656 ( N_VDD_M115_noxref_s N_noxref_19_c_6215_n ) capacitor c=0.00363031f \
 //x=58.375 //y=5.02 //x2=62.785 //y2=4.07
cc_1657 ( N_VDD_c_960_p N_noxref_19_c_6222_n ) capacitor c=0.00172491f \
 //x=73.63 //y=7.4 //x2=57.095 //y2=4.07
cc_1658 ( N_VDD_c_954_n N_noxref_19_c_6222_n ) capacitor c=0.00104972f \
 //x=57.72 //y=7.4 //x2=57.095 //y2=4.07
cc_1659 ( N_VDD_M114_noxref_d N_noxref_19_c_6222_n ) capacitor c=5.14736e-19 \
 //x=56.795 //y=5.02 //x2=57.095 //y2=4.07
cc_1660 ( N_VDD_c_960_p N_noxref_19_c_6190_n ) capacitor c=9.10347e-19 \
 //x=73.63 //y=7.4 //x2=44.03 //y2=2.08
cc_1661 ( N_VDD_c_950_n N_noxref_19_c_6190_n ) capacitor c=0.0137129f \
 //x=42.92 //y=7.4 //x2=44.03 //y2=2.08
cc_1662 ( N_VDD_M97_noxref_s N_noxref_19_c_6190_n ) capacitor c=0.0120327f \
 //x=43.875 //y=5.02 //x2=44.03 //y2=2.08
cc_1663 ( N_VDD_c_952_n N_noxref_19_c_6191_n ) capacitor c=4.57806e-19 \
 //x=51.06 //y=7.4 //x2=52.91 //y2=2.08
cc_1664 ( N_VDD_c_953_n N_noxref_19_c_6191_n ) capacitor c=3.69525e-19 \
 //x=54.39 //y=7.4 //x2=52.91 //y2=2.08
cc_1665 ( N_VDD_c_960_p N_noxref_19_c_6230_n ) capacitor c=0.00453473f \
 //x=73.63 //y=7.4 //x2=56.415 //y2=5.2
cc_1666 ( N_VDD_c_1427_p N_noxref_19_c_6230_n ) capacitor c=4.48391e-19 \
 //x=55.975 //y=7.4 //x2=56.415 //y2=5.2
cc_1667 ( N_VDD_c_1576_p N_noxref_19_c_6230_n ) capacitor c=4.48377e-19 \
 //x=56.855 //y=7.4 //x2=56.415 //y2=5.2
cc_1668 ( N_VDD_M112_noxref_d N_noxref_19_c_6230_n ) capacitor c=0.0124506f \
 //x=55.915 //y=5.02 //x2=56.415 //y2=5.2
cc_1669 ( N_VDD_c_953_n N_noxref_19_c_6234_n ) capacitor c=0.00985474f \
 //x=54.39 //y=7.4 //x2=55.705 //y2=5.2
cc_1670 ( N_VDD_M111_noxref_s N_noxref_19_c_6234_n ) capacitor c=0.087833f \
 //x=55.045 //y=5.02 //x2=55.705 //y2=5.2
cc_1671 ( N_VDD_c_960_p N_noxref_19_c_6236_n ) capacitor c=0.00307016f \
 //x=73.63 //y=7.4 //x2=56.895 //y2=5.2
cc_1672 ( N_VDD_c_1576_p N_noxref_19_c_6236_n ) capacitor c=7.73167e-19 \
 //x=56.855 //y=7.4 //x2=56.895 //y2=5.2
cc_1673 ( N_VDD_M114_noxref_d N_noxref_19_c_6236_n ) capacitor c=0.016133f \
 //x=56.795 //y=5.02 //x2=56.895 //y2=5.2
cc_1674 ( N_VDD_M115_noxref_s N_noxref_19_c_6236_n ) capacitor c=2.44532e-19 \
 //x=58.375 //y=5.02 //x2=56.895 //y2=5.2
cc_1675 ( N_VDD_c_953_n N_noxref_19_c_6194_n ) capacitor c=0.00151618f \
 //x=54.39 //y=7.4 //x2=56.98 //y2=4.07
cc_1676 ( N_VDD_c_954_n N_noxref_19_c_6194_n ) capacitor c=0.0448479f \
 //x=57.72 //y=7.4 //x2=56.98 //y2=4.07
cc_1677 ( N_VDD_c_955_n N_noxref_19_c_6195_n ) capacitor c=7.9392e-19 \
 //x=61.05 //y=7.4 //x2=62.9 //y2=2.08
cc_1678 ( N_VDD_c_956_n N_noxref_19_c_6195_n ) capacitor c=0.00120485f \
 //x=64.38 //y=7.4 //x2=62.9 //y2=2.08
cc_1679 ( N_VDD_c_1512_p N_noxref_19_M97_noxref_g ) capacitor c=0.00749687f \
 //x=44.805 //y=7.4 //x2=44.23 //y2=6.02
cc_1680 ( N_VDD_M97_noxref_s N_noxref_19_M97_noxref_g ) capacitor c=0.0477201f \
 //x=43.875 //y=5.02 //x2=44.23 //y2=6.02
cc_1681 ( N_VDD_c_1512_p N_noxref_19_M98_noxref_g ) capacitor c=0.00675175f \
 //x=44.805 //y=7.4 //x2=44.67 //y2=6.02
cc_1682 ( N_VDD_M98_noxref_d N_noxref_19_M98_noxref_g ) capacitor c=0.015318f \
 //x=44.745 //y=5.02 //x2=44.67 //y2=6.02
cc_1683 ( N_VDD_c_1416_p N_noxref_19_M109_noxref_g ) capacitor c=0.00673971f \
 //x=53.525 //y=7.4 //x2=52.95 //y2=6.02
cc_1684 ( N_VDD_M108_noxref_d N_noxref_19_M109_noxref_g ) capacitor \
 c=0.015318f //x=52.585 //y=5.02 //x2=52.95 //y2=6.02
cc_1685 ( N_VDD_c_1416_p N_noxref_19_M110_noxref_g ) capacitor c=0.00672952f \
 //x=53.525 //y=7.4 //x2=53.39 //y2=6.02
cc_1686 ( N_VDD_c_953_n N_noxref_19_M110_noxref_g ) capacitor c=0.00864163f \
 //x=54.39 //y=7.4 //x2=53.39 //y2=6.02
cc_1687 ( N_VDD_M110_noxref_d N_noxref_19_M110_noxref_g ) capacitor \
 c=0.0430452f //x=53.465 //y=5.02 //x2=53.39 //y2=6.02
cc_1688 ( N_VDD_c_1710_p N_noxref_19_M121_noxref_g ) capacitor c=0.00673971f \
 //x=63.515 //y=7.4 //x2=62.94 //y2=6.02
cc_1689 ( N_VDD_M120_noxref_d N_noxref_19_M121_noxref_g ) capacitor \
 c=0.015318f //x=62.575 //y=5.02 //x2=62.94 //y2=6.02
cc_1690 ( N_VDD_c_1710_p N_noxref_19_M122_noxref_g ) capacitor c=0.00672952f \
 //x=63.515 //y=7.4 //x2=63.38 //y2=6.02
cc_1691 ( N_VDD_c_956_n N_noxref_19_M122_noxref_g ) capacitor c=0.00814158f \
 //x=64.38 //y=7.4 //x2=63.38 //y2=6.02
cc_1692 ( N_VDD_M122_noxref_d N_noxref_19_M122_noxref_g ) capacitor \
 c=0.0430452f //x=63.455 //y=5.02 //x2=63.38 //y2=6.02
cc_1693 ( N_VDD_c_950_n N_noxref_19_c_6258_n ) capacitor c=0.00757682f \
 //x=42.92 //y=7.4 //x2=44.305 //y2=4.79
cc_1694 ( N_VDD_M97_noxref_s N_noxref_19_c_6258_n ) capacitor c=0.00444914f \
 //x=43.875 //y=5.02 //x2=44.305 //y2=4.79
cc_1695 ( N_VDD_c_960_p N_noxref_19_M111_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=55.475 //y2=5.02
cc_1696 ( N_VDD_c_1427_p N_noxref_19_M111_noxref_d ) capacitor c=0.0140317f \
 //x=55.975 //y=7.4 //x2=55.475 //y2=5.02
cc_1697 ( N_VDD_c_954_n N_noxref_19_M111_noxref_d ) capacitor c=6.94454e-19 \
 //x=57.72 //y=7.4 //x2=55.475 //y2=5.02
cc_1698 ( N_VDD_M112_noxref_d N_noxref_19_M111_noxref_d ) capacitor \
 c=0.0664752f //x=55.915 //y=5.02 //x2=55.475 //y2=5.02
cc_1699 ( N_VDD_c_960_p N_noxref_19_M113_noxref_d ) capacitor c=0.00285083f \
 //x=73.63 //y=7.4 //x2=56.355 //y2=5.02
cc_1700 ( N_VDD_c_1576_p N_noxref_19_M113_noxref_d ) capacitor c=0.0140984f \
 //x=56.855 //y=7.4 //x2=56.355 //y2=5.02
cc_1701 ( N_VDD_c_954_n N_noxref_19_M113_noxref_d ) capacitor c=0.0120541f \
 //x=57.72 //y=7.4 //x2=56.355 //y2=5.02
cc_1702 ( N_VDD_M111_noxref_s N_noxref_19_M113_noxref_d ) capacitor \
 c=0.00111971f //x=55.045 //y=5.02 //x2=56.355 //y2=5.02
cc_1703 ( N_VDD_M112_noxref_d N_noxref_19_M113_noxref_d ) capacitor \
 c=0.0664752f //x=55.915 //y=5.02 //x2=56.355 //y2=5.02
cc_1704 ( N_VDD_M114_noxref_d N_noxref_19_M113_noxref_d ) capacitor \
 c=0.0664752f //x=56.795 //y=5.02 //x2=56.355 //y2=5.02
cc_1705 ( N_VDD_M115_noxref_s N_noxref_19_M113_noxref_d ) capacitor \
 c=4.54516e-19 //x=58.375 //y=5.02 //x2=56.355 //y2=5.02
cc_1706 ( N_VDD_c_960_p N_noxref_20_c_6592_n ) capacitor c=0.00858137f \
 //x=73.63 //y=7.4 //x2=63.525 //y2=3.7
cc_1707 ( N_VDD_c_960_p N_noxref_20_c_6593_n ) capacitor c=0.00807586f \
 //x=73.63 //y=7.4 //x2=65.005 //y2=3.7
cc_1708 ( N_VDD_c_956_n N_noxref_20_c_6593_n ) capacitor c=0.0109524f \
 //x=64.38 //y=7.4 //x2=65.005 //y2=3.7
cc_1709 ( N_VDD_c_960_p N_noxref_20_c_6595_n ) capacitor c=0.00154061f \
 //x=73.63 //y=7.4 //x2=63.755 //y2=3.7
cc_1710 ( N_VDD_M122_noxref_d N_noxref_20_c_6595_n ) capacitor c=4.05358e-19 \
 //x=63.455 //y=5.02 //x2=63.755 //y2=3.7
cc_1711 ( N_VDD_c_960_p N_noxref_20_c_6597_n ) capacitor c=0.014626f //x=73.63 \
 //y=7.4 //x2=68.705 //y2=4.44
cc_1712 ( N_VDD_c_1734_p N_noxref_20_c_6597_n ) capacitor c=0.00134165f \
 //x=65.965 //y=7.4 //x2=68.705 //y2=4.44
cc_1713 ( N_VDD_c_957_n N_noxref_20_c_6597_n ) capacitor c=0.03415f //x=67.71 \
 //y=7.4 //x2=68.705 //y2=4.44
cc_1714 ( N_VDD_M123_noxref_s N_noxref_20_c_6597_n ) capacitor c=6.29527e-19 \
 //x=65.035 //y=5.025 //x2=68.705 //y2=4.44
cc_1715 ( N_VDD_M126_noxref_d N_noxref_20_c_6597_n ) capacitor c=0.0033086f \
 //x=66.785 //y=5.025 //x2=68.705 //y2=4.44
cc_1716 ( N_VDD_c_960_p N_noxref_20_c_6602_n ) capacitor c=0.00166343f \
 //x=73.63 //y=7.4 //x2=65.235 //y2=4.44
cc_1717 ( N_VDD_c_1739_p N_noxref_20_c_6602_n ) capacitor c=4.53049e-19 \
 //x=65.085 //y=7.4 //x2=65.235 //y2=4.44
cc_1718 ( N_VDD_c_956_n N_noxref_20_c_6602_n ) capacitor c=0.00560881f \
 //x=64.38 //y=7.4 //x2=65.235 //y2=4.44
cc_1719 ( N_VDD_M123_noxref_s N_noxref_20_c_6602_n ) capacitor c=0.00225389f \
 //x=65.035 //y=5.025 //x2=65.235 //y2=4.44
cc_1720 ( N_VDD_c_954_n N_noxref_20_c_6560_n ) capacitor c=0.00111716f \
 //x=57.72 //y=7.4 //x2=59.57 //y2=2.08
cc_1721 ( N_VDD_c_955_n N_noxref_20_c_6560_n ) capacitor c=6.86445e-19 \
 //x=61.05 //y=7.4 //x2=59.57 //y2=2.08
cc_1722 ( N_VDD_c_960_p N_noxref_20_c_6608_n ) capacitor c=0.00459955f \
 //x=73.63 //y=7.4 //x2=63.075 //y2=5.2
cc_1723 ( N_VDD_c_1630_p N_noxref_20_c_6608_n ) capacitor c=4.48705e-19 \
 //x=62.635 //y=7.4 //x2=63.075 //y2=5.2
cc_1724 ( N_VDD_c_1710_p N_noxref_20_c_6608_n ) capacitor c=4.48693e-19 \
 //x=63.515 //y=7.4 //x2=63.075 //y2=5.2
cc_1725 ( N_VDD_M120_noxref_d N_noxref_20_c_6608_n ) capacitor c=0.01269f \
 //x=62.575 //y=5.02 //x2=63.075 //y2=5.2
cc_1726 ( N_VDD_c_955_n N_noxref_20_c_6612_n ) capacitor c=0.00985474f \
 //x=61.05 //y=7.4 //x2=62.365 //y2=5.2
cc_1727 ( N_VDD_M119_noxref_s N_noxref_20_c_6612_n ) capacitor c=0.087833f \
 //x=61.705 //y=5.02 //x2=62.365 //y2=5.2
cc_1728 ( N_VDD_c_960_p N_noxref_20_c_6614_n ) capacitor c=0.00311875f \
 //x=73.63 //y=7.4 //x2=63.555 //y2=5.2
cc_1729 ( N_VDD_c_1710_p N_noxref_20_c_6614_n ) capacitor c=7.21492e-19 \
 //x=63.515 //y=7.4 //x2=63.555 //y2=5.2
cc_1730 ( N_VDD_M122_noxref_d N_noxref_20_c_6614_n ) capacitor c=0.0163364f \
 //x=63.455 //y=5.02 //x2=63.555 //y2=5.2
cc_1731 ( N_VDD_M123_noxref_s N_noxref_20_c_6614_n ) capacitor c=5.34061e-19 \
 //x=65.035 //y=5.025 //x2=63.555 //y2=5.2
cc_1732 ( N_VDD_c_955_n N_noxref_20_c_6563_n ) capacitor c=0.00151618f \
 //x=61.05 //y=7.4 //x2=63.64 //y2=3.7
cc_1733 ( N_VDD_c_956_n N_noxref_20_c_6563_n ) capacitor c=0.0445019f \
 //x=64.38 //y=7.4 //x2=63.64 //y2=3.7
cc_1734 ( N_VDD_c_960_p N_noxref_20_c_6564_n ) capacitor c=0.00142825f \
 //x=73.63 //y=7.4 //x2=65.12 //y2=2.08
cc_1735 ( N_VDD_c_956_n N_noxref_20_c_6564_n ) capacitor c=0.0257873f \
 //x=64.38 //y=7.4 //x2=65.12 //y2=2.08
cc_1736 ( N_VDD_c_957_n N_noxref_20_c_6564_n ) capacitor c=4.17679e-19 \
 //x=67.71 //y=7.4 //x2=65.12 //y2=2.08
cc_1737 ( N_VDD_M123_noxref_s N_noxref_20_c_6564_n ) capacitor c=0.0113998f \
 //x=65.035 //y=5.025 //x2=65.12 //y2=2.08
cc_1738 ( N_VDD_c_957_n N_noxref_20_c_6567_n ) capacitor c=0.0131686f \
 //x=67.71 //y=7.4 //x2=68.82 //y2=2.08
cc_1739 ( N_VDD_c_958_n N_noxref_20_c_6567_n ) capacitor c=0.00133861f \
 //x=71.04 //y=7.4 //x2=68.82 //y2=2.08
cc_1740 ( N_VDD_c_1638_p N_noxref_20_M117_noxref_g ) capacitor c=0.00673971f \
 //x=60.185 //y=7.4 //x2=59.61 //y2=6.02
cc_1741 ( N_VDD_M116_noxref_d N_noxref_20_M117_noxref_g ) capacitor \
 c=0.015318f //x=59.245 //y=5.02 //x2=59.61 //y2=6.02
cc_1742 ( N_VDD_c_1638_p N_noxref_20_M118_noxref_g ) capacitor c=0.00672952f \
 //x=60.185 //y=7.4 //x2=60.05 //y2=6.02
cc_1743 ( N_VDD_c_955_n N_noxref_20_M118_noxref_g ) capacitor c=0.00864163f \
 //x=61.05 //y=7.4 //x2=60.05 //y2=6.02
cc_1744 ( N_VDD_M118_noxref_d N_noxref_20_M118_noxref_g ) capacitor \
 c=0.0430452f //x=60.125 //y=5.02 //x2=60.05 //y2=6.02
cc_1745 ( N_VDD_c_1734_p N_noxref_20_M123_noxref_g ) capacitor c=0.00754867f \
 //x=65.965 //y=7.4 //x2=65.39 //y2=6.025
cc_1746 ( N_VDD_c_956_n N_noxref_20_M123_noxref_g ) capacitor c=0.00684066f \
 //x=64.38 //y=7.4 //x2=65.39 //y2=6.025
cc_1747 ( N_VDD_M123_noxref_s N_noxref_20_M123_noxref_g ) capacitor \
 c=0.0547553f //x=65.035 //y=5.025 //x2=65.39 //y2=6.025
cc_1748 ( N_VDD_c_1734_p N_noxref_20_M124_noxref_g ) capacitor c=0.00678153f \
 //x=65.965 //y=7.4 //x2=65.83 //y2=6.025
cc_1749 ( N_VDD_M124_noxref_d N_noxref_20_M124_noxref_g ) capacitor \
 c=0.015501f //x=65.905 //y=5.025 //x2=65.83 //y2=6.025
cc_1750 ( N_VDD_c_1772_p N_noxref_20_M127_noxref_g ) capacitor c=0.00513227f \
 //x=70.87 //y=7.4 //x2=68.71 //y2=6.025
cc_1751 ( N_VDD_c_957_n N_noxref_20_M127_noxref_g ) capacitor c=0.00316281f \
 //x=67.71 //y=7.4 //x2=68.71 //y2=6.025
cc_1752 ( N_VDD_c_1772_p N_noxref_20_M128_noxref_g ) capacitor c=0.00512552f \
 //x=70.87 //y=7.4 //x2=69.15 //y2=6.025
cc_1753 ( N_VDD_c_956_n N_noxref_20_c_6639_n ) capacitor c=0.0110236f \
 //x=64.38 //y=7.4 //x2=65.465 //y2=4.795
cc_1754 ( N_VDD_M123_noxref_s N_noxref_20_c_6639_n ) capacitor c=0.00628155f \
 //x=65.035 //y=5.025 //x2=65.465 //y2=4.795
cc_1755 ( N_VDD_c_957_n N_noxref_20_c_6641_n ) capacitor c=0.0115029f \
 //x=67.71 //y=7.4 //x2=68.82 //y2=4.705
cc_1756 ( N_VDD_c_960_p N_noxref_20_M119_noxref_d ) capacitor c=0.00278311f \
 //x=73.63 //y=7.4 //x2=62.135 //y2=5.02
cc_1757 ( N_VDD_c_1630_p N_noxref_20_M119_noxref_d ) capacitor c=0.0140526f \
 //x=62.635 //y=7.4 //x2=62.135 //y2=5.02
cc_1758 ( N_VDD_c_956_n N_noxref_20_M119_noxref_d ) capacitor c=6.94454e-19 \
 //x=64.38 //y=7.4 //x2=62.135 //y2=5.02
cc_1759 ( N_VDD_M120_noxref_d N_noxref_20_M119_noxref_d ) capacitor \
 c=0.0664752f //x=62.575 //y=5.02 //x2=62.135 //y2=5.02
cc_1760 ( N_VDD_c_960_p N_noxref_20_M121_noxref_d ) capacitor c=0.00294217f \
 //x=73.63 //y=7.4 //x2=63.015 //y2=5.02
cc_1761 ( N_VDD_c_1710_p N_noxref_20_M121_noxref_d ) capacitor c=0.0138379f \
 //x=63.515 //y=7.4 //x2=63.015 //y2=5.02
cc_1762 ( N_VDD_c_956_n N_noxref_20_M121_noxref_d ) capacitor c=0.0120518f \
 //x=64.38 //y=7.4 //x2=63.015 //y2=5.02
cc_1763 ( N_VDD_M119_noxref_s N_noxref_20_M121_noxref_d ) capacitor \
 c=0.00111971f //x=61.705 //y=5.02 //x2=63.015 //y2=5.02
cc_1764 ( N_VDD_M120_noxref_d N_noxref_20_M121_noxref_d ) capacitor \
 c=0.0664752f //x=62.575 //y=5.02 //x2=63.015 //y2=5.02
cc_1765 ( N_VDD_M122_noxref_d N_noxref_20_M121_noxref_d ) capacitor \
 c=0.0664752f //x=63.455 //y=5.02 //x2=63.015 //y2=5.02
cc_1766 ( N_VDD_M123_noxref_s N_noxref_20_M121_noxref_d ) capacitor \
 c=4.54243e-19 //x=65.035 //y=5.025 //x2=63.015 //y2=5.02
cc_1767 ( N_VDD_c_960_p N_noxref_21_c_6938_n ) capacitor c=0.0151699f \
 //x=73.63 //y=7.4 //x2=72.775 //y2=4.07
cc_1768 ( N_VDD_c_938_n N_noxref_21_c_6938_n ) capacitor c=4.075e-19 //x=73.63 \
 //y=7.4 //x2=72.775 //y2=4.07
cc_1769 ( N_VDD_c_957_n N_noxref_21_c_6938_n ) capacitor c=0.0150456f \
 //x=67.71 //y=7.4 //x2=72.775 //y2=4.07
cc_1770 ( N_VDD_c_958_n N_noxref_21_c_6938_n ) capacitor c=0.0225025f \
 //x=71.04 //y=7.4 //x2=72.775 //y2=4.07
cc_1771 ( N_VDD_c_957_n N_noxref_21_c_6956_n ) capacitor c=5.4458e-19 \
 //x=67.71 //y=7.4 //x2=66.345 //y2=4.07
cc_1772 ( N_VDD_c_948_n N_noxref_21_c_6939_n ) capacitor c=5.3048e-19 \
 //x=36.26 //y=7.4 //x2=38.11 //y2=2.08
cc_1773 ( N_VDD_c_949_n N_noxref_21_c_6939_n ) capacitor c=3.37458e-19 \
 //x=39.59 //y=7.4 //x2=38.11 //y2=2.08
cc_1774 ( N_VDD_c_960_p N_noxref_21_c_6959_n ) capacitor c=0.00453663f \
 //x=73.63 //y=7.4 //x2=41.615 //y2=5.2
cc_1775 ( N_VDD_c_1286_p N_noxref_21_c_6959_n ) capacitor c=4.48391e-19 \
 //x=41.175 //y=7.4 //x2=41.615 //y2=5.2
cc_1776 ( N_VDD_c_1339_p N_noxref_21_c_6959_n ) capacitor c=4.48391e-19 \
 //x=42.055 //y=7.4 //x2=41.615 //y2=5.2
cc_1777 ( N_VDD_M94_noxref_d N_noxref_21_c_6959_n ) capacitor c=0.0124542f \
 //x=41.115 //y=5.02 //x2=41.615 //y2=5.2
cc_1778 ( N_VDD_c_949_n N_noxref_21_c_6963_n ) capacitor c=0.00985474f \
 //x=39.59 //y=7.4 //x2=40.905 //y2=5.2
cc_1779 ( N_VDD_M93_noxref_s N_noxref_21_c_6963_n ) capacitor c=0.087833f \
 //x=40.245 //y=5.02 //x2=40.905 //y2=5.2
cc_1780 ( N_VDD_c_960_p N_noxref_21_c_6965_n ) capacitor c=0.00301575f \
 //x=73.63 //y=7.4 //x2=42.095 //y2=5.2
cc_1781 ( N_VDD_c_1339_p N_noxref_21_c_6965_n ) capacitor c=7.72068e-19 \
 //x=42.055 //y=7.4 //x2=42.095 //y2=5.2
cc_1782 ( N_VDD_M96_noxref_d N_noxref_21_c_6965_n ) capacitor c=0.0158515f \
 //x=41.995 //y=5.02 //x2=42.095 //y2=5.2
cc_1783 ( N_VDD_c_949_n N_noxref_21_c_6942_n ) capacitor c=0.00151618f \
 //x=39.59 //y=7.4 //x2=42.18 //y2=2.22
cc_1784 ( N_VDD_c_950_n N_noxref_21_c_6942_n ) capacitor c=0.0433069f \
 //x=42.92 //y=7.4 //x2=42.18 //y2=2.22
cc_1785 ( N_VDD_c_957_n N_noxref_21_c_6970_n ) capacitor c=0.00491684f \
 //x=67.71 //y=7.4 //x2=66.23 //y2=4.54
cc_1786 ( N_VDD_c_956_n N_noxref_21_c_6944_n ) capacitor c=0.00113585f \
 //x=64.38 //y=7.4 //x2=66.23 //y2=2.08
cc_1787 ( N_VDD_c_957_n N_noxref_21_c_6944_n ) capacitor c=0.0042566f \
 //x=67.71 //y=7.4 //x2=66.23 //y2=2.08
cc_1788 ( N_VDD_c_938_n N_noxref_21_c_6946_n ) capacitor c=6.69172e-19 \
 //x=73.63 //y=7.4 //x2=72.89 //y2=2.08
cc_1789 ( N_VDD_c_958_n N_noxref_21_c_6946_n ) capacitor c=0.00116377f \
 //x=71.04 //y=7.4 //x2=72.89 //y2=2.08
cc_1790 ( N_VDD_c_1275_p N_noxref_21_M91_noxref_g ) capacitor c=0.00673971f \
 //x=38.725 //y=7.4 //x2=38.15 //y2=6.02
cc_1791 ( N_VDD_M90_noxref_d N_noxref_21_M91_noxref_g ) capacitor c=0.015318f \
 //x=37.785 //y=5.02 //x2=38.15 //y2=6.02
cc_1792 ( N_VDD_c_1275_p N_noxref_21_M92_noxref_g ) capacitor c=0.00672952f \
 //x=38.725 //y=7.4 //x2=38.59 //y2=6.02
cc_1793 ( N_VDD_c_949_n N_noxref_21_M92_noxref_g ) capacitor c=0.00864163f \
 //x=39.59 //y=7.4 //x2=38.59 //y2=6.02
cc_1794 ( N_VDD_M92_noxref_d N_noxref_21_M92_noxref_g ) capacitor c=0.0430452f \
 //x=38.665 //y=5.02 //x2=38.59 //y2=6.02
cc_1795 ( N_VDD_c_1817_p N_noxref_21_M125_noxref_g ) capacitor c=0.0067918f \
 //x=66.845 //y=7.4 //x2=66.27 //y2=6.025
cc_1796 ( N_VDD_M124_noxref_d N_noxref_21_M125_noxref_g ) capacitor \
 c=0.015526f //x=65.905 //y=5.025 //x2=66.27 //y2=6.025
cc_1797 ( N_VDD_c_1817_p N_noxref_21_M126_noxref_g ) capacitor c=0.00754867f \
 //x=66.845 //y=7.4 //x2=66.71 //y2=6.025
cc_1798 ( N_VDD_M126_noxref_d N_noxref_21_M126_noxref_g ) capacitor \
 c=0.0537676f //x=66.785 //y=5.025 //x2=66.71 //y2=6.025
cc_1799 ( N_VDD_c_938_n N_noxref_21_M133_noxref_g ) capacitor c=0.00513565f \
 //x=73.63 //y=7.4 //x2=72.93 //y2=6.025
cc_1800 ( N_VDD_c_938_n N_noxref_21_M134_noxref_g ) capacitor c=0.0309137f \
 //x=73.63 //y=7.4 //x2=73.37 //y2=6.025
cc_1801 ( N_VDD_c_957_n N_noxref_21_c_6986_n ) capacitor c=0.00985898f \
 //x=67.71 //y=7.4 //x2=66.635 //y2=4.795
cc_1802 ( N_VDD_c_957_n N_noxref_21_c_6987_n ) capacitor c=2.76772e-19 \
 //x=67.71 //y=7.4 //x2=66.27 //y2=4.705
cc_1803 ( N_VDD_c_960_p N_noxref_21_M93_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=40.675 //y2=5.02
cc_1804 ( N_VDD_c_1286_p N_noxref_21_M93_noxref_d ) capacitor c=0.0140317f \
 //x=41.175 //y=7.4 //x2=40.675 //y2=5.02
cc_1805 ( N_VDD_c_950_n N_noxref_21_M93_noxref_d ) capacitor c=6.94454e-19 \
 //x=42.92 //y=7.4 //x2=40.675 //y2=5.02
cc_1806 ( N_VDD_M94_noxref_d N_noxref_21_M93_noxref_d ) capacitor c=0.0664752f \
 //x=41.115 //y=5.02 //x2=40.675 //y2=5.02
cc_1807 ( N_VDD_c_960_p N_noxref_21_M95_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=41.555 //y2=5.02
cc_1808 ( N_VDD_c_1339_p N_noxref_21_M95_noxref_d ) capacitor c=0.0140317f \
 //x=42.055 //y=7.4 //x2=41.555 //y2=5.02
cc_1809 ( N_VDD_c_950_n N_noxref_21_M95_noxref_d ) capacitor c=0.0120541f \
 //x=42.92 //y=7.4 //x2=41.555 //y2=5.02
cc_1810 ( N_VDD_M93_noxref_s N_noxref_21_M95_noxref_d ) capacitor \
 c=0.00111971f //x=40.245 //y=5.02 //x2=41.555 //y2=5.02
cc_1811 ( N_VDD_M94_noxref_d N_noxref_21_M95_noxref_d ) capacitor c=0.0664752f \
 //x=41.115 //y=5.02 //x2=41.555 //y2=5.02
cc_1812 ( N_VDD_M96_noxref_d N_noxref_21_M95_noxref_d ) capacitor c=0.0664752f \
 //x=41.995 //y=5.02 //x2=41.555 //y2=5.02
cc_1813 ( N_VDD_M97_noxref_s N_noxref_21_M95_noxref_d ) capacitor \
 c=3.73257e-19 //x=43.875 //y=5.02 //x2=41.555 //y2=5.02
cc_1814 ( N_VDD_c_960_p N_noxref_22_c_7406_n ) capacitor c=0.0206457f \
 //x=73.63 //y=7.4 //x2=68.375 //y2=5.21
cc_1815 ( N_VDD_c_1817_p N_noxref_22_c_7406_n ) capacitor c=0.00213763f \
 //x=66.845 //y=7.4 //x2=68.375 //y2=5.21
cc_1816 ( N_VDD_c_1838_p N_noxref_22_c_7406_n ) capacitor c=0.003172f \
 //x=67.54 //y=7.4 //x2=68.375 //y2=5.21
cc_1817 ( N_VDD_c_1772_p N_noxref_22_c_7406_n ) capacitor c=0.00424633f \
 //x=70.87 //y=7.4 //x2=68.375 //y2=5.21
cc_1818 ( N_VDD_c_957_n N_noxref_22_c_7406_n ) capacitor c=0.0430305f \
 //x=67.71 //y=7.4 //x2=68.375 //y2=5.21
cc_1819 ( N_VDD_M126_noxref_d N_noxref_22_c_7406_n ) capacitor c=0.0197937f \
 //x=66.785 //y=5.025 //x2=68.375 //y2=5.21
cc_1820 ( N_VDD_c_960_p N_noxref_22_c_7412_n ) capacitor c=0.00274812f \
 //x=73.63 //y=7.4 //x2=66.605 //y2=5.21
cc_1821 ( N_VDD_c_1817_p N_noxref_22_c_7412_n ) capacitor c=0.00107267f \
 //x=66.845 //y=7.4 //x2=66.605 //y2=5.21
cc_1822 ( N_VDD_c_956_n N_noxref_22_c_7412_n ) capacitor c=2.89592e-19 \
 //x=64.38 //y=7.4 //x2=66.605 //y2=5.21
cc_1823 ( N_VDD_c_957_n N_noxref_22_c_7412_n ) capacitor c=3.35418e-19 \
 //x=67.71 //y=7.4 //x2=66.605 //y2=5.21
cc_1824 ( N_VDD_M126_noxref_d N_noxref_22_c_7412_n ) capacitor c=6.02701e-19 \
 //x=66.785 //y=5.025 //x2=66.605 //y2=5.21
cc_1825 ( N_VDD_c_960_p N_noxref_22_c_7417_n ) capacitor c=0.00453889f \
 //x=73.63 //y=7.4 //x2=66.405 //y2=5.21
cc_1826 ( N_VDD_c_1734_p N_noxref_22_c_7417_n ) capacitor c=4.52207e-19 \
 //x=65.965 //y=7.4 //x2=66.405 //y2=5.21
cc_1827 ( N_VDD_c_1817_p N_noxref_22_c_7417_n ) capacitor c=4.11408e-19 \
 //x=66.845 //y=7.4 //x2=66.405 //y2=5.21
cc_1828 ( N_VDD_M124_noxref_d N_noxref_22_c_7417_n ) capacitor c=0.0127968f \
 //x=65.905 //y=5.025 //x2=66.405 //y2=5.21
cc_1829 ( N_VDD_c_956_n N_noxref_22_c_7421_n ) capacitor c=0.00914165f \
 //x=64.38 //y=7.4 //x2=65.695 //y2=5.21
cc_1830 ( N_VDD_M123_noxref_s N_noxref_22_c_7421_n ) capacitor c=0.0872987f \
 //x=65.035 //y=5.025 //x2=65.695 //y2=5.21
cc_1831 ( N_VDD_c_956_n N_noxref_22_c_7423_n ) capacitor c=6.3991e-19 \
 //x=64.38 //y=7.4 //x2=66.49 //y2=5.295
cc_1832 ( N_VDD_c_957_n N_noxref_22_c_7423_n ) capacitor c=0.00985441f \
 //x=67.71 //y=7.4 //x2=66.49 //y2=5.295
cc_1833 ( N_VDD_M126_noxref_d N_noxref_22_c_7423_n ) capacitor c=0.0873334f \
 //x=66.785 //y=5.025 //x2=66.49 //y2=5.295
cc_1834 ( N_VDD_c_957_n N_noxref_22_c_7426_n ) capacitor c=0.0674112f \
 //x=67.71 //y=7.4 //x2=68.49 //y2=5.21
cc_1835 ( N_VDD_M126_noxref_d N_noxref_22_c_7426_n ) capacitor c=0.00235009f \
 //x=66.785 //y=5.025 //x2=68.49 //y2=5.21
cc_1836 ( N_VDD_c_960_p N_noxref_22_c_7428_n ) capacitor c=0.0296174f \
 //x=73.63 //y=7.4 //x2=68.575 //y2=6.91
cc_1837 ( N_VDD_c_1772_p N_noxref_22_c_7428_n ) capacitor c=0.109938f \
 //x=70.87 //y=7.4 //x2=68.575 //y2=6.91
cc_1838 ( N_VDD_c_960_p N_noxref_22_M123_noxref_d ) capacitor c=0.00291898f \
 //x=73.63 //y=7.4 //x2=65.465 //y2=5.025
cc_1839 ( N_VDD_c_1734_p N_noxref_22_M123_noxref_d ) capacitor c=0.0137097f \
 //x=65.965 //y=7.4 //x2=65.465 //y2=5.025
cc_1840 ( N_VDD_M124_noxref_d N_noxref_22_M123_noxref_d ) capacitor \
 c=0.067695f //x=65.905 //y=5.025 //x2=65.465 //y2=5.025
cc_1841 ( N_VDD_M126_noxref_d N_noxref_22_M123_noxref_d ) capacitor \
 c=0.00105738f //x=66.785 //y=5.025 //x2=65.465 //y2=5.025
cc_1842 ( N_VDD_c_960_p N_noxref_22_M125_noxref_d ) capacitor c=0.00241371f \
 //x=73.63 //y=7.4 //x2=66.345 //y2=5.025
cc_1843 ( N_VDD_c_1817_p N_noxref_22_M125_noxref_d ) capacitor c=0.01268f \
 //x=66.845 //y=7.4 //x2=66.345 //y2=5.025
cc_1844 ( N_VDD_M123_noxref_s N_noxref_22_M125_noxref_d ) capacitor \
 c=0.00103189f //x=65.035 //y=5.025 //x2=66.345 //y2=5.025
cc_1845 ( N_VDD_M124_noxref_d N_noxref_22_M125_noxref_d ) capacitor \
 c=0.0653408f //x=65.905 //y=5.025 //x2=66.345 //y2=5.025
cc_1846 ( N_VDD_c_957_n N_noxref_22_M128_noxref_d ) capacitor c=8.96067e-19 \
 //x=67.71 //y=7.4 //x2=69.225 //y2=5.025
cc_1847 ( N_VDD_c_958_n N_noxref_22_M128_noxref_d ) capacitor c=8.88629e-19 \
 //x=71.04 //y=7.4 //x2=69.225 //y2=5.025
cc_1848 ( N_VDD_c_958_n N_noxref_22_M130_noxref_d ) capacitor c=0.0575594f \
 //x=71.04 //y=7.4 //x2=70.105 //y2=5.025
cc_1849 ( N_VDD_c_944_n N_noxref_23_c_7498_n ) capacitor c=0.00315988f \
 //x=21.46 //y=7.4 //x2=70.185 //y2=2.96
cc_1850 ( N_VDD_c_950_n N_noxref_23_c_7498_n ) capacitor c=0.00315988f \
 //x=42.92 //y=7.4 //x2=70.185 //y2=2.96
cc_1851 ( N_VDD_c_942_n N_noxref_23_c_7515_n ) capacitor c=5.6016e-19 //x=14.8 \
 //y=7.4 //x2=16.65 //y2=2.08
cc_1852 ( N_VDD_c_943_n N_noxref_23_c_7515_n ) capacitor c=3.59368e-19 \
 //x=18.13 //y=7.4 //x2=16.65 //y2=2.08
cc_1853 ( N_VDD_c_960_p N_noxref_23_c_7540_n ) capacitor c=0.00453663f \
 //x=73.63 //y=7.4 //x2=20.155 //y2=5.2
cc_1854 ( N_VDD_c_1085_p N_noxref_23_c_7540_n ) capacitor c=4.48391e-19 \
 //x=19.715 //y=7.4 //x2=20.155 //y2=5.2
cc_1855 ( N_VDD_c_1142_p N_noxref_23_c_7540_n ) capacitor c=4.48391e-19 \
 //x=20.595 //y=7.4 //x2=20.155 //y2=5.2
cc_1856 ( N_VDD_M68_noxref_d N_noxref_23_c_7540_n ) capacitor c=0.0124542f \
 //x=19.655 //y=5.02 //x2=20.155 //y2=5.2
cc_1857 ( N_VDD_c_943_n N_noxref_23_c_7544_n ) capacitor c=0.00985474f \
 //x=18.13 //y=7.4 //x2=19.445 //y2=5.2
cc_1858 ( N_VDD_M67_noxref_s N_noxref_23_c_7544_n ) capacitor c=0.087833f \
 //x=18.785 //y=5.02 //x2=19.445 //y2=5.2
cc_1859 ( N_VDD_c_960_p N_noxref_23_c_7546_n ) capacitor c=0.00301575f \
 //x=73.63 //y=7.4 //x2=20.635 //y2=5.2
cc_1860 ( N_VDD_c_1142_p N_noxref_23_c_7546_n ) capacitor c=7.72068e-19 \
 //x=20.595 //y=7.4 //x2=20.635 //y2=5.2
cc_1861 ( N_VDD_M70_noxref_d N_noxref_23_c_7546_n ) capacitor c=0.0158515f \
 //x=20.535 //y=5.02 //x2=20.635 //y2=5.2
cc_1862 ( N_VDD_c_943_n N_noxref_23_c_7518_n ) capacitor c=0.00151618f \
 //x=18.13 //y=7.4 //x2=20.72 //y2=2.96
cc_1863 ( N_VDD_c_944_n N_noxref_23_c_7518_n ) capacitor c=0.0433069f \
 //x=21.46 //y=7.4 //x2=20.72 //y2=2.96
cc_1864 ( N_VDD_c_957_n N_noxref_23_c_7519_n ) capacitor c=7.57423e-19 \
 //x=67.71 //y=7.4 //x2=70.3 //y2=2.08
cc_1865 ( N_VDD_c_958_n N_noxref_23_c_7519_n ) capacitor c=0.0263215f \
 //x=71.04 //y=7.4 //x2=70.3 //y2=2.08
cc_1866 ( N_VDD_c_958_n N_noxref_23_c_7521_n ) capacitor c=0.0263871f \
 //x=71.04 //y=7.4 //x2=71.78 //y2=2.08
cc_1867 ( N_VDD_c_1074_p N_noxref_23_M65_noxref_g ) capacitor c=0.00673971f \
 //x=17.265 //y=7.4 //x2=16.69 //y2=6.02
cc_1868 ( N_VDD_M64_noxref_d N_noxref_23_M65_noxref_g ) capacitor c=0.015318f \
 //x=16.325 //y=5.02 //x2=16.69 //y2=6.02
cc_1869 ( N_VDD_c_1074_p N_noxref_23_M66_noxref_g ) capacitor c=0.00672952f \
 //x=17.265 //y=7.4 //x2=17.13 //y2=6.02
cc_1870 ( N_VDD_c_943_n N_noxref_23_M66_noxref_g ) capacitor c=0.00864163f \
 //x=18.13 //y=7.4 //x2=17.13 //y2=6.02
cc_1871 ( N_VDD_M66_noxref_d N_noxref_23_M66_noxref_g ) capacitor c=0.0430452f \
 //x=17.205 //y=5.02 //x2=17.13 //y2=6.02
cc_1872 ( N_VDD_c_1772_p N_noxref_23_M129_noxref_g ) capacitor c=0.00512552f \
 //x=70.87 //y=7.4 //x2=69.59 //y2=6.025
cc_1873 ( N_VDD_c_1772_p N_noxref_23_M130_noxref_g ) capacitor c=0.00512552f \
 //x=70.87 //y=7.4 //x2=70.03 //y2=6.025
cc_1874 ( N_VDD_c_958_n N_noxref_23_M130_noxref_g ) capacitor c=0.010355f \
 //x=71.04 //y=7.4 //x2=70.03 //y2=6.025
cc_1875 ( N_VDD_c_938_n N_noxref_23_M131_noxref_g ) capacitor c=0.00512552f \
 //x=73.63 //y=7.4 //x2=72.05 //y2=6.025
cc_1876 ( N_VDD_c_958_n N_noxref_23_M131_noxref_g ) capacitor c=0.00767856f \
 //x=71.04 //y=7.4 //x2=72.05 //y2=6.025
cc_1877 ( N_VDD_c_938_n N_noxref_23_M132_noxref_g ) capacitor c=0.00512552f \
 //x=73.63 //y=7.4 //x2=72.49 //y2=6.025
cc_1878 ( N_VDD_c_958_n N_noxref_23_c_7565_n ) capacitor c=0.00803198f \
 //x=71.04 //y=7.4 //x2=70.03 //y2=4.87
cc_1879 ( N_VDD_c_958_n N_noxref_23_c_7566_n ) capacitor c=0.00803198f \
 //x=71.04 //y=7.4 //x2=72.125 //y2=4.795
cc_1880 ( N_VDD_c_960_p N_noxref_23_M67_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=19.215 //y2=5.02
cc_1881 ( N_VDD_c_1085_p N_noxref_23_M67_noxref_d ) capacitor c=0.0140317f \
 //x=19.715 //y=7.4 //x2=19.215 //y2=5.02
cc_1882 ( N_VDD_c_944_n N_noxref_23_M67_noxref_d ) capacitor c=6.94454e-19 \
 //x=21.46 //y=7.4 //x2=19.215 //y2=5.02
cc_1883 ( N_VDD_M68_noxref_d N_noxref_23_M67_noxref_d ) capacitor c=0.0664752f \
 //x=19.655 //y=5.02 //x2=19.215 //y2=5.02
cc_1884 ( N_VDD_c_960_p N_noxref_23_M69_noxref_d ) capacitor c=0.00275225f \
 //x=73.63 //y=7.4 //x2=20.095 //y2=5.02
cc_1885 ( N_VDD_c_1142_p N_noxref_23_M69_noxref_d ) capacitor c=0.0140317f \
 //x=20.595 //y=7.4 //x2=20.095 //y2=5.02
cc_1886 ( N_VDD_c_944_n N_noxref_23_M69_noxref_d ) capacitor c=0.0120541f \
 //x=21.46 //y=7.4 //x2=20.095 //y2=5.02
cc_1887 ( N_VDD_M67_noxref_s N_noxref_23_M69_noxref_d ) capacitor \
 c=0.00111971f //x=18.785 //y=5.02 //x2=20.095 //y2=5.02
cc_1888 ( N_VDD_M68_noxref_d N_noxref_23_M69_noxref_d ) capacitor c=0.0664752f \
 //x=19.655 //y=5.02 //x2=20.095 //y2=5.02
cc_1889 ( N_VDD_M70_noxref_d N_noxref_23_M69_noxref_d ) capacitor c=0.0664752f \
 //x=20.535 //y=5.02 //x2=20.095 //y2=5.02
cc_1890 ( N_VDD_M71_noxref_s N_noxref_23_M69_noxref_d ) capacitor \
 c=3.73257e-19 //x=22.415 //y=5.02 //x2=20.095 //y2=5.02
cc_1891 ( N_VDD_c_960_p N_noxref_24_c_7956_n ) capacitor c=0.0212729f \
 //x=73.63 //y=7.4 //x2=71.715 //y2=5.21
cc_1892 ( N_VDD_c_1772_p N_noxref_24_c_7956_n ) capacitor c=0.00386143f \
 //x=70.87 //y=7.4 //x2=71.715 //y2=5.21
cc_1893 ( N_VDD_c_938_n N_noxref_24_c_7956_n ) capacitor c=0.00403412f \
 //x=73.63 //y=7.4 //x2=71.715 //y2=5.21
cc_1894 ( N_VDD_c_958_n N_noxref_24_c_7956_n ) capacitor c=0.0473381f \
 //x=71.04 //y=7.4 //x2=71.715 //y2=5.21
cc_1895 ( N_VDD_c_960_p N_noxref_24_c_7960_n ) capacitor c=0.00264311f \
 //x=73.63 //y=7.4 //x2=69.925 //y2=5.21
cc_1896 ( N_VDD_c_958_n N_noxref_24_c_7960_n ) capacitor c=6.67754e-19 \
 //x=71.04 //y=7.4 //x2=69.925 //y2=5.21
cc_1897 ( N_VDD_c_957_n N_noxref_24_c_7962_n ) capacitor c=0.00662411f \
 //x=67.71 //y=7.4 //x2=69.015 //y2=5.21
cc_1898 ( N_VDD_c_958_n N_noxref_24_c_7963_n ) capacitor c=0.00999961f \
 //x=71.04 //y=7.4 //x2=69.81 //y2=5.295
cc_1899 ( N_VDD_c_938_n N_noxref_24_c_7964_n ) capacitor c=6.48751e-19 \
 //x=73.63 //y=7.4 //x2=71.83 //y2=5.21
cc_1900 ( N_VDD_c_958_n N_noxref_24_c_7964_n ) capacitor c=0.0664301f \
 //x=71.04 //y=7.4 //x2=71.83 //y2=5.21
cc_1901 ( N_VDD_c_960_p N_noxref_24_c_7966_n ) capacitor c=0.043423f //x=73.63 \
 //y=7.4 //x2=71.915 //y2=6.91
cc_1902 ( N_VDD_c_938_n N_noxref_24_c_7966_n ) capacitor c=0.108124f //x=73.63 \
 //y=7.4 //x2=71.915 //y2=6.91
cc_1903 ( N_VDD_c_938_n N_noxref_24_M132_noxref_d ) capacitor c=8.96067e-19 \
 //x=73.63 //y=7.4 //x2=72.565 //y2=5.025
cc_1904 ( N_VDD_c_958_n N_noxref_24_M132_noxref_d ) capacitor c=8.88629e-19 \
 //x=71.04 //y=7.4 //x2=72.565 //y2=5.025
cc_1905 ( N_VDD_c_938_n N_noxref_24_M134_noxref_d ) capacitor c=0.0529764f \
 //x=73.63 //y=7.4 //x2=73.445 //y2=5.025
cc_1906 ( N_VDD_c_938_n QN ) capacitor c=0.0470629f //x=73.63 //y=7.4 \
 //x2=73.63 //y2=2.22
cc_1907 ( N_VDD_c_958_n QN ) capacitor c=0.00147633f //x=71.04 //y=7.4 \
 //x2=73.63 //y2=2.22
cc_1908 ( N_VDD_c_958_n N_QN_c_8074_n ) capacitor c=0.00660621f //x=71.04 \
 //y=7.4 //x2=72.355 //y2=5.21
cc_1909 ( N_VDD_c_960_p N_QN_c_8075_n ) capacitor c=0.00240012f //x=73.63 \
 //y=7.4 //x2=73.545 //y2=5.21
cc_1910 ( N_VDD_c_938_n N_QN_c_8075_n ) capacitor c=0.00136974f //x=73.63 \
 //y=7.4 //x2=73.545 //y2=5.21
cc_1911 ( N_VDD_c_938_n N_QN_M131_noxref_d ) capacitor c=6.67979e-19 //x=73.63 \
 //y=7.4 //x2=72.125 //y2=5.025
cc_1912 ( N_VDD_c_938_n N_QN_M133_noxref_d ) capacitor c=0.0099096f //x=73.63 \
 //y=7.4 //x2=73.005 //y2=5.025
cc_1913 ( N_noxref_3_c_1940_n N_noxref_4_c_2215_n ) capacitor c=0.011463f \
 //x=9.135 //y=3.33 //x2=10.845 //y2=3.33
cc_1914 ( N_noxref_3_M56_noxref_g N_noxref_4_c_2184_n ) capacitor c=0.0169521f \
 //x=9.59 //y=6.02 //x2=10.165 //y2=5.2
cc_1915 ( N_noxref_3_c_1944_n N_noxref_4_c_2188_n ) capacitor c=0.00539951f \
 //x=9.25 //y=2.08 //x2=9.455 //y2=5.2
cc_1916 ( N_noxref_3_M55_noxref_g N_noxref_4_c_2188_n ) capacitor c=0.0177326f \
 //x=9.15 //y=6.02 //x2=9.455 //y2=5.2
cc_1917 ( N_noxref_3_c_1982_n N_noxref_4_c_2188_n ) capacitor c=0.00581252f \
 //x=9.25 //y=4.7 //x2=9.455 //y2=5.2
cc_1918 ( N_noxref_3_c_1943_n N_noxref_4_c_2169_n ) capacitor c=3.49822e-19 \
 //x=7.4 //y=3.33 //x2=10.73 //y2=3.33
cc_1919 ( N_noxref_3_c_1944_n N_noxref_4_c_2169_n ) capacitor c=0.00297939f \
 //x=9.25 //y=2.08 //x2=10.73 //y2=3.33
cc_1920 ( N_noxref_3_M56_noxref_g N_noxref_4_M55_noxref_d ) capacitor \
 c=0.0173476f //x=9.59 //y=6.02 //x2=9.225 //y2=5.02
cc_1921 ( N_noxref_3_c_1935_n N_noxref_5_c_2388_n ) capacitor c=0.146341f \
 //x=7.285 //y=3.33 //x2=5.805 //y2=3.7
cc_1922 ( N_noxref_3_c_1935_n N_noxref_5_c_2389_n ) capacitor c=0.0294746f \
 //x=7.285 //y=3.33 //x2=4.185 //y2=3.7
cc_1923 ( N_noxref_3_c_1941_n N_noxref_5_c_2389_n ) capacitor c=0.00687545f \
 //x=3.33 //y=2.08 //x2=4.185 //y2=3.7
cc_1924 ( N_noxref_3_c_1935_n N_noxref_5_c_2317_n ) capacitor c=0.108749f \
 //x=7.285 //y=3.33 //x2=15.795 //y2=3.7
cc_1925 ( N_noxref_3_c_1940_n N_noxref_5_c_2317_n ) capacitor c=0.175696f \
 //x=9.135 //y=3.33 //x2=15.795 //y2=3.7
cc_1926 ( N_noxref_3_c_2007_p N_noxref_5_c_2317_n ) capacitor c=0.0267668f \
 //x=7.515 //y=3.33 //x2=15.795 //y2=3.7
cc_1927 ( N_noxref_3_c_1943_n N_noxref_5_c_2317_n ) capacitor c=0.0206034f \
 //x=7.4 //y=3.33 //x2=15.795 //y2=3.7
cc_1928 ( N_noxref_3_c_1944_n N_noxref_5_c_2317_n ) capacitor c=0.0205831f \
 //x=9.25 //y=2.08 //x2=15.795 //y2=3.7
cc_1929 ( N_noxref_3_c_1935_n N_noxref_5_c_2396_n ) capacitor c=0.0266674f \
 //x=7.285 //y=3.33 //x2=6.035 //y2=3.7
cc_1930 ( N_noxref_3_M49_noxref_g N_noxref_5_c_2348_n ) capacitor c=0.01736f \
 //x=3.07 //y=6.02 //x2=3.205 //y2=5.155
cc_1931 ( N_noxref_3_M50_noxref_g N_noxref_5_c_2352_n ) capacitor c=0.0194981f \
 //x=3.51 //y=6.02 //x2=3.985 //y2=5.155
cc_1932 ( N_noxref_3_c_2013_p N_noxref_5_c_2352_n ) capacitor c=0.00201851f \
 //x=3.33 //y=4.7 //x2=3.985 //y2=5.155
cc_1933 ( N_noxref_3_c_2014_p N_noxref_5_c_2318_n ) capacitor c=0.00359704f \
 //x=3.695 //y=1.415 //x2=3.985 //y2=1.665
cc_1934 ( N_noxref_3_c_2015_p N_noxref_5_c_2318_n ) capacitor c=0.00457401f \
 //x=3.85 //y=1.26 //x2=3.985 //y2=1.665
cc_1935 ( N_noxref_3_c_1935_n N_noxref_5_c_2402_n ) capacitor c=0.00628992f \
 //x=7.285 //y=3.33 //x2=3.67 //y2=1.665
cc_1936 ( N_noxref_3_c_1935_n N_noxref_5_c_2356_n ) capacitor c=0.0260398f \
 //x=7.285 //y=3.33 //x2=4.07 //y2=3.7
cc_1937 ( N_noxref_3_c_1939_n N_noxref_5_c_2356_n ) capacitor c=0.00117715f \
 //x=3.445 //y=3.33 //x2=4.07 //y2=3.7
cc_1938 ( N_noxref_3_c_1941_n N_noxref_5_c_2356_n ) capacitor c=0.0828498f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_1939 ( N_noxref_3_c_1943_n N_noxref_5_c_2356_n ) capacitor c=3.52729e-19 \
 //x=7.4 //y=3.33 //x2=4.07 //y2=3.7
cc_1940 ( N_noxref_3_c_2021_p N_noxref_5_c_2356_n ) capacitor c=0.00877984f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_1941 ( N_noxref_3_c_2022_p N_noxref_5_c_2356_n ) capacitor c=0.00283672f \
 //x=3.33 //y=1.915 //x2=4.07 //y2=3.7
cc_1942 ( N_noxref_3_c_2013_p N_noxref_5_c_2356_n ) capacitor c=0.013693f \
 //x=3.33 //y=4.7 //x2=4.07 //y2=3.7
cc_1943 ( N_noxref_3_c_1935_n N_noxref_5_c_2319_n ) capacitor c=0.0257693f \
 //x=7.285 //y=3.33 //x2=5.92 //y2=2.08
cc_1944 ( N_noxref_3_c_1941_n N_noxref_5_c_2319_n ) capacitor c=9.66956e-19 \
 //x=3.33 //y=2.08 //x2=5.92 //y2=2.08
cc_1945 ( N_noxref_3_c_1963_n N_noxref_5_c_2319_n ) capacitor c=0.00521572f \
 //x=6.125 //y=5.2 //x2=5.92 //y2=2.08
cc_1946 ( N_noxref_3_c_1943_n N_noxref_5_c_2319_n ) capacitor c=0.00336482f \
 //x=7.4 //y=3.33 //x2=5.92 //y2=2.08
cc_1947 ( N_noxref_3_c_1941_n N_noxref_5_c_2414_n ) capacitor c=0.0171303f \
 //x=3.33 //y=2.08 //x2=3.29 //y2=5.155
cc_1948 ( N_noxref_3_c_2013_p N_noxref_5_c_2414_n ) capacitor c=0.00475601f \
 //x=3.33 //y=4.7 //x2=3.29 //y2=5.155
cc_1949 ( N_noxref_3_c_1963_n N_noxref_5_M51_noxref_g ) capacitor c=0.0177326f \
 //x=6.125 //y=5.2 //x2=5.82 //y2=6.02
cc_1950 ( N_noxref_3_c_1959_n N_noxref_5_M52_noxref_g ) capacitor c=0.0169521f \
 //x=6.835 //y=5.2 //x2=6.26 //y2=6.02
cc_1951 ( N_noxref_3_M51_noxref_d N_noxref_5_M52_noxref_g ) capacitor \
 c=0.0173476f //x=5.895 //y=5.02 //x2=6.26 //y2=6.02
cc_1952 ( N_noxref_3_c_1963_n N_noxref_5_c_2371_n ) capacitor c=0.00581252f \
 //x=6.125 //y=5.2 //x2=5.92 //y2=4.7
cc_1953 ( N_noxref_3_c_2034_p N_noxref_5_M2_noxref_d ) capacitor c=0.00217566f \
 //x=3.32 //y=0.915 //x2=3.395 //y2=0.915
cc_1954 ( N_noxref_3_c_2035_p N_noxref_5_M2_noxref_d ) capacitor c=0.0034598f \
 //x=3.32 //y=1.26 //x2=3.395 //y2=0.915
cc_1955 ( N_noxref_3_c_2036_p N_noxref_5_M2_noxref_d ) capacitor c=0.00544291f \
 //x=3.32 //y=1.57 //x2=3.395 //y2=0.915
cc_1956 ( N_noxref_3_c_2037_p N_noxref_5_M2_noxref_d ) capacitor c=0.00241102f \
 //x=3.695 //y=0.76 //x2=3.395 //y2=0.915
cc_1957 ( N_noxref_3_c_2014_p N_noxref_5_M2_noxref_d ) capacitor c=0.0140297f \
 //x=3.695 //y=1.415 //x2=3.395 //y2=0.915
cc_1958 ( N_noxref_3_c_2039_p N_noxref_5_M2_noxref_d ) capacitor c=0.00219619f \
 //x=3.85 //y=0.915 //x2=3.395 //y2=0.915
cc_1959 ( N_noxref_3_c_2015_p N_noxref_5_M2_noxref_d ) capacitor c=0.00603828f \
 //x=3.85 //y=1.26 //x2=3.395 //y2=0.915
cc_1960 ( N_noxref_3_c_2022_p N_noxref_5_M2_noxref_d ) capacitor c=0.00661782f \
 //x=3.33 //y=1.915 //x2=3.395 //y2=0.915
cc_1961 ( N_noxref_3_M49_noxref_g N_noxref_5_M49_noxref_d ) capacitor \
 c=0.0180032f //x=3.07 //y=6.02 //x2=3.145 //y2=5.02
cc_1962 ( N_noxref_3_M50_noxref_g N_noxref_5_M49_noxref_d ) capacitor \
 c=0.0194246f //x=3.51 //y=6.02 //x2=3.145 //y2=5.02
cc_1963 ( N_noxref_3_c_1935_n N_noxref_7_c_2715_n ) capacitor c=0.0428508f \
 //x=7.285 //y=3.33 //x2=9.875 //y2=4.07
cc_1964 ( N_noxref_3_c_1939_n N_noxref_7_c_2715_n ) capacitor c=0.0135672f \
 //x=3.445 //y=3.33 //x2=9.875 //y2=4.07
cc_1965 ( N_noxref_3_c_1940_n N_noxref_7_c_2715_n ) capacitor c=0.0110241f \
 //x=9.135 //y=3.33 //x2=9.875 //y2=4.07
cc_1966 ( N_noxref_3_c_2007_p N_noxref_7_c_2715_n ) capacitor c=5.70661e-19 \
 //x=7.515 //y=3.33 //x2=9.875 //y2=4.07
cc_1967 ( N_noxref_3_c_1941_n N_noxref_7_c_2715_n ) capacitor c=0.0206302f \
 //x=3.33 //y=2.08 //x2=9.875 //y2=4.07
cc_1968 ( N_noxref_3_c_1943_n N_noxref_7_c_2715_n ) capacitor c=0.0181936f \
 //x=7.4 //y=3.33 //x2=9.875 //y2=4.07
cc_1969 ( N_noxref_3_c_1944_n N_noxref_7_c_2715_n ) capacitor c=0.0184765f \
 //x=9.25 //y=2.08 //x2=9.875 //y2=4.07
cc_1970 ( N_noxref_3_c_1944_n N_noxref_7_c_2801_n ) capacitor c=0.00179385f \
 //x=9.25 //y=2.08 //x2=10.105 //y2=4.07
cc_1971 ( N_noxref_3_c_1941_n N_noxref_7_c_2717_n ) capacitor c=0.00175117f \
 //x=3.33 //y=2.08 //x2=1.11 //y2=2.08
cc_1972 ( N_noxref_3_c_1944_n N_noxref_7_c_2803_n ) capacitor c=0.00400249f \
 //x=9.25 //y=2.08 //x2=9.99 //y2=4.535
cc_1973 ( N_noxref_3_c_1982_n N_noxref_7_c_2803_n ) capacitor c=0.00417994f \
 //x=9.25 //y=4.7 //x2=9.99 //y2=4.535
cc_1974 ( N_noxref_3_c_1940_n N_noxref_7_c_2718_n ) capacitor c=0.00318578f \
 //x=9.135 //y=3.33 //x2=9.99 //y2=2.08
cc_1975 ( N_noxref_3_c_1943_n N_noxref_7_c_2718_n ) capacitor c=9.69022e-19 \
 //x=7.4 //y=3.33 //x2=9.99 //y2=2.08
cc_1976 ( N_noxref_3_c_1944_n N_noxref_7_c_2718_n ) capacitor c=0.0768945f \
 //x=9.25 //y=2.08 //x2=9.99 //y2=2.08
cc_1977 ( N_noxref_3_c_1949_n N_noxref_7_c_2718_n ) capacitor c=0.00308814f \
 //x=9.055 //y=1.915 //x2=9.99 //y2=2.08
cc_1978 ( N_noxref_3_M55_noxref_g N_noxref_7_M57_noxref_g ) capacitor \
 c=0.0104611f //x=9.15 //y=6.02 //x2=10.03 //y2=6.02
cc_1979 ( N_noxref_3_M56_noxref_g N_noxref_7_M57_noxref_g ) capacitor \
 c=0.106811f //x=9.59 //y=6.02 //x2=10.03 //y2=6.02
cc_1980 ( N_noxref_3_M56_noxref_g N_noxref_7_M58_noxref_g ) capacitor \
 c=0.0100341f //x=9.59 //y=6.02 //x2=10.47 //y2=6.02
cc_1981 ( N_noxref_3_c_1945_n N_noxref_7_c_2812_n ) capacitor c=4.86506e-19 \
 //x=9.055 //y=0.865 //x2=10.025 //y2=0.905
cc_1982 ( N_noxref_3_c_1947_n N_noxref_7_c_2812_n ) capacitor c=0.00152104f \
 //x=9.055 //y=1.21 //x2=10.025 //y2=0.905
cc_1983 ( N_noxref_3_c_1952_n N_noxref_7_c_2812_n ) capacitor c=0.0151475f \
 //x=9.585 //y=0.865 //x2=10.025 //y2=0.905
cc_1984 ( N_noxref_3_c_1948_n N_noxref_7_c_2815_n ) capacitor c=0.00109982f \
 //x=9.055 //y=1.52 //x2=10.025 //y2=1.25
cc_1985 ( N_noxref_3_c_1954_n N_noxref_7_c_2815_n ) capacitor c=0.0111064f \
 //x=9.585 //y=1.21 //x2=10.025 //y2=1.25
cc_1986 ( N_noxref_3_c_1948_n N_noxref_7_c_2817_n ) capacitor c=9.57794e-19 \
 //x=9.055 //y=1.52 //x2=10.025 //y2=1.56
cc_1987 ( N_noxref_3_c_1949_n N_noxref_7_c_2817_n ) capacitor c=0.00662747f \
 //x=9.055 //y=1.915 //x2=10.025 //y2=1.56
cc_1988 ( N_noxref_3_c_1954_n N_noxref_7_c_2817_n ) capacitor c=0.00862358f \
 //x=9.585 //y=1.21 //x2=10.025 //y2=1.56
cc_1989 ( N_noxref_3_c_1952_n N_noxref_7_c_2820_n ) capacitor c=0.00124821f \
 //x=9.585 //y=0.865 //x2=10.555 //y2=0.905
cc_1990 ( N_noxref_3_c_1954_n N_noxref_7_c_2821_n ) capacitor c=0.00200715f \
 //x=9.585 //y=1.21 //x2=10.555 //y2=1.25
cc_1991 ( N_noxref_3_c_1944_n N_noxref_7_c_2822_n ) capacitor c=0.00307062f \
 //x=9.25 //y=2.08 //x2=9.99 //y2=2.08
cc_1992 ( N_noxref_3_c_1949_n N_noxref_7_c_2822_n ) capacitor c=0.0179092f \
 //x=9.055 //y=1.915 //x2=9.99 //y2=2.08
cc_1993 ( N_noxref_3_c_1944_n N_noxref_7_c_2824_n ) capacitor c=0.00344981f \
 //x=9.25 //y=2.08 //x2=10.02 //y2=4.7
cc_1994 ( N_noxref_3_c_1982_n N_noxref_7_c_2824_n ) capacitor c=0.0293367f \
 //x=9.25 //y=4.7 //x2=10.02 //y2=4.7
cc_1995 ( N_noxref_3_c_1935_n N_D_c_4217_n ) capacitor c=0.0214765f //x=7.285 \
 //y=3.33 //x2=28.005 //y2=2.59
cc_1996 ( N_noxref_3_c_1940_n N_D_c_4217_n ) capacitor c=0.083897f //x=9.135 \
 //y=3.33 //x2=28.005 //y2=2.59
cc_1997 ( N_noxref_3_c_2007_p N_D_c_4217_n ) capacitor c=0.0120757f //x=7.515 \
 //y=3.33 //x2=28.005 //y2=2.59
cc_1998 ( N_noxref_3_c_2079_p N_D_c_4217_n ) capacitor c=0.0102711f //x=7.045 \
 //y=1.655 //x2=28.005 //y2=2.59
cc_1999 ( N_noxref_3_c_1943_n N_D_c_4217_n ) capacitor c=0.0237178f //x=7.4 \
 //y=3.33 //x2=28.005 //y2=2.59
cc_2000 ( N_noxref_3_c_1944_n N_D_c_4217_n ) capacitor c=0.0239823f //x=9.25 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2001 ( N_noxref_3_c_1949_n N_D_c_4217_n ) capacitor c=0.00424331f //x=9.055 \
 //y=1.915 //x2=28.005 //y2=2.59
cc_2002 ( N_noxref_3_c_1935_n N_D_c_4236_n ) capacitor c=0.0132679f //x=7.285 \
 //y=3.33 //x2=6.775 //y2=2.59
cc_2003 ( N_noxref_3_c_1943_n N_D_c_4236_n ) capacitor c=0.00179385f //x=7.4 \
 //y=3.33 //x2=6.775 //y2=2.59
cc_2004 ( N_noxref_3_c_1959_n N_D_c_4289_n ) capacitor c=0.0127676f //x=6.835 \
 //y=5.2 //x2=6.66 //y2=4.535
cc_2005 ( N_noxref_3_c_1943_n N_D_c_4289_n ) capacitor c=0.0101284f //x=7.4 \
 //y=3.33 //x2=6.66 //y2=4.535
cc_2006 ( N_noxref_3_c_1935_n N_D_c_4253_n ) capacitor c=0.0196365f //x=7.285 \
 //y=3.33 //x2=6.66 //y2=2.08
cc_2007 ( N_noxref_3_c_2007_p N_D_c_4253_n ) capacitor c=0.00117715f //x=7.515 \
 //y=3.33 //x2=6.66 //y2=2.08
cc_2008 ( N_noxref_3_c_1943_n N_D_c_4253_n ) capacitor c=0.0702997f //x=7.4 \
 //y=3.33 //x2=6.66 //y2=2.08
cc_2009 ( N_noxref_3_c_1944_n N_D_c_4253_n ) capacitor c=7.76771e-19 //x=9.25 \
 //y=2.08 //x2=6.66 //y2=2.08
cc_2010 ( N_noxref_3_c_1959_n N_D_M53_noxref_g ) capacitor c=0.0166421f \
 //x=6.835 //y=5.2 //x2=6.7 //y2=6.02
cc_2011 ( N_noxref_3_M53_noxref_d N_D_M53_noxref_g ) capacitor c=0.0173476f \
 //x=6.775 //y=5.02 //x2=6.7 //y2=6.02
cc_2012 ( N_noxref_3_c_1965_n N_D_M54_noxref_g ) capacitor c=0.018922f \
 //x=7.315 //y=5.2 //x2=7.14 //y2=6.02
cc_2013 ( N_noxref_3_M53_noxref_d N_D_M54_noxref_g ) capacitor c=0.0179769f \
 //x=6.775 //y=5.02 //x2=7.14 //y2=6.02
cc_2014 ( N_noxref_3_M4_noxref_d N_D_c_4299_n ) capacitor c=0.00217566f \
 //x=6.77 //y=0.905 //x2=6.695 //y2=0.905
cc_2015 ( N_noxref_3_M4_noxref_d N_D_c_4300_n ) capacitor c=0.0034598f \
 //x=6.77 //y=0.905 //x2=6.695 //y2=1.25
cc_2016 ( N_noxref_3_M4_noxref_d N_D_c_4301_n ) capacitor c=0.00656319f \
 //x=6.77 //y=0.905 //x2=6.695 //y2=1.56
cc_2017 ( N_noxref_3_c_1943_n N_D_c_4302_n ) capacitor c=0.0142673f //x=7.4 \
 //y=3.33 //x2=7.065 //y2=4.79
cc_2018 ( N_noxref_3_c_2099_p N_D_c_4302_n ) capacitor c=0.00407665f //x=6.92 \
 //y=5.2 //x2=7.065 //y2=4.79
cc_2019 ( N_noxref_3_M4_noxref_d N_D_c_4304_n ) capacitor c=0.00241102f \
 //x=6.77 //y=0.905 //x2=7.07 //y2=0.75
cc_2020 ( N_noxref_3_c_1942_n N_D_c_4305_n ) capacitor c=0.00359704f //x=7.315 \
 //y=1.655 //x2=7.07 //y2=1.405
cc_2021 ( N_noxref_3_M4_noxref_d N_D_c_4305_n ) capacitor c=0.0138845f \
 //x=6.77 //y=0.905 //x2=7.07 //y2=1.405
cc_2022 ( N_noxref_3_M4_noxref_d N_D_c_4307_n ) capacitor c=0.00132245f \
 //x=6.77 //y=0.905 //x2=7.225 //y2=0.905
cc_2023 ( N_noxref_3_c_1942_n N_D_c_4308_n ) capacitor c=0.00457401f //x=7.315 \
 //y=1.655 //x2=7.225 //y2=1.25
cc_2024 ( N_noxref_3_M4_noxref_d N_D_c_4308_n ) capacitor c=0.00566463f \
 //x=6.77 //y=0.905 //x2=7.225 //y2=1.25
cc_2025 ( N_noxref_3_c_1943_n N_D_c_4310_n ) capacitor c=0.00877984f //x=7.4 \
 //y=3.33 //x2=6.66 //y2=2.08
cc_2026 ( N_noxref_3_c_1943_n N_D_c_4311_n ) capacitor c=0.00306024f //x=7.4 \
 //y=3.33 //x2=6.66 //y2=1.915
cc_2027 ( N_noxref_3_M4_noxref_d N_D_c_4311_n ) capacitor c=0.00660593f \
 //x=6.77 //y=0.905 //x2=6.66 //y2=1.915
cc_2028 ( N_noxref_3_c_1959_n N_D_c_4313_n ) capacitor c=0.00346527f //x=6.835 \
 //y=5.2 //x2=6.69 //y2=4.7
cc_2029 ( N_noxref_3_c_1943_n N_D_c_4313_n ) capacitor c=0.00533692f //x=7.4 \
 //y=3.33 //x2=6.69 //y2=4.7
cc_2030 ( N_noxref_3_c_1935_n N_CLK_c_5034_n ) capacitor c=0.00360213f \
 //x=7.285 //y=3.33 //x2=13.205 //y2=4.44
cc_2031 ( N_noxref_3_c_1939_n N_CLK_c_5034_n ) capacitor c=4.49102e-19 \
 //x=3.445 //y=3.33 //x2=13.205 //y2=4.44
cc_2032 ( N_noxref_3_c_1941_n N_CLK_c_5034_n ) capacitor c=0.0200057f //x=3.33 \
 //y=2.08 //x2=13.205 //y2=4.44
cc_2033 ( N_noxref_3_c_1959_n N_CLK_c_5034_n ) capacitor c=0.0185297f \
 //x=6.835 //y=5.2 //x2=13.205 //y2=4.44
cc_2034 ( N_noxref_3_c_1963_n N_CLK_c_5034_n ) capacitor c=0.0181237f \
 //x=6.125 //y=5.2 //x2=13.205 //y2=4.44
cc_2035 ( N_noxref_3_c_1943_n N_CLK_c_5034_n ) capacitor c=0.0208321f //x=7.4 \
 //y=3.33 //x2=13.205 //y2=4.44
cc_2036 ( N_noxref_3_c_1944_n N_CLK_c_5034_n ) capacitor c=0.0198304f //x=9.25 \
 //y=2.08 //x2=13.205 //y2=4.44
cc_2037 ( N_noxref_3_c_2013_p N_CLK_c_5034_n ) capacitor c=0.0111881f //x=3.33 \
 //y=4.7 //x2=13.205 //y2=4.44
cc_2038 ( N_noxref_3_c_1982_n N_CLK_c_5034_n ) capacitor c=0.0107057f //x=9.25 \
 //y=4.7 //x2=13.205 //y2=4.44
cc_2039 ( N_noxref_3_c_1941_n N_CLK_c_5052_n ) capacitor c=0.00153281f \
 //x=3.33 //y=2.08 //x2=2.335 //y2=4.44
cc_2040 ( N_noxref_3_c_1939_n N_CLK_c_5025_n ) capacitor c=0.00526349f \
 //x=3.445 //y=3.33 //x2=2.22 //y2=2.08
cc_2041 ( N_noxref_3_c_1941_n N_CLK_c_5025_n ) capacitor c=0.0511464f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_2042 ( N_noxref_3_c_2021_p N_CLK_c_5025_n ) capacitor c=0.00228632f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=2.08
cc_2043 ( N_noxref_3_c_2013_p N_CLK_c_5025_n ) capacitor c=0.00218014f \
 //x=3.33 //y=4.7 //x2=2.22 //y2=2.08
cc_2044 ( N_noxref_3_M49_noxref_g N_CLK_M47_noxref_g ) capacitor c=0.0101598f \
 //x=3.07 //y=6.02 //x2=2.19 //y2=6.02
cc_2045 ( N_noxref_3_M49_noxref_g N_CLK_M48_noxref_g ) capacitor c=0.0602553f \
 //x=3.07 //y=6.02 //x2=2.63 //y2=6.02
cc_2046 ( N_noxref_3_M50_noxref_g N_CLK_M48_noxref_g ) capacitor c=0.0101598f \
 //x=3.51 //y=6.02 //x2=2.63 //y2=6.02
cc_2047 ( N_noxref_3_c_2034_p N_CLK_c_5187_n ) capacitor c=0.00456962f \
 //x=3.32 //y=0.915 //x2=2.31 //y2=0.91
cc_2048 ( N_noxref_3_c_2035_p N_CLK_c_5188_n ) capacitor c=0.00438372f \
 //x=3.32 //y=1.26 //x2=2.31 //y2=1.22
cc_2049 ( N_noxref_3_c_2036_p N_CLK_c_5189_n ) capacitor c=0.00438372f \
 //x=3.32 //y=1.57 //x2=2.31 //y2=1.45
cc_2050 ( N_noxref_3_c_1941_n N_CLK_c_5190_n ) capacitor c=0.0023343f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_2051 ( N_noxref_3_c_2021_p N_CLK_c_5190_n ) capacitor c=0.00933826f \
 //x=3.33 //y=2.08 //x2=2.31 //y2=1.915
cc_2052 ( N_noxref_3_c_2022_p N_CLK_c_5190_n ) capacitor c=0.00438372f \
 //x=3.33 //y=1.915 //x2=2.31 //y2=1.915
cc_2053 ( N_noxref_3_c_2013_p N_CLK_c_5193_n ) capacitor c=0.0611812f //x=3.33 \
 //y=4.7 //x2=2.555 //y2=4.79
cc_2054 ( N_noxref_3_c_1941_n N_CLK_c_5194_n ) capacitor c=0.00142741f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=4.7
cc_2055 ( N_noxref_3_c_2013_p N_CLK_c_5194_n ) capacitor c=0.00487508f \
 //x=3.33 //y=4.7 //x2=2.22 //y2=4.7
cc_2056 ( N_noxref_3_c_1935_n N_noxref_27_c_8266_n ) capacitor c=2.45218e-19 \
 //x=7.285 //y=3.33 //x2=3.985 //y2=0.54
cc_2057 ( N_noxref_3_c_1941_n N_noxref_27_c_8266_n ) capacitor c=0.00208521f \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_2058 ( N_noxref_3_c_2034_p N_noxref_27_c_8266_n ) capacitor c=0.0194423f \
 //x=3.32 //y=0.915 //x2=3.985 //y2=0.54
cc_2059 ( N_noxref_3_c_2039_p N_noxref_27_c_8266_n ) capacitor c=0.00656458f \
 //x=3.85 //y=0.915 //x2=3.985 //y2=0.54
cc_2060 ( N_noxref_3_c_2021_p N_noxref_27_c_8266_n ) capacitor c=2.20712e-19 \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_2061 ( N_noxref_3_c_2035_p N_noxref_27_c_8280_n ) capacitor c=0.00538829f \
 //x=3.32 //y=1.26 //x2=3.1 //y2=0.995
cc_2062 ( N_noxref_3_c_2034_p N_noxref_27_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=0.915 //x2=2.965 //y2=0.375
cc_2063 ( N_noxref_3_c_2036_p N_noxref_27_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=1.57 //x2=2.965 //y2=0.375
cc_2064 ( N_noxref_3_c_2039_p N_noxref_27_M2_noxref_s ) capacitor c=0.0143002f \
 //x=3.85 //y=0.915 //x2=2.965 //y2=0.375
cc_2065 ( N_noxref_3_c_2015_p N_noxref_27_M2_noxref_s ) capacitor \
 c=0.00290153f //x=3.85 //y=1.26 //x2=2.965 //y2=0.375
cc_2066 ( N_noxref_3_c_1935_n N_noxref_28_c_8333_n ) capacitor c=0.00241565f \
 //x=7.285 //y=3.33 //x2=5.505 //y2=1.495
cc_2067 ( N_noxref_3_c_2079_p N_noxref_28_c_8333_n ) capacitor c=3.15806e-19 \
 //x=7.045 //y=1.655 //x2=5.505 //y2=1.495
cc_2068 ( N_noxref_3_c_1935_n N_noxref_28_c_8314_n ) capacitor c=0.010299f \
 //x=7.285 //y=3.33 //x2=6.39 //y2=1.58
cc_2069 ( N_noxref_3_c_1935_n N_noxref_28_c_8321_n ) capacitor c=0.00177621f \
 //x=7.285 //y=3.33 //x2=6.475 //y2=1.495
cc_2070 ( N_noxref_3_c_2079_p N_noxref_28_c_8321_n ) capacitor c=0.020324f \
 //x=7.045 //y=1.655 //x2=6.475 //y2=1.495
cc_2071 ( N_noxref_3_c_1942_n N_noxref_28_c_8322_n ) capacitor c=0.00461444f \
 //x=7.315 //y=1.655 //x2=7.36 //y2=0.53
cc_2072 ( N_noxref_3_M4_noxref_d N_noxref_28_c_8322_n ) capacitor c=0.0116735f \
 //x=6.77 //y=0.905 //x2=7.36 //y2=0.53
cc_2073 ( N_noxref_3_c_1942_n N_noxref_28_M3_noxref_s ) capacitor c=0.0137901f \
 //x=7.315 //y=1.655 //x2=5.37 //y2=0.365
cc_2074 ( N_noxref_3_M4_noxref_d N_noxref_28_M3_noxref_s ) capacitor \
 c=0.0439476f //x=6.77 //y=0.905 //x2=5.37 //y2=0.365
cc_2075 ( N_noxref_3_c_1942_n N_noxref_29_c_8387_n ) capacitor c=3.22188e-19 \
 //x=7.315 //y=1.655 //x2=8.835 //y2=1.495
cc_2076 ( N_noxref_3_c_1949_n N_noxref_29_c_8387_n ) capacitor c=0.0034165f \
 //x=9.055 //y=1.915 //x2=8.835 //y2=1.495
cc_2077 ( N_noxref_3_c_1944_n N_noxref_29_c_8368_n ) capacitor c=0.0118762f \
 //x=9.25 //y=2.08 //x2=9.72 //y2=1.58
cc_2078 ( N_noxref_3_c_1948_n N_noxref_29_c_8368_n ) capacitor c=0.00703567f \
 //x=9.055 //y=1.52 //x2=9.72 //y2=1.58
cc_2079 ( N_noxref_3_c_1949_n N_noxref_29_c_8368_n ) capacitor c=0.018562f \
 //x=9.055 //y=1.915 //x2=9.72 //y2=1.58
cc_2080 ( N_noxref_3_c_1951_n N_noxref_29_c_8368_n ) capacitor c=0.00780629f \
 //x=9.43 //y=1.365 //x2=9.72 //y2=1.58
cc_2081 ( N_noxref_3_c_1954_n N_noxref_29_c_8368_n ) capacitor c=0.00339872f \
 //x=9.585 //y=1.21 //x2=9.72 //y2=1.58
cc_2082 ( N_noxref_3_c_1949_n N_noxref_29_c_8375_n ) capacitor c=6.71402e-19 \
 //x=9.055 //y=1.915 //x2=9.805 //y2=1.495
cc_2083 ( N_noxref_3_c_1945_n N_noxref_29_M5_noxref_s ) capacitor c=0.0326577f \
 //x=9.055 //y=0.865 //x2=8.7 //y2=0.365
cc_2084 ( N_noxref_3_c_1948_n N_noxref_29_M5_noxref_s ) capacitor \
 c=3.48408e-19 //x=9.055 //y=1.52 //x2=8.7 //y2=0.365
cc_2085 ( N_noxref_3_c_1952_n N_noxref_29_M5_noxref_s ) capacitor c=0.0120759f \
 //x=9.585 //y=0.865 //x2=8.7 //y2=0.365
cc_2086 ( N_noxref_4_c_2167_n N_noxref_5_c_2317_n ) capacitor c=0.175696f \
 //x=12.465 //y=3.33 //x2=15.795 //y2=3.7
cc_2087 ( N_noxref_4_c_2215_n N_noxref_5_c_2317_n ) capacitor c=0.0293967f \
 //x=10.845 //y=3.33 //x2=15.795 //y2=3.7
cc_2088 ( N_noxref_4_c_2169_n N_noxref_5_c_2317_n ) capacitor c=0.0206034f \
 //x=10.73 //y=3.33 //x2=15.795 //y2=3.7
cc_2089 ( N_noxref_4_c_2170_n N_noxref_5_c_2317_n ) capacitor c=0.0205831f \
 //x=12.58 //y=2.08 //x2=15.795 //y2=3.7
cc_2090 ( N_noxref_4_c_2167_n N_noxref_7_c_2744_n ) capacitor c=0.0110241f \
 //x=12.465 //y=3.33 //x2=13.945 //y2=4.07
cc_2091 ( N_noxref_4_c_2215_n N_noxref_7_c_2744_n ) capacitor c=8.88358e-19 \
 //x=10.845 //y=3.33 //x2=13.945 //y2=4.07
cc_2092 ( N_noxref_4_c_2169_n N_noxref_7_c_2744_n ) capacitor c=0.0181936f \
 //x=10.73 //y=3.33 //x2=13.945 //y2=4.07
cc_2093 ( N_noxref_4_c_2170_n N_noxref_7_c_2744_n ) capacitor c=0.0184765f \
 //x=12.58 //y=2.08 //x2=13.945 //y2=4.07
cc_2094 ( N_noxref_4_c_2169_n N_noxref_7_c_2801_n ) capacitor c=0.00117715f \
 //x=10.73 //y=3.33 //x2=10.105 //y2=4.07
cc_2095 ( N_noxref_4_c_2184_n N_noxref_7_c_2803_n ) capacitor c=0.0126603f \
 //x=10.165 //y=5.2 //x2=9.99 //y2=4.535
cc_2096 ( N_noxref_4_c_2169_n N_noxref_7_c_2803_n ) capacitor c=0.0101319f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=4.535
cc_2097 ( N_noxref_4_c_2215_n N_noxref_7_c_2718_n ) capacitor c=0.00329059f \
 //x=10.845 //y=3.33 //x2=9.99 //y2=2.08
cc_2098 ( N_noxref_4_c_2169_n N_noxref_7_c_2718_n ) capacitor c=0.0717703f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=2.08
cc_2099 ( N_noxref_4_c_2170_n N_noxref_7_c_2718_n ) capacitor c=9.69022e-19 \
 //x=12.58 //y=2.08 //x2=9.99 //y2=2.08
cc_2100 ( N_noxref_4_M60_noxref_g N_noxref_7_c_2753_n ) capacitor c=0.0169521f \
 //x=12.92 //y=6.02 //x2=13.495 //y2=5.2
cc_2101 ( N_noxref_4_c_2170_n N_noxref_7_c_2757_n ) capacitor c=0.00539951f \
 //x=12.58 //y=2.08 //x2=12.785 //y2=5.2
cc_2102 ( N_noxref_4_M59_noxref_g N_noxref_7_c_2757_n ) capacitor c=0.0177326f \
 //x=12.48 //y=6.02 //x2=12.785 //y2=5.2
cc_2103 ( N_noxref_4_c_2203_n N_noxref_7_c_2757_n ) capacitor c=0.00581252f \
 //x=12.58 //y=4.7 //x2=12.785 //y2=5.2
cc_2104 ( N_noxref_4_c_2169_n N_noxref_7_c_2721_n ) capacitor c=3.49822e-19 \
 //x=10.73 //y=3.33 //x2=14.06 //y2=4.07
cc_2105 ( N_noxref_4_c_2170_n N_noxref_7_c_2721_n ) capacitor c=0.0034438f \
 //x=12.58 //y=2.08 //x2=14.06 //y2=4.07
cc_2106 ( N_noxref_4_c_2184_n N_noxref_7_M57_noxref_g ) capacitor c=0.0166421f \
 //x=10.165 //y=5.2 //x2=10.03 //y2=6.02
cc_2107 ( N_noxref_4_M57_noxref_d N_noxref_7_M57_noxref_g ) capacitor \
 c=0.0173476f //x=10.105 //y=5.02 //x2=10.03 //y2=6.02
cc_2108 ( N_noxref_4_c_2190_n N_noxref_7_M58_noxref_g ) capacitor c=0.018922f \
 //x=10.645 //y=5.2 //x2=10.47 //y2=6.02
cc_2109 ( N_noxref_4_M57_noxref_d N_noxref_7_M58_noxref_g ) capacitor \
 c=0.0179769f //x=10.105 //y=5.02 //x2=10.47 //y2=6.02
cc_2110 ( N_noxref_4_M6_noxref_d N_noxref_7_c_2812_n ) capacitor c=0.00217566f \
 //x=10.1 //y=0.905 //x2=10.025 //y2=0.905
cc_2111 ( N_noxref_4_M6_noxref_d N_noxref_7_c_2815_n ) capacitor c=0.0034598f \
 //x=10.1 //y=0.905 //x2=10.025 //y2=1.25
cc_2112 ( N_noxref_4_M6_noxref_d N_noxref_7_c_2817_n ) capacitor c=0.00656319f \
 //x=10.1 //y=0.905 //x2=10.025 //y2=1.56
cc_2113 ( N_noxref_4_c_2169_n N_noxref_7_c_2849_n ) capacitor c=0.0142673f \
 //x=10.73 //y=3.33 //x2=10.395 //y2=4.79
cc_2114 ( N_noxref_4_c_2251_p N_noxref_7_c_2849_n ) capacitor c=0.00407665f \
 //x=10.25 //y=5.2 //x2=10.395 //y2=4.79
cc_2115 ( N_noxref_4_M6_noxref_d N_noxref_7_c_2851_n ) capacitor c=0.00241102f \
 //x=10.1 //y=0.905 //x2=10.4 //y2=0.75
cc_2116 ( N_noxref_4_c_2168_n N_noxref_7_c_2852_n ) capacitor c=0.00359704f \
 //x=10.645 //y=1.655 //x2=10.4 //y2=1.405
cc_2117 ( N_noxref_4_M6_noxref_d N_noxref_7_c_2852_n ) capacitor c=0.0138845f \
 //x=10.1 //y=0.905 //x2=10.4 //y2=1.405
cc_2118 ( N_noxref_4_M6_noxref_d N_noxref_7_c_2820_n ) capacitor c=0.00132245f \
 //x=10.1 //y=0.905 //x2=10.555 //y2=0.905
cc_2119 ( N_noxref_4_c_2168_n N_noxref_7_c_2821_n ) capacitor c=0.00457401f \
 //x=10.645 //y=1.655 //x2=10.555 //y2=1.25
cc_2120 ( N_noxref_4_M6_noxref_d N_noxref_7_c_2821_n ) capacitor c=0.00566463f \
 //x=10.1 //y=0.905 //x2=10.555 //y2=1.25
cc_2121 ( N_noxref_4_c_2169_n N_noxref_7_c_2822_n ) capacitor c=0.00877984f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=2.08
cc_2122 ( N_noxref_4_c_2169_n N_noxref_7_c_2858_n ) capacitor c=0.00306024f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=1.915
cc_2123 ( N_noxref_4_M6_noxref_d N_noxref_7_c_2858_n ) capacitor c=0.00660593f \
 //x=10.1 //y=0.905 //x2=9.99 //y2=1.915
cc_2124 ( N_noxref_4_c_2184_n N_noxref_7_c_2824_n ) capacitor c=0.00346527f \
 //x=10.165 //y=5.2 //x2=10.02 //y2=4.7
cc_2125 ( N_noxref_4_c_2169_n N_noxref_7_c_2824_n ) capacitor c=0.00517969f \
 //x=10.73 //y=3.33 //x2=10.02 //y2=4.7
cc_2126 ( N_noxref_4_M60_noxref_g N_noxref_7_M59_noxref_d ) capacitor \
 c=0.0173476f //x=12.92 //y=6.02 //x2=12.555 //y2=5.02
cc_2127 ( N_noxref_4_c_2167_n N_D_c_4217_n ) capacitor c=0.083897f //x=12.465 \
 //y=3.33 //x2=28.005 //y2=2.59
cc_2128 ( N_noxref_4_c_2215_n N_D_c_4217_n ) capacitor c=0.0133398f //x=10.845 \
 //y=3.33 //x2=28.005 //y2=2.59
cc_2129 ( N_noxref_4_c_2266_p N_D_c_4217_n ) capacitor c=0.0102711f //x=10.375 \
 //y=1.655 //x2=28.005 //y2=2.59
cc_2130 ( N_noxref_4_c_2169_n N_D_c_4217_n ) capacitor c=0.0237178f //x=10.73 \
 //y=3.33 //x2=28.005 //y2=2.59
cc_2131 ( N_noxref_4_c_2170_n N_D_c_4217_n ) capacitor c=0.0239823f //x=12.58 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2132 ( N_noxref_4_c_2175_n N_D_c_4217_n ) capacitor c=0.00424331f \
 //x=12.385 //y=1.915 //x2=28.005 //y2=2.59
cc_2133 ( N_noxref_4_c_2184_n N_CLK_c_5034_n ) capacitor c=0.0185297f \
 //x=10.165 //y=5.2 //x2=13.205 //y2=4.44
cc_2134 ( N_noxref_4_c_2188_n N_CLK_c_5034_n ) capacitor c=0.018142f //x=9.455 \
 //y=5.2 //x2=13.205 //y2=4.44
cc_2135 ( N_noxref_4_c_2169_n N_CLK_c_5034_n ) capacitor c=0.0208321f \
 //x=10.73 //y=3.33 //x2=13.205 //y2=4.44
cc_2136 ( N_noxref_4_c_2170_n N_CLK_c_5034_n ) capacitor c=0.0198304f \
 //x=12.58 //y=2.08 //x2=13.205 //y2=4.44
cc_2137 ( N_noxref_4_c_2203_n N_CLK_c_5034_n ) capacitor c=0.0107057f \
 //x=12.58 //y=4.7 //x2=13.205 //y2=4.44
cc_2138 ( N_noxref_4_c_2170_n N_CLK_c_5060_n ) capacitor c=0.00168329f \
 //x=12.58 //y=2.08 //x2=13.465 //y2=4.442
cc_2139 ( N_noxref_4_c_2203_n N_CLK_c_5060_n ) capacitor c=2.91071e-19 \
 //x=12.58 //y=4.7 //x2=13.465 //y2=4.442
cc_2140 ( N_noxref_4_c_2170_n N_CLK_c_5203_n ) capacitor c=0.00400249f \
 //x=12.58 //y=2.08 //x2=13.32 //y2=4.535
cc_2141 ( N_noxref_4_c_2203_n N_CLK_c_5203_n ) capacitor c=0.00415951f \
 //x=12.58 //y=4.7 //x2=13.32 //y2=4.535
cc_2142 ( N_noxref_4_c_2167_n N_CLK_c_5026_n ) capacitor c=0.00720056f \
 //x=12.465 //y=3.33 //x2=13.32 //y2=2.08
cc_2143 ( N_noxref_4_c_2169_n N_CLK_c_5026_n ) capacitor c=0.00102338f \
 //x=10.73 //y=3.33 //x2=13.32 //y2=2.08
cc_2144 ( N_noxref_4_c_2170_n N_CLK_c_5026_n ) capacitor c=0.0760595f \
 //x=12.58 //y=2.08 //x2=13.32 //y2=2.08
cc_2145 ( N_noxref_4_c_2175_n N_CLK_c_5026_n ) capacitor c=0.00308814f \
 //x=12.385 //y=1.915 //x2=13.32 //y2=2.08
cc_2146 ( N_noxref_4_M59_noxref_g N_CLK_M61_noxref_g ) capacitor c=0.0104611f \
 //x=12.48 //y=6.02 //x2=13.36 //y2=6.02
cc_2147 ( N_noxref_4_M60_noxref_g N_CLK_M61_noxref_g ) capacitor c=0.106811f \
 //x=12.92 //y=6.02 //x2=13.36 //y2=6.02
cc_2148 ( N_noxref_4_M60_noxref_g N_CLK_M62_noxref_g ) capacitor c=0.0100341f \
 //x=12.92 //y=6.02 //x2=13.8 //y2=6.02
cc_2149 ( N_noxref_4_c_2171_n N_CLK_c_5212_n ) capacitor c=4.86506e-19 \
 //x=12.385 //y=0.865 //x2=13.355 //y2=0.905
cc_2150 ( N_noxref_4_c_2173_n N_CLK_c_5212_n ) capacitor c=0.00152104f \
 //x=12.385 //y=1.21 //x2=13.355 //y2=0.905
cc_2151 ( N_noxref_4_c_2178_n N_CLK_c_5212_n ) capacitor c=0.0151475f \
 //x=12.915 //y=0.865 //x2=13.355 //y2=0.905
cc_2152 ( N_noxref_4_c_2174_n N_CLK_c_5215_n ) capacitor c=0.00109982f \
 //x=12.385 //y=1.52 //x2=13.355 //y2=1.25
cc_2153 ( N_noxref_4_c_2180_n N_CLK_c_5215_n ) capacitor c=0.0111064f \
 //x=12.915 //y=1.21 //x2=13.355 //y2=1.25
cc_2154 ( N_noxref_4_c_2174_n N_CLK_c_5217_n ) capacitor c=9.57794e-19 \
 //x=12.385 //y=1.52 //x2=13.355 //y2=1.56
cc_2155 ( N_noxref_4_c_2175_n N_CLK_c_5217_n ) capacitor c=0.00662747f \
 //x=12.385 //y=1.915 //x2=13.355 //y2=1.56
cc_2156 ( N_noxref_4_c_2180_n N_CLK_c_5217_n ) capacitor c=0.00862358f \
 //x=12.915 //y=1.21 //x2=13.355 //y2=1.56
cc_2157 ( N_noxref_4_c_2178_n N_CLK_c_5220_n ) capacitor c=0.00124821f \
 //x=12.915 //y=0.865 //x2=13.885 //y2=0.905
cc_2158 ( N_noxref_4_c_2180_n N_CLK_c_5221_n ) capacitor c=0.00200715f \
 //x=12.915 //y=1.21 //x2=13.885 //y2=1.25
cc_2159 ( N_noxref_4_c_2170_n N_CLK_c_5222_n ) capacitor c=0.00307062f \
 //x=12.58 //y=2.08 //x2=13.32 //y2=2.08
cc_2160 ( N_noxref_4_c_2175_n N_CLK_c_5222_n ) capacitor c=0.0179092f \
 //x=12.385 //y=1.915 //x2=13.32 //y2=2.08
cc_2161 ( N_noxref_4_c_2170_n N_CLK_c_5224_n ) capacitor c=0.00342116f \
 //x=12.58 //y=2.08 //x2=13.35 //y2=4.7
cc_2162 ( N_noxref_4_c_2203_n N_CLK_c_5224_n ) capacitor c=0.0292158f \
 //x=12.58 //y=4.7 //x2=13.35 //y2=4.7
cc_2163 ( N_noxref_4_c_2266_p N_noxref_29_c_8387_n ) capacitor c=3.15806e-19 \
 //x=10.375 //y=1.655 //x2=8.835 //y2=1.495
cc_2164 ( N_noxref_4_c_2266_p N_noxref_29_c_8375_n ) capacitor c=0.0203424f \
 //x=10.375 //y=1.655 //x2=9.805 //y2=1.495
cc_2165 ( N_noxref_4_c_2168_n N_noxref_29_c_8376_n ) capacitor c=0.00461444f \
 //x=10.645 //y=1.655 //x2=10.69 //y2=0.53
cc_2166 ( N_noxref_4_M6_noxref_d N_noxref_29_c_8376_n ) capacitor c=0.0116735f \
 //x=10.1 //y=0.905 //x2=10.69 //y2=0.53
cc_2167 ( N_noxref_4_c_2168_n N_noxref_29_M5_noxref_s ) capacitor c=0.0137901f \
 //x=10.645 //y=1.655 //x2=8.7 //y2=0.365
cc_2168 ( N_noxref_4_M6_noxref_d N_noxref_29_M5_noxref_s ) capacitor \
 c=0.043966f //x=10.1 //y=0.905 //x2=8.7 //y2=0.365
cc_2169 ( N_noxref_4_c_2168_n N_noxref_30_c_8439_n ) capacitor c=3.22188e-19 \
 //x=10.645 //y=1.655 //x2=12.165 //y2=1.495
cc_2170 ( N_noxref_4_c_2175_n N_noxref_30_c_8439_n ) capacitor c=0.0034165f \
 //x=12.385 //y=1.915 //x2=12.165 //y2=1.495
cc_2171 ( N_noxref_4_c_2170_n N_noxref_30_c_8420_n ) capacitor c=0.0118762f \
 //x=12.58 //y=2.08 //x2=13.05 //y2=1.58
cc_2172 ( N_noxref_4_c_2174_n N_noxref_30_c_8420_n ) capacitor c=0.00703567f \
 //x=12.385 //y=1.52 //x2=13.05 //y2=1.58
cc_2173 ( N_noxref_4_c_2175_n N_noxref_30_c_8420_n ) capacitor c=0.018562f \
 //x=12.385 //y=1.915 //x2=13.05 //y2=1.58
cc_2174 ( N_noxref_4_c_2177_n N_noxref_30_c_8420_n ) capacitor c=0.00780629f \
 //x=12.76 //y=1.365 //x2=13.05 //y2=1.58
cc_2175 ( N_noxref_4_c_2180_n N_noxref_30_c_8420_n ) capacitor c=0.00339872f \
 //x=12.915 //y=1.21 //x2=13.05 //y2=1.58
cc_2176 ( N_noxref_4_c_2175_n N_noxref_30_c_8427_n ) capacitor c=6.71402e-19 \
 //x=12.385 //y=1.915 //x2=13.135 //y2=1.495
cc_2177 ( N_noxref_4_c_2171_n N_noxref_30_M7_noxref_s ) capacitor c=0.0326577f \
 //x=12.385 //y=0.865 //x2=12.03 //y2=0.365
cc_2178 ( N_noxref_4_c_2174_n N_noxref_30_M7_noxref_s ) capacitor \
 c=3.48408e-19 //x=12.385 //y=1.52 //x2=12.03 //y2=0.365
cc_2179 ( N_noxref_4_c_2178_n N_noxref_30_M7_noxref_s ) capacitor c=0.0120759f \
 //x=12.915 //y=0.865 //x2=12.03 //y2=0.365
cc_2180 ( N_noxref_5_c_2317_n N_noxref_6_c_2612_n ) capacitor c=0.0114735f \
 //x=15.795 //y=3.7 //x2=17.505 //y2=3.7
cc_2181 ( N_noxref_5_M64_noxref_g N_noxref_6_c_2581_n ) capacitor c=0.0169675f \
 //x=16.25 //y=6.02 //x2=16.825 //y2=5.2
cc_2182 ( N_noxref_5_c_2320_n N_noxref_6_c_2585_n ) capacitor c=0.00521711f \
 //x=15.91 //y=2.08 //x2=16.115 //y2=5.2
cc_2183 ( N_noxref_5_M63_noxref_g N_noxref_6_c_2585_n ) capacitor c=0.0177326f \
 //x=15.81 //y=6.02 //x2=16.115 //y2=5.2
cc_2184 ( N_noxref_5_c_2372_n N_noxref_6_c_2585_n ) capacitor c=0.00581264f \
 //x=15.91 //y=4.7 //x2=16.115 //y2=5.2
cc_2185 ( N_noxref_5_c_2320_n N_noxref_6_c_2566_n ) capacitor c=0.00334373f \
 //x=15.91 //y=2.08 //x2=17.39 //y2=3.7
cc_2186 ( N_noxref_5_M64_noxref_g N_noxref_6_M63_noxref_d ) capacitor \
 c=0.0173476f //x=16.25 //y=6.02 //x2=15.885 //y2=5.02
cc_2187 ( N_noxref_5_c_2388_n N_noxref_7_c_2715_n ) capacitor c=0.147021f \
 //x=5.805 //y=3.7 //x2=9.875 //y2=4.07
cc_2188 ( N_noxref_5_c_2389_n N_noxref_7_c_2715_n ) capacitor c=0.0294294f \
 //x=4.185 //y=3.7 //x2=9.875 //y2=4.07
cc_2189 ( N_noxref_5_c_2317_n N_noxref_7_c_2715_n ) capacitor c=0.338937f \
 //x=15.795 //y=3.7 //x2=9.875 //y2=4.07
cc_2190 ( N_noxref_5_c_2396_n N_noxref_7_c_2715_n ) capacitor c=0.0264478f \
 //x=6.035 //y=3.7 //x2=9.875 //y2=4.07
cc_2191 ( N_noxref_5_c_2346_n N_noxref_7_c_2715_n ) capacitor c=0.0154449f \
 //x=1.615 //y=5.155 //x2=9.875 //y2=4.07
cc_2192 ( N_noxref_5_c_2356_n N_noxref_7_c_2715_n ) capacitor c=0.0200328f \
 //x=4.07 //y=3.7 //x2=9.875 //y2=4.07
cc_2193 ( N_noxref_5_c_2319_n N_noxref_7_c_2715_n ) capacitor c=0.0203111f \
 //x=5.92 //y=2.08 //x2=9.875 //y2=4.07
cc_2194 ( N_noxref_5_c_2317_n N_noxref_7_c_2744_n ) capacitor c=0.339146f \
 //x=15.795 //y=3.7 //x2=13.945 //y2=4.07
cc_2195 ( N_noxref_5_c_2317_n N_noxref_7_c_2801_n ) capacitor c=0.0267832f \
 //x=15.795 //y=3.7 //x2=10.105 //y2=4.07
cc_2196 ( N_noxref_5_c_2317_n N_noxref_7_c_2745_n ) capacitor c=0.176049f \
 //x=15.795 //y=3.7 //x2=19.865 //y2=4.07
cc_2197 ( N_noxref_5_c_2320_n N_noxref_7_c_2745_n ) capacitor c=0.0203675f \
 //x=15.91 //y=2.08 //x2=19.865 //y2=4.07
cc_2198 ( N_noxref_5_c_2317_n N_noxref_7_c_2747_n ) capacitor c=0.0266833f \
 //x=15.795 //y=3.7 //x2=14.175 //y2=4.07
cc_2199 ( N_noxref_5_c_2320_n N_noxref_7_c_2747_n ) capacitor c=3.50683e-19 \
 //x=15.91 //y=2.08 //x2=14.175 //y2=4.07
cc_2200 ( N_noxref_5_c_2317_n N_noxref_7_c_2718_n ) capacitor c=0.0226566f \
 //x=15.795 //y=3.7 //x2=9.99 //y2=2.08
cc_2201 ( N_noxref_5_c_2317_n N_noxref_7_c_2721_n ) capacitor c=0.0250326f \
 //x=15.795 //y=3.7 //x2=14.06 //y2=4.07
cc_2202 ( N_noxref_5_c_2320_n N_noxref_7_c_2721_n ) capacitor c=0.0139373f \
 //x=15.91 //y=2.08 //x2=14.06 //y2=4.07
cc_2203 ( N_noxref_5_c_2346_n N_noxref_7_M45_noxref_g ) capacitor c=0.0213876f \
 //x=1.615 //y=5.155 //x2=1.31 //y2=6.02
cc_2204 ( N_noxref_5_c_2342_n N_noxref_7_M46_noxref_g ) capacitor c=0.0178794f \
 //x=2.325 //y=5.155 //x2=1.75 //y2=6.02
cc_2205 ( N_noxref_5_M45_noxref_d N_noxref_7_M46_noxref_g ) capacitor \
 c=0.0180032f //x=1.385 //y=5.02 //x2=1.75 //y2=6.02
cc_2206 ( N_noxref_5_c_2346_n N_noxref_7_c_2882_n ) capacitor c=0.00429591f \
 //x=1.615 //y=5.155 //x2=1.675 //y2=4.79
cc_2207 ( N_noxref_5_c_2317_n N_D_c_4217_n ) capacitor c=0.146448f //x=15.795 \
 //y=3.7 //x2=28.005 //y2=2.59
cc_2208 ( N_noxref_5_c_2320_n N_D_c_4217_n ) capacitor c=0.025277f //x=15.91 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2209 ( N_noxref_5_c_2335_n N_D_c_4217_n ) capacitor c=0.00396741f \
 //x=15.715 //y=1.915 //x2=28.005 //y2=2.59
cc_2210 ( N_noxref_5_c_2317_n N_D_c_4236_n ) capacitor c=6.75065e-19 \
 //x=15.795 //y=3.7 //x2=6.775 //y2=2.59
cc_2211 ( N_noxref_5_c_2319_n N_D_c_4236_n ) capacitor c=0.00735597f //x=5.92 \
 //y=2.08 //x2=6.775 //y2=2.59
cc_2212 ( N_noxref_5_c_2319_n N_D_c_4289_n ) capacitor c=0.00400249f //x=5.92 \
 //y=2.08 //x2=6.66 //y2=4.535
cc_2213 ( N_noxref_5_c_2371_n N_D_c_4289_n ) capacitor c=0.00417994f //x=5.92 \
 //y=4.7 //x2=6.66 //y2=4.535
cc_2214 ( N_noxref_5_c_2317_n N_D_c_4253_n ) capacitor c=0.0169594f //x=15.795 \
 //y=3.7 //x2=6.66 //y2=2.08
cc_2215 ( N_noxref_5_c_2396_n N_D_c_4253_n ) capacitor c=0.00131333f //x=6.035 \
 //y=3.7 //x2=6.66 //y2=2.08
cc_2216 ( N_noxref_5_c_2356_n N_D_c_4253_n ) capacitor c=8.12815e-19 //x=4.07 \
 //y=3.7 //x2=6.66 //y2=2.08
cc_2217 ( N_noxref_5_c_2319_n N_D_c_4253_n ) capacitor c=0.0761047f //x=5.92 \
 //y=2.08 //x2=6.66 //y2=2.08
cc_2218 ( N_noxref_5_c_2325_n N_D_c_4253_n ) capacitor c=0.00308814f //x=5.725 \
 //y=1.915 //x2=6.66 //y2=2.08
cc_2219 ( N_noxref_5_M51_noxref_g N_D_M53_noxref_g ) capacitor c=0.0104611f \
 //x=5.82 //y=6.02 //x2=6.7 //y2=6.02
cc_2220 ( N_noxref_5_M52_noxref_g N_D_M53_noxref_g ) capacitor c=0.106811f \
 //x=6.26 //y=6.02 //x2=6.7 //y2=6.02
cc_2221 ( N_noxref_5_M52_noxref_g N_D_M54_noxref_g ) capacitor c=0.0100341f \
 //x=6.26 //y=6.02 //x2=7.14 //y2=6.02
cc_2222 ( N_noxref_5_c_2321_n N_D_c_4299_n ) capacitor c=4.86506e-19 //x=5.725 \
 //y=0.865 //x2=6.695 //y2=0.905
cc_2223 ( N_noxref_5_c_2323_n N_D_c_4299_n ) capacitor c=0.00152104f //x=5.725 \
 //y=1.21 //x2=6.695 //y2=0.905
cc_2224 ( N_noxref_5_c_2328_n N_D_c_4299_n ) capacitor c=0.0151475f //x=6.255 \
 //y=0.865 //x2=6.695 //y2=0.905
cc_2225 ( N_noxref_5_c_2324_n N_D_c_4300_n ) capacitor c=0.00109982f //x=5.725 \
 //y=1.52 //x2=6.695 //y2=1.25
cc_2226 ( N_noxref_5_c_2330_n N_D_c_4300_n ) capacitor c=0.0111064f //x=6.255 \
 //y=1.21 //x2=6.695 //y2=1.25
cc_2227 ( N_noxref_5_c_2324_n N_D_c_4301_n ) capacitor c=9.57794e-19 //x=5.725 \
 //y=1.52 //x2=6.695 //y2=1.56
cc_2228 ( N_noxref_5_c_2325_n N_D_c_4301_n ) capacitor c=0.00662747f //x=5.725 \
 //y=1.915 //x2=6.695 //y2=1.56
cc_2229 ( N_noxref_5_c_2330_n N_D_c_4301_n ) capacitor c=0.00862358f //x=6.255 \
 //y=1.21 //x2=6.695 //y2=1.56
cc_2230 ( N_noxref_5_c_2328_n N_D_c_4307_n ) capacitor c=0.00124821f //x=6.255 \
 //y=0.865 //x2=7.225 //y2=0.905
cc_2231 ( N_noxref_5_c_2330_n N_D_c_4308_n ) capacitor c=0.00200715f //x=6.255 \
 //y=1.21 //x2=7.225 //y2=1.25
cc_2232 ( N_noxref_5_c_2319_n N_D_c_4310_n ) capacitor c=0.00307062f //x=5.92 \
 //y=2.08 //x2=6.66 //y2=2.08
cc_2233 ( N_noxref_5_c_2325_n N_D_c_4310_n ) capacitor c=0.0179092f //x=5.725 \
 //y=1.915 //x2=6.66 //y2=2.08
cc_2234 ( N_noxref_5_c_2319_n N_D_c_4313_n ) capacitor c=0.00344981f //x=5.92 \
 //y=2.08 //x2=6.69 //y2=4.7
cc_2235 ( N_noxref_5_c_2371_n N_D_c_4313_n ) capacitor c=0.0293367f //x=5.92 \
 //y=4.7 //x2=6.69 //y2=4.7
cc_2236 ( N_noxref_5_c_2388_n N_CLK_c_5034_n ) capacitor c=0.00940379f \
 //x=5.805 //y=3.7 //x2=13.205 //y2=4.44
cc_2237 ( N_noxref_5_c_2389_n N_CLK_c_5034_n ) capacitor c=7.95009e-19 \
 //x=4.185 //y=3.7 //x2=13.205 //y2=4.44
cc_2238 ( N_noxref_5_c_2317_n N_CLK_c_5034_n ) capacitor c=0.0485341f \
 //x=15.795 //y=3.7 //x2=13.205 //y2=4.44
cc_2239 ( N_noxref_5_c_2396_n N_CLK_c_5034_n ) capacitor c=6.59192e-19 \
 //x=6.035 //y=3.7 //x2=13.205 //y2=4.44
cc_2240 ( N_noxref_5_c_2352_n N_CLK_c_5034_n ) capacitor c=0.0183122f \
 //x=3.985 //y=5.155 //x2=13.205 //y2=4.44
cc_2241 ( N_noxref_5_c_2356_n N_CLK_c_5034_n ) capacitor c=0.0210274f //x=4.07 \
 //y=3.7 //x2=13.205 //y2=4.44
cc_2242 ( N_noxref_5_c_2319_n N_CLK_c_5034_n ) capacitor c=0.0198304f //x=5.92 \
 //y=2.08 //x2=13.205 //y2=4.44
cc_2243 ( N_noxref_5_c_2497_p N_CLK_c_5034_n ) capacitor c=0.0311227f //x=2.41 \
 //y=5.155 //x2=13.205 //y2=4.44
cc_2244 ( N_noxref_5_c_2371_n N_CLK_c_5034_n ) capacitor c=0.0107057f //x=5.92 \
 //y=4.7 //x2=13.205 //y2=4.44
cc_2245 ( N_noxref_5_c_2342_n N_CLK_c_5052_n ) capacitor c=0.00330099f \
 //x=2.325 //y=5.155 //x2=2.335 //y2=4.44
cc_2246 ( N_noxref_5_c_2317_n N_CLK_c_5053_n ) capacitor c=0.0155891f \
 //x=15.795 //y=3.7 //x2=16.745 //y2=4.442
cc_2247 ( N_noxref_5_c_2320_n N_CLK_c_5053_n ) capacitor c=0.0187387f \
 //x=15.91 //y=2.08 //x2=16.745 //y2=4.442
cc_2248 ( N_noxref_5_c_2372_n N_CLK_c_5053_n ) capacitor c=0.0104218f \
 //x=15.91 //y=4.7 //x2=16.745 //y2=4.442
cc_2249 ( N_noxref_5_c_2317_n N_CLK_c_5060_n ) capacitor c=7.37075e-19 \
 //x=15.795 //y=3.7 //x2=13.465 //y2=4.442
cc_2250 ( N_noxref_5_c_2342_n N_CLK_c_5025_n ) capacitor c=0.014564f //x=2.325 \
 //y=5.155 //x2=2.22 //y2=2.08
cc_2251 ( N_noxref_5_c_2356_n N_CLK_c_5025_n ) capacitor c=0.00319363f \
 //x=4.07 //y=3.7 //x2=2.22 //y2=2.08
cc_2252 ( N_noxref_5_c_2317_n N_CLK_c_5026_n ) capacitor c=0.0208196f \
 //x=15.795 //y=3.7 //x2=13.32 //y2=2.08
cc_2253 ( N_noxref_5_c_2320_n N_CLK_c_5026_n ) capacitor c=0.00128802f \
 //x=15.91 //y=2.08 //x2=13.32 //y2=2.08
cc_2254 ( N_noxref_5_c_2342_n N_CLK_M47_noxref_g ) capacitor c=0.016514f \
 //x=2.325 //y=5.155 //x2=2.19 //y2=6.02
cc_2255 ( N_noxref_5_M47_noxref_d N_CLK_M47_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.19 //y2=6.02
cc_2256 ( N_noxref_5_c_2348_n N_CLK_M48_noxref_g ) capacitor c=0.01736f \
 //x=3.205 //y=5.155 //x2=2.63 //y2=6.02
cc_2257 ( N_noxref_5_M47_noxref_d N_CLK_M48_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.63 //y2=6.02
cc_2258 ( N_noxref_5_c_2497_p N_CLK_c_5193_n ) capacitor c=0.00426767f \
 //x=2.41 //y=5.155 //x2=2.555 //y2=4.79
cc_2259 ( N_noxref_5_c_2342_n N_CLK_c_5194_n ) capacitor c=0.00322046f \
 //x=2.325 //y=5.155 //x2=2.22 //y2=4.7
cc_2260 ( N_noxref_5_c_2320_n N_noxref_23_c_7578_n ) capacitor c=0.00735597f \
 //x=15.91 //y=2.08 //x2=16.765 //y2=2.96
cc_2261 ( N_noxref_5_c_2320_n N_noxref_23_c_7579_n ) capacitor c=0.00400249f \
 //x=15.91 //y=2.08 //x2=16.65 //y2=4.535
cc_2262 ( N_noxref_5_c_2372_n N_noxref_23_c_7579_n ) capacitor c=0.00417994f \
 //x=15.91 //y=4.7 //x2=16.65 //y2=4.535
cc_2263 ( N_noxref_5_c_2317_n N_noxref_23_c_7515_n ) capacitor c=0.00318578f \
 //x=15.795 //y=3.7 //x2=16.65 //y2=2.08
cc_2264 ( N_noxref_5_c_2320_n N_noxref_23_c_7515_n ) capacitor c=0.0776595f \
 //x=15.91 //y=2.08 //x2=16.65 //y2=2.08
cc_2265 ( N_noxref_5_c_2335_n N_noxref_23_c_7515_n ) capacitor c=0.00308814f \
 //x=15.715 //y=1.915 //x2=16.65 //y2=2.08
cc_2266 ( N_noxref_5_M63_noxref_g N_noxref_23_M65_noxref_g ) capacitor \
 c=0.0104611f //x=15.81 //y=6.02 //x2=16.69 //y2=6.02
cc_2267 ( N_noxref_5_M64_noxref_g N_noxref_23_M65_noxref_g ) capacitor \
 c=0.106811f //x=16.25 //y=6.02 //x2=16.69 //y2=6.02
cc_2268 ( N_noxref_5_M64_noxref_g N_noxref_23_M66_noxref_g ) capacitor \
 c=0.0100341f //x=16.25 //y=6.02 //x2=17.13 //y2=6.02
cc_2269 ( N_noxref_5_c_2331_n N_noxref_23_c_7587_n ) capacitor c=4.86506e-19 \
 //x=15.715 //y=0.865 //x2=16.685 //y2=0.905
cc_2270 ( N_noxref_5_c_2333_n N_noxref_23_c_7587_n ) capacitor c=0.00152104f \
 //x=15.715 //y=1.21 //x2=16.685 //y2=0.905
cc_2271 ( N_noxref_5_c_2338_n N_noxref_23_c_7587_n ) capacitor c=0.0151475f \
 //x=16.245 //y=0.865 //x2=16.685 //y2=0.905
cc_2272 ( N_noxref_5_c_2334_n N_noxref_23_c_7590_n ) capacitor c=0.00109982f \
 //x=15.715 //y=1.52 //x2=16.685 //y2=1.25
cc_2273 ( N_noxref_5_c_2340_n N_noxref_23_c_7590_n ) capacitor c=0.0111064f \
 //x=16.245 //y=1.21 //x2=16.685 //y2=1.25
cc_2274 ( N_noxref_5_c_2334_n N_noxref_23_c_7592_n ) capacitor c=9.57794e-19 \
 //x=15.715 //y=1.52 //x2=16.685 //y2=1.56
cc_2275 ( N_noxref_5_c_2335_n N_noxref_23_c_7592_n ) capacitor c=0.00662747f \
 //x=15.715 //y=1.915 //x2=16.685 //y2=1.56
cc_2276 ( N_noxref_5_c_2340_n N_noxref_23_c_7592_n ) capacitor c=0.00862358f \
 //x=16.245 //y=1.21 //x2=16.685 //y2=1.56
cc_2277 ( N_noxref_5_c_2338_n N_noxref_23_c_7595_n ) capacitor c=0.00124821f \
 //x=16.245 //y=0.865 //x2=17.215 //y2=0.905
cc_2278 ( N_noxref_5_c_2340_n N_noxref_23_c_7596_n ) capacitor c=0.00200715f \
 //x=16.245 //y=1.21 //x2=17.215 //y2=1.25
cc_2279 ( N_noxref_5_c_2320_n N_noxref_23_c_7597_n ) capacitor c=0.00307062f \
 //x=15.91 //y=2.08 //x2=16.65 //y2=2.08
cc_2280 ( N_noxref_5_c_2335_n N_noxref_23_c_7597_n ) capacitor c=0.0179092f \
 //x=15.715 //y=1.915 //x2=16.65 //y2=2.08
cc_2281 ( N_noxref_5_c_2320_n N_noxref_23_c_7599_n ) capacitor c=0.00344981f \
 //x=15.91 //y=2.08 //x2=16.68 //y2=4.7
cc_2282 ( N_noxref_5_c_2372_n N_noxref_23_c_7599_n ) capacitor c=0.0293367f \
 //x=15.91 //y=4.7 //x2=16.68 //y2=4.7
cc_2283 ( N_noxref_5_M2_noxref_d N_noxref_26_M0_noxref_s ) capacitor \
 c=0.00309936f //x=3.395 //y=0.915 //x2=0.455 //y2=0.375
cc_2284 ( N_noxref_5_c_2318_n N_noxref_27_c_8266_n ) capacitor c=0.00466084f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_2285 ( N_noxref_5_M2_noxref_d N_noxref_27_c_8266_n ) capacitor c=0.0117786f \
 //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_2286 ( N_noxref_5_c_2402_n N_noxref_27_c_8280_n ) capacitor c=0.020048f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_2287 ( N_noxref_5_M2_noxref_d N_noxref_27_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_2288 ( N_noxref_5_c_2318_n N_noxref_27_M2_noxref_s ) capacitor c=0.0207678f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_2289 ( N_noxref_5_M2_noxref_d N_noxref_27_M2_noxref_s ) capacitor \
 c=0.0426444f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
cc_2290 ( N_noxref_5_c_2318_n N_noxref_28_c_8333_n ) capacitor c=3.04182e-19 \
 //x=3.985 //y=1.665 //x2=5.505 //y2=1.495
cc_2291 ( N_noxref_5_c_2325_n N_noxref_28_c_8333_n ) capacitor c=0.0034165f \
 //x=5.725 //y=1.915 //x2=5.505 //y2=1.495
cc_2292 ( N_noxref_5_c_2319_n N_noxref_28_c_8314_n ) capacitor c=0.0116993f \
 //x=5.92 //y=2.08 //x2=6.39 //y2=1.58
cc_2293 ( N_noxref_5_c_2324_n N_noxref_28_c_8314_n ) capacitor c=0.00703567f \
 //x=5.725 //y=1.52 //x2=6.39 //y2=1.58
cc_2294 ( N_noxref_5_c_2325_n N_noxref_28_c_8314_n ) capacitor c=0.0203514f \
 //x=5.725 //y=1.915 //x2=6.39 //y2=1.58
cc_2295 ( N_noxref_5_c_2327_n N_noxref_28_c_8314_n ) capacitor c=0.00780629f \
 //x=6.1 //y=1.365 //x2=6.39 //y2=1.58
cc_2296 ( N_noxref_5_c_2330_n N_noxref_28_c_8314_n ) capacitor c=0.00339872f \
 //x=6.255 //y=1.21 //x2=6.39 //y2=1.58
cc_2297 ( N_noxref_5_c_2325_n N_noxref_28_c_8321_n ) capacitor c=6.71402e-19 \
 //x=5.725 //y=1.915 //x2=6.475 //y2=1.495
cc_2298 ( N_noxref_5_c_2321_n N_noxref_28_M3_noxref_s ) capacitor c=0.0327502f \
 //x=5.725 //y=0.865 //x2=5.37 //y2=0.365
cc_2299 ( N_noxref_5_c_2324_n N_noxref_28_M3_noxref_s ) capacitor \
 c=3.48408e-19 //x=5.725 //y=1.52 //x2=5.37 //y2=0.365
cc_2300 ( N_noxref_5_c_2328_n N_noxref_28_M3_noxref_s ) capacitor c=0.0120759f \
 //x=6.255 //y=0.865 //x2=5.37 //y2=0.365
cc_2301 ( N_noxref_5_c_2335_n N_noxref_31_c_8491_n ) capacitor c=0.0034165f \
 //x=15.715 //y=1.915 //x2=15.495 //y2=1.495
cc_2302 ( N_noxref_5_c_2320_n N_noxref_31_c_8472_n ) capacitor c=0.011424f \
 //x=15.91 //y=2.08 //x2=16.38 //y2=1.58
cc_2303 ( N_noxref_5_c_2334_n N_noxref_31_c_8472_n ) capacitor c=0.00703567f \
 //x=15.715 //y=1.52 //x2=16.38 //y2=1.58
cc_2304 ( N_noxref_5_c_2335_n N_noxref_31_c_8472_n ) capacitor c=0.018562f \
 //x=15.715 //y=1.915 //x2=16.38 //y2=1.58
cc_2305 ( N_noxref_5_c_2337_n N_noxref_31_c_8472_n ) capacitor c=0.00780629f \
 //x=16.09 //y=1.365 //x2=16.38 //y2=1.58
cc_2306 ( N_noxref_5_c_2340_n N_noxref_31_c_8472_n ) capacitor c=0.00339872f \
 //x=16.245 //y=1.21 //x2=16.38 //y2=1.58
cc_2307 ( N_noxref_5_c_2335_n N_noxref_31_c_8479_n ) capacitor c=6.71402e-19 \
 //x=15.715 //y=1.915 //x2=16.465 //y2=1.495
cc_2308 ( N_noxref_5_c_2331_n N_noxref_31_M9_noxref_s ) capacitor c=0.0326577f \
 //x=15.715 //y=0.865 //x2=15.36 //y2=0.365
cc_2309 ( N_noxref_5_c_2334_n N_noxref_31_M9_noxref_s ) capacitor \
 c=3.48408e-19 //x=15.715 //y=1.52 //x2=15.36 //y2=0.365
cc_2310 ( N_noxref_5_c_2338_n N_noxref_31_M9_noxref_s ) capacitor c=0.0120759f \
 //x=16.245 //y=0.865 //x2=15.36 //y2=0.365
cc_2311 ( N_noxref_6_c_2619_p N_noxref_7_c_2745_n ) capacitor c=0.176046f \
 //x=19.125 //y=3.7 //x2=19.865 //y2=4.07
cc_2312 ( N_noxref_6_c_2612_n N_noxref_7_c_2745_n ) capacitor c=0.0293656f \
 //x=17.505 //y=3.7 //x2=19.865 //y2=4.07
cc_2313 ( N_noxref_6_c_2566_n N_noxref_7_c_2745_n ) capacitor c=0.0200089f \
 //x=17.39 //y=3.7 //x2=19.865 //y2=4.07
cc_2314 ( N_noxref_6_c_2567_n N_noxref_7_c_2745_n ) capacitor c=0.0216244f \
 //x=19.24 //y=2.08 //x2=19.865 //y2=4.07
cc_2315 ( N_noxref_6_c_2566_n N_noxref_7_c_2721_n ) capacitor c=3.49822e-19 \
 //x=17.39 //y=3.7 //x2=14.06 //y2=4.07
cc_2316 ( N_noxref_6_c_2567_n N_noxref_7_c_2888_n ) capacitor c=0.00400249f \
 //x=19.24 //y=2.08 //x2=19.98 //y2=4.535
cc_2317 ( N_noxref_6_c_2600_n N_noxref_7_c_2888_n ) capacitor c=0.00417994f \
 //x=19.24 //y=4.7 //x2=19.98 //y2=4.535
cc_2318 ( N_noxref_6_c_2619_p N_noxref_7_c_2722_n ) capacitor c=0.00720056f \
 //x=19.125 //y=3.7 //x2=19.98 //y2=2.08
cc_2319 ( N_noxref_6_c_2566_n N_noxref_7_c_2722_n ) capacitor c=0.00107361f \
 //x=17.39 //y=3.7 //x2=19.98 //y2=2.08
cc_2320 ( N_noxref_6_c_2567_n N_noxref_7_c_2722_n ) capacitor c=0.0761047f \
 //x=19.24 //y=2.08 //x2=19.98 //y2=2.08
cc_2321 ( N_noxref_6_c_2572_n N_noxref_7_c_2722_n ) capacitor c=0.00308814f \
 //x=19.045 //y=1.915 //x2=19.98 //y2=2.08
cc_2322 ( N_noxref_6_M67_noxref_g N_noxref_7_M69_noxref_g ) capacitor \
 c=0.0104611f //x=19.14 //y=6.02 //x2=20.02 //y2=6.02
cc_2323 ( N_noxref_6_M68_noxref_g N_noxref_7_M69_noxref_g ) capacitor \
 c=0.106811f //x=19.58 //y=6.02 //x2=20.02 //y2=6.02
cc_2324 ( N_noxref_6_M68_noxref_g N_noxref_7_M70_noxref_g ) capacitor \
 c=0.0100341f //x=19.58 //y=6.02 //x2=20.46 //y2=6.02
cc_2325 ( N_noxref_6_c_2568_n N_noxref_7_c_2897_n ) capacitor c=4.86506e-19 \
 //x=19.045 //y=0.865 //x2=20.015 //y2=0.905
cc_2326 ( N_noxref_6_c_2570_n N_noxref_7_c_2897_n ) capacitor c=0.00152104f \
 //x=19.045 //y=1.21 //x2=20.015 //y2=0.905
cc_2327 ( N_noxref_6_c_2575_n N_noxref_7_c_2897_n ) capacitor c=0.0151475f \
 //x=19.575 //y=0.865 //x2=20.015 //y2=0.905
cc_2328 ( N_noxref_6_c_2571_n N_noxref_7_c_2900_n ) capacitor c=0.00109982f \
 //x=19.045 //y=1.52 //x2=20.015 //y2=1.25
cc_2329 ( N_noxref_6_c_2577_n N_noxref_7_c_2900_n ) capacitor c=0.0111064f \
 //x=19.575 //y=1.21 //x2=20.015 //y2=1.25
cc_2330 ( N_noxref_6_c_2571_n N_noxref_7_c_2902_n ) capacitor c=9.57794e-19 \
 //x=19.045 //y=1.52 //x2=20.015 //y2=1.56
cc_2331 ( N_noxref_6_c_2572_n N_noxref_7_c_2902_n ) capacitor c=0.00662747f \
 //x=19.045 //y=1.915 //x2=20.015 //y2=1.56
cc_2332 ( N_noxref_6_c_2577_n N_noxref_7_c_2902_n ) capacitor c=0.00862358f \
 //x=19.575 //y=1.21 //x2=20.015 //y2=1.56
cc_2333 ( N_noxref_6_c_2575_n N_noxref_7_c_2905_n ) capacitor c=0.00124821f \
 //x=19.575 //y=0.865 //x2=20.545 //y2=0.905
cc_2334 ( N_noxref_6_c_2577_n N_noxref_7_c_2906_n ) capacitor c=0.00200715f \
 //x=19.575 //y=1.21 //x2=20.545 //y2=1.25
cc_2335 ( N_noxref_6_c_2567_n N_noxref_7_c_2907_n ) capacitor c=0.00307062f \
 //x=19.24 //y=2.08 //x2=19.98 //y2=2.08
cc_2336 ( N_noxref_6_c_2572_n N_noxref_7_c_2907_n ) capacitor c=0.0179092f \
 //x=19.045 //y=1.915 //x2=19.98 //y2=2.08
cc_2337 ( N_noxref_6_c_2567_n N_noxref_7_c_2909_n ) capacitor c=0.00344981f \
 //x=19.24 //y=2.08 //x2=20.01 //y2=4.7
cc_2338 ( N_noxref_6_c_2600_n N_noxref_7_c_2909_n ) capacitor c=0.0293367f \
 //x=19.24 //y=4.7 //x2=20.01 //y2=4.7
cc_2339 ( N_noxref_6_c_2619_p N_D_c_4217_n ) capacitor c=0.00669561f \
 //x=19.125 //y=3.7 //x2=28.005 //y2=2.59
cc_2340 ( N_noxref_6_c_2612_n N_D_c_4217_n ) capacitor c=6.305e-19 //x=17.505 \
 //y=3.7 //x2=28.005 //y2=2.59
cc_2341 ( N_noxref_6_c_2649_p N_D_c_4217_n ) capacitor c=0.0102711f //x=17.035 \
 //y=1.655 //x2=28.005 //y2=2.59
cc_2342 ( N_noxref_6_c_2566_n N_D_c_4217_n ) capacitor c=0.0210598f //x=17.39 \
 //y=3.7 //x2=28.005 //y2=2.59
cc_2343 ( N_noxref_6_c_2567_n N_D_c_4217_n ) capacitor c=0.0213243f //x=19.24 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2344 ( N_noxref_6_c_2572_n N_D_c_4217_n ) capacitor c=0.0052136f //x=19.045 \
 //y=1.915 //x2=28.005 //y2=2.59
cc_2345 ( N_noxref_6_c_2581_n N_CLK_c_5053_n ) capacitor c=0.00115095f \
 //x=16.825 //y=5.2 //x2=16.745 //y2=4.442
cc_2346 ( N_noxref_6_c_2585_n N_CLK_c_5053_n ) capacitor c=0.0179906f \
 //x=16.115 //y=5.2 //x2=16.745 //y2=4.442
cc_2347 ( N_noxref_6_c_2619_p N_CLK_c_5079_n ) capacitor c=0.0104236f \
 //x=19.125 //y=3.7 //x2=23.795 //y2=4.44
cc_2348 ( N_noxref_6_c_2612_n N_CLK_c_5079_n ) capacitor c=8.86008e-19 \
 //x=17.505 //y=3.7 //x2=23.795 //y2=4.44
cc_2349 ( N_noxref_6_c_2581_n N_CLK_c_5079_n ) capacitor c=0.0173718f \
 //x=16.825 //y=5.2 //x2=23.795 //y2=4.44
cc_2350 ( N_noxref_6_c_2566_n N_CLK_c_5079_n ) capacitor c=0.0208251f \
 //x=17.39 //y=3.7 //x2=23.795 //y2=4.44
cc_2351 ( N_noxref_6_c_2567_n N_CLK_c_5079_n ) capacitor c=0.0198304f \
 //x=19.24 //y=2.08 //x2=23.795 //y2=4.44
cc_2352 ( N_noxref_6_c_2600_n N_CLK_c_5079_n ) capacitor c=0.0107057f \
 //x=19.24 //y=4.7 //x2=23.795 //y2=4.44
cc_2353 ( N_noxref_6_c_2619_p N_noxref_23_c_7497_n ) capacitor c=0.0868505f \
 //x=19.125 //y=3.7 //x2=20.605 //y2=2.96
cc_2354 ( N_noxref_6_c_2612_n N_noxref_23_c_7497_n ) capacitor c=0.0133597f \
 //x=17.505 //y=3.7 //x2=20.605 //y2=2.96
cc_2355 ( N_noxref_6_c_2566_n N_noxref_23_c_7497_n ) capacitor c=0.0214247f \
 //x=17.39 //y=3.7 //x2=20.605 //y2=2.96
cc_2356 ( N_noxref_6_c_2567_n N_noxref_23_c_7497_n ) capacitor c=0.0213728f \
 //x=19.24 //y=2.08 //x2=20.605 //y2=2.96
cc_2357 ( N_noxref_6_c_2566_n N_noxref_23_c_7578_n ) capacitor c=0.00117715f \
 //x=17.39 //y=3.7 //x2=16.765 //y2=2.96
cc_2358 ( N_noxref_6_c_2581_n N_noxref_23_c_7579_n ) capacitor c=0.0127216f \
 //x=16.825 //y=5.2 //x2=16.65 //y2=4.535
cc_2359 ( N_noxref_6_c_2566_n N_noxref_23_c_7579_n ) capacitor c=0.0101284f \
 //x=17.39 //y=3.7 //x2=16.65 //y2=4.535
cc_2360 ( N_noxref_6_c_2612_n N_noxref_23_c_7515_n ) capacitor c=0.00329059f \
 //x=17.505 //y=3.7 //x2=16.65 //y2=2.08
cc_2361 ( N_noxref_6_c_2566_n N_noxref_23_c_7515_n ) capacitor c=0.071705f \
 //x=17.39 //y=3.7 //x2=16.65 //y2=2.08
cc_2362 ( N_noxref_6_c_2567_n N_noxref_23_c_7515_n ) capacitor c=0.001003f \
 //x=19.24 //y=2.08 //x2=16.65 //y2=2.08
cc_2363 ( N_noxref_6_M68_noxref_g N_noxref_23_c_7540_n ) capacitor \
 c=0.0169521f //x=19.58 //y=6.02 //x2=20.155 //y2=5.2
cc_2364 ( N_noxref_6_c_2567_n N_noxref_23_c_7544_n ) capacitor c=0.00521572f \
 //x=19.24 //y=2.08 //x2=19.445 //y2=5.2
cc_2365 ( N_noxref_6_M67_noxref_g N_noxref_23_c_7544_n ) capacitor \
 c=0.0177326f //x=19.14 //y=6.02 //x2=19.445 //y2=5.2
cc_2366 ( N_noxref_6_c_2600_n N_noxref_23_c_7544_n ) capacitor c=0.00581252f \
 //x=19.24 //y=4.7 //x2=19.445 //y2=5.2
cc_2367 ( N_noxref_6_c_2566_n N_noxref_23_c_7518_n ) capacitor c=3.49822e-19 \
 //x=17.39 //y=3.7 //x2=20.72 //y2=2.96
cc_2368 ( N_noxref_6_c_2567_n N_noxref_23_c_7518_n ) capacitor c=0.00365805f \
 //x=19.24 //y=2.08 //x2=20.72 //y2=2.96
cc_2369 ( N_noxref_6_c_2581_n N_noxref_23_M65_noxref_g ) capacitor \
 c=0.0166421f //x=16.825 //y=5.2 //x2=16.69 //y2=6.02
cc_2370 ( N_noxref_6_M65_noxref_d N_noxref_23_M65_noxref_g ) capacitor \
 c=0.0173476f //x=16.765 //y=5.02 //x2=16.69 //y2=6.02
cc_2371 ( N_noxref_6_c_2587_n N_noxref_23_M66_noxref_g ) capacitor c=0.018922f \
 //x=17.305 //y=5.2 //x2=17.13 //y2=6.02
cc_2372 ( N_noxref_6_M65_noxref_d N_noxref_23_M66_noxref_g ) capacitor \
 c=0.0179769f //x=16.765 //y=5.02 //x2=17.13 //y2=6.02
cc_2373 ( N_noxref_6_M10_noxref_d N_noxref_23_c_7587_n ) capacitor \
 c=0.00217566f //x=16.76 //y=0.905 //x2=16.685 //y2=0.905
cc_2374 ( N_noxref_6_M10_noxref_d N_noxref_23_c_7590_n ) capacitor \
 c=0.0034598f //x=16.76 //y=0.905 //x2=16.685 //y2=1.25
cc_2375 ( N_noxref_6_M10_noxref_d N_noxref_23_c_7592_n ) capacitor \
 c=0.00656319f //x=16.76 //y=0.905 //x2=16.685 //y2=1.56
cc_2376 ( N_noxref_6_c_2566_n N_noxref_23_c_7624_n ) capacitor c=0.0142673f \
 //x=17.39 //y=3.7 //x2=17.055 //y2=4.79
cc_2377 ( N_noxref_6_c_2685_p N_noxref_23_c_7624_n ) capacitor c=0.00407665f \
 //x=16.91 //y=5.2 //x2=17.055 //y2=4.79
cc_2378 ( N_noxref_6_M10_noxref_d N_noxref_23_c_7626_n ) capacitor \
 c=0.00241102f //x=16.76 //y=0.905 //x2=17.06 //y2=0.75
cc_2379 ( N_noxref_6_c_2565_n N_noxref_23_c_7627_n ) capacitor c=0.00359704f \
 //x=17.305 //y=1.655 //x2=17.06 //y2=1.405
cc_2380 ( N_noxref_6_M10_noxref_d N_noxref_23_c_7627_n ) capacitor \
 c=0.0138845f //x=16.76 //y=0.905 //x2=17.06 //y2=1.405
cc_2381 ( N_noxref_6_M10_noxref_d N_noxref_23_c_7595_n ) capacitor \
 c=0.00132245f //x=16.76 //y=0.905 //x2=17.215 //y2=0.905
cc_2382 ( N_noxref_6_c_2565_n N_noxref_23_c_7596_n ) capacitor c=0.00457401f \
 //x=17.305 //y=1.655 //x2=17.215 //y2=1.25
cc_2383 ( N_noxref_6_M10_noxref_d N_noxref_23_c_7596_n ) capacitor \
 c=0.00566463f //x=16.76 //y=0.905 //x2=17.215 //y2=1.25
cc_2384 ( N_noxref_6_c_2566_n N_noxref_23_c_7597_n ) capacitor c=0.00877984f \
 //x=17.39 //y=3.7 //x2=16.65 //y2=2.08
cc_2385 ( N_noxref_6_c_2566_n N_noxref_23_c_7633_n ) capacitor c=0.00306024f \
 //x=17.39 //y=3.7 //x2=16.65 //y2=1.915
cc_2386 ( N_noxref_6_M10_noxref_d N_noxref_23_c_7633_n ) capacitor \
 c=0.00660593f //x=16.76 //y=0.905 //x2=16.65 //y2=1.915
cc_2387 ( N_noxref_6_c_2581_n N_noxref_23_c_7599_n ) capacitor c=0.00346528f \
 //x=16.825 //y=5.2 //x2=16.68 //y2=4.7
cc_2388 ( N_noxref_6_c_2566_n N_noxref_23_c_7599_n ) capacitor c=0.00533692f \
 //x=17.39 //y=3.7 //x2=16.68 //y2=4.7
cc_2389 ( N_noxref_6_M68_noxref_g N_noxref_23_M67_noxref_d ) capacitor \
 c=0.0173476f //x=19.58 //y=6.02 //x2=19.215 //y2=5.02
cc_2390 ( N_noxref_6_c_2649_p N_noxref_31_c_8491_n ) capacitor c=3.15806e-19 \
 //x=17.035 //y=1.655 //x2=15.495 //y2=1.495
cc_2391 ( N_noxref_6_c_2649_p N_noxref_31_c_8479_n ) capacitor c=0.0203424f \
 //x=17.035 //y=1.655 //x2=16.465 //y2=1.495
cc_2392 ( N_noxref_6_c_2565_n N_noxref_31_c_8480_n ) capacitor c=0.00461444f \
 //x=17.305 //y=1.655 //x2=17.35 //y2=0.53
cc_2393 ( N_noxref_6_M10_noxref_d N_noxref_31_c_8480_n ) capacitor \
 c=0.0116735f //x=16.76 //y=0.905 //x2=17.35 //y2=0.53
cc_2394 ( N_noxref_6_c_2565_n N_noxref_31_M9_noxref_s ) capacitor c=0.0137901f \
 //x=17.305 //y=1.655 //x2=15.36 //y2=0.365
cc_2395 ( N_noxref_6_M10_noxref_d N_noxref_31_M9_noxref_s ) capacitor \
 c=0.043966f //x=16.76 //y=0.905 //x2=15.36 //y2=0.365
cc_2396 ( N_noxref_6_c_2565_n N_noxref_32_c_8543_n ) capacitor c=3.22188e-19 \
 //x=17.305 //y=1.655 //x2=18.825 //y2=1.495
cc_2397 ( N_noxref_6_c_2572_n N_noxref_32_c_8543_n ) capacitor c=0.0034165f \
 //x=19.045 //y=1.915 //x2=18.825 //y2=1.495
cc_2398 ( N_noxref_6_c_2567_n N_noxref_32_c_8524_n ) capacitor c=0.0118762f \
 //x=19.24 //y=2.08 //x2=19.71 //y2=1.58
cc_2399 ( N_noxref_6_c_2571_n N_noxref_32_c_8524_n ) capacitor c=0.00703567f \
 //x=19.045 //y=1.52 //x2=19.71 //y2=1.58
cc_2400 ( N_noxref_6_c_2572_n N_noxref_32_c_8524_n ) capacitor c=0.018562f \
 //x=19.045 //y=1.915 //x2=19.71 //y2=1.58
cc_2401 ( N_noxref_6_c_2574_n N_noxref_32_c_8524_n ) capacitor c=0.00780629f \
 //x=19.42 //y=1.365 //x2=19.71 //y2=1.58
cc_2402 ( N_noxref_6_c_2577_n N_noxref_32_c_8524_n ) capacitor c=0.00339872f \
 //x=19.575 //y=1.21 //x2=19.71 //y2=1.58
cc_2403 ( N_noxref_6_c_2572_n N_noxref_32_c_8531_n ) capacitor c=6.71402e-19 \
 //x=19.045 //y=1.915 //x2=19.795 //y2=1.495
cc_2404 ( N_noxref_6_c_2568_n N_noxref_32_M11_noxref_s ) capacitor \
 c=0.0326577f //x=19.045 //y=0.865 //x2=18.69 //y2=0.365
cc_2405 ( N_noxref_6_c_2571_n N_noxref_32_M11_noxref_s ) capacitor \
 c=3.48408e-19 //x=19.045 //y=1.52 //x2=18.69 //y2=0.365
cc_2406 ( N_noxref_6_c_2575_n N_noxref_32_M11_noxref_s ) capacitor \
 c=0.0120759f //x=19.575 //y=0.865 //x2=18.69 //y2=0.365
cc_2407 ( N_noxref_7_c_2745_n N_noxref_12_c_3884_n ) capacitor c=0.00649178f \
 //x=19.865 //y=4.07 //x2=22.685 //y2=4.07
cc_2408 ( N_noxref_7_c_2722_n N_noxref_12_c_3862_n ) capacitor c=9.69916e-19 \
 //x=19.98 //y=2.08 //x2=22.57 //y2=2.08
cc_2409 ( N_noxref_7_c_2715_n N_D_c_4217_n ) capacitor c=0.00334753f //x=9.875 \
 //y=4.07 //x2=28.005 //y2=2.59
cc_2410 ( N_noxref_7_c_2744_n N_D_c_4217_n ) capacitor c=0.00994417f \
 //x=13.945 //y=4.07 //x2=28.005 //y2=2.59
cc_2411 ( N_noxref_7_c_2801_n N_D_c_4217_n ) capacitor c=3.04562e-19 \
 //x=10.105 //y=4.07 //x2=28.005 //y2=2.59
cc_2412 ( N_noxref_7_c_2745_n N_D_c_4217_n ) capacitor c=0.0235271f //x=19.865 \
 //y=4.07 //x2=28.005 //y2=2.59
cc_2413 ( N_noxref_7_c_2747_n N_D_c_4217_n ) capacitor c=4.12718e-19 \
 //x=14.175 //y=4.07 //x2=28.005 //y2=2.59
cc_2414 ( N_noxref_7_c_2718_n N_D_c_4217_n ) capacitor c=0.024321f //x=9.99 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2415 ( N_noxref_7_c_2919_p N_D_c_4217_n ) capacitor c=0.0102711f //x=13.705 \
 //y=1.655 //x2=28.005 //y2=2.59
cc_2416 ( N_noxref_7_c_2721_n N_D_c_4217_n ) capacitor c=0.0249199f //x=14.06 \
 //y=4.07 //x2=28.005 //y2=2.59
cc_2417 ( N_noxref_7_c_2722_n N_D_c_4217_n ) capacitor c=0.0204615f //x=19.98 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2418 ( N_noxref_7_c_2822_n N_D_c_4217_n ) capacitor c=0.00217166f //x=9.99 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2419 ( N_noxref_7_c_2907_n N_D_c_4217_n ) capacitor c=0.00219932f //x=19.98 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2420 ( N_noxref_7_c_2715_n N_D_c_4253_n ) capacitor c=0.0169317f //x=9.875 \
 //y=4.07 //x2=6.66 //y2=2.08
cc_2421 ( N_noxref_7_c_2715_n N_CLK_c_5034_n ) capacitor c=0.656956f //x=9.875 \
 //y=4.07 //x2=13.205 //y2=4.44
cc_2422 ( N_noxref_7_c_2744_n N_CLK_c_5034_n ) capacitor c=0.270915f \
 //x=13.945 //y=4.07 //x2=13.205 //y2=4.44
cc_2423 ( N_noxref_7_c_2801_n N_CLK_c_5034_n ) capacitor c=0.0263375f \
 //x=10.105 //y=4.07 //x2=13.205 //y2=4.44
cc_2424 ( N_noxref_7_c_2803_n N_CLK_c_5034_n ) capacitor c=0.0016972f //x=9.99 \
 //y=4.535 //x2=13.205 //y2=4.44
cc_2425 ( N_noxref_7_c_2718_n N_CLK_c_5034_n ) capacitor c=0.0207534f //x=9.99 \
 //y=2.08 //x2=13.205 //y2=4.44
cc_2426 ( N_noxref_7_c_2757_n N_CLK_c_5034_n ) capacitor c=0.0172877f \
 //x=12.785 //y=5.2 //x2=13.205 //y2=4.44
cc_2427 ( N_noxref_7_c_2849_n N_CLK_c_5034_n ) capacitor c=0.00960248f \
 //x=10.395 //y=4.79 //x2=13.205 //y2=4.44
cc_2428 ( N_noxref_7_c_2824_n N_CLK_c_5034_n ) capacitor c=0.00203982f \
 //x=10.02 //y=4.7 //x2=13.205 //y2=4.44
cc_2429 ( N_noxref_7_c_2715_n N_CLK_c_5052_n ) capacitor c=0.0291328f \
 //x=9.875 //y=4.07 //x2=2.335 //y2=4.44
cc_2430 ( N_noxref_7_c_2717_n N_CLK_c_5052_n ) capacitor c=0.00551083f \
 //x=1.11 //y=2.08 //x2=2.335 //y2=4.44
cc_2431 ( N_noxref_7_c_2744_n N_CLK_c_5053_n ) capacitor c=0.0406398f \
 //x=13.945 //y=4.07 //x2=16.745 //y2=4.442
cc_2432 ( N_noxref_7_c_2745_n N_CLK_c_5053_n ) capacitor c=0.218547f \
 //x=19.865 //y=4.07 //x2=16.745 //y2=4.442
cc_2433 ( N_noxref_7_c_2747_n N_CLK_c_5053_n ) capacitor c=0.0258275f \
 //x=14.175 //y=4.07 //x2=16.745 //y2=4.442
cc_2434 ( N_noxref_7_c_2753_n N_CLK_c_5053_n ) capacitor c=0.0163436f \
 //x=13.495 //y=5.2 //x2=16.745 //y2=4.442
cc_2435 ( N_noxref_7_c_2721_n N_CLK_c_5053_n ) capacitor c=0.0216361f \
 //x=14.06 //y=4.07 //x2=16.745 //y2=4.442
cc_2436 ( N_noxref_7_c_2744_n N_CLK_c_5060_n ) capacitor c=0.0293862f \
 //x=13.945 //y=4.07 //x2=13.465 //y2=4.442
cc_2437 ( N_noxref_7_c_2753_n N_CLK_c_5060_n ) capacitor c=0.00325337f \
 //x=13.495 //y=5.2 //x2=13.465 //y2=4.442
cc_2438 ( N_noxref_7_c_2721_n N_CLK_c_5060_n ) capacitor c=0.00183349f \
 //x=14.06 //y=4.07 //x2=13.465 //y2=4.442
cc_2439 ( N_noxref_7_c_2745_n N_CLK_c_5079_n ) capacitor c=0.301708f \
 //x=19.865 //y=4.07 //x2=23.795 //y2=4.44
cc_2440 ( N_noxref_7_c_2888_n N_CLK_c_5079_n ) capacitor c=0.0016972f \
 //x=19.98 //y=4.535 //x2=23.795 //y2=4.44
cc_2441 ( N_noxref_7_c_2722_n N_CLK_c_5079_n ) capacitor c=0.0207534f \
 //x=19.98 //y=2.08 //x2=23.795 //y2=4.44
cc_2442 ( N_noxref_7_c_2946_p N_CLK_c_5079_n ) capacitor c=0.00720343f \
 //x=20.385 //y=4.79 //x2=23.795 //y2=4.44
cc_2443 ( N_noxref_7_c_2909_n N_CLK_c_5079_n ) capacitor c=0.0019199f \
 //x=20.01 //y=4.7 //x2=23.795 //y2=4.44
cc_2444 ( N_noxref_7_c_2715_n N_CLK_c_5025_n ) capacitor c=0.0265867f \
 //x=9.875 //y=4.07 //x2=2.22 //y2=2.08
cc_2445 ( N_noxref_7_c_2716_n N_CLK_c_5025_n ) capacitor c=0.00128547f \
 //x=1.225 //y=4.07 //x2=2.22 //y2=2.08
cc_2446 ( N_noxref_7_c_2717_n N_CLK_c_5025_n ) capacitor c=0.0535714f //x=1.11 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_2447 ( N_noxref_7_c_2728_n N_CLK_c_5025_n ) capacitor c=0.00238338f \
 //x=0.81 //y=1.915 //x2=2.22 //y2=2.08
cc_2448 ( N_noxref_7_c_2882_n N_CLK_c_5025_n ) capacitor c=0.00147352f \
 //x=1.675 //y=4.79 //x2=2.22 //y2=2.08
cc_2449 ( N_noxref_7_c_2781_n N_CLK_c_5025_n ) capacitor c=0.00141297f \
 //x=1.385 //y=4.79 //x2=2.22 //y2=2.08
cc_2450 ( N_noxref_7_c_2753_n N_CLK_c_5203_n ) capacitor c=0.0126974f \
 //x=13.495 //y=5.2 //x2=13.32 //y2=4.535
cc_2451 ( N_noxref_7_c_2721_n N_CLK_c_5203_n ) capacitor c=0.00923416f \
 //x=14.06 //y=4.07 //x2=13.32 //y2=4.535
cc_2452 ( N_noxref_7_c_2744_n N_CLK_c_5026_n ) capacitor c=0.0187718f \
 //x=13.945 //y=4.07 //x2=13.32 //y2=2.08
cc_2453 ( N_noxref_7_c_2747_n N_CLK_c_5026_n ) capacitor c=0.00117715f \
 //x=14.175 //y=4.07 //x2=13.32 //y2=2.08
cc_2454 ( N_noxref_7_c_2753_n N_CLK_c_5026_n ) capacitor c=3.74769e-19 \
 //x=13.495 //y=5.2 //x2=13.32 //y2=2.08
cc_2455 ( N_noxref_7_c_2721_n N_CLK_c_5026_n ) capacitor c=0.0723779f \
 //x=14.06 //y=4.07 //x2=13.32 //y2=2.08
cc_2456 ( N_noxref_7_M45_noxref_g N_CLK_M47_noxref_g ) capacitor c=0.0105869f \
 //x=1.31 //y=6.02 //x2=2.19 //y2=6.02
cc_2457 ( N_noxref_7_M46_noxref_g N_CLK_M47_noxref_g ) capacitor c=0.10632f \
 //x=1.75 //y=6.02 //x2=2.19 //y2=6.02
cc_2458 ( N_noxref_7_M46_noxref_g N_CLK_M48_noxref_g ) capacitor c=0.0101598f \
 //x=1.75 //y=6.02 //x2=2.63 //y2=6.02
cc_2459 ( N_noxref_7_c_2753_n N_CLK_M61_noxref_g ) capacitor c=0.0166421f \
 //x=13.495 //y=5.2 //x2=13.36 //y2=6.02
cc_2460 ( N_noxref_7_M61_noxref_d N_CLK_M61_noxref_g ) capacitor c=0.0173476f \
 //x=13.435 //y=5.02 //x2=13.36 //y2=6.02
cc_2461 ( N_noxref_7_c_2759_n N_CLK_M62_noxref_g ) capacitor c=0.0189374f \
 //x=13.975 //y=5.2 //x2=13.8 //y2=6.02
cc_2462 ( N_noxref_7_M61_noxref_d N_CLK_M62_noxref_g ) capacitor c=0.0179769f \
 //x=13.435 //y=5.02 //x2=13.8 //y2=6.02
cc_2463 ( N_noxref_7_c_2724_n N_CLK_c_5300_n ) capacitor c=5.72482e-19 \
 //x=0.81 //y=0.875 //x2=1.785 //y2=0.91
cc_2464 ( N_noxref_7_c_2726_n N_CLK_c_5300_n ) capacitor c=0.00149976f \
 //x=0.81 //y=1.22 //x2=1.785 //y2=0.91
cc_2465 ( N_noxref_7_c_2731_n N_CLK_c_5300_n ) capacitor c=0.0160123f //x=1.34 \
 //y=0.875 //x2=1.785 //y2=0.91
cc_2466 ( N_noxref_7_c_2727_n N_CLK_c_5303_n ) capacitor c=0.00111227f \
 //x=0.81 //y=1.53 //x2=1.785 //y2=1.22
cc_2467 ( N_noxref_7_c_2733_n N_CLK_c_5303_n ) capacitor c=0.0124075f //x=1.34 \
 //y=1.22 //x2=1.785 //y2=1.22
cc_2468 ( N_noxref_7_c_2731_n N_CLK_c_5187_n ) capacitor c=0.00103227f \
 //x=1.34 //y=0.875 //x2=2.31 //y2=0.91
cc_2469 ( N_noxref_7_c_2733_n N_CLK_c_5188_n ) capacitor c=0.0010154f //x=1.34 \
 //y=1.22 //x2=2.31 //y2=1.22
cc_2470 ( N_noxref_7_c_2733_n N_CLK_c_5189_n ) capacitor c=9.23422e-19 \
 //x=1.34 //y=1.22 //x2=2.31 //y2=1.45
cc_2471 ( N_noxref_7_c_2717_n N_CLK_c_5190_n ) capacitor c=0.00231304f \
 //x=1.11 //y=2.08 //x2=2.31 //y2=1.915
cc_2472 ( N_noxref_7_c_2728_n N_CLK_c_5190_n ) capacitor c=0.00964411f \
 //x=0.81 //y=1.915 //x2=2.31 //y2=1.915
cc_2473 ( N_noxref_7_M8_noxref_d N_CLK_c_5212_n ) capacitor c=0.00217566f \
 //x=13.43 //y=0.905 //x2=13.355 //y2=0.905
cc_2474 ( N_noxref_7_M8_noxref_d N_CLK_c_5215_n ) capacitor c=0.0034598f \
 //x=13.43 //y=0.905 //x2=13.355 //y2=1.25
cc_2475 ( N_noxref_7_M8_noxref_d N_CLK_c_5217_n ) capacitor c=0.00656319f \
 //x=13.43 //y=0.905 //x2=13.355 //y2=1.56
cc_2476 ( N_noxref_7_c_2721_n N_CLK_c_5313_n ) capacitor c=0.0142673f \
 //x=14.06 //y=4.07 //x2=13.725 //y2=4.79
cc_2477 ( N_noxref_7_c_2981_p N_CLK_c_5313_n ) capacitor c=0.00407678f \
 //x=13.58 //y=5.2 //x2=13.725 //y2=4.79
cc_2478 ( N_noxref_7_M8_noxref_d N_CLK_c_5315_n ) capacitor c=0.00241102f \
 //x=13.43 //y=0.905 //x2=13.73 //y2=0.75
cc_2479 ( N_noxref_7_c_2720_n N_CLK_c_5316_n ) capacitor c=0.00359704f \
 //x=13.975 //y=1.655 //x2=13.73 //y2=1.405
cc_2480 ( N_noxref_7_M8_noxref_d N_CLK_c_5316_n ) capacitor c=0.0138845f \
 //x=13.43 //y=0.905 //x2=13.73 //y2=1.405
cc_2481 ( N_noxref_7_M8_noxref_d N_CLK_c_5220_n ) capacitor c=0.00132245f \
 //x=13.43 //y=0.905 //x2=13.885 //y2=0.905
cc_2482 ( N_noxref_7_c_2720_n N_CLK_c_5221_n ) capacitor c=0.00457401f \
 //x=13.975 //y=1.655 //x2=13.885 //y2=1.25
cc_2483 ( N_noxref_7_M8_noxref_d N_CLK_c_5221_n ) capacitor c=0.00566463f \
 //x=13.43 //y=0.905 //x2=13.885 //y2=1.25
cc_2484 ( N_noxref_7_c_2715_n N_CLK_c_5194_n ) capacitor c=6.38735e-19 \
 //x=9.875 //y=4.07 //x2=2.22 //y2=4.7
cc_2485 ( N_noxref_7_c_2717_n N_CLK_c_5194_n ) capacitor c=0.00183762f \
 //x=1.11 //y=2.08 //x2=2.22 //y2=4.7
cc_2486 ( N_noxref_7_c_2882_n N_CLK_c_5194_n ) capacitor c=0.0168581f \
 //x=1.675 //y=4.79 //x2=2.22 //y2=4.7
cc_2487 ( N_noxref_7_c_2781_n N_CLK_c_5194_n ) capacitor c=0.00484466f \
 //x=1.385 //y=4.79 //x2=2.22 //y2=4.7
cc_2488 ( N_noxref_7_c_2721_n N_CLK_c_5222_n ) capacitor c=0.00877984f \
 //x=14.06 //y=4.07 //x2=13.32 //y2=2.08
cc_2489 ( N_noxref_7_c_2721_n N_CLK_c_5326_n ) capacitor c=0.00306024f \
 //x=14.06 //y=4.07 //x2=13.32 //y2=1.915
cc_2490 ( N_noxref_7_M8_noxref_d N_CLK_c_5326_n ) capacitor c=0.00660593f \
 //x=13.43 //y=0.905 //x2=13.32 //y2=1.915
cc_2491 ( N_noxref_7_c_2753_n N_CLK_c_5224_n ) capacitor c=0.00346519f \
 //x=13.495 //y=5.2 //x2=13.35 //y2=4.7
cc_2492 ( N_noxref_7_c_2721_n N_CLK_c_5224_n ) capacitor c=0.00518077f \
 //x=14.06 //y=4.07 //x2=13.35 //y2=4.7
cc_2493 ( N_noxref_7_c_2745_n N_noxref_23_c_7497_n ) capacitor c=0.0433611f \
 //x=19.865 //y=4.07 //x2=20.605 //y2=2.96
cc_2494 ( N_noxref_7_c_2722_n N_noxref_23_c_7497_n ) capacitor c=0.0209015f \
 //x=19.98 //y=2.08 //x2=20.605 //y2=2.96
cc_2495 ( N_noxref_7_c_2745_n N_noxref_23_c_7578_n ) capacitor c=0.0076696f \
 //x=19.865 //y=4.07 //x2=16.765 //y2=2.96
cc_2496 ( N_noxref_7_c_2722_n N_noxref_23_c_7641_n ) capacitor c=0.00117715f \
 //x=19.98 //y=2.08 //x2=20.835 //y2=2.96
cc_2497 ( N_noxref_7_c_2745_n N_noxref_23_c_7515_n ) capacitor c=0.0209602f \
 //x=19.865 //y=4.07 //x2=16.65 //y2=2.08
cc_2498 ( N_noxref_7_c_2721_n N_noxref_23_c_7515_n ) capacitor c=0.00114594f \
 //x=14.06 //y=4.07 //x2=16.65 //y2=2.08
cc_2499 ( N_noxref_7_c_2888_n N_noxref_23_c_7540_n ) capacitor c=0.0127164f \
 //x=19.98 //y=4.535 //x2=20.155 //y2=5.2
cc_2500 ( N_noxref_7_M69_noxref_g N_noxref_23_c_7540_n ) capacitor \
 c=0.0166421f //x=20.02 //y=6.02 //x2=20.155 //y2=5.2
cc_2501 ( N_noxref_7_c_2909_n N_noxref_23_c_7540_n ) capacitor c=0.00346527f \
 //x=20.01 //y=4.7 //x2=20.155 //y2=5.2
cc_2502 ( N_noxref_7_M70_noxref_g N_noxref_23_c_7546_n ) capacitor c=0.018922f \
 //x=20.46 //y=6.02 //x2=20.635 //y2=5.2
cc_2503 ( N_noxref_7_c_3007_p N_noxref_23_c_7517_n ) capacitor c=0.00359704f \
 //x=20.39 //y=1.405 //x2=20.635 //y2=1.655
cc_2504 ( N_noxref_7_c_2906_n N_noxref_23_c_7517_n ) capacitor c=0.00457401f \
 //x=20.545 //y=1.25 //x2=20.635 //y2=1.655
cc_2505 ( N_noxref_7_c_2745_n N_noxref_23_c_7518_n ) capacitor c=0.00423741f \
 //x=19.865 //y=4.07 //x2=20.72 //y2=2.96
cc_2506 ( N_noxref_7_c_2888_n N_noxref_23_c_7518_n ) capacitor c=0.0101115f \
 //x=19.98 //y=4.535 //x2=20.72 //y2=2.96
cc_2507 ( N_noxref_7_c_2722_n N_noxref_23_c_7518_n ) capacitor c=0.073972f \
 //x=19.98 //y=2.08 //x2=20.72 //y2=2.96
cc_2508 ( N_noxref_7_c_2946_p N_noxref_23_c_7518_n ) capacitor c=0.0142673f \
 //x=20.385 //y=4.79 //x2=20.72 //y2=2.96
cc_2509 ( N_noxref_7_c_2907_n N_noxref_23_c_7518_n ) capacitor c=0.00877984f \
 //x=19.98 //y=2.08 //x2=20.72 //y2=2.96
cc_2510 ( N_noxref_7_c_3014_p N_noxref_23_c_7518_n ) capacitor c=0.00306024f \
 //x=19.98 //y=1.915 //x2=20.72 //y2=2.96
cc_2511 ( N_noxref_7_c_2909_n N_noxref_23_c_7518_n ) capacitor c=0.00517969f \
 //x=20.01 //y=4.7 //x2=20.72 //y2=2.96
cc_2512 ( N_noxref_7_c_2946_p N_noxref_23_c_7657_n ) capacitor c=0.00407665f \
 //x=20.385 //y=4.79 //x2=20.24 //y2=5.2
cc_2513 ( N_noxref_7_c_2897_n N_noxref_23_M12_noxref_d ) capacitor \
 c=0.00217566f //x=20.015 //y=0.905 //x2=20.09 //y2=0.905
cc_2514 ( N_noxref_7_c_2900_n N_noxref_23_M12_noxref_d ) capacitor \
 c=0.0034598f //x=20.015 //y=1.25 //x2=20.09 //y2=0.905
cc_2515 ( N_noxref_7_c_2902_n N_noxref_23_M12_noxref_d ) capacitor \
 c=0.00656319f //x=20.015 //y=1.56 //x2=20.09 //y2=0.905
cc_2516 ( N_noxref_7_c_3020_p N_noxref_23_M12_noxref_d ) capacitor \
 c=0.00241102f //x=20.39 //y=0.75 //x2=20.09 //y2=0.905
cc_2517 ( N_noxref_7_c_3007_p N_noxref_23_M12_noxref_d ) capacitor \
 c=0.0138845f //x=20.39 //y=1.405 //x2=20.09 //y2=0.905
cc_2518 ( N_noxref_7_c_2905_n N_noxref_23_M12_noxref_d ) capacitor \
 c=0.00132245f //x=20.545 //y=0.905 //x2=20.09 //y2=0.905
cc_2519 ( N_noxref_7_c_2906_n N_noxref_23_M12_noxref_d ) capacitor \
 c=0.00566463f //x=20.545 //y=1.25 //x2=20.09 //y2=0.905
cc_2520 ( N_noxref_7_c_3014_p N_noxref_23_M12_noxref_d ) capacitor \
 c=0.00660593f //x=19.98 //y=1.915 //x2=20.09 //y2=0.905
cc_2521 ( N_noxref_7_M69_noxref_g N_noxref_23_M69_noxref_d ) capacitor \
 c=0.0173476f //x=20.02 //y=6.02 //x2=20.095 //y2=5.02
cc_2522 ( N_noxref_7_M70_noxref_g N_noxref_23_M69_noxref_d ) capacitor \
 c=0.0179769f //x=20.46 //y=6.02 //x2=20.095 //y2=5.02
cc_2523 ( N_noxref_7_c_2728_n N_noxref_26_c_8231_n ) capacitor c=0.0034165f \
 //x=0.81 //y=1.915 //x2=0.59 //y2=1.505
cc_2524 ( N_noxref_7_c_2715_n N_noxref_26_c_8214_n ) capacitor c=0.00179505f \
 //x=9.875 //y=4.07 //x2=1.475 //y2=1.59
cc_2525 ( N_noxref_7_c_2716_n N_noxref_26_c_8214_n ) capacitor c=0.00102628f \
 //x=1.225 //y=4.07 //x2=1.475 //y2=1.59
cc_2526 ( N_noxref_7_c_2717_n N_noxref_26_c_8214_n ) capacitor c=0.0122033f \
 //x=1.11 //y=2.08 //x2=1.475 //y2=1.59
cc_2527 ( N_noxref_7_c_2727_n N_noxref_26_c_8214_n ) capacitor c=0.00703864f \
 //x=0.81 //y=1.53 //x2=1.475 //y2=1.59
cc_2528 ( N_noxref_7_c_2728_n N_noxref_26_c_8214_n ) capacitor c=0.0259045f \
 //x=0.81 //y=1.915 //x2=1.475 //y2=1.59
cc_2529 ( N_noxref_7_c_2730_n N_noxref_26_c_8214_n ) capacitor c=0.00708583f \
 //x=1.185 //y=1.375 //x2=1.475 //y2=1.59
cc_2530 ( N_noxref_7_c_2733_n N_noxref_26_c_8214_n ) capacitor c=0.00698822f \
 //x=1.34 //y=1.22 //x2=1.475 //y2=1.59
cc_2531 ( N_noxref_7_c_2715_n N_noxref_26_c_8239_n ) capacitor c=0.0058169f \
 //x=9.875 //y=4.07 //x2=2.445 //y2=1.59
cc_2532 ( N_noxref_7_c_2715_n N_noxref_26_M0_noxref_s ) capacitor \
 c=0.00262629f //x=9.875 //y=4.07 //x2=0.455 //y2=0.375
cc_2533 ( N_noxref_7_c_2724_n N_noxref_26_M0_noxref_s ) capacitor c=0.0327271f \
 //x=0.81 //y=0.875 //x2=0.455 //y2=0.375
cc_2534 ( N_noxref_7_c_2727_n N_noxref_26_M0_noxref_s ) capacitor \
 c=7.99997e-19 //x=0.81 //y=1.53 //x2=0.455 //y2=0.375
cc_2535 ( N_noxref_7_c_2728_n N_noxref_26_M0_noxref_s ) capacitor \
 c=0.00122123f //x=0.81 //y=1.915 //x2=0.455 //y2=0.375
cc_2536 ( N_noxref_7_c_2731_n N_noxref_26_M0_noxref_s ) capacitor c=0.0121427f \
 //x=1.34 //y=0.875 //x2=0.455 //y2=0.375
cc_2537 ( N_noxref_7_c_2715_n N_noxref_27_c_8261_n ) capacitor c=0.0020922f \
 //x=9.875 //y=4.07 //x2=3.015 //y2=0.995
cc_2538 ( N_noxref_7_c_2715_n N_noxref_27_M2_noxref_s ) capacitor \
 c=0.00143334f //x=9.875 //y=4.07 //x2=2.965 //y2=0.375
cc_2539 ( N_noxref_7_c_2817_n N_noxref_29_c_8375_n ) capacitor c=0.00623646f \
 //x=10.025 //y=1.56 //x2=9.805 //y2=1.495
cc_2540 ( N_noxref_7_c_2822_n N_noxref_29_c_8375_n ) capacitor c=0.00174019f \
 //x=9.99 //y=2.08 //x2=9.805 //y2=1.495
cc_2541 ( N_noxref_7_c_2718_n N_noxref_29_c_8376_n ) capacitor c=0.00158203f \
 //x=9.99 //y=2.08 //x2=10.69 //y2=0.53
cc_2542 ( N_noxref_7_c_2812_n N_noxref_29_c_8376_n ) capacitor c=0.0188655f \
 //x=10.025 //y=0.905 //x2=10.69 //y2=0.53
cc_2543 ( N_noxref_7_c_2820_n N_noxref_29_c_8376_n ) capacitor c=0.00656458f \
 //x=10.555 //y=0.905 //x2=10.69 //y2=0.53
cc_2544 ( N_noxref_7_c_2822_n N_noxref_29_c_8376_n ) capacitor c=2.1838e-19 \
 //x=9.99 //y=2.08 //x2=10.69 //y2=0.53
cc_2545 ( N_noxref_7_c_2812_n N_noxref_29_M5_noxref_s ) capacitor \
 c=0.00623646f //x=10.025 //y=0.905 //x2=8.7 //y2=0.365
cc_2546 ( N_noxref_7_c_2820_n N_noxref_29_M5_noxref_s ) capacitor c=0.0143002f \
 //x=10.555 //y=0.905 //x2=8.7 //y2=0.365
cc_2547 ( N_noxref_7_c_2821_n N_noxref_29_M5_noxref_s ) capacitor \
 c=0.00290153f //x=10.555 //y=1.25 //x2=8.7 //y2=0.365
cc_2548 ( N_noxref_7_c_2919_p N_noxref_30_c_8439_n ) capacitor c=3.15806e-19 \
 //x=13.705 //y=1.655 //x2=12.165 //y2=1.495
cc_2549 ( N_noxref_7_c_2919_p N_noxref_30_c_8427_n ) capacitor c=0.0203424f \
 //x=13.705 //y=1.655 //x2=13.135 //y2=1.495
cc_2550 ( N_noxref_7_c_2720_n N_noxref_30_c_8428_n ) capacitor c=0.00461444f \
 //x=13.975 //y=1.655 //x2=14.02 //y2=0.53
cc_2551 ( N_noxref_7_M8_noxref_d N_noxref_30_c_8428_n ) capacitor c=0.0116735f \
 //x=13.43 //y=0.905 //x2=14.02 //y2=0.53
cc_2552 ( N_noxref_7_c_2720_n N_noxref_30_M7_noxref_s ) capacitor c=0.0137901f \
 //x=13.975 //y=1.655 //x2=12.03 //y2=0.365
cc_2553 ( N_noxref_7_M8_noxref_d N_noxref_30_M7_noxref_s ) capacitor \
 c=0.043966f //x=13.43 //y=0.905 //x2=12.03 //y2=0.365
cc_2554 ( N_noxref_7_c_2720_n N_noxref_31_c_8491_n ) capacitor c=3.22188e-19 \
 //x=13.975 //y=1.655 //x2=15.495 //y2=1.495
cc_2555 ( N_noxref_7_c_2902_n N_noxref_32_c_8531_n ) capacitor c=0.00623646f \
 //x=20.015 //y=1.56 //x2=19.795 //y2=1.495
cc_2556 ( N_noxref_7_c_2907_n N_noxref_32_c_8531_n ) capacitor c=0.00174019f \
 //x=19.98 //y=2.08 //x2=19.795 //y2=1.495
cc_2557 ( N_noxref_7_c_2722_n N_noxref_32_c_8532_n ) capacitor c=0.00158203f \
 //x=19.98 //y=2.08 //x2=20.68 //y2=0.53
cc_2558 ( N_noxref_7_c_2897_n N_noxref_32_c_8532_n ) capacitor c=0.0188655f \
 //x=20.015 //y=0.905 //x2=20.68 //y2=0.53
cc_2559 ( N_noxref_7_c_2905_n N_noxref_32_c_8532_n ) capacitor c=0.00656458f \
 //x=20.545 //y=0.905 //x2=20.68 //y2=0.53
cc_2560 ( N_noxref_7_c_2907_n N_noxref_32_c_8532_n ) capacitor c=2.1838e-19 \
 //x=19.98 //y=2.08 //x2=20.68 //y2=0.53
cc_2561 ( N_noxref_7_c_2897_n N_noxref_32_M11_noxref_s ) capacitor \
 c=0.00623646f //x=20.015 //y=0.905 //x2=18.69 //y2=0.365
cc_2562 ( N_noxref_7_c_2905_n N_noxref_32_M11_noxref_s ) capacitor \
 c=0.0143002f //x=20.545 //y=0.905 //x2=18.69 //y2=0.365
cc_2563 ( N_noxref_7_c_2906_n N_noxref_32_M11_noxref_s ) capacitor \
 c=0.00290153f //x=20.545 //y=1.25 //x2=18.69 //y2=0.365
cc_2564 ( N_noxref_8_c_3121_p N_noxref_9_c_3347_n ) capacitor c=0.011463f \
 //x=30.595 //y=3.33 //x2=32.305 //y2=3.33
cc_2565 ( N_noxref_8_M82_noxref_g N_noxref_9_c_3316_n ) capacitor c=0.0169521f \
 //x=31.05 //y=6.02 //x2=31.625 //y2=5.2
cc_2566 ( N_noxref_8_c_3071_n N_noxref_9_c_3320_n ) capacitor c=0.00539951f \
 //x=30.71 //y=2.08 //x2=30.915 //y2=5.2
cc_2567 ( N_noxref_8_M81_noxref_g N_noxref_9_c_3320_n ) capacitor c=0.0177326f \
 //x=30.61 //y=6.02 //x2=30.915 //y2=5.2
cc_2568 ( N_noxref_8_c_3109_n N_noxref_9_c_3320_n ) capacitor c=0.00581252f \
 //x=30.71 //y=4.7 //x2=30.915 //y2=5.2
cc_2569 ( N_noxref_8_c_3070_n N_noxref_9_c_3301_n ) capacitor c=3.49822e-19 \
 //x=28.86 //y=3.33 //x2=32.19 //y2=3.33
cc_2570 ( N_noxref_8_c_3071_n N_noxref_9_c_3301_n ) capacitor c=0.00277094f \
 //x=30.71 //y=2.08 //x2=32.19 //y2=3.33
cc_2571 ( N_noxref_8_M82_noxref_g N_noxref_9_M81_noxref_d ) capacitor \
 c=0.0173476f //x=31.05 //y=6.02 //x2=30.685 //y2=5.02
cc_2572 ( N_noxref_8_c_3129_p N_noxref_10_c_3523_n ) capacitor c=0.146341f \
 //x=28.745 //y=3.33 //x2=27.265 //y2=3.7
cc_2573 ( N_noxref_8_c_3129_p N_noxref_10_c_3524_n ) capacitor c=0.0294746f \
 //x=28.745 //y=3.33 //x2=25.645 //y2=3.7
cc_2574 ( N_noxref_8_c_3068_n N_noxref_10_c_3524_n ) capacitor c=0.00687545f \
 //x=24.79 //y=2.08 //x2=25.645 //y2=3.7
cc_2575 ( N_noxref_8_c_3129_p N_noxref_10_c_3526_n ) capacitor c=0.108749f \
 //x=28.745 //y=3.33 //x2=37.255 //y2=3.7
cc_2576 ( N_noxref_8_c_3121_p N_noxref_10_c_3526_n ) capacitor c=0.175696f \
 //x=30.595 //y=3.33 //x2=37.255 //y2=3.7
cc_2577 ( N_noxref_8_c_3134_p N_noxref_10_c_3526_n ) capacitor c=0.0267668f \
 //x=28.975 //y=3.33 //x2=37.255 //y2=3.7
cc_2578 ( N_noxref_8_c_3070_n N_noxref_10_c_3526_n ) capacitor c=0.0206034f \
 //x=28.86 //y=3.33 //x2=37.255 //y2=3.7
cc_2579 ( N_noxref_8_c_3071_n N_noxref_10_c_3526_n ) capacitor c=0.0205831f \
 //x=30.71 //y=2.08 //x2=37.255 //y2=3.7
cc_2580 ( N_noxref_8_c_3129_p N_noxref_10_c_3531_n ) capacitor c=0.0266674f \
 //x=28.745 //y=3.33 //x2=27.495 //y2=3.7
cc_2581 ( N_noxref_8_M75_noxref_g N_noxref_10_c_3483_n ) capacitor c=0.01736f \
 //x=24.53 //y=6.02 //x2=24.665 //y2=5.155
cc_2582 ( N_noxref_8_M76_noxref_g N_noxref_10_c_3487_n ) capacitor \
 c=0.0194981f //x=24.97 //y=6.02 //x2=25.445 //y2=5.155
cc_2583 ( N_noxref_8_c_3140_p N_noxref_10_c_3487_n ) capacitor c=0.00201851f \
 //x=24.79 //y=4.7 //x2=25.445 //y2=5.155
cc_2584 ( N_noxref_8_c_3141_p N_noxref_10_c_3453_n ) capacitor c=0.00359704f \
 //x=25.155 //y=1.415 //x2=25.445 //y2=1.665
cc_2585 ( N_noxref_8_c_3142_p N_noxref_10_c_3453_n ) capacitor c=0.00457401f \
 //x=25.31 //y=1.26 //x2=25.445 //y2=1.665
cc_2586 ( N_noxref_8_c_3129_p N_noxref_10_c_3491_n ) capacitor c=0.0206036f \
 //x=28.745 //y=3.33 //x2=25.53 //y2=3.7
cc_2587 ( N_noxref_8_c_3144_p N_noxref_10_c_3491_n ) capacitor c=0.00117715f \
 //x=24.905 //y=3.33 //x2=25.53 //y2=3.7
cc_2588 ( N_noxref_8_c_3068_n N_noxref_10_c_3491_n ) capacitor c=0.0780861f \
 //x=24.79 //y=2.08 //x2=25.53 //y2=3.7
cc_2589 ( N_noxref_8_c_3070_n N_noxref_10_c_3491_n ) capacitor c=3.52729e-19 \
 //x=28.86 //y=3.33 //x2=25.53 //y2=3.7
cc_2590 ( N_noxref_8_c_3147_p N_noxref_10_c_3491_n ) capacitor c=0.00877984f \
 //x=24.79 //y=2.08 //x2=25.53 //y2=3.7
cc_2591 ( N_noxref_8_c_3148_p N_noxref_10_c_3491_n ) capacitor c=0.00283672f \
 //x=24.79 //y=1.915 //x2=25.53 //y2=3.7
cc_2592 ( N_noxref_8_c_3140_p N_noxref_10_c_3491_n ) capacitor c=0.013693f \
 //x=24.79 //y=4.7 //x2=25.53 //y2=3.7
cc_2593 ( N_noxref_8_c_3129_p N_noxref_10_c_3454_n ) capacitor c=0.020575f \
 //x=28.745 //y=3.33 //x2=27.38 //y2=2.08
cc_2594 ( N_noxref_8_c_3068_n N_noxref_10_c_3454_n ) capacitor c=8.46099e-19 \
 //x=24.79 //y=2.08 //x2=27.38 //y2=2.08
cc_2595 ( N_noxref_8_c_3090_n N_noxref_10_c_3454_n ) capacitor c=0.00521572f \
 //x=27.585 //y=5.2 //x2=27.38 //y2=2.08
cc_2596 ( N_noxref_8_c_3070_n N_noxref_10_c_3454_n ) capacitor c=0.00288966f \
 //x=28.86 //y=3.33 //x2=27.38 //y2=2.08
cc_2597 ( N_noxref_8_c_3068_n N_noxref_10_c_3548_n ) capacitor c=0.0171303f \
 //x=24.79 //y=2.08 //x2=24.75 //y2=5.155
cc_2598 ( N_noxref_8_c_3140_p N_noxref_10_c_3548_n ) capacitor c=0.00475601f \
 //x=24.79 //y=4.7 //x2=24.75 //y2=5.155
cc_2599 ( N_noxref_8_c_3090_n N_noxref_10_M77_noxref_g ) capacitor \
 c=0.0177326f //x=27.585 //y=5.2 //x2=27.28 //y2=6.02
cc_2600 ( N_noxref_8_c_3086_n N_noxref_10_M78_noxref_g ) capacitor \
 c=0.0169521f //x=28.295 //y=5.2 //x2=27.72 //y2=6.02
cc_2601 ( N_noxref_8_M77_noxref_d N_noxref_10_M78_noxref_g ) capacitor \
 c=0.0173476f //x=27.355 //y=5.02 //x2=27.72 //y2=6.02
cc_2602 ( N_noxref_8_c_3090_n N_noxref_10_c_3506_n ) capacitor c=0.00581252f \
 //x=27.585 //y=5.2 //x2=27.38 //y2=4.7
cc_2603 ( N_noxref_8_c_3160_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00217566f //x=24.78 //y=0.915 //x2=24.855 //y2=0.915
cc_2604 ( N_noxref_8_c_3161_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.0034598f //x=24.78 //y=1.26 //x2=24.855 //y2=0.915
cc_2605 ( N_noxref_8_c_3162_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00544291f //x=24.78 //y=1.57 //x2=24.855 //y2=0.915
cc_2606 ( N_noxref_8_c_3163_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00241102f //x=25.155 //y=0.76 //x2=24.855 //y2=0.915
cc_2607 ( N_noxref_8_c_3141_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.0140297f //x=25.155 //y=1.415 //x2=24.855 //y2=0.915
cc_2608 ( N_noxref_8_c_3165_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00219619f //x=25.31 //y=0.915 //x2=24.855 //y2=0.915
cc_2609 ( N_noxref_8_c_3142_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00603828f //x=25.31 //y=1.26 //x2=24.855 //y2=0.915
cc_2610 ( N_noxref_8_c_3148_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00661782f //x=24.79 //y=1.915 //x2=24.855 //y2=0.915
cc_2611 ( N_noxref_8_M75_noxref_g N_noxref_10_M75_noxref_d ) capacitor \
 c=0.0180032f //x=24.53 //y=6.02 //x2=24.605 //y2=5.02
cc_2612 ( N_noxref_8_M76_noxref_g N_noxref_10_M75_noxref_d ) capacitor \
 c=0.0194246f //x=24.97 //y=6.02 //x2=24.605 //y2=5.02
cc_2613 ( N_noxref_8_c_3129_p N_noxref_12_c_3882_n ) capacitor c=0.0428508f \
 //x=28.745 //y=3.33 //x2=31.335 //y2=4.07
cc_2614 ( N_noxref_8_c_3144_p N_noxref_12_c_3882_n ) capacitor c=0.0135672f \
 //x=24.905 //y=3.33 //x2=31.335 //y2=4.07
cc_2615 ( N_noxref_8_c_3121_p N_noxref_12_c_3882_n ) capacitor c=0.0110241f \
 //x=30.595 //y=3.33 //x2=31.335 //y2=4.07
cc_2616 ( N_noxref_8_c_3134_p N_noxref_12_c_3882_n ) capacitor c=5.70661e-19 \
 //x=28.975 //y=3.33 //x2=31.335 //y2=4.07
cc_2617 ( N_noxref_8_c_3068_n N_noxref_12_c_3882_n ) capacitor c=0.0206302f \
 //x=24.79 //y=2.08 //x2=31.335 //y2=4.07
cc_2618 ( N_noxref_8_c_3070_n N_noxref_12_c_3882_n ) capacitor c=0.0181936f \
 //x=28.86 //y=3.33 //x2=31.335 //y2=4.07
cc_2619 ( N_noxref_8_c_3071_n N_noxref_12_c_3882_n ) capacitor c=0.0184765f \
 //x=30.71 //y=2.08 //x2=31.335 //y2=4.07
cc_2620 ( N_noxref_8_c_3071_n N_noxref_12_c_3944_n ) capacitor c=0.00179385f \
 //x=30.71 //y=2.08 //x2=31.565 //y2=4.07
cc_2621 ( N_noxref_8_c_3068_n N_noxref_12_c_3862_n ) capacitor c=0.00137085f \
 //x=24.79 //y=2.08 //x2=22.57 //y2=2.08
cc_2622 ( N_noxref_8_c_3071_n N_noxref_12_c_3946_n ) capacitor c=0.00400249f \
 //x=30.71 //y=2.08 //x2=31.45 //y2=4.535
cc_2623 ( N_noxref_8_c_3109_n N_noxref_12_c_3946_n ) capacitor c=0.00417994f \
 //x=30.71 //y=4.7 //x2=31.45 //y2=4.535
cc_2624 ( N_noxref_8_c_3121_p N_noxref_12_c_3863_n ) capacitor c=0.00318578f \
 //x=30.595 //y=3.33 //x2=31.45 //y2=2.08
cc_2625 ( N_noxref_8_c_3070_n N_noxref_12_c_3863_n ) capacitor c=8.48165e-19 \
 //x=28.86 //y=3.33 //x2=31.45 //y2=2.08
cc_2626 ( N_noxref_8_c_3071_n N_noxref_12_c_3863_n ) capacitor c=0.0743975f \
 //x=30.71 //y=2.08 //x2=31.45 //y2=2.08
cc_2627 ( N_noxref_8_c_3076_n N_noxref_12_c_3863_n ) capacitor c=0.00308814f \
 //x=30.515 //y=1.915 //x2=31.45 //y2=2.08
cc_2628 ( N_noxref_8_M81_noxref_g N_noxref_12_M83_noxref_g ) capacitor \
 c=0.0104611f //x=30.61 //y=6.02 //x2=31.49 //y2=6.02
cc_2629 ( N_noxref_8_M82_noxref_g N_noxref_12_M83_noxref_g ) capacitor \
 c=0.106811f //x=31.05 //y=6.02 //x2=31.49 //y2=6.02
cc_2630 ( N_noxref_8_M82_noxref_g N_noxref_12_M84_noxref_g ) capacitor \
 c=0.0100341f //x=31.05 //y=6.02 //x2=31.93 //y2=6.02
cc_2631 ( N_noxref_8_c_3072_n N_noxref_12_c_3955_n ) capacitor c=4.86506e-19 \
 //x=30.515 //y=0.865 //x2=31.485 //y2=0.905
cc_2632 ( N_noxref_8_c_3074_n N_noxref_12_c_3955_n ) capacitor c=0.00152104f \
 //x=30.515 //y=1.21 //x2=31.485 //y2=0.905
cc_2633 ( N_noxref_8_c_3079_n N_noxref_12_c_3955_n ) capacitor c=0.0151475f \
 //x=31.045 //y=0.865 //x2=31.485 //y2=0.905
cc_2634 ( N_noxref_8_c_3075_n N_noxref_12_c_3958_n ) capacitor c=0.00109982f \
 //x=30.515 //y=1.52 //x2=31.485 //y2=1.25
cc_2635 ( N_noxref_8_c_3081_n N_noxref_12_c_3958_n ) capacitor c=0.0111064f \
 //x=31.045 //y=1.21 //x2=31.485 //y2=1.25
cc_2636 ( N_noxref_8_c_3075_n N_noxref_12_c_3960_n ) capacitor c=9.57794e-19 \
 //x=30.515 //y=1.52 //x2=31.485 //y2=1.56
cc_2637 ( N_noxref_8_c_3076_n N_noxref_12_c_3960_n ) capacitor c=0.00662747f \
 //x=30.515 //y=1.915 //x2=31.485 //y2=1.56
cc_2638 ( N_noxref_8_c_3081_n N_noxref_12_c_3960_n ) capacitor c=0.00862358f \
 //x=31.045 //y=1.21 //x2=31.485 //y2=1.56
cc_2639 ( N_noxref_8_c_3079_n N_noxref_12_c_3963_n ) capacitor c=0.00124821f \
 //x=31.045 //y=0.865 //x2=32.015 //y2=0.905
cc_2640 ( N_noxref_8_c_3081_n N_noxref_12_c_3964_n ) capacitor c=0.00200715f \
 //x=31.045 //y=1.21 //x2=32.015 //y2=1.25
cc_2641 ( N_noxref_8_c_3071_n N_noxref_12_c_3965_n ) capacitor c=0.00307062f \
 //x=30.71 //y=2.08 //x2=31.45 //y2=2.08
cc_2642 ( N_noxref_8_c_3076_n N_noxref_12_c_3965_n ) capacitor c=0.0179092f \
 //x=30.515 //y=1.915 //x2=31.45 //y2=2.08
cc_2643 ( N_noxref_8_c_3071_n N_noxref_12_c_3967_n ) capacitor c=0.00344981f \
 //x=30.71 //y=2.08 //x2=31.48 //y2=4.7
cc_2644 ( N_noxref_8_c_3109_n N_noxref_12_c_3967_n ) capacitor c=0.0293367f \
 //x=30.71 //y=4.7 //x2=31.48 //y2=4.7
cc_2645 ( N_noxref_8_c_3129_p N_D_c_4217_n ) capacitor c=0.0235344f //x=28.745 \
 //y=3.33 //x2=28.005 //y2=2.59
cc_2646 ( N_noxref_8_c_3144_p N_D_c_4217_n ) capacitor c=9.8111e-19 //x=24.905 \
 //y=3.33 //x2=28.005 //y2=2.59
cc_2647 ( N_noxref_8_c_3068_n N_D_c_4217_n ) capacitor c=0.021502f //x=24.79 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2648 ( N_noxref_8_c_3147_p N_D_c_4217_n ) capacitor c=0.0021022f //x=24.79 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2649 ( N_noxref_8_c_3129_p N_D_c_4238_n ) capacitor c=0.00538961f \
 //x=28.745 //y=3.33 //x2=49.465 //y2=2.59
cc_2650 ( N_noxref_8_c_3121_p N_D_c_4238_n ) capacitor c=0.0125396f //x=30.595 \
 //y=3.33 //x2=49.465 //y2=2.59
cc_2651 ( N_noxref_8_c_3134_p N_D_c_4238_n ) capacitor c=5.75258e-19 \
 //x=28.975 //y=3.33 //x2=49.465 //y2=2.59
cc_2652 ( N_noxref_8_c_3209_p N_D_c_4238_n ) capacitor c=0.0102711f //x=28.505 \
 //y=1.655 //x2=49.465 //y2=2.59
cc_2653 ( N_noxref_8_c_3070_n N_D_c_4238_n ) capacitor c=0.0210598f //x=28.86 \
 //y=3.33 //x2=49.465 //y2=2.59
cc_2654 ( N_noxref_8_c_3071_n N_D_c_4238_n ) capacitor c=0.0213243f //x=30.71 \
 //y=2.08 //x2=49.465 //y2=2.59
cc_2655 ( N_noxref_8_c_3076_n N_D_c_4238_n ) capacitor c=0.0052136f //x=30.515 \
 //y=1.915 //x2=49.465 //y2=2.59
cc_2656 ( N_noxref_8_c_3129_p N_D_c_4251_n ) capacitor c=6.67046e-19 \
 //x=28.745 //y=3.33 //x2=28.235 //y2=2.59
cc_2657 ( N_noxref_8_c_3070_n N_D_c_4251_n ) capacitor c=0.00179385f //x=28.86 \
 //y=3.33 //x2=28.235 //y2=2.59
cc_2658 ( N_noxref_8_c_3086_n N_D_c_4381_n ) capacitor c=0.0127164f //x=28.295 \
 //y=5.2 //x2=28.12 //y2=4.535
cc_2659 ( N_noxref_8_c_3070_n N_D_c_4381_n ) capacitor c=0.0101284f //x=28.86 \
 //y=3.33 //x2=28.12 //y2=4.535
cc_2660 ( N_noxref_8_c_3129_p N_D_c_4255_n ) capacitor c=0.0169786f //x=28.745 \
 //y=3.33 //x2=28.12 //y2=2.08
cc_2661 ( N_noxref_8_c_3134_p N_D_c_4255_n ) capacitor c=0.00117715f \
 //x=28.975 //y=3.33 //x2=28.12 //y2=2.08
cc_2662 ( N_noxref_8_c_3070_n N_D_c_4255_n ) capacitor c=0.0678027f //x=28.86 \
 //y=3.33 //x2=28.12 //y2=2.08
cc_2663 ( N_noxref_8_c_3071_n N_D_c_4255_n ) capacitor c=6.55913e-19 //x=30.71 \
 //y=2.08 //x2=28.12 //y2=2.08
cc_2664 ( N_noxref_8_c_3086_n N_D_M79_noxref_g ) capacitor c=0.0166421f \
 //x=28.295 //y=5.2 //x2=28.16 //y2=6.02
cc_2665 ( N_noxref_8_M79_noxref_d N_D_M79_noxref_g ) capacitor c=0.0173476f \
 //x=28.235 //y=5.02 //x2=28.16 //y2=6.02
cc_2666 ( N_noxref_8_c_3092_n N_D_M80_noxref_g ) capacitor c=0.018922f \
 //x=28.775 //y=5.2 //x2=28.6 //y2=6.02
cc_2667 ( N_noxref_8_M79_noxref_d N_D_M80_noxref_g ) capacitor c=0.0179769f \
 //x=28.235 //y=5.02 //x2=28.6 //y2=6.02
cc_2668 ( N_noxref_8_M17_noxref_d N_D_c_4391_n ) capacitor c=0.00217566f \
 //x=28.23 //y=0.905 //x2=28.155 //y2=0.905
cc_2669 ( N_noxref_8_M17_noxref_d N_D_c_4392_n ) capacitor c=0.0034598f \
 //x=28.23 //y=0.905 //x2=28.155 //y2=1.25
cc_2670 ( N_noxref_8_M17_noxref_d N_D_c_4393_n ) capacitor c=0.00656319f \
 //x=28.23 //y=0.905 //x2=28.155 //y2=1.56
cc_2671 ( N_noxref_8_c_3070_n N_D_c_4394_n ) capacitor c=0.0142673f //x=28.86 \
 //y=3.33 //x2=28.525 //y2=4.79
cc_2672 ( N_noxref_8_c_3229_p N_D_c_4394_n ) capacitor c=0.00407665f //x=28.38 \
 //y=5.2 //x2=28.525 //y2=4.79
cc_2673 ( N_noxref_8_M17_noxref_d N_D_c_4396_n ) capacitor c=0.00241102f \
 //x=28.23 //y=0.905 //x2=28.53 //y2=0.75
cc_2674 ( N_noxref_8_c_3069_n N_D_c_4397_n ) capacitor c=0.00359704f \
 //x=28.775 //y=1.655 //x2=28.53 //y2=1.405
cc_2675 ( N_noxref_8_M17_noxref_d N_D_c_4397_n ) capacitor c=0.0138845f \
 //x=28.23 //y=0.905 //x2=28.53 //y2=1.405
cc_2676 ( N_noxref_8_M17_noxref_d N_D_c_4399_n ) capacitor c=0.00132245f \
 //x=28.23 //y=0.905 //x2=28.685 //y2=0.905
cc_2677 ( N_noxref_8_c_3069_n N_D_c_4400_n ) capacitor c=0.00457401f \
 //x=28.775 //y=1.655 //x2=28.685 //y2=1.25
cc_2678 ( N_noxref_8_M17_noxref_d N_D_c_4400_n ) capacitor c=0.00566463f \
 //x=28.23 //y=0.905 //x2=28.685 //y2=1.25
cc_2679 ( N_noxref_8_c_3070_n N_D_c_4402_n ) capacitor c=0.00877984f //x=28.86 \
 //y=3.33 //x2=28.12 //y2=2.08
cc_2680 ( N_noxref_8_c_3070_n N_D_c_4403_n ) capacitor c=0.00306024f //x=28.86 \
 //y=3.33 //x2=28.12 //y2=1.915
cc_2681 ( N_noxref_8_M17_noxref_d N_D_c_4403_n ) capacitor c=0.00660593f \
 //x=28.23 //y=0.905 //x2=28.12 //y2=1.915
cc_2682 ( N_noxref_8_c_3086_n N_D_c_4405_n ) capacitor c=0.00346527f \
 //x=28.295 //y=5.2 //x2=28.15 //y2=4.7
cc_2683 ( N_noxref_8_c_3070_n N_D_c_4405_n ) capacitor c=0.00533692f //x=28.86 \
 //y=3.33 //x2=28.15 //y2=4.7
cc_2684 ( N_noxref_8_c_3129_p N_CLK_c_5061_n ) capacitor c=0.00360213f \
 //x=28.745 //y=3.33 //x2=34.665 //y2=4.44
cc_2685 ( N_noxref_8_c_3144_p N_CLK_c_5061_n ) capacitor c=4.49102e-19 \
 //x=24.905 //y=3.33 //x2=34.665 //y2=4.44
cc_2686 ( N_noxref_8_c_3068_n N_CLK_c_5061_n ) capacitor c=0.0200057f \
 //x=24.79 //y=2.08 //x2=34.665 //y2=4.44
cc_2687 ( N_noxref_8_c_3086_n N_CLK_c_5061_n ) capacitor c=0.0185297f \
 //x=28.295 //y=5.2 //x2=34.665 //y2=4.44
cc_2688 ( N_noxref_8_c_3090_n N_CLK_c_5061_n ) capacitor c=0.0181237f \
 //x=27.585 //y=5.2 //x2=34.665 //y2=4.44
cc_2689 ( N_noxref_8_c_3070_n N_CLK_c_5061_n ) capacitor c=0.0208321f \
 //x=28.86 //y=3.33 //x2=34.665 //y2=4.44
cc_2690 ( N_noxref_8_c_3071_n N_CLK_c_5061_n ) capacitor c=0.0198304f \
 //x=30.71 //y=2.08 //x2=34.665 //y2=4.44
cc_2691 ( N_noxref_8_c_3140_p N_CLK_c_5061_n ) capacitor c=0.0111881f \
 //x=24.79 //y=4.7 //x2=34.665 //y2=4.44
cc_2692 ( N_noxref_8_c_3109_n N_CLK_c_5061_n ) capacitor c=0.0107057f \
 //x=30.71 //y=4.7 //x2=34.665 //y2=4.44
cc_2693 ( N_noxref_8_c_3068_n N_CLK_c_5079_n ) capacitor c=0.00153281f \
 //x=24.79 //y=2.08 //x2=23.795 //y2=4.44
cc_2694 ( N_noxref_8_c_3144_p N_CLK_c_5028_n ) capacitor c=0.00526349f \
 //x=24.905 //y=3.33 //x2=23.68 //y2=2.08
cc_2695 ( N_noxref_8_c_3068_n N_CLK_c_5028_n ) capacitor c=0.0463871f \
 //x=24.79 //y=2.08 //x2=23.68 //y2=2.08
cc_2696 ( N_noxref_8_c_3147_p N_CLK_c_5028_n ) capacitor c=0.00228632f \
 //x=24.79 //y=2.08 //x2=23.68 //y2=2.08
cc_2697 ( N_noxref_8_c_3140_p N_CLK_c_5028_n ) capacitor c=0.00218014f \
 //x=24.79 //y=4.7 //x2=23.68 //y2=2.08
cc_2698 ( N_noxref_8_M75_noxref_g N_CLK_M73_noxref_g ) capacitor c=0.0101598f \
 //x=24.53 //y=6.02 //x2=23.65 //y2=6.02
cc_2699 ( N_noxref_8_M75_noxref_g N_CLK_M74_noxref_g ) capacitor c=0.0602553f \
 //x=24.53 //y=6.02 //x2=24.09 //y2=6.02
cc_2700 ( N_noxref_8_M76_noxref_g N_CLK_M74_noxref_g ) capacitor c=0.0101598f \
 //x=24.97 //y=6.02 //x2=24.09 //y2=6.02
cc_2701 ( N_noxref_8_c_3160_p N_CLK_c_5347_n ) capacitor c=0.00456962f \
 //x=24.78 //y=0.915 //x2=23.77 //y2=0.91
cc_2702 ( N_noxref_8_c_3161_p N_CLK_c_5348_n ) capacitor c=0.00438372f \
 //x=24.78 //y=1.26 //x2=23.77 //y2=1.22
cc_2703 ( N_noxref_8_c_3162_p N_CLK_c_5349_n ) capacitor c=0.00438372f \
 //x=24.78 //y=1.57 //x2=23.77 //y2=1.45
cc_2704 ( N_noxref_8_c_3068_n N_CLK_c_5350_n ) capacitor c=0.0023343f \
 //x=24.79 //y=2.08 //x2=23.77 //y2=1.915
cc_2705 ( N_noxref_8_c_3147_p N_CLK_c_5350_n ) capacitor c=0.00933826f \
 //x=24.79 //y=2.08 //x2=23.77 //y2=1.915
cc_2706 ( N_noxref_8_c_3148_p N_CLK_c_5350_n ) capacitor c=0.00438372f \
 //x=24.79 //y=1.915 //x2=23.77 //y2=1.915
cc_2707 ( N_noxref_8_c_3140_p N_CLK_c_5353_n ) capacitor c=0.0611812f \
 //x=24.79 //y=4.7 //x2=24.015 //y2=4.79
cc_2708 ( N_noxref_8_c_3068_n N_CLK_c_5354_n ) capacitor c=0.00142741f \
 //x=24.79 //y=2.08 //x2=23.68 //y2=4.7
cc_2709 ( N_noxref_8_c_3140_p N_CLK_c_5354_n ) capacitor c=0.00487508f \
 //x=24.79 //y=4.7 //x2=23.68 //y2=4.7
cc_2710 ( N_noxref_8_c_3129_p N_noxref_23_c_7498_n ) capacitor c=0.336622f \
 //x=28.745 //y=3.33 //x2=70.185 //y2=2.96
cc_2711 ( N_noxref_8_c_3144_p N_noxref_23_c_7498_n ) capacitor c=0.0291389f \
 //x=24.905 //y=3.33 //x2=70.185 //y2=2.96
cc_2712 ( N_noxref_8_c_3121_p N_noxref_23_c_7498_n ) capacitor c=0.173509f \
 //x=30.595 //y=3.33 //x2=70.185 //y2=2.96
cc_2713 ( N_noxref_8_c_3134_p N_noxref_23_c_7498_n ) capacitor c=0.0266415f \
 //x=28.975 //y=3.33 //x2=70.185 //y2=2.96
cc_2714 ( N_noxref_8_c_3068_n N_noxref_23_c_7498_n ) capacitor c=0.0198264f \
 //x=24.79 //y=2.08 //x2=70.185 //y2=2.96
cc_2715 ( N_noxref_8_c_3070_n N_noxref_23_c_7498_n ) capacitor c=0.0206014f \
 //x=28.86 //y=3.33 //x2=70.185 //y2=2.96
cc_2716 ( N_noxref_8_c_3071_n N_noxref_23_c_7498_n ) capacitor c=0.0205758f \
 //x=30.71 //y=2.08 //x2=70.185 //y2=2.96
cc_2717 ( N_noxref_8_c_3068_n N_noxref_34_c_8631_n ) capacitor c=0.0020642f \
 //x=24.79 //y=2.08 //x2=25.445 //y2=0.54
cc_2718 ( N_noxref_8_c_3160_p N_noxref_34_c_8631_n ) capacitor c=0.0194423f \
 //x=24.78 //y=0.915 //x2=25.445 //y2=0.54
cc_2719 ( N_noxref_8_c_3165_p N_noxref_34_c_8631_n ) capacitor c=0.00656458f \
 //x=25.31 //y=0.915 //x2=25.445 //y2=0.54
cc_2720 ( N_noxref_8_c_3147_p N_noxref_34_c_8631_n ) capacitor c=2.20712e-19 \
 //x=24.79 //y=2.08 //x2=25.445 //y2=0.54
cc_2721 ( N_noxref_8_c_3161_p N_noxref_34_c_8644_n ) capacitor c=0.00538829f \
 //x=24.78 //y=1.26 //x2=24.56 //y2=0.995
cc_2722 ( N_noxref_8_c_3160_p N_noxref_34_M15_noxref_s ) capacitor \
 c=0.00538829f //x=24.78 //y=0.915 //x2=24.425 //y2=0.375
cc_2723 ( N_noxref_8_c_3162_p N_noxref_34_M15_noxref_s ) capacitor \
 c=0.00538829f //x=24.78 //y=1.57 //x2=24.425 //y2=0.375
cc_2724 ( N_noxref_8_c_3165_p N_noxref_34_M15_noxref_s ) capacitor \
 c=0.0143002f //x=25.31 //y=0.915 //x2=24.425 //y2=0.375
cc_2725 ( N_noxref_8_c_3142_p N_noxref_34_M15_noxref_s ) capacitor \
 c=0.00290153f //x=25.31 //y=1.26 //x2=24.425 //y2=0.375
cc_2726 ( N_noxref_8_c_3209_p N_noxref_35_c_8698_n ) capacitor c=3.15806e-19 \
 //x=28.505 //y=1.655 //x2=26.965 //y2=1.495
cc_2727 ( N_noxref_8_c_3209_p N_noxref_35_c_8686_n ) capacitor c=0.020324f \
 //x=28.505 //y=1.655 //x2=27.935 //y2=1.495
cc_2728 ( N_noxref_8_c_3069_n N_noxref_35_c_8687_n ) capacitor c=0.00461444f \
 //x=28.775 //y=1.655 //x2=28.82 //y2=0.53
cc_2729 ( N_noxref_8_M17_noxref_d N_noxref_35_c_8687_n ) capacitor \
 c=0.0116735f //x=28.23 //y=0.905 //x2=28.82 //y2=0.53
cc_2730 ( N_noxref_8_c_3069_n N_noxref_35_M16_noxref_s ) capacitor \
 c=0.0137901f //x=28.775 //y=1.655 //x2=26.83 //y2=0.365
cc_2731 ( N_noxref_8_M17_noxref_d N_noxref_35_M16_noxref_s ) capacitor \
 c=0.0439476f //x=28.23 //y=0.905 //x2=26.83 //y2=0.365
cc_2732 ( N_noxref_8_c_3069_n N_noxref_36_c_8752_n ) capacitor c=3.22188e-19 \
 //x=28.775 //y=1.655 //x2=30.295 //y2=1.495
cc_2733 ( N_noxref_8_c_3076_n N_noxref_36_c_8752_n ) capacitor c=0.0034165f \
 //x=30.515 //y=1.915 //x2=30.295 //y2=1.495
cc_2734 ( N_noxref_8_c_3071_n N_noxref_36_c_8733_n ) capacitor c=0.0118762f \
 //x=30.71 //y=2.08 //x2=31.18 //y2=1.58
cc_2735 ( N_noxref_8_c_3075_n N_noxref_36_c_8733_n ) capacitor c=0.00703567f \
 //x=30.515 //y=1.52 //x2=31.18 //y2=1.58
cc_2736 ( N_noxref_8_c_3076_n N_noxref_36_c_8733_n ) capacitor c=0.018562f \
 //x=30.515 //y=1.915 //x2=31.18 //y2=1.58
cc_2737 ( N_noxref_8_c_3078_n N_noxref_36_c_8733_n ) capacitor c=0.00780629f \
 //x=30.89 //y=1.365 //x2=31.18 //y2=1.58
cc_2738 ( N_noxref_8_c_3081_n N_noxref_36_c_8733_n ) capacitor c=0.00339872f \
 //x=31.045 //y=1.21 //x2=31.18 //y2=1.58
cc_2739 ( N_noxref_8_c_3076_n N_noxref_36_c_8740_n ) capacitor c=6.71402e-19 \
 //x=30.515 //y=1.915 //x2=31.265 //y2=1.495
cc_2740 ( N_noxref_8_c_3072_n N_noxref_36_M18_noxref_s ) capacitor \
 c=0.0326577f //x=30.515 //y=0.865 //x2=30.16 //y2=0.365
cc_2741 ( N_noxref_8_c_3075_n N_noxref_36_M18_noxref_s ) capacitor \
 c=3.48408e-19 //x=30.515 //y=1.52 //x2=30.16 //y2=0.365
cc_2742 ( N_noxref_8_c_3079_n N_noxref_36_M18_noxref_s ) capacitor \
 c=0.0120759f //x=31.045 //y=0.865 //x2=30.16 //y2=0.365
cc_2743 ( N_noxref_9_c_3355_p N_noxref_10_c_3526_n ) capacitor c=0.175696f \
 //x=33.925 //y=3.33 //x2=37.255 //y2=3.7
cc_2744 ( N_noxref_9_c_3347_n N_noxref_10_c_3526_n ) capacitor c=0.0293967f \
 //x=32.305 //y=3.33 //x2=37.255 //y2=3.7
cc_2745 ( N_noxref_9_c_3301_n N_noxref_10_c_3526_n ) capacitor c=0.0206034f \
 //x=32.19 //y=3.33 //x2=37.255 //y2=3.7
cc_2746 ( N_noxref_9_c_3302_n N_noxref_10_c_3526_n ) capacitor c=0.0205831f \
 //x=34.04 //y=2.08 //x2=37.255 //y2=3.7
cc_2747 ( N_noxref_9_c_3355_p N_noxref_12_c_3885_n ) capacitor c=0.0110241f \
 //x=33.925 //y=3.33 //x2=35.405 //y2=4.07
cc_2748 ( N_noxref_9_c_3347_n N_noxref_12_c_3885_n ) capacitor c=8.88358e-19 \
 //x=32.305 //y=3.33 //x2=35.405 //y2=4.07
cc_2749 ( N_noxref_9_c_3301_n N_noxref_12_c_3885_n ) capacitor c=0.0181936f \
 //x=32.19 //y=3.33 //x2=35.405 //y2=4.07
cc_2750 ( N_noxref_9_c_3302_n N_noxref_12_c_3885_n ) capacitor c=0.0184765f \
 //x=34.04 //y=2.08 //x2=35.405 //y2=4.07
cc_2751 ( N_noxref_9_c_3301_n N_noxref_12_c_3944_n ) capacitor c=0.00117715f \
 //x=32.19 //y=3.33 //x2=31.565 //y2=4.07
cc_2752 ( N_noxref_9_c_3316_n N_noxref_12_c_3946_n ) capacitor c=0.0126603f \
 //x=31.625 //y=5.2 //x2=31.45 //y2=4.535
cc_2753 ( N_noxref_9_c_3301_n N_noxref_12_c_3946_n ) capacitor c=0.0101319f \
 //x=32.19 //y=3.33 //x2=31.45 //y2=4.535
cc_2754 ( N_noxref_9_c_3347_n N_noxref_12_c_3863_n ) capacitor c=0.00329059f \
 //x=32.305 //y=3.33 //x2=31.45 //y2=2.08
cc_2755 ( N_noxref_9_c_3301_n N_noxref_12_c_3863_n ) capacitor c=0.0692733f \
 //x=32.19 //y=3.33 //x2=31.45 //y2=2.08
cc_2756 ( N_noxref_9_c_3302_n N_noxref_12_c_3863_n ) capacitor c=8.48165e-19 \
 //x=34.04 //y=2.08 //x2=31.45 //y2=2.08
cc_2757 ( N_noxref_9_M86_noxref_g N_noxref_12_c_3894_n ) capacitor \
 c=0.0169521f //x=34.38 //y=6.02 //x2=34.955 //y2=5.2
cc_2758 ( N_noxref_9_c_3302_n N_noxref_12_c_3898_n ) capacitor c=0.00539951f \
 //x=34.04 //y=2.08 //x2=34.245 //y2=5.2
cc_2759 ( N_noxref_9_M85_noxref_g N_noxref_12_c_3898_n ) capacitor \
 c=0.0177326f //x=33.94 //y=6.02 //x2=34.245 //y2=5.2
cc_2760 ( N_noxref_9_c_3335_n N_noxref_12_c_3898_n ) capacitor c=0.00581252f \
 //x=34.04 //y=4.7 //x2=34.245 //y2=5.2
cc_2761 ( N_noxref_9_c_3301_n N_noxref_12_c_3866_n ) capacitor c=3.49822e-19 \
 //x=32.19 //y=3.33 //x2=35.52 //y2=4.07
cc_2762 ( N_noxref_9_c_3302_n N_noxref_12_c_3866_n ) capacitor c=0.00321182f \
 //x=34.04 //y=2.08 //x2=35.52 //y2=4.07
cc_2763 ( N_noxref_9_c_3316_n N_noxref_12_M83_noxref_g ) capacitor \
 c=0.0166421f //x=31.625 //y=5.2 //x2=31.49 //y2=6.02
cc_2764 ( N_noxref_9_M83_noxref_d N_noxref_12_M83_noxref_g ) capacitor \
 c=0.0173476f //x=31.565 //y=5.02 //x2=31.49 //y2=6.02
cc_2765 ( N_noxref_9_c_3322_n N_noxref_12_M84_noxref_g ) capacitor c=0.018922f \
 //x=32.105 //y=5.2 //x2=31.93 //y2=6.02
cc_2766 ( N_noxref_9_M83_noxref_d N_noxref_12_M84_noxref_g ) capacitor \
 c=0.0179769f //x=31.565 //y=5.02 //x2=31.93 //y2=6.02
cc_2767 ( N_noxref_9_M19_noxref_d N_noxref_12_c_3955_n ) capacitor \
 c=0.00217566f //x=31.56 //y=0.905 //x2=31.485 //y2=0.905
cc_2768 ( N_noxref_9_M19_noxref_d N_noxref_12_c_3958_n ) capacitor \
 c=0.0034598f //x=31.56 //y=0.905 //x2=31.485 //y2=1.25
cc_2769 ( N_noxref_9_M19_noxref_d N_noxref_12_c_3960_n ) capacitor \
 c=0.00656319f //x=31.56 //y=0.905 //x2=31.485 //y2=1.56
cc_2770 ( N_noxref_9_c_3301_n N_noxref_12_c_3992_n ) capacitor c=0.0142673f \
 //x=32.19 //y=3.33 //x2=31.855 //y2=4.79
cc_2771 ( N_noxref_9_c_3383_p N_noxref_12_c_3992_n ) capacitor c=0.00407665f \
 //x=31.71 //y=5.2 //x2=31.855 //y2=4.79
cc_2772 ( N_noxref_9_M19_noxref_d N_noxref_12_c_3994_n ) capacitor \
 c=0.00241102f //x=31.56 //y=0.905 //x2=31.86 //y2=0.75
cc_2773 ( N_noxref_9_c_3300_n N_noxref_12_c_3995_n ) capacitor c=0.00359704f \
 //x=32.105 //y=1.655 //x2=31.86 //y2=1.405
cc_2774 ( N_noxref_9_M19_noxref_d N_noxref_12_c_3995_n ) capacitor \
 c=0.0138845f //x=31.56 //y=0.905 //x2=31.86 //y2=1.405
cc_2775 ( N_noxref_9_M19_noxref_d N_noxref_12_c_3963_n ) capacitor \
 c=0.00132245f //x=31.56 //y=0.905 //x2=32.015 //y2=0.905
cc_2776 ( N_noxref_9_c_3300_n N_noxref_12_c_3964_n ) capacitor c=0.00457401f \
 //x=32.105 //y=1.655 //x2=32.015 //y2=1.25
cc_2777 ( N_noxref_9_M19_noxref_d N_noxref_12_c_3964_n ) capacitor \
 c=0.00566463f //x=31.56 //y=0.905 //x2=32.015 //y2=1.25
cc_2778 ( N_noxref_9_c_3301_n N_noxref_12_c_3965_n ) capacitor c=0.00877984f \
 //x=32.19 //y=3.33 //x2=31.45 //y2=2.08
cc_2779 ( N_noxref_9_c_3301_n N_noxref_12_c_4001_n ) capacitor c=0.00306024f \
 //x=32.19 //y=3.33 //x2=31.45 //y2=1.915
cc_2780 ( N_noxref_9_M19_noxref_d N_noxref_12_c_4001_n ) capacitor \
 c=0.00660593f //x=31.56 //y=0.905 //x2=31.45 //y2=1.915
cc_2781 ( N_noxref_9_c_3316_n N_noxref_12_c_3967_n ) capacitor c=0.00346527f \
 //x=31.625 //y=5.2 //x2=31.48 //y2=4.7
cc_2782 ( N_noxref_9_c_3301_n N_noxref_12_c_3967_n ) capacitor c=0.00517969f \
 //x=32.19 //y=3.33 //x2=31.48 //y2=4.7
cc_2783 ( N_noxref_9_M86_noxref_g N_noxref_12_M85_noxref_d ) capacitor \
 c=0.0173476f //x=34.38 //y=6.02 //x2=34.015 //y2=5.02
cc_2784 ( N_noxref_9_c_3355_p N_D_c_4238_n ) capacitor c=0.0125396f //x=33.925 \
 //y=3.33 //x2=49.465 //y2=2.59
cc_2785 ( N_noxref_9_c_3347_n N_D_c_4238_n ) capacitor c=8.92472e-19 \
 //x=32.305 //y=3.33 //x2=49.465 //y2=2.59
cc_2786 ( N_noxref_9_c_3398_p N_D_c_4238_n ) capacitor c=0.0102711f //x=31.835 \
 //y=1.655 //x2=49.465 //y2=2.59
cc_2787 ( N_noxref_9_c_3301_n N_D_c_4238_n ) capacitor c=0.0210598f //x=32.19 \
 //y=3.33 //x2=49.465 //y2=2.59
cc_2788 ( N_noxref_9_c_3302_n N_D_c_4238_n ) capacitor c=0.0213243f //x=34.04 \
 //y=2.08 //x2=49.465 //y2=2.59
cc_2789 ( N_noxref_9_c_3307_n N_D_c_4238_n ) capacitor c=0.0052136f //x=33.845 \
 //y=1.915 //x2=49.465 //y2=2.59
cc_2790 ( N_noxref_9_c_3316_n N_CLK_c_5061_n ) capacitor c=0.0185297f \
 //x=31.625 //y=5.2 //x2=34.665 //y2=4.44
cc_2791 ( N_noxref_9_c_3320_n N_CLK_c_5061_n ) capacitor c=0.018142f \
 //x=30.915 //y=5.2 //x2=34.665 //y2=4.44
cc_2792 ( N_noxref_9_c_3301_n N_CLK_c_5061_n ) capacitor c=0.0208321f \
 //x=32.19 //y=3.33 //x2=34.665 //y2=4.44
cc_2793 ( N_noxref_9_c_3302_n N_CLK_c_5061_n ) capacitor c=0.0198304f \
 //x=34.04 //y=2.08 //x2=34.665 //y2=4.44
cc_2794 ( N_noxref_9_c_3335_n N_CLK_c_5061_n ) capacitor c=0.0107057f \
 //x=34.04 //y=4.7 //x2=34.665 //y2=4.44
cc_2795 ( N_noxref_9_c_3302_n N_CLK_c_5111_n ) capacitor c=0.00168329f \
 //x=34.04 //y=2.08 //x2=34.895 //y2=4.44
cc_2796 ( N_noxref_9_c_3335_n N_CLK_c_5111_n ) capacitor c=2.91071e-19 \
 //x=34.04 //y=4.7 //x2=34.895 //y2=4.44
cc_2797 ( N_noxref_9_c_3302_n N_CLK_c_5363_n ) capacitor c=0.00400249f \
 //x=34.04 //y=2.08 //x2=34.78 //y2=4.535
cc_2798 ( N_noxref_9_c_3335_n N_CLK_c_5363_n ) capacitor c=0.00415951f \
 //x=34.04 //y=4.7 //x2=34.78 //y2=4.535
cc_2799 ( N_noxref_9_c_3355_p N_CLK_c_5029_n ) capacitor c=0.00720056f \
 //x=33.925 //y=3.33 //x2=34.78 //y2=2.08
cc_2800 ( N_noxref_9_c_3301_n N_CLK_c_5029_n ) capacitor c=9.02527e-19 \
 //x=32.19 //y=3.33 //x2=34.78 //y2=2.08
cc_2801 ( N_noxref_9_c_3302_n N_CLK_c_5029_n ) capacitor c=0.0735625f \
 //x=34.04 //y=2.08 //x2=34.78 //y2=2.08
cc_2802 ( N_noxref_9_c_3307_n N_CLK_c_5029_n ) capacitor c=0.00308814f \
 //x=33.845 //y=1.915 //x2=34.78 //y2=2.08
cc_2803 ( N_noxref_9_M85_noxref_g N_CLK_M87_noxref_g ) capacitor c=0.0104611f \
 //x=33.94 //y=6.02 //x2=34.82 //y2=6.02
cc_2804 ( N_noxref_9_M86_noxref_g N_CLK_M87_noxref_g ) capacitor c=0.106811f \
 //x=34.38 //y=6.02 //x2=34.82 //y2=6.02
cc_2805 ( N_noxref_9_M86_noxref_g N_CLK_M88_noxref_g ) capacitor c=0.0100341f \
 //x=34.38 //y=6.02 //x2=35.26 //y2=6.02
cc_2806 ( N_noxref_9_c_3303_n N_CLK_c_5372_n ) capacitor c=4.86506e-19 \
 //x=33.845 //y=0.865 //x2=34.815 //y2=0.905
cc_2807 ( N_noxref_9_c_3305_n N_CLK_c_5372_n ) capacitor c=0.00152104f \
 //x=33.845 //y=1.21 //x2=34.815 //y2=0.905
cc_2808 ( N_noxref_9_c_3310_n N_CLK_c_5372_n ) capacitor c=0.0151475f \
 //x=34.375 //y=0.865 //x2=34.815 //y2=0.905
cc_2809 ( N_noxref_9_c_3306_n N_CLK_c_5375_n ) capacitor c=0.00109982f \
 //x=33.845 //y=1.52 //x2=34.815 //y2=1.25
cc_2810 ( N_noxref_9_c_3312_n N_CLK_c_5375_n ) capacitor c=0.0111064f \
 //x=34.375 //y=1.21 //x2=34.815 //y2=1.25
cc_2811 ( N_noxref_9_c_3306_n N_CLK_c_5377_n ) capacitor c=9.57794e-19 \
 //x=33.845 //y=1.52 //x2=34.815 //y2=1.56
cc_2812 ( N_noxref_9_c_3307_n N_CLK_c_5377_n ) capacitor c=0.00662747f \
 //x=33.845 //y=1.915 //x2=34.815 //y2=1.56
cc_2813 ( N_noxref_9_c_3312_n N_CLK_c_5377_n ) capacitor c=0.00862358f \
 //x=34.375 //y=1.21 //x2=34.815 //y2=1.56
cc_2814 ( N_noxref_9_c_3310_n N_CLK_c_5380_n ) capacitor c=0.00124821f \
 //x=34.375 //y=0.865 //x2=35.345 //y2=0.905
cc_2815 ( N_noxref_9_c_3312_n N_CLK_c_5381_n ) capacitor c=0.00200715f \
 //x=34.375 //y=1.21 //x2=35.345 //y2=1.25
cc_2816 ( N_noxref_9_c_3302_n N_CLK_c_5382_n ) capacitor c=0.00307062f \
 //x=34.04 //y=2.08 //x2=34.78 //y2=2.08
cc_2817 ( N_noxref_9_c_3307_n N_CLK_c_5382_n ) capacitor c=0.0179092f \
 //x=33.845 //y=1.915 //x2=34.78 //y2=2.08
cc_2818 ( N_noxref_9_c_3302_n N_CLK_c_5384_n ) capacitor c=0.00342116f \
 //x=34.04 //y=2.08 //x2=34.81 //y2=4.7
cc_2819 ( N_noxref_9_c_3335_n N_CLK_c_5384_n ) capacitor c=0.0292158f \
 //x=34.04 //y=4.7 //x2=34.81 //y2=4.7
cc_2820 ( N_noxref_9_c_3355_p N_noxref_23_c_7498_n ) capacitor c=0.173509f \
 //x=33.925 //y=3.33 //x2=70.185 //y2=2.96
cc_2821 ( N_noxref_9_c_3347_n N_noxref_23_c_7498_n ) capacitor c=0.0292689f \
 //x=32.305 //y=3.33 //x2=70.185 //y2=2.96
cc_2822 ( N_noxref_9_c_3301_n N_noxref_23_c_7498_n ) capacitor c=0.0206014f \
 //x=32.19 //y=3.33 //x2=70.185 //y2=2.96
cc_2823 ( N_noxref_9_c_3302_n N_noxref_23_c_7498_n ) capacitor c=0.0205758f \
 //x=34.04 //y=2.08 //x2=70.185 //y2=2.96
cc_2824 ( N_noxref_9_c_3398_p N_noxref_36_c_8752_n ) capacitor c=3.15806e-19 \
 //x=31.835 //y=1.655 //x2=30.295 //y2=1.495
cc_2825 ( N_noxref_9_c_3398_p N_noxref_36_c_8740_n ) capacitor c=0.0203424f \
 //x=31.835 //y=1.655 //x2=31.265 //y2=1.495
cc_2826 ( N_noxref_9_c_3300_n N_noxref_36_c_8741_n ) capacitor c=0.00461444f \
 //x=32.105 //y=1.655 //x2=32.15 //y2=0.53
cc_2827 ( N_noxref_9_M19_noxref_d N_noxref_36_c_8741_n ) capacitor \
 c=0.0116735f //x=31.56 //y=0.905 //x2=32.15 //y2=0.53
cc_2828 ( N_noxref_9_c_3300_n N_noxref_36_M18_noxref_s ) capacitor \
 c=0.0137901f //x=32.105 //y=1.655 //x2=30.16 //y2=0.365
cc_2829 ( N_noxref_9_M19_noxref_d N_noxref_36_M18_noxref_s ) capacitor \
 c=0.043966f //x=31.56 //y=0.905 //x2=30.16 //y2=0.365
cc_2830 ( N_noxref_9_c_3300_n N_noxref_37_c_8804_n ) capacitor c=3.22188e-19 \
 //x=32.105 //y=1.655 //x2=33.625 //y2=1.495
cc_2831 ( N_noxref_9_c_3307_n N_noxref_37_c_8804_n ) capacitor c=0.0034165f \
 //x=33.845 //y=1.915 //x2=33.625 //y2=1.495
cc_2832 ( N_noxref_9_c_3302_n N_noxref_37_c_8785_n ) capacitor c=0.0118762f \
 //x=34.04 //y=2.08 //x2=34.51 //y2=1.58
cc_2833 ( N_noxref_9_c_3306_n N_noxref_37_c_8785_n ) capacitor c=0.00703567f \
 //x=33.845 //y=1.52 //x2=34.51 //y2=1.58
cc_2834 ( N_noxref_9_c_3307_n N_noxref_37_c_8785_n ) capacitor c=0.018562f \
 //x=33.845 //y=1.915 //x2=34.51 //y2=1.58
cc_2835 ( N_noxref_9_c_3309_n N_noxref_37_c_8785_n ) capacitor c=0.00780629f \
 //x=34.22 //y=1.365 //x2=34.51 //y2=1.58
cc_2836 ( N_noxref_9_c_3312_n N_noxref_37_c_8785_n ) capacitor c=0.00339872f \
 //x=34.375 //y=1.21 //x2=34.51 //y2=1.58
cc_2837 ( N_noxref_9_c_3307_n N_noxref_37_c_8792_n ) capacitor c=6.71402e-19 \
 //x=33.845 //y=1.915 //x2=34.595 //y2=1.495
cc_2838 ( N_noxref_9_c_3303_n N_noxref_37_M20_noxref_s ) capacitor \
 c=0.0326577f //x=33.845 //y=0.865 //x2=33.49 //y2=0.365
cc_2839 ( N_noxref_9_c_3306_n N_noxref_37_M20_noxref_s ) capacitor \
 c=3.48408e-19 //x=33.845 //y=1.52 //x2=33.49 //y2=0.365
cc_2840 ( N_noxref_9_c_3310_n N_noxref_37_M20_noxref_s ) capacitor \
 c=0.0120759f //x=34.375 //y=0.865 //x2=33.49 //y2=0.365
cc_2841 ( N_noxref_10_c_3526_n N_noxref_11_c_3758_n ) capacitor c=0.0114735f \
 //x=37.255 //y=3.7 //x2=38.965 //y2=3.7
cc_2842 ( N_noxref_10_M90_noxref_g N_noxref_11_c_3727_n ) capacitor \
 c=0.0169521f //x=37.71 //y=6.02 //x2=38.285 //y2=5.2
cc_2843 ( N_noxref_10_c_3455_n N_noxref_11_c_3731_n ) capacitor c=0.00521572f \
 //x=37.37 //y=2.08 //x2=37.575 //y2=5.2
cc_2844 ( N_noxref_10_M89_noxref_g N_noxref_11_c_3731_n ) capacitor \
 c=0.0177326f //x=37.27 //y=6.02 //x2=37.575 //y2=5.2
cc_2845 ( N_noxref_10_c_3507_n N_noxref_11_c_3731_n ) capacitor c=0.00581252f \
 //x=37.37 //y=4.7 //x2=37.575 //y2=5.2
cc_2846 ( N_noxref_10_c_3455_n N_noxref_11_c_3712_n ) capacitor c=0.00281709f \
 //x=37.37 //y=2.08 //x2=38.85 //y2=3.7
cc_2847 ( N_noxref_10_M90_noxref_g N_noxref_11_M89_noxref_d ) capacitor \
 c=0.0173476f //x=37.71 //y=6.02 //x2=37.345 //y2=5.02
cc_2848 ( N_noxref_10_c_3523_n N_noxref_12_c_3882_n ) capacitor c=0.147021f \
 //x=27.265 //y=3.7 //x2=31.335 //y2=4.07
cc_2849 ( N_noxref_10_c_3524_n N_noxref_12_c_3882_n ) capacitor c=0.0294294f \
 //x=25.645 //y=3.7 //x2=31.335 //y2=4.07
cc_2850 ( N_noxref_10_c_3526_n N_noxref_12_c_3882_n ) capacitor c=0.338937f \
 //x=37.255 //y=3.7 //x2=31.335 //y2=4.07
cc_2851 ( N_noxref_10_c_3531_n N_noxref_12_c_3882_n ) capacitor c=0.0264478f \
 //x=27.495 //y=3.7 //x2=31.335 //y2=4.07
cc_2852 ( N_noxref_10_c_3491_n N_noxref_12_c_3882_n ) capacitor c=0.0200328f \
 //x=25.53 //y=3.7 //x2=31.335 //y2=4.07
cc_2853 ( N_noxref_10_c_3454_n N_noxref_12_c_3882_n ) capacitor c=0.0203111f \
 //x=27.38 //y=2.08 //x2=31.335 //y2=4.07
cc_2854 ( N_noxref_10_c_3526_n N_noxref_12_c_3885_n ) capacitor c=0.339146f \
 //x=37.255 //y=3.7 //x2=35.405 //y2=4.07
cc_2855 ( N_noxref_10_c_3526_n N_noxref_12_c_3944_n ) capacitor c=0.0267832f \
 //x=37.255 //y=3.7 //x2=31.565 //y2=4.07
cc_2856 ( N_noxref_10_c_3526_n N_noxref_12_c_3886_n ) capacitor c=0.176049f \
 //x=37.255 //y=3.7 //x2=41.325 //y2=4.07
cc_2857 ( N_noxref_10_c_3455_n N_noxref_12_c_3886_n ) capacitor c=0.0202919f \
 //x=37.37 //y=2.08 //x2=41.325 //y2=4.07
cc_2858 ( N_noxref_10_c_3526_n N_noxref_12_c_3888_n ) capacitor c=0.0266833f \
 //x=37.255 //y=3.7 //x2=35.635 //y2=4.07
cc_2859 ( N_noxref_10_c_3455_n N_noxref_12_c_3888_n ) capacitor c=3.50683e-19 \
 //x=37.37 //y=2.08 //x2=35.635 //y2=4.07
cc_2860 ( N_noxref_10_c_3526_n N_noxref_12_c_3863_n ) capacitor c=0.0211371f \
 //x=37.255 //y=3.7 //x2=31.45 //y2=2.08
cc_2861 ( N_noxref_10_c_3526_n N_noxref_12_c_3866_n ) capacitor c=0.0235138f \
 //x=37.255 //y=3.7 //x2=35.52 //y2=4.07
cc_2862 ( N_noxref_10_c_3455_n N_noxref_12_c_3866_n ) capacitor c=0.0125822f \
 //x=37.37 //y=2.08 //x2=35.52 //y2=4.07
cc_2863 ( N_noxref_10_c_3481_n N_noxref_12_M71_noxref_g ) capacitor \
 c=0.0213876f //x=23.075 //y=5.155 //x2=22.77 //y2=6.02
cc_2864 ( N_noxref_10_c_3477_n N_noxref_12_M72_noxref_g ) capacitor \
 c=0.0168349f //x=23.785 //y=5.155 //x2=23.21 //y2=6.02
cc_2865 ( N_noxref_10_M71_noxref_d N_noxref_12_M72_noxref_g ) capacitor \
 c=0.0180032f //x=22.845 //y=5.02 //x2=23.21 //y2=6.02
cc_2866 ( N_noxref_10_c_3481_n N_noxref_12_c_4024_n ) capacitor c=0.00428486f \
 //x=23.075 //y=5.155 //x2=23.135 //y2=4.79
cc_2867 ( N_noxref_10_c_3594_p N_D_c_4217_n ) capacitor c=0.0115788f //x=25.13 \
 //y=1.665 //x2=28.005 //y2=2.59
cc_2868 ( N_noxref_10_c_3491_n N_D_c_4217_n ) capacitor c=0.0209737f //x=25.53 \
 //y=3.7 //x2=28.005 //y2=2.59
cc_2869 ( N_noxref_10_c_3454_n N_D_c_4217_n ) capacitor c=0.0213243f //x=27.38 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_2870 ( N_noxref_10_c_3460_n N_D_c_4217_n ) capacitor c=0.0052136f \
 //x=27.185 //y=1.915 //x2=28.005 //y2=2.59
cc_2871 ( N_noxref_10_c_3526_n N_D_c_4238_n ) capacitor c=0.023303f //x=37.255 \
 //y=3.7 //x2=49.465 //y2=2.59
cc_2872 ( N_noxref_10_c_3455_n N_D_c_4238_n ) capacitor c=0.0213243f //x=37.37 \
 //y=2.08 //x2=49.465 //y2=2.59
cc_2873 ( N_noxref_10_c_3470_n N_D_c_4238_n ) capacitor c=0.0052136f \
 //x=37.175 //y=1.915 //x2=49.465 //y2=2.59
cc_2874 ( N_noxref_10_c_3454_n N_D_c_4251_n ) capacitor c=0.00179385f \
 //x=27.38 //y=2.08 //x2=28.235 //y2=2.59
cc_2875 ( N_noxref_10_c_3454_n N_D_c_4381_n ) capacitor c=0.00400249f \
 //x=27.38 //y=2.08 //x2=28.12 //y2=4.535
cc_2876 ( N_noxref_10_c_3506_n N_D_c_4381_n ) capacitor c=0.00417994f \
 //x=27.38 //y=4.7 //x2=28.12 //y2=4.535
cc_2877 ( N_noxref_10_c_3526_n N_D_c_4255_n ) capacitor c=0.0169594f \
 //x=37.255 //y=3.7 //x2=28.12 //y2=2.08
cc_2878 ( N_noxref_10_c_3531_n N_D_c_4255_n ) capacitor c=0.00131333f \
 //x=27.495 //y=3.7 //x2=28.12 //y2=2.08
cc_2879 ( N_noxref_10_c_3491_n N_D_c_4255_n ) capacitor c=6.91957e-19 \
 //x=25.53 //y=3.7 //x2=28.12 //y2=2.08
cc_2880 ( N_noxref_10_c_3454_n N_D_c_4255_n ) capacitor c=0.0729553f //x=27.38 \
 //y=2.08 //x2=28.12 //y2=2.08
cc_2881 ( N_noxref_10_c_3460_n N_D_c_4255_n ) capacitor c=0.00308814f \
 //x=27.185 //y=1.915 //x2=28.12 //y2=2.08
cc_2882 ( N_noxref_10_M77_noxref_g N_D_M79_noxref_g ) capacitor c=0.0104611f \
 //x=27.28 //y=6.02 //x2=28.16 //y2=6.02
cc_2883 ( N_noxref_10_M78_noxref_g N_D_M79_noxref_g ) capacitor c=0.106811f \
 //x=27.72 //y=6.02 //x2=28.16 //y2=6.02
cc_2884 ( N_noxref_10_M78_noxref_g N_D_M80_noxref_g ) capacitor c=0.0100341f \
 //x=27.72 //y=6.02 //x2=28.6 //y2=6.02
cc_2885 ( N_noxref_10_c_3456_n N_D_c_4391_n ) capacitor c=4.86506e-19 \
 //x=27.185 //y=0.865 //x2=28.155 //y2=0.905
cc_2886 ( N_noxref_10_c_3458_n N_D_c_4391_n ) capacitor c=0.00152104f \
 //x=27.185 //y=1.21 //x2=28.155 //y2=0.905
cc_2887 ( N_noxref_10_c_3463_n N_D_c_4391_n ) capacitor c=0.0151475f \
 //x=27.715 //y=0.865 //x2=28.155 //y2=0.905
cc_2888 ( N_noxref_10_c_3459_n N_D_c_4392_n ) capacitor c=0.00109982f \
 //x=27.185 //y=1.52 //x2=28.155 //y2=1.25
cc_2889 ( N_noxref_10_c_3465_n N_D_c_4392_n ) capacitor c=0.0111064f \
 //x=27.715 //y=1.21 //x2=28.155 //y2=1.25
cc_2890 ( N_noxref_10_c_3459_n N_D_c_4393_n ) capacitor c=9.57794e-19 \
 //x=27.185 //y=1.52 //x2=28.155 //y2=1.56
cc_2891 ( N_noxref_10_c_3460_n N_D_c_4393_n ) capacitor c=0.00662747f \
 //x=27.185 //y=1.915 //x2=28.155 //y2=1.56
cc_2892 ( N_noxref_10_c_3465_n N_D_c_4393_n ) capacitor c=0.00862358f \
 //x=27.715 //y=1.21 //x2=28.155 //y2=1.56
cc_2893 ( N_noxref_10_c_3463_n N_D_c_4399_n ) capacitor c=0.00124821f \
 //x=27.715 //y=0.865 //x2=28.685 //y2=0.905
cc_2894 ( N_noxref_10_c_3465_n N_D_c_4400_n ) capacitor c=0.00200715f \
 //x=27.715 //y=1.21 //x2=28.685 //y2=1.25
cc_2895 ( N_noxref_10_c_3454_n N_D_c_4402_n ) capacitor c=0.00307062f \
 //x=27.38 //y=2.08 //x2=28.12 //y2=2.08
cc_2896 ( N_noxref_10_c_3460_n N_D_c_4402_n ) capacitor c=0.0179092f \
 //x=27.185 //y=1.915 //x2=28.12 //y2=2.08
cc_2897 ( N_noxref_10_c_3454_n N_D_c_4405_n ) capacitor c=0.00344981f \
 //x=27.38 //y=2.08 //x2=28.15 //y2=4.7
cc_2898 ( N_noxref_10_c_3506_n N_D_c_4405_n ) capacitor c=0.0293367f //x=27.38 \
 //y=4.7 //x2=28.15 //y2=4.7
cc_2899 ( N_noxref_10_c_3523_n N_CLK_c_5061_n ) capacitor c=0.00940379f \
 //x=27.265 //y=3.7 //x2=34.665 //y2=4.44
cc_2900 ( N_noxref_10_c_3524_n N_CLK_c_5061_n ) capacitor c=7.95009e-19 \
 //x=25.645 //y=3.7 //x2=34.665 //y2=4.44
cc_2901 ( N_noxref_10_c_3526_n N_CLK_c_5061_n ) capacitor c=0.0485341f \
 //x=37.255 //y=3.7 //x2=34.665 //y2=4.44
cc_2902 ( N_noxref_10_c_3531_n N_CLK_c_5061_n ) capacitor c=6.59192e-19 \
 //x=27.495 //y=3.7 //x2=34.665 //y2=4.44
cc_2903 ( N_noxref_10_c_3487_n N_CLK_c_5061_n ) capacitor c=0.0183122f \
 //x=25.445 //y=5.155 //x2=34.665 //y2=4.44
cc_2904 ( N_noxref_10_c_3491_n N_CLK_c_5061_n ) capacitor c=0.0210274f \
 //x=25.53 //y=3.7 //x2=34.665 //y2=4.44
cc_2905 ( N_noxref_10_c_3454_n N_CLK_c_5061_n ) capacitor c=0.0198304f \
 //x=27.38 //y=2.08 //x2=34.665 //y2=4.44
cc_2906 ( N_noxref_10_c_3633_p N_CLK_c_5061_n ) capacitor c=0.0311227f \
 //x=23.87 //y=5.155 //x2=34.665 //y2=4.44
cc_2907 ( N_noxref_10_c_3506_n N_CLK_c_5061_n ) capacitor c=0.0107057f \
 //x=27.38 //y=4.7 //x2=34.665 //y2=4.44
cc_2908 ( N_noxref_10_c_3477_n N_CLK_c_5079_n ) capacitor c=0.00241768f \
 //x=23.785 //y=5.155 //x2=23.795 //y2=4.44
cc_2909 ( N_noxref_10_c_3481_n N_CLK_c_5079_n ) capacitor c=0.0219242f \
 //x=23.075 //y=5.155 //x2=23.795 //y2=4.44
cc_2910 ( N_noxref_10_c_3526_n N_CLK_c_5092_n ) capacitor c=0.0160726f \
 //x=37.255 //y=3.7 //x2=45.025 //y2=4.44
cc_2911 ( N_noxref_10_c_3455_n N_CLK_c_5092_n ) capacitor c=0.0198304f \
 //x=37.37 //y=2.08 //x2=45.025 //y2=4.44
cc_2912 ( N_noxref_10_c_3507_n N_CLK_c_5092_n ) capacitor c=0.0107057f \
 //x=37.37 //y=4.7 //x2=45.025 //y2=4.44
cc_2913 ( N_noxref_10_c_3526_n N_CLK_c_5111_n ) capacitor c=5.12294e-19 \
 //x=37.255 //y=3.7 //x2=34.895 //y2=4.44
cc_2914 ( N_noxref_10_c_3477_n N_CLK_c_5028_n ) capacitor c=0.0143918f \
 //x=23.785 //y=5.155 //x2=23.68 //y2=2.08
cc_2915 ( N_noxref_10_c_3491_n N_CLK_c_5028_n ) capacitor c=0.00288484f \
 //x=25.53 //y=3.7 //x2=23.68 //y2=2.08
cc_2916 ( N_noxref_10_c_3526_n N_CLK_c_5029_n ) capacitor c=0.0193001f \
 //x=37.255 //y=3.7 //x2=34.78 //y2=2.08
cc_2917 ( N_noxref_10_c_3455_n N_CLK_c_5029_n ) capacitor c=8.90899e-19 \
 //x=37.37 //y=2.08 //x2=34.78 //y2=2.08
cc_2918 ( N_noxref_10_c_3477_n N_CLK_M73_noxref_g ) capacitor c=0.016514f \
 //x=23.785 //y=5.155 //x2=23.65 //y2=6.02
cc_2919 ( N_noxref_10_M73_noxref_d N_CLK_M73_noxref_g ) capacitor c=0.0180032f \
 //x=23.725 //y=5.02 //x2=23.65 //y2=6.02
cc_2920 ( N_noxref_10_c_3483_n N_CLK_M74_noxref_g ) capacitor c=0.01736f \
 //x=24.665 //y=5.155 //x2=24.09 //y2=6.02
cc_2921 ( N_noxref_10_M73_noxref_d N_CLK_M74_noxref_g ) capacitor c=0.0180032f \
 //x=23.725 //y=5.02 //x2=24.09 //y2=6.02
cc_2922 ( N_noxref_10_c_3633_p N_CLK_c_5353_n ) capacitor c=0.00426767f \
 //x=23.87 //y=5.155 //x2=24.015 //y2=4.79
cc_2923 ( N_noxref_10_c_3477_n N_CLK_c_5354_n ) capacitor c=0.00322046f \
 //x=23.785 //y=5.155 //x2=23.68 //y2=4.7
cc_2924 ( N_noxref_10_c_3455_n N_noxref_21_c_6909_n ) capacitor c=0.00689524f \
 //x=37.37 //y=2.08 //x2=38.225 //y2=2.22
cc_2925 ( N_noxref_10_c_3470_n N_noxref_21_c_6909_n ) capacitor c=0.00226803f \
 //x=37.175 //y=1.915 //x2=38.225 //y2=2.22
cc_2926 ( N_noxref_10_c_3455_n N_noxref_21_c_7001_n ) capacitor c=0.00400249f \
 //x=37.37 //y=2.08 //x2=38.11 //y2=4.535
cc_2927 ( N_noxref_10_c_3507_n N_noxref_21_c_7001_n ) capacitor c=0.00417994f \
 //x=37.37 //y=4.7 //x2=38.11 //y2=4.535
cc_2928 ( N_noxref_10_c_3526_n N_noxref_21_c_6939_n ) capacitor c=0.00318578f \
 //x=37.255 //y=3.7 //x2=38.11 //y2=2.08
cc_2929 ( N_noxref_10_c_3455_n N_noxref_21_c_6939_n ) capacitor c=0.0750332f \
 //x=37.37 //y=2.08 //x2=38.11 //y2=2.08
cc_2930 ( N_noxref_10_c_3470_n N_noxref_21_c_6939_n ) capacitor c=0.00296726f \
 //x=37.175 //y=1.915 //x2=38.11 //y2=2.08
cc_2931 ( N_noxref_10_M89_noxref_g N_noxref_21_M91_noxref_g ) capacitor \
 c=0.0104611f //x=37.27 //y=6.02 //x2=38.15 //y2=6.02
cc_2932 ( N_noxref_10_M90_noxref_g N_noxref_21_M91_noxref_g ) capacitor \
 c=0.106811f //x=37.71 //y=6.02 //x2=38.15 //y2=6.02
cc_2933 ( N_noxref_10_M90_noxref_g N_noxref_21_M92_noxref_g ) capacitor \
 c=0.0100341f //x=37.71 //y=6.02 //x2=38.59 //y2=6.02
cc_2934 ( N_noxref_10_c_3466_n N_noxref_21_c_7009_n ) capacitor c=4.86506e-19 \
 //x=37.175 //y=0.865 //x2=38.145 //y2=0.905
cc_2935 ( N_noxref_10_c_3468_n N_noxref_21_c_7009_n ) capacitor c=0.00152104f \
 //x=37.175 //y=1.21 //x2=38.145 //y2=0.905
cc_2936 ( N_noxref_10_c_3473_n N_noxref_21_c_7009_n ) capacitor c=0.0151475f \
 //x=37.705 //y=0.865 //x2=38.145 //y2=0.905
cc_2937 ( N_noxref_10_c_3469_n N_noxref_21_c_7012_n ) capacitor c=0.00109982f \
 //x=37.175 //y=1.52 //x2=38.145 //y2=1.25
cc_2938 ( N_noxref_10_c_3475_n N_noxref_21_c_7012_n ) capacitor c=0.0111064f \
 //x=37.705 //y=1.21 //x2=38.145 //y2=1.25
cc_2939 ( N_noxref_10_c_3469_n N_noxref_21_c_7014_n ) capacitor c=9.57794e-19 \
 //x=37.175 //y=1.52 //x2=38.145 //y2=1.56
cc_2940 ( N_noxref_10_c_3470_n N_noxref_21_c_7014_n ) capacitor c=0.00662747f \
 //x=37.175 //y=1.915 //x2=38.145 //y2=1.56
cc_2941 ( N_noxref_10_c_3475_n N_noxref_21_c_7014_n ) capacitor c=0.00862358f \
 //x=37.705 //y=1.21 //x2=38.145 //y2=1.56
cc_2942 ( N_noxref_10_c_3473_n N_noxref_21_c_7017_n ) capacitor c=0.00124821f \
 //x=37.705 //y=0.865 //x2=38.675 //y2=0.905
cc_2943 ( N_noxref_10_c_3475_n N_noxref_21_c_7018_n ) capacitor c=0.00200715f \
 //x=37.705 //y=1.21 //x2=38.675 //y2=1.25
cc_2944 ( N_noxref_10_c_3455_n N_noxref_21_c_7019_n ) capacitor c=0.00291775f \
 //x=37.37 //y=2.08 //x2=38.11 //y2=2.08
cc_2945 ( N_noxref_10_c_3470_n N_noxref_21_c_7019_n ) capacitor c=0.0174866f \
 //x=37.175 //y=1.915 //x2=38.11 //y2=2.08
cc_2946 ( N_noxref_10_c_3455_n N_noxref_21_c_7021_n ) capacitor c=0.00344981f \
 //x=37.37 //y=2.08 //x2=38.14 //y2=4.7
cc_2947 ( N_noxref_10_c_3507_n N_noxref_21_c_7021_n ) capacitor c=0.0293367f \
 //x=37.37 //y=4.7 //x2=38.14 //y2=4.7
cc_2948 ( N_noxref_10_c_3523_n N_noxref_23_c_7498_n ) capacitor c=0.0110781f \
 //x=27.265 //y=3.7 //x2=70.185 //y2=2.96
cc_2949 ( N_noxref_10_c_3524_n N_noxref_23_c_7498_n ) capacitor c=7.98411e-19 \
 //x=25.645 //y=3.7 //x2=70.185 //y2=2.96
cc_2950 ( N_noxref_10_c_3526_n N_noxref_23_c_7498_n ) capacitor c=0.232839f \
 //x=37.255 //y=3.7 //x2=70.185 //y2=2.96
cc_2951 ( N_noxref_10_c_3531_n N_noxref_23_c_7498_n ) capacitor c=5.76555e-19 \
 //x=27.495 //y=3.7 //x2=70.185 //y2=2.96
cc_2952 ( N_noxref_10_c_3491_n N_noxref_23_c_7498_n ) capacitor c=0.0187656f \
 //x=25.53 //y=3.7 //x2=70.185 //y2=2.96
cc_2953 ( N_noxref_10_c_3454_n N_noxref_23_c_7498_n ) capacitor c=0.0187412f \
 //x=27.38 //y=2.08 //x2=70.185 //y2=2.96
cc_2954 ( N_noxref_10_c_3455_n N_noxref_23_c_7498_n ) capacitor c=0.0213728f \
 //x=37.37 //y=2.08 //x2=70.185 //y2=2.96
cc_2955 ( N_noxref_10_c_3481_n N_noxref_23_c_7518_n ) capacitor c=2.97874e-19 \
 //x=23.075 //y=5.155 //x2=20.72 //y2=2.96
cc_2956 ( N_noxref_10_M15_noxref_d N_noxref_33_M13_noxref_s ) capacitor \
 c=0.00309936f //x=24.855 //y=0.915 //x2=21.915 //y2=0.375
cc_2957 ( N_noxref_10_c_3453_n N_noxref_34_c_8631_n ) capacitor c=0.00461497f \
 //x=25.445 //y=1.665 //x2=25.445 //y2=0.54
cc_2958 ( N_noxref_10_M15_noxref_d N_noxref_34_c_8631_n ) capacitor \
 c=0.0116817f //x=24.855 //y=0.915 //x2=25.445 //y2=0.54
cc_2959 ( N_noxref_10_c_3594_p N_noxref_34_c_8644_n ) capacitor c=0.020048f \
 //x=25.13 //y=1.665 //x2=24.56 //y2=0.995
cc_2960 ( N_noxref_10_M15_noxref_d N_noxref_34_M14_noxref_d ) capacitor \
 c=5.27807e-19 //x=24.855 //y=0.915 //x2=23.32 //y2=0.91
cc_2961 ( N_noxref_10_c_3453_n N_noxref_34_M15_noxref_s ) capacitor \
 c=0.0201579f //x=25.445 //y=1.665 //x2=24.425 //y2=0.375
cc_2962 ( N_noxref_10_M15_noxref_d N_noxref_34_M15_noxref_s ) capacitor \
 c=0.0426444f //x=24.855 //y=0.915 //x2=24.425 //y2=0.375
cc_2963 ( N_noxref_10_c_3453_n N_noxref_35_c_8698_n ) capacitor c=3.04182e-19 \
 //x=25.445 //y=1.665 //x2=26.965 //y2=1.495
cc_2964 ( N_noxref_10_c_3460_n N_noxref_35_c_8698_n ) capacitor c=0.0034165f \
 //x=27.185 //y=1.915 //x2=26.965 //y2=1.495
cc_2965 ( N_noxref_10_c_3454_n N_noxref_35_c_8679_n ) capacitor c=0.0118762f \
 //x=27.38 //y=2.08 //x2=27.85 //y2=1.58
cc_2966 ( N_noxref_10_c_3459_n N_noxref_35_c_8679_n ) capacitor c=0.00703567f \
 //x=27.185 //y=1.52 //x2=27.85 //y2=1.58
cc_2967 ( N_noxref_10_c_3460_n N_noxref_35_c_8679_n ) capacitor c=0.018562f \
 //x=27.185 //y=1.915 //x2=27.85 //y2=1.58
cc_2968 ( N_noxref_10_c_3462_n N_noxref_35_c_8679_n ) capacitor c=0.00780629f \
 //x=27.56 //y=1.365 //x2=27.85 //y2=1.58
cc_2969 ( N_noxref_10_c_3465_n N_noxref_35_c_8679_n ) capacitor c=0.00339872f \
 //x=27.715 //y=1.21 //x2=27.85 //y2=1.58
cc_2970 ( N_noxref_10_c_3460_n N_noxref_35_c_8686_n ) capacitor c=6.71402e-19 \
 //x=27.185 //y=1.915 //x2=27.935 //y2=1.495
cc_2971 ( N_noxref_10_c_3456_n N_noxref_35_M16_noxref_s ) capacitor \
 c=0.0327502f //x=27.185 //y=0.865 //x2=26.83 //y2=0.365
cc_2972 ( N_noxref_10_c_3459_n N_noxref_35_M16_noxref_s ) capacitor \
 c=3.48408e-19 //x=27.185 //y=1.52 //x2=26.83 //y2=0.365
cc_2973 ( N_noxref_10_c_3463_n N_noxref_35_M16_noxref_s ) capacitor \
 c=0.0120759f //x=27.715 //y=0.865 //x2=26.83 //y2=0.365
cc_2974 ( N_noxref_10_c_3470_n N_noxref_38_c_8856_n ) capacitor c=0.0034165f \
 //x=37.175 //y=1.915 //x2=36.955 //y2=1.495
cc_2975 ( N_noxref_10_c_3455_n N_noxref_38_c_8837_n ) capacitor c=0.0118762f \
 //x=37.37 //y=2.08 //x2=37.84 //y2=1.58
cc_2976 ( N_noxref_10_c_3469_n N_noxref_38_c_8837_n ) capacitor c=0.00703567f \
 //x=37.175 //y=1.52 //x2=37.84 //y2=1.58
cc_2977 ( N_noxref_10_c_3470_n N_noxref_38_c_8837_n ) capacitor c=0.018562f \
 //x=37.175 //y=1.915 //x2=37.84 //y2=1.58
cc_2978 ( N_noxref_10_c_3472_n N_noxref_38_c_8837_n ) capacitor c=0.00780629f \
 //x=37.55 //y=1.365 //x2=37.84 //y2=1.58
cc_2979 ( N_noxref_10_c_3475_n N_noxref_38_c_8837_n ) capacitor c=0.00339872f \
 //x=37.705 //y=1.21 //x2=37.84 //y2=1.58
cc_2980 ( N_noxref_10_c_3470_n N_noxref_38_c_8844_n ) capacitor c=6.71402e-19 \
 //x=37.175 //y=1.915 //x2=37.925 //y2=1.495
cc_2981 ( N_noxref_10_c_3466_n N_noxref_38_M22_noxref_s ) capacitor \
 c=0.0326577f //x=37.175 //y=0.865 //x2=36.82 //y2=0.365
cc_2982 ( N_noxref_10_c_3469_n N_noxref_38_M22_noxref_s ) capacitor \
 c=3.48408e-19 //x=37.175 //y=1.52 //x2=36.82 //y2=0.365
cc_2983 ( N_noxref_10_c_3473_n N_noxref_38_M22_noxref_s ) capacitor \
 c=0.0120759f //x=37.705 //y=0.865 //x2=36.82 //y2=0.365
cc_2984 ( N_noxref_11_c_3765_p N_noxref_12_c_3886_n ) capacitor c=0.176046f \
 //x=40.585 //y=3.7 //x2=41.325 //y2=4.07
cc_2985 ( N_noxref_11_c_3758_n N_noxref_12_c_3886_n ) capacitor c=0.0293656f \
 //x=38.965 //y=3.7 //x2=41.325 //y2=4.07
cc_2986 ( N_noxref_11_c_3712_n N_noxref_12_c_3886_n ) capacitor c=0.0200089f \
 //x=38.85 //y=3.7 //x2=41.325 //y2=4.07
cc_2987 ( N_noxref_11_c_3713_n N_noxref_12_c_3886_n ) capacitor c=0.0216244f \
 //x=40.7 //y=2.08 //x2=41.325 //y2=4.07
cc_2988 ( N_noxref_11_c_3712_n N_noxref_12_c_3866_n ) capacitor c=3.49822e-19 \
 //x=38.85 //y=3.7 //x2=35.52 //y2=4.07
cc_2989 ( N_noxref_11_c_3713_n N_noxref_12_c_4030_n ) capacitor c=0.00400249f \
 //x=40.7 //y=2.08 //x2=41.44 //y2=4.535
cc_2990 ( N_noxref_11_c_3746_n N_noxref_12_c_4030_n ) capacitor c=0.00417994f \
 //x=40.7 //y=4.7 //x2=41.44 //y2=4.535
cc_2991 ( N_noxref_11_c_3765_p N_noxref_12_c_3867_n ) capacitor c=0.00720056f \
 //x=40.585 //y=3.7 //x2=41.44 //y2=2.08
cc_2992 ( N_noxref_11_c_3712_n N_noxref_12_c_3867_n ) capacitor c=9.69022e-19 \
 //x=38.85 //y=3.7 //x2=41.44 //y2=2.08
cc_2993 ( N_noxref_11_c_3713_n N_noxref_12_c_3867_n ) capacitor c=0.0739033f \
 //x=40.7 //y=2.08 //x2=41.44 //y2=2.08
cc_2994 ( N_noxref_11_c_3718_n N_noxref_12_c_3867_n ) capacitor c=0.00284029f \
 //x=40.505 //y=1.915 //x2=41.44 //y2=2.08
cc_2995 ( N_noxref_11_M93_noxref_g N_noxref_12_M95_noxref_g ) capacitor \
 c=0.0104611f //x=40.6 //y=6.02 //x2=41.48 //y2=6.02
cc_2996 ( N_noxref_11_M94_noxref_g N_noxref_12_M95_noxref_g ) capacitor \
 c=0.106811f //x=41.04 //y=6.02 //x2=41.48 //y2=6.02
cc_2997 ( N_noxref_11_M94_noxref_g N_noxref_12_M96_noxref_g ) capacitor \
 c=0.0100341f //x=41.04 //y=6.02 //x2=41.92 //y2=6.02
cc_2998 ( N_noxref_11_c_3714_n N_noxref_12_c_4039_n ) capacitor c=4.86506e-19 \
 //x=40.505 //y=0.865 //x2=41.475 //y2=0.905
cc_2999 ( N_noxref_11_c_3716_n N_noxref_12_c_4039_n ) capacitor c=0.00152104f \
 //x=40.505 //y=1.21 //x2=41.475 //y2=0.905
cc_3000 ( N_noxref_11_c_3721_n N_noxref_12_c_4039_n ) capacitor c=0.0151475f \
 //x=41.035 //y=0.865 //x2=41.475 //y2=0.905
cc_3001 ( N_noxref_11_c_3717_n N_noxref_12_c_4042_n ) capacitor c=0.00109982f \
 //x=40.505 //y=1.52 //x2=41.475 //y2=1.25
cc_3002 ( N_noxref_11_c_3723_n N_noxref_12_c_4042_n ) capacitor c=0.0111064f \
 //x=41.035 //y=1.21 //x2=41.475 //y2=1.25
cc_3003 ( N_noxref_11_c_3717_n N_noxref_12_c_4044_n ) capacitor c=9.57794e-19 \
 //x=40.505 //y=1.52 //x2=41.475 //y2=1.56
cc_3004 ( N_noxref_11_c_3718_n N_noxref_12_c_4044_n ) capacitor c=0.00662747f \
 //x=40.505 //y=1.915 //x2=41.475 //y2=1.56
cc_3005 ( N_noxref_11_c_3723_n N_noxref_12_c_4044_n ) capacitor c=0.00862358f \
 //x=41.035 //y=1.21 //x2=41.475 //y2=1.56
cc_3006 ( N_noxref_11_c_3721_n N_noxref_12_c_4047_n ) capacitor c=0.00124821f \
 //x=41.035 //y=0.865 //x2=42.005 //y2=0.905
cc_3007 ( N_noxref_11_c_3723_n N_noxref_12_c_4048_n ) capacitor c=0.00200715f \
 //x=41.035 //y=1.21 //x2=42.005 //y2=1.25
cc_3008 ( N_noxref_11_c_3713_n N_noxref_12_c_4049_n ) capacitor c=0.00282278f \
 //x=40.7 //y=2.08 //x2=41.44 //y2=2.08
cc_3009 ( N_noxref_11_c_3718_n N_noxref_12_c_4049_n ) capacitor c=0.0172771f \
 //x=40.505 //y=1.915 //x2=41.44 //y2=2.08
cc_3010 ( N_noxref_11_c_3713_n N_noxref_12_c_4051_n ) capacitor c=0.00344981f \
 //x=40.7 //y=2.08 //x2=41.47 //y2=4.7
cc_3011 ( N_noxref_11_c_3746_n N_noxref_12_c_4051_n ) capacitor c=0.0293367f \
 //x=40.7 //y=4.7 //x2=41.47 //y2=4.7
cc_3012 ( N_noxref_11_c_3765_p N_D_c_4238_n ) capacitor c=0.00669561f \
 //x=40.585 //y=3.7 //x2=49.465 //y2=2.59
cc_3013 ( N_noxref_11_c_3758_n N_D_c_4238_n ) capacitor c=6.305e-19 //x=38.965 \
 //y=3.7 //x2=49.465 //y2=2.59
cc_3014 ( N_noxref_11_c_3712_n N_D_c_4238_n ) capacitor c=0.0165961f //x=38.85 \
 //y=3.7 //x2=49.465 //y2=2.59
cc_3015 ( N_noxref_11_c_3713_n N_D_c_4238_n ) capacitor c=0.0177872f //x=40.7 \
 //y=2.08 //x2=49.465 //y2=2.59
cc_3016 ( N_noxref_11_c_3765_p N_CLK_c_5092_n ) capacitor c=0.0104236f \
 //x=40.585 //y=3.7 //x2=45.025 //y2=4.44
cc_3017 ( N_noxref_11_c_3758_n N_CLK_c_5092_n ) capacitor c=8.86008e-19 \
 //x=38.965 //y=3.7 //x2=45.025 //y2=4.44
cc_3018 ( N_noxref_11_c_3727_n N_CLK_c_5092_n ) capacitor c=0.0185297f \
 //x=38.285 //y=5.2 //x2=45.025 //y2=4.44
cc_3019 ( N_noxref_11_c_3731_n N_CLK_c_5092_n ) capacitor c=0.018142f \
 //x=37.575 //y=5.2 //x2=45.025 //y2=4.44
cc_3020 ( N_noxref_11_c_3712_n N_CLK_c_5092_n ) capacitor c=0.0208321f \
 //x=38.85 //y=3.7 //x2=45.025 //y2=4.44
cc_3021 ( N_noxref_11_c_3713_n N_CLK_c_5092_n ) capacitor c=0.0198304f \
 //x=40.7 //y=2.08 //x2=45.025 //y2=4.44
cc_3022 ( N_noxref_11_c_3746_n N_CLK_c_5092_n ) capacitor c=0.0107057f \
 //x=40.7 //y=4.7 //x2=45.025 //y2=4.44
cc_3023 ( N_noxref_11_c_3804_p N_noxref_21_c_6904_n ) capacitor c=0.0146822f \
 //x=38.495 //y=1.655 //x2=42.065 //y2=2.22
cc_3024 ( N_noxref_11_c_3712_n N_noxref_21_c_6904_n ) capacitor c=0.0199049f \
 //x=38.85 //y=3.7 //x2=42.065 //y2=2.22
cc_3025 ( N_noxref_11_c_3713_n N_noxref_21_c_6904_n ) capacitor c=0.0185012f \
 //x=40.7 //y=2.08 //x2=42.065 //y2=2.22
cc_3026 ( N_noxref_11_c_3718_n N_noxref_21_c_6904_n ) capacitor c=0.00894156f \
 //x=40.505 //y=1.915 //x2=42.065 //y2=2.22
cc_3027 ( N_noxref_11_c_3712_n N_noxref_21_c_6909_n ) capacitor c=0.00122089f \
 //x=38.85 //y=3.7 //x2=38.225 //y2=2.22
cc_3028 ( N_noxref_11_c_3727_n N_noxref_21_c_7001_n ) capacitor c=0.0127164f \
 //x=38.285 //y=5.2 //x2=38.11 //y2=4.535
cc_3029 ( N_noxref_11_c_3712_n N_noxref_21_c_7001_n ) capacitor c=0.0101284f \
 //x=38.85 //y=3.7 //x2=38.11 //y2=4.535
cc_3030 ( N_noxref_11_c_3758_n N_noxref_21_c_6939_n ) capacitor c=0.00329059f \
 //x=38.965 //y=3.7 //x2=38.11 //y2=2.08
cc_3031 ( N_noxref_11_c_3712_n N_noxref_21_c_6939_n ) capacitor c=0.0696008f \
 //x=38.85 //y=3.7 //x2=38.11 //y2=2.08
cc_3032 ( N_noxref_11_c_3713_n N_noxref_21_c_6939_n ) capacitor c=0.00100713f \
 //x=40.7 //y=2.08 //x2=38.11 //y2=2.08
cc_3033 ( N_noxref_11_M94_noxref_g N_noxref_21_c_6959_n ) capacitor \
 c=0.0169521f //x=41.04 //y=6.02 //x2=41.615 //y2=5.2
cc_3034 ( N_noxref_11_c_3713_n N_noxref_21_c_6963_n ) capacitor c=0.00521572f \
 //x=40.7 //y=2.08 //x2=40.905 //y2=5.2
cc_3035 ( N_noxref_11_M93_noxref_g N_noxref_21_c_6963_n ) capacitor \
 c=0.0177326f //x=40.6 //y=6.02 //x2=40.905 //y2=5.2
cc_3036 ( N_noxref_11_c_3746_n N_noxref_21_c_6963_n ) capacitor c=0.00581252f \
 //x=40.7 //y=4.7 //x2=40.905 //y2=5.2
cc_3037 ( N_noxref_11_c_3712_n N_noxref_21_c_6942_n ) capacitor c=3.49822e-19 \
 //x=38.85 //y=3.7 //x2=42.18 //y2=2.22
cc_3038 ( N_noxref_11_c_3713_n N_noxref_21_c_6942_n ) capacitor c=0.00332679f \
 //x=40.7 //y=2.08 //x2=42.18 //y2=2.22
cc_3039 ( N_noxref_11_c_3727_n N_noxref_21_M91_noxref_g ) capacitor \
 c=0.0166421f //x=38.285 //y=5.2 //x2=38.15 //y2=6.02
cc_3040 ( N_noxref_11_M91_noxref_d N_noxref_21_M91_noxref_g ) capacitor \
 c=0.0173476f //x=38.225 //y=5.02 //x2=38.15 //y2=6.02
cc_3041 ( N_noxref_11_c_3733_n N_noxref_21_M92_noxref_g ) capacitor \
 c=0.018922f //x=38.765 //y=5.2 //x2=38.59 //y2=6.02
cc_3042 ( N_noxref_11_M91_noxref_d N_noxref_21_M92_noxref_g ) capacitor \
 c=0.0179769f //x=38.225 //y=5.02 //x2=38.59 //y2=6.02
cc_3043 ( N_noxref_11_M23_noxref_d N_noxref_21_c_7009_n ) capacitor \
 c=0.00217566f //x=38.22 //y=0.905 //x2=38.145 //y2=0.905
cc_3044 ( N_noxref_11_M23_noxref_d N_noxref_21_c_7012_n ) capacitor \
 c=0.0034598f //x=38.22 //y=0.905 //x2=38.145 //y2=1.25
cc_3045 ( N_noxref_11_M23_noxref_d N_noxref_21_c_7014_n ) capacitor \
 c=0.0066953f //x=38.22 //y=0.905 //x2=38.145 //y2=1.56
cc_3046 ( N_noxref_11_c_3712_n N_noxref_21_c_7046_n ) capacitor c=0.0142673f \
 //x=38.85 //y=3.7 //x2=38.515 //y2=4.79
cc_3047 ( N_noxref_11_c_3828_p N_noxref_21_c_7046_n ) capacitor c=0.00407665f \
 //x=38.37 //y=5.2 //x2=38.515 //y2=4.79
cc_3048 ( N_noxref_11_M23_noxref_d N_noxref_21_c_7048_n ) capacitor \
 c=0.00241102f //x=38.22 //y=0.905 //x2=38.52 //y2=0.75
cc_3049 ( N_noxref_11_c_3711_n N_noxref_21_c_7049_n ) capacitor c=0.00371277f \
 //x=38.765 //y=1.655 //x2=38.52 //y2=1.405
cc_3050 ( N_noxref_11_M23_noxref_d N_noxref_21_c_7049_n ) capacitor \
 c=0.0137169f //x=38.22 //y=0.905 //x2=38.52 //y2=1.405
cc_3051 ( N_noxref_11_M23_noxref_d N_noxref_21_c_7017_n ) capacitor \
 c=0.00132245f //x=38.22 //y=0.905 //x2=38.675 //y2=0.905
cc_3052 ( N_noxref_11_c_3711_n N_noxref_21_c_7018_n ) capacitor c=0.00457401f \
 //x=38.765 //y=1.655 //x2=38.675 //y2=1.25
cc_3053 ( N_noxref_11_M23_noxref_d N_noxref_21_c_7018_n ) capacitor \
 c=0.00566463f //x=38.22 //y=0.905 //x2=38.675 //y2=1.25
cc_3054 ( N_noxref_11_c_3712_n N_noxref_21_c_7019_n ) capacitor c=0.00709342f \
 //x=38.85 //y=3.7 //x2=38.11 //y2=2.08
cc_3055 ( N_noxref_11_c_3712_n N_noxref_21_c_7055_n ) capacitor c=0.00306024f \
 //x=38.85 //y=3.7 //x2=38.11 //y2=1.915
cc_3056 ( N_noxref_11_M23_noxref_d N_noxref_21_c_7055_n ) capacitor \
 c=0.00660593f //x=38.22 //y=0.905 //x2=38.11 //y2=1.915
cc_3057 ( N_noxref_11_c_3727_n N_noxref_21_c_7021_n ) capacitor c=0.00346527f \
 //x=38.285 //y=5.2 //x2=38.14 //y2=4.7
cc_3058 ( N_noxref_11_c_3712_n N_noxref_21_c_7021_n ) capacitor c=0.00533692f \
 //x=38.85 //y=3.7 //x2=38.14 //y2=4.7
cc_3059 ( N_noxref_11_M94_noxref_g N_noxref_21_M93_noxref_d ) capacitor \
 c=0.0173476f //x=41.04 //y=6.02 //x2=40.675 //y2=5.02
cc_3060 ( N_noxref_11_c_3765_p N_noxref_23_c_7498_n ) capacitor c=0.0868505f \
 //x=40.585 //y=3.7 //x2=70.185 //y2=2.96
cc_3061 ( N_noxref_11_c_3758_n N_noxref_23_c_7498_n ) capacitor c=0.0133597f \
 //x=38.965 //y=3.7 //x2=70.185 //y2=2.96
cc_3062 ( N_noxref_11_c_3712_n N_noxref_23_c_7498_n ) capacitor c=0.0214247f \
 //x=38.85 //y=3.7 //x2=70.185 //y2=2.96
cc_3063 ( N_noxref_11_c_3713_n N_noxref_23_c_7498_n ) capacitor c=0.021399f \
 //x=40.7 //y=2.08 //x2=70.185 //y2=2.96
cc_3064 ( N_noxref_11_c_3804_p N_noxref_38_c_8856_n ) capacitor c=3.15806e-19 \
 //x=38.495 //y=1.655 //x2=36.955 //y2=1.495
cc_3065 ( N_noxref_11_c_3804_p N_noxref_38_c_8844_n ) capacitor c=0.0203424f \
 //x=38.495 //y=1.655 //x2=37.925 //y2=1.495
cc_3066 ( N_noxref_11_c_3711_n N_noxref_38_c_8845_n ) capacitor c=0.00457164f \
 //x=38.765 //y=1.655 //x2=38.81 //y2=0.53
cc_3067 ( N_noxref_11_M23_noxref_d N_noxref_38_c_8845_n ) capacitor \
 c=0.0115831f //x=38.22 //y=0.905 //x2=38.81 //y2=0.53
cc_3068 ( N_noxref_11_c_3711_n N_noxref_38_M22_noxref_s ) capacitor \
 c=0.013435f //x=38.765 //y=1.655 //x2=36.82 //y2=0.365
cc_3069 ( N_noxref_11_M23_noxref_d N_noxref_38_M22_noxref_s ) capacitor \
 c=0.043966f //x=38.22 //y=0.905 //x2=36.82 //y2=0.365
cc_3070 ( N_noxref_11_c_3711_n N_noxref_39_c_8910_n ) capacitor c=3.22188e-19 \
 //x=38.765 //y=1.655 //x2=40.285 //y2=1.495
cc_3071 ( N_noxref_11_c_3718_n N_noxref_39_c_8910_n ) capacitor c=0.0034165f \
 //x=40.505 //y=1.915 //x2=40.285 //y2=1.495
cc_3072 ( N_noxref_11_c_3713_n N_noxref_39_c_8891_n ) capacitor c=0.011618f \
 //x=40.7 //y=2.08 //x2=41.17 //y2=1.58
cc_3073 ( N_noxref_11_c_3717_n N_noxref_39_c_8891_n ) capacitor c=0.00696403f \
 //x=40.505 //y=1.52 //x2=41.17 //y2=1.58
cc_3074 ( N_noxref_11_c_3718_n N_noxref_39_c_8891_n ) capacitor c=0.0174694f \
 //x=40.505 //y=1.915 //x2=41.17 //y2=1.58
cc_3075 ( N_noxref_11_c_3720_n N_noxref_39_c_8891_n ) capacitor c=0.00776811f \
 //x=40.88 //y=1.365 //x2=41.17 //y2=1.58
cc_3076 ( N_noxref_11_c_3723_n N_noxref_39_c_8891_n ) capacitor c=0.00339872f \
 //x=41.035 //y=1.21 //x2=41.17 //y2=1.58
cc_3077 ( N_noxref_11_c_3718_n N_noxref_39_c_8898_n ) capacitor c=6.71402e-19 \
 //x=40.505 //y=1.915 //x2=41.255 //y2=1.495
cc_3078 ( N_noxref_11_c_3714_n N_noxref_39_M24_noxref_s ) capacitor \
 c=0.0326577f //x=40.505 //y=0.865 //x2=40.15 //y2=0.365
cc_3079 ( N_noxref_11_c_3717_n N_noxref_39_M24_noxref_s ) capacitor \
 c=3.48408e-19 //x=40.505 //y=1.52 //x2=40.15 //y2=0.365
cc_3080 ( N_noxref_11_c_3721_n N_noxref_39_M24_noxref_s ) capacitor \
 c=0.0120759f //x=41.035 //y=0.865 //x2=40.15 //y2=0.365
cc_3081 ( N_noxref_12_c_3882_n N_D_c_4217_n ) capacitor c=0.011848f //x=31.335 \
 //y=4.07 //x2=28.005 //y2=2.59
cc_3082 ( N_noxref_12_c_3884_n N_D_c_4217_n ) capacitor c=4.25679e-19 \
 //x=22.685 //y=4.07 //x2=28.005 //y2=2.59
cc_3083 ( N_noxref_12_c_3862_n N_D_c_4217_n ) capacitor c=0.0223514f //x=22.57 \
 //y=2.08 //x2=28.005 //y2=2.59
cc_3084 ( N_noxref_12_c_3873_n N_D_c_4217_n ) capacitor c=0.00712164f \
 //x=22.27 //y=1.915 //x2=28.005 //y2=2.59
cc_3085 ( N_noxref_12_c_3886_n N_D_c_4238_n ) capacitor c=0.0108438f \
 //x=41.325 //y=4.07 //x2=49.465 //y2=2.59
cc_3086 ( N_noxref_12_c_3863_n N_D_c_4238_n ) capacitor c=0.0204615f //x=31.45 \
 //y=2.08 //x2=49.465 //y2=2.59
cc_3087 ( N_noxref_12_c_4059_p N_D_c_4238_n ) capacitor c=0.0102711f \
 //x=35.165 //y=1.655 //x2=49.465 //y2=2.59
cc_3088 ( N_noxref_12_c_3866_n N_D_c_4238_n ) capacitor c=0.0210598f //x=35.52 \
 //y=4.07 //x2=49.465 //y2=2.59
cc_3089 ( N_noxref_12_c_3867_n N_D_c_4238_n ) capacitor c=0.0169223f //x=41.44 \
 //y=2.08 //x2=49.465 //y2=2.59
cc_3090 ( N_noxref_12_c_3965_n N_D_c_4238_n ) capacitor c=0.00219932f \
 //x=31.45 //y=2.08 //x2=49.465 //y2=2.59
cc_3091 ( N_noxref_12_c_3882_n N_D_c_4255_n ) capacitor c=0.0169317f \
 //x=31.335 //y=4.07 //x2=28.12 //y2=2.08
cc_3092 ( N_noxref_12_c_3882_n N_CLK_c_5061_n ) capacitor c=0.656956f \
 //x=31.335 //y=4.07 //x2=34.665 //y2=4.44
cc_3093 ( N_noxref_12_c_3885_n N_CLK_c_5061_n ) capacitor c=0.270915f \
 //x=35.405 //y=4.07 //x2=34.665 //y2=4.44
cc_3094 ( N_noxref_12_c_3944_n N_CLK_c_5061_n ) capacitor c=0.0263375f \
 //x=31.565 //y=4.07 //x2=34.665 //y2=4.44
cc_3095 ( N_noxref_12_c_3946_n N_CLK_c_5061_n ) capacitor c=0.0016972f \
 //x=31.45 //y=4.535 //x2=34.665 //y2=4.44
cc_3096 ( N_noxref_12_c_3863_n N_CLK_c_5061_n ) capacitor c=0.0207534f \
 //x=31.45 //y=2.08 //x2=34.665 //y2=4.44
cc_3097 ( N_noxref_12_c_3898_n N_CLK_c_5061_n ) capacitor c=0.0172877f \
 //x=34.245 //y=5.2 //x2=34.665 //y2=4.44
cc_3098 ( N_noxref_12_c_3992_n N_CLK_c_5061_n ) capacitor c=0.00960248f \
 //x=31.855 //y=4.79 //x2=34.665 //y2=4.44
cc_3099 ( N_noxref_12_c_3967_n N_CLK_c_5061_n ) capacitor c=0.00203982f \
 //x=31.48 //y=4.7 //x2=34.665 //y2=4.44
cc_3100 ( N_noxref_12_c_3882_n N_CLK_c_5079_n ) capacitor c=0.102795f \
 //x=31.335 //y=4.07 //x2=23.795 //y2=4.44
cc_3101 ( N_noxref_12_c_3884_n N_CLK_c_5079_n ) capacitor c=0.0290178f \
 //x=22.685 //y=4.07 //x2=23.795 //y2=4.44
cc_3102 ( N_noxref_12_c_3862_n N_CLK_c_5079_n ) capacitor c=0.0242383f \
 //x=22.57 //y=2.08 //x2=23.795 //y2=4.44
cc_3103 ( N_noxref_12_c_3922_n N_CLK_c_5079_n ) capacitor c=0.0168514f \
 //x=22.845 //y=4.79 //x2=23.795 //y2=4.44
cc_3104 ( N_noxref_12_c_3885_n N_CLK_c_5092_n ) capacitor c=0.0444029f \
 //x=35.405 //y=4.07 //x2=45.025 //y2=4.44
cc_3105 ( N_noxref_12_c_3886_n N_CLK_c_5092_n ) capacitor c=0.526398f \
 //x=41.325 //y=4.07 //x2=45.025 //y2=4.44
cc_3106 ( N_noxref_12_c_3888_n N_CLK_c_5092_n ) capacitor c=0.0265844f \
 //x=35.635 //y=4.07 //x2=45.025 //y2=4.44
cc_3107 ( N_noxref_12_c_3894_n N_CLK_c_5092_n ) capacitor c=0.0173598f \
 //x=34.955 //y=5.2 //x2=45.025 //y2=4.44
cc_3108 ( N_noxref_12_c_3866_n N_CLK_c_5092_n ) capacitor c=0.0226667f \
 //x=35.52 //y=4.07 //x2=45.025 //y2=4.44
cc_3109 ( N_noxref_12_c_4030_n N_CLK_c_5092_n ) capacitor c=0.0016972f \
 //x=41.44 //y=4.535 //x2=45.025 //y2=4.44
cc_3110 ( N_noxref_12_c_3867_n N_CLK_c_5092_n ) capacitor c=0.0207534f \
 //x=41.44 //y=2.08 //x2=45.025 //y2=4.44
cc_3111 ( N_noxref_12_c_4083_p N_CLK_c_5092_n ) capacitor c=0.00720343f \
 //x=41.845 //y=4.79 //x2=45.025 //y2=4.44
cc_3112 ( N_noxref_12_c_4051_n N_CLK_c_5092_n ) capacitor c=0.0019199f \
 //x=41.47 //y=4.7 //x2=45.025 //y2=4.44
cc_3113 ( N_noxref_12_c_3885_n N_CLK_c_5111_n ) capacitor c=0.0267161f \
 //x=35.405 //y=4.07 //x2=34.895 //y2=4.44
cc_3114 ( N_noxref_12_c_3894_n N_CLK_c_5111_n ) capacitor c=0.0023575f \
 //x=34.955 //y=5.2 //x2=34.895 //y2=4.44
cc_3115 ( N_noxref_12_c_3866_n N_CLK_c_5111_n ) capacitor c=0.00151334f \
 //x=35.52 //y=4.07 //x2=34.895 //y2=4.44
cc_3116 ( N_noxref_12_c_3882_n N_CLK_c_5028_n ) capacitor c=0.0247116f \
 //x=31.335 //y=4.07 //x2=23.68 //y2=2.08
cc_3117 ( N_noxref_12_c_3884_n N_CLK_c_5028_n ) capacitor c=0.00128547f \
 //x=22.685 //y=4.07 //x2=23.68 //y2=2.08
cc_3118 ( N_noxref_12_c_3862_n N_CLK_c_5028_n ) capacitor c=0.0476719f \
 //x=22.57 //y=2.08 //x2=23.68 //y2=2.08
cc_3119 ( N_noxref_12_c_3873_n N_CLK_c_5028_n ) capacitor c=0.00238338f \
 //x=22.27 //y=1.915 //x2=23.68 //y2=2.08
cc_3120 ( N_noxref_12_c_4024_n N_CLK_c_5028_n ) capacitor c=0.00147352f \
 //x=23.135 //y=4.79 //x2=23.68 //y2=2.08
cc_3121 ( N_noxref_12_c_3922_n N_CLK_c_5028_n ) capacitor c=0.00141297f \
 //x=22.845 //y=4.79 //x2=23.68 //y2=2.08
cc_3122 ( N_noxref_12_c_3894_n N_CLK_c_5363_n ) capacitor c=0.0126416f \
 //x=34.955 //y=5.2 //x2=34.78 //y2=4.535
cc_3123 ( N_noxref_12_c_3866_n N_CLK_c_5363_n ) capacitor c=0.00923416f \
 //x=35.52 //y=4.07 //x2=34.78 //y2=4.535
cc_3124 ( N_noxref_12_c_3885_n N_CLK_c_5029_n ) capacitor c=0.0187718f \
 //x=35.405 //y=4.07 //x2=34.78 //y2=2.08
cc_3125 ( N_noxref_12_c_3888_n N_CLK_c_5029_n ) capacitor c=0.00117715f \
 //x=35.635 //y=4.07 //x2=34.78 //y2=2.08
cc_3126 ( N_noxref_12_c_3894_n N_CLK_c_5029_n ) capacitor c=3.74769e-19 \
 //x=34.955 //y=5.2 //x2=34.78 //y2=2.08
cc_3127 ( N_noxref_12_c_3866_n N_CLK_c_5029_n ) capacitor c=0.0700213f \
 //x=35.52 //y=4.07 //x2=34.78 //y2=2.08
cc_3128 ( N_noxref_12_M71_noxref_g N_CLK_M73_noxref_g ) capacitor c=0.0105869f \
 //x=22.77 //y=6.02 //x2=23.65 //y2=6.02
cc_3129 ( N_noxref_12_M72_noxref_g N_CLK_M73_noxref_g ) capacitor c=0.10632f \
 //x=23.21 //y=6.02 //x2=23.65 //y2=6.02
cc_3130 ( N_noxref_12_M72_noxref_g N_CLK_M74_noxref_g ) capacitor c=0.0101598f \
 //x=23.21 //y=6.02 //x2=24.09 //y2=6.02
cc_3131 ( N_noxref_12_c_3894_n N_CLK_M87_noxref_g ) capacitor c=0.0166421f \
 //x=34.955 //y=5.2 //x2=34.82 //y2=6.02
cc_3132 ( N_noxref_12_M87_noxref_d N_CLK_M87_noxref_g ) capacitor c=0.0173476f \
 //x=34.895 //y=5.02 //x2=34.82 //y2=6.02
cc_3133 ( N_noxref_12_c_3900_n N_CLK_M88_noxref_g ) capacitor c=0.018922f \
 //x=35.435 //y=5.2 //x2=35.26 //y2=6.02
cc_3134 ( N_noxref_12_M87_noxref_d N_CLK_M88_noxref_g ) capacitor c=0.0179769f \
 //x=34.895 //y=5.02 //x2=35.26 //y2=6.02
cc_3135 ( N_noxref_12_c_3869_n N_CLK_c_5461_n ) capacitor c=5.72482e-19 \
 //x=22.27 //y=0.875 //x2=23.245 //y2=0.91
cc_3136 ( N_noxref_12_c_3871_n N_CLK_c_5461_n ) capacitor c=0.00149976f \
 //x=22.27 //y=1.22 //x2=23.245 //y2=0.91
cc_3137 ( N_noxref_12_c_3876_n N_CLK_c_5461_n ) capacitor c=0.0160123f \
 //x=22.8 //y=0.875 //x2=23.245 //y2=0.91
cc_3138 ( N_noxref_12_c_3872_n N_CLK_c_5464_n ) capacitor c=0.00111227f \
 //x=22.27 //y=1.53 //x2=23.245 //y2=1.22
cc_3139 ( N_noxref_12_c_3878_n N_CLK_c_5464_n ) capacitor c=0.0124075f \
 //x=22.8 //y=1.22 //x2=23.245 //y2=1.22
cc_3140 ( N_noxref_12_c_3876_n N_CLK_c_5347_n ) capacitor c=0.00103227f \
 //x=22.8 //y=0.875 //x2=23.77 //y2=0.91
cc_3141 ( N_noxref_12_c_3878_n N_CLK_c_5348_n ) capacitor c=0.0010154f \
 //x=22.8 //y=1.22 //x2=23.77 //y2=1.22
cc_3142 ( N_noxref_12_c_3878_n N_CLK_c_5349_n ) capacitor c=9.23422e-19 \
 //x=22.8 //y=1.22 //x2=23.77 //y2=1.45
cc_3143 ( N_noxref_12_c_3862_n N_CLK_c_5350_n ) capacitor c=0.00231304f \
 //x=22.57 //y=2.08 //x2=23.77 //y2=1.915
cc_3144 ( N_noxref_12_c_3873_n N_CLK_c_5350_n ) capacitor c=0.00964411f \
 //x=22.27 //y=1.915 //x2=23.77 //y2=1.915
cc_3145 ( N_noxref_12_M21_noxref_d N_CLK_c_5372_n ) capacitor c=0.00217566f \
 //x=34.89 //y=0.905 //x2=34.815 //y2=0.905
cc_3146 ( N_noxref_12_M21_noxref_d N_CLK_c_5375_n ) capacitor c=0.0034598f \
 //x=34.89 //y=0.905 //x2=34.815 //y2=1.25
cc_3147 ( N_noxref_12_M21_noxref_d N_CLK_c_5377_n ) capacitor c=0.00656319f \
 //x=34.89 //y=0.905 //x2=34.815 //y2=1.56
cc_3148 ( N_noxref_12_c_3866_n N_CLK_c_5474_n ) capacitor c=0.0142673f \
 //x=35.52 //y=4.07 //x2=35.185 //y2=4.79
cc_3149 ( N_noxref_12_c_4121_p N_CLK_c_5474_n ) capacitor c=0.00407665f \
 //x=35.04 //y=5.2 //x2=35.185 //y2=4.79
cc_3150 ( N_noxref_12_M21_noxref_d N_CLK_c_5476_n ) capacitor c=0.00241102f \
 //x=34.89 //y=0.905 //x2=35.19 //y2=0.75
cc_3151 ( N_noxref_12_c_3865_n N_CLK_c_5477_n ) capacitor c=0.00359704f \
 //x=35.435 //y=1.655 //x2=35.19 //y2=1.405
cc_3152 ( N_noxref_12_M21_noxref_d N_CLK_c_5477_n ) capacitor c=0.0138845f \
 //x=34.89 //y=0.905 //x2=35.19 //y2=1.405
cc_3153 ( N_noxref_12_M21_noxref_d N_CLK_c_5380_n ) capacitor c=0.00132245f \
 //x=34.89 //y=0.905 //x2=35.345 //y2=0.905
cc_3154 ( N_noxref_12_c_3865_n N_CLK_c_5381_n ) capacitor c=0.00457401f \
 //x=35.435 //y=1.655 //x2=35.345 //y2=1.25
cc_3155 ( N_noxref_12_M21_noxref_d N_CLK_c_5381_n ) capacitor c=0.00566463f \
 //x=34.89 //y=0.905 //x2=35.345 //y2=1.25
cc_3156 ( N_noxref_12_c_3862_n N_CLK_c_5354_n ) capacitor c=0.00183762f \
 //x=22.57 //y=2.08 //x2=23.68 //y2=4.7
cc_3157 ( N_noxref_12_c_4024_n N_CLK_c_5354_n ) capacitor c=0.0168581f \
 //x=23.135 //y=4.79 //x2=23.68 //y2=4.7
cc_3158 ( N_noxref_12_c_3922_n N_CLK_c_5354_n ) capacitor c=0.00484466f \
 //x=22.845 //y=4.79 //x2=23.68 //y2=4.7
cc_3159 ( N_noxref_12_c_3866_n N_CLK_c_5382_n ) capacitor c=0.00772308f \
 //x=35.52 //y=4.07 //x2=34.78 //y2=2.08
cc_3160 ( N_noxref_12_c_3866_n N_CLK_c_5486_n ) capacitor c=0.00306024f \
 //x=35.52 //y=4.07 //x2=34.78 //y2=1.915
cc_3161 ( N_noxref_12_M21_noxref_d N_CLK_c_5486_n ) capacitor c=0.00660593f \
 //x=34.89 //y=0.905 //x2=34.78 //y2=1.915
cc_3162 ( N_noxref_12_c_3894_n N_CLK_c_5384_n ) capacitor c=0.00346519f \
 //x=34.955 //y=5.2 //x2=34.81 //y2=4.7
cc_3163 ( N_noxref_12_c_3866_n N_CLK_c_5384_n ) capacitor c=0.00518077f \
 //x=35.52 //y=4.07 //x2=34.81 //y2=4.7
cc_3164 ( N_noxref_12_c_3886_n N_noxref_19_c_6212_n ) capacitor c=0.00649178f \
 //x=41.325 //y=4.07 //x2=44.145 //y2=4.07
cc_3165 ( N_noxref_12_c_3867_n N_noxref_19_c_6190_n ) capacitor c=8.8171e-19 \
 //x=41.44 //y=2.08 //x2=44.03 //y2=2.08
cc_3166 ( N_noxref_12_c_3867_n N_noxref_21_c_6904_n ) capacitor c=0.0178519f \
 //x=41.44 //y=2.08 //x2=42.065 //y2=2.22
cc_3167 ( N_noxref_12_c_4139_p N_noxref_21_c_6904_n ) capacitor c=3.11115e-19 \
 //x=41.85 //y=1.405 //x2=42.065 //y2=2.22
cc_3168 ( N_noxref_12_c_4049_n N_noxref_21_c_6904_n ) capacitor c=0.00570799f \
 //x=41.44 //y=2.08 //x2=42.065 //y2=2.22
cc_3169 ( N_noxref_12_c_3867_n N_noxref_21_c_6935_n ) capacitor c=0.00125295f \
 //x=41.44 //y=2.08 //x2=42.295 //y2=2.22
cc_3170 ( N_noxref_12_c_4049_n N_noxref_21_c_6935_n ) capacitor c=6.64454e-19 \
 //x=41.44 //y=2.08 //x2=42.295 //y2=2.22
cc_3171 ( N_noxref_12_c_3886_n N_noxref_21_c_6939_n ) capacitor c=0.0207919f \
 //x=41.325 //y=4.07 //x2=38.11 //y2=2.08
cc_3172 ( N_noxref_12_c_3866_n N_noxref_21_c_6939_n ) capacitor c=0.00104099f \
 //x=35.52 //y=4.07 //x2=38.11 //y2=2.08
cc_3173 ( N_noxref_12_c_4030_n N_noxref_21_c_6959_n ) capacitor c=0.0126603f \
 //x=41.44 //y=4.535 //x2=41.615 //y2=5.2
cc_3174 ( N_noxref_12_M95_noxref_g N_noxref_21_c_6959_n ) capacitor \
 c=0.0166421f //x=41.48 //y=6.02 //x2=41.615 //y2=5.2
cc_3175 ( N_noxref_12_c_4051_n N_noxref_21_c_6959_n ) capacitor c=0.00346527f \
 //x=41.47 //y=4.7 //x2=41.615 //y2=5.2
cc_3176 ( N_noxref_12_M96_noxref_g N_noxref_21_c_6965_n ) capacitor \
 c=0.018922f //x=41.92 //y=6.02 //x2=42.095 //y2=5.2
cc_3177 ( N_noxref_12_c_4139_p N_noxref_21_c_6941_n ) capacitor c=0.00371277f \
 //x=41.85 //y=1.405 //x2=42.095 //y2=1.655
cc_3178 ( N_noxref_12_c_4048_n N_noxref_21_c_6941_n ) capacitor c=0.00457401f \
 //x=42.005 //y=1.25 //x2=42.095 //y2=1.655
cc_3179 ( N_noxref_12_c_3886_n N_noxref_21_c_6942_n ) capacitor c=0.00423741f \
 //x=41.325 //y=4.07 //x2=42.18 //y2=2.22
cc_3180 ( N_noxref_12_c_4030_n N_noxref_21_c_6942_n ) capacitor c=0.0101115f \
 //x=41.44 //y=4.535 //x2=42.18 //y2=2.22
cc_3181 ( N_noxref_12_c_3867_n N_noxref_21_c_6942_n ) capacitor c=0.0718861f \
 //x=41.44 //y=2.08 //x2=42.18 //y2=2.22
cc_3182 ( N_noxref_12_c_4083_p N_noxref_21_c_6942_n ) capacitor c=0.0142673f \
 //x=41.845 //y=4.79 //x2=42.18 //y2=2.22
cc_3183 ( N_noxref_12_c_4049_n N_noxref_21_c_6942_n ) capacitor c=0.00708548f \
 //x=41.44 //y=2.08 //x2=42.18 //y2=2.22
cc_3184 ( N_noxref_12_c_4156_p N_noxref_21_c_6942_n ) capacitor c=0.00306024f \
 //x=41.44 //y=1.915 //x2=42.18 //y2=2.22
cc_3185 ( N_noxref_12_c_4051_n N_noxref_21_c_6942_n ) capacitor c=0.00517969f \
 //x=41.47 //y=4.7 //x2=42.18 //y2=2.22
cc_3186 ( N_noxref_12_c_4083_p N_noxref_21_c_7080_n ) capacitor c=0.00407665f \
 //x=41.845 //y=4.79 //x2=41.7 //y2=5.2
cc_3187 ( N_noxref_12_c_4039_n N_noxref_21_M25_noxref_d ) capacitor \
 c=0.00217566f //x=41.475 //y=0.905 //x2=41.55 //y2=0.905
cc_3188 ( N_noxref_12_c_4042_n N_noxref_21_M25_noxref_d ) capacitor \
 c=0.0034598f //x=41.475 //y=1.25 //x2=41.55 //y2=0.905
cc_3189 ( N_noxref_12_c_4044_n N_noxref_21_M25_noxref_d ) capacitor \
 c=0.0066953f //x=41.475 //y=1.56 //x2=41.55 //y2=0.905
cc_3190 ( N_noxref_12_c_4162_p N_noxref_21_M25_noxref_d ) capacitor \
 c=0.00241102f //x=41.85 //y=0.75 //x2=41.55 //y2=0.905
cc_3191 ( N_noxref_12_c_4139_p N_noxref_21_M25_noxref_d ) capacitor \
 c=0.0137169f //x=41.85 //y=1.405 //x2=41.55 //y2=0.905
cc_3192 ( N_noxref_12_c_4047_n N_noxref_21_M25_noxref_d ) capacitor \
 c=0.00132245f //x=42.005 //y=0.905 //x2=41.55 //y2=0.905
cc_3193 ( N_noxref_12_c_4048_n N_noxref_21_M25_noxref_d ) capacitor \
 c=0.00566463f //x=42.005 //y=1.25 //x2=41.55 //y2=0.905
cc_3194 ( N_noxref_12_c_4156_p N_noxref_21_M25_noxref_d ) capacitor \
 c=0.00660593f //x=41.44 //y=1.915 //x2=41.55 //y2=0.905
cc_3195 ( N_noxref_12_M95_noxref_g N_noxref_21_M95_noxref_d ) capacitor \
 c=0.0173476f //x=41.48 //y=6.02 //x2=41.555 //y2=5.02
cc_3196 ( N_noxref_12_M96_noxref_g N_noxref_21_M95_noxref_d ) capacitor \
 c=0.0179769f //x=41.92 //y=6.02 //x2=41.555 //y2=5.02
cc_3197 ( N_noxref_12_c_3882_n N_noxref_23_c_7498_n ) capacitor c=0.0615741f \
 //x=31.335 //y=4.07 //x2=70.185 //y2=2.96
cc_3198 ( N_noxref_12_c_3884_n N_noxref_23_c_7498_n ) capacitor c=0.00776275f \
 //x=22.685 //y=4.07 //x2=70.185 //y2=2.96
cc_3199 ( N_noxref_12_c_3885_n N_noxref_23_c_7498_n ) capacitor c=0.0112822f \
 //x=35.405 //y=4.07 //x2=70.185 //y2=2.96
cc_3200 ( N_noxref_12_c_3944_n N_noxref_23_c_7498_n ) capacitor c=3.56521e-19 \
 //x=31.565 //y=4.07 //x2=70.185 //y2=2.96
cc_3201 ( N_noxref_12_c_3886_n N_noxref_23_c_7498_n ) capacitor c=0.0695653f \
 //x=41.325 //y=4.07 //x2=70.185 //y2=2.96
cc_3202 ( N_noxref_12_c_3888_n N_noxref_23_c_7498_n ) capacitor c=4.50823e-19 \
 //x=35.635 //y=4.07 //x2=70.185 //y2=2.96
cc_3203 ( N_noxref_12_c_3862_n N_noxref_23_c_7498_n ) capacitor c=0.0237066f \
 //x=22.57 //y=2.08 //x2=70.185 //y2=2.96
cc_3204 ( N_noxref_12_c_3863_n N_noxref_23_c_7498_n ) capacitor c=0.019291f \
 //x=31.45 //y=2.08 //x2=70.185 //y2=2.96
cc_3205 ( N_noxref_12_c_3866_n N_noxref_23_c_7498_n ) capacitor c=0.0210811f \
 //x=35.52 //y=4.07 //x2=70.185 //y2=2.96
cc_3206 ( N_noxref_12_c_3867_n N_noxref_23_c_7498_n ) capacitor c=0.0209015f \
 //x=41.44 //y=2.08 //x2=70.185 //y2=2.96
cc_3207 ( N_noxref_12_c_3862_n N_noxref_23_c_7641_n ) capacitor c=7.01366e-19 \
 //x=22.57 //y=2.08 //x2=20.835 //y2=2.96
cc_3208 ( N_noxref_12_c_3884_n N_noxref_23_c_7518_n ) capacitor c=0.00103915f \
 //x=22.685 //y=4.07 //x2=20.72 //y2=2.96
cc_3209 ( N_noxref_12_c_3862_n N_noxref_23_c_7518_n ) capacitor c=0.0148997f \
 //x=22.57 //y=2.08 //x2=20.72 //y2=2.96
cc_3210 ( N_noxref_12_c_3873_n N_noxref_33_c_8593_n ) capacitor c=0.0034165f \
 //x=22.27 //y=1.915 //x2=22.05 //y2=1.505
cc_3211 ( N_noxref_12_c_3862_n N_noxref_33_c_8576_n ) capacitor c=0.0122624f \
 //x=22.57 //y=2.08 //x2=22.935 //y2=1.59
cc_3212 ( N_noxref_12_c_3872_n N_noxref_33_c_8576_n ) capacitor c=0.00703864f \
 //x=22.27 //y=1.53 //x2=22.935 //y2=1.59
cc_3213 ( N_noxref_12_c_3873_n N_noxref_33_c_8576_n ) capacitor c=0.0215834f \
 //x=22.27 //y=1.915 //x2=22.935 //y2=1.59
cc_3214 ( N_noxref_12_c_3875_n N_noxref_33_c_8576_n ) capacitor c=0.00708583f \
 //x=22.645 //y=1.375 //x2=22.935 //y2=1.59
cc_3215 ( N_noxref_12_c_3878_n N_noxref_33_c_8576_n ) capacitor c=0.00698822f \
 //x=22.8 //y=1.22 //x2=22.935 //y2=1.59
cc_3216 ( N_noxref_12_c_3869_n N_noxref_33_M13_noxref_s ) capacitor \
 c=0.0327271f //x=22.27 //y=0.875 //x2=21.915 //y2=0.375
cc_3217 ( N_noxref_12_c_3872_n N_noxref_33_M13_noxref_s ) capacitor \
 c=7.99997e-19 //x=22.27 //y=1.53 //x2=21.915 //y2=0.375
cc_3218 ( N_noxref_12_c_3873_n N_noxref_33_M13_noxref_s ) capacitor \
 c=0.00122123f //x=22.27 //y=1.915 //x2=21.915 //y2=0.375
cc_3219 ( N_noxref_12_c_3876_n N_noxref_33_M13_noxref_s ) capacitor \
 c=0.0121427f //x=22.8 //y=0.875 //x2=21.915 //y2=0.375
cc_3220 ( N_noxref_12_c_3960_n N_noxref_36_c_8740_n ) capacitor c=0.00623646f \
 //x=31.485 //y=1.56 //x2=31.265 //y2=1.495
cc_3221 ( N_noxref_12_c_3965_n N_noxref_36_c_8740_n ) capacitor c=0.00174019f \
 //x=31.45 //y=2.08 //x2=31.265 //y2=1.495
cc_3222 ( N_noxref_12_c_3863_n N_noxref_36_c_8741_n ) capacitor c=0.00158203f \
 //x=31.45 //y=2.08 //x2=32.15 //y2=0.53
cc_3223 ( N_noxref_12_c_3955_n N_noxref_36_c_8741_n ) capacitor c=0.0188655f \
 //x=31.485 //y=0.905 //x2=32.15 //y2=0.53
cc_3224 ( N_noxref_12_c_3963_n N_noxref_36_c_8741_n ) capacitor c=0.00656458f \
 //x=32.015 //y=0.905 //x2=32.15 //y2=0.53
cc_3225 ( N_noxref_12_c_3965_n N_noxref_36_c_8741_n ) capacitor c=2.1838e-19 \
 //x=31.45 //y=2.08 //x2=32.15 //y2=0.53
cc_3226 ( N_noxref_12_c_3955_n N_noxref_36_M18_noxref_s ) capacitor \
 c=0.00623646f //x=31.485 //y=0.905 //x2=30.16 //y2=0.365
cc_3227 ( N_noxref_12_c_3963_n N_noxref_36_M18_noxref_s ) capacitor \
 c=0.0143002f //x=32.015 //y=0.905 //x2=30.16 //y2=0.365
cc_3228 ( N_noxref_12_c_3964_n N_noxref_36_M18_noxref_s ) capacitor \
 c=0.00290153f //x=32.015 //y=1.25 //x2=30.16 //y2=0.365
cc_3229 ( N_noxref_12_c_4059_p N_noxref_37_c_8804_n ) capacitor c=3.15806e-19 \
 //x=35.165 //y=1.655 //x2=33.625 //y2=1.495
cc_3230 ( N_noxref_12_c_4059_p N_noxref_37_c_8792_n ) capacitor c=0.0203424f \
 //x=35.165 //y=1.655 //x2=34.595 //y2=1.495
cc_3231 ( N_noxref_12_c_3865_n N_noxref_37_c_8793_n ) capacitor c=0.00461444f \
 //x=35.435 //y=1.655 //x2=35.48 //y2=0.53
cc_3232 ( N_noxref_12_M21_noxref_d N_noxref_37_c_8793_n ) capacitor \
 c=0.0116735f //x=34.89 //y=0.905 //x2=35.48 //y2=0.53
cc_3233 ( N_noxref_12_c_3865_n N_noxref_37_M20_noxref_s ) capacitor \
 c=0.0137901f //x=35.435 //y=1.655 //x2=33.49 //y2=0.365
cc_3234 ( N_noxref_12_M21_noxref_d N_noxref_37_M20_noxref_s ) capacitor \
 c=0.043966f //x=34.89 //y=0.905 //x2=33.49 //y2=0.365
cc_3235 ( N_noxref_12_c_3865_n N_noxref_38_c_8856_n ) capacitor c=3.22188e-19 \
 //x=35.435 //y=1.655 //x2=36.955 //y2=1.495
cc_3236 ( N_noxref_12_c_4044_n N_noxref_39_c_8898_n ) capacitor c=0.00623646f \
 //x=41.475 //y=1.56 //x2=41.255 //y2=1.495
cc_3237 ( N_noxref_12_c_4049_n N_noxref_39_c_8898_n ) capacitor c=0.00173579f \
 //x=41.44 //y=2.08 //x2=41.255 //y2=1.495
cc_3238 ( N_noxref_12_c_3867_n N_noxref_39_c_8899_n ) capacitor c=0.00156605f \
 //x=41.44 //y=2.08 //x2=42.14 //y2=0.53
cc_3239 ( N_noxref_12_c_4039_n N_noxref_39_c_8899_n ) capacitor c=0.0188655f \
 //x=41.475 //y=0.905 //x2=42.14 //y2=0.53
cc_3240 ( N_noxref_12_c_4047_n N_noxref_39_c_8899_n ) capacitor c=0.00656458f \
 //x=42.005 //y=0.905 //x2=42.14 //y2=0.53
cc_3241 ( N_noxref_12_c_4049_n N_noxref_39_c_8899_n ) capacitor c=2.1838e-19 \
 //x=41.44 //y=2.08 //x2=42.14 //y2=0.53
cc_3242 ( N_noxref_12_c_4039_n N_noxref_39_M24_noxref_s ) capacitor \
 c=0.00623646f //x=41.475 //y=0.905 //x2=40.15 //y2=0.365
cc_3243 ( N_noxref_12_c_4047_n N_noxref_39_M24_noxref_s ) capacitor \
 c=0.0143002f //x=42.005 //y=0.905 //x2=40.15 //y2=0.365
cc_3244 ( N_noxref_12_c_4048_n N_noxref_39_M24_noxref_s ) capacitor \
 c=0.00290153f //x=42.005 //y=1.25 //x2=40.15 //y2=0.365
cc_3245 ( N_D_c_4238_n N_noxref_14_c_4694_n ) capacitor c=0.0245209f \
 //x=49.465 //y=2.59 //x2=50.205 //y2=3.33
cc_3246 ( N_D_c_4257_n N_noxref_14_c_4694_n ) capacitor c=0.0169786f //x=49.58 \
 //y=2.08 //x2=50.205 //y2=3.33
cc_3247 ( N_D_c_4238_n N_noxref_14_c_4696_n ) capacitor c=9.8111e-19 \
 //x=49.465 //y=2.59 //x2=46.365 //y2=3.33
cc_3248 ( N_D_c_4257_n N_noxref_14_c_4697_n ) capacitor c=0.00117715f \
 //x=49.58 //y=2.08 //x2=50.435 //y2=3.33
cc_3249 ( N_D_c_4238_n N_noxref_14_c_4641_n ) capacitor c=0.0179628f \
 //x=49.465 //y=2.59 //x2=46.25 //y2=2.08
cc_3250 ( N_D_c_4465_p N_noxref_14_c_4659_n ) capacitor c=0.0127676f //x=49.58 \
 //y=4.535 //x2=49.755 //y2=5.2
cc_3251 ( N_D_M105_noxref_g N_noxref_14_c_4659_n ) capacitor c=0.0166421f \
 //x=49.62 //y=6.02 //x2=49.755 //y2=5.2
cc_3252 ( N_D_c_4467_p N_noxref_14_c_4659_n ) capacitor c=0.00346527f \
 //x=49.61 //y=4.7 //x2=49.755 //y2=5.2
cc_3253 ( N_D_M106_noxref_g N_noxref_14_c_4665_n ) capacitor c=0.018922f \
 //x=50.06 //y=6.02 //x2=50.235 //y2=5.2
cc_3254 ( N_D_c_4469_p N_noxref_14_c_4642_n ) capacitor c=0.00371277f \
 //x=49.99 //y=1.405 //x2=50.235 //y2=1.655
cc_3255 ( N_D_c_4470_p N_noxref_14_c_4642_n ) capacitor c=0.00457401f \
 //x=50.145 //y=1.25 //x2=50.235 //y2=1.655
cc_3256 ( N_D_c_4238_n N_noxref_14_c_4643_n ) capacitor c=0.00735597f \
 //x=49.465 //y=2.59 //x2=50.32 //y2=3.33
cc_3257 ( N_D_c_4465_p N_noxref_14_c_4643_n ) capacitor c=0.0101284f //x=49.58 \
 //y=4.535 //x2=50.32 //y2=3.33
cc_3258 ( N_D_c_4257_n N_noxref_14_c_4643_n ) capacitor c=0.0663198f //x=49.58 \
 //y=2.08 //x2=50.32 //y2=3.33
cc_3259 ( N_D_c_4474_p N_noxref_14_c_4643_n ) capacitor c=0.0142673f \
 //x=49.985 //y=4.79 //x2=50.32 //y2=3.33
cc_3260 ( N_D_c_4475_p N_noxref_14_c_4643_n ) capacitor c=0.00731987f \
 //x=49.58 //y=2.08 //x2=50.32 //y2=3.33
cc_3261 ( N_D_c_4476_p N_noxref_14_c_4643_n ) capacitor c=0.00306024f \
 //x=49.58 //y=1.915 //x2=50.32 //y2=3.33
cc_3262 ( N_D_c_4467_p N_noxref_14_c_4643_n ) capacitor c=0.00533692f \
 //x=49.61 //y=4.7 //x2=50.32 //y2=3.33
cc_3263 ( N_D_c_4257_n N_noxref_14_c_4644_n ) capacitor c=6.55913e-19 \
 //x=49.58 //y=2.08 //x2=52.17 //y2=2.08
cc_3264 ( N_D_c_4474_p N_noxref_14_c_4713_n ) capacitor c=0.00407665f \
 //x=49.985 //y=4.79 //x2=49.84 //y2=5.2
cc_3265 ( N_D_c_4480_p N_noxref_14_M30_noxref_d ) capacitor c=0.00217566f \
 //x=49.615 //y=0.905 //x2=49.69 //y2=0.905
cc_3266 ( N_D_c_4481_p N_noxref_14_M30_noxref_d ) capacitor c=0.0034598f \
 //x=49.615 //y=1.25 //x2=49.69 //y2=0.905
cc_3267 ( N_D_c_4482_p N_noxref_14_M30_noxref_d ) capacitor c=0.0066953f \
 //x=49.615 //y=1.56 //x2=49.69 //y2=0.905
cc_3268 ( N_D_c_4483_p N_noxref_14_M30_noxref_d ) capacitor c=0.00241102f \
 //x=49.99 //y=0.75 //x2=49.69 //y2=0.905
cc_3269 ( N_D_c_4469_p N_noxref_14_M30_noxref_d ) capacitor c=0.0137169f \
 //x=49.99 //y=1.405 //x2=49.69 //y2=0.905
cc_3270 ( N_D_c_4485_p N_noxref_14_M30_noxref_d ) capacitor c=0.00132245f \
 //x=50.145 //y=0.905 //x2=49.69 //y2=0.905
cc_3271 ( N_D_c_4470_p N_noxref_14_M30_noxref_d ) capacitor c=0.00566463f \
 //x=50.145 //y=1.25 //x2=49.69 //y2=0.905
cc_3272 ( N_D_c_4476_p N_noxref_14_M30_noxref_d ) capacitor c=0.00660593f \
 //x=49.58 //y=1.915 //x2=49.69 //y2=0.905
cc_3273 ( N_D_M105_noxref_g N_noxref_14_M105_noxref_d ) capacitor c=0.0173476f \
 //x=49.62 //y=6.02 //x2=49.695 //y2=5.02
cc_3274 ( N_D_M106_noxref_g N_noxref_14_M105_noxref_d ) capacitor c=0.0179769f \
 //x=50.06 //y=6.02 //x2=49.695 //y2=5.02
cc_3275 ( N_D_c_4289_n N_CLK_c_5034_n ) capacitor c=0.0016972f //x=6.66 \
 //y=4.535 //x2=13.205 //y2=4.44
cc_3276 ( N_D_c_4253_n N_CLK_c_5034_n ) capacitor c=0.0189188f //x=6.66 \
 //y=2.08 //x2=13.205 //y2=4.44
cc_3277 ( N_D_c_4302_n N_CLK_c_5034_n ) capacitor c=0.00960248f //x=7.065 \
 //y=4.79 //x2=13.205 //y2=4.44
cc_3278 ( N_D_c_4313_n N_CLK_c_5034_n ) capacitor c=0.00203982f //x=6.69 \
 //y=4.7 //x2=13.205 //y2=4.44
cc_3279 ( N_D_c_4217_n N_CLK_c_5053_n ) capacitor c=0.00288787f //x=28.005 \
 //y=2.59 //x2=16.745 //y2=4.442
cc_3280 ( N_D_c_4381_n N_CLK_c_5061_n ) capacitor c=0.0016972f //x=28.12 \
 //y=4.535 //x2=34.665 //y2=4.44
cc_3281 ( N_D_c_4255_n N_CLK_c_5061_n ) capacitor c=0.0189188f //x=28.12 \
 //y=2.08 //x2=34.665 //y2=4.44
cc_3282 ( N_D_c_4394_n N_CLK_c_5061_n ) capacitor c=0.00960248f //x=28.525 \
 //y=4.79 //x2=34.665 //y2=4.44
cc_3283 ( N_D_c_4405_n N_CLK_c_5061_n ) capacitor c=0.00203982f //x=28.15 \
 //y=4.7 //x2=34.665 //y2=4.44
cc_3284 ( N_D_c_4217_n N_CLK_c_5079_n ) capacitor c=0.00711882f //x=28.005 \
 //y=2.59 //x2=23.795 //y2=4.44
cc_3285 ( N_D_c_4238_n N_CLK_c_5092_n ) capacitor c=0.00710187f //x=49.465 \
 //y=2.59 //x2=45.025 //y2=4.44
cc_3286 ( N_D_c_4465_p N_CLK_c_5112_n ) capacitor c=0.0016972f //x=49.58 \
 //y=4.535 //x2=56.125 //y2=4.44
cc_3287 ( N_D_c_4257_n N_CLK_c_5112_n ) capacitor c=0.0189188f //x=49.58 \
 //y=2.08 //x2=56.125 //y2=4.44
cc_3288 ( N_D_c_4474_p N_CLK_c_5112_n ) capacitor c=0.00960248f //x=49.985 \
 //y=4.79 //x2=56.125 //y2=4.44
cc_3289 ( N_D_c_4467_p N_CLK_c_5112_n ) capacitor c=0.00203982f //x=49.61 \
 //y=4.7 //x2=56.125 //y2=4.44
cc_3290 ( N_D_c_4217_n N_CLK_c_5026_n ) capacitor c=0.024321f //x=28.005 \
 //y=2.59 //x2=13.32 //y2=2.08
cc_3291 ( N_D_c_4217_n N_CLK_c_5028_n ) capacitor c=0.0225267f //x=28.005 \
 //y=2.59 //x2=23.68 //y2=2.08
cc_3292 ( N_D_c_4238_n N_CLK_c_5029_n ) capacitor c=0.0204615f //x=49.465 \
 //y=2.59 //x2=34.78 //y2=2.08
cc_3293 ( N_D_c_4238_n N_CLK_c_5031_n ) capacitor c=0.0190006f //x=49.465 \
 //y=2.59 //x2=45.14 //y2=2.08
cc_3294 ( N_D_c_4217_n N_CLK_c_5350_n ) capacitor c=0.0030046f //x=28.005 \
 //y=2.59 //x2=23.77 //y2=1.915
cc_3295 ( N_D_c_4217_n N_CLK_c_5222_n ) capacitor c=0.00217166f //x=28.005 \
 //y=2.59 //x2=13.32 //y2=2.08
cc_3296 ( N_D_c_4238_n N_CLK_c_5382_n ) capacitor c=0.00219932f //x=49.465 \
 //y=2.59 //x2=34.78 //y2=2.08
cc_3297 ( N_D_c_4257_n N_noxref_17_c_5847_n ) capacitor c=0.0169594f //x=49.58 \
 //y=2.08 //x2=58.715 //y2=3.7
cc_3298 ( N_D_c_4257_n N_noxref_17_c_5848_n ) capacitor c=0.00131333f \
 //x=49.58 //y=2.08 //x2=48.955 //y2=3.7
cc_3299 ( N_D_c_4238_n N_noxref_17_c_5815_n ) capacitor c=0.0165903f \
 //x=49.465 //y=2.59 //x2=46.99 //y2=3.7
cc_3300 ( N_D_c_4257_n N_noxref_17_c_5815_n ) capacitor c=6.91957e-19 \
 //x=49.58 //y=2.08 //x2=46.99 //y2=3.7
cc_3301 ( N_D_c_4238_n N_noxref_17_c_5778_n ) capacitor c=0.019581f //x=49.465 \
 //y=2.59 //x2=48.84 //y2=2.08
cc_3302 ( N_D_c_4465_p N_noxref_17_c_5778_n ) capacitor c=0.00400249f \
 //x=49.58 //y=4.535 //x2=48.84 //y2=2.08
cc_3303 ( N_D_c_4257_n N_noxref_17_c_5778_n ) capacitor c=0.0706876f //x=49.58 \
 //y=2.08 //x2=48.84 //y2=2.08
cc_3304 ( N_D_c_4475_p N_noxref_17_c_5778_n ) capacitor c=0.00282278f \
 //x=49.58 //y=2.08 //x2=48.84 //y2=2.08
cc_3305 ( N_D_c_4467_p N_noxref_17_c_5778_n ) capacitor c=0.00344981f \
 //x=49.61 //y=4.7 //x2=48.84 //y2=2.08
cc_3306 ( N_D_M105_noxref_g N_noxref_17_M103_noxref_g ) capacitor c=0.0104611f \
 //x=49.62 //y=6.02 //x2=48.74 //y2=6.02
cc_3307 ( N_D_M105_noxref_g N_noxref_17_M104_noxref_g ) capacitor c=0.106811f \
 //x=49.62 //y=6.02 //x2=49.18 //y2=6.02
cc_3308 ( N_D_M106_noxref_g N_noxref_17_M104_noxref_g ) capacitor c=0.0100341f \
 //x=50.06 //y=6.02 //x2=49.18 //y2=6.02
cc_3309 ( N_D_c_4480_p N_noxref_17_c_5780_n ) capacitor c=4.86506e-19 \
 //x=49.615 //y=0.905 //x2=48.645 //y2=0.865
cc_3310 ( N_D_c_4480_p N_noxref_17_c_5782_n ) capacitor c=0.00152104f \
 //x=49.615 //y=0.905 //x2=48.645 //y2=1.21
cc_3311 ( N_D_c_4481_p N_noxref_17_c_5783_n ) capacitor c=0.00109982f \
 //x=49.615 //y=1.25 //x2=48.645 //y2=1.52
cc_3312 ( N_D_c_4482_p N_noxref_17_c_5783_n ) capacitor c=9.57794e-19 \
 //x=49.615 //y=1.56 //x2=48.645 //y2=1.52
cc_3313 ( N_D_c_4257_n N_noxref_17_c_5784_n ) capacitor c=0.00284029f \
 //x=49.58 //y=2.08 //x2=48.645 //y2=1.915
cc_3314 ( N_D_c_4482_p N_noxref_17_c_5784_n ) capacitor c=0.00662747f \
 //x=49.615 //y=1.56 //x2=48.645 //y2=1.915
cc_3315 ( N_D_c_4475_p N_noxref_17_c_5784_n ) capacitor c=0.0172771f //x=49.58 \
 //y=2.08 //x2=48.645 //y2=1.915
cc_3316 ( N_D_c_4480_p N_noxref_17_c_5787_n ) capacitor c=0.0151475f \
 //x=49.615 //y=0.905 //x2=49.175 //y2=0.865
cc_3317 ( N_D_c_4485_p N_noxref_17_c_5787_n ) capacitor c=0.00124821f \
 //x=50.145 //y=0.905 //x2=49.175 //y2=0.865
cc_3318 ( N_D_c_4481_p N_noxref_17_c_5789_n ) capacitor c=0.0111064f \
 //x=49.615 //y=1.25 //x2=49.175 //y2=1.21
cc_3319 ( N_D_c_4482_p N_noxref_17_c_5789_n ) capacitor c=0.00862358f \
 //x=49.615 //y=1.56 //x2=49.175 //y2=1.21
cc_3320 ( N_D_c_4470_p N_noxref_17_c_5789_n ) capacitor c=0.00200715f \
 //x=50.145 //y=1.25 //x2=49.175 //y2=1.21
cc_3321 ( N_D_c_4465_p N_noxref_17_c_5830_n ) capacitor c=0.00417994f \
 //x=49.58 //y=4.535 //x2=48.84 //y2=4.7
cc_3322 ( N_D_c_4467_p N_noxref_17_c_5830_n ) capacitor c=0.0293367f //x=49.61 \
 //y=4.7 //x2=48.84 //y2=4.7
cc_3323 ( N_D_c_4238_n N_noxref_19_c_6210_n ) capacitor c=0.011848f //x=49.465 \
 //y=2.59 //x2=52.795 //y2=4.07
cc_3324 ( N_D_c_4257_n N_noxref_19_c_6210_n ) capacitor c=0.0169317f //x=49.58 \
 //y=2.08 //x2=52.795 //y2=4.07
cc_3325 ( N_D_c_4238_n N_noxref_19_c_6212_n ) capacitor c=4.25679e-19 \
 //x=49.465 //y=2.59 //x2=44.145 //y2=4.07
cc_3326 ( N_D_c_4238_n N_noxref_19_c_6190_n ) capacitor c=0.0188253f \
 //x=49.465 //y=2.59 //x2=44.03 //y2=2.08
cc_3327 ( N_D_c_4238_n N_noxref_21_c_6904_n ) capacitor c=0.333585f //x=49.465 \
 //y=2.59 //x2=42.065 //y2=2.22
cc_3328 ( N_D_c_4238_n N_noxref_21_c_6909_n ) capacitor c=0.0291005f \
 //x=49.465 //y=2.59 //x2=38.225 //y2=2.22
cc_3329 ( N_D_c_4238_n N_noxref_21_c_6911_n ) capacitor c=0.653602f //x=49.465 \
 //y=2.59 //x2=66.115 //y2=2.22
cc_3330 ( N_D_c_4257_n N_noxref_21_c_6911_n ) capacitor c=0.0196864f //x=49.58 \
 //y=2.08 //x2=66.115 //y2=2.22
cc_3331 ( N_D_c_4469_p N_noxref_21_c_6911_n ) capacitor c=3.11115e-19 \
 //x=49.99 //y=1.405 //x2=66.115 //y2=2.22
cc_3332 ( N_D_c_4475_p N_noxref_21_c_6911_n ) capacitor c=0.00570799f \
 //x=49.58 //y=2.08 //x2=66.115 //y2=2.22
cc_3333 ( N_D_c_4238_n N_noxref_21_c_6935_n ) capacitor c=0.0267062f \
 //x=49.465 //y=2.59 //x2=42.295 //y2=2.22
cc_3334 ( N_D_c_4238_n N_noxref_21_c_6939_n ) capacitor c=0.0187633f \
 //x=49.465 //y=2.59 //x2=38.11 //y2=2.08
cc_3335 ( N_D_c_4238_n N_noxref_21_c_6942_n ) capacitor c=0.0184323f \
 //x=49.465 //y=2.59 //x2=42.18 //y2=2.22
cc_3336 ( N_D_c_4217_n N_noxref_23_c_7497_n ) capacitor c=0.334621f //x=28.005 \
 //y=2.59 //x2=20.605 //y2=2.96
cc_3337 ( N_D_c_4217_n N_noxref_23_c_7578_n ) capacitor c=0.0290247f \
 //x=28.005 //y=2.59 //x2=16.765 //y2=2.96
cc_3338 ( N_D_c_4217_n N_noxref_23_c_7498_n ) capacitor c=0.626458f //x=28.005 \
 //y=2.59 //x2=70.185 //y2=2.96
cc_3339 ( N_D_c_4238_n N_noxref_23_c_7498_n ) capacitor c=1.88026f //x=49.465 \
 //y=2.59 //x2=70.185 //y2=2.96
cc_3340 ( N_D_c_4251_n N_noxref_23_c_7498_n ) capacitor c=0.0265274f \
 //x=28.235 //y=2.59 //x2=70.185 //y2=2.96
cc_3341 ( N_D_c_4255_n N_noxref_23_c_7498_n ) capacitor c=0.0187892f //x=28.12 \
 //y=2.08 //x2=70.185 //y2=2.96
cc_3342 ( N_D_c_4257_n N_noxref_23_c_7498_n ) capacitor c=0.0187892f //x=49.58 \
 //y=2.08 //x2=70.185 //y2=2.96
cc_3343 ( N_D_c_4217_n N_noxref_23_c_7641_n ) capacitor c=0.0265752f \
 //x=28.005 //y=2.59 //x2=20.835 //y2=2.96
cc_3344 ( N_D_c_4217_n N_noxref_23_c_7515_n ) capacitor c=0.0222961f \
 //x=28.005 //y=2.59 //x2=16.65 //y2=2.08
cc_3345 ( N_D_c_4217_n N_noxref_23_c_7713_n ) capacitor c=0.0102711f \
 //x=28.005 //y=2.59 //x2=20.365 //y2=1.655
cc_3346 ( N_D_c_4217_n N_noxref_23_c_7518_n ) capacitor c=0.0228944f \
 //x=28.005 //y=2.59 //x2=20.72 //y2=2.96
cc_3347 ( N_D_c_4217_n N_noxref_23_c_7597_n ) capacitor c=0.00219618f \
 //x=28.005 //y=2.59 //x2=16.65 //y2=2.08
cc_3348 ( N_D_c_4236_n N_noxref_28_c_8321_n ) capacitor c=0.00121262f \
 //x=6.775 //y=2.59 //x2=6.475 //y2=1.495
cc_3349 ( N_D_c_4301_n N_noxref_28_c_8321_n ) capacitor c=0.00623646f \
 //x=6.695 //y=1.56 //x2=6.475 //y2=1.495
cc_3350 ( N_D_c_4310_n N_noxref_28_c_8321_n ) capacitor c=0.00174002f //x=6.66 \
 //y=2.08 //x2=6.475 //y2=1.495
cc_3351 ( N_D_c_4217_n N_noxref_28_c_8322_n ) capacitor c=8.64573e-19 \
 //x=28.005 //y=2.59 //x2=7.36 //y2=0.53
cc_3352 ( N_D_c_4236_n N_noxref_28_c_8322_n ) capacitor c=2.73833e-19 \
 //x=6.775 //y=2.59 //x2=7.36 //y2=0.53
cc_3353 ( N_D_c_4253_n N_noxref_28_c_8322_n ) capacitor c=0.00158098f //x=6.66 \
 //y=2.08 //x2=7.36 //y2=0.53
cc_3354 ( N_D_c_4299_n N_noxref_28_c_8322_n ) capacitor c=0.0188655f //x=6.695 \
 //y=0.905 //x2=7.36 //y2=0.53
cc_3355 ( N_D_c_4307_n N_noxref_28_c_8322_n ) capacitor c=0.00656458f \
 //x=7.225 //y=0.905 //x2=7.36 //y2=0.53
cc_3356 ( N_D_c_4310_n N_noxref_28_c_8322_n ) capacitor c=2.1838e-19 //x=6.66 \
 //y=2.08 //x2=7.36 //y2=0.53
cc_3357 ( N_D_c_4217_n N_noxref_28_M3_noxref_s ) capacitor c=8.24206e-19 \
 //x=28.005 //y=2.59 //x2=5.37 //y2=0.365
cc_3358 ( N_D_c_4299_n N_noxref_28_M3_noxref_s ) capacitor c=0.00623646f \
 //x=6.695 //y=0.905 //x2=5.37 //y2=0.365
cc_3359 ( N_D_c_4307_n N_noxref_28_M3_noxref_s ) capacitor c=0.0143002f \
 //x=7.225 //y=0.905 //x2=5.37 //y2=0.365
cc_3360 ( N_D_c_4308_n N_noxref_28_M3_noxref_s ) capacitor c=0.00290153f \
 //x=7.225 //y=1.25 //x2=5.37 //y2=0.365
cc_3361 ( N_D_c_4217_n N_noxref_29_c_8387_n ) capacitor c=0.00444239f \
 //x=28.005 //y=2.59 //x2=8.835 //y2=1.495
cc_3362 ( N_D_c_4217_n N_noxref_29_c_8368_n ) capacitor c=0.0162171f \
 //x=28.005 //y=2.59 //x2=9.72 //y2=1.58
cc_3363 ( N_D_c_4217_n N_noxref_29_c_8375_n ) capacitor c=0.00444239f \
 //x=28.005 //y=2.59 //x2=9.805 //y2=1.495
cc_3364 ( N_D_c_4217_n N_noxref_29_c_8376_n ) capacitor c=0.00112749f \
 //x=28.005 //y=2.59 //x2=10.69 //y2=0.53
cc_3365 ( N_D_c_4217_n N_noxref_29_M5_noxref_s ) capacitor c=8.24206e-19 \
 //x=28.005 //y=2.59 //x2=8.7 //y2=0.365
cc_3366 ( N_D_c_4217_n N_noxref_30_c_8439_n ) capacitor c=0.00444239f \
 //x=28.005 //y=2.59 //x2=12.165 //y2=1.495
cc_3367 ( N_D_c_4217_n N_noxref_30_c_8420_n ) capacitor c=0.0162171f \
 //x=28.005 //y=2.59 //x2=13.05 //y2=1.58
cc_3368 ( N_D_c_4217_n N_noxref_30_c_8427_n ) capacitor c=0.00444239f \
 //x=28.005 //y=2.59 //x2=13.135 //y2=1.495
cc_3369 ( N_D_c_4217_n N_noxref_30_c_8428_n ) capacitor c=0.00112749f \
 //x=28.005 //y=2.59 //x2=14.02 //y2=0.53
cc_3370 ( N_D_c_4217_n N_noxref_30_M7_noxref_s ) capacitor c=8.24206e-19 \
 //x=28.005 //y=2.59 //x2=12.03 //y2=0.365
cc_3371 ( N_D_c_4217_n N_noxref_31_c_8491_n ) capacitor c=0.00444239f \
 //x=28.005 //y=2.59 //x2=15.495 //y2=1.495
cc_3372 ( N_D_c_4217_n N_noxref_31_c_8472_n ) capacitor c=0.0162171f \
 //x=28.005 //y=2.59 //x2=16.38 //y2=1.58
cc_3373 ( N_D_c_4217_n N_noxref_31_c_8479_n ) capacitor c=0.00444239f \
 //x=28.005 //y=2.59 //x2=16.465 //y2=1.495
cc_3374 ( N_D_c_4217_n N_noxref_31_c_8480_n ) capacitor c=0.00112749f \
 //x=28.005 //y=2.59 //x2=17.35 //y2=0.53
cc_3375 ( N_D_c_4217_n N_noxref_31_M9_noxref_s ) capacitor c=8.24206e-19 \
 //x=28.005 //y=2.59 //x2=15.36 //y2=0.365
cc_3376 ( N_D_c_4217_n N_noxref_32_c_8543_n ) capacitor c=0.00444239f \
 //x=28.005 //y=2.59 //x2=18.825 //y2=1.495
cc_3377 ( N_D_c_4217_n N_noxref_32_c_8524_n ) capacitor c=0.0162171f \
 //x=28.005 //y=2.59 //x2=19.71 //y2=1.58
cc_3378 ( N_D_c_4217_n N_noxref_32_c_8531_n ) capacitor c=0.00444239f \
 //x=28.005 //y=2.59 //x2=19.795 //y2=1.495
cc_3379 ( N_D_c_4217_n N_noxref_32_c_8532_n ) capacitor c=0.00112749f \
 //x=28.005 //y=2.59 //x2=20.68 //y2=0.53
cc_3380 ( N_D_c_4217_n N_noxref_32_M11_noxref_s ) capacitor c=8.24206e-19 \
 //x=28.005 //y=2.59 //x2=18.69 //y2=0.365
cc_3381 ( N_D_c_4217_n N_noxref_33_c_8593_n ) capacitor c=0.00448771f \
 //x=28.005 //y=2.59 //x2=22.05 //y2=1.505
cc_3382 ( N_D_c_4217_n N_noxref_33_c_8576_n ) capacitor c=0.0163649f \
 //x=28.005 //y=2.59 //x2=22.935 //y2=1.59
cc_3383 ( N_D_c_4217_n N_noxref_33_c_8605_n ) capacitor c=0.0144126f \
 //x=28.005 //y=2.59 //x2=23.905 //y2=1.59
cc_3384 ( N_D_c_4217_n N_noxref_33_M13_noxref_s ) capacitor c=0.00867201f \
 //x=28.005 //y=2.59 //x2=21.915 //y2=0.375
cc_3385 ( N_D_c_4217_n N_noxref_34_c_8626_n ) capacitor c=0.00494691f \
 //x=28.005 //y=2.59 //x2=24.475 //y2=0.995
cc_3386 ( N_D_c_4217_n N_noxref_34_c_8631_n ) capacitor c=8.29806e-19 \
 //x=28.005 //y=2.59 //x2=25.445 //y2=0.54
cc_3387 ( N_D_c_4217_n N_noxref_34_M15_noxref_s ) capacitor c=0.00448771f \
 //x=28.005 //y=2.59 //x2=24.425 //y2=0.375
cc_3388 ( N_D_c_4217_n N_noxref_35_c_8698_n ) capacitor c=0.00444239f \
 //x=28.005 //y=2.59 //x2=26.965 //y2=1.495
cc_3389 ( N_D_c_4217_n N_noxref_35_c_8679_n ) capacitor c=0.0162171f \
 //x=28.005 //y=2.59 //x2=27.85 //y2=1.58
cc_3390 ( N_D_c_4217_n N_noxref_35_c_8686_n ) capacitor c=0.00404008f \
 //x=28.005 //y=2.59 //x2=27.935 //y2=1.495
cc_3391 ( N_D_c_4251_n N_noxref_35_c_8686_n ) capacitor c=4.2867e-19 \
 //x=28.235 //y=2.59 //x2=27.935 //y2=1.495
cc_3392 ( N_D_c_4393_n N_noxref_35_c_8686_n ) capacitor c=0.00623646f \
 //x=28.155 //y=1.56 //x2=27.935 //y2=1.495
cc_3393 ( N_D_c_4402_n N_noxref_35_c_8686_n ) capacitor c=0.00174002f \
 //x=28.12 //y=2.08 //x2=27.935 //y2=1.495
cc_3394 ( N_D_c_4238_n N_noxref_35_c_8687_n ) capacitor c=8.64573e-19 \
 //x=49.465 //y=2.59 //x2=28.82 //y2=0.53
cc_3395 ( N_D_c_4251_n N_noxref_35_c_8687_n ) capacitor c=2.73833e-19 \
 //x=28.235 //y=2.59 //x2=28.82 //y2=0.53
cc_3396 ( N_D_c_4255_n N_noxref_35_c_8687_n ) capacitor c=0.00158098f \
 //x=28.12 //y=2.08 //x2=28.82 //y2=0.53
cc_3397 ( N_D_c_4391_n N_noxref_35_c_8687_n ) capacitor c=0.0188655f \
 //x=28.155 //y=0.905 //x2=28.82 //y2=0.53
cc_3398 ( N_D_c_4399_n N_noxref_35_c_8687_n ) capacitor c=0.00656458f \
 //x=28.685 //y=0.905 //x2=28.82 //y2=0.53
cc_3399 ( N_D_c_4402_n N_noxref_35_c_8687_n ) capacitor c=2.1838e-19 //x=28.12 \
 //y=2.08 //x2=28.82 //y2=0.53
cc_3400 ( N_D_c_4238_n N_noxref_35_M16_noxref_s ) capacitor c=8.24206e-19 \
 //x=49.465 //y=2.59 //x2=26.83 //y2=0.365
cc_3401 ( N_D_c_4391_n N_noxref_35_M16_noxref_s ) capacitor c=0.00623646f \
 //x=28.155 //y=0.905 //x2=26.83 //y2=0.365
cc_3402 ( N_D_c_4399_n N_noxref_35_M16_noxref_s ) capacitor c=0.0143002f \
 //x=28.685 //y=0.905 //x2=26.83 //y2=0.365
cc_3403 ( N_D_c_4400_n N_noxref_35_M16_noxref_s ) capacitor c=0.00290153f \
 //x=28.685 //y=1.25 //x2=26.83 //y2=0.365
cc_3404 ( N_D_c_4238_n N_noxref_36_c_8752_n ) capacitor c=0.00444239f \
 //x=49.465 //y=2.59 //x2=30.295 //y2=1.495
cc_3405 ( N_D_c_4238_n N_noxref_36_c_8733_n ) capacitor c=0.0162171f \
 //x=49.465 //y=2.59 //x2=31.18 //y2=1.58
cc_3406 ( N_D_c_4238_n N_noxref_36_c_8740_n ) capacitor c=0.00444239f \
 //x=49.465 //y=2.59 //x2=31.265 //y2=1.495
cc_3407 ( N_D_c_4238_n N_noxref_36_c_8741_n ) capacitor c=0.00112749f \
 //x=49.465 //y=2.59 //x2=32.15 //y2=0.53
cc_3408 ( N_D_c_4238_n N_noxref_36_M18_noxref_s ) capacitor c=8.24206e-19 \
 //x=49.465 //y=2.59 //x2=30.16 //y2=0.365
cc_3409 ( N_D_c_4238_n N_noxref_37_c_8804_n ) capacitor c=0.00444239f \
 //x=49.465 //y=2.59 //x2=33.625 //y2=1.495
cc_3410 ( N_D_c_4238_n N_noxref_37_c_8785_n ) capacitor c=0.0162171f \
 //x=49.465 //y=2.59 //x2=34.51 //y2=1.58
cc_3411 ( N_D_c_4238_n N_noxref_37_c_8792_n ) capacitor c=0.00444239f \
 //x=49.465 //y=2.59 //x2=34.595 //y2=1.495
cc_3412 ( N_D_c_4238_n N_noxref_37_c_8793_n ) capacitor c=0.00112749f \
 //x=49.465 //y=2.59 //x2=35.48 //y2=0.53
cc_3413 ( N_D_c_4238_n N_noxref_37_M20_noxref_s ) capacitor c=8.24206e-19 \
 //x=49.465 //y=2.59 //x2=33.49 //y2=0.365
cc_3414 ( N_D_c_4238_n N_noxref_38_c_8856_n ) capacitor c=0.00444239f \
 //x=49.465 //y=2.59 //x2=36.955 //y2=1.495
cc_3415 ( N_D_c_4238_n N_noxref_38_c_8837_n ) capacitor c=0.0162171f \
 //x=49.465 //y=2.59 //x2=37.84 //y2=1.58
cc_3416 ( N_D_c_4238_n N_noxref_38_c_8844_n ) capacitor c=0.00326646f \
 //x=49.465 //y=2.59 //x2=37.925 //y2=1.495
cc_3417 ( N_D_c_4482_p N_noxref_42_c_9055_n ) capacitor c=0.00623646f \
 //x=49.615 //y=1.56 //x2=49.395 //y2=1.495
cc_3418 ( N_D_c_4475_p N_noxref_42_c_9055_n ) capacitor c=0.00173579f \
 //x=49.58 //y=2.08 //x2=49.395 //y2=1.495
cc_3419 ( N_D_c_4257_n N_noxref_42_c_9056_n ) capacitor c=0.00156605f \
 //x=49.58 //y=2.08 //x2=50.28 //y2=0.53
cc_3420 ( N_D_c_4480_p N_noxref_42_c_9056_n ) capacitor c=0.0188655f \
 //x=49.615 //y=0.905 //x2=50.28 //y2=0.53
cc_3421 ( N_D_c_4485_p N_noxref_42_c_9056_n ) capacitor c=0.00656458f \
 //x=50.145 //y=0.905 //x2=50.28 //y2=0.53
cc_3422 ( N_D_c_4475_p N_noxref_42_c_9056_n ) capacitor c=2.1838e-19 //x=49.58 \
 //y=2.08 //x2=50.28 //y2=0.53
cc_3423 ( N_D_c_4480_p N_noxref_42_M29_noxref_s ) capacitor c=0.00623646f \
 //x=49.615 //y=0.905 //x2=48.29 //y2=0.365
cc_3424 ( N_D_c_4485_p N_noxref_42_M29_noxref_s ) capacitor c=0.0143002f \
 //x=50.145 //y=0.905 //x2=48.29 //y2=0.365
cc_3425 ( N_D_c_4470_p N_noxref_42_M29_noxref_s ) capacitor c=0.00290153f \
 //x=50.145 //y=1.25 //x2=48.29 //y2=0.365
cc_3426 ( N_noxref_14_c_4724_p N_noxref_15_c_4921_n ) capacitor c=0.011463f \
 //x=52.055 //y=3.33 //x2=53.765 //y2=3.33
cc_3427 ( N_noxref_14_M108_noxref_g N_noxref_15_c_4890_n ) capacitor \
 c=0.0169521f //x=52.51 //y=6.02 //x2=53.085 //y2=5.2
cc_3428 ( N_noxref_14_c_4644_n N_noxref_15_c_4894_n ) capacitor c=0.00539951f \
 //x=52.17 //y=2.08 //x2=52.375 //y2=5.2
cc_3429 ( N_noxref_14_M107_noxref_g N_noxref_15_c_4894_n ) capacitor \
 c=0.0177326f //x=52.07 //y=6.02 //x2=52.375 //y2=5.2
cc_3430 ( N_noxref_14_c_4682_n N_noxref_15_c_4894_n ) capacitor c=0.00581252f \
 //x=52.17 //y=4.7 //x2=52.375 //y2=5.2
cc_3431 ( N_noxref_14_c_4643_n N_noxref_15_c_4875_n ) capacitor c=3.49822e-19 \
 //x=50.32 //y=3.33 //x2=53.65 //y2=3.33
cc_3432 ( N_noxref_14_c_4644_n N_noxref_15_c_4875_n ) capacitor c=0.0027152f \
 //x=52.17 //y=2.08 //x2=53.65 //y2=3.33
cc_3433 ( N_noxref_14_M108_noxref_g N_noxref_15_M107_noxref_d ) capacitor \
 c=0.0173476f //x=52.51 //y=6.02 //x2=52.145 //y2=5.02
cc_3434 ( N_noxref_14_c_4694_n N_CLK_c_5112_n ) capacitor c=0.00360213f \
 //x=50.205 //y=3.33 //x2=56.125 //y2=4.44
cc_3435 ( N_noxref_14_c_4696_n N_CLK_c_5112_n ) capacitor c=4.49102e-19 \
 //x=46.365 //y=3.33 //x2=56.125 //y2=4.44
cc_3436 ( N_noxref_14_c_4641_n N_CLK_c_5112_n ) capacitor c=0.0200057f \
 //x=46.25 //y=2.08 //x2=56.125 //y2=4.44
cc_3437 ( N_noxref_14_c_4659_n N_CLK_c_5112_n ) capacitor c=0.0185677f \
 //x=49.755 //y=5.2 //x2=56.125 //y2=4.44
cc_3438 ( N_noxref_14_c_4663_n N_CLK_c_5112_n ) capacitor c=0.0181237f \
 //x=49.045 //y=5.2 //x2=56.125 //y2=4.44
cc_3439 ( N_noxref_14_c_4643_n N_CLK_c_5112_n ) capacitor c=0.0208321f \
 //x=50.32 //y=3.33 //x2=56.125 //y2=4.44
cc_3440 ( N_noxref_14_c_4644_n N_CLK_c_5112_n ) capacitor c=0.0198304f \
 //x=52.17 //y=2.08 //x2=56.125 //y2=4.44
cc_3441 ( N_noxref_14_c_4739_p N_CLK_c_5112_n ) capacitor c=0.0111881f \
 //x=46.25 //y=4.7 //x2=56.125 //y2=4.44
cc_3442 ( N_noxref_14_c_4682_n N_CLK_c_5112_n ) capacitor c=0.0107057f \
 //x=52.17 //y=4.7 //x2=56.125 //y2=4.44
cc_3443 ( N_noxref_14_c_4641_n N_CLK_c_5130_n ) capacitor c=0.00153281f \
 //x=46.25 //y=2.08 //x2=45.255 //y2=4.44
cc_3444 ( N_noxref_14_c_4696_n N_CLK_c_5031_n ) capacitor c=0.00526349f \
 //x=46.365 //y=3.33 //x2=45.14 //y2=2.08
cc_3445 ( N_noxref_14_c_4641_n N_CLK_c_5031_n ) capacitor c=0.0443839f \
 //x=46.25 //y=2.08 //x2=45.14 //y2=2.08
cc_3446 ( N_noxref_14_c_4744_p N_CLK_c_5031_n ) capacitor c=0.00201097f \
 //x=46.25 //y=2.08 //x2=45.14 //y2=2.08
cc_3447 ( N_noxref_14_c_4739_p N_CLK_c_5031_n ) capacitor c=0.00218014f \
 //x=46.25 //y=4.7 //x2=45.14 //y2=2.08
cc_3448 ( N_noxref_14_M101_noxref_g N_CLK_M99_noxref_g ) capacitor \
 c=0.0101598f //x=45.99 //y=6.02 //x2=45.11 //y2=6.02
cc_3449 ( N_noxref_14_M101_noxref_g N_CLK_M100_noxref_g ) capacitor \
 c=0.0602553f //x=45.99 //y=6.02 //x2=45.55 //y2=6.02
cc_3450 ( N_noxref_14_M102_noxref_g N_CLK_M100_noxref_g ) capacitor \
 c=0.0101598f //x=46.43 //y=6.02 //x2=45.55 //y2=6.02
cc_3451 ( N_noxref_14_c_4749_p N_CLK_c_5529_n ) capacitor c=0.00456962f \
 //x=46.24 //y=0.915 //x2=45.23 //y2=0.91
cc_3452 ( N_noxref_14_c_4750_p N_CLK_c_5530_n ) capacitor c=0.00438372f \
 //x=46.24 //y=1.26 //x2=45.23 //y2=1.22
cc_3453 ( N_noxref_14_c_4751_p N_CLK_c_5531_n ) capacitor c=0.00438372f \
 //x=46.24 //y=1.57 //x2=45.23 //y2=1.45
cc_3454 ( N_noxref_14_c_4641_n N_CLK_c_5532_n ) capacitor c=0.00205895f \
 //x=46.25 //y=2.08 //x2=45.23 //y2=1.915
cc_3455 ( N_noxref_14_c_4744_p N_CLK_c_5532_n ) capacitor c=0.00828003f \
 //x=46.25 //y=2.08 //x2=45.23 //y2=1.915
cc_3456 ( N_noxref_14_c_4754_p N_CLK_c_5532_n ) capacitor c=0.00438372f \
 //x=46.25 //y=1.915 //x2=45.23 //y2=1.915
cc_3457 ( N_noxref_14_c_4739_p N_CLK_c_5535_n ) capacitor c=0.0611812f \
 //x=46.25 //y=4.7 //x2=45.475 //y2=4.79
cc_3458 ( N_noxref_14_c_4641_n N_CLK_c_5536_n ) capacitor c=0.00142741f \
 //x=46.25 //y=2.08 //x2=45.14 //y2=4.7
cc_3459 ( N_noxref_14_c_4739_p N_CLK_c_5536_n ) capacitor c=0.00487508f \
 //x=46.25 //y=4.7 //x2=45.14 //y2=4.7
cc_3460 ( N_noxref_14_c_4694_n N_noxref_17_c_5873_n ) capacitor c=0.146341f \
 //x=50.205 //y=3.33 //x2=48.725 //y2=3.7
cc_3461 ( N_noxref_14_c_4694_n N_noxref_17_c_5874_n ) capacitor c=0.0294746f \
 //x=50.205 //y=3.33 //x2=47.105 //y2=3.7
cc_3462 ( N_noxref_14_c_4641_n N_noxref_17_c_5874_n ) capacitor c=0.00687545f \
 //x=46.25 //y=2.08 //x2=47.105 //y2=3.7
cc_3463 ( N_noxref_14_c_4694_n N_noxref_17_c_5847_n ) capacitor c=0.108749f \
 //x=50.205 //y=3.33 //x2=58.715 //y2=3.7
cc_3464 ( N_noxref_14_c_4724_p N_noxref_17_c_5847_n ) capacitor c=0.175696f \
 //x=52.055 //y=3.33 //x2=58.715 //y2=3.7
cc_3465 ( N_noxref_14_c_4697_n N_noxref_17_c_5847_n ) capacitor c=0.0267668f \
 //x=50.435 //y=3.33 //x2=58.715 //y2=3.7
cc_3466 ( N_noxref_14_c_4643_n N_noxref_17_c_5847_n ) capacitor c=0.0206034f \
 //x=50.32 //y=3.33 //x2=58.715 //y2=3.7
cc_3467 ( N_noxref_14_c_4644_n N_noxref_17_c_5847_n ) capacitor c=0.0205831f \
 //x=52.17 //y=2.08 //x2=58.715 //y2=3.7
cc_3468 ( N_noxref_14_c_4694_n N_noxref_17_c_5848_n ) capacitor c=0.0266674f \
 //x=50.205 //y=3.33 //x2=48.955 //y2=3.7
cc_3469 ( N_noxref_14_M101_noxref_g N_noxref_17_c_5807_n ) capacitor \
 c=0.01736f //x=45.99 //y=6.02 //x2=46.125 //y2=5.155
cc_3470 ( N_noxref_14_M102_noxref_g N_noxref_17_c_5811_n ) capacitor \
 c=0.0194981f //x=46.43 //y=6.02 //x2=46.905 //y2=5.155
cc_3471 ( N_noxref_14_c_4739_p N_noxref_17_c_5811_n ) capacitor c=0.00201851f \
 //x=46.25 //y=4.7 //x2=46.905 //y2=5.155
cc_3472 ( N_noxref_14_c_4770_p N_noxref_17_c_5777_n ) capacitor c=0.00371277f \
 //x=46.615 //y=1.415 //x2=46.905 //y2=1.665
cc_3473 ( N_noxref_14_c_4771_p N_noxref_17_c_5777_n ) capacitor c=0.00457401f \
 //x=46.77 //y=1.26 //x2=46.905 //y2=1.665
cc_3474 ( N_noxref_14_c_4694_n N_noxref_17_c_5815_n ) capacitor c=0.0206036f \
 //x=50.205 //y=3.33 //x2=46.99 //y2=3.7
cc_3475 ( N_noxref_14_c_4696_n N_noxref_17_c_5815_n ) capacitor c=0.00117715f \
 //x=46.365 //y=3.33 //x2=46.99 //y2=3.7
cc_3476 ( N_noxref_14_c_4641_n N_noxref_17_c_5815_n ) capacitor c=0.0759508f \
 //x=46.25 //y=2.08 //x2=46.99 //y2=3.7
cc_3477 ( N_noxref_14_c_4643_n N_noxref_17_c_5815_n ) capacitor c=3.52729e-19 \
 //x=50.32 //y=3.33 //x2=46.99 //y2=3.7
cc_3478 ( N_noxref_14_c_4744_p N_noxref_17_c_5815_n ) capacitor c=0.00731987f \
 //x=46.25 //y=2.08 //x2=46.99 //y2=3.7
cc_3479 ( N_noxref_14_c_4754_p N_noxref_17_c_5815_n ) capacitor c=0.00283672f \
 //x=46.25 //y=1.915 //x2=46.99 //y2=3.7
cc_3480 ( N_noxref_14_c_4739_p N_noxref_17_c_5815_n ) capacitor c=0.013693f \
 //x=46.25 //y=4.7 //x2=46.99 //y2=3.7
cc_3481 ( N_noxref_14_c_4694_n N_noxref_17_c_5778_n ) capacitor c=0.020575f \
 //x=50.205 //y=3.33 //x2=48.84 //y2=2.08
cc_3482 ( N_noxref_14_c_4641_n N_noxref_17_c_5778_n ) capacitor c=8.46099e-19 \
 //x=46.25 //y=2.08 //x2=48.84 //y2=2.08
cc_3483 ( N_noxref_14_c_4663_n N_noxref_17_c_5778_n ) capacitor c=0.00521572f \
 //x=49.045 //y=5.2 //x2=48.84 //y2=2.08
cc_3484 ( N_noxref_14_c_4643_n N_noxref_17_c_5778_n ) capacitor c=0.00289219f \
 //x=50.32 //y=3.33 //x2=48.84 //y2=2.08
cc_3485 ( N_noxref_14_c_4641_n N_noxref_17_c_5898_n ) capacitor c=0.0166016f \
 //x=46.25 //y=2.08 //x2=46.21 //y2=5.155
cc_3486 ( N_noxref_14_c_4739_p N_noxref_17_c_5898_n ) capacitor c=0.00475601f \
 //x=46.25 //y=4.7 //x2=46.21 //y2=5.155
cc_3487 ( N_noxref_14_c_4663_n N_noxref_17_M103_noxref_g ) capacitor \
 c=0.0177326f //x=49.045 //y=5.2 //x2=48.74 //y2=6.02
cc_3488 ( N_noxref_14_c_4659_n N_noxref_17_M104_noxref_g ) capacitor \
 c=0.0169521f //x=49.755 //y=5.2 //x2=49.18 //y2=6.02
cc_3489 ( N_noxref_14_M103_noxref_d N_noxref_17_M104_noxref_g ) capacitor \
 c=0.0173476f //x=48.815 //y=5.02 //x2=49.18 //y2=6.02
cc_3490 ( N_noxref_14_c_4663_n N_noxref_17_c_5830_n ) capacitor c=0.00581252f \
 //x=49.045 //y=5.2 //x2=48.84 //y2=4.7
cc_3491 ( N_noxref_14_c_4749_p N_noxref_17_M28_noxref_d ) capacitor \
 c=0.00217566f //x=46.24 //y=0.915 //x2=46.315 //y2=0.915
cc_3492 ( N_noxref_14_c_4750_p N_noxref_17_M28_noxref_d ) capacitor \
 c=0.0034598f //x=46.24 //y=1.26 //x2=46.315 //y2=0.915
cc_3493 ( N_noxref_14_c_4751_p N_noxref_17_M28_noxref_d ) capacitor \
 c=0.00546784f //x=46.24 //y=1.57 //x2=46.315 //y2=0.915
cc_3494 ( N_noxref_14_c_4792_p N_noxref_17_M28_noxref_d ) capacitor \
 c=0.00241102f //x=46.615 //y=0.76 //x2=46.315 //y2=0.915
cc_3495 ( N_noxref_14_c_4770_p N_noxref_17_M28_noxref_d ) capacitor \
 c=0.0138621f //x=46.615 //y=1.415 //x2=46.315 //y2=0.915
cc_3496 ( N_noxref_14_c_4794_p N_noxref_17_M28_noxref_d ) capacitor \
 c=0.00219619f //x=46.77 //y=0.915 //x2=46.315 //y2=0.915
cc_3497 ( N_noxref_14_c_4771_p N_noxref_17_M28_noxref_d ) capacitor \
 c=0.00603828f //x=46.77 //y=1.26 //x2=46.315 //y2=0.915
cc_3498 ( N_noxref_14_c_4754_p N_noxref_17_M28_noxref_d ) capacitor \
 c=0.00661782f //x=46.25 //y=1.915 //x2=46.315 //y2=0.915
cc_3499 ( N_noxref_14_M101_noxref_g N_noxref_17_M101_noxref_d ) capacitor \
 c=0.0180032f //x=45.99 //y=6.02 //x2=46.065 //y2=5.02
cc_3500 ( N_noxref_14_M102_noxref_g N_noxref_17_M101_noxref_d ) capacitor \
 c=0.0194246f //x=46.43 //y=6.02 //x2=46.065 //y2=5.02
cc_3501 ( N_noxref_14_c_4694_n N_noxref_19_c_6210_n ) capacitor c=0.0428508f \
 //x=50.205 //y=3.33 //x2=52.795 //y2=4.07
cc_3502 ( N_noxref_14_c_4696_n N_noxref_19_c_6210_n ) capacitor c=0.0135672f \
 //x=46.365 //y=3.33 //x2=52.795 //y2=4.07
cc_3503 ( N_noxref_14_c_4724_p N_noxref_19_c_6210_n ) capacitor c=0.0110241f \
 //x=52.055 //y=3.33 //x2=52.795 //y2=4.07
cc_3504 ( N_noxref_14_c_4697_n N_noxref_19_c_6210_n ) capacitor c=5.70661e-19 \
 //x=50.435 //y=3.33 //x2=52.795 //y2=4.07
cc_3505 ( N_noxref_14_c_4641_n N_noxref_19_c_6210_n ) capacitor c=0.0206302f \
 //x=46.25 //y=2.08 //x2=52.795 //y2=4.07
cc_3506 ( N_noxref_14_c_4643_n N_noxref_19_c_6210_n ) capacitor c=0.0181936f \
 //x=50.32 //y=3.33 //x2=52.795 //y2=4.07
cc_3507 ( N_noxref_14_c_4644_n N_noxref_19_c_6210_n ) capacitor c=0.0184765f \
 //x=52.17 //y=2.08 //x2=52.795 //y2=4.07
cc_3508 ( N_noxref_14_c_4644_n N_noxref_19_c_6284_n ) capacitor c=0.00179385f \
 //x=52.17 //y=2.08 //x2=53.025 //y2=4.07
cc_3509 ( N_noxref_14_c_4641_n N_noxref_19_c_6190_n ) capacitor c=0.00133538f \
 //x=46.25 //y=2.08 //x2=44.03 //y2=2.08
cc_3510 ( N_noxref_14_c_4644_n N_noxref_19_c_6286_n ) capacitor c=0.00400249f \
 //x=52.17 //y=2.08 //x2=52.91 //y2=4.535
cc_3511 ( N_noxref_14_c_4682_n N_noxref_19_c_6286_n ) capacitor c=0.00417994f \
 //x=52.17 //y=4.7 //x2=52.91 //y2=4.535
cc_3512 ( N_noxref_14_c_4724_p N_noxref_19_c_6191_n ) capacitor c=0.00318578f \
 //x=52.055 //y=3.33 //x2=52.91 //y2=2.08
cc_3513 ( N_noxref_14_c_4643_n N_noxref_19_c_6191_n ) capacitor c=8.48165e-19 \
 //x=50.32 //y=3.33 //x2=52.91 //y2=2.08
cc_3514 ( N_noxref_14_c_4644_n N_noxref_19_c_6191_n ) capacitor c=0.0743965f \
 //x=52.17 //y=2.08 //x2=52.91 //y2=2.08
cc_3515 ( N_noxref_14_c_4649_n N_noxref_19_c_6191_n ) capacitor c=0.00284029f \
 //x=51.975 //y=1.915 //x2=52.91 //y2=2.08
cc_3516 ( N_noxref_14_M107_noxref_g N_noxref_19_M109_noxref_g ) capacitor \
 c=0.0104611f //x=52.07 //y=6.02 //x2=52.95 //y2=6.02
cc_3517 ( N_noxref_14_M108_noxref_g N_noxref_19_M109_noxref_g ) capacitor \
 c=0.106811f //x=52.51 //y=6.02 //x2=52.95 //y2=6.02
cc_3518 ( N_noxref_14_M108_noxref_g N_noxref_19_M110_noxref_g ) capacitor \
 c=0.0100341f //x=52.51 //y=6.02 //x2=53.39 //y2=6.02
cc_3519 ( N_noxref_14_c_4645_n N_noxref_19_c_6295_n ) capacitor c=4.86506e-19 \
 //x=51.975 //y=0.865 //x2=52.945 //y2=0.905
cc_3520 ( N_noxref_14_c_4647_n N_noxref_19_c_6295_n ) capacitor c=0.00152104f \
 //x=51.975 //y=1.21 //x2=52.945 //y2=0.905
cc_3521 ( N_noxref_14_c_4652_n N_noxref_19_c_6295_n ) capacitor c=0.0151475f \
 //x=52.505 //y=0.865 //x2=52.945 //y2=0.905
cc_3522 ( N_noxref_14_c_4648_n N_noxref_19_c_6298_n ) capacitor c=0.00109982f \
 //x=51.975 //y=1.52 //x2=52.945 //y2=1.25
cc_3523 ( N_noxref_14_c_4654_n N_noxref_19_c_6298_n ) capacitor c=0.0111064f \
 //x=52.505 //y=1.21 //x2=52.945 //y2=1.25
cc_3524 ( N_noxref_14_c_4648_n N_noxref_19_c_6300_n ) capacitor c=9.57794e-19 \
 //x=51.975 //y=1.52 //x2=52.945 //y2=1.56
cc_3525 ( N_noxref_14_c_4649_n N_noxref_19_c_6300_n ) capacitor c=0.00662747f \
 //x=51.975 //y=1.915 //x2=52.945 //y2=1.56
cc_3526 ( N_noxref_14_c_4654_n N_noxref_19_c_6300_n ) capacitor c=0.00862358f \
 //x=52.505 //y=1.21 //x2=52.945 //y2=1.56
cc_3527 ( N_noxref_14_c_4652_n N_noxref_19_c_6303_n ) capacitor c=0.00124821f \
 //x=52.505 //y=0.865 //x2=53.475 //y2=0.905
cc_3528 ( N_noxref_14_c_4654_n N_noxref_19_c_6304_n ) capacitor c=0.00200715f \
 //x=52.505 //y=1.21 //x2=53.475 //y2=1.25
cc_3529 ( N_noxref_14_c_4644_n N_noxref_19_c_6305_n ) capacitor c=0.00282278f \
 //x=52.17 //y=2.08 //x2=52.91 //y2=2.08
cc_3530 ( N_noxref_14_c_4649_n N_noxref_19_c_6305_n ) capacitor c=0.0172771f \
 //x=51.975 //y=1.915 //x2=52.91 //y2=2.08
cc_3531 ( N_noxref_14_c_4644_n N_noxref_19_c_6307_n ) capacitor c=0.00344981f \
 //x=52.17 //y=2.08 //x2=52.94 //y2=4.7
cc_3532 ( N_noxref_14_c_4682_n N_noxref_19_c_6307_n ) capacitor c=0.0293367f \
 //x=52.17 //y=4.7 //x2=52.94 //y2=4.7
cc_3533 ( N_noxref_14_c_4694_n N_noxref_21_c_6911_n ) capacitor c=0.00374806f \
 //x=50.205 //y=3.33 //x2=66.115 //y2=2.22
cc_3534 ( N_noxref_14_c_4724_p N_noxref_21_c_6911_n ) capacitor c=0.0102155f \
 //x=52.055 //y=3.33 //x2=66.115 //y2=2.22
cc_3535 ( N_noxref_14_c_4697_n N_noxref_21_c_6911_n ) capacitor c=4.47816e-19 \
 //x=50.435 //y=3.33 //x2=66.115 //y2=2.22
cc_3536 ( N_noxref_14_c_4641_n N_noxref_21_c_6911_n ) capacitor c=0.0186201f \
 //x=46.25 //y=2.08 //x2=66.115 //y2=2.22
cc_3537 ( N_noxref_14_c_4835_p N_noxref_21_c_6911_n ) capacitor c=0.0146822f \
 //x=49.965 //y=1.655 //x2=66.115 //y2=2.22
cc_3538 ( N_noxref_14_c_4643_n N_noxref_21_c_6911_n ) capacitor c=0.0222456f \
 //x=50.32 //y=3.33 //x2=66.115 //y2=2.22
cc_3539 ( N_noxref_14_c_4644_n N_noxref_21_c_6911_n ) capacitor c=0.0208418f \
 //x=52.17 //y=2.08 //x2=66.115 //y2=2.22
cc_3540 ( N_noxref_14_c_4770_p N_noxref_21_c_6911_n ) capacitor c=3.13485e-19 \
 //x=46.615 //y=1.415 //x2=66.115 //y2=2.22
cc_3541 ( N_noxref_14_c_4649_n N_noxref_21_c_6911_n ) capacitor c=0.00894156f \
 //x=51.975 //y=1.915 //x2=66.115 //y2=2.22
cc_3542 ( N_noxref_14_c_4744_p N_noxref_21_c_6911_n ) capacitor c=0.00584491f \
 //x=46.25 //y=2.08 //x2=66.115 //y2=2.22
cc_3543 ( N_noxref_14_c_4694_n N_noxref_23_c_7498_n ) capacitor c=0.336622f \
 //x=50.205 //y=3.33 //x2=70.185 //y2=2.96
cc_3544 ( N_noxref_14_c_4696_n N_noxref_23_c_7498_n ) capacitor c=0.0291389f \
 //x=46.365 //y=3.33 //x2=70.185 //y2=2.96
cc_3545 ( N_noxref_14_c_4724_p N_noxref_23_c_7498_n ) capacitor c=0.173509f \
 //x=52.055 //y=3.33 //x2=70.185 //y2=2.96
cc_3546 ( N_noxref_14_c_4697_n N_noxref_23_c_7498_n ) capacitor c=0.0266415f \
 //x=50.435 //y=3.33 //x2=70.185 //y2=2.96
cc_3547 ( N_noxref_14_c_4641_n N_noxref_23_c_7498_n ) capacitor c=0.0198264f \
 //x=46.25 //y=2.08 //x2=70.185 //y2=2.96
cc_3548 ( N_noxref_14_c_4643_n N_noxref_23_c_7498_n ) capacitor c=0.0229357f \
 //x=50.32 //y=3.33 //x2=70.185 //y2=2.96
cc_3549 ( N_noxref_14_c_4644_n N_noxref_23_c_7498_n ) capacitor c=0.0228696f \
 //x=52.17 //y=2.08 //x2=70.185 //y2=2.96
cc_3550 ( N_noxref_14_c_4641_n N_noxref_41_c_9000_n ) capacitor c=0.00204385f \
 //x=46.25 //y=2.08 //x2=46.905 //y2=0.54
cc_3551 ( N_noxref_14_c_4749_p N_noxref_41_c_9000_n ) capacitor c=0.0194423f \
 //x=46.24 //y=0.915 //x2=46.905 //y2=0.54
cc_3552 ( N_noxref_14_c_4794_p N_noxref_41_c_9000_n ) capacitor c=0.00656458f \
 //x=46.77 //y=0.915 //x2=46.905 //y2=0.54
cc_3553 ( N_noxref_14_c_4744_p N_noxref_41_c_9000_n ) capacitor c=2.20712e-19 \
 //x=46.25 //y=2.08 //x2=46.905 //y2=0.54
cc_3554 ( N_noxref_14_c_4750_p N_noxref_41_c_9013_n ) capacitor c=0.00538829f \
 //x=46.24 //y=1.26 //x2=46.02 //y2=0.995
cc_3555 ( N_noxref_14_c_4749_p N_noxref_41_M28_noxref_s ) capacitor \
 c=0.00538829f //x=46.24 //y=0.915 //x2=45.885 //y2=0.375
cc_3556 ( N_noxref_14_c_4751_p N_noxref_41_M28_noxref_s ) capacitor \
 c=0.00538829f //x=46.24 //y=1.57 //x2=45.885 //y2=0.375
cc_3557 ( N_noxref_14_c_4794_p N_noxref_41_M28_noxref_s ) capacitor \
 c=0.0143002f //x=46.77 //y=0.915 //x2=45.885 //y2=0.375
cc_3558 ( N_noxref_14_c_4771_p N_noxref_41_M28_noxref_s ) capacitor \
 c=0.00290153f //x=46.77 //y=1.26 //x2=45.885 //y2=0.375
cc_3559 ( N_noxref_14_c_4835_p N_noxref_42_c_9076_n ) capacitor c=3.15806e-19 \
 //x=49.965 //y=1.655 //x2=48.425 //y2=1.495
cc_3560 ( N_noxref_14_c_4835_p N_noxref_42_c_9055_n ) capacitor c=0.020324f \
 //x=49.965 //y=1.655 //x2=49.395 //y2=1.495
cc_3561 ( N_noxref_14_c_4642_n N_noxref_42_c_9056_n ) capacitor c=0.00457164f \
 //x=50.235 //y=1.655 //x2=50.28 //y2=0.53
cc_3562 ( N_noxref_14_M30_noxref_d N_noxref_42_c_9056_n ) capacitor \
 c=0.0115831f //x=49.69 //y=0.905 //x2=50.28 //y2=0.53
cc_3563 ( N_noxref_14_c_4642_n N_noxref_42_M29_noxref_s ) capacitor \
 c=0.013435f //x=50.235 //y=1.655 //x2=48.29 //y2=0.365
cc_3564 ( N_noxref_14_M30_noxref_d N_noxref_42_M29_noxref_s ) capacitor \
 c=0.0439476f //x=49.69 //y=0.905 //x2=48.29 //y2=0.365
cc_3565 ( N_noxref_14_c_4642_n N_noxref_43_c_9119_n ) capacitor c=3.22188e-19 \
 //x=50.235 //y=1.655 //x2=51.755 //y2=1.495
cc_3566 ( N_noxref_14_c_4649_n N_noxref_43_c_9119_n ) capacitor c=0.0034165f \
 //x=51.975 //y=1.915 //x2=51.755 //y2=1.495
cc_3567 ( N_noxref_14_c_4644_n N_noxref_43_c_9100_n ) capacitor c=0.011618f \
 //x=52.17 //y=2.08 //x2=52.64 //y2=1.58
cc_3568 ( N_noxref_14_c_4648_n N_noxref_43_c_9100_n ) capacitor c=0.00696403f \
 //x=51.975 //y=1.52 //x2=52.64 //y2=1.58
cc_3569 ( N_noxref_14_c_4649_n N_noxref_43_c_9100_n ) capacitor c=0.0174694f \
 //x=51.975 //y=1.915 //x2=52.64 //y2=1.58
cc_3570 ( N_noxref_14_c_4651_n N_noxref_43_c_9100_n ) capacitor c=0.00776811f \
 //x=52.35 //y=1.365 //x2=52.64 //y2=1.58
cc_3571 ( N_noxref_14_c_4654_n N_noxref_43_c_9100_n ) capacitor c=0.00339872f \
 //x=52.505 //y=1.21 //x2=52.64 //y2=1.58
cc_3572 ( N_noxref_14_c_4649_n N_noxref_43_c_9107_n ) capacitor c=6.71402e-19 \
 //x=51.975 //y=1.915 //x2=52.725 //y2=1.495
cc_3573 ( N_noxref_14_c_4645_n N_noxref_43_M31_noxref_s ) capacitor \
 c=0.0326577f //x=51.975 //y=0.865 //x2=51.62 //y2=0.365
cc_3574 ( N_noxref_14_c_4648_n N_noxref_43_M31_noxref_s ) capacitor \
 c=3.48408e-19 //x=51.975 //y=1.52 //x2=51.62 //y2=0.365
cc_3575 ( N_noxref_14_c_4652_n N_noxref_43_M31_noxref_s ) capacitor \
 c=0.0120759f //x=52.505 //y=0.865 //x2=51.62 //y2=0.365
cc_3576 ( N_noxref_15_c_4890_n N_CLK_c_5112_n ) capacitor c=0.0185297f \
 //x=53.085 //y=5.2 //x2=56.125 //y2=4.44
cc_3577 ( N_noxref_15_c_4894_n N_CLK_c_5112_n ) capacitor c=0.018142f \
 //x=52.375 //y=5.2 //x2=56.125 //y2=4.44
cc_3578 ( N_noxref_15_c_4875_n N_CLK_c_5112_n ) capacitor c=0.0208321f \
 //x=53.65 //y=3.33 //x2=56.125 //y2=4.44
cc_3579 ( N_noxref_15_c_4876_n N_CLK_c_5112_n ) capacitor c=0.0215137f \
 //x=55.5 //y=2.08 //x2=56.125 //y2=4.44
cc_3580 ( N_noxref_15_c_4909_n N_CLK_c_5112_n ) capacitor c=0.0109968f \
 //x=55.5 //y=4.7 //x2=56.125 //y2=4.44
cc_3581 ( N_noxref_15_c_4876_n N_CLK_c_5543_n ) capacitor c=0.00400249f \
 //x=55.5 //y=2.08 //x2=56.24 //y2=4.535
cc_3582 ( N_noxref_15_c_4909_n N_CLK_c_5543_n ) capacitor c=0.00415951f \
 //x=55.5 //y=4.7 //x2=56.24 //y2=4.535
cc_3583 ( N_noxref_15_c_4936_p N_CLK_c_5032_n ) capacitor c=0.00720056f \
 //x=55.385 //y=3.33 //x2=56.24 //y2=2.08
cc_3584 ( N_noxref_15_c_4875_n N_CLK_c_5032_n ) capacitor c=9.02527e-19 \
 //x=53.65 //y=3.33 //x2=56.24 //y2=2.08
cc_3585 ( N_noxref_15_c_4876_n N_CLK_c_5032_n ) capacitor c=0.0737918f \
 //x=55.5 //y=2.08 //x2=56.24 //y2=2.08
cc_3586 ( N_noxref_15_c_4881_n N_CLK_c_5032_n ) capacitor c=0.00284029f \
 //x=55.305 //y=1.915 //x2=56.24 //y2=2.08
cc_3587 ( N_noxref_15_M111_noxref_g N_CLK_M113_noxref_g ) capacitor \
 c=0.0104611f //x=55.4 //y=6.02 //x2=56.28 //y2=6.02
cc_3588 ( N_noxref_15_M112_noxref_g N_CLK_M113_noxref_g ) capacitor \
 c=0.106811f //x=55.84 //y=6.02 //x2=56.28 //y2=6.02
cc_3589 ( N_noxref_15_M112_noxref_g N_CLK_M114_noxref_g ) capacitor \
 c=0.0100341f //x=55.84 //y=6.02 //x2=56.72 //y2=6.02
cc_3590 ( N_noxref_15_c_4877_n N_CLK_c_5552_n ) capacitor c=4.86506e-19 \
 //x=55.305 //y=0.865 //x2=56.275 //y2=0.905
cc_3591 ( N_noxref_15_c_4879_n N_CLK_c_5552_n ) capacitor c=0.00152104f \
 //x=55.305 //y=1.21 //x2=56.275 //y2=0.905
cc_3592 ( N_noxref_15_c_4884_n N_CLK_c_5552_n ) capacitor c=0.0151475f \
 //x=55.835 //y=0.865 //x2=56.275 //y2=0.905
cc_3593 ( N_noxref_15_c_4880_n N_CLK_c_5555_n ) capacitor c=0.00109982f \
 //x=55.305 //y=1.52 //x2=56.275 //y2=1.25
cc_3594 ( N_noxref_15_c_4886_n N_CLK_c_5555_n ) capacitor c=0.0111064f \
 //x=55.835 //y=1.21 //x2=56.275 //y2=1.25
cc_3595 ( N_noxref_15_c_4880_n N_CLK_c_5557_n ) capacitor c=9.57794e-19 \
 //x=55.305 //y=1.52 //x2=56.275 //y2=1.56
cc_3596 ( N_noxref_15_c_4881_n N_CLK_c_5557_n ) capacitor c=0.00662747f \
 //x=55.305 //y=1.915 //x2=56.275 //y2=1.56
cc_3597 ( N_noxref_15_c_4886_n N_CLK_c_5557_n ) capacitor c=0.00862358f \
 //x=55.835 //y=1.21 //x2=56.275 //y2=1.56
cc_3598 ( N_noxref_15_c_4884_n N_CLK_c_5560_n ) capacitor c=0.00124821f \
 //x=55.835 //y=0.865 //x2=56.805 //y2=0.905
cc_3599 ( N_noxref_15_c_4886_n N_CLK_c_5561_n ) capacitor c=0.00200715f \
 //x=55.835 //y=1.21 //x2=56.805 //y2=1.25
cc_3600 ( N_noxref_15_c_4876_n N_CLK_c_5562_n ) capacitor c=0.00282278f \
 //x=55.5 //y=2.08 //x2=56.24 //y2=2.08
cc_3601 ( N_noxref_15_c_4881_n N_CLK_c_5562_n ) capacitor c=0.0172771f \
 //x=55.305 //y=1.915 //x2=56.24 //y2=2.08
cc_3602 ( N_noxref_15_c_4876_n N_CLK_c_5564_n ) capacitor c=0.00342116f \
 //x=55.5 //y=2.08 //x2=56.27 //y2=4.7
cc_3603 ( N_noxref_15_c_4909_n N_CLK_c_5564_n ) capacitor c=0.0292158f \
 //x=55.5 //y=4.7 //x2=56.27 //y2=4.7
cc_3604 ( N_noxref_15_c_4936_p N_noxref_17_c_5847_n ) capacitor c=0.175696f \
 //x=55.385 //y=3.33 //x2=58.715 //y2=3.7
cc_3605 ( N_noxref_15_c_4921_n N_noxref_17_c_5847_n ) capacitor c=0.0293967f \
 //x=53.765 //y=3.33 //x2=58.715 //y2=3.7
cc_3606 ( N_noxref_15_c_4875_n N_noxref_17_c_5847_n ) capacitor c=0.0206034f \
 //x=53.65 //y=3.33 //x2=58.715 //y2=3.7
cc_3607 ( N_noxref_15_c_4876_n N_noxref_17_c_5847_n ) capacitor c=0.0205831f \
 //x=55.5 //y=2.08 //x2=58.715 //y2=3.7
cc_3608 ( N_noxref_15_c_4936_p N_noxref_19_c_6213_n ) capacitor c=0.0110241f \
 //x=55.385 //y=3.33 //x2=56.865 //y2=4.07
cc_3609 ( N_noxref_15_c_4921_n N_noxref_19_c_6213_n ) capacitor c=8.88358e-19 \
 //x=53.765 //y=3.33 //x2=56.865 //y2=4.07
cc_3610 ( N_noxref_15_c_4875_n N_noxref_19_c_6213_n ) capacitor c=0.0181936f \
 //x=53.65 //y=3.33 //x2=56.865 //y2=4.07
cc_3611 ( N_noxref_15_c_4876_n N_noxref_19_c_6213_n ) capacitor c=0.0184765f \
 //x=55.5 //y=2.08 //x2=56.865 //y2=4.07
cc_3612 ( N_noxref_15_c_4875_n N_noxref_19_c_6284_n ) capacitor c=0.00117715f \
 //x=53.65 //y=3.33 //x2=53.025 //y2=4.07
cc_3613 ( N_noxref_15_c_4890_n N_noxref_19_c_6286_n ) capacitor c=0.0126603f \
 //x=53.085 //y=5.2 //x2=52.91 //y2=4.535
cc_3614 ( N_noxref_15_c_4875_n N_noxref_19_c_6286_n ) capacitor c=0.0101319f \
 //x=53.65 //y=3.33 //x2=52.91 //y2=4.535
cc_3615 ( N_noxref_15_c_4921_n N_noxref_19_c_6191_n ) capacitor c=0.00329059f \
 //x=53.765 //y=3.33 //x2=52.91 //y2=2.08
cc_3616 ( N_noxref_15_c_4875_n N_noxref_19_c_6191_n ) capacitor c=0.069635f \
 //x=53.65 //y=3.33 //x2=52.91 //y2=2.08
cc_3617 ( N_noxref_15_c_4876_n N_noxref_19_c_6191_n ) capacitor c=8.48165e-19 \
 //x=55.5 //y=2.08 //x2=52.91 //y2=2.08
cc_3618 ( N_noxref_15_M112_noxref_g N_noxref_19_c_6230_n ) capacitor \
 c=0.0169521f //x=55.84 //y=6.02 //x2=56.415 //y2=5.2
cc_3619 ( N_noxref_15_c_4876_n N_noxref_19_c_6234_n ) capacitor c=0.00539951f \
 //x=55.5 //y=2.08 //x2=55.705 //y2=5.2
cc_3620 ( N_noxref_15_M111_noxref_g N_noxref_19_c_6234_n ) capacitor \
 c=0.0177326f //x=55.4 //y=6.02 //x2=55.705 //y2=5.2
cc_3621 ( N_noxref_15_c_4909_n N_noxref_19_c_6234_n ) capacitor c=0.00581252f \
 //x=55.5 //y=4.7 //x2=55.705 //y2=5.2
cc_3622 ( N_noxref_15_c_4875_n N_noxref_19_c_6194_n ) capacitor c=3.49822e-19 \
 //x=53.65 //y=3.33 //x2=56.98 //y2=4.07
cc_3623 ( N_noxref_15_c_4876_n N_noxref_19_c_6194_n ) capacitor c=0.0034228f \
 //x=55.5 //y=2.08 //x2=56.98 //y2=4.07
cc_3624 ( N_noxref_15_c_4890_n N_noxref_19_M109_noxref_g ) capacitor \
 c=0.0166421f //x=53.085 //y=5.2 //x2=52.95 //y2=6.02
cc_3625 ( N_noxref_15_M109_noxref_d N_noxref_19_M109_noxref_g ) capacitor \
 c=0.0173476f //x=53.025 //y=5.02 //x2=52.95 //y2=6.02
cc_3626 ( N_noxref_15_c_4896_n N_noxref_19_M110_noxref_g ) capacitor \
 c=0.018922f //x=53.565 //y=5.2 //x2=53.39 //y2=6.02
cc_3627 ( N_noxref_15_M109_noxref_d N_noxref_19_M110_noxref_g ) capacitor \
 c=0.0179769f //x=53.025 //y=5.02 //x2=53.39 //y2=6.02
cc_3628 ( N_noxref_15_M32_noxref_d N_noxref_19_c_6295_n ) capacitor \
 c=0.00217566f //x=53.02 //y=0.905 //x2=52.945 //y2=0.905
cc_3629 ( N_noxref_15_M32_noxref_d N_noxref_19_c_6298_n ) capacitor \
 c=0.0034598f //x=53.02 //y=0.905 //x2=52.945 //y2=1.25
cc_3630 ( N_noxref_15_M32_noxref_d N_noxref_19_c_6300_n ) capacitor \
 c=0.00669531f //x=53.02 //y=0.905 //x2=52.945 //y2=1.56
cc_3631 ( N_noxref_15_c_4875_n N_noxref_19_c_6332_n ) capacitor c=0.0142673f \
 //x=53.65 //y=3.33 //x2=53.315 //y2=4.79
cc_3632 ( N_noxref_15_c_4985_p N_noxref_19_c_6332_n ) capacitor c=0.00407665f \
 //x=53.17 //y=5.2 //x2=53.315 //y2=4.79
cc_3633 ( N_noxref_15_M32_noxref_d N_noxref_19_c_6334_n ) capacitor \
 c=0.00241102f //x=53.02 //y=0.905 //x2=53.32 //y2=0.75
cc_3634 ( N_noxref_15_c_4874_n N_noxref_19_c_6335_n ) capacitor c=0.00371277f \
 //x=53.565 //y=1.655 //x2=53.32 //y2=1.405
cc_3635 ( N_noxref_15_M32_noxref_d N_noxref_19_c_6335_n ) capacitor \
 c=0.0137169f //x=53.02 //y=0.905 //x2=53.32 //y2=1.405
cc_3636 ( N_noxref_15_M32_noxref_d N_noxref_19_c_6303_n ) capacitor \
 c=0.00132245f //x=53.02 //y=0.905 //x2=53.475 //y2=0.905
cc_3637 ( N_noxref_15_c_4874_n N_noxref_19_c_6304_n ) capacitor c=0.00457401f \
 //x=53.565 //y=1.655 //x2=53.475 //y2=1.25
cc_3638 ( N_noxref_15_M32_noxref_d N_noxref_19_c_6304_n ) capacitor \
 c=0.00566463f //x=53.02 //y=0.905 //x2=53.475 //y2=1.25
cc_3639 ( N_noxref_15_c_4875_n N_noxref_19_c_6305_n ) capacitor c=0.00731987f \
 //x=53.65 //y=3.33 //x2=52.91 //y2=2.08
cc_3640 ( N_noxref_15_c_4875_n N_noxref_19_c_6341_n ) capacitor c=0.00306024f \
 //x=53.65 //y=3.33 //x2=52.91 //y2=1.915
cc_3641 ( N_noxref_15_M32_noxref_d N_noxref_19_c_6341_n ) capacitor \
 c=0.00660593f //x=53.02 //y=0.905 //x2=52.91 //y2=1.915
cc_3642 ( N_noxref_15_c_4890_n N_noxref_19_c_6307_n ) capacitor c=0.00346527f \
 //x=53.085 //y=5.2 //x2=52.94 //y2=4.7
cc_3643 ( N_noxref_15_c_4875_n N_noxref_19_c_6307_n ) capacitor c=0.00517969f \
 //x=53.65 //y=3.33 //x2=52.94 //y2=4.7
cc_3644 ( N_noxref_15_M112_noxref_g N_noxref_19_M111_noxref_d ) capacitor \
 c=0.0173476f //x=55.84 //y=6.02 //x2=55.475 //y2=5.02
cc_3645 ( N_noxref_15_c_4936_p N_noxref_21_c_6911_n ) capacitor c=0.0102155f \
 //x=55.385 //y=3.33 //x2=66.115 //y2=2.22
cc_3646 ( N_noxref_15_c_4921_n N_noxref_21_c_6911_n ) capacitor c=6.82068e-19 \
 //x=53.765 //y=3.33 //x2=66.115 //y2=2.22
cc_3647 ( N_noxref_15_c_5000_p N_noxref_21_c_6911_n ) capacitor c=0.0146822f \
 //x=53.295 //y=1.655 //x2=66.115 //y2=2.22
cc_3648 ( N_noxref_15_c_4875_n N_noxref_21_c_6911_n ) capacitor c=0.0222456f \
 //x=53.65 //y=3.33 //x2=66.115 //y2=2.22
cc_3649 ( N_noxref_15_c_4876_n N_noxref_21_c_6911_n ) capacitor c=0.0208418f \
 //x=55.5 //y=2.08 //x2=66.115 //y2=2.22
cc_3650 ( N_noxref_15_c_4881_n N_noxref_21_c_6911_n ) capacitor c=0.00894156f \
 //x=55.305 //y=1.915 //x2=66.115 //y2=2.22
cc_3651 ( N_noxref_15_c_4936_p N_noxref_23_c_7498_n ) capacitor c=0.173509f \
 //x=55.385 //y=3.33 //x2=70.185 //y2=2.96
cc_3652 ( N_noxref_15_c_4921_n N_noxref_23_c_7498_n ) capacitor c=0.0292689f \
 //x=53.765 //y=3.33 //x2=70.185 //y2=2.96
cc_3653 ( N_noxref_15_c_4875_n N_noxref_23_c_7498_n ) capacitor c=0.0229357f \
 //x=53.65 //y=3.33 //x2=70.185 //y2=2.96
cc_3654 ( N_noxref_15_c_4876_n N_noxref_23_c_7498_n ) capacitor c=0.0228696f \
 //x=55.5 //y=2.08 //x2=70.185 //y2=2.96
cc_3655 ( N_noxref_15_c_5000_p N_noxref_43_c_9119_n ) capacitor c=3.15806e-19 \
 //x=53.295 //y=1.655 //x2=51.755 //y2=1.495
cc_3656 ( N_noxref_15_c_5000_p N_noxref_43_c_9107_n ) capacitor c=0.0203424f \
 //x=53.295 //y=1.655 //x2=52.725 //y2=1.495
cc_3657 ( N_noxref_15_c_4874_n N_noxref_43_c_9108_n ) capacitor c=0.00457164f \
 //x=53.565 //y=1.655 //x2=53.61 //y2=0.53
cc_3658 ( N_noxref_15_M32_noxref_d N_noxref_43_c_9108_n ) capacitor \
 c=0.0115831f //x=53.02 //y=0.905 //x2=53.61 //y2=0.53
cc_3659 ( N_noxref_15_c_4874_n N_noxref_43_M31_noxref_s ) capacitor \
 c=0.013435f //x=53.565 //y=1.655 //x2=51.62 //y2=0.365
cc_3660 ( N_noxref_15_M32_noxref_d N_noxref_43_M31_noxref_s ) capacitor \
 c=0.043966f //x=53.02 //y=0.905 //x2=51.62 //y2=0.365
cc_3661 ( N_noxref_15_c_4874_n N_noxref_44_c_9171_n ) capacitor c=3.22188e-19 \
 //x=53.565 //y=1.655 //x2=55.085 //y2=1.495
cc_3662 ( N_noxref_15_c_4881_n N_noxref_44_c_9171_n ) capacitor c=0.0034165f \
 //x=55.305 //y=1.915 //x2=55.085 //y2=1.495
cc_3663 ( N_noxref_15_c_4876_n N_noxref_44_c_9152_n ) capacitor c=0.011618f \
 //x=55.5 //y=2.08 //x2=55.97 //y2=1.58
cc_3664 ( N_noxref_15_c_4880_n N_noxref_44_c_9152_n ) capacitor c=0.00696403f \
 //x=55.305 //y=1.52 //x2=55.97 //y2=1.58
cc_3665 ( N_noxref_15_c_4881_n N_noxref_44_c_9152_n ) capacitor c=0.0174694f \
 //x=55.305 //y=1.915 //x2=55.97 //y2=1.58
cc_3666 ( N_noxref_15_c_4883_n N_noxref_44_c_9152_n ) capacitor c=0.00776811f \
 //x=55.68 //y=1.365 //x2=55.97 //y2=1.58
cc_3667 ( N_noxref_15_c_4886_n N_noxref_44_c_9152_n ) capacitor c=0.00339872f \
 //x=55.835 //y=1.21 //x2=55.97 //y2=1.58
cc_3668 ( N_noxref_15_c_4881_n N_noxref_44_c_9159_n ) capacitor c=6.71402e-19 \
 //x=55.305 //y=1.915 //x2=56.055 //y2=1.495
cc_3669 ( N_noxref_15_c_4877_n N_noxref_44_M33_noxref_s ) capacitor \
 c=0.0326577f //x=55.305 //y=0.865 //x2=54.95 //y2=0.365
cc_3670 ( N_noxref_15_c_4880_n N_noxref_44_M33_noxref_s ) capacitor \
 c=3.48408e-19 //x=55.305 //y=1.52 //x2=54.95 //y2=0.365
cc_3671 ( N_noxref_15_c_4884_n N_noxref_44_M33_noxref_s ) capacitor \
 c=0.0120759f //x=55.835 //y=0.865 //x2=54.95 //y2=0.365
cc_3672 ( N_CLK_c_5112_n N_noxref_17_c_5873_n ) capacitor c=0.00940379f \
 //x=56.125 //y=4.44 //x2=48.725 //y2=3.7
cc_3673 ( N_CLK_c_5112_n N_noxref_17_c_5874_n ) capacitor c=7.95009e-19 \
 //x=56.125 //y=4.44 //x2=47.105 //y2=3.7
cc_3674 ( N_CLK_c_5112_n N_noxref_17_c_5847_n ) capacitor c=0.0492712f \
 //x=56.125 //y=4.44 //x2=58.715 //y2=3.7
cc_3675 ( N_CLK_c_5032_n N_noxref_17_c_5847_n ) capacitor c=0.0193001f \
 //x=56.24 //y=2.08 //x2=58.715 //y2=3.7
cc_3676 ( N_CLK_c_5112_n N_noxref_17_c_5848_n ) capacitor c=6.59192e-19 \
 //x=56.125 //y=4.44 //x2=48.955 //y2=3.7
cc_3677 ( N_CLK_c_5130_n N_noxref_17_c_5801_n ) capacitor c=0.00241768f \
 //x=45.255 //y=4.44 //x2=45.245 //y2=5.155
cc_3678 ( N_CLK_c_5031_n N_noxref_17_c_5801_n ) capacitor c=0.0143918f \
 //x=45.14 //y=2.08 //x2=45.245 //y2=5.155
cc_3679 ( N_CLK_M99_noxref_g N_noxref_17_c_5801_n ) capacitor c=0.016514f \
 //x=45.11 //y=6.02 //x2=45.245 //y2=5.155
cc_3680 ( N_CLK_c_5536_n N_noxref_17_c_5801_n ) capacitor c=0.00322046f \
 //x=45.14 //y=4.7 //x2=45.245 //y2=5.155
cc_3681 ( N_CLK_c_5092_n N_noxref_17_c_5805_n ) capacitor c=0.0219114f \
 //x=45.025 //y=4.44 //x2=44.535 //y2=5.155
cc_3682 ( N_CLK_M100_noxref_g N_noxref_17_c_5807_n ) capacitor c=0.01736f \
 //x=45.55 //y=6.02 //x2=46.125 //y2=5.155
cc_3683 ( N_CLK_c_5112_n N_noxref_17_c_5811_n ) capacitor c=0.0183122f \
 //x=56.125 //y=4.44 //x2=46.905 //y2=5.155
cc_3684 ( N_CLK_c_5112_n N_noxref_17_c_5815_n ) capacitor c=0.0210274f \
 //x=56.125 //y=4.44 //x2=46.99 //y2=3.7
cc_3685 ( N_CLK_c_5031_n N_noxref_17_c_5815_n ) capacitor c=0.00264025f \
 //x=45.14 //y=2.08 //x2=46.99 //y2=3.7
cc_3686 ( N_CLK_c_5112_n N_noxref_17_c_5778_n ) capacitor c=0.0198304f \
 //x=56.125 //y=4.44 //x2=48.84 //y2=2.08
cc_3687 ( N_CLK_c_5032_n N_noxref_17_c_5779_n ) capacitor c=8.90899e-19 \
 //x=56.24 //y=2.08 //x2=58.83 //y2=2.08
cc_3688 ( N_CLK_c_5112_n N_noxref_17_c_5934_n ) capacitor c=0.0311227f \
 //x=56.125 //y=4.44 //x2=45.33 //y2=5.155
cc_3689 ( N_CLK_c_5535_n N_noxref_17_c_5934_n ) capacitor c=0.00426767f \
 //x=45.475 //y=4.79 //x2=45.33 //y2=5.155
cc_3690 ( N_CLK_c_5112_n N_noxref_17_c_5830_n ) capacitor c=0.0107057f \
 //x=56.125 //y=4.44 //x2=48.84 //y2=4.7
cc_3691 ( N_CLK_M99_noxref_g N_noxref_17_M99_noxref_d ) capacitor c=0.0180032f \
 //x=45.11 //y=6.02 //x2=45.185 //y2=5.02
cc_3692 ( N_CLK_M100_noxref_g N_noxref_17_M99_noxref_d ) capacitor \
 c=0.0180032f //x=45.55 //y=6.02 //x2=45.185 //y2=5.02
cc_3693 ( N_CLK_c_5112_n N_noxref_18_c_6054_n ) capacitor c=0.0035313f \
 //x=56.125 //y=4.44 //x2=60.425 //y2=4.44
cc_3694 ( N_CLK_c_5092_n N_noxref_19_c_6210_n ) capacitor c=0.076217f \
 //x=45.025 //y=4.44 //x2=52.795 //y2=4.07
cc_3695 ( N_CLK_c_5112_n N_noxref_19_c_6210_n ) capacitor c=0.656956f \
 //x=56.125 //y=4.44 //x2=52.795 //y2=4.07
cc_3696 ( N_CLK_c_5130_n N_noxref_19_c_6210_n ) capacitor c=0.026534f \
 //x=45.255 //y=4.44 //x2=52.795 //y2=4.07
cc_3697 ( N_CLK_c_5031_n N_noxref_19_c_6210_n ) capacitor c=0.0247116f \
 //x=45.14 //y=2.08 //x2=52.795 //y2=4.07
cc_3698 ( N_CLK_c_5092_n N_noxref_19_c_6212_n ) capacitor c=0.0290178f \
 //x=45.025 //y=4.44 //x2=44.145 //y2=4.07
cc_3699 ( N_CLK_c_5031_n N_noxref_19_c_6212_n ) capacitor c=0.00128547f \
 //x=45.14 //y=2.08 //x2=44.145 //y2=4.07
cc_3700 ( N_CLK_c_5112_n N_noxref_19_c_6213_n ) capacitor c=0.300301f \
 //x=56.125 //y=4.44 //x2=56.865 //y2=4.07
cc_3701 ( N_CLK_c_5032_n N_noxref_19_c_6213_n ) capacitor c=0.0187718f \
 //x=56.24 //y=2.08 //x2=56.865 //y2=4.07
cc_3702 ( N_CLK_c_5596_p N_noxref_19_c_6213_n ) capacitor c=0.00756255f \
 //x=56.645 //y=4.79 //x2=56.865 //y2=4.07
cc_3703 ( N_CLK_c_5564_n N_noxref_19_c_6213_n ) capacitor c=4.6185e-19 \
 //x=56.27 //y=4.7 //x2=56.865 //y2=4.07
cc_3704 ( N_CLK_c_5112_n N_noxref_19_c_6284_n ) capacitor c=0.0263375f \
 //x=56.125 //y=4.44 //x2=53.025 //y2=4.07
cc_3705 ( N_CLK_c_5032_n N_noxref_19_c_6222_n ) capacitor c=0.00117715f \
 //x=56.24 //y=2.08 //x2=57.095 //y2=4.07
cc_3706 ( N_CLK_c_5092_n N_noxref_19_c_6190_n ) capacitor c=0.0227055f \
 //x=45.025 //y=4.44 //x2=44.03 //y2=2.08
cc_3707 ( N_CLK_c_5130_n N_noxref_19_c_6190_n ) capacitor c=0.00153281f \
 //x=45.255 //y=4.44 //x2=44.03 //y2=2.08
cc_3708 ( N_CLK_c_5031_n N_noxref_19_c_6190_n ) capacitor c=0.0456878f \
 //x=45.14 //y=2.08 //x2=44.03 //y2=2.08
cc_3709 ( N_CLK_c_5532_n N_noxref_19_c_6190_n ) capacitor c=0.00203769f \
 //x=45.23 //y=1.915 //x2=44.03 //y2=2.08
cc_3710 ( N_CLK_c_5536_n N_noxref_19_c_6190_n ) capacitor c=0.00183762f \
 //x=45.14 //y=4.7 //x2=44.03 //y2=2.08
cc_3711 ( N_CLK_c_5112_n N_noxref_19_c_6286_n ) capacitor c=0.0016972f \
 //x=56.125 //y=4.44 //x2=52.91 //y2=4.535
cc_3712 ( N_CLK_c_5112_n N_noxref_19_c_6191_n ) capacitor c=0.0207534f \
 //x=56.125 //y=4.44 //x2=52.91 //y2=2.08
cc_3713 ( N_CLK_c_5112_n N_noxref_19_c_6230_n ) capacitor c=0.00325337f \
 //x=56.125 //y=4.44 //x2=56.415 //y2=5.2
cc_3714 ( N_CLK_c_5543_n N_noxref_19_c_6230_n ) capacitor c=0.0126974f \
 //x=56.24 //y=4.535 //x2=56.415 //y2=5.2
cc_3715 ( N_CLK_c_5032_n N_noxref_19_c_6230_n ) capacitor c=3.74769e-19 \
 //x=56.24 //y=2.08 //x2=56.415 //y2=5.2
cc_3716 ( N_CLK_M113_noxref_g N_noxref_19_c_6230_n ) capacitor c=0.0166421f \
 //x=56.28 //y=6.02 //x2=56.415 //y2=5.2
cc_3717 ( N_CLK_c_5564_n N_noxref_19_c_6230_n ) capacitor c=0.00346519f \
 //x=56.27 //y=4.7 //x2=56.415 //y2=5.2
cc_3718 ( N_CLK_c_5112_n N_noxref_19_c_6234_n ) capacitor c=0.0172877f \
 //x=56.125 //y=4.44 //x2=55.705 //y2=5.2
cc_3719 ( N_CLK_M114_noxref_g N_noxref_19_c_6236_n ) capacitor c=0.0199348f \
 //x=56.72 //y=6.02 //x2=56.895 //y2=5.2
cc_3720 ( N_CLK_c_5614_p N_noxref_19_c_6193_n ) capacitor c=0.00371277f \
 //x=56.65 //y=1.405 //x2=56.895 //y2=1.655
cc_3721 ( N_CLK_c_5561_n N_noxref_19_c_6193_n ) capacitor c=0.00457401f \
 //x=56.805 //y=1.25 //x2=56.895 //y2=1.655
cc_3722 ( N_CLK_c_5112_n N_noxref_19_c_6194_n ) capacitor c=0.0047845f \
 //x=56.125 //y=4.44 //x2=56.98 //y2=4.07
cc_3723 ( N_CLK_c_5543_n N_noxref_19_c_6194_n ) capacitor c=0.00923416f \
 //x=56.24 //y=4.535 //x2=56.98 //y2=4.07
cc_3724 ( N_CLK_c_5032_n N_noxref_19_c_6194_n ) capacitor c=0.0711489f \
 //x=56.24 //y=2.08 //x2=56.98 //y2=4.07
cc_3725 ( N_CLK_c_5596_p N_noxref_19_c_6194_n ) capacitor c=0.0142673f \
 //x=56.645 //y=4.79 //x2=56.98 //y2=4.07
cc_3726 ( N_CLK_c_5562_n N_noxref_19_c_6194_n ) capacitor c=0.00731987f \
 //x=56.24 //y=2.08 //x2=56.98 //y2=4.07
cc_3727 ( N_CLK_c_5621_p N_noxref_19_c_6194_n ) capacitor c=0.00306024f \
 //x=56.24 //y=1.915 //x2=56.98 //y2=4.07
cc_3728 ( N_CLK_c_5564_n N_noxref_19_c_6194_n ) capacitor c=0.00518077f \
 //x=56.27 //y=4.7 //x2=56.98 //y2=4.07
cc_3729 ( N_CLK_c_5596_p N_noxref_19_c_6381_n ) capacitor c=0.00408717f \
 //x=56.645 //y=4.79 //x2=56.5 //y2=5.2
cc_3730 ( N_CLK_M99_noxref_g N_noxref_19_M97_noxref_g ) capacitor c=0.0105869f \
 //x=45.11 //y=6.02 //x2=44.23 //y2=6.02
cc_3731 ( N_CLK_M99_noxref_g N_noxref_19_M98_noxref_g ) capacitor c=0.10632f \
 //x=45.11 //y=6.02 //x2=44.67 //y2=6.02
cc_3732 ( N_CLK_M100_noxref_g N_noxref_19_M98_noxref_g ) capacitor \
 c=0.0101598f //x=45.55 //y=6.02 //x2=44.67 //y2=6.02
cc_3733 ( N_CLK_c_5627_p N_noxref_19_c_6197_n ) capacitor c=5.72482e-19 \
 //x=44.705 //y=0.91 //x2=43.73 //y2=0.875
cc_3734 ( N_CLK_c_5627_p N_noxref_19_c_6199_n ) capacitor c=0.00149976f \
 //x=44.705 //y=0.91 //x2=43.73 //y2=1.22
cc_3735 ( N_CLK_c_5629_p N_noxref_19_c_6200_n ) capacitor c=0.00111227f \
 //x=44.705 //y=1.22 //x2=43.73 //y2=1.53
cc_3736 ( N_CLK_c_5031_n N_noxref_19_c_6201_n ) capacitor c=0.00210802f \
 //x=45.14 //y=2.08 //x2=43.73 //y2=1.915
cc_3737 ( N_CLK_c_5532_n N_noxref_19_c_6201_n ) capacitor c=0.00834532f \
 //x=45.23 //y=1.915 //x2=43.73 //y2=1.915
cc_3738 ( N_CLK_c_5627_p N_noxref_19_c_6204_n ) capacitor c=0.0160123f \
 //x=44.705 //y=0.91 //x2=44.26 //y2=0.875
cc_3739 ( N_CLK_c_5529_n N_noxref_19_c_6204_n ) capacitor c=0.00103227f \
 //x=45.23 //y=0.91 //x2=44.26 //y2=0.875
cc_3740 ( N_CLK_c_5629_p N_noxref_19_c_6206_n ) capacitor c=0.0124075f \
 //x=44.705 //y=1.22 //x2=44.26 //y2=1.22
cc_3741 ( N_CLK_c_5530_n N_noxref_19_c_6206_n ) capacitor c=0.0010154f \
 //x=45.23 //y=1.22 //x2=44.26 //y2=1.22
cc_3742 ( N_CLK_c_5531_n N_noxref_19_c_6206_n ) capacitor c=9.23422e-19 \
 //x=45.23 //y=1.45 //x2=44.26 //y2=1.22
cc_3743 ( N_CLK_c_5031_n N_noxref_19_c_6395_n ) capacitor c=0.00147352f \
 //x=45.14 //y=2.08 //x2=44.595 //y2=4.79
cc_3744 ( N_CLK_c_5536_n N_noxref_19_c_6395_n ) capacitor c=0.0168581f \
 //x=45.14 //y=4.7 //x2=44.595 //y2=4.79
cc_3745 ( N_CLK_c_5092_n N_noxref_19_c_6258_n ) capacitor c=0.0166959f \
 //x=45.025 //y=4.44 //x2=44.305 //y2=4.79
cc_3746 ( N_CLK_c_5031_n N_noxref_19_c_6258_n ) capacitor c=0.00141297f \
 //x=45.14 //y=2.08 //x2=44.305 //y2=4.79
cc_3747 ( N_CLK_c_5536_n N_noxref_19_c_6258_n ) capacitor c=0.00484466f \
 //x=45.14 //y=4.7 //x2=44.305 //y2=4.79
cc_3748 ( N_CLK_c_5112_n N_noxref_19_c_6332_n ) capacitor c=0.00960248f \
 //x=56.125 //y=4.44 //x2=53.315 //y2=4.79
cc_3749 ( N_CLK_c_5112_n N_noxref_19_c_6307_n ) capacitor c=0.00203982f \
 //x=56.125 //y=4.44 //x2=52.94 //y2=4.7
cc_3750 ( N_CLK_c_5552_n N_noxref_19_M34_noxref_d ) capacitor c=0.00217566f \
 //x=56.275 //y=0.905 //x2=56.35 //y2=0.905
cc_3751 ( N_CLK_c_5555_n N_noxref_19_M34_noxref_d ) capacitor c=0.0034598f \
 //x=56.275 //y=1.25 //x2=56.35 //y2=0.905
cc_3752 ( N_CLK_c_5557_n N_noxref_19_M34_noxref_d ) capacitor c=0.00669531f \
 //x=56.275 //y=1.56 //x2=56.35 //y2=0.905
cc_3753 ( N_CLK_c_5647_p N_noxref_19_M34_noxref_d ) capacitor c=0.00241102f \
 //x=56.65 //y=0.75 //x2=56.35 //y2=0.905
cc_3754 ( N_CLK_c_5614_p N_noxref_19_M34_noxref_d ) capacitor c=0.0137169f \
 //x=56.65 //y=1.405 //x2=56.35 //y2=0.905
cc_3755 ( N_CLK_c_5560_n N_noxref_19_M34_noxref_d ) capacitor c=0.00132245f \
 //x=56.805 //y=0.905 //x2=56.35 //y2=0.905
cc_3756 ( N_CLK_c_5561_n N_noxref_19_M34_noxref_d ) capacitor c=0.00566463f \
 //x=56.805 //y=1.25 //x2=56.35 //y2=0.905
cc_3757 ( N_CLK_c_5621_p N_noxref_19_M34_noxref_d ) capacitor c=0.00660593f \
 //x=56.24 //y=1.915 //x2=56.35 //y2=0.905
cc_3758 ( N_CLK_M113_noxref_g N_noxref_19_M113_noxref_d ) capacitor \
 c=0.0173476f //x=56.28 //y=6.02 //x2=56.355 //y2=5.02
cc_3759 ( N_CLK_M114_noxref_g N_noxref_19_M113_noxref_d ) capacitor \
 c=0.0179769f //x=56.72 //y=6.02 //x2=56.355 //y2=5.02
cc_3760 ( N_CLK_c_5031_n N_noxref_21_c_6911_n ) capacitor c=0.0193884f \
 //x=45.14 //y=2.08 //x2=66.115 //y2=2.22
cc_3761 ( N_CLK_c_5032_n N_noxref_21_c_6911_n ) capacitor c=0.0201924f \
 //x=56.24 //y=2.08 //x2=66.115 //y2=2.22
cc_3762 ( N_CLK_c_5532_n N_noxref_21_c_6911_n ) capacitor c=0.00583058f \
 //x=45.23 //y=1.915 //x2=66.115 //y2=2.22
cc_3763 ( N_CLK_c_5614_p N_noxref_21_c_6911_n ) capacitor c=3.11115e-19 \
 //x=56.65 //y=1.405 //x2=66.115 //y2=2.22
cc_3764 ( N_CLK_c_5562_n N_noxref_21_c_6911_n ) capacitor c=0.00568402f \
 //x=56.24 //y=2.08 //x2=66.115 //y2=2.22
cc_3765 ( N_CLK_c_5092_n N_noxref_21_c_7001_n ) capacitor c=0.0016972f \
 //x=45.025 //y=4.44 //x2=38.11 //y2=4.535
cc_3766 ( N_CLK_c_5092_n N_noxref_21_c_6939_n ) capacitor c=0.0189188f \
 //x=45.025 //y=4.44 //x2=38.11 //y2=2.08
cc_3767 ( N_CLK_c_5092_n N_noxref_21_c_6959_n ) capacitor c=0.0185677f \
 //x=45.025 //y=4.44 //x2=41.615 //y2=5.2
cc_3768 ( N_CLK_c_5092_n N_noxref_21_c_6963_n ) capacitor c=0.018142f \
 //x=45.025 //y=4.44 //x2=40.905 //y2=5.2
cc_3769 ( N_CLK_c_5092_n N_noxref_21_c_6942_n ) capacitor c=0.0256789f \
 //x=45.025 //y=4.44 //x2=42.18 //y2=2.22
cc_3770 ( N_CLK_c_5031_n N_noxref_21_c_6942_n ) capacitor c=5.45205e-19 \
 //x=45.14 //y=2.08 //x2=42.18 //y2=2.22
cc_3771 ( N_CLK_c_5092_n N_noxref_21_c_7046_n ) capacitor c=0.00960248f \
 //x=45.025 //y=4.44 //x2=38.515 //y2=4.79
cc_3772 ( N_CLK_c_5092_n N_noxref_21_c_7021_n ) capacitor c=0.00203982f \
 //x=45.025 //y=4.44 //x2=38.14 //y2=4.7
cc_3773 ( N_CLK_c_5079_n N_noxref_23_c_7497_n ) capacitor c=0.0170511f \
 //x=23.795 //y=4.44 //x2=20.605 //y2=2.96
cc_3774 ( N_CLK_c_5053_n N_noxref_23_c_7578_n ) capacitor c=4.06095e-19 \
 //x=16.745 //y=4.442 //x2=16.765 //y2=2.96
cc_3775 ( N_CLK_c_5061_n N_noxref_23_c_7498_n ) capacitor c=0.00594004f \
 //x=34.665 //y=4.44 //x2=70.185 //y2=2.96
cc_3776 ( N_CLK_c_5079_n N_noxref_23_c_7498_n ) capacitor c=0.042751f \
 //x=23.795 //y=4.44 //x2=70.185 //y2=2.96
cc_3777 ( N_CLK_c_5092_n N_noxref_23_c_7498_n ) capacitor c=0.0662424f \
 //x=45.025 //y=4.44 //x2=70.185 //y2=2.96
cc_3778 ( N_CLK_c_5112_n N_noxref_23_c_7498_n ) capacitor c=0.00594004f \
 //x=56.125 //y=4.44 //x2=70.185 //y2=2.96
cc_3779 ( N_CLK_c_5130_n N_noxref_23_c_7498_n ) capacitor c=4.4954e-19 \
 //x=45.255 //y=4.44 //x2=70.185 //y2=2.96
cc_3780 ( N_CLK_c_5028_n N_noxref_23_c_7498_n ) capacitor c=0.0228892f \
 //x=23.68 //y=2.08 //x2=70.185 //y2=2.96
cc_3781 ( N_CLK_c_5029_n N_noxref_23_c_7498_n ) capacitor c=0.019291f \
 //x=34.78 //y=2.08 //x2=70.185 //y2=2.96
cc_3782 ( N_CLK_c_5031_n N_noxref_23_c_7498_n ) capacitor c=0.0228892f \
 //x=45.14 //y=2.08 //x2=70.185 //y2=2.96
cc_3783 ( N_CLK_c_5032_n N_noxref_23_c_7498_n ) capacitor c=0.0215847f \
 //x=56.24 //y=2.08 //x2=70.185 //y2=2.96
cc_3784 ( N_CLK_c_5079_n N_noxref_23_c_7641_n ) capacitor c=0.00454388f \
 //x=23.795 //y=4.44 //x2=20.835 //y2=2.96
cc_3785 ( N_CLK_c_5053_n N_noxref_23_c_7579_n ) capacitor c=5.33303e-19 \
 //x=16.745 //y=4.442 //x2=16.65 //y2=4.535
cc_3786 ( N_CLK_c_5079_n N_noxref_23_c_7579_n ) capacitor c=0.00113146f \
 //x=23.795 //y=4.44 //x2=16.65 //y2=4.535
cc_3787 ( N_CLK_c_5053_n N_noxref_23_c_7515_n ) capacitor c=0.0179078f \
 //x=16.745 //y=4.442 //x2=16.65 //y2=2.08
cc_3788 ( N_CLK_c_5079_n N_noxref_23_c_7515_n ) capacitor c=6.30528e-19 \
 //x=23.795 //y=4.44 //x2=16.65 //y2=2.08
cc_3789 ( N_CLK_c_5079_n N_noxref_23_c_7540_n ) capacitor c=0.0185677f \
 //x=23.795 //y=4.44 //x2=20.155 //y2=5.2
cc_3790 ( N_CLK_c_5079_n N_noxref_23_c_7544_n ) capacitor c=0.018142f \
 //x=23.795 //y=4.44 //x2=19.445 //y2=5.2
cc_3791 ( N_CLK_c_5079_n N_noxref_23_c_7518_n ) capacitor c=0.0257082f \
 //x=23.795 //y=4.44 //x2=20.72 //y2=2.96
cc_3792 ( N_CLK_c_5028_n N_noxref_23_c_7518_n ) capacitor c=5.89489e-19 \
 //x=23.68 //y=2.08 //x2=20.72 //y2=2.96
cc_3793 ( N_CLK_c_5079_n N_noxref_23_c_7624_n ) capacitor c=0.00960248f \
 //x=23.795 //y=4.44 //x2=17.055 //y2=4.79
cc_3794 ( N_CLK_c_5053_n N_noxref_23_c_7599_n ) capacitor c=5.57952e-19 \
 //x=16.745 //y=4.442 //x2=16.68 //y2=4.7
cc_3795 ( N_CLK_c_5079_n N_noxref_23_c_7599_n ) capacitor c=0.00146858f \
 //x=23.795 //y=4.44 //x2=16.68 //y2=4.7
cc_3796 ( N_CLK_c_5300_n N_noxref_26_c_8221_n ) capacitor c=0.0167228f \
 //x=1.785 //y=0.91 //x2=2.445 //y2=0.54
cc_3797 ( N_CLK_c_5187_n N_noxref_26_c_8221_n ) capacitor c=0.00534519f \
 //x=2.31 //y=0.91 //x2=2.445 //y2=0.54
cc_3798 ( N_CLK_c_5025_n N_noxref_26_c_8239_n ) capacitor c=0.012357f //x=2.22 \
 //y=2.08 //x2=2.445 //y2=1.59
cc_3799 ( N_CLK_c_5303_n N_noxref_26_c_8239_n ) capacitor c=0.0153476f \
 //x=1.785 //y=1.22 //x2=2.445 //y2=1.59
cc_3800 ( N_CLK_c_5190_n N_noxref_26_c_8239_n ) capacitor c=0.0230663f \
 //x=2.31 //y=1.915 //x2=2.445 //y2=1.59
cc_3801 ( N_CLK_c_5300_n N_noxref_26_M0_noxref_s ) capacitor c=0.00798959f \
 //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_3802 ( N_CLK_c_5189_n N_noxref_26_M0_noxref_s ) capacitor c=0.00212176f \
 //x=2.31 //y=1.45 //x2=0.455 //y2=0.375
cc_3803 ( N_CLK_c_5190_n N_noxref_26_M0_noxref_s ) capacitor c=0.00298115f \
 //x=2.31 //y=1.915 //x2=0.455 //y2=0.375
cc_3804 ( N_CLK_c_5698_p N_noxref_27_c_8261_n ) capacitor c=2.14837e-19 \
 //x=2.155 //y=0.755 //x2=3.015 //y2=0.995
cc_3805 ( N_CLK_c_5187_n N_noxref_27_c_8261_n ) capacitor c=0.00123426f \
 //x=2.31 //y=0.91 //x2=3.015 //y2=0.995
cc_3806 ( N_CLK_c_5188_n N_noxref_27_c_8261_n ) capacitor c=0.0129288f \
 //x=2.31 //y=1.22 //x2=3.015 //y2=0.995
cc_3807 ( N_CLK_c_5189_n N_noxref_27_c_8261_n ) capacitor c=0.00142359f \
 //x=2.31 //y=1.45 //x2=3.015 //y2=0.995
cc_3808 ( N_CLK_c_5300_n N_noxref_27_M1_noxref_d ) capacitor c=0.00223875f \
 //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_3809 ( N_CLK_c_5303_n N_noxref_27_M1_noxref_d ) capacitor c=0.00262485f \
 //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_3810 ( N_CLK_c_5698_p N_noxref_27_M1_noxref_d ) capacitor c=0.00220746f \
 //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_3811 ( N_CLK_c_5705_p N_noxref_27_M1_noxref_d ) capacitor c=0.00194798f \
 //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_3812 ( N_CLK_c_5187_n N_noxref_27_M1_noxref_d ) capacitor c=0.00198465f \
 //x=2.31 //y=0.91 //x2=1.86 //y2=0.91
cc_3813 ( N_CLK_c_5188_n N_noxref_27_M1_noxref_d ) capacitor c=0.00128384f \
 //x=2.31 //y=1.22 //x2=1.86 //y2=0.91
cc_3814 ( N_CLK_c_5187_n N_noxref_27_M2_noxref_s ) capacitor c=7.21316e-19 \
 //x=2.31 //y=0.91 //x2=2.965 //y2=0.375
cc_3815 ( N_CLK_c_5188_n N_noxref_27_M2_noxref_s ) capacitor c=0.00348171f \
 //x=2.31 //y=1.22 //x2=2.965 //y2=0.375
cc_3816 ( N_CLK_c_5217_n N_noxref_30_c_8427_n ) capacitor c=0.00623646f \
 //x=13.355 //y=1.56 //x2=13.135 //y2=1.495
cc_3817 ( N_CLK_c_5222_n N_noxref_30_c_8427_n ) capacitor c=0.00174019f \
 //x=13.32 //y=2.08 //x2=13.135 //y2=1.495
cc_3818 ( N_CLK_c_5026_n N_noxref_30_c_8428_n ) capacitor c=0.00158203f \
 //x=13.32 //y=2.08 //x2=14.02 //y2=0.53
cc_3819 ( N_CLK_c_5212_n N_noxref_30_c_8428_n ) capacitor c=0.0188655f \
 //x=13.355 //y=0.905 //x2=14.02 //y2=0.53
cc_3820 ( N_CLK_c_5220_n N_noxref_30_c_8428_n ) capacitor c=0.00656458f \
 //x=13.885 //y=0.905 //x2=14.02 //y2=0.53
cc_3821 ( N_CLK_c_5222_n N_noxref_30_c_8428_n ) capacitor c=2.1838e-19 \
 //x=13.32 //y=2.08 //x2=14.02 //y2=0.53
cc_3822 ( N_CLK_c_5212_n N_noxref_30_M7_noxref_s ) capacitor c=0.00623646f \
 //x=13.355 //y=0.905 //x2=12.03 //y2=0.365
cc_3823 ( N_CLK_c_5220_n N_noxref_30_M7_noxref_s ) capacitor c=0.0143002f \
 //x=13.885 //y=0.905 //x2=12.03 //y2=0.365
cc_3824 ( N_CLK_c_5221_n N_noxref_30_M7_noxref_s ) capacitor c=0.00290153f \
 //x=13.885 //y=1.25 //x2=12.03 //y2=0.365
cc_3825 ( N_CLK_c_5461_n N_noxref_33_c_8583_n ) capacitor c=0.0167228f \
 //x=23.245 //y=0.91 //x2=23.905 //y2=0.54
cc_3826 ( N_CLK_c_5347_n N_noxref_33_c_8583_n ) capacitor c=0.00534519f \
 //x=23.77 //y=0.91 //x2=23.905 //y2=0.54
cc_3827 ( N_CLK_c_5028_n N_noxref_33_c_8605_n ) capacitor c=0.012334f \
 //x=23.68 //y=2.08 //x2=23.905 //y2=1.59
cc_3828 ( N_CLK_c_5464_n N_noxref_33_c_8605_n ) capacitor c=0.0153476f \
 //x=23.245 //y=1.22 //x2=23.905 //y2=1.59
cc_3829 ( N_CLK_c_5350_n N_noxref_33_c_8605_n ) capacitor c=0.0219329f \
 //x=23.77 //y=1.915 //x2=23.905 //y2=1.59
cc_3830 ( N_CLK_c_5461_n N_noxref_33_M13_noxref_s ) capacitor c=0.00798959f \
 //x=23.245 //y=0.91 //x2=21.915 //y2=0.375
cc_3831 ( N_CLK_c_5349_n N_noxref_33_M13_noxref_s ) capacitor c=0.00212176f \
 //x=23.77 //y=1.45 //x2=21.915 //y2=0.375
cc_3832 ( N_CLK_c_5350_n N_noxref_33_M13_noxref_s ) capacitor c=0.00298115f \
 //x=23.77 //y=1.915 //x2=21.915 //y2=0.375
cc_3833 ( N_CLK_c_5727_p N_noxref_34_c_8626_n ) capacitor c=2.14837e-19 \
 //x=23.615 //y=0.755 //x2=24.475 //y2=0.995
cc_3834 ( N_CLK_c_5347_n N_noxref_34_c_8626_n ) capacitor c=0.00123426f \
 //x=23.77 //y=0.91 //x2=24.475 //y2=0.995
cc_3835 ( N_CLK_c_5348_n N_noxref_34_c_8626_n ) capacitor c=0.0129288f \
 //x=23.77 //y=1.22 //x2=24.475 //y2=0.995
cc_3836 ( N_CLK_c_5349_n N_noxref_34_c_8626_n ) capacitor c=0.00142359f \
 //x=23.77 //y=1.45 //x2=24.475 //y2=0.995
cc_3837 ( N_CLK_c_5461_n N_noxref_34_M14_noxref_d ) capacitor c=0.00223875f \
 //x=23.245 //y=0.91 //x2=23.32 //y2=0.91
cc_3838 ( N_CLK_c_5464_n N_noxref_34_M14_noxref_d ) capacitor c=0.00262485f \
 //x=23.245 //y=1.22 //x2=23.32 //y2=0.91
cc_3839 ( N_CLK_c_5727_p N_noxref_34_M14_noxref_d ) capacitor c=0.00220746f \
 //x=23.615 //y=0.755 //x2=23.32 //y2=0.91
cc_3840 ( N_CLK_c_5734_p N_noxref_34_M14_noxref_d ) capacitor c=0.00194798f \
 //x=23.615 //y=1.375 //x2=23.32 //y2=0.91
cc_3841 ( N_CLK_c_5347_n N_noxref_34_M14_noxref_d ) capacitor c=0.00198465f \
 //x=23.77 //y=0.91 //x2=23.32 //y2=0.91
cc_3842 ( N_CLK_c_5348_n N_noxref_34_M14_noxref_d ) capacitor c=0.00128384f \
 //x=23.77 //y=1.22 //x2=23.32 //y2=0.91
cc_3843 ( N_CLK_c_5347_n N_noxref_34_M15_noxref_s ) capacitor c=7.21316e-19 \
 //x=23.77 //y=0.91 //x2=24.425 //y2=0.375
cc_3844 ( N_CLK_c_5348_n N_noxref_34_M15_noxref_s ) capacitor c=0.00348171f \
 //x=23.77 //y=1.22 //x2=24.425 //y2=0.375
cc_3845 ( N_CLK_c_5377_n N_noxref_37_c_8792_n ) capacitor c=0.00623646f \
 //x=34.815 //y=1.56 //x2=34.595 //y2=1.495
cc_3846 ( N_CLK_c_5382_n N_noxref_37_c_8792_n ) capacitor c=0.00174019f \
 //x=34.78 //y=2.08 //x2=34.595 //y2=1.495
cc_3847 ( N_CLK_c_5029_n N_noxref_37_c_8793_n ) capacitor c=0.00158203f \
 //x=34.78 //y=2.08 //x2=35.48 //y2=0.53
cc_3848 ( N_CLK_c_5372_n N_noxref_37_c_8793_n ) capacitor c=0.0188655f \
 //x=34.815 //y=0.905 //x2=35.48 //y2=0.53
cc_3849 ( N_CLK_c_5380_n N_noxref_37_c_8793_n ) capacitor c=0.00656458f \
 //x=35.345 //y=0.905 //x2=35.48 //y2=0.53
cc_3850 ( N_CLK_c_5382_n N_noxref_37_c_8793_n ) capacitor c=2.1838e-19 \
 //x=34.78 //y=2.08 //x2=35.48 //y2=0.53
cc_3851 ( N_CLK_c_5372_n N_noxref_37_M20_noxref_s ) capacitor c=0.00623646f \
 //x=34.815 //y=0.905 //x2=33.49 //y2=0.365
cc_3852 ( N_CLK_c_5380_n N_noxref_37_M20_noxref_s ) capacitor c=0.0143002f \
 //x=35.345 //y=0.905 //x2=33.49 //y2=0.365
cc_3853 ( N_CLK_c_5381_n N_noxref_37_M20_noxref_s ) capacitor c=0.00290153f \
 //x=35.345 //y=1.25 //x2=33.49 //y2=0.365
cc_3854 ( N_CLK_c_5627_p N_noxref_40_c_8952_n ) capacitor c=0.0167228f \
 //x=44.705 //y=0.91 //x2=45.365 //y2=0.54
cc_3855 ( N_CLK_c_5529_n N_noxref_40_c_8952_n ) capacitor c=0.00534519f \
 //x=45.23 //y=0.91 //x2=45.365 //y2=0.54
cc_3856 ( N_CLK_c_5031_n N_noxref_40_c_8963_n ) capacitor c=0.0117694f \
 //x=45.14 //y=2.08 //x2=45.365 //y2=1.59
cc_3857 ( N_CLK_c_5629_p N_noxref_40_c_8963_n ) capacitor c=0.0157358f \
 //x=44.705 //y=1.22 //x2=45.365 //y2=1.59
cc_3858 ( N_CLK_c_5532_n N_noxref_40_c_8963_n ) capacitor c=0.021347f \
 //x=45.23 //y=1.915 //x2=45.365 //y2=1.59
cc_3859 ( N_CLK_c_5627_p N_noxref_40_M26_noxref_s ) capacitor c=0.00798959f \
 //x=44.705 //y=0.91 //x2=43.375 //y2=0.375
cc_3860 ( N_CLK_c_5531_n N_noxref_40_M26_noxref_s ) capacitor c=0.00212176f \
 //x=45.23 //y=1.45 //x2=43.375 //y2=0.375
cc_3861 ( N_CLK_c_5532_n N_noxref_40_M26_noxref_s ) capacitor c=0.00298115f \
 //x=45.23 //y=1.915 //x2=43.375 //y2=0.375
cc_3862 ( N_CLK_c_5756_p N_noxref_41_c_8995_n ) capacitor c=2.14837e-19 \
 //x=45.075 //y=0.755 //x2=45.935 //y2=0.995
cc_3863 ( N_CLK_c_5529_n N_noxref_41_c_8995_n ) capacitor c=0.00123426f \
 //x=45.23 //y=0.91 //x2=45.935 //y2=0.995
cc_3864 ( N_CLK_c_5530_n N_noxref_41_c_8995_n ) capacitor c=0.0129288f \
 //x=45.23 //y=1.22 //x2=45.935 //y2=0.995
cc_3865 ( N_CLK_c_5531_n N_noxref_41_c_8995_n ) capacitor c=0.00142359f \
 //x=45.23 //y=1.45 //x2=45.935 //y2=0.995
cc_3866 ( N_CLK_c_5627_p N_noxref_41_M27_noxref_d ) capacitor c=0.00223875f \
 //x=44.705 //y=0.91 //x2=44.78 //y2=0.91
cc_3867 ( N_CLK_c_5629_p N_noxref_41_M27_noxref_d ) capacitor c=0.00262485f \
 //x=44.705 //y=1.22 //x2=44.78 //y2=0.91
cc_3868 ( N_CLK_c_5756_p N_noxref_41_M27_noxref_d ) capacitor c=0.00220746f \
 //x=45.075 //y=0.755 //x2=44.78 //y2=0.91
cc_3869 ( N_CLK_c_5763_p N_noxref_41_M27_noxref_d ) capacitor c=0.00194798f \
 //x=45.075 //y=1.375 //x2=44.78 //y2=0.91
cc_3870 ( N_CLK_c_5529_n N_noxref_41_M27_noxref_d ) capacitor c=0.00198465f \
 //x=45.23 //y=0.91 //x2=44.78 //y2=0.91
cc_3871 ( N_CLK_c_5530_n N_noxref_41_M27_noxref_d ) capacitor c=0.00128384f \
 //x=45.23 //y=1.22 //x2=44.78 //y2=0.91
cc_3872 ( N_CLK_c_5529_n N_noxref_41_M28_noxref_s ) capacitor c=7.21316e-19 \
 //x=45.23 //y=0.91 //x2=45.885 //y2=0.375
cc_3873 ( N_CLK_c_5530_n N_noxref_41_M28_noxref_s ) capacitor c=0.00348171f \
 //x=45.23 //y=1.22 //x2=45.885 //y2=0.375
cc_3874 ( N_CLK_c_5557_n N_noxref_44_c_9159_n ) capacitor c=0.00623646f \
 //x=56.275 //y=1.56 //x2=56.055 //y2=1.495
cc_3875 ( N_CLK_c_5562_n N_noxref_44_c_9159_n ) capacitor c=0.00173579f \
 //x=56.24 //y=2.08 //x2=56.055 //y2=1.495
cc_3876 ( N_CLK_c_5032_n N_noxref_44_c_9160_n ) capacitor c=0.00156605f \
 //x=56.24 //y=2.08 //x2=56.94 //y2=0.53
cc_3877 ( N_CLK_c_5552_n N_noxref_44_c_9160_n ) capacitor c=0.0188655f \
 //x=56.275 //y=0.905 //x2=56.94 //y2=0.53
cc_3878 ( N_CLK_c_5560_n N_noxref_44_c_9160_n ) capacitor c=0.00656458f \
 //x=56.805 //y=0.905 //x2=56.94 //y2=0.53
cc_3879 ( N_CLK_c_5562_n N_noxref_44_c_9160_n ) capacitor c=2.1838e-19 \
 //x=56.24 //y=2.08 //x2=56.94 //y2=0.53
cc_3880 ( N_CLK_c_5552_n N_noxref_44_M33_noxref_s ) capacitor c=0.00623646f \
 //x=56.275 //y=0.905 //x2=54.95 //y2=0.365
cc_3881 ( N_CLK_c_5560_n N_noxref_44_M33_noxref_s ) capacitor c=0.0143002f \
 //x=56.805 //y=0.905 //x2=54.95 //y2=0.365
cc_3882 ( N_CLK_c_5561_n N_noxref_44_M33_noxref_s ) capacitor c=0.00290153f \
 //x=56.805 //y=1.25 //x2=54.95 //y2=0.365
cc_3883 ( N_noxref_17_M116_noxref_g N_noxref_18_c_6057_n ) capacitor \
 c=0.017965f //x=59.17 //y=6.02 //x2=59.745 //y2=5.2
cc_3884 ( N_noxref_17_c_5779_n N_noxref_18_c_6061_n ) capacitor c=0.00530485f \
 //x=58.83 //y=2.08 //x2=59.035 //y2=5.2
cc_3885 ( N_noxref_17_M115_noxref_g N_noxref_18_c_6061_n ) capacitor \
 c=0.0177326f //x=58.73 //y=6.02 //x2=59.035 //y2=5.2
cc_3886 ( N_noxref_17_c_5831_n N_noxref_18_c_6061_n ) capacitor c=0.00582246f \
 //x=58.83 //y=4.7 //x2=59.035 //y2=5.2
cc_3887 ( N_noxref_17_c_5779_n N_noxref_18_c_6033_n ) capacitor c=0.00323781f \
 //x=58.83 //y=2.08 //x2=60.31 //y2=4.44
cc_3888 ( N_noxref_17_M116_noxref_g N_noxref_18_M115_noxref_d ) capacitor \
 c=0.0173476f //x=59.17 //y=6.02 //x2=58.805 //y2=5.02
cc_3889 ( N_noxref_17_c_5873_n N_noxref_19_c_6210_n ) capacitor c=0.147021f \
 //x=48.725 //y=3.7 //x2=52.795 //y2=4.07
cc_3890 ( N_noxref_17_c_5874_n N_noxref_19_c_6210_n ) capacitor c=0.0294294f \
 //x=47.105 //y=3.7 //x2=52.795 //y2=4.07
cc_3891 ( N_noxref_17_c_5847_n N_noxref_19_c_6210_n ) capacitor c=0.338937f \
 //x=58.715 //y=3.7 //x2=52.795 //y2=4.07
cc_3892 ( N_noxref_17_c_5848_n N_noxref_19_c_6210_n ) capacitor c=0.0264478f \
 //x=48.955 //y=3.7 //x2=52.795 //y2=4.07
cc_3893 ( N_noxref_17_c_5815_n N_noxref_19_c_6210_n ) capacitor c=0.0200328f \
 //x=46.99 //y=3.7 //x2=52.795 //y2=4.07
cc_3894 ( N_noxref_17_c_5778_n N_noxref_19_c_6210_n ) capacitor c=0.0203111f \
 //x=48.84 //y=2.08 //x2=52.795 //y2=4.07
cc_3895 ( N_noxref_17_c_5847_n N_noxref_19_c_6213_n ) capacitor c=0.339146f \
 //x=58.715 //y=3.7 //x2=56.865 //y2=4.07
cc_3896 ( N_noxref_17_c_5847_n N_noxref_19_c_6284_n ) capacitor c=0.0267832f \
 //x=58.715 //y=3.7 //x2=53.025 //y2=4.07
cc_3897 ( N_noxref_17_c_5847_n N_noxref_19_c_6215_n ) capacitor c=0.176049f \
 //x=58.715 //y=3.7 //x2=62.785 //y2=4.07
cc_3898 ( N_noxref_17_c_5779_n N_noxref_19_c_6215_n ) capacitor c=0.0242341f \
 //x=58.83 //y=2.08 //x2=62.785 //y2=4.07
cc_3899 ( N_noxref_17_c_5831_n N_noxref_19_c_6215_n ) capacitor c=0.00703556f \
 //x=58.83 //y=4.7 //x2=62.785 //y2=4.07
cc_3900 ( N_noxref_17_c_5847_n N_noxref_19_c_6222_n ) capacitor c=0.0266833f \
 //x=58.715 //y=3.7 //x2=57.095 //y2=4.07
cc_3901 ( N_noxref_17_c_5779_n N_noxref_19_c_6222_n ) capacitor c=3.50683e-19 \
 //x=58.83 //y=2.08 //x2=57.095 //y2=4.07
cc_3902 ( N_noxref_17_c_5847_n N_noxref_19_c_6191_n ) capacitor c=0.0211371f \
 //x=58.715 //y=3.7 //x2=52.91 //y2=2.08
cc_3903 ( N_noxref_17_c_5847_n N_noxref_19_c_6194_n ) capacitor c=0.0235138f \
 //x=58.715 //y=3.7 //x2=56.98 //y2=4.07
cc_3904 ( N_noxref_17_c_5779_n N_noxref_19_c_6194_n ) capacitor c=0.0129673f \
 //x=58.83 //y=2.08 //x2=56.98 //y2=4.07
cc_3905 ( N_noxref_17_c_5805_n N_noxref_19_M97_noxref_g ) capacitor \
 c=0.0213876f //x=44.535 //y=5.155 //x2=44.23 //y2=6.02
cc_3906 ( N_noxref_17_c_5801_n N_noxref_19_M98_noxref_g ) capacitor \
 c=0.0168349f //x=45.245 //y=5.155 //x2=44.67 //y2=6.02
cc_3907 ( N_noxref_17_M97_noxref_d N_noxref_19_M98_noxref_g ) capacitor \
 c=0.0180032f //x=44.305 //y=5.02 //x2=44.67 //y2=6.02
cc_3908 ( N_noxref_17_c_5805_n N_noxref_19_c_6395_n ) capacitor c=0.00428486f \
 //x=44.535 //y=5.155 //x2=44.595 //y2=4.79
cc_3909 ( N_noxref_17_c_5847_n N_noxref_20_c_6653_n ) capacitor c=0.0244534f \
 //x=58.715 //y=3.7 //x2=59.685 //y2=3.7
cc_3910 ( N_noxref_17_c_5779_n N_noxref_20_c_6653_n ) capacitor c=0.00246068f \
 //x=58.83 //y=2.08 //x2=59.685 //y2=3.7
cc_3911 ( N_noxref_17_c_5779_n N_noxref_20_c_6655_n ) capacitor c=0.00400249f \
 //x=58.83 //y=2.08 //x2=59.57 //y2=4.535
cc_3912 ( N_noxref_17_c_5831_n N_noxref_20_c_6655_n ) capacitor c=0.00417994f \
 //x=58.83 //y=4.7 //x2=59.57 //y2=4.535
cc_3913 ( N_noxref_17_c_5847_n N_noxref_20_c_6560_n ) capacitor c=0.00246068f \
 //x=58.715 //y=3.7 //x2=59.57 //y2=2.08
cc_3914 ( N_noxref_17_c_5779_n N_noxref_20_c_6560_n ) capacitor c=0.0790324f \
 //x=58.83 //y=2.08 //x2=59.57 //y2=2.08
cc_3915 ( N_noxref_17_c_5794_n N_noxref_20_c_6560_n ) capacitor c=0.00284029f \
 //x=58.635 //y=1.915 //x2=59.57 //y2=2.08
cc_3916 ( N_noxref_17_M115_noxref_g N_noxref_20_M117_noxref_g ) capacitor \
 c=0.0104611f //x=58.73 //y=6.02 //x2=59.61 //y2=6.02
cc_3917 ( N_noxref_17_M116_noxref_g N_noxref_20_M117_noxref_g ) capacitor \
 c=0.106811f //x=59.17 //y=6.02 //x2=59.61 //y2=6.02
cc_3918 ( N_noxref_17_M116_noxref_g N_noxref_20_M118_noxref_g ) capacitor \
 c=0.0100341f //x=59.17 //y=6.02 //x2=60.05 //y2=6.02
cc_3919 ( N_noxref_17_c_5790_n N_noxref_20_c_6663_n ) capacitor c=4.86506e-19 \
 //x=58.635 //y=0.865 //x2=59.605 //y2=0.905
cc_3920 ( N_noxref_17_c_5792_n N_noxref_20_c_6663_n ) capacitor c=0.00152104f \
 //x=58.635 //y=1.21 //x2=59.605 //y2=0.905
cc_3921 ( N_noxref_17_c_5797_n N_noxref_20_c_6663_n ) capacitor c=0.0151475f \
 //x=59.165 //y=0.865 //x2=59.605 //y2=0.905
cc_3922 ( N_noxref_17_c_5793_n N_noxref_20_c_6666_n ) capacitor c=0.00109982f \
 //x=58.635 //y=1.52 //x2=59.605 //y2=1.25
cc_3923 ( N_noxref_17_c_5799_n N_noxref_20_c_6666_n ) capacitor c=0.0111064f \
 //x=59.165 //y=1.21 //x2=59.605 //y2=1.25
cc_3924 ( N_noxref_17_c_5793_n N_noxref_20_c_6668_n ) capacitor c=9.57794e-19 \
 //x=58.635 //y=1.52 //x2=59.605 //y2=1.56
cc_3925 ( N_noxref_17_c_5794_n N_noxref_20_c_6668_n ) capacitor c=0.00662747f \
 //x=58.635 //y=1.915 //x2=59.605 //y2=1.56
cc_3926 ( N_noxref_17_c_5799_n N_noxref_20_c_6668_n ) capacitor c=0.00862358f \
 //x=59.165 //y=1.21 //x2=59.605 //y2=1.56
cc_3927 ( N_noxref_17_c_5797_n N_noxref_20_c_6671_n ) capacitor c=0.00124821f \
 //x=59.165 //y=0.865 //x2=60.135 //y2=0.905
cc_3928 ( N_noxref_17_c_5799_n N_noxref_20_c_6672_n ) capacitor c=0.00200715f \
 //x=59.165 //y=1.21 //x2=60.135 //y2=1.25
cc_3929 ( N_noxref_17_c_5779_n N_noxref_20_c_6673_n ) capacitor c=0.00282278f \
 //x=58.83 //y=2.08 //x2=59.57 //y2=2.08
cc_3930 ( N_noxref_17_c_5794_n N_noxref_20_c_6673_n ) capacitor c=0.0172771f \
 //x=58.635 //y=1.915 //x2=59.57 //y2=2.08
cc_3931 ( N_noxref_17_c_5779_n N_noxref_20_c_6675_n ) capacitor c=0.00344981f \
 //x=58.83 //y=2.08 //x2=59.6 //y2=4.7
cc_3932 ( N_noxref_17_c_5831_n N_noxref_20_c_6675_n ) capacitor c=0.0293367f \
 //x=58.83 //y=4.7 //x2=59.6 //y2=4.7
cc_3933 ( N_noxref_17_c_5847_n N_noxref_21_c_6911_n ) capacitor c=0.0151374f \
 //x=58.715 //y=3.7 //x2=66.115 //y2=2.22
cc_3934 ( N_noxref_17_c_5990_p N_noxref_21_c_6911_n ) capacitor c=0.016327f \
 //x=46.59 //y=1.665 //x2=66.115 //y2=2.22
cc_3935 ( N_noxref_17_c_5815_n N_noxref_21_c_6911_n ) capacitor c=0.0197307f \
 //x=46.99 //y=3.7 //x2=66.115 //y2=2.22
cc_3936 ( N_noxref_17_c_5778_n N_noxref_21_c_6911_n ) capacitor c=0.0185012f \
 //x=48.84 //y=2.08 //x2=66.115 //y2=2.22
cc_3937 ( N_noxref_17_c_5779_n N_noxref_21_c_6911_n ) capacitor c=0.0208418f \
 //x=58.83 //y=2.08 //x2=66.115 //y2=2.22
cc_3938 ( N_noxref_17_c_5784_n N_noxref_21_c_6911_n ) capacitor c=0.00894156f \
 //x=48.645 //y=1.915 //x2=66.115 //y2=2.22
cc_3939 ( N_noxref_17_c_5794_n N_noxref_21_c_6911_n ) capacitor c=0.00894156f \
 //x=58.635 //y=1.915 //x2=66.115 //y2=2.22
cc_3940 ( N_noxref_17_c_5805_n N_noxref_21_c_6942_n ) capacitor c=2.97874e-19 \
 //x=44.535 //y=5.155 //x2=42.18 //y2=2.22
cc_3941 ( N_noxref_17_c_5873_n N_noxref_23_c_7498_n ) capacitor c=0.0110781f \
 //x=48.725 //y=3.7 //x2=70.185 //y2=2.96
cc_3942 ( N_noxref_17_c_5874_n N_noxref_23_c_7498_n ) capacitor c=7.98411e-19 \
 //x=47.105 //y=3.7 //x2=70.185 //y2=2.96
cc_3943 ( N_noxref_17_c_5847_n N_noxref_23_c_7498_n ) capacitor c=0.232839f \
 //x=58.715 //y=3.7 //x2=70.185 //y2=2.96
cc_3944 ( N_noxref_17_c_5848_n N_noxref_23_c_7498_n ) capacitor c=5.76555e-19 \
 //x=48.955 //y=3.7 //x2=70.185 //y2=2.96
cc_3945 ( N_noxref_17_c_5815_n N_noxref_23_c_7498_n ) capacitor c=0.0187656f \
 //x=46.99 //y=3.7 //x2=70.185 //y2=2.96
cc_3946 ( N_noxref_17_c_5778_n N_noxref_23_c_7498_n ) capacitor c=0.0187412f \
 //x=48.84 //y=2.08 //x2=70.185 //y2=2.96
cc_3947 ( N_noxref_17_c_5779_n N_noxref_23_c_7498_n ) capacitor c=0.0236665f \
 //x=58.83 //y=2.08 //x2=70.185 //y2=2.96
cc_3948 ( N_noxref_17_M28_noxref_d N_noxref_40_M26_noxref_s ) capacitor \
 c=0.00309936f //x=46.315 //y=0.915 //x2=43.375 //y2=0.375
cc_3949 ( N_noxref_17_c_5777_n N_noxref_41_c_9000_n ) capacitor c=0.00457167f \
 //x=46.905 //y=1.665 //x2=46.905 //y2=0.54
cc_3950 ( N_noxref_17_M28_noxref_d N_noxref_41_c_9000_n ) capacitor \
 c=0.0115903f //x=46.315 //y=0.915 //x2=46.905 //y2=0.54
cc_3951 ( N_noxref_17_c_5990_p N_noxref_41_c_9013_n ) capacitor c=0.020048f \
 //x=46.59 //y=1.665 //x2=46.02 //y2=0.995
cc_3952 ( N_noxref_17_M28_noxref_d N_noxref_41_M27_noxref_d ) capacitor \
 c=5.27807e-19 //x=46.315 //y=0.915 //x2=44.78 //y2=0.91
cc_3953 ( N_noxref_17_c_5777_n N_noxref_41_M28_noxref_s ) capacitor \
 c=0.0196084f //x=46.905 //y=1.665 //x2=45.885 //y2=0.375
cc_3954 ( N_noxref_17_M28_noxref_d N_noxref_41_M28_noxref_s ) capacitor \
 c=0.0426444f //x=46.315 //y=0.915 //x2=45.885 //y2=0.375
cc_3955 ( N_noxref_17_c_5777_n N_noxref_42_c_9076_n ) capacitor c=3.04182e-19 \
 //x=46.905 //y=1.665 //x2=48.425 //y2=1.495
cc_3956 ( N_noxref_17_c_5784_n N_noxref_42_c_9076_n ) capacitor c=0.0034165f \
 //x=48.645 //y=1.915 //x2=48.425 //y2=1.495
cc_3957 ( N_noxref_17_c_5778_n N_noxref_42_c_9048_n ) capacitor c=0.0111916f \
 //x=48.84 //y=2.08 //x2=49.31 //y2=1.58
cc_3958 ( N_noxref_17_c_5783_n N_noxref_42_c_9048_n ) capacitor c=0.00696403f \
 //x=48.645 //y=1.52 //x2=49.31 //y2=1.58
cc_3959 ( N_noxref_17_c_5784_n N_noxref_42_c_9048_n ) capacitor c=0.0174694f \
 //x=48.645 //y=1.915 //x2=49.31 //y2=1.58
cc_3960 ( N_noxref_17_c_5786_n N_noxref_42_c_9048_n ) capacitor c=0.00776811f \
 //x=49.02 //y=1.365 //x2=49.31 //y2=1.58
cc_3961 ( N_noxref_17_c_5789_n N_noxref_42_c_9048_n ) capacitor c=0.00339872f \
 //x=49.175 //y=1.21 //x2=49.31 //y2=1.58
cc_3962 ( N_noxref_17_c_5784_n N_noxref_42_c_9055_n ) capacitor c=6.71402e-19 \
 //x=48.645 //y=1.915 //x2=49.395 //y2=1.495
cc_3963 ( N_noxref_17_c_5780_n N_noxref_42_M29_noxref_s ) capacitor \
 c=0.0327502f //x=48.645 //y=0.865 //x2=48.29 //y2=0.365
cc_3964 ( N_noxref_17_c_5783_n N_noxref_42_M29_noxref_s ) capacitor \
 c=3.48408e-19 //x=48.645 //y=1.52 //x2=48.29 //y2=0.365
cc_3965 ( N_noxref_17_c_5787_n N_noxref_42_M29_noxref_s ) capacitor \
 c=0.0120759f //x=49.175 //y=0.865 //x2=48.29 //y2=0.365
cc_3966 ( N_noxref_17_c_5794_n N_noxref_45_c_9223_n ) capacitor c=0.0034165f \
 //x=58.635 //y=1.915 //x2=58.415 //y2=1.495
cc_3967 ( N_noxref_17_c_5779_n N_noxref_45_c_9204_n ) capacitor c=0.0111916f \
 //x=58.83 //y=2.08 //x2=59.3 //y2=1.58
cc_3968 ( N_noxref_17_c_5793_n N_noxref_45_c_9204_n ) capacitor c=0.00696403f \
 //x=58.635 //y=1.52 //x2=59.3 //y2=1.58
cc_3969 ( N_noxref_17_c_5794_n N_noxref_45_c_9204_n ) capacitor c=0.0174694f \
 //x=58.635 //y=1.915 //x2=59.3 //y2=1.58
cc_3970 ( N_noxref_17_c_5796_n N_noxref_45_c_9204_n ) capacitor c=0.00776811f \
 //x=59.01 //y=1.365 //x2=59.3 //y2=1.58
cc_3971 ( N_noxref_17_c_5799_n N_noxref_45_c_9204_n ) capacitor c=0.00339872f \
 //x=59.165 //y=1.21 //x2=59.3 //y2=1.58
cc_3972 ( N_noxref_17_c_5794_n N_noxref_45_c_9211_n ) capacitor c=6.71402e-19 \
 //x=58.635 //y=1.915 //x2=59.385 //y2=1.495
cc_3973 ( N_noxref_17_c_5790_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.0326577f //x=58.635 //y=0.865 //x2=58.28 //y2=0.365
cc_3974 ( N_noxref_17_c_5793_n N_noxref_45_M35_noxref_s ) capacitor \
 c=3.48408e-19 //x=58.635 //y=1.52 //x2=58.28 //y2=0.365
cc_3975 ( N_noxref_17_c_5797_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.0120759f //x=59.165 //y=0.865 //x2=58.28 //y2=0.365
cc_3976 ( N_noxref_18_c_6048_n N_noxref_19_c_6215_n ) capacitor c=0.172652f \
 //x=62.045 //y=4.44 //x2=62.785 //y2=4.07
cc_3977 ( N_noxref_18_c_6054_n N_noxref_19_c_6215_n ) capacitor c=0.0292297f \
 //x=60.425 //y=4.44 //x2=62.785 //y2=4.07
cc_3978 ( N_noxref_18_c_6057_n N_noxref_19_c_6215_n ) capacitor c=0.0128589f \
 //x=59.745 //y=5.2 //x2=62.785 //y2=4.07
cc_3979 ( N_noxref_18_c_6061_n N_noxref_19_c_6215_n ) capacitor c=0.013796f \
 //x=59.035 //y=5.2 //x2=62.785 //y2=4.07
cc_3980 ( N_noxref_18_c_6033_n N_noxref_19_c_6215_n ) capacitor c=0.0200095f \
 //x=60.31 //y=4.44 //x2=62.785 //y2=4.07
cc_3981 ( N_noxref_18_c_6034_n N_noxref_19_c_6215_n ) capacitor c=0.0221104f \
 //x=62.16 //y=2.08 //x2=62.785 //y2=4.07
cc_3982 ( N_noxref_18_c_6076_n N_noxref_19_c_6215_n ) capacitor c=0.00536694f \
 //x=62.16 //y=4.7 //x2=62.785 //y2=4.07
cc_3983 ( N_noxref_18_c_6033_n N_noxref_19_c_6194_n ) capacitor c=3.49822e-19 \
 //x=60.31 //y=4.44 //x2=56.98 //y2=4.07
cc_3984 ( N_noxref_18_c_6034_n N_noxref_19_c_6440_n ) capacitor c=0.00400249f \
 //x=62.16 //y=2.08 //x2=62.9 //y2=4.535
cc_3985 ( N_noxref_18_c_6076_n N_noxref_19_c_6440_n ) capacitor c=0.00417994f \
 //x=62.16 //y=4.7 //x2=62.9 //y2=4.535
cc_3986 ( N_noxref_18_c_6048_n N_noxref_19_c_6195_n ) capacitor c=0.00467582f \
 //x=62.045 //y=4.44 //x2=62.9 //y2=2.08
cc_3987 ( N_noxref_18_c_6033_n N_noxref_19_c_6195_n ) capacitor c=7.60135e-19 \
 //x=60.31 //y=4.44 //x2=62.9 //y2=2.08
cc_3988 ( N_noxref_18_c_6034_n N_noxref_19_c_6195_n ) capacitor c=0.0771278f \
 //x=62.16 //y=2.08 //x2=62.9 //y2=2.08
cc_3989 ( N_noxref_18_c_6039_n N_noxref_19_c_6195_n ) capacitor c=0.00284029f \
 //x=61.965 //y=1.915 //x2=62.9 //y2=2.08
cc_3990 ( N_noxref_18_M119_noxref_g N_noxref_19_M121_noxref_g ) capacitor \
 c=0.0104611f //x=62.06 //y=6.02 //x2=62.94 //y2=6.02
cc_3991 ( N_noxref_18_M120_noxref_g N_noxref_19_M121_noxref_g ) capacitor \
 c=0.106811f //x=62.5 //y=6.02 //x2=62.94 //y2=6.02
cc_3992 ( N_noxref_18_M120_noxref_g N_noxref_19_M122_noxref_g ) capacitor \
 c=0.0100341f //x=62.5 //y=6.02 //x2=63.38 //y2=6.02
cc_3993 ( N_noxref_18_c_6035_n N_noxref_19_c_6449_n ) capacitor c=4.86506e-19 \
 //x=61.965 //y=0.865 //x2=62.935 //y2=0.905
cc_3994 ( N_noxref_18_c_6037_n N_noxref_19_c_6449_n ) capacitor c=0.00152104f \
 //x=61.965 //y=1.21 //x2=62.935 //y2=0.905
cc_3995 ( N_noxref_18_c_6042_n N_noxref_19_c_6449_n ) capacitor c=0.0151475f \
 //x=62.495 //y=0.865 //x2=62.935 //y2=0.905
cc_3996 ( N_noxref_18_c_6038_n N_noxref_19_c_6452_n ) capacitor c=0.00109982f \
 //x=61.965 //y=1.52 //x2=62.935 //y2=1.25
cc_3997 ( N_noxref_18_c_6044_n N_noxref_19_c_6452_n ) capacitor c=0.0111064f \
 //x=62.495 //y=1.21 //x2=62.935 //y2=1.25
cc_3998 ( N_noxref_18_c_6038_n N_noxref_19_c_6454_n ) capacitor c=9.57794e-19 \
 //x=61.965 //y=1.52 //x2=62.935 //y2=1.56
cc_3999 ( N_noxref_18_c_6039_n N_noxref_19_c_6454_n ) capacitor c=0.00662747f \
 //x=61.965 //y=1.915 //x2=62.935 //y2=1.56
cc_4000 ( N_noxref_18_c_6044_n N_noxref_19_c_6454_n ) capacitor c=0.00862358f \
 //x=62.495 //y=1.21 //x2=62.935 //y2=1.56
cc_4001 ( N_noxref_18_c_6042_n N_noxref_19_c_6457_n ) capacitor c=0.00124821f \
 //x=62.495 //y=0.865 //x2=63.465 //y2=0.905
cc_4002 ( N_noxref_18_c_6044_n N_noxref_19_c_6458_n ) capacitor c=0.00200715f \
 //x=62.495 //y=1.21 //x2=63.465 //y2=1.25
cc_4003 ( N_noxref_18_c_6034_n N_noxref_19_c_6459_n ) capacitor c=0.00282278f \
 //x=62.16 //y=2.08 //x2=62.9 //y2=2.08
cc_4004 ( N_noxref_18_c_6039_n N_noxref_19_c_6459_n ) capacitor c=0.0172771f \
 //x=61.965 //y=1.915 //x2=62.9 //y2=2.08
cc_4005 ( N_noxref_18_c_6034_n N_noxref_19_c_6461_n ) capacitor c=0.00343287f \
 //x=62.16 //y=2.08 //x2=62.93 //y2=4.7
cc_4006 ( N_noxref_18_c_6076_n N_noxref_19_c_6461_n ) capacitor c=0.0293367f \
 //x=62.16 //y=4.7 //x2=62.93 //y2=4.7
cc_4007 ( N_noxref_18_c_6048_n N_noxref_20_c_6592_n ) capacitor c=0.0104216f \
 //x=62.045 //y=4.44 //x2=63.525 //y2=3.7
cc_4008 ( N_noxref_18_c_6054_n N_noxref_20_c_6592_n ) capacitor c=8.92918e-19 \
 //x=60.425 //y=4.44 //x2=63.525 //y2=3.7
cc_4009 ( N_noxref_18_c_6033_n N_noxref_20_c_6592_n ) capacitor c=0.0211091f \
 //x=60.31 //y=4.44 //x2=63.525 //y2=3.7
cc_4010 ( N_noxref_18_c_6034_n N_noxref_20_c_6592_n ) capacitor c=0.0210613f \
 //x=62.16 //y=2.08 //x2=63.525 //y2=3.7
cc_4011 ( N_noxref_18_c_6033_n N_noxref_20_c_6653_n ) capacitor c=0.00117715f \
 //x=60.31 //y=4.44 //x2=59.685 //y2=3.7
cc_4012 ( N_noxref_18_c_6048_n N_noxref_20_c_6602_n ) capacitor c=0.00550845f \
 //x=62.045 //y=4.44 //x2=65.235 //y2=4.44
cc_4013 ( N_noxref_18_c_6054_n N_noxref_20_c_6655_n ) capacitor c=4.57222e-19 \
 //x=60.425 //y=4.44 //x2=59.57 //y2=4.535
cc_4014 ( N_noxref_18_c_6057_n N_noxref_20_c_6655_n ) capacitor c=0.0129336f \
 //x=59.745 //y=5.2 //x2=59.57 //y2=4.535
cc_4015 ( N_noxref_18_c_6033_n N_noxref_20_c_6655_n ) capacitor c=0.00985792f \
 //x=60.31 //y=4.44 //x2=59.57 //y2=4.535
cc_4016 ( N_noxref_18_c_6054_n N_noxref_20_c_6560_n ) capacitor c=0.00463722f \
 //x=60.425 //y=4.44 //x2=59.57 //y2=2.08
cc_4017 ( N_noxref_18_c_6033_n N_noxref_20_c_6560_n ) capacitor c=0.0715836f \
 //x=60.31 //y=4.44 //x2=59.57 //y2=2.08
cc_4018 ( N_noxref_18_c_6034_n N_noxref_20_c_6560_n ) capacitor c=6.89521e-19 \
 //x=62.16 //y=2.08 //x2=59.57 //y2=2.08
cc_4019 ( N_noxref_18_M120_noxref_g N_noxref_20_c_6608_n ) capacitor \
 c=0.017965f //x=62.5 //y=6.02 //x2=63.075 //y2=5.2
cc_4020 ( N_noxref_18_c_6048_n N_noxref_20_c_6612_n ) capacitor c=0.00218812f \
 //x=62.045 //y=4.44 //x2=62.365 //y2=5.2
cc_4021 ( N_noxref_18_c_6034_n N_noxref_20_c_6612_n ) capacitor c=0.00520726f \
 //x=62.16 //y=2.08 //x2=62.365 //y2=5.2
cc_4022 ( N_noxref_18_M119_noxref_g N_noxref_20_c_6612_n ) capacitor \
 c=0.0177326f //x=62.06 //y=6.02 //x2=62.365 //y2=5.2
cc_4023 ( N_noxref_18_c_6076_n N_noxref_20_c_6612_n ) capacitor c=0.00581512f \
 //x=62.16 //y=4.7 //x2=62.365 //y2=5.2
cc_4024 ( N_noxref_18_c_6033_n N_noxref_20_c_6563_n ) capacitor c=3.49822e-19 \
 //x=60.31 //y=4.44 //x2=63.64 //y2=3.7
cc_4025 ( N_noxref_18_c_6034_n N_noxref_20_c_6563_n ) capacitor c=0.00358999f \
 //x=62.16 //y=2.08 //x2=63.64 //y2=3.7
cc_4026 ( N_noxref_18_c_6057_n N_noxref_20_M117_noxref_g ) capacitor \
 c=0.0166421f //x=59.745 //y=5.2 //x2=59.61 //y2=6.02
cc_4027 ( N_noxref_18_M117_noxref_d N_noxref_20_M117_noxref_g ) capacitor \
 c=0.0173476f //x=59.685 //y=5.02 //x2=59.61 //y2=6.02
cc_4028 ( N_noxref_18_c_6063_n N_noxref_20_M118_noxref_g ) capacitor \
 c=0.0199348f //x=60.225 //y=5.2 //x2=60.05 //y2=6.02
cc_4029 ( N_noxref_18_M117_noxref_d N_noxref_20_M118_noxref_g ) capacitor \
 c=0.0179769f //x=59.685 //y=5.02 //x2=60.05 //y2=6.02
cc_4030 ( N_noxref_18_M36_noxref_d N_noxref_20_c_6663_n ) capacitor \
 c=0.00217566f //x=59.68 //y=0.905 //x2=59.605 //y2=0.905
cc_4031 ( N_noxref_18_M36_noxref_d N_noxref_20_c_6666_n ) capacitor \
 c=0.0034598f //x=59.68 //y=0.905 //x2=59.605 //y2=1.25
cc_4032 ( N_noxref_18_M36_noxref_d N_noxref_20_c_6668_n ) capacitor \
 c=0.00669531f //x=59.68 //y=0.905 //x2=59.605 //y2=1.56
cc_4033 ( N_noxref_18_c_6033_n N_noxref_20_c_6703_n ) capacitor c=0.0142673f \
 //x=60.31 //y=4.44 //x2=59.975 //y2=4.79
cc_4034 ( N_noxref_18_c_6153_p N_noxref_20_c_6703_n ) capacitor c=0.00408717f \
 //x=59.83 //y=5.2 //x2=59.975 //y2=4.79
cc_4035 ( N_noxref_18_M36_noxref_d N_noxref_20_c_6705_n ) capacitor \
 c=0.00241102f //x=59.68 //y=0.905 //x2=59.98 //y2=0.75
cc_4036 ( N_noxref_18_c_6032_n N_noxref_20_c_6706_n ) capacitor c=0.00371277f \
 //x=60.225 //y=1.655 //x2=59.98 //y2=1.405
cc_4037 ( N_noxref_18_M36_noxref_d N_noxref_20_c_6706_n ) capacitor \
 c=0.0137169f //x=59.68 //y=0.905 //x2=59.98 //y2=1.405
cc_4038 ( N_noxref_18_M36_noxref_d N_noxref_20_c_6671_n ) capacitor \
 c=0.00132245f //x=59.68 //y=0.905 //x2=60.135 //y2=0.905
cc_4039 ( N_noxref_18_c_6032_n N_noxref_20_c_6672_n ) capacitor c=0.00457401f \
 //x=60.225 //y=1.655 //x2=60.135 //y2=1.25
cc_4040 ( N_noxref_18_M36_noxref_d N_noxref_20_c_6672_n ) capacitor \
 c=0.00566463f //x=59.68 //y=0.905 //x2=60.135 //y2=1.25
cc_4041 ( N_noxref_18_c_6033_n N_noxref_20_c_6673_n ) capacitor c=0.00731987f \
 //x=60.31 //y=4.44 //x2=59.57 //y2=2.08
cc_4042 ( N_noxref_18_c_6033_n N_noxref_20_c_6712_n ) capacitor c=0.00306024f \
 //x=60.31 //y=4.44 //x2=59.57 //y2=1.915
cc_4043 ( N_noxref_18_M36_noxref_d N_noxref_20_c_6712_n ) capacitor \
 c=0.00660593f //x=59.68 //y=0.905 //x2=59.57 //y2=1.915
cc_4044 ( N_noxref_18_c_6054_n N_noxref_20_c_6675_n ) capacitor c=4.521e-19 \
 //x=60.425 //y=4.44 //x2=59.6 //y2=4.7
cc_4045 ( N_noxref_18_c_6057_n N_noxref_20_c_6675_n ) capacitor c=0.00346635f \
 //x=59.745 //y=5.2 //x2=59.6 //y2=4.7
cc_4046 ( N_noxref_18_c_6033_n N_noxref_20_c_6675_n ) capacitor c=0.00517603f \
 //x=60.31 //y=4.44 //x2=59.6 //y2=4.7
cc_4047 ( N_noxref_18_M120_noxref_g N_noxref_20_M119_noxref_d ) capacitor \
 c=0.0173476f //x=62.5 //y=6.02 //x2=62.135 //y2=5.02
cc_4048 ( N_noxref_18_c_6167_p N_noxref_21_c_6911_n ) capacitor c=0.0146822f \
 //x=59.955 //y=1.655 //x2=66.115 //y2=2.22
cc_4049 ( N_noxref_18_c_6033_n N_noxref_21_c_6911_n ) capacitor c=0.0222456f \
 //x=60.31 //y=4.44 //x2=66.115 //y2=2.22
cc_4050 ( N_noxref_18_c_6034_n N_noxref_21_c_6911_n ) capacitor c=0.0208418f \
 //x=62.16 //y=2.08 //x2=66.115 //y2=2.22
cc_4051 ( N_noxref_18_c_6039_n N_noxref_21_c_6911_n ) capacitor c=0.00894156f \
 //x=61.965 //y=1.915 //x2=66.115 //y2=2.22
cc_4052 ( N_noxref_18_c_6033_n N_noxref_23_c_7498_n ) capacitor c=0.0234416f \
 //x=60.31 //y=4.44 //x2=70.185 //y2=2.96
cc_4053 ( N_noxref_18_c_6034_n N_noxref_23_c_7498_n ) capacitor c=0.0233753f \
 //x=62.16 //y=2.08 //x2=70.185 //y2=2.96
cc_4054 ( N_noxref_18_c_6167_p N_noxref_45_c_9223_n ) capacitor c=3.15806e-19 \
 //x=59.955 //y=1.655 //x2=58.415 //y2=1.495
cc_4055 ( N_noxref_18_c_6167_p N_noxref_45_c_9211_n ) capacitor c=0.0203424f \
 //x=59.955 //y=1.655 //x2=59.385 //y2=1.495
cc_4056 ( N_noxref_18_c_6032_n N_noxref_45_c_9212_n ) capacitor c=0.00457164f \
 //x=60.225 //y=1.655 //x2=60.27 //y2=0.53
cc_4057 ( N_noxref_18_M36_noxref_d N_noxref_45_c_9212_n ) capacitor \
 c=0.0115831f //x=59.68 //y=0.905 //x2=60.27 //y2=0.53
cc_4058 ( N_noxref_18_c_6032_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.013435f //x=60.225 //y=1.655 //x2=58.28 //y2=0.365
cc_4059 ( N_noxref_18_M36_noxref_d N_noxref_45_M35_noxref_s ) capacitor \
 c=0.043966f //x=59.68 //y=0.905 //x2=58.28 //y2=0.365
cc_4060 ( N_noxref_18_c_6032_n N_noxref_46_c_9275_n ) capacitor c=3.22188e-19 \
 //x=60.225 //y=1.655 //x2=61.745 //y2=1.495
cc_4061 ( N_noxref_18_c_6039_n N_noxref_46_c_9275_n ) capacitor c=0.0034165f \
 //x=61.965 //y=1.915 //x2=61.745 //y2=1.495
cc_4062 ( N_noxref_18_c_6034_n N_noxref_46_c_9256_n ) capacitor c=0.011618f \
 //x=62.16 //y=2.08 //x2=62.63 //y2=1.58
cc_4063 ( N_noxref_18_c_6038_n N_noxref_46_c_9256_n ) capacitor c=0.00696403f \
 //x=61.965 //y=1.52 //x2=62.63 //y2=1.58
cc_4064 ( N_noxref_18_c_6039_n N_noxref_46_c_9256_n ) capacitor c=0.0174694f \
 //x=61.965 //y=1.915 //x2=62.63 //y2=1.58
cc_4065 ( N_noxref_18_c_6041_n N_noxref_46_c_9256_n ) capacitor c=0.00776811f \
 //x=62.34 //y=1.365 //x2=62.63 //y2=1.58
cc_4066 ( N_noxref_18_c_6044_n N_noxref_46_c_9256_n ) capacitor c=0.00339872f \
 //x=62.495 //y=1.21 //x2=62.63 //y2=1.58
cc_4067 ( N_noxref_18_c_6039_n N_noxref_46_c_9263_n ) capacitor c=6.71402e-19 \
 //x=61.965 //y=1.915 //x2=62.715 //y2=1.495
cc_4068 ( N_noxref_18_c_6035_n N_noxref_46_M37_noxref_s ) capacitor \
 c=0.0326577f //x=61.965 //y=0.865 //x2=61.61 //y2=0.365
cc_4069 ( N_noxref_18_c_6038_n N_noxref_46_M37_noxref_s ) capacitor \
 c=3.48408e-19 //x=61.965 //y=1.52 //x2=61.61 //y2=0.365
cc_4070 ( N_noxref_18_c_6042_n N_noxref_46_M37_noxref_s ) capacitor \
 c=0.0120759f //x=62.495 //y=0.865 //x2=61.61 //y2=0.365
cc_4071 ( N_noxref_19_c_6215_n N_noxref_20_c_6592_n ) capacitor c=0.304477f \
 //x=62.785 //y=4.07 //x2=63.525 //y2=3.7
cc_4072 ( N_noxref_19_c_6195_n N_noxref_20_c_6592_n ) capacitor c=0.0211371f \
 //x=62.9 //y=2.08 //x2=63.525 //y2=3.7
cc_4073 ( N_noxref_19_c_6465_p N_noxref_20_c_6592_n ) capacitor c=0.00624857f \
 //x=63.305 //y=4.79 //x2=63.525 //y2=3.7
cc_4074 ( N_noxref_19_c_6461_n N_noxref_20_c_6592_n ) capacitor c=2.85902e-19 \
 //x=62.93 //y=4.7 //x2=63.525 //y2=3.7
cc_4075 ( N_noxref_19_c_6215_n N_noxref_20_c_6653_n ) capacitor c=0.0291169f \
 //x=62.785 //y=4.07 //x2=59.685 //y2=3.7
cc_4076 ( N_noxref_19_c_6195_n N_noxref_20_c_6595_n ) capacitor c=0.00117715f \
 //x=62.9 //y=2.08 //x2=63.755 //y2=3.7
cc_4077 ( N_noxref_19_c_6215_n N_noxref_20_c_6655_n ) capacitor c=0.00135863f \
 //x=62.785 //y=4.07 //x2=59.57 //y2=4.535
cc_4078 ( N_noxref_19_c_6215_n N_noxref_20_c_6560_n ) capacitor c=0.022647f \
 //x=62.785 //y=4.07 //x2=59.57 //y2=2.08
cc_4079 ( N_noxref_19_c_6194_n N_noxref_20_c_6560_n ) capacitor c=6.84853e-19 \
 //x=56.98 //y=4.07 //x2=59.57 //y2=2.08
cc_4080 ( N_noxref_19_c_6215_n N_noxref_20_c_6608_n ) capacitor c=0.00208151f \
 //x=62.785 //y=4.07 //x2=63.075 //y2=5.2
cc_4081 ( N_noxref_19_c_6440_n N_noxref_20_c_6608_n ) capacitor c=0.0129794f \
 //x=62.9 //y=4.535 //x2=63.075 //y2=5.2
cc_4082 ( N_noxref_19_M121_noxref_g N_noxref_20_c_6608_n ) capacitor \
 c=0.0166421f //x=62.94 //y=6.02 //x2=63.075 //y2=5.2
cc_4083 ( N_noxref_19_c_6461_n N_noxref_20_c_6608_n ) capacitor c=0.00346627f \
 //x=62.93 //y=4.7 //x2=63.075 //y2=5.2
cc_4084 ( N_noxref_19_c_6215_n N_noxref_20_c_6612_n ) capacitor c=0.0118122f \
 //x=62.785 //y=4.07 //x2=62.365 //y2=5.2
cc_4085 ( N_noxref_19_M122_noxref_g N_noxref_20_c_6614_n ) capacitor \
 c=0.0206783f //x=63.38 //y=6.02 //x2=63.555 //y2=5.2
cc_4086 ( N_noxref_19_c_6478_p N_noxref_20_c_6562_n ) capacitor c=0.00371277f \
 //x=63.31 //y=1.405 //x2=63.555 //y2=1.655
cc_4087 ( N_noxref_19_c_6458_n N_noxref_20_c_6562_n ) capacitor c=0.00457401f \
 //x=63.465 //y=1.25 //x2=63.555 //y2=1.655
cc_4088 ( N_noxref_19_c_6215_n N_noxref_20_c_6563_n ) capacitor c=0.00465962f \
 //x=62.785 //y=4.07 //x2=63.64 //y2=3.7
cc_4089 ( N_noxref_19_c_6440_n N_noxref_20_c_6563_n ) capacitor c=0.010101f \
 //x=62.9 //y=4.535 //x2=63.64 //y2=3.7
cc_4090 ( N_noxref_19_c_6195_n N_noxref_20_c_6563_n ) capacitor c=0.0740686f \
 //x=62.9 //y=2.08 //x2=63.64 //y2=3.7
cc_4091 ( N_noxref_19_c_6465_p N_noxref_20_c_6563_n ) capacitor c=0.0142673f \
 //x=63.305 //y=4.79 //x2=63.64 //y2=3.7
cc_4092 ( N_noxref_19_c_6459_n N_noxref_20_c_6563_n ) capacitor c=0.00709342f \
 //x=62.9 //y=2.08 //x2=63.64 //y2=3.7
cc_4093 ( N_noxref_19_c_6485_p N_noxref_20_c_6563_n ) capacitor c=0.00306024f \
 //x=62.9 //y=1.915 //x2=63.64 //y2=3.7
cc_4094 ( N_noxref_19_c_6461_n N_noxref_20_c_6563_n ) capacitor c=0.00517969f \
 //x=62.93 //y=4.7 //x2=63.64 //y2=3.7
cc_4095 ( N_noxref_19_c_6195_n N_noxref_20_c_6564_n ) capacitor c=8.75643e-19 \
 //x=62.9 //y=2.08 //x2=65.12 //y2=2.08
cc_4096 ( N_noxref_19_c_6465_p N_noxref_20_c_6743_n ) capacitor c=0.00421574f \
 //x=63.305 //y=4.79 //x2=63.16 //y2=5.2
cc_4097 ( N_noxref_19_c_6215_n N_noxref_20_c_6703_n ) capacitor c=0.00756255f \
 //x=62.785 //y=4.07 //x2=59.975 //y2=4.79
cc_4098 ( N_noxref_19_c_6215_n N_noxref_20_c_6675_n ) capacitor c=0.00160199f \
 //x=62.785 //y=4.07 //x2=59.6 //y2=4.7
cc_4099 ( N_noxref_19_c_6449_n N_noxref_20_M38_noxref_d ) capacitor \
 c=0.00217566f //x=62.935 //y=0.905 //x2=63.01 //y2=0.905
cc_4100 ( N_noxref_19_c_6452_n N_noxref_20_M38_noxref_d ) capacitor \
 c=0.0034598f //x=62.935 //y=1.25 //x2=63.01 //y2=0.905
cc_4101 ( N_noxref_19_c_6454_n N_noxref_20_M38_noxref_d ) capacitor \
 c=0.00669531f //x=62.935 //y=1.56 //x2=63.01 //y2=0.905
cc_4102 ( N_noxref_19_c_6494_p N_noxref_20_M38_noxref_d ) capacitor \
 c=0.00241102f //x=63.31 //y=0.75 //x2=63.01 //y2=0.905
cc_4103 ( N_noxref_19_c_6478_p N_noxref_20_M38_noxref_d ) capacitor \
 c=0.0137169f //x=63.31 //y=1.405 //x2=63.01 //y2=0.905
cc_4104 ( N_noxref_19_c_6457_n N_noxref_20_M38_noxref_d ) capacitor \
 c=0.00132245f //x=63.465 //y=0.905 //x2=63.01 //y2=0.905
cc_4105 ( N_noxref_19_c_6458_n N_noxref_20_M38_noxref_d ) capacitor \
 c=0.00566463f //x=63.465 //y=1.25 //x2=63.01 //y2=0.905
cc_4106 ( N_noxref_19_c_6485_p N_noxref_20_M38_noxref_d ) capacitor \
 c=0.00660593f //x=62.9 //y=1.915 //x2=63.01 //y2=0.905
cc_4107 ( N_noxref_19_M121_noxref_g N_noxref_20_M121_noxref_d ) capacitor \
 c=0.0173477f //x=62.94 //y=6.02 //x2=63.015 //y2=5.02
cc_4108 ( N_noxref_19_M122_noxref_g N_noxref_20_M121_noxref_d ) capacitor \
 c=0.0179769f //x=63.38 //y=6.02 //x2=63.015 //y2=5.02
cc_4109 ( N_noxref_19_c_6215_n N_noxref_21_c_6911_n ) capacitor c=0.00190245f \
 //x=62.785 //y=4.07 //x2=66.115 //y2=2.22
cc_4110 ( N_noxref_19_c_6190_n N_noxref_21_c_6911_n ) capacitor c=0.0192695f \
 //x=44.03 //y=2.08 //x2=66.115 //y2=2.22
cc_4111 ( N_noxref_19_c_6191_n N_noxref_21_c_6911_n ) capacitor c=0.0201924f \
 //x=52.91 //y=2.08 //x2=66.115 //y2=2.22
cc_4112 ( N_noxref_19_c_6504_p N_noxref_21_c_6911_n ) capacitor c=0.0146822f \
 //x=56.625 //y=1.655 //x2=66.115 //y2=2.22
cc_4113 ( N_noxref_19_c_6194_n N_noxref_21_c_6911_n ) capacitor c=0.0222456f \
 //x=56.98 //y=4.07 //x2=66.115 //y2=2.22
cc_4114 ( N_noxref_19_c_6195_n N_noxref_21_c_6911_n ) capacitor c=0.0201924f \
 //x=62.9 //y=2.08 //x2=66.115 //y2=2.22
cc_4115 ( N_noxref_19_c_6201_n N_noxref_21_c_6911_n ) capacitor c=0.011987f \
 //x=43.73 //y=1.915 //x2=66.115 //y2=2.22
cc_4116 ( N_noxref_19_c_6335_n N_noxref_21_c_6911_n ) capacitor c=3.11115e-19 \
 //x=53.32 //y=1.405 //x2=66.115 //y2=2.22
cc_4117 ( N_noxref_19_c_6478_p N_noxref_21_c_6911_n ) capacitor c=3.11115e-19 \
 //x=63.31 //y=1.405 //x2=66.115 //y2=2.22
cc_4118 ( N_noxref_19_c_6305_n N_noxref_21_c_6911_n ) capacitor c=0.00570799f \
 //x=52.91 //y=2.08 //x2=66.115 //y2=2.22
cc_4119 ( N_noxref_19_c_6459_n N_noxref_21_c_6911_n ) capacitor c=0.00570799f \
 //x=62.9 //y=2.08 //x2=66.115 //y2=2.22
cc_4120 ( N_noxref_19_c_6215_n N_noxref_21_c_6956_n ) capacitor c=0.0048081f \
 //x=62.785 //y=4.07 //x2=66.345 //y2=4.07
cc_4121 ( N_noxref_19_c_6212_n N_noxref_21_c_6942_n ) capacitor c=0.00103915f \
 //x=44.145 //y=4.07 //x2=42.18 //y2=2.22
cc_4122 ( N_noxref_19_c_6190_n N_noxref_21_c_6942_n ) capacitor c=0.0150916f \
 //x=44.03 //y=2.08 //x2=42.18 //y2=2.22
cc_4123 ( N_noxref_19_c_6210_n N_noxref_23_c_7498_n ) capacitor c=0.0615741f \
 //x=52.795 //y=4.07 //x2=70.185 //y2=2.96
cc_4124 ( N_noxref_19_c_6212_n N_noxref_23_c_7498_n ) capacitor c=0.00776275f \
 //x=44.145 //y=4.07 //x2=70.185 //y2=2.96
cc_4125 ( N_noxref_19_c_6213_n N_noxref_23_c_7498_n ) capacitor c=0.0112822f \
 //x=56.865 //y=4.07 //x2=70.185 //y2=2.96
cc_4126 ( N_noxref_19_c_6284_n N_noxref_23_c_7498_n ) capacitor c=3.56521e-19 \
 //x=53.025 //y=4.07 //x2=70.185 //y2=2.96
cc_4127 ( N_noxref_19_c_6215_n N_noxref_23_c_7498_n ) capacitor c=0.037151f \
 //x=62.785 //y=4.07 //x2=70.185 //y2=2.96
cc_4128 ( N_noxref_19_c_6222_n N_noxref_23_c_7498_n ) capacitor c=4.50823e-19 \
 //x=57.095 //y=4.07 //x2=70.185 //y2=2.96
cc_4129 ( N_noxref_19_c_6190_n N_noxref_23_c_7498_n ) capacitor c=0.0237066f \
 //x=44.03 //y=2.08 //x2=70.185 //y2=2.96
cc_4130 ( N_noxref_19_c_6191_n N_noxref_23_c_7498_n ) capacitor c=0.0215847f \
 //x=52.91 //y=2.08 //x2=70.185 //y2=2.96
cc_4131 ( N_noxref_19_c_6194_n N_noxref_23_c_7498_n ) capacitor c=0.0234154f \
 //x=56.98 //y=4.07 //x2=70.185 //y2=2.96
cc_4132 ( N_noxref_19_c_6195_n N_noxref_23_c_7498_n ) capacitor c=0.0215847f \
 //x=62.9 //y=2.08 //x2=70.185 //y2=2.96
cc_4133 ( N_noxref_19_c_6201_n N_noxref_40_c_8970_n ) capacitor c=0.0034165f \
 //x=43.73 //y=1.915 //x2=43.51 //y2=1.505
cc_4134 ( N_noxref_19_c_6190_n N_noxref_40_c_8945_n ) capacitor c=0.0115578f \
 //x=44.03 //y=2.08 //x2=44.395 //y2=1.59
cc_4135 ( N_noxref_19_c_6200_n N_noxref_40_c_8945_n ) capacitor c=0.00697148f \
 //x=43.73 //y=1.53 //x2=44.395 //y2=1.59
cc_4136 ( N_noxref_19_c_6201_n N_noxref_40_c_8945_n ) capacitor c=0.0204849f \
 //x=43.73 //y=1.915 //x2=44.395 //y2=1.59
cc_4137 ( N_noxref_19_c_6203_n N_noxref_40_c_8945_n ) capacitor c=0.00610316f \
 //x=44.105 //y=1.375 //x2=44.395 //y2=1.59
cc_4138 ( N_noxref_19_c_6206_n N_noxref_40_c_8945_n ) capacitor c=0.00698822f \
 //x=44.26 //y=1.22 //x2=44.395 //y2=1.59
cc_4139 ( N_noxref_19_c_6197_n N_noxref_40_M26_noxref_s ) capacitor \
 c=0.0327271f //x=43.73 //y=0.875 //x2=43.375 //y2=0.375
cc_4140 ( N_noxref_19_c_6200_n N_noxref_40_M26_noxref_s ) capacitor \
 c=7.99997e-19 //x=43.73 //y=1.53 //x2=43.375 //y2=0.375
cc_4141 ( N_noxref_19_c_6201_n N_noxref_40_M26_noxref_s ) capacitor \
 c=0.00122123f //x=43.73 //y=1.915 //x2=43.375 //y2=0.375
cc_4142 ( N_noxref_19_c_6204_n N_noxref_40_M26_noxref_s ) capacitor \
 c=0.0121427f //x=44.26 //y=0.875 //x2=43.375 //y2=0.375
cc_4143 ( N_noxref_19_c_6300_n N_noxref_43_c_9107_n ) capacitor c=0.00623646f \
 //x=52.945 //y=1.56 //x2=52.725 //y2=1.495
cc_4144 ( N_noxref_19_c_6305_n N_noxref_43_c_9107_n ) capacitor c=0.00173579f \
 //x=52.91 //y=2.08 //x2=52.725 //y2=1.495
cc_4145 ( N_noxref_19_c_6191_n N_noxref_43_c_9108_n ) capacitor c=0.00156605f \
 //x=52.91 //y=2.08 //x2=53.61 //y2=0.53
cc_4146 ( N_noxref_19_c_6295_n N_noxref_43_c_9108_n ) capacitor c=0.0188655f \
 //x=52.945 //y=0.905 //x2=53.61 //y2=0.53
cc_4147 ( N_noxref_19_c_6303_n N_noxref_43_c_9108_n ) capacitor c=0.00656458f \
 //x=53.475 //y=0.905 //x2=53.61 //y2=0.53
cc_4148 ( N_noxref_19_c_6305_n N_noxref_43_c_9108_n ) capacitor c=2.1838e-19 \
 //x=52.91 //y=2.08 //x2=53.61 //y2=0.53
cc_4149 ( N_noxref_19_c_6295_n N_noxref_43_M31_noxref_s ) capacitor \
 c=0.00623646f //x=52.945 //y=0.905 //x2=51.62 //y2=0.365
cc_4150 ( N_noxref_19_c_6303_n N_noxref_43_M31_noxref_s ) capacitor \
 c=0.0143002f //x=53.475 //y=0.905 //x2=51.62 //y2=0.365
cc_4151 ( N_noxref_19_c_6304_n N_noxref_43_M31_noxref_s ) capacitor \
 c=0.00290153f //x=53.475 //y=1.25 //x2=51.62 //y2=0.365
cc_4152 ( N_noxref_19_c_6504_p N_noxref_44_c_9171_n ) capacitor c=3.15806e-19 \
 //x=56.625 //y=1.655 //x2=55.085 //y2=1.495
cc_4153 ( N_noxref_19_c_6504_p N_noxref_44_c_9159_n ) capacitor c=0.0203424f \
 //x=56.625 //y=1.655 //x2=56.055 //y2=1.495
cc_4154 ( N_noxref_19_c_6193_n N_noxref_44_c_9160_n ) capacitor c=0.00457164f \
 //x=56.895 //y=1.655 //x2=56.94 //y2=0.53
cc_4155 ( N_noxref_19_M34_noxref_d N_noxref_44_c_9160_n ) capacitor \
 c=0.0115831f //x=56.35 //y=0.905 //x2=56.94 //y2=0.53
cc_4156 ( N_noxref_19_c_6193_n N_noxref_44_M33_noxref_s ) capacitor \
 c=0.013435f //x=56.895 //y=1.655 //x2=54.95 //y2=0.365
cc_4157 ( N_noxref_19_M34_noxref_d N_noxref_44_M33_noxref_s ) capacitor \
 c=0.043966f //x=56.35 //y=0.905 //x2=54.95 //y2=0.365
cc_4158 ( N_noxref_19_c_6193_n N_noxref_45_c_9223_n ) capacitor c=3.22188e-19 \
 //x=56.895 //y=1.655 //x2=58.415 //y2=1.495
cc_4159 ( N_noxref_19_c_6454_n N_noxref_46_c_9263_n ) capacitor c=0.00623646f \
 //x=62.935 //y=1.56 //x2=62.715 //y2=1.495
cc_4160 ( N_noxref_19_c_6459_n N_noxref_46_c_9263_n ) capacitor c=0.00173579f \
 //x=62.9 //y=2.08 //x2=62.715 //y2=1.495
cc_4161 ( N_noxref_19_c_6195_n N_noxref_46_c_9264_n ) capacitor c=0.00156605f \
 //x=62.9 //y=2.08 //x2=63.6 //y2=0.53
cc_4162 ( N_noxref_19_c_6449_n N_noxref_46_c_9264_n ) capacitor c=0.0188655f \
 //x=62.935 //y=0.905 //x2=63.6 //y2=0.53
cc_4163 ( N_noxref_19_c_6457_n N_noxref_46_c_9264_n ) capacitor c=0.00656458f \
 //x=63.465 //y=0.905 //x2=63.6 //y2=0.53
cc_4164 ( N_noxref_19_c_6459_n N_noxref_46_c_9264_n ) capacitor c=2.1838e-19 \
 //x=62.9 //y=2.08 //x2=63.6 //y2=0.53
cc_4165 ( N_noxref_19_c_6449_n N_noxref_46_M37_noxref_s ) capacitor \
 c=0.00623646f //x=62.935 //y=0.905 //x2=61.61 //y2=0.365
cc_4166 ( N_noxref_19_c_6457_n N_noxref_46_M37_noxref_s ) capacitor \
 c=0.0143002f //x=63.465 //y=0.905 //x2=61.61 //y2=0.365
cc_4167 ( N_noxref_19_c_6458_n N_noxref_46_M37_noxref_s ) capacitor \
 c=0.00290153f //x=63.465 //y=1.25 //x2=61.61 //y2=0.365
cc_4168 ( N_noxref_20_c_6592_n N_noxref_21_c_6911_n ) capacitor c=0.0125472f \
 //x=63.525 //y=3.7 //x2=66.115 //y2=2.22
cc_4169 ( N_noxref_20_c_6653_n N_noxref_21_c_6911_n ) capacitor c=4.44747e-19 \
 //x=59.685 //y=3.7 //x2=66.115 //y2=2.22
cc_4170 ( N_noxref_20_c_6593_n N_noxref_21_c_6911_n ) capacitor c=0.00281503f \
 //x=65.005 //y=3.7 //x2=66.115 //y2=2.22
cc_4171 ( N_noxref_20_c_6595_n N_noxref_21_c_6911_n ) capacitor c=2.67441e-19 \
 //x=63.755 //y=3.7 //x2=66.115 //y2=2.22
cc_4172 ( N_noxref_20_c_6597_n N_noxref_21_c_6911_n ) capacitor c=0.00268543f \
 //x=68.705 //y=4.44 //x2=66.115 //y2=2.22
cc_4173 ( N_noxref_20_c_6560_n N_noxref_21_c_6911_n ) capacitor c=0.0201924f \
 //x=59.57 //y=2.08 //x2=66.115 //y2=2.22
cc_4174 ( N_noxref_20_c_6762_p N_noxref_21_c_6911_n ) capacitor c=0.0146822f \
 //x=63.285 //y=1.655 //x2=66.115 //y2=2.22
cc_4175 ( N_noxref_20_c_6563_n N_noxref_21_c_6911_n ) capacitor c=0.0222456f \
 //x=63.64 //y=3.7 //x2=66.115 //y2=2.22
cc_4176 ( N_noxref_20_c_6564_n N_noxref_21_c_6911_n ) capacitor c=0.0223124f \
 //x=65.12 //y=2.08 //x2=66.115 //y2=2.22
cc_4177 ( N_noxref_20_c_6706_n N_noxref_21_c_6911_n ) capacitor c=3.11115e-19 \
 //x=59.98 //y=1.405 //x2=66.115 //y2=2.22
cc_4178 ( N_noxref_20_c_6673_n N_noxref_21_c_6911_n ) capacitor c=0.00570799f \
 //x=59.57 //y=2.08 //x2=66.115 //y2=2.22
cc_4179 ( N_noxref_20_c_6588_n N_noxref_21_c_6911_n ) capacitor c=0.00891908f \
 //x=65.12 //y=2.08 //x2=66.115 //y2=2.22
cc_4180 ( N_noxref_20_c_6597_n N_noxref_21_c_6938_n ) capacitor c=0.23799f \
 //x=68.705 //y=4.44 //x2=72.775 //y2=4.07
cc_4181 ( N_noxref_20_c_6567_n N_noxref_21_c_6938_n ) capacitor c=0.0258036f \
 //x=68.82 //y=2.08 //x2=72.775 //y2=4.07
cc_4182 ( N_noxref_20_c_6641_n N_noxref_21_c_6938_n ) capacitor c=0.00381677f \
 //x=68.82 //y=4.705 //x2=72.775 //y2=4.07
cc_4183 ( N_noxref_20_c_6597_n N_noxref_21_c_6956_n ) capacitor c=0.0289488f \
 //x=68.705 //y=4.44 //x2=66.345 //y2=4.07
cc_4184 ( N_noxref_20_c_6564_n N_noxref_21_c_6956_n ) capacitor c=0.0032662f \
 //x=65.12 //y=2.08 //x2=66.345 //y2=4.07
cc_4185 ( N_noxref_20_c_6597_n N_noxref_21_c_6970_n ) capacitor c=0.00210648f \
 //x=68.705 //y=4.44 //x2=66.23 //y2=4.54
cc_4186 ( N_noxref_20_c_6564_n N_noxref_21_c_6970_n ) capacitor c=0.00227044f \
 //x=65.12 //y=2.08 //x2=66.23 //y2=4.54
cc_4187 ( N_noxref_20_c_6775_p N_noxref_21_c_6970_n ) capacitor c=0.00155256f \
 //x=65.755 //y=4.795 //x2=66.23 //y2=4.54
cc_4188 ( N_noxref_20_c_6639_n N_noxref_21_c_6970_n ) capacitor c=0.00180548f \
 //x=65.465 //y=4.795 //x2=66.23 //y2=4.54
cc_4189 ( N_noxref_20_c_6593_n N_noxref_21_c_6944_n ) capacitor c=0.00402215f \
 //x=65.005 //y=3.7 //x2=66.23 //y2=2.08
cc_4190 ( N_noxref_20_c_6597_n N_noxref_21_c_6944_n ) capacitor c=0.0232321f \
 //x=68.705 //y=4.44 //x2=66.23 //y2=2.08
cc_4191 ( N_noxref_20_c_6602_n N_noxref_21_c_6944_n ) capacitor c=9.10428e-19 \
 //x=65.235 //y=4.44 //x2=66.23 //y2=2.08
cc_4192 ( N_noxref_20_c_6563_n N_noxref_21_c_6944_n ) capacitor c=7.58505e-19 \
 //x=63.64 //y=3.7 //x2=66.23 //y2=2.08
cc_4193 ( N_noxref_20_c_6564_n N_noxref_21_c_6944_n ) capacitor c=0.0458192f \
 //x=65.12 //y=2.08 //x2=66.23 //y2=2.08
cc_4194 ( N_noxref_20_c_6567_n N_noxref_21_c_6944_n ) capacitor c=0.00969589f \
 //x=68.82 //y=2.08 //x2=66.23 //y2=2.08
cc_4195 ( N_noxref_20_c_6588_n N_noxref_21_c_6944_n ) capacitor c=0.00207026f \
 //x=65.12 //y=2.08 //x2=66.23 //y2=2.08
cc_4196 ( N_noxref_20_M123_noxref_g N_noxref_21_M125_noxref_g ) capacitor \
 c=0.010584f //x=65.39 //y=6.025 //x2=66.27 //y2=6.025
cc_4197 ( N_noxref_20_M124_noxref_g N_noxref_21_M125_noxref_g ) capacitor \
 c=0.106414f //x=65.83 //y=6.025 //x2=66.27 //y2=6.025
cc_4198 ( N_noxref_20_M124_noxref_g N_noxref_21_M126_noxref_g ) capacitor \
 c=0.0102479f //x=65.83 //y=6.025 //x2=66.71 //y2=6.025
cc_4199 ( N_noxref_20_c_6569_n N_noxref_21_c_7186_n ) capacitor c=4.86506e-19 \
 //x=65.295 //y=0.865 //x2=66.265 //y2=0.905
cc_4200 ( N_noxref_20_c_6571_n N_noxref_21_c_7186_n ) capacitor c=0.00152104f \
 //x=65.295 //y=1.21 //x2=66.265 //y2=0.905
cc_4201 ( N_noxref_20_c_6576_n N_noxref_21_c_7186_n ) capacitor c=0.0151475f \
 //x=65.825 //y=0.865 //x2=66.265 //y2=0.905
cc_4202 ( N_noxref_20_c_6572_n N_noxref_21_c_7189_n ) capacitor c=0.00109982f \
 //x=65.295 //y=1.52 //x2=66.265 //y2=1.25
cc_4203 ( N_noxref_20_c_6578_n N_noxref_21_c_7189_n ) capacitor c=0.0111064f \
 //x=65.825 //y=1.21 //x2=66.265 //y2=1.25
cc_4204 ( N_noxref_20_c_6572_n N_noxref_21_c_7191_n ) capacitor c=0.00182948f \
 //x=65.295 //y=1.52 //x2=66.265 //y2=1.56
cc_4205 ( N_noxref_20_c_6573_n N_noxref_21_c_7191_n ) capacitor c=0.00662747f \
 //x=65.295 //y=1.915 //x2=66.265 //y2=1.56
cc_4206 ( N_noxref_20_c_6578_n N_noxref_21_c_7191_n ) capacitor c=0.00862358f \
 //x=65.825 //y=1.21 //x2=66.265 //y2=1.56
cc_4207 ( N_noxref_20_c_6597_n N_noxref_21_c_6986_n ) capacitor c=0.0069773f \
 //x=68.705 //y=4.44 //x2=66.635 //y2=4.795
cc_4208 ( N_noxref_20_c_6576_n N_noxref_21_c_7195_n ) capacitor c=0.00124846f \
 //x=65.825 //y=0.865 //x2=66.795 //y2=0.905
cc_4209 ( N_noxref_20_c_6578_n N_noxref_21_c_7196_n ) capacitor c=0.00168739f \
 //x=65.825 //y=1.21 //x2=66.795 //y2=1.25
cc_4210 ( N_noxref_20_c_6564_n N_noxref_21_c_6948_n ) capacitor c=0.00197072f \
 //x=65.12 //y=2.08 //x2=66.23 //y2=2.08
cc_4211 ( N_noxref_20_c_6588_n N_noxref_21_c_6948_n ) capacitor c=0.00836805f \
 //x=65.12 //y=2.08 //x2=66.23 //y2=2.08
cc_4212 ( N_noxref_20_c_6597_n N_noxref_21_c_6987_n ) capacitor c=0.0014023f \
 //x=68.705 //y=4.44 //x2=66.27 //y2=4.705
cc_4213 ( N_noxref_20_c_6564_n N_noxref_21_c_6987_n ) capacitor c=0.00228787f \
 //x=65.12 //y=2.08 //x2=66.27 //y2=4.705
cc_4214 ( N_noxref_20_c_6775_p N_noxref_21_c_6987_n ) capacitor c=0.0201611f \
 //x=65.755 //y=4.795 //x2=66.27 //y2=4.705
cc_4215 ( N_noxref_20_c_6639_n N_noxref_21_c_6987_n ) capacitor c=0.00447195f \
 //x=65.465 //y=4.795 //x2=66.27 //y2=4.705
cc_4216 ( N_noxref_20_c_6597_n N_noxref_22_c_7406_n ) capacitor c=0.0856654f \
 //x=68.705 //y=4.44 //x2=68.375 //y2=5.21
cc_4217 ( N_noxref_20_M127_noxref_g N_noxref_22_c_7406_n ) capacitor \
 c=0.00503498f //x=68.71 //y=6.025 //x2=68.375 //y2=5.21
cc_4218 ( N_noxref_20_c_6597_n N_noxref_22_c_7412_n ) capacitor c=0.0130311f \
 //x=68.705 //y=4.44 //x2=66.605 //y2=5.21
cc_4219 ( N_noxref_20_c_6597_n N_noxref_22_c_7417_n ) capacitor c=0.00145992f \
 //x=68.705 //y=4.44 //x2=66.405 //y2=5.21
cc_4220 ( N_noxref_20_M124_noxref_g N_noxref_22_c_7417_n ) capacitor \
 c=0.0169795f //x=65.83 //y=6.025 //x2=66.405 //y2=5.21
cc_4221 ( N_noxref_20_c_6597_n N_noxref_22_c_7421_n ) capacitor c=0.0197096f \
 //x=68.705 //y=4.44 //x2=65.695 //y2=5.21
cc_4222 ( N_noxref_20_M123_noxref_g N_noxref_22_c_7421_n ) capacitor \
 c=0.0172236f //x=65.39 //y=6.025 //x2=65.695 //y2=5.21
cc_4223 ( N_noxref_20_c_6775_p N_noxref_22_c_7421_n ) capacitor c=0.00405363f \
 //x=65.755 //y=4.795 //x2=65.695 //y2=5.21
cc_4224 ( N_noxref_20_c_6597_n N_noxref_22_c_7423_n ) capacitor c=0.00467548f \
 //x=68.705 //y=4.44 //x2=66.49 //y2=5.295
cc_4225 ( N_noxref_20_c_6597_n N_noxref_22_c_7426_n ) capacitor c=0.00439121f \
 //x=68.705 //y=4.44 //x2=68.49 //y2=5.21
cc_4226 ( N_noxref_20_M127_noxref_g N_noxref_22_c_7426_n ) capacitor \
 c=0.0481665f //x=68.71 //y=6.025 //x2=68.49 //y2=5.21
cc_4227 ( N_noxref_20_c_6597_n N_noxref_22_c_7452_n ) capacitor c=0.00249667f \
 //x=68.705 //y=4.44 //x2=69.285 //y2=6.91
cc_4228 ( N_noxref_20_c_6567_n N_noxref_22_c_7452_n ) capacitor c=8.81369e-19 \
 //x=68.82 //y=2.08 //x2=69.285 //y2=6.91
cc_4229 ( N_noxref_20_M127_noxref_g N_noxref_22_c_7452_n ) capacitor \
 c=0.0163949f //x=68.71 //y=6.025 //x2=69.285 //y2=6.91
cc_4230 ( N_noxref_20_M128_noxref_g N_noxref_22_c_7452_n ) capacitor \
 c=0.0150104f //x=69.15 //y=6.025 //x2=69.285 //y2=6.91
cc_4231 ( N_noxref_20_M124_noxref_g N_noxref_22_M123_noxref_d ) capacitor \
 c=0.0169879f //x=65.83 //y=6.025 //x2=65.465 //y2=5.025
cc_4232 ( N_noxref_20_M128_noxref_g N_noxref_22_M128_noxref_d ) capacitor \
 c=0.0130327f //x=69.15 //y=6.025 //x2=69.225 //y2=5.025
cc_4233 ( N_noxref_20_c_6592_n N_noxref_23_c_7498_n ) capacitor c=0.164827f \
 //x=63.525 //y=3.7 //x2=70.185 //y2=2.96
cc_4234 ( N_noxref_20_c_6653_n N_noxref_23_c_7498_n ) capacitor c=0.0133752f \
 //x=59.685 //y=3.7 //x2=70.185 //y2=2.96
cc_4235 ( N_noxref_20_c_6593_n N_noxref_23_c_7498_n ) capacitor c=0.0706939f \
 //x=65.005 //y=3.7 //x2=70.185 //y2=2.96
cc_4236 ( N_noxref_20_c_6595_n N_noxref_23_c_7498_n ) capacitor c=0.0120929f \
 //x=63.755 //y=3.7 //x2=70.185 //y2=2.96
cc_4237 ( N_noxref_20_c_6597_n N_noxref_23_c_7498_n ) capacitor c=0.0280807f \
 //x=68.705 //y=4.44 //x2=70.185 //y2=2.96
cc_4238 ( N_noxref_20_c_6602_n N_noxref_23_c_7498_n ) capacitor c=3.57796e-19 \
 //x=65.235 //y=4.44 //x2=70.185 //y2=2.96
cc_4239 ( N_noxref_20_c_6560_n N_noxref_23_c_7498_n ) capacitor c=0.0219022f \
 //x=59.57 //y=2.08 //x2=70.185 //y2=2.96
cc_4240 ( N_noxref_20_c_6563_n N_noxref_23_c_7498_n ) capacitor c=0.0235216f \
 //x=63.64 //y=3.7 //x2=70.185 //y2=2.96
cc_4241 ( N_noxref_20_c_6564_n N_noxref_23_c_7498_n ) capacitor c=0.0244953f \
 //x=65.12 //y=2.08 //x2=70.185 //y2=2.96
cc_4242 ( N_noxref_20_c_6567_n N_noxref_23_c_7498_n ) capacitor c=0.0289771f \
 //x=68.82 //y=2.08 //x2=70.185 //y2=2.96
cc_4243 ( N_noxref_20_c_6582_n N_noxref_23_c_7498_n ) capacitor c=0.00383621f \
 //x=68.625 //y=1.915 //x2=70.185 //y2=2.96
cc_4244 ( N_noxref_20_c_6567_n N_noxref_23_c_7514_n ) capacitor c=0.00557744f \
 //x=68.82 //y=2.08 //x2=70.415 //y2=2.08
cc_4245 ( N_noxref_20_c_6597_n N_noxref_23_c_7519_n ) capacitor c=0.00408068f \
 //x=68.705 //y=4.44 //x2=70.3 //y2=2.08
cc_4246 ( N_noxref_20_c_6567_n N_noxref_23_c_7519_n ) capacitor c=0.0343626f \
 //x=68.82 //y=2.08 //x2=70.3 //y2=2.08
cc_4247 ( N_noxref_20_c_6582_n N_noxref_23_c_7519_n ) capacitor c=2.35599e-19 \
 //x=68.625 //y=1.915 //x2=70.3 //y2=2.08
cc_4248 ( N_noxref_20_c_6641_n N_noxref_23_c_7519_n ) capacitor c=2.35599e-19 \
 //x=68.82 //y=4.705 //x2=70.3 //y2=2.08
cc_4249 ( N_noxref_20_c_6567_n N_noxref_23_c_7521_n ) capacitor c=5.76627e-19 \
 //x=68.82 //y=2.08 //x2=71.78 //y2=2.08
cc_4250 ( N_noxref_20_M127_noxref_g N_noxref_23_M129_noxref_g ) capacitor \
 c=0.009459f //x=68.71 //y=6.025 //x2=69.59 //y2=6.025
cc_4251 ( N_noxref_20_M128_noxref_g N_noxref_23_M129_noxref_g ) capacitor \
 c=0.0626756f //x=69.15 //y=6.025 //x2=69.59 //y2=6.025
cc_4252 ( N_noxref_20_M128_noxref_g N_noxref_23_M130_noxref_g ) capacitor \
 c=0.00899012f //x=69.15 //y=6.025 //x2=70.03 //y2=6.025
cc_4253 ( N_noxref_20_c_6579_n N_noxref_23_c_7789_n ) capacitor c=4.86506e-19 \
 //x=68.625 //y=0.865 //x2=69.595 //y2=0.905
cc_4254 ( N_noxref_20_c_6581_n N_noxref_23_c_7789_n ) capacitor c=0.00101233f \
 //x=68.625 //y=1.21 //x2=69.595 //y2=0.905
cc_4255 ( N_noxref_20_c_6585_n N_noxref_23_c_7789_n ) capacitor c=0.0168844f \
 //x=69.155 //y=0.865 //x2=69.595 //y2=0.905
cc_4256 ( N_noxref_20_c_6844_p N_noxref_23_c_7792_n ) capacitor c=7.88071e-19 \
 //x=68.625 //y=1.52 //x2=69.595 //y2=1.25
cc_4257 ( N_noxref_20_c_6587_n N_noxref_23_c_7792_n ) capacitor c=0.0168218f \
 //x=69.155 //y=1.21 //x2=69.595 //y2=1.25
cc_4258 ( N_noxref_20_c_6567_n N_noxref_23_c_7794_n ) capacitor c=9.39431e-19 \
 //x=68.82 //y=2.08 //x2=69.665 //y2=4.795
cc_4259 ( N_noxref_20_c_6641_n N_noxref_23_c_7794_n ) capacitor c=0.0634092f \
 //x=68.82 //y=4.705 //x2=69.665 //y2=4.795
cc_4260 ( N_noxref_20_c_6567_n N_noxref_23_c_7565_n ) capacitor c=2.35599e-19 \
 //x=68.82 //y=2.08 //x2=70.03 //y2=4.87
cc_4261 ( N_noxref_20_c_6641_n N_noxref_23_c_7565_n ) capacitor c=5.35364e-19 \
 //x=68.82 //y=4.705 //x2=70.03 //y2=4.87
cc_4262 ( N_noxref_20_c_6585_n N_noxref_23_c_7798_n ) capacitor c=0.00124821f \
 //x=69.155 //y=0.865 //x2=70.125 //y2=0.905
cc_4263 ( N_noxref_20_c_6587_n N_noxref_23_c_7799_n ) capacitor c=8.19575e-19 \
 //x=69.155 //y=1.21 //x2=70.125 //y2=1.25
cc_4264 ( N_noxref_20_c_6587_n N_noxref_23_c_7800_n ) capacitor c=3.60397e-19 \
 //x=69.155 //y=1.21 //x2=70.125 //y2=1.56
cc_4265 ( N_noxref_20_c_6582_n N_noxref_23_c_7522_n ) capacitor c=4.61972e-19 \
 //x=68.625 //y=1.915 //x2=70.125 //y2=1.915
cc_4266 ( N_noxref_20_M128_noxref_g N_noxref_24_c_7971_n ) capacitor \
 c=0.0179287f //x=69.15 //y=6.025 //x2=69.725 //y2=5.21
cc_4267 ( N_noxref_20_c_6597_n N_noxref_24_c_7962_n ) capacitor c=0.0021588f \
 //x=68.705 //y=4.44 //x2=69.015 //y2=5.21
cc_4268 ( N_noxref_20_c_6567_n N_noxref_24_c_7962_n ) capacitor c=0.0056513f \
 //x=68.82 //y=2.08 //x2=69.015 //y2=5.21
cc_4269 ( N_noxref_20_M127_noxref_g N_noxref_24_c_7962_n ) capacitor \
 c=0.0132827f //x=68.71 //y=6.025 //x2=69.015 //y2=5.21
cc_4270 ( N_noxref_20_c_6641_n N_noxref_24_c_7962_n ) capacitor c=0.00554802f \
 //x=68.82 //y=4.705 //x2=69.015 //y2=5.21
cc_4271 ( N_noxref_20_M128_noxref_g N_noxref_24_M127_noxref_d ) capacitor \
 c=0.0130327f //x=69.15 //y=6.025 //x2=68.785 //y2=5.025
cc_4272 ( N_noxref_20_c_6581_n N_QN_c_8045_n ) capacitor c=0.00500281f \
 //x=68.625 //y=1.21 //x2=69.745 //y2=1.18
cc_4273 ( N_noxref_20_c_6844_p N_QN_c_8045_n ) capacitor c=0.00342096f \
 //x=68.625 //y=1.52 //x2=69.745 //y2=1.18
cc_4274 ( N_noxref_20_c_6583_n N_QN_c_8045_n ) capacitor c=4.02408e-19 //x=69 \
 //y=0.71 //x2=69.745 //y2=1.18
cc_4275 ( N_noxref_20_c_6584_n N_QN_c_8045_n ) capacitor c=0.0032199f //x=69 \
 //y=1.365 //x2=69.745 //y2=1.18
cc_4276 ( N_noxref_20_c_6587_n N_QN_c_8045_n ) capacitor c=0.00735559f \
 //x=69.155 //y=1.21 //x2=69.745 //y2=1.18
cc_4277 ( N_noxref_20_c_6668_n N_noxref_45_c_9211_n ) capacitor c=0.00623646f \
 //x=59.605 //y=1.56 //x2=59.385 //y2=1.495
cc_4278 ( N_noxref_20_c_6673_n N_noxref_45_c_9211_n ) capacitor c=0.00173579f \
 //x=59.57 //y=2.08 //x2=59.385 //y2=1.495
cc_4279 ( N_noxref_20_c_6560_n N_noxref_45_c_9212_n ) capacitor c=0.00156605f \
 //x=59.57 //y=2.08 //x2=60.27 //y2=0.53
cc_4280 ( N_noxref_20_c_6663_n N_noxref_45_c_9212_n ) capacitor c=0.0188655f \
 //x=59.605 //y=0.905 //x2=60.27 //y2=0.53
cc_4281 ( N_noxref_20_c_6671_n N_noxref_45_c_9212_n ) capacitor c=0.00656458f \
 //x=60.135 //y=0.905 //x2=60.27 //y2=0.53
cc_4282 ( N_noxref_20_c_6673_n N_noxref_45_c_9212_n ) capacitor c=2.1838e-19 \
 //x=59.57 //y=2.08 //x2=60.27 //y2=0.53
cc_4283 ( N_noxref_20_c_6663_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.00623646f //x=59.605 //y=0.905 //x2=58.28 //y2=0.365
cc_4284 ( N_noxref_20_c_6671_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.0143002f //x=60.135 //y=0.905 //x2=58.28 //y2=0.365
cc_4285 ( N_noxref_20_c_6672_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.00290153f //x=60.135 //y=1.25 //x2=58.28 //y2=0.365
cc_4286 ( N_noxref_20_c_6762_p N_noxref_46_c_9275_n ) capacitor c=3.15806e-19 \
 //x=63.285 //y=1.655 //x2=61.745 //y2=1.495
cc_4287 ( N_noxref_20_c_6762_p N_noxref_46_c_9263_n ) capacitor c=0.0203424f \
 //x=63.285 //y=1.655 //x2=62.715 //y2=1.495
cc_4288 ( N_noxref_20_c_6562_n N_noxref_46_c_9264_n ) capacitor c=0.00457164f \
 //x=63.555 //y=1.655 //x2=63.6 //y2=0.53
cc_4289 ( N_noxref_20_M38_noxref_d N_noxref_46_c_9264_n ) capacitor \
 c=0.0115831f //x=63.01 //y=0.905 //x2=63.6 //y2=0.53
cc_4290 ( N_noxref_20_c_6562_n N_noxref_46_M37_noxref_s ) capacitor \
 c=0.013435f //x=63.555 //y=1.655 //x2=61.61 //y2=0.365
cc_4291 ( N_noxref_20_M38_noxref_d N_noxref_46_M37_noxref_s ) capacitor \
 c=0.0439333f //x=63.01 //y=0.905 //x2=61.61 //y2=0.365
cc_4292 ( N_noxref_20_c_6562_n N_noxref_47_c_9327_n ) capacitor c=3.22188e-19 \
 //x=63.555 //y=1.655 //x2=65.075 //y2=1.495
cc_4293 ( N_noxref_20_c_6564_n N_noxref_47_c_9327_n ) capacitor c=0.015296f \
 //x=65.12 //y=2.08 //x2=65.075 //y2=1.495
cc_4294 ( N_noxref_20_c_6573_n N_noxref_47_c_9327_n ) capacitor c=0.0034165f \
 //x=65.295 //y=1.915 //x2=65.075 //y2=1.495
cc_4295 ( N_noxref_20_c_6588_n N_noxref_47_c_9327_n ) capacitor c=0.00780881f \
 //x=65.12 //y=2.08 //x2=65.075 //y2=1.495
cc_4296 ( N_noxref_20_c_6564_n N_noxref_47_c_9308_n ) capacitor c=0.00497226f \
 //x=65.12 //y=2.08 //x2=65.96 //y2=1.58
cc_4297 ( N_noxref_20_c_6572_n N_noxref_47_c_9308_n ) capacitor c=0.00700766f \
 //x=65.295 //y=1.52 //x2=65.96 //y2=1.58
cc_4298 ( N_noxref_20_c_6573_n N_noxref_47_c_9308_n ) capacitor c=0.0121133f \
 //x=65.295 //y=1.915 //x2=65.96 //y2=1.58
cc_4299 ( N_noxref_20_c_6575_n N_noxref_47_c_9308_n ) capacitor c=0.0103505f \
 //x=65.67 //y=1.365 //x2=65.96 //y2=1.58
cc_4300 ( N_noxref_20_c_6578_n N_noxref_47_c_9308_n ) capacitor c=0.00339872f \
 //x=65.825 //y=1.21 //x2=65.96 //y2=1.58
cc_4301 ( N_noxref_20_c_6588_n N_noxref_47_c_9308_n ) capacitor c=0.00324269f \
 //x=65.12 //y=2.08 //x2=65.96 //y2=1.58
cc_4302 ( N_noxref_20_c_6573_n N_noxref_47_c_9315_n ) capacitor c=6.71402e-19 \
 //x=65.295 //y=1.915 //x2=66.045 //y2=1.495
cc_4303 ( N_noxref_20_c_6569_n N_noxref_47_M39_noxref_s ) capacitor \
 c=0.0326001f //x=65.295 //y=0.865 //x2=64.94 //y2=0.365
cc_4304 ( N_noxref_20_c_6572_n N_noxref_47_M39_noxref_s ) capacitor \
 c=0.00110192f //x=65.295 //y=1.52 //x2=64.94 //y2=0.365
cc_4305 ( N_noxref_20_c_6576_n N_noxref_47_M39_noxref_s ) capacitor \
 c=0.0120759f //x=65.825 //y=0.865 //x2=64.94 //y2=0.365
cc_4306 ( N_noxref_20_c_6582_n N_noxref_48_c_9384_n ) capacitor c=0.0034165f \
 //x=68.625 //y=1.915 //x2=68.405 //y2=1.495
cc_4307 ( N_noxref_20_c_6567_n N_noxref_48_c_9366_n ) capacitor c=0.011159f \
 //x=68.82 //y=2.08 //x2=69.29 //y2=1.58
cc_4308 ( N_noxref_20_c_6844_p N_noxref_48_c_9366_n ) capacitor c=0.00598984f \
 //x=68.625 //y=1.52 //x2=69.29 //y2=1.58
cc_4309 ( N_noxref_20_c_6582_n N_noxref_48_c_9366_n ) capacitor c=0.0197952f \
 //x=68.625 //y=1.915 //x2=69.29 //y2=1.58
cc_4310 ( N_noxref_20_c_6584_n N_noxref_48_c_9366_n ) capacitor c=0.00767729f \
 //x=69 //y=1.365 //x2=69.29 //y2=1.58
cc_4311 ( N_noxref_20_c_6587_n N_noxref_48_c_9366_n ) capacitor c=0.0059368f \
 //x=69.155 //y=1.21 //x2=69.29 //y2=1.58
cc_4312 ( N_noxref_20_c_6582_n N_noxref_48_c_9372_n ) capacitor c=0.00122123f \
 //x=68.625 //y=1.915 //x2=69.375 //y2=1.495
cc_4313 ( N_noxref_20_c_6579_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.0312776f //x=68.625 //y=0.865 //x2=68.27 //y2=0.365
cc_4314 ( N_noxref_20_c_6844_p N_noxref_48_M41_noxref_s ) capacitor \
 c=3.48408e-19 //x=68.625 //y=1.52 //x2=68.27 //y2=0.365
cc_4315 ( N_noxref_20_c_6585_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.0132463f //x=69.155 //y=0.865 //x2=68.27 //y2=0.365
cc_4316 ( N_noxref_21_c_6938_n N_noxref_22_c_7406_n ) capacitor c=0.00923886f \
 //x=72.775 //y=4.07 //x2=68.375 //y2=5.21
cc_4317 ( N_noxref_21_M126_noxref_g N_noxref_22_c_7406_n ) capacitor \
 c=0.0104371f //x=66.71 //y=6.025 //x2=68.375 //y2=5.21
cc_4318 ( N_noxref_21_c_6938_n N_noxref_22_c_7412_n ) capacitor c=0.00122833f \
 //x=72.775 //y=4.07 //x2=66.605 //y2=5.21
cc_4319 ( N_noxref_21_M125_noxref_g N_noxref_22_c_7412_n ) capacitor \
 c=0.0010118f //x=66.27 //y=6.025 //x2=66.605 //y2=5.21
cc_4320 ( N_noxref_21_M126_noxref_g N_noxref_22_c_7412_n ) capacitor \
 c=8.30848e-19 //x=66.71 //y=6.025 //x2=66.605 //y2=5.21
cc_4321 ( N_noxref_21_c_6970_n N_noxref_22_c_7417_n ) capacitor c=0.012748f \
 //x=66.23 //y=4.54 //x2=66.405 //y2=5.21
cc_4322 ( N_noxref_21_M125_noxref_g N_noxref_22_c_7417_n ) capacitor \
 c=0.0161605f //x=66.27 //y=6.025 //x2=66.405 //y2=5.21
cc_4323 ( N_noxref_21_c_6987_n N_noxref_22_c_7417_n ) capacitor c=0.00307538f \
 //x=66.27 //y=4.705 //x2=66.405 //y2=5.21
cc_4324 ( N_noxref_21_M125_noxref_g N_noxref_22_c_7423_n ) capacitor \
 c=0.00226657f //x=66.27 //y=6.025 //x2=66.49 //y2=5.295
cc_4325 ( N_noxref_21_M126_noxref_g N_noxref_22_c_7423_n ) capacitor \
 c=0.0197448f //x=66.71 //y=6.025 //x2=66.49 //y2=5.295
cc_4326 ( N_noxref_21_c_6986_n N_noxref_22_c_7423_n ) capacitor c=0.00458101f \
 //x=66.635 //y=4.795 //x2=66.49 //y2=5.295
cc_4327 ( N_noxref_21_M125_noxref_g N_noxref_22_M125_noxref_d ) capacitor \
 c=0.016914f //x=66.27 //y=6.025 //x2=66.345 //y2=5.025
cc_4328 ( N_noxref_21_c_6904_n N_noxref_23_c_7498_n ) capacitor c=0.0293744f \
 //x=42.065 //y=2.22 //x2=70.185 //y2=2.96
cc_4329 ( N_noxref_21_c_6909_n N_noxref_23_c_7498_n ) capacitor c=9.7346e-19 \
 //x=38.225 //y=2.22 //x2=70.185 //y2=2.96
cc_4330 ( N_noxref_21_c_6911_n N_noxref_23_c_7498_n ) capacitor c=0.756304f \
 //x=66.115 //y=2.22 //x2=70.185 //y2=2.96
cc_4331 ( N_noxref_21_c_6935_n N_noxref_23_c_7498_n ) capacitor c=5.66322e-19 \
 //x=42.295 //y=2.22 //x2=70.185 //y2=2.96
cc_4332 ( N_noxref_21_c_6938_n N_noxref_23_c_7498_n ) capacitor c=0.123798f \
 //x=72.775 //y=4.07 //x2=70.185 //y2=2.96
cc_4333 ( N_noxref_21_c_6956_n N_noxref_23_c_7498_n ) capacitor c=0.00784775f \
 //x=66.345 //y=4.07 //x2=70.185 //y2=2.96
cc_4334 ( N_noxref_21_c_6939_n N_noxref_23_c_7498_n ) capacitor c=0.0208087f \
 //x=38.11 //y=2.08 //x2=70.185 //y2=2.96
cc_4335 ( N_noxref_21_c_6942_n N_noxref_23_c_7498_n ) capacitor c=0.0235867f \
 //x=42.18 //y=2.22 //x2=70.185 //y2=2.96
cc_4336 ( N_noxref_21_c_6944_n N_noxref_23_c_7498_n ) capacitor c=0.0264768f \
 //x=66.23 //y=2.08 //x2=70.185 //y2=2.96
cc_4337 ( N_noxref_21_c_6938_n N_noxref_23_c_7513_n ) capacitor c=0.0234111f \
 //x=72.775 //y=4.07 //x2=71.665 //y2=2.08
cc_4338 ( N_noxref_21_c_6946_n N_noxref_23_c_7513_n ) capacitor c=0.00668632f \
 //x=72.89 //y=2.08 //x2=71.665 //y2=2.08
cc_4339 ( N_noxref_21_c_7226_p N_noxref_23_c_7513_n ) capacitor c=0.00319611f \
 //x=72.89 //y=2.08 //x2=71.665 //y2=2.08
cc_4340 ( N_noxref_21_c_6911_n N_noxref_23_c_7514_n ) capacitor c=0.00135454f \
 //x=66.115 //y=2.22 //x2=70.415 //y2=2.08
cc_4341 ( N_noxref_21_c_6938_n N_noxref_23_c_7519_n ) capacitor c=0.0261405f \
 //x=72.775 //y=4.07 //x2=70.3 //y2=2.08
cc_4342 ( N_noxref_21_c_6946_n N_noxref_23_c_7519_n ) capacitor c=7.56813e-19 \
 //x=72.89 //y=2.08 //x2=70.3 //y2=2.08
cc_4343 ( N_noxref_21_c_6938_n N_noxref_23_c_7521_n ) capacitor c=0.0285749f \
 //x=72.775 //y=4.07 //x2=71.78 //y2=2.08
cc_4344 ( N_noxref_21_c_6946_n N_noxref_23_c_7521_n ) capacitor c=0.0538261f \
 //x=72.89 //y=2.08 //x2=71.78 //y2=2.08
cc_4345 ( N_noxref_21_c_7226_p N_noxref_23_c_7521_n ) capacitor c=0.00207994f \
 //x=72.89 //y=2.08 //x2=71.78 //y2=2.08
cc_4346 ( N_noxref_21_c_7233_p N_noxref_23_c_7521_n ) capacitor c=0.00196222f \
 //x=72.91 //y=4.705 //x2=71.78 //y2=2.08
cc_4347 ( N_noxref_21_M133_noxref_g N_noxref_23_M131_noxref_g ) capacitor \
 c=0.00932631f //x=72.93 //y=6.025 //x2=72.05 //y2=6.025
cc_4348 ( N_noxref_21_M133_noxref_g N_noxref_23_M132_noxref_g ) capacitor \
 c=0.110179f //x=72.93 //y=6.025 //x2=72.49 //y2=6.025
cc_4349 ( N_noxref_21_M134_noxref_g N_noxref_23_M132_noxref_g ) capacitor \
 c=0.00876656f //x=73.37 //y=6.025 //x2=72.49 //y2=6.025
cc_4350 ( N_noxref_21_c_6938_n N_noxref_23_c_7794_n ) capacitor c=0.00791694f \
 //x=72.775 //y=4.07 //x2=69.665 //y2=4.795
cc_4351 ( N_noxref_21_c_6938_n N_noxref_23_c_7565_n ) capacitor c=0.0014567f \
 //x=72.775 //y=4.07 //x2=70.03 //y2=4.87
cc_4352 ( N_noxref_21_c_7239_p N_noxref_23_c_7523_n ) capacitor c=4.86506e-19 \
 //x=72.925 //y=0.905 //x2=71.955 //y2=0.865
cc_4353 ( N_noxref_21_c_7239_p N_noxref_23_c_7525_n ) capacitor c=0.00101233f \
 //x=72.925 //y=0.905 //x2=71.955 //y2=1.21
cc_4354 ( N_noxref_21_c_7241_p N_noxref_23_c_7828_n ) capacitor c=0.00257836f \
 //x=72.925 //y=1.56 //x2=71.955 //y2=1.52
cc_4355 ( N_noxref_21_c_7241_p N_noxref_23_c_7526_n ) capacitor c=0.00662747f \
 //x=72.925 //y=1.56 //x2=71.955 //y2=1.915
cc_4356 ( N_noxref_21_c_7243_p N_noxref_23_c_7830_n ) capacitor c=0.00168516f \
 //x=72.91 //y=4.705 //x2=72.415 //y2=4.795
cc_4357 ( N_noxref_21_c_7233_p N_noxref_23_c_7830_n ) capacitor c=0.0225854f \
 //x=72.91 //y=4.705 //x2=72.415 //y2=4.795
cc_4358 ( N_noxref_21_c_6938_n N_noxref_23_c_7566_n ) capacitor c=0.0117386f \
 //x=72.775 //y=4.07 //x2=72.125 //y2=4.795
cc_4359 ( N_noxref_21_c_7243_p N_noxref_23_c_7566_n ) capacitor c=0.00143876f \
 //x=72.91 //y=4.705 //x2=72.125 //y2=4.795
cc_4360 ( N_noxref_21_c_7233_p N_noxref_23_c_7566_n ) capacitor c=0.00469886f \
 //x=72.91 //y=4.705 //x2=72.125 //y2=4.795
cc_4361 ( N_noxref_21_c_7239_p N_noxref_23_c_7529_n ) capacitor c=0.0161138f \
 //x=72.925 //y=0.905 //x2=72.485 //y2=0.865
cc_4362 ( N_noxref_21_c_7249_p N_noxref_23_c_7529_n ) capacitor c=0.00130607f \
 //x=73.455 //y=0.905 //x2=72.485 //y2=0.865
cc_4363 ( N_noxref_21_c_7250_p N_noxref_23_c_7531_n ) capacitor c=0.0120728f \
 //x=72.925 //y=1.255 //x2=72.485 //y2=1.21
cc_4364 ( N_noxref_21_c_7241_p N_noxref_23_c_7531_n ) capacitor c=0.00862358f \
 //x=72.925 //y=1.56 //x2=72.485 //y2=1.21
cc_4365 ( N_noxref_21_c_7252_p N_noxref_23_c_7531_n ) capacitor c=4.4593e-19 \
 //x=73.3 //y=1.405 //x2=72.485 //y2=1.21
cc_4366 ( N_noxref_21_c_7253_p N_noxref_23_c_7531_n ) capacitor c=0.00111855f \
 //x=73.455 //y=1.255 //x2=72.485 //y2=1.21
cc_4367 ( N_noxref_21_c_6946_n N_noxref_23_c_7532_n ) capacitor c=0.00218919f \
 //x=72.89 //y=2.08 //x2=71.78 //y2=2.08
cc_4368 ( N_noxref_21_c_7226_p N_noxref_23_c_7532_n ) capacitor c=0.00908973f \
 //x=72.89 //y=2.08 //x2=71.78 //y2=2.08
cc_4369 ( N_noxref_21_c_6938_n N_noxref_24_c_7956_n ) capacitor c=0.0535575f \
 //x=72.775 //y=4.07 //x2=71.715 //y2=5.21
cc_4370 ( N_noxref_21_c_6938_n N_noxref_24_c_7960_n ) capacitor c=0.008149f \
 //x=72.775 //y=4.07 //x2=69.925 //y2=5.21
cc_4371 ( N_noxref_21_c_6938_n N_noxref_24_c_7971_n ) capacitor c=3.2507e-19 \
 //x=72.775 //y=4.07 //x2=69.725 //y2=5.21
cc_4372 ( N_noxref_21_c_6938_n N_noxref_24_c_7962_n ) capacitor c=0.0181202f \
 //x=72.775 //y=4.07 //x2=69.015 //y2=5.21
cc_4373 ( N_noxref_21_c_6938_n N_noxref_24_c_7963_n ) capacitor c=0.00337443f \
 //x=72.775 //y=4.07 //x2=69.81 //y2=5.295
cc_4374 ( N_noxref_21_c_6938_n N_noxref_24_c_7964_n ) capacitor c=0.0011253f \
 //x=72.775 //y=4.07 //x2=71.83 //y2=5.21
cc_4375 ( N_noxref_21_c_6938_n N_noxref_24_c_7983_n ) capacitor c=0.00358031f \
 //x=72.775 //y=4.07 //x2=72.625 //y2=6.91
cc_4376 ( N_noxref_21_M133_noxref_g N_noxref_24_c_7984_n ) capacitor \
 c=0.0150104f //x=72.93 //y=6.025 //x2=73.505 //y2=6.91
cc_4377 ( N_noxref_21_M134_noxref_g N_noxref_24_c_7984_n ) capacitor \
 c=0.0163361f //x=73.37 //y=6.025 //x2=73.505 //y2=6.91
cc_4378 ( N_noxref_21_M133_noxref_g N_noxref_24_M132_noxref_d ) capacitor \
 c=0.0130327f //x=72.93 //y=6.025 //x2=72.565 //y2=5.025
cc_4379 ( N_noxref_21_M134_noxref_g N_noxref_24_M134_noxref_d ) capacitor \
 c=0.0351101f //x=73.37 //y=6.025 //x2=73.445 //y2=5.025
cc_4380 ( N_noxref_21_c_6938_n N_QN_c_8045_n ) capacitor c=0.00322521f \
 //x=72.775 //y=4.07 //x2=69.745 //y2=1.18
cc_4381 ( N_noxref_21_c_7195_n N_QN_c_8045_n ) capacitor c=4.67724e-19 \
 //x=66.795 //y=0.905 //x2=69.745 //y2=1.18
cc_4382 ( N_noxref_21_c_7196_n N_QN_c_8045_n ) capacitor c=0.00732681f \
 //x=66.795 //y=1.25 //x2=69.745 //y2=1.18
cc_4383 ( N_noxref_21_c_6938_n N_QN_c_8052_n ) capacitor c=4.20225e-19 \
 //x=72.775 //y=4.07 //x2=66.645 //y2=1.18
cc_4384 ( N_noxref_21_c_7186_n N_QN_c_8052_n ) capacitor c=3.66947e-19 \
 //x=66.265 //y=0.905 //x2=66.645 //y2=1.18
cc_4385 ( N_noxref_21_c_7189_n N_QN_c_8052_n ) capacitor c=0.00353233f \
 //x=66.265 //y=1.25 //x2=66.645 //y2=1.18
cc_4386 ( N_noxref_21_c_7191_n N_QN_c_8052_n ) capacitor c=0.00289074f \
 //x=66.265 //y=1.56 //x2=66.645 //y2=1.18
cc_4387 ( N_noxref_21_c_7274_p N_QN_c_8052_n ) capacitor c=4.06815e-19 \
 //x=66.64 //y=0.75 //x2=66.645 //y2=1.18
cc_4388 ( N_noxref_21_c_7275_p N_QN_c_8052_n ) capacitor c=7.42023e-19 \
 //x=66.64 //y=1.405 //x2=66.645 //y2=1.18
cc_4389 ( N_noxref_21_c_7196_n N_QN_c_8052_n ) capacitor c=0.00133904f \
 //x=66.795 //y=1.25 //x2=66.645 //y2=1.18
cc_4390 ( N_noxref_21_c_6938_n N_QN_c_8053_n ) capacitor c=0.0113709f \
 //x=72.775 //y=4.07 //x2=73.075 //y2=1.18
cc_4391 ( N_noxref_21_c_6946_n N_QN_c_8053_n ) capacitor c=0.00449159f \
 //x=72.89 //y=2.08 //x2=73.075 //y2=1.18
cc_4392 ( N_noxref_21_c_7239_p N_QN_c_8053_n ) capacitor c=6.33948e-19 \
 //x=72.925 //y=0.905 //x2=73.075 //y2=1.18
cc_4393 ( N_noxref_21_c_7250_p N_QN_c_8053_n ) capacitor c=0.0043333f \
 //x=72.925 //y=1.255 //x2=73.075 //y2=1.18
cc_4394 ( N_noxref_21_c_7241_p N_QN_c_8053_n ) capacitor c=0.0040799f \
 //x=72.925 //y=1.56 //x2=73.075 //y2=1.18
cc_4395 ( N_noxref_21_c_7282_p N_QN_c_8053_n ) capacitor c=4.52813e-19 \
 //x=73.3 //y=0.75 //x2=73.075 //y2=1.18
cc_4396 ( N_noxref_21_c_7252_p N_QN_c_8053_n ) capacitor c=0.00296491f \
 //x=73.3 //y=1.405 //x2=73.075 //y2=1.18
cc_4397 ( N_noxref_21_c_7249_p N_QN_c_8053_n ) capacitor c=2.65983e-19 \
 //x=73.455 //y=0.905 //x2=73.075 //y2=1.18
cc_4398 ( N_noxref_21_c_7253_p N_QN_c_8053_n ) capacitor c=0.00362989f \
 //x=73.455 //y=1.255 //x2=73.075 //y2=1.18
cc_4399 ( N_noxref_21_c_7226_p N_QN_c_8053_n ) capacitor c=5.89141e-19 \
 //x=72.89 //y=2.08 //x2=73.075 //y2=1.18
cc_4400 ( N_noxref_21_c_6938_n N_QN_c_8059_n ) capacitor c=3.74512e-19 \
 //x=72.775 //y=4.07 //x2=69.975 //y2=1.18
cc_4401 ( N_noxref_21_c_6938_n QN ) capacitor c=0.00642908f //x=72.775 \
 //y=4.07 //x2=73.63 //y2=2.22
cc_4402 ( N_noxref_21_c_6946_n QN ) capacitor c=0.0816497f //x=72.89 //y=2.08 \
 //x2=73.63 //y2=2.22
cc_4403 ( N_noxref_21_c_7243_p QN ) capacitor c=0.00998395f //x=72.91 \
 //y=4.705 //x2=73.63 //y2=2.22
cc_4404 ( N_noxref_21_c_7291_p QN ) capacitor c=0.0143966f //x=73.295 \
 //y=4.795 //x2=73.63 //y2=2.22
cc_4405 ( N_noxref_21_c_7226_p QN ) capacitor c=0.00704374f //x=72.89 //y=2.08 \
 //x2=73.63 //y2=2.22
cc_4406 ( N_noxref_21_c_7293_p QN ) capacitor c=0.0033061f //x=72.89 //y=1.915 \
 //x2=73.63 //y2=2.22
cc_4407 ( N_noxref_21_c_7233_p QN ) capacitor c=0.00526987f //x=72.91 \
 //y=4.705 //x2=73.63 //y2=2.22
cc_4408 ( N_noxref_21_c_6938_n N_QN_c_8112_n ) capacitor c=0.00154966f \
 //x=72.775 //y=4.07 //x2=73.065 //y2=5.21
cc_4409 ( N_noxref_21_c_7243_p N_QN_c_8112_n ) capacitor c=0.0128151f \
 //x=72.91 //y=4.705 //x2=73.065 //y2=5.21
cc_4410 ( N_noxref_21_M133_noxref_g N_QN_c_8112_n ) capacitor c=0.0167296f \
 //x=72.93 //y=6.025 //x2=73.065 //y2=5.21
cc_4411 ( N_noxref_21_c_7233_p N_QN_c_8112_n ) capacitor c=0.00368327f \
 //x=72.91 //y=4.705 //x2=73.065 //y2=5.21
cc_4412 ( N_noxref_21_c_6938_n N_QN_c_8074_n ) capacitor c=0.0138451f \
 //x=72.775 //y=4.07 //x2=72.355 //y2=5.21
cc_4413 ( N_noxref_21_M134_noxref_g N_QN_c_8075_n ) capacitor c=0.0222938f \
 //x=73.37 //y=6.025 //x2=73.545 //y2=5.21
cc_4414 ( N_noxref_21_c_7252_p N_QN_c_8061_n ) capacitor c=0.00810194f \
 //x=73.3 //y=1.405 //x2=73.545 //y2=1.645
cc_4415 ( N_noxref_21_c_7293_p N_QN_c_8119_n ) capacitor c=0.00671029f \
 //x=72.89 //y=1.915 //x2=73.275 //y2=1.645
cc_4416 ( N_noxref_21_c_7291_p N_QN_c_8120_n ) capacitor c=0.00410596f \
 //x=73.295 //y=4.795 //x2=73.15 //y2=5.21
cc_4417 ( N_noxref_21_c_7186_n N_QN_M40_noxref_d ) capacitor c=0.00218556f \
 //x=66.265 //y=0.905 //x2=66.34 //y2=0.905
cc_4418 ( N_noxref_21_c_7189_n N_QN_M40_noxref_d ) capacitor c=0.00327871f \
 //x=66.265 //y=1.25 //x2=66.34 //y2=0.905
cc_4419 ( N_noxref_21_c_7191_n N_QN_M40_noxref_d ) capacitor c=0.00292542f \
 //x=66.265 //y=1.56 //x2=66.34 //y2=0.905
cc_4420 ( N_noxref_21_c_7274_p N_QN_M40_noxref_d ) capacitor c=0.00235569f \
 //x=66.64 //y=0.75 //x2=66.34 //y2=0.905
cc_4421 ( N_noxref_21_c_7275_p N_QN_M40_noxref_d ) capacitor c=0.00613695f \
 //x=66.64 //y=1.405 //x2=66.34 //y2=0.905
cc_4422 ( N_noxref_21_c_7195_n N_QN_M40_noxref_d ) capacitor c=0.00131413f \
 //x=66.795 //y=0.905 //x2=66.34 //y2=0.905
cc_4423 ( N_noxref_21_c_7196_n N_QN_M40_noxref_d ) capacitor c=0.00676348f \
 //x=66.795 //y=1.25 //x2=66.34 //y2=0.905
cc_4424 ( N_noxref_21_c_7239_p N_QN_M44_noxref_d ) capacitor c=0.00226395f \
 //x=72.925 //y=0.905 //x2=73 //y2=0.905
cc_4425 ( N_noxref_21_c_7250_p N_QN_M44_noxref_d ) capacitor c=0.004517f \
 //x=72.925 //y=1.255 //x2=73 //y2=0.905
cc_4426 ( N_noxref_21_c_7241_p N_QN_M44_noxref_d ) capacitor c=0.00655125f \
 //x=72.925 //y=1.56 //x2=73 //y2=0.905
cc_4427 ( N_noxref_21_c_7282_p N_QN_M44_noxref_d ) capacitor c=0.00241003f \
 //x=73.3 //y=0.75 //x2=73 //y2=0.905
cc_4428 ( N_noxref_21_c_7252_p N_QN_M44_noxref_d ) capacitor c=0.0159024f \
 //x=73.3 //y=1.405 //x2=73 //y2=0.905
cc_4429 ( N_noxref_21_c_7249_p N_QN_M44_noxref_d ) capacitor c=0.00132831f \
 //x=73.455 //y=0.905 //x2=73 //y2=0.905
cc_4430 ( N_noxref_21_c_7253_p N_QN_M44_noxref_d ) capacitor c=0.00330743f \
 //x=73.455 //y=1.255 //x2=73 //y2=0.905
cc_4431 ( N_noxref_21_M133_noxref_g N_QN_M133_noxref_d ) capacitor \
 c=0.0130327f //x=72.93 //y=6.025 //x2=73.005 //y2=5.025
cc_4432 ( N_noxref_21_M134_noxref_g N_QN_M133_noxref_d ) capacitor \
 c=0.0136385f //x=73.37 //y=6.025 //x2=73.005 //y2=5.025
cc_4433 ( N_noxref_21_c_6909_n N_noxref_38_c_8844_n ) capacitor c=0.00185188f \
 //x=38.225 //y=2.22 //x2=37.925 //y2=1.495
cc_4434 ( N_noxref_21_c_7014_n N_noxref_38_c_8844_n ) capacitor c=0.00623646f \
 //x=38.145 //y=1.56 //x2=37.925 //y2=1.495
cc_4435 ( N_noxref_21_c_7019_n N_noxref_38_c_8844_n ) capacitor c=0.00173568f \
 //x=38.11 //y=2.08 //x2=37.925 //y2=1.495
cc_4436 ( N_noxref_21_c_6904_n N_noxref_38_c_8845_n ) capacitor c=0.00123263f \
 //x=42.065 //y=2.22 //x2=38.81 //y2=0.53
cc_4437 ( N_noxref_21_c_6909_n N_noxref_38_c_8845_n ) capacitor c=5.55767e-19 \
 //x=38.225 //y=2.22 //x2=38.81 //y2=0.53
cc_4438 ( N_noxref_21_c_6939_n N_noxref_38_c_8845_n ) capacitor c=0.00156443f \
 //x=38.11 //y=2.08 //x2=38.81 //y2=0.53
cc_4439 ( N_noxref_21_c_7009_n N_noxref_38_c_8845_n ) capacitor c=0.0188655f \
 //x=38.145 //y=0.905 //x2=38.81 //y2=0.53
cc_4440 ( N_noxref_21_c_7017_n N_noxref_38_c_8845_n ) capacitor c=0.00656458f \
 //x=38.675 //y=0.905 //x2=38.81 //y2=0.53
cc_4441 ( N_noxref_21_c_7019_n N_noxref_38_c_8845_n ) capacitor c=2.1838e-19 \
 //x=38.11 //y=2.08 //x2=38.81 //y2=0.53
cc_4442 ( N_noxref_21_c_6904_n N_noxref_38_M22_noxref_s ) capacitor \
 c=0.00113237f //x=42.065 //y=2.22 //x2=36.82 //y2=0.365
cc_4443 ( N_noxref_21_c_7009_n N_noxref_38_M22_noxref_s ) capacitor \
 c=0.00623646f //x=38.145 //y=0.905 //x2=36.82 //y2=0.365
cc_4444 ( N_noxref_21_c_7017_n N_noxref_38_M22_noxref_s ) capacitor \
 c=0.0143002f //x=38.675 //y=0.905 //x2=36.82 //y2=0.365
cc_4445 ( N_noxref_21_c_7018_n N_noxref_38_M22_noxref_s ) capacitor \
 c=0.00290153f //x=38.675 //y=1.25 //x2=36.82 //y2=0.365
cc_4446 ( N_noxref_21_c_6904_n N_noxref_39_c_8910_n ) capacitor c=0.00635755f \
 //x=42.065 //y=2.22 //x2=40.285 //y2=1.495
cc_4447 ( N_noxref_21_c_7334_p N_noxref_39_c_8910_n ) capacitor c=3.15806e-19 \
 //x=41.825 //y=1.655 //x2=40.285 //y2=1.495
cc_4448 ( N_noxref_21_c_6904_n N_noxref_39_c_8891_n ) capacitor c=0.0223494f \
 //x=42.065 //y=2.22 //x2=41.17 //y2=1.58
cc_4449 ( N_noxref_21_c_6904_n N_noxref_39_c_8898_n ) capacitor c=0.00649228f \
 //x=42.065 //y=2.22 //x2=41.255 //y2=1.495
cc_4450 ( N_noxref_21_c_7334_p N_noxref_39_c_8898_n ) capacitor c=0.0203424f \
 //x=41.825 //y=1.655 //x2=41.255 //y2=1.495
cc_4451 ( N_noxref_21_c_6904_n N_noxref_39_c_8899_n ) capacitor c=0.00178534f \
 //x=42.065 //y=2.22 //x2=42.14 //y2=0.53
cc_4452 ( N_noxref_21_c_6941_n N_noxref_39_c_8899_n ) capacitor c=0.00457122f \
 //x=42.095 //y=1.655 //x2=42.14 //y2=0.53
cc_4453 ( N_noxref_21_M25_noxref_d N_noxref_39_c_8899_n ) capacitor \
 c=0.0115831f //x=41.55 //y=0.905 //x2=42.14 //y2=0.53
cc_4454 ( N_noxref_21_c_6911_n N_noxref_39_M24_noxref_s ) capacitor \
 c=3.68089e-19 //x=66.115 //y=2.22 //x2=40.15 //y2=0.365
cc_4455 ( N_noxref_21_c_6935_n N_noxref_39_M24_noxref_s ) capacitor \
 c=8.2308e-19 //x=42.295 //y=2.22 //x2=40.15 //y2=0.365
cc_4456 ( N_noxref_21_c_6941_n N_noxref_39_M24_noxref_s ) capacitor \
 c=0.0130338f //x=42.095 //y=1.655 //x2=40.15 //y2=0.365
cc_4457 ( N_noxref_21_c_6942_n N_noxref_39_M24_noxref_s ) capacitor \
 c=2.31582e-19 //x=42.18 //y=2.22 //x2=40.15 //y2=0.365
cc_4458 ( N_noxref_21_M25_noxref_d N_noxref_39_M24_noxref_s ) capacitor \
 c=0.043966f //x=41.55 //y=0.905 //x2=40.15 //y2=0.365
cc_4459 ( N_noxref_21_c_6911_n N_noxref_40_c_8970_n ) capacitor c=0.00642985f \
 //x=66.115 //y=2.22 //x2=43.51 //y2=1.505
cc_4460 ( N_noxref_21_c_6941_n N_noxref_40_c_8970_n ) capacitor c=4.08644e-19 \
 //x=42.095 //y=1.655 //x2=43.51 //y2=1.505
cc_4461 ( N_noxref_21_c_6911_n N_noxref_40_c_8945_n ) capacitor c=0.0225733f \
 //x=66.115 //y=2.22 //x2=44.395 //y2=1.59
cc_4462 ( N_noxref_21_c_6911_n N_noxref_40_c_8963_n ) capacitor c=0.0203655f \
 //x=66.115 //y=2.22 //x2=45.365 //y2=1.59
cc_4463 ( N_noxref_21_c_6911_n N_noxref_40_M26_noxref_s ) capacitor \
 c=0.012425f //x=66.115 //y=2.22 //x2=43.375 //y2=0.375
cc_4464 ( N_noxref_21_M25_noxref_d N_noxref_40_M26_noxref_s ) capacitor \
 c=2.53688e-19 //x=41.55 //y=0.905 //x2=43.375 //y2=0.375
cc_4465 ( N_noxref_21_c_6911_n N_noxref_41_c_8995_n ) capacitor c=0.00657782f \
 //x=66.115 //y=2.22 //x2=45.935 //y2=0.995
cc_4466 ( N_noxref_21_c_6911_n N_noxref_41_c_9000_n ) capacitor c=0.00147946f \
 //x=66.115 //y=2.22 //x2=46.905 //y2=0.54
cc_4467 ( N_noxref_21_c_6911_n N_noxref_41_M28_noxref_s ) capacitor \
 c=0.00642985f //x=66.115 //y=2.22 //x2=45.885 //y2=0.375
cc_4468 ( N_noxref_21_c_6911_n N_noxref_42_c_9076_n ) capacitor c=0.00635755f \
 //x=66.115 //y=2.22 //x2=48.425 //y2=1.495
cc_4469 ( N_noxref_21_c_6911_n N_noxref_42_c_9048_n ) capacitor c=0.0223494f \
 //x=66.115 //y=2.22 //x2=49.31 //y2=1.58
cc_4470 ( N_noxref_21_c_6911_n N_noxref_42_c_9055_n ) capacitor c=0.00649228f \
 //x=66.115 //y=2.22 //x2=49.395 //y2=1.495
cc_4471 ( N_noxref_21_c_6911_n N_noxref_42_c_9056_n ) capacitor c=0.00178534f \
 //x=66.115 //y=2.22 //x2=50.28 //y2=0.53
cc_4472 ( N_noxref_21_c_6911_n N_noxref_42_M29_noxref_s ) capacitor \
 c=0.00113237f //x=66.115 //y=2.22 //x2=48.29 //y2=0.365
cc_4473 ( N_noxref_21_c_6911_n N_noxref_43_c_9119_n ) capacitor c=0.00635755f \
 //x=66.115 //y=2.22 //x2=51.755 //y2=1.495
cc_4474 ( N_noxref_21_c_6911_n N_noxref_43_c_9100_n ) capacitor c=0.0223494f \
 //x=66.115 //y=2.22 //x2=52.64 //y2=1.58
cc_4475 ( N_noxref_21_c_6911_n N_noxref_43_c_9107_n ) capacitor c=0.00649228f \
 //x=66.115 //y=2.22 //x2=52.725 //y2=1.495
cc_4476 ( N_noxref_21_c_6911_n N_noxref_43_c_9108_n ) capacitor c=0.00178534f \
 //x=66.115 //y=2.22 //x2=53.61 //y2=0.53
cc_4477 ( N_noxref_21_c_6911_n N_noxref_43_M31_noxref_s ) capacitor \
 c=0.00113237f //x=66.115 //y=2.22 //x2=51.62 //y2=0.365
cc_4478 ( N_noxref_21_c_6911_n N_noxref_44_c_9171_n ) capacitor c=0.00635755f \
 //x=66.115 //y=2.22 //x2=55.085 //y2=1.495
cc_4479 ( N_noxref_21_c_6911_n N_noxref_44_c_9152_n ) capacitor c=0.0223494f \
 //x=66.115 //y=2.22 //x2=55.97 //y2=1.58
cc_4480 ( N_noxref_21_c_6911_n N_noxref_44_c_9159_n ) capacitor c=0.00649228f \
 //x=66.115 //y=2.22 //x2=56.055 //y2=1.495
cc_4481 ( N_noxref_21_c_6911_n N_noxref_44_c_9160_n ) capacitor c=0.00178534f \
 //x=66.115 //y=2.22 //x2=56.94 //y2=0.53
cc_4482 ( N_noxref_21_c_6911_n N_noxref_44_M33_noxref_s ) capacitor \
 c=0.00113237f //x=66.115 //y=2.22 //x2=54.95 //y2=0.365
cc_4483 ( N_noxref_21_c_6911_n N_noxref_45_c_9223_n ) capacitor c=0.00635755f \
 //x=66.115 //y=2.22 //x2=58.415 //y2=1.495
cc_4484 ( N_noxref_21_c_6911_n N_noxref_45_c_9204_n ) capacitor c=0.0223494f \
 //x=66.115 //y=2.22 //x2=59.3 //y2=1.58
cc_4485 ( N_noxref_21_c_6911_n N_noxref_45_c_9211_n ) capacitor c=0.00649228f \
 //x=66.115 //y=2.22 //x2=59.385 //y2=1.495
cc_4486 ( N_noxref_21_c_6911_n N_noxref_45_c_9212_n ) capacitor c=0.00178534f \
 //x=66.115 //y=2.22 //x2=60.27 //y2=0.53
cc_4487 ( N_noxref_21_c_6911_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.00113237f //x=66.115 //y=2.22 //x2=58.28 //y2=0.365
cc_4488 ( N_noxref_21_c_6911_n N_noxref_46_c_9275_n ) capacitor c=0.00635755f \
 //x=66.115 //y=2.22 //x2=61.745 //y2=1.495
cc_4489 ( N_noxref_21_c_6911_n N_noxref_46_c_9256_n ) capacitor c=0.0223494f \
 //x=66.115 //y=2.22 //x2=62.63 //y2=1.58
cc_4490 ( N_noxref_21_c_6911_n N_noxref_46_c_9263_n ) capacitor c=0.00649228f \
 //x=66.115 //y=2.22 //x2=62.715 //y2=1.495
cc_4491 ( N_noxref_21_c_6911_n N_noxref_46_c_9264_n ) capacitor c=0.00178534f \
 //x=66.115 //y=2.22 //x2=63.6 //y2=0.53
cc_4492 ( N_noxref_21_c_6911_n N_noxref_46_M37_noxref_s ) capacitor \
 c=0.00113237f //x=66.115 //y=2.22 //x2=61.61 //y2=0.365
cc_4493 ( N_noxref_21_c_6911_n N_noxref_47_c_9327_n ) capacitor c=0.0018561f \
 //x=66.115 //y=2.22 //x2=65.075 //y2=1.495
cc_4494 ( N_noxref_21_c_6911_n N_noxref_47_c_9308_n ) capacitor c=0.024432f \
 //x=66.115 //y=2.22 //x2=65.96 //y2=1.58
cc_4495 ( N_noxref_21_c_6911_n N_noxref_47_c_9315_n ) capacitor c=0.00650742f \
 //x=66.115 //y=2.22 //x2=66.045 //y2=1.495
cc_4496 ( N_noxref_21_c_7191_n N_noxref_47_c_9315_n ) capacitor c=0.00746306f \
 //x=66.265 //y=1.56 //x2=66.045 //y2=1.495
cc_4497 ( N_noxref_21_c_6948_n N_noxref_47_c_9315_n ) capacitor c=0.00173568f \
 //x=66.23 //y=2.08 //x2=66.045 //y2=1.495
cc_4498 ( N_noxref_21_c_6911_n N_noxref_47_c_9316_n ) capacitor c=0.00102746f \
 //x=66.115 //y=2.22 //x2=66.93 //y2=0.53
cc_4499 ( N_noxref_21_c_6944_n N_noxref_47_c_9316_n ) capacitor c=0.00156442f \
 //x=66.23 //y=2.08 //x2=66.93 //y2=0.53
cc_4500 ( N_noxref_21_c_7186_n N_noxref_47_c_9316_n ) capacitor c=0.0200006f \
 //x=66.265 //y=0.905 //x2=66.93 //y2=0.53
cc_4501 ( N_noxref_21_c_7195_n N_noxref_47_c_9316_n ) capacitor c=0.00825432f \
 //x=66.795 //y=0.905 //x2=66.93 //y2=0.53
cc_4502 ( N_noxref_21_c_6948_n N_noxref_47_c_9316_n ) capacitor c=2.1838e-19 \
 //x=66.23 //y=2.08 //x2=66.93 //y2=0.53
cc_4503 ( N_noxref_21_c_7186_n N_noxref_47_M39_noxref_s ) capacitor \
 c=0.00746306f //x=66.265 //y=0.905 //x2=64.94 //y2=0.365
cc_4504 ( N_noxref_21_c_7191_n N_noxref_47_M39_noxref_s ) capacitor \
 c=0.00213023f //x=66.265 //y=1.56 //x2=64.94 //y2=0.365
cc_4505 ( N_noxref_21_c_7195_n N_noxref_47_M39_noxref_s ) capacitor \
 c=0.0133026f //x=66.795 //y=0.905 //x2=64.94 //y2=0.365
cc_4506 ( N_noxref_21_c_7196_n N_noxref_47_M39_noxref_s ) capacitor \
 c=0.00793126f //x=66.795 //y=1.25 //x2=64.94 //y2=0.365
cc_4507 ( N_noxref_21_c_7394_p N_noxref_47_M39_noxref_s ) capacitor \
 c=0.00392195f //x=66.23 //y=1.915 //x2=64.94 //y2=0.365
cc_4508 ( N_noxref_21_c_6938_n N_noxref_49_c_9422_n ) capacitor c=0.00631223f \
 //x=72.775 //y=4.07 //x2=72.62 //y2=1.58
cc_4509 ( N_noxref_21_c_6938_n N_noxref_49_c_9428_n ) capacitor c=0.00108825f \
 //x=72.775 //y=4.07 //x2=72.705 //y2=1.495
cc_4510 ( N_noxref_21_c_7241_p N_noxref_49_c_9428_n ) capacitor c=0.00698471f \
 //x=72.925 //y=1.56 //x2=72.705 //y2=1.495
cc_4511 ( N_noxref_21_c_7226_p N_noxref_49_c_9428_n ) capacitor c=0.00171785f \
 //x=72.89 //y=2.08 //x2=72.705 //y2=1.495
cc_4512 ( N_noxref_21_c_6946_n N_noxref_49_c_9429_n ) capacitor c=0.00118117f \
 //x=72.89 //y=2.08 //x2=73.59 //y2=0.53
cc_4513 ( N_noxref_21_c_7239_p N_noxref_49_c_9429_n ) capacitor c=0.0191024f \
 //x=72.925 //y=0.905 //x2=73.59 //y2=0.53
cc_4514 ( N_noxref_21_c_7249_p N_noxref_49_c_9429_n ) capacitor c=0.00655165f \
 //x=73.455 //y=0.905 //x2=73.59 //y2=0.53
cc_4515 ( N_noxref_21_c_7226_p N_noxref_49_c_9429_n ) capacitor c=2.1838e-19 \
 //x=72.89 //y=2.08 //x2=73.59 //y2=0.53
cc_4516 ( N_noxref_21_c_7239_p N_noxref_49_M43_noxref_s ) capacitor \
 c=0.00698471f //x=72.925 //y=0.905 //x2=71.6 //y2=0.365
cc_4517 ( N_noxref_21_c_7252_p N_noxref_49_M43_noxref_s ) capacitor \
 c=0.00316186f //x=73.3 //y=1.405 //x2=71.6 //y2=0.365
cc_4518 ( N_noxref_21_c_7249_p N_noxref_49_M43_noxref_s ) capacitor \
 c=0.0142835f //x=73.455 //y=0.905 //x2=71.6 //y2=0.365
cc_4519 ( N_noxref_22_M130_noxref_d N_noxref_23_c_7519_n ) capacitor \
 c=0.00496677f //x=70.105 //y=5.025 //x2=70.3 //y2=2.08
cc_4520 ( N_noxref_22_c_7471_p N_noxref_23_M129_noxref_g ) capacitor \
 c=0.0150104f //x=70.165 //y=6.91 //x2=69.59 //y2=6.025
cc_4521 ( N_noxref_22_M128_noxref_d N_noxref_23_M129_noxref_g ) capacitor \
 c=0.0130327f //x=69.225 //y=5.025 //x2=69.59 //y2=6.025
cc_4522 ( N_noxref_22_c_7471_p N_noxref_23_M130_noxref_g ) capacitor \
 c=0.0155183f //x=70.165 //y=6.91 //x2=70.03 //y2=6.025
cc_4523 ( N_noxref_22_M130_noxref_d N_noxref_23_M130_noxref_g ) capacitor \
 c=0.0398886f //x=70.105 //y=5.025 //x2=70.03 //y2=6.025
cc_4524 ( N_noxref_22_M130_noxref_d N_noxref_23_c_7565_n ) capacitor \
 c=0.00411435f //x=70.105 //y=5.025 //x2=70.03 //y2=4.87
cc_4525 ( N_noxref_22_c_7471_p N_noxref_24_c_7956_n ) capacitor c=0.00546043f \
 //x=70.165 //y=6.91 //x2=71.715 //y2=5.21
cc_4526 ( N_noxref_22_M130_noxref_d N_noxref_24_c_7956_n ) capacitor \
 c=0.00675852f //x=70.105 //y=5.025 //x2=71.715 //y2=5.21
cc_4527 ( N_noxref_22_c_7406_n N_noxref_24_c_7960_n ) capacitor c=0.0086908f \
 //x=68.375 //y=5.21 //x2=69.925 //y2=5.21
cc_4528 ( N_noxref_22_c_7471_p N_noxref_24_c_7960_n ) capacitor c=9.39989e-19 \
 //x=70.165 //y=6.91 //x2=69.925 //y2=5.21
cc_4529 ( N_noxref_22_c_7452_n N_noxref_24_c_7971_n ) capacitor c=0.00102709f \
 //x=69.285 //y=6.91 //x2=69.725 //y2=5.21
cc_4530 ( N_noxref_22_c_7471_p N_noxref_24_c_7971_n ) capacitor c=9.89472e-19 \
 //x=70.165 //y=6.91 //x2=69.725 //y2=5.21
cc_4531 ( N_noxref_22_M128_noxref_d N_noxref_24_c_7971_n ) capacitor \
 c=0.0124612f //x=69.225 //y=5.025 //x2=69.725 //y2=5.21
cc_4532 ( N_noxref_22_c_7406_n N_noxref_24_c_7962_n ) capacitor c=0.00638395f \
 //x=68.375 //y=5.21 //x2=69.015 //y2=5.21
cc_4533 ( N_noxref_22_c_7426_n N_noxref_24_c_7962_n ) capacitor c=0.0682565f \
 //x=68.49 //y=5.21 //x2=69.015 //y2=5.21
cc_4534 ( N_noxref_22_c_7426_n N_noxref_24_c_7963_n ) capacitor c=9.46973e-19 \
 //x=68.49 //y=5.21 //x2=69.81 //y2=5.295
cc_4535 ( N_noxref_22_M130_noxref_d N_noxref_24_c_7964_n ) capacitor \
 c=0.001104f //x=70.105 //y=5.025 //x2=71.83 //y2=5.21
cc_4536 ( N_noxref_22_c_7471_p N_noxref_24_c_7966_n ) capacitor c=0.001104f \
 //x=70.165 //y=6.91 //x2=71.915 //y2=6.91
cc_4537 ( N_noxref_22_c_7406_n N_noxref_24_M127_noxref_d ) capacitor \
 c=4.76678e-19 //x=68.375 //y=5.21 //x2=68.785 //y2=5.025
cc_4538 ( N_noxref_22_c_7452_n N_noxref_24_M127_noxref_d ) capacitor \
 c=0.0115421f //x=69.285 //y=6.91 //x2=68.785 //y2=5.025
cc_4539 ( N_noxref_22_M128_noxref_d N_noxref_24_M127_noxref_d ) capacitor \
 c=0.0458293f //x=69.225 //y=5.025 //x2=68.785 //y2=5.025
cc_4540 ( N_noxref_22_M130_noxref_d N_noxref_24_M127_noxref_d ) capacitor \
 c=7.47391e-19 //x=70.105 //y=5.025 //x2=68.785 //y2=5.025
cc_4541 ( N_noxref_22_c_7426_n N_noxref_24_M129_noxref_d ) capacitor \
 c=9.55e-19 //x=68.49 //y=5.21 //x2=69.665 //y2=5.025
cc_4542 ( N_noxref_22_c_7471_p N_noxref_24_M129_noxref_d ) capacitor \
 c=0.0115693f //x=70.165 //y=6.91 //x2=69.665 //y2=5.025
cc_4543 ( N_noxref_22_M128_noxref_d N_noxref_24_M129_noxref_d ) capacitor \
 c=0.0458293f //x=69.225 //y=5.025 //x2=69.665 //y2=5.025
cc_4544 ( N_noxref_22_M130_noxref_d N_noxref_24_M129_noxref_d ) capacitor \
 c=0.0550393f //x=70.105 //y=5.025 //x2=69.665 //y2=5.025
cc_4545 ( N_noxref_22_c_7426_n N_noxref_48_c_9384_n ) capacitor c=0.00109479f \
 //x=68.49 //y=5.21 //x2=68.405 //y2=1.495
cc_4546 ( N_noxref_23_c_7498_n N_noxref_24_c_7956_n ) capacitor c=7.38711e-19 \
 //x=70.185 //y=2.96 //x2=71.715 //y2=5.21
cc_4547 ( N_noxref_23_c_7513_n N_noxref_24_c_7956_n ) capacitor c=5.48246e-19 \
 //x=71.665 //y=2.08 //x2=71.715 //y2=5.21
cc_4548 ( N_noxref_23_c_7519_n N_noxref_24_c_7956_n ) capacitor c=0.00419026f \
 //x=70.3 //y=2.08 //x2=71.715 //y2=5.21
cc_4549 ( N_noxref_23_c_7521_n N_noxref_24_c_7956_n ) capacitor c=0.0031527f \
 //x=71.78 //y=2.08 //x2=71.715 //y2=5.21
cc_4550 ( N_noxref_23_M130_noxref_g N_noxref_24_c_7956_n ) capacitor \
 c=0.0109874f //x=70.03 //y=6.025 //x2=71.715 //y2=5.21
cc_4551 ( N_noxref_23_M131_noxref_g N_noxref_24_c_7956_n ) capacitor \
 c=0.00645933f //x=72.05 //y=6.025 //x2=71.715 //y2=5.21
cc_4552 ( N_noxref_23_c_7565_n N_noxref_24_c_7956_n ) capacitor c=0.00270424f \
 //x=70.03 //y=4.87 //x2=71.715 //y2=5.21
cc_4553 ( N_noxref_23_c_7566_n N_noxref_24_c_7956_n ) capacitor c=0.00176728f \
 //x=72.125 //y=4.795 //x2=71.715 //y2=5.21
cc_4554 ( N_noxref_23_c_7498_n N_noxref_24_c_7960_n ) capacitor c=3.75024e-19 \
 //x=70.185 //y=2.96 //x2=69.925 //y2=5.21
cc_4555 ( N_noxref_23_M129_noxref_g N_noxref_24_c_7960_n ) capacitor \
 c=6.87102e-19 //x=69.59 //y=6.025 //x2=69.925 //y2=5.21
cc_4556 ( N_noxref_23_M130_noxref_g N_noxref_24_c_7960_n ) capacitor \
 c=8.33934e-19 //x=70.03 //y=6.025 //x2=69.925 //y2=5.21
cc_4557 ( N_noxref_23_M129_noxref_g N_noxref_24_c_7971_n ) capacitor \
 c=0.0179287f //x=69.59 //y=6.025 //x2=69.725 //y2=5.21
cc_4558 ( N_noxref_23_M129_noxref_g N_noxref_24_c_7963_n ) capacitor \
 c=0.0019882f //x=69.59 //y=6.025 //x2=69.81 //y2=5.295
cc_4559 ( N_noxref_23_M130_noxref_g N_noxref_24_c_7963_n ) capacitor \
 c=0.0159381f //x=70.03 //y=6.025 //x2=69.81 //y2=5.295
cc_4560 ( N_noxref_23_c_7863_p N_noxref_24_c_7963_n ) capacitor c=0.00456817f \
 //x=69.955 //y=4.795 //x2=69.81 //y2=5.295
cc_4561 ( N_noxref_23_c_7521_n N_noxref_24_c_7964_n ) capacitor c=0.0184695f \
 //x=71.78 //y=2.08 //x2=71.83 //y2=5.21
cc_4562 ( N_noxref_23_M131_noxref_g N_noxref_24_c_7964_n ) capacitor \
 c=0.0484795f //x=72.05 //y=6.025 //x2=71.83 //y2=5.21
cc_4563 ( N_noxref_23_c_7566_n N_noxref_24_c_7964_n ) capacitor c=0.0078825f \
 //x=72.125 //y=4.795 //x2=71.83 //y2=5.21
cc_4564 ( N_noxref_23_M131_noxref_g N_noxref_24_c_7983_n ) capacitor \
 c=0.0164606f //x=72.05 //y=6.025 //x2=72.625 //y2=6.91
cc_4565 ( N_noxref_23_M132_noxref_g N_noxref_24_c_7983_n ) capacitor \
 c=0.0150104f //x=72.49 //y=6.025 //x2=72.625 //y2=6.91
cc_4566 ( N_noxref_23_M129_noxref_g N_noxref_24_M129_noxref_d ) capacitor \
 c=0.0129738f //x=69.59 //y=6.025 //x2=69.665 //y2=5.025
cc_4567 ( N_noxref_23_M132_noxref_g N_noxref_24_M132_noxref_d ) capacitor \
 c=0.0130327f //x=72.49 //y=6.025 //x2=72.565 //y2=5.025
cc_4568 ( N_noxref_23_c_7498_n N_QN_c_8045_n ) capacitor c=0.0489549f \
 //x=70.185 //y=2.96 //x2=69.745 //y2=1.18
cc_4569 ( N_noxref_23_c_7789_n N_QN_c_8045_n ) capacitor c=5.17481e-19 \
 //x=69.595 //y=0.905 //x2=69.745 //y2=1.18
cc_4570 ( N_noxref_23_c_7792_n N_QN_c_8045_n ) capacitor c=0.00609699f \
 //x=69.595 //y=1.25 //x2=69.745 //y2=1.18
cc_4571 ( N_noxref_23_c_7498_n N_QN_c_8052_n ) capacitor c=0.00467724f \
 //x=70.185 //y=2.96 //x2=66.645 //y2=1.18
cc_4572 ( N_noxref_23_c_7498_n N_QN_c_8053_n ) capacitor c=0.00337366f \
 //x=70.185 //y=2.96 //x2=73.075 //y2=1.18
cc_4573 ( N_noxref_23_c_7513_n N_QN_c_8053_n ) capacitor c=0.053129f \
 //x=71.665 //y=2.08 //x2=73.075 //y2=1.18
cc_4574 ( N_noxref_23_c_7514_n N_QN_c_8053_n ) capacitor c=0.0102038f \
 //x=70.415 //y=2.08 //x2=73.075 //y2=1.18
cc_4575 ( N_noxref_23_c_7519_n N_QN_c_8053_n ) capacitor c=0.00189559f \
 //x=70.3 //y=2.08 //x2=73.075 //y2=1.18
cc_4576 ( N_noxref_23_c_7521_n N_QN_c_8053_n ) capacitor c=0.00134607f \
 //x=71.78 //y=2.08 //x2=73.075 //y2=1.18
cc_4577 ( N_noxref_23_c_7798_n N_QN_c_8053_n ) capacitor c=4.67724e-19 \
 //x=70.125 //y=0.905 //x2=73.075 //y2=1.18
cc_4578 ( N_noxref_23_c_7799_n N_QN_c_8053_n ) capacitor c=0.00591245f \
 //x=70.125 //y=1.25 //x2=73.075 //y2=1.18
cc_4579 ( N_noxref_23_c_7800_n N_QN_c_8053_n ) capacitor c=0.00326119f \
 //x=70.125 //y=1.56 //x2=73.075 //y2=1.18
cc_4580 ( N_noxref_23_c_7522_n N_QN_c_8053_n ) capacitor c=2.04565e-19 \
 //x=70.125 //y=1.915 //x2=73.075 //y2=1.18
cc_4581 ( N_noxref_23_c_7525_n N_QN_c_8053_n ) capacitor c=0.00500281f \
 //x=71.955 //y=1.21 //x2=73.075 //y2=1.18
cc_4582 ( N_noxref_23_c_7828_n N_QN_c_8053_n ) capacitor c=0.00361177f \
 //x=71.955 //y=1.52 //x2=73.075 //y2=1.18
cc_4583 ( N_noxref_23_c_7527_n N_QN_c_8053_n ) capacitor c=4.02408e-19 \
 //x=72.33 //y=0.71 //x2=73.075 //y2=1.18
cc_4584 ( N_noxref_23_c_7528_n N_QN_c_8053_n ) capacitor c=0.0036677f \
 //x=72.33 //y=1.365 //x2=73.075 //y2=1.18
cc_4585 ( N_noxref_23_c_7531_n N_QN_c_8053_n ) capacitor c=0.00776505f \
 //x=72.485 //y=1.21 //x2=73.075 //y2=1.18
cc_4586 ( N_noxref_23_c_7498_n N_QN_c_8059_n ) capacitor c=0.00413336f \
 //x=70.185 //y=2.96 //x2=69.975 //y2=1.18
cc_4587 ( N_noxref_23_c_7792_n N_QN_c_8059_n ) capacitor c=0.0015439f \
 //x=69.595 //y=1.25 //x2=69.975 //y2=1.18
cc_4588 ( N_noxref_23_c_7891_p N_QN_c_8059_n ) capacitor c=4.52813e-19 \
 //x=69.97 //y=0.75 //x2=69.975 //y2=1.18
cc_4589 ( N_noxref_23_c_7892_p N_QN_c_8059_n ) capacitor c=7.42023e-19 \
 //x=69.97 //y=1.405 //x2=69.975 //y2=1.18
cc_4590 ( N_noxref_23_c_7799_n N_QN_c_8059_n ) capacitor c=4.79299e-19 \
 //x=70.125 //y=1.25 //x2=69.975 //y2=1.18
cc_4591 ( N_noxref_23_c_7800_n N_QN_c_8059_n ) capacitor c=9.64184e-19 \
 //x=70.125 //y=1.56 //x2=69.975 //y2=1.18
cc_4592 ( N_noxref_23_c_7521_n QN ) capacitor c=0.00370801f //x=71.78 //y=2.08 \
 //x2=73.63 //y2=2.22
cc_4593 ( N_noxref_23_M132_noxref_g N_QN_c_8112_n ) capacitor c=0.0179287f \
 //x=72.49 //y=6.025 //x2=73.065 //y2=5.21
cc_4594 ( N_noxref_23_M131_noxref_g N_QN_c_8074_n ) capacitor c=0.0132916f \
 //x=72.05 //y=6.025 //x2=72.355 //y2=5.21
cc_4595 ( N_noxref_23_c_7830_n N_QN_c_8074_n ) capacitor c=0.00405122f \
 //x=72.415 //y=4.795 //x2=72.355 //y2=5.21
cc_4596 ( N_noxref_23_c_7498_n N_QN_M40_noxref_d ) capacitor c=0.00446326f \
 //x=70.185 //y=2.96 //x2=66.34 //y2=0.905
cc_4597 ( N_noxref_23_c_7498_n N_QN_M42_noxref_d ) capacitor c=0.00446423f \
 //x=70.185 //y=2.96 //x2=69.67 //y2=0.905
cc_4598 ( N_noxref_23_c_7789_n N_QN_M42_noxref_d ) capacitor c=0.00217566f \
 //x=69.595 //y=0.905 //x2=69.67 //y2=0.905
cc_4599 ( N_noxref_23_c_7792_n N_QN_M42_noxref_d ) capacitor c=0.00711747f \
 //x=69.595 //y=1.25 //x2=69.67 //y2=0.905
cc_4600 ( N_noxref_23_c_7891_p N_QN_M42_noxref_d ) capacitor c=0.00234223f \
 //x=69.97 //y=0.75 //x2=69.67 //y2=0.905
cc_4601 ( N_noxref_23_c_7892_p N_QN_M42_noxref_d ) capacitor c=0.00602848f \
 //x=69.97 //y=1.405 //x2=69.67 //y2=0.905
cc_4602 ( N_noxref_23_c_7798_n N_QN_M42_noxref_d ) capacitor c=0.00132245f \
 //x=70.125 //y=0.905 //x2=69.67 //y2=0.905
cc_4603 ( N_noxref_23_c_7799_n N_QN_M42_noxref_d ) capacitor c=0.004434f \
 //x=70.125 //y=1.25 //x2=69.67 //y2=0.905
cc_4604 ( N_noxref_23_c_7800_n N_QN_M42_noxref_d ) capacitor c=0.00270197f \
 //x=70.125 //y=1.56 //x2=69.67 //y2=0.905
cc_4605 ( N_noxref_23_M132_noxref_g N_QN_M131_noxref_d ) capacitor \
 c=0.0130327f //x=72.49 //y=6.025 //x2=72.125 //y2=5.025
cc_4606 ( N_noxref_23_c_7592_n N_noxref_31_c_8479_n ) capacitor c=0.00623646f \
 //x=16.685 //y=1.56 //x2=16.465 //y2=1.495
cc_4607 ( N_noxref_23_c_7597_n N_noxref_31_c_8479_n ) capacitor c=0.00174019f \
 //x=16.65 //y=2.08 //x2=16.465 //y2=1.495
cc_4608 ( N_noxref_23_c_7515_n N_noxref_31_c_8480_n ) capacitor c=0.00158203f \
 //x=16.65 //y=2.08 //x2=17.35 //y2=0.53
cc_4609 ( N_noxref_23_c_7587_n N_noxref_31_c_8480_n ) capacitor c=0.0188655f \
 //x=16.685 //y=0.905 //x2=17.35 //y2=0.53
cc_4610 ( N_noxref_23_c_7595_n N_noxref_31_c_8480_n ) capacitor c=0.00656458f \
 //x=17.215 //y=0.905 //x2=17.35 //y2=0.53
cc_4611 ( N_noxref_23_c_7597_n N_noxref_31_c_8480_n ) capacitor c=2.1838e-19 \
 //x=16.65 //y=2.08 //x2=17.35 //y2=0.53
cc_4612 ( N_noxref_23_c_7587_n N_noxref_31_M9_noxref_s ) capacitor \
 c=0.00623646f //x=16.685 //y=0.905 //x2=15.36 //y2=0.365
cc_4613 ( N_noxref_23_c_7595_n N_noxref_31_M9_noxref_s ) capacitor \
 c=0.0143002f //x=17.215 //y=0.905 //x2=15.36 //y2=0.365
cc_4614 ( N_noxref_23_c_7596_n N_noxref_31_M9_noxref_s ) capacitor \
 c=0.00290153f //x=17.215 //y=1.25 //x2=15.36 //y2=0.365
cc_4615 ( N_noxref_23_c_7713_n N_noxref_32_c_8543_n ) capacitor c=3.15806e-19 \
 //x=20.365 //y=1.655 //x2=18.825 //y2=1.495
cc_4616 ( N_noxref_23_c_7713_n N_noxref_32_c_8531_n ) capacitor c=0.0203424f \
 //x=20.365 //y=1.655 //x2=19.795 //y2=1.495
cc_4617 ( N_noxref_23_c_7517_n N_noxref_32_c_8532_n ) capacitor c=0.00461444f \
 //x=20.635 //y=1.655 //x2=20.68 //y2=0.53
cc_4618 ( N_noxref_23_M12_noxref_d N_noxref_32_c_8532_n ) capacitor \
 c=0.0116735f //x=20.09 //y=0.905 //x2=20.68 //y2=0.53
cc_4619 ( N_noxref_23_c_7517_n N_noxref_32_M11_noxref_s ) capacitor \
 c=0.0137901f //x=20.635 //y=1.655 //x2=18.69 //y2=0.365
cc_4620 ( N_noxref_23_M12_noxref_d N_noxref_32_M11_noxref_s ) capacitor \
 c=0.043966f //x=20.09 //y=0.905 //x2=18.69 //y2=0.365
cc_4621 ( N_noxref_23_c_7517_n N_noxref_33_c_8593_n ) capacitor c=4.08644e-19 \
 //x=20.635 //y=1.655 //x2=22.05 //y2=1.505
cc_4622 ( N_noxref_23_M12_noxref_d N_noxref_33_M13_noxref_s ) capacitor \
 c=2.53688e-19 //x=20.09 //y=0.905 //x2=21.915 //y2=0.375
cc_4623 ( N_noxref_23_c_7498_n N_noxref_47_M39_noxref_s ) capacitor \
 c=0.00285734f //x=70.185 //y=2.96 //x2=64.94 //y2=0.365
cc_4624 ( N_noxref_23_c_7498_n N_noxref_48_c_9384_n ) capacitor c=0.00256304f \
 //x=70.185 //y=2.96 //x2=68.405 //y2=1.495
cc_4625 ( N_noxref_23_c_7498_n N_noxref_48_c_9366_n ) capacitor c=0.0114954f \
 //x=70.185 //y=2.96 //x2=69.29 //y2=1.58
cc_4626 ( N_noxref_23_c_7498_n N_noxref_48_c_9372_n ) capacitor c=0.00285734f \
 //x=70.185 //y=2.96 //x2=69.375 //y2=1.495
cc_4627 ( N_noxref_23_c_7522_n N_noxref_48_c_9372_n ) capacitor c=0.0028747f \
 //x=70.125 //y=1.915 //x2=69.375 //y2=1.495
cc_4628 ( N_noxref_23_c_7789_n N_noxref_48_c_9373_n ) capacitor c=0.021566f \
 //x=69.595 //y=0.905 //x2=70.26 //y2=0.53
cc_4629 ( N_noxref_23_c_7798_n N_noxref_48_c_9373_n ) capacitor c=0.00781103f \
 //x=70.125 //y=0.905 //x2=70.26 //y2=0.53
cc_4630 ( N_noxref_23_c_7513_n N_noxref_48_M41_noxref_s ) capacitor \
 c=5.34178e-19 //x=71.665 //y=2.08 //x2=68.27 //y2=0.365
cc_4631 ( N_noxref_23_c_7514_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.00116116f //x=70.415 //y=2.08 //x2=68.27 //y2=0.365
cc_4632 ( N_noxref_23_c_7519_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.0149616f //x=70.3 //y=2.08 //x2=68.27 //y2=0.365
cc_4633 ( N_noxref_23_c_7789_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.0064603f //x=69.595 //y=0.905 //x2=68.27 //y2=0.365
cc_4634 ( N_noxref_23_c_7792_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.00602248f //x=69.595 //y=1.25 //x2=68.27 //y2=0.365
cc_4635 ( N_noxref_23_c_7798_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.0321601f //x=70.125 //y=0.905 //x2=68.27 //y2=0.365
cc_4636 ( N_noxref_23_c_7800_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.00239072f //x=70.125 //y=1.56 //x2=68.27 //y2=0.365
cc_4637 ( N_noxref_23_c_7522_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.00784558f //x=70.125 //y=1.915 //x2=68.27 //y2=0.365
cc_4638 ( N_noxref_23_c_7513_n N_noxref_49_c_9449_n ) capacitor c=0.00169534f \
 //x=71.665 //y=2.08 //x2=71.735 //y2=1.495
cc_4639 ( N_noxref_23_c_7521_n N_noxref_49_c_9449_n ) capacitor c=0.016698f \
 //x=71.78 //y=2.08 //x2=71.735 //y2=1.495
cc_4640 ( N_noxref_23_c_7526_n N_noxref_49_c_9449_n ) capacitor c=0.0034165f \
 //x=71.955 //y=1.915 //x2=71.735 //y2=1.495
cc_4641 ( N_noxref_23_c_7532_n N_noxref_49_c_9449_n ) capacitor c=0.00531095f \
 //x=71.78 //y=2.08 //x2=71.735 //y2=1.495
cc_4642 ( N_noxref_23_c_7513_n N_noxref_49_c_9422_n ) capacitor c=0.00222439f \
 //x=71.665 //y=2.08 //x2=72.62 //y2=1.58
cc_4643 ( N_noxref_23_c_7521_n N_noxref_49_c_9422_n ) capacitor c=0.00587616f \
 //x=71.78 //y=2.08 //x2=72.62 //y2=1.58
cc_4644 ( N_noxref_23_c_7828_n N_noxref_49_c_9422_n ) capacitor c=0.0061593f \
 //x=71.955 //y=1.52 //x2=72.62 //y2=1.58
cc_4645 ( N_noxref_23_c_7526_n N_noxref_49_c_9422_n ) capacitor c=0.0142098f \
 //x=71.955 //y=1.915 //x2=72.62 //y2=1.58
cc_4646 ( N_noxref_23_c_7528_n N_noxref_49_c_9422_n ) capacitor c=0.00991953f \
 //x=72.33 //y=1.365 //x2=72.62 //y2=1.58
cc_4647 ( N_noxref_23_c_7531_n N_noxref_49_c_9422_n ) capacitor c=0.00339872f \
 //x=72.485 //y=1.21 //x2=72.62 //y2=1.58
cc_4648 ( N_noxref_23_c_7532_n N_noxref_49_c_9422_n ) capacitor c=0.00147967f \
 //x=71.78 //y=2.08 //x2=72.62 //y2=1.58
cc_4649 ( N_noxref_23_c_7526_n N_noxref_49_c_9428_n ) capacitor c=6.71402e-19 \
 //x=71.955 //y=1.915 //x2=72.705 //y2=1.495
cc_4650 ( N_noxref_23_c_7523_n N_noxref_49_M43_noxref_s ) capacitor \
 c=0.0314164f //x=71.955 //y=0.865 //x2=71.6 //y2=0.365
cc_4651 ( N_noxref_23_c_7828_n N_noxref_49_M43_noxref_s ) capacitor \
 c=0.00110192f //x=71.955 //y=1.52 //x2=71.6 //y2=0.365
cc_4652 ( N_noxref_23_c_7529_n N_noxref_49_M43_noxref_s ) capacitor \
 c=0.0132463f //x=72.485 //y=0.865 //x2=71.6 //y2=0.365
cc_4653 ( N_noxref_24_c_7964_n QN ) capacitor c=3.02032e-19 //x=71.83 //y=5.21 \
 //x2=73.63 //y2=2.22
cc_4654 ( N_noxref_24_c_7983_n N_QN_c_8112_n ) capacitor c=0.00102709f \
 //x=72.625 //y=6.91 //x2=73.065 //y2=5.21
cc_4655 ( N_noxref_24_c_7984_n N_QN_c_8112_n ) capacitor c=0.00101874f \
 //x=73.505 //y=6.91 //x2=73.065 //y2=5.21
cc_4656 ( N_noxref_24_M132_noxref_d N_QN_c_8112_n ) capacitor c=0.012404f \
 //x=72.565 //y=5.025 //x2=73.065 //y2=5.21
cc_4657 ( N_noxref_24_c_7956_n N_QN_c_8074_n ) capacitor c=0.00602307f \
 //x=71.715 //y=5.21 //x2=72.355 //y2=5.21
cc_4658 ( N_noxref_24_c_7964_n N_QN_c_8074_n ) capacitor c=0.0683084f \
 //x=71.83 //y=5.21 //x2=72.355 //y2=5.21
cc_4659 ( N_noxref_24_c_7984_n N_QN_c_8075_n ) capacitor c=0.00173777f \
 //x=73.505 //y=6.91 //x2=73.545 //y2=5.21
cc_4660 ( N_noxref_24_M134_noxref_d N_QN_c_8075_n ) capacitor c=0.0159033f \
 //x=73.445 //y=5.025 //x2=73.545 //y2=5.21
cc_4661 ( N_noxref_24_c_7956_n N_QN_M131_noxref_d ) capacitor c=8.04912e-19 \
 //x=71.715 //y=5.21 //x2=72.125 //y2=5.025
cc_4662 ( N_noxref_24_c_7983_n N_QN_M131_noxref_d ) capacitor c=0.0117542f \
 //x=72.625 //y=6.91 //x2=72.125 //y2=5.025
cc_4663 ( N_noxref_24_M132_noxref_d N_QN_M131_noxref_d ) capacitor \
 c=0.0458293f //x=72.565 //y=5.025 //x2=72.125 //y2=5.025
cc_4664 ( N_noxref_24_c_7964_n N_QN_M133_noxref_d ) capacitor c=9.91979e-19 \
 //x=71.83 //y=5.21 //x2=73.005 //y2=5.025
cc_4665 ( N_noxref_24_c_7984_n N_QN_M133_noxref_d ) capacitor c=0.0118172f \
 //x=73.505 //y=6.91 //x2=73.005 //y2=5.025
cc_4666 ( N_noxref_24_M132_noxref_d N_QN_M133_noxref_d ) capacitor \
 c=0.0458293f //x=72.565 //y=5.025 //x2=73.005 //y2=5.025
cc_4667 ( N_noxref_24_M134_noxref_d N_QN_M133_noxref_d ) capacitor \
 c=0.0458293f //x=73.445 //y=5.025 //x2=73.005 //y2=5.025
cc_4668 ( N_QN_c_8045_n N_noxref_47_c_9316_n ) capacitor c=0.00641749f \
 //x=69.745 //y=1.18 //x2=66.93 //y2=0.53
cc_4669 ( N_QN_c_8052_n N_noxref_47_c_9316_n ) capacitor c=0.00219859f \
 //x=66.645 //y=1.18 //x2=66.93 //y2=0.53
cc_4670 ( N_QN_M40_noxref_d N_noxref_47_c_9316_n ) capacitor c=0.0136817f \
 //x=66.34 //y=0.905 //x2=66.93 //y2=0.53
cc_4671 ( N_QN_c_8045_n N_noxref_47_M39_noxref_s ) capacitor c=0.0207977f \
 //x=69.745 //y=1.18 //x2=64.94 //y2=0.365
cc_4672 ( N_QN_c_8052_n N_noxref_47_M39_noxref_s ) capacitor c=0.00804471f \
 //x=66.645 //y=1.18 //x2=64.94 //y2=0.365
cc_4673 ( N_QN_M40_noxref_d N_noxref_47_M39_noxref_s ) capacitor c=0.0458734f \
 //x=66.34 //y=0.905 //x2=64.94 //y2=0.365
cc_4674 ( N_QN_c_8045_n N_noxref_48_c_9366_n ) capacitor c=0.0224452f \
 //x=69.745 //y=1.18 //x2=69.29 //y2=1.58
cc_4675 ( N_QN_c_8045_n N_noxref_48_c_9373_n ) capacitor c=0.00641749f \
 //x=69.745 //y=1.18 //x2=70.26 //y2=0.53
cc_4676 ( N_QN_c_8053_n N_noxref_48_c_9373_n ) capacitor c=0.00641749f \
 //x=73.075 //y=1.18 //x2=70.26 //y2=0.53
cc_4677 ( N_QN_c_8059_n N_noxref_48_c_9373_n ) capacitor c=0.0015838f \
 //x=69.975 //y=1.18 //x2=70.26 //y2=0.53
cc_4678 ( N_QN_M42_noxref_d N_noxref_48_c_9373_n ) capacitor c=0.0130616f \
 //x=69.67 //y=0.905 //x2=70.26 //y2=0.53
cc_4679 ( N_QN_c_8045_n N_noxref_48_M41_noxref_s ) capacitor c=0.0443893f \
 //x=69.745 //y=1.18 //x2=68.27 //y2=0.365
cc_4680 ( N_QN_c_8053_n N_noxref_48_M41_noxref_s ) capacitor c=0.019112f \
 //x=73.075 //y=1.18 //x2=68.27 //y2=0.365
cc_4681 ( N_QN_c_8059_n N_noxref_48_M41_noxref_s ) capacitor c=0.00279707f \
 //x=69.975 //y=1.18 //x2=68.27 //y2=0.365
cc_4682 ( N_QN_M42_noxref_d N_noxref_48_M41_noxref_s ) capacitor c=0.0444718f \
 //x=69.67 //y=0.905 //x2=68.27 //y2=0.365
cc_4683 ( N_QN_c_8119_n N_noxref_49_c_9449_n ) capacitor c=2.73698e-19 \
 //x=73.275 //y=1.645 //x2=71.735 //y2=1.495
cc_4684 ( N_QN_c_8053_n N_noxref_49_c_9422_n ) capacitor c=0.0234642f \
 //x=73.075 //y=1.18 //x2=72.62 //y2=1.58
cc_4685 ( N_QN_c_8119_n N_noxref_49_c_9428_n ) capacitor c=0.0195484f \
 //x=73.275 //y=1.645 //x2=72.705 //y2=1.495
cc_4686 ( N_QN_c_8053_n N_noxref_49_c_9429_n ) capacitor c=0.0069137f \
 //x=73.075 //y=1.18 //x2=73.59 //y2=0.53
cc_4687 ( N_QN_c_8061_n N_noxref_49_c_9429_n ) capacitor c=0.00458011f \
 //x=73.545 //y=1.645 //x2=73.59 //y2=0.53
cc_4688 ( N_QN_M44_noxref_d N_noxref_49_c_9429_n ) capacitor c=0.0132979f \
 //x=73 //y=0.905 //x2=73.59 //y2=0.53
cc_4689 ( N_QN_c_8053_n N_noxref_49_M43_noxref_s ) capacitor c=0.0513705f \
 //x=73.075 //y=1.18 //x2=71.6 //y2=0.365
cc_4690 ( N_QN_c_8061_n N_noxref_49_M43_noxref_s ) capacitor c=0.0155576f \
 //x=73.545 //y=1.645 //x2=71.6 //y2=0.365
cc_4691 ( N_QN_M44_noxref_d N_noxref_49_M43_noxref_s ) capacitor c=0.0438441f \
 //x=73 //y=0.905 //x2=71.6 //y2=0.365
cc_4692 ( N_noxref_26_c_8221_n N_noxref_27_c_8261_n ) capacitor c=0.0136048f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_4693 ( N_noxref_26_c_8239_n N_noxref_27_c_8261_n ) capacitor c=0.0102225f \
 //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_4694 ( N_noxref_26_M0_noxref_s N_noxref_27_c_8261_n ) capacitor \
 c=0.0228676f //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_4695 ( N_noxref_26_M0_noxref_s N_noxref_27_c_8263_n ) capacitor \
 c=0.0180035f //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_4696 ( N_noxref_26_c_8221_n N_noxref_27_M1_noxref_d ) capacitor \
 c=0.0129526f //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_4697 ( N_noxref_26_c_8239_n N_noxref_27_M1_noxref_d ) capacitor \
 c=0.00908243f //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_4698 ( N_noxref_26_M0_noxref_s N_noxref_27_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_4699 ( N_noxref_26_M0_noxref_s N_noxref_27_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_4700 ( N_noxref_27_c_8269_n N_noxref_28_M3_noxref_s ) capacitor \
 c=0.00164795f //x=4.07 //y=0.625 //x2=5.37 //y2=0.365
cc_4701 ( N_noxref_28_c_8325_n N_noxref_29_M5_noxref_s ) capacitor \
 c=0.00174327f //x=7.445 //y=0.615 //x2=8.7 //y2=0.365
cc_4702 ( N_noxref_29_c_8379_n N_noxref_30_M7_noxref_s ) capacitor \
 c=0.00174327f //x=10.775 //y=0.615 //x2=12.03 //y2=0.365
cc_4703 ( N_noxref_30_c_8431_n N_noxref_31_M9_noxref_s ) capacitor \
 c=0.00174327f //x=14.105 //y=0.615 //x2=15.36 //y2=0.365
cc_4704 ( N_noxref_31_c_8483_n N_noxref_32_M11_noxref_s ) capacitor \
 c=0.00174327f //x=17.435 //y=0.615 //x2=18.69 //y2=0.365
cc_4705 ( N_noxref_32_c_8535_n N_noxref_33_M13_noxref_s ) capacitor \
 c=0.00199452f //x=20.765 //y=0.615 //x2=21.915 //y2=0.375
cc_4706 ( N_noxref_33_c_8583_n N_noxref_34_c_8626_n ) capacitor c=0.0133059f \
 //x=23.905 //y=0.54 //x2=24.475 //y2=0.995
cc_4707 ( N_noxref_33_c_8605_n N_noxref_34_c_8626_n ) capacitor c=0.0100097f \
 //x=23.905 //y=1.59 //x2=24.475 //y2=0.995
cc_4708 ( N_noxref_33_M13_noxref_s N_noxref_34_c_8626_n ) capacitor \
 c=0.0224457f //x=21.915 //y=0.375 //x2=24.475 //y2=0.995
cc_4709 ( N_noxref_33_M13_noxref_s N_noxref_34_c_8628_n ) capacitor \
 c=0.0180035f //x=21.915 //y=0.375 //x2=24.56 //y2=0.625
cc_4710 ( N_noxref_33_c_8583_n N_noxref_34_M14_noxref_d ) capacitor \
 c=0.0128027f //x=23.905 //y=0.54 //x2=23.32 //y2=0.91
cc_4711 ( N_noxref_33_c_8605_n N_noxref_34_M14_noxref_d ) capacitor \
 c=0.00879751f //x=23.905 //y=1.59 //x2=23.32 //y2=0.91
cc_4712 ( N_noxref_33_M13_noxref_s N_noxref_34_M14_noxref_d ) capacitor \
 c=0.0159202f //x=21.915 //y=0.375 //x2=23.32 //y2=0.91
cc_4713 ( N_noxref_33_M13_noxref_s N_noxref_34_M15_noxref_s ) capacitor \
 c=0.0213553f //x=21.915 //y=0.375 //x2=24.425 //y2=0.375
cc_4714 ( N_noxref_34_c_8634_n N_noxref_35_M16_noxref_s ) capacitor \
 c=0.00164795f //x=25.53 //y=0.625 //x2=26.83 //y2=0.365
cc_4715 ( N_noxref_35_c_8690_n N_noxref_36_M18_noxref_s ) capacitor \
 c=0.00174327f //x=28.905 //y=0.615 //x2=30.16 //y2=0.365
cc_4716 ( N_noxref_36_c_8744_n N_noxref_37_M20_noxref_s ) capacitor \
 c=0.00174327f //x=32.235 //y=0.615 //x2=33.49 //y2=0.365
cc_4717 ( N_noxref_37_c_8796_n N_noxref_38_M22_noxref_s ) capacitor \
 c=0.00174327f //x=35.565 //y=0.615 //x2=36.82 //y2=0.365
cc_4718 ( N_noxref_38_c_8848_n N_noxref_39_M24_noxref_s ) capacitor \
 c=0.00174327f //x=38.895 //y=0.615 //x2=40.15 //y2=0.365
cc_4719 ( N_noxref_39_c_8902_n N_noxref_40_M26_noxref_s ) capacitor \
 c=0.00199452f //x=42.225 //y=0.615 //x2=43.375 //y2=0.375
cc_4720 ( N_noxref_40_c_8952_n N_noxref_41_c_8995_n ) capacitor c=0.0131877f \
 //x=45.365 //y=0.54 //x2=45.935 //y2=0.995
cc_4721 ( N_noxref_40_c_8963_n N_noxref_41_c_8995_n ) capacitor c=0.00981707f \
 //x=45.365 //y=1.59 //x2=45.935 //y2=0.995
cc_4722 ( N_noxref_40_M26_noxref_s N_noxref_41_c_8995_n ) capacitor \
 c=0.0221661f //x=43.375 //y=0.375 //x2=45.935 //y2=0.995
cc_4723 ( N_noxref_40_M26_noxref_s N_noxref_41_c_8997_n ) capacitor \
 c=0.0180035f //x=43.375 //y=0.375 //x2=46.02 //y2=0.625
cc_4724 ( N_noxref_40_c_8952_n N_noxref_41_M27_noxref_d ) capacitor \
 c=0.0127191f //x=45.365 //y=0.54 //x2=44.78 //y2=0.91
cc_4725 ( N_noxref_40_c_8963_n N_noxref_41_M27_noxref_d ) capacitor \
 c=0.00861161f //x=45.365 //y=1.59 //x2=44.78 //y2=0.91
cc_4726 ( N_noxref_40_M26_noxref_s N_noxref_41_M27_noxref_d ) capacitor \
 c=0.0159202f //x=43.375 //y=0.375 //x2=44.78 //y2=0.91
cc_4727 ( N_noxref_40_M26_noxref_s N_noxref_41_M28_noxref_s ) capacitor \
 c=0.0213553f //x=43.375 //y=0.375 //x2=45.885 //y2=0.375
cc_4728 ( N_noxref_41_c_9003_n N_noxref_42_M29_noxref_s ) capacitor \
 c=0.00164795f //x=46.99 //y=0.625 //x2=48.29 //y2=0.365
cc_4729 ( N_noxref_42_c_9059_n N_noxref_43_M31_noxref_s ) capacitor \
 c=0.00174327f //x=50.365 //y=0.615 //x2=51.62 //y2=0.365
cc_4730 ( N_noxref_43_c_9111_n N_noxref_44_M33_noxref_s ) capacitor \
 c=0.00174327f //x=53.695 //y=0.615 //x2=54.95 //y2=0.365
cc_4731 ( N_noxref_44_c_9163_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.00174327f //x=57.025 //y=0.615 //x2=58.28 //y2=0.365
cc_4732 ( N_noxref_45_c_9215_n N_noxref_46_M37_noxref_s ) capacitor \
 c=0.00174327f //x=60.355 //y=0.615 //x2=61.61 //y2=0.365
cc_4733 ( N_noxref_46_c_9267_n N_noxref_47_M39_noxref_s ) capacitor \
 c=0.00205929f //x=63.685 //y=0.615 //x2=64.94 //y2=0.365
cc_4734 ( N_noxref_47_M39_noxref_s N_noxref_48_c_9384_n ) capacitor \
 c=0.0011299f //x=64.94 //y=0.365 //x2=68.405 //y2=1.495
cc_4735 ( N_noxref_47_c_9319_n N_noxref_48_M41_noxref_s ) capacitor \
 c=0.0011299f //x=67.015 //y=0.615 //x2=68.27 //y2=0.365
cc_4736 ( N_noxref_48_M41_noxref_s N_noxref_49_c_9449_n ) capacitor \
 c=0.0011299f //x=68.27 //y=0.365 //x2=71.735 //y2=1.495
cc_4737 ( N_noxref_48_c_9376_n N_noxref_49_M43_noxref_s ) capacitor \
 c=0.0011299f //x=70.345 //y=0.615 //x2=71.6 //y2=0.365
