* SPICE3 file created from DLATCHN.ext - technology: sky130A

.subckt DLATCHN Q D GATE_N VDD VSS
X0 VDD a_1771_1050 a_2405_209 VDD sky130_fd_pr__pfet_01v8 ad=0.00892 pd=7.292 as=0 ps=0 w=2 l=0.15 M=2
X1 Q a_3007_411 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.003582 pd=3.15 as=0.0087946 ps=6.142 w=3 l=0.15
X2 VDD D a_1771_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X3 a_185_209 D VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X4 a_1295_209 a_661_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X5 a_1771_1050 D a_1666_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X6 a_661_1050 a_n259_209 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X7 VSS a_185_209 a_556_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X8 a_185_209 D VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X9 Q a_3007_411 a_2795_1051 VDD sky130_fd_pr__pfet_01v8 ad=0.0058 pd=4.58 as=0 ps=0 w=2 l=0.15 M=2
X10 a_3461_1051 a_2405_209 a_3007_411 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X11 a_661_1050 a_185_209 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X12 a_1771_1050 a_n259_209 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X13 a_2795_1051 a_1295_209 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X14 VDD Q a_3461_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X15 VDD GATE_N a_n259_209 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X16 a_3007_411 Q VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X17 a_661_1050 a_n259_209 a_556_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X18 VSS a_n259_209 a_1666_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X19 a_n259_209 GATE_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X20 a_1295_209 a_661_1050 VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X21 a_3007_411 a_2405_209 VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X22 Q a_1295_209 VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X23 a_2405_209 a_1771_1050 VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 a_661_1050 VDD 2.27f
C1 a_1771_1050 VDD 2.27f
C2 VDD VSS 7.44f
.ends
