// File: AOA4X1.spi.AOA4X1.pxi
// Created: Tue Oct 15 15:44:57 2024
// 
simulator lang=spectre
x_PM_AOA4X1\%GND ( GND N_GND_c_14_p N_GND_c_90_p N_GND_c_1_p N_GND_c_97_p \
 N_GND_c_116_p N_GND_c_6_p N_GND_c_22_p N_GND_c_34_p N_GND_c_37_p \
 N_GND_c_154_p N_GND_c_43_p N_GND_c_50_p N_GND_c_150_p N_GND_c_62_p \
 N_GND_c_79_p N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p N_GND_c_5_p \
 N_GND_M0_noxref_d N_GND_M2_noxref_s N_GND_M4_noxref_d N_GND_M6_noxref_s )  \
 PM_AOA4X1\%GND
x_PM_AOA4X1\%VDD ( VDD N_VDD_c_194_p N_VDD_c_176_p N_VDD_c_177_p N_VDD_c_188_p \
 N_VDD_c_191_p N_VDD_c_212_p N_VDD_c_224_p N_VDD_c_235_p N_VDD_c_170_n \
 N_VDD_c_171_n N_VDD_c_172_n N_VDD_c_173_n N_VDD_c_174_n N_VDD_M7_noxref_s \
 N_VDD_M8_noxref_d N_VDD_M10_noxref_d N_VDD_M11_noxref_d N_VDD_M15_noxref_s \
 N_VDD_M16_noxref_d N_VDD_M18_noxref_d N_VDD_M19_noxref_s N_VDD_M20_noxref_d ) \
 PM_AOA4X1\%VDD
x_PM_AOA4X1\%noxref_3 ( N_noxref_3_c_311_n N_noxref_3_c_314_n \
 N_noxref_3_c_334_n N_noxref_3_c_337_n N_noxref_3_c_339_n N_noxref_3_c_315_n \
 N_noxref_3_c_410_p N_noxref_3_c_317_n N_noxref_3_c_319_n N_noxref_3_c_398_p \
 N_noxref_3_c_344_n N_noxref_3_M2_noxref_g N_noxref_3_M11_noxref_g \
 N_noxref_3_M12_noxref_g N_noxref_3_c_322_n N_noxref_3_c_372_p \
 N_noxref_3_c_373_p N_noxref_3_c_324_n N_noxref_3_c_326_n N_noxref_3_c_376_p \
 N_noxref_3_c_419_p N_noxref_3_c_327_n N_noxref_3_c_329_n N_noxref_3_c_351_n \
 N_noxref_3_M1_noxref_d N_noxref_3_M7_noxref_d N_noxref_3_M9_noxref_d )  \
 PM_AOA4X1\%noxref_3
x_PM_AOA4X1\%noxref_4 ( N_noxref_4_c_455_n N_noxref_4_c_457_n \
 N_noxref_4_c_459_n N_noxref_4_c_507_n N_noxref_4_c_490_n N_noxref_4_c_492_n \
 N_noxref_4_c_463_n N_noxref_4_c_467_n N_noxref_4_c_469_n \
 N_noxref_4_M4_noxref_g N_noxref_4_M15_noxref_g N_noxref_4_M16_noxref_g \
 N_noxref_4_c_470_n N_noxref_4_c_472_n N_noxref_4_c_473_n N_noxref_4_c_474_n \
 N_noxref_4_c_475_n N_noxref_4_c_476_n N_noxref_4_c_477_n N_noxref_4_c_479_n \
 N_noxref_4_c_501_n N_noxref_4_M2_noxref_d N_noxref_4_M3_noxref_d \
 N_noxref_4_M13_noxref_d )  PM_AOA4X1\%noxref_4
x_PM_AOA4X1\%noxref_5 ( N_noxref_5_c_597_n N_noxref_5_c_600_n \
 N_noxref_5_c_625_n N_noxref_5_c_628_n N_noxref_5_c_630_n N_noxref_5_c_601_n \
 N_noxref_5_c_691_p N_noxref_5_c_603_n N_noxref_5_c_605_n N_noxref_5_c_679_p \
 N_noxref_5_M6_noxref_g N_noxref_5_M19_noxref_g N_noxref_5_M20_noxref_g \
 N_noxref_5_c_610_n N_noxref_5_c_711_p N_noxref_5_c_712_p N_noxref_5_c_612_n \
 N_noxref_5_c_642_n N_noxref_5_c_643_n N_noxref_5_c_613_n N_noxref_5_c_703_p \
 N_noxref_5_c_614_n N_noxref_5_c_616_n N_noxref_5_c_617_n \
 N_noxref_5_M5_noxref_d N_noxref_5_M15_noxref_d N_noxref_5_M17_noxref_d )  \
 PM_AOA4X1\%noxref_5
x_PM_AOA4X1\%A ( A A A A A A A N_A_c_723_n N_A_M0_noxref_g N_A_M7_noxref_g \
 N_A_M8_noxref_g N_A_c_724_n N_A_c_726_n N_A_c_727_n N_A_c_728_n N_A_c_729_n \
 N_A_c_730_n N_A_c_731_n N_A_c_733_n N_A_c_740_n )  PM_AOA4X1\%A
x_PM_AOA4X1\%B ( B B B B B B B N_B_c_787_n N_B_c_778_n N_B_M1_noxref_g \
 N_B_M9_noxref_g N_B_M10_noxref_g N_B_c_796_n N_B_c_797_n N_B_c_798_n \
 N_B_c_799_n N_B_c_801_n N_B_c_802_n N_B_c_804_n N_B_c_805_n N_B_c_807_n \
 N_B_c_808_n N_B_c_810_n )  PM_AOA4X1\%B
x_PM_AOA4X1\%noxref_8 ( N_noxref_8_c_866_n N_noxref_8_c_842_n \
 N_noxref_8_c_846_n N_noxref_8_c_850_n N_noxref_8_c_851_n N_noxref_8_c_854_n \
 N_noxref_8_M0_noxref_s )  PM_AOA4X1\%noxref_8
x_PM_AOA4X1\%C ( C C C C C C C N_C_c_906_n N_C_c_893_n N_C_M3_noxref_g \
 N_C_M13_noxref_g N_C_M14_noxref_g N_C_c_895_n N_C_c_918_n N_C_c_921_n \
 N_C_c_945_n N_C_c_897_n N_C_c_898_n N_C_c_899_n N_C_c_925_n N_C_c_926_n \
 N_C_c_928_n N_C_c_929_n )  PM_AOA4X1\%C
x_PM_AOA4X1\%noxref_10 ( N_noxref_10_c_964_n N_noxref_10_c_968_n \
 N_noxref_10_c_969_n N_noxref_10_c_970_n N_noxref_10_M11_noxref_s \
 N_noxref_10_M12_noxref_d N_noxref_10_M14_noxref_d )  PM_AOA4X1\%noxref_10
x_PM_AOA4X1\%D ( D D D D D D D N_D_c_1016_n N_D_c_1007_n N_D_M5_noxref_g \
 N_D_M17_noxref_g N_D_M18_noxref_g N_D_c_1025_n N_D_c_1028_n N_D_c_1030_n \
 N_D_c_1051_n N_D_c_1053_n N_D_c_1054_n N_D_c_1033_n N_D_c_1034_n N_D_c_1035_n \
 N_D_c_1060_n N_D_c_1037_n )  PM_AOA4X1\%D
x_PM_AOA4X1\%noxref_12 ( N_noxref_12_c_1098_n N_noxref_12_c_1073_n \
 N_noxref_12_c_1077_n N_noxref_12_c_1081_n N_noxref_12_c_1082_n \
 N_noxref_12_c_1085_n N_noxref_12_M4_noxref_s )  PM_AOA4X1\%noxref_12
x_PM_AOA4X1\%Y ( Y Y Y Y Y Y Y N_Y_c_1129_n N_Y_c_1152_n N_Y_c_1139_n \
 N_Y_c_1141_n N_Y_M6_noxref_d N_Y_M19_noxref_d )  PM_AOA4X1\%Y
cc_1 ( N_GND_c_1_p N_VDD_c_170_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_171_n ) capacitor c=0.00962895f //x=3.33 //y=0 \
 //x2=3.33 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_172_n ) capacitor c=0.00962895f //x=6.66 //y=0 \
 //x2=6.66 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_173_n ) capacitor c=0.00962895f //x=9.99 //y=0 \
 //x2=9.99 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_174_n ) capacitor c=0.00989031f //x=11.59 //y=0 \
 //x2=11.47 //y2=7.4
cc_6 ( N_GND_c_6_p N_noxref_3_c_311_n ) capacitor c=7.22787e-19 //x=4.425 \
 //y=0.53 //x2=4.325 //y2=2.59
cc_7 ( N_GND_c_2_p N_noxref_3_c_311_n ) capacitor c=0.0435449f //x=3.33 //y=0 \
 //x2=4.325 //y2=2.59
cc_8 ( N_GND_M2_noxref_s N_noxref_3_c_311_n ) capacitor c=0.00494344f //x=3.89 \
 //y=0.365 //x2=4.325 //y2=2.59
cc_9 ( N_GND_c_2_p N_noxref_3_c_314_n ) capacitor c=0.00102529f //x=3.33 //y=0 \
 //x2=2.705 //y2=2.59
cc_10 ( N_GND_c_2_p N_noxref_3_c_315_n ) capacitor c=0.0431271f //x=3.33 //y=0 \
 //x2=2.505 //y2=1.655
cc_11 ( N_GND_M2_noxref_s N_noxref_3_c_315_n ) capacitor c=3.00901e-19 \
 //x=3.89 //y=0.365 //x2=2.505 //y2=1.655
cc_12 ( N_GND_c_1_p N_noxref_3_c_317_n ) capacitor c=0.00101801f //x=0.74 \
 //y=0 //x2=2.59 //y2=2.59
cc_13 ( N_GND_c_2_p N_noxref_3_c_317_n ) capacitor c=5.56859e-19 //x=3.33 \
 //y=0 //x2=2.59 //y2=2.59
cc_14 ( N_GND_c_14_p N_noxref_3_c_319_n ) capacitor c=6.7762e-19 //x=11.47 \
 //y=0 //x2=4.44 //y2=2.08
cc_15 ( N_GND_c_6_p N_noxref_3_c_319_n ) capacitor c=0.00133118f //x=4.425 \
 //y=0.53 //x2=4.44 //y2=2.08
cc_16 ( N_GND_c_2_p N_noxref_3_c_319_n ) capacitor c=0.0147015f //x=3.33 //y=0 \
 //x2=4.44 //y2=2.08
cc_17 ( N_GND_c_6_p N_noxref_3_c_322_n ) capacitor c=0.0122561f //x=4.425 \
 //y=0.53 //x2=4.245 //y2=0.905
cc_18 ( N_GND_M2_noxref_s N_noxref_3_c_322_n ) capacitor c=0.0318086f //x=3.89 \
 //y=0.365 //x2=4.245 //y2=0.905
cc_19 ( N_GND_c_6_p N_noxref_3_c_324_n ) capacitor c=2.1838e-19 //x=4.425 \
 //y=0.53 //x2=4.245 //y2=1.915
cc_20 ( N_GND_c_2_p N_noxref_3_c_324_n ) capacitor c=0.0131707f //x=3.33 //y=0 \
 //x2=4.245 //y2=1.915
cc_21 ( N_GND_M2_noxref_s N_noxref_3_c_326_n ) capacitor c=0.00476335f \
 //x=3.89 //y=0.365 //x2=4.62 //y2=0.75
cc_22 ( N_GND_c_22_p N_noxref_3_c_327_n ) capacitor c=0.0113279f //x=4.91 \
 //y=0.53 //x2=4.775 //y2=0.905
cc_23 ( N_GND_M2_noxref_s N_noxref_3_c_327_n ) capacitor c=0.00514143f \
 //x=3.89 //y=0.365 //x2=4.775 //y2=0.905
cc_24 ( N_GND_M2_noxref_s N_noxref_3_c_329_n ) capacitor c=8.33128e-19 \
 //x=3.89 //y=0.365 //x2=4.775 //y2=1.25
cc_25 ( N_GND_c_1_p N_noxref_3_M1_noxref_d ) capacitor c=8.58106e-19 //x=0.74 \
 //y=0 //x2=1.96 //y2=0.905
cc_26 ( N_GND_c_2_p N_noxref_3_M1_noxref_d ) capacitor c=0.00616547f //x=3.33 \
 //y=0 //x2=1.96 //y2=0.905
cc_27 ( N_GND_M0_noxref_d N_noxref_3_M1_noxref_d ) capacitor c=0.00143464f \
 //x=0.99 //y=0.865 //x2=1.96 //y2=0.905
cc_28 ( N_GND_c_3_p N_noxref_4_c_455_n ) capacitor c=0.0435449f //x=6.66 //y=0 \
 //x2=7.655 //y2=2.59
cc_29 ( N_GND_M2_noxref_s N_noxref_4_c_455_n ) capacitor c=3.07321e-19 \
 //x=3.89 //y=0.365 //x2=7.655 //y2=2.59
cc_30 ( N_GND_c_3_p N_noxref_4_c_457_n ) capacitor c=0.00102529f //x=6.66 \
 //y=0 //x2=6.035 //y2=2.59
cc_31 ( N_GND_M2_noxref_s N_noxref_4_c_457_n ) capacitor c=0.00162156f \
 //x=3.89 //y=0.365 //x2=6.035 //y2=2.59
cc_32 ( N_GND_c_14_p N_noxref_4_c_459_n ) capacitor c=0.00359057f //x=11.47 \
 //y=0 //x2=5.395 //y2=1.655
cc_33 ( N_GND_c_22_p N_noxref_4_c_459_n ) capacitor c=0.00381844f //x=4.91 \
 //y=0.53 //x2=5.395 //y2=1.655
cc_34 ( N_GND_c_34_p N_noxref_4_c_459_n ) capacitor c=0.00323369f //x=5.395 \
 //y=0.53 //x2=5.395 //y2=1.655
cc_35 ( N_GND_M2_noxref_s N_noxref_4_c_459_n ) capacitor c=0.0173679f //x=3.89 \
 //y=0.365 //x2=5.395 //y2=1.655
cc_36 ( N_GND_c_14_p N_noxref_4_c_463_n ) capacitor c=0.00232664f //x=11.47 \
 //y=0 //x2=5.835 //y2=1.655
cc_37 ( N_GND_c_37_p N_noxref_4_c_463_n ) capacitor c=0.0047903f //x=5.88 \
 //y=0.53 //x2=5.835 //y2=1.655
cc_38 ( N_GND_c_3_p N_noxref_4_c_463_n ) capacitor c=0.04345f //x=6.66 //y=0 \
 //x2=5.835 //y2=1.655
cc_39 ( N_GND_M2_noxref_s N_noxref_4_c_463_n ) capacitor c=0.0145566f //x=3.89 \
 //y=0.365 //x2=5.835 //y2=1.655
cc_40 ( N_GND_c_2_p N_noxref_4_c_467_n ) capacitor c=9.64732e-19 //x=3.33 \
 //y=0 //x2=5.92 //y2=2.59
cc_41 ( N_GND_c_3_p N_noxref_4_c_467_n ) capacitor c=5.56859e-19 //x=6.66 \
 //y=0 //x2=5.92 //y2=2.59
cc_42 ( N_GND_c_3_p N_noxref_4_c_469_n ) capacitor c=0.0150626f //x=6.66 //y=0 \
 //x2=7.77 //y2=2.08
cc_43 ( N_GND_c_43_p N_noxref_4_c_470_n ) capacitor c=0.00135046f //x=7.755 \
 //y=0 //x2=7.575 //y2=0.865
cc_44 ( N_GND_M4_noxref_d N_noxref_4_c_470_n ) capacitor c=0.00220047f \
 //x=7.65 //y=0.865 //x2=7.575 //y2=0.865
cc_45 ( N_GND_M4_noxref_d N_noxref_4_c_472_n ) capacitor c=0.00255985f \
 //x=7.65 //y=0.865 //x2=7.575 //y2=1.21
cc_46 ( N_GND_c_3_p N_noxref_4_c_473_n ) capacitor c=0.0018059f //x=6.66 //y=0 \
 //x2=7.575 //y2=1.52
cc_47 ( N_GND_c_3_p N_noxref_4_c_474_n ) capacitor c=0.0114883f //x=6.66 //y=0 \
 //x2=7.575 //y2=1.915
cc_48 ( N_GND_M4_noxref_d N_noxref_4_c_475_n ) capacitor c=0.0131326f //x=7.65 \
 //y=0.865 //x2=7.95 //y2=0.71
cc_49 ( N_GND_M4_noxref_d N_noxref_4_c_476_n ) capacitor c=0.00193127f \
 //x=7.65 //y=0.865 //x2=7.95 //y2=1.365
cc_50 ( N_GND_c_50_p N_noxref_4_c_477_n ) capacitor c=0.00130622f //x=9.82 \
 //y=0 //x2=8.105 //y2=0.865
cc_51 ( N_GND_M4_noxref_d N_noxref_4_c_477_n ) capacitor c=0.00257848f \
 //x=7.65 //y=0.865 //x2=8.105 //y2=0.865
cc_52 ( N_GND_M4_noxref_d N_noxref_4_c_479_n ) capacitor c=0.00255985f \
 //x=7.65 //y=0.865 //x2=8.105 //y2=1.21
cc_53 ( N_GND_c_14_p N_noxref_4_M2_noxref_d ) capacitor c=0.00175924f \
 //x=11.47 //y=0 //x2=4.32 //y2=0.905
cc_54 ( N_GND_c_2_p N_noxref_4_M2_noxref_d ) capacitor c=0.00416273f //x=3.33 \
 //y=0 //x2=4.32 //y2=0.905
cc_55 ( N_GND_c_3_p N_noxref_4_M2_noxref_d ) capacitor c=2.57516e-19 //x=6.66 \
 //y=0 //x2=4.32 //y2=0.905
cc_56 ( N_GND_c_5_p N_noxref_4_M2_noxref_d ) capacitor c=2.31043e-19 //x=11.59 \
 //y=0 //x2=4.32 //y2=0.905
cc_57 ( N_GND_M2_noxref_s N_noxref_4_M2_noxref_d ) capacitor c=0.0769466f \
 //x=3.89 //y=0.365 //x2=4.32 //y2=0.905
cc_58 ( N_GND_c_14_p N_noxref_4_M3_noxref_d ) capacitor c=0.00195394f \
 //x=11.47 //y=0 //x2=5.29 //y2=0.905
cc_59 ( N_GND_c_3_p N_noxref_4_M3_noxref_d ) capacitor c=0.00609243f //x=6.66 \
 //y=0 //x2=5.29 //y2=0.905
cc_60 ( N_GND_c_5_p N_noxref_4_M3_noxref_d ) capacitor c=2.31043e-19 //x=11.59 \
 //y=0 //x2=5.29 //y2=0.905
cc_61 ( N_GND_M2_noxref_s N_noxref_4_M3_noxref_d ) capacitor c=0.0610175f \
 //x=3.89 //y=0.365 //x2=5.29 //y2=0.905
cc_62 ( N_GND_c_62_p N_noxref_5_c_597_n ) capacitor c=2.8021e-19 //x=11.02 \
 //y=0.535 //x2=10.615 //y2=2.59
cc_63 ( N_GND_c_4_p N_noxref_5_c_597_n ) capacitor c=0.0424932f //x=9.99 //y=0 \
 //x2=10.615 //y2=2.59
cc_64 ( N_GND_M6_noxref_s N_noxref_5_c_597_n ) capacitor c=0.00380483f \
 //x=10.485 //y=0.37 //x2=10.615 //y2=2.59
cc_65 ( N_GND_c_4_p N_noxref_5_c_600_n ) capacitor c=9.11674e-19 //x=9.99 \
 //y=0 //x2=9.365 //y2=2.59
cc_66 ( N_GND_c_4_p N_noxref_5_c_601_n ) capacitor c=0.0429465f //x=9.99 //y=0 \
 //x2=9.165 //y2=1.655
cc_67 ( N_GND_M6_noxref_s N_noxref_5_c_601_n ) capacitor c=3.37896e-19 \
 //x=10.485 //y=0.37 //x2=9.165 //y2=1.655
cc_68 ( N_GND_c_3_p N_noxref_5_c_603_n ) capacitor c=9.64732e-19 //x=6.66 \
 //y=0 //x2=9.25 //y2=2.59
cc_69 ( N_GND_c_4_p N_noxref_5_c_603_n ) capacitor c=5.56859e-19 //x=9.99 \
 //y=0 //x2=9.25 //y2=2.59
cc_70 ( N_GND_c_14_p N_noxref_5_c_605_n ) capacitor c=0.00203213f //x=11.47 \
 //y=0 //x2=10.73 //y2=2.085
cc_71 ( N_GND_c_62_p N_noxref_5_c_605_n ) capacitor c=7.79915e-19 //x=11.02 \
 //y=0.535 //x2=10.73 //y2=2.085
cc_72 ( N_GND_c_4_p N_noxref_5_c_605_n ) capacitor c=0.0264037f //x=9.99 //y=0 \
 //x2=10.73 //y2=2.085
cc_73 ( N_GND_c_5_p N_noxref_5_c_605_n ) capacitor c=0.00135052f //x=11.59 \
 //y=0 //x2=10.73 //y2=2.085
cc_74 ( N_GND_M6_noxref_s N_noxref_5_c_605_n ) capacitor c=0.0105356f \
 //x=10.485 //y=0.37 //x2=10.73 //y2=2.085
cc_75 ( N_GND_c_62_p N_noxref_5_c_610_n ) capacitor c=0.0121126f //x=11.02 \
 //y=0.535 //x2=10.84 //y2=0.91
cc_76 ( N_GND_M6_noxref_s N_noxref_5_c_610_n ) capacitor c=0.0317792f \
 //x=10.485 //y=0.37 //x2=10.84 //y2=0.91
cc_77 ( N_GND_c_4_p N_noxref_5_c_612_n ) capacitor c=0.0056248f //x=9.99 //y=0 \
 //x2=10.84 //y2=1.92
cc_78 ( N_GND_M6_noxref_s N_noxref_5_c_613_n ) capacitor c=0.00483274f \
 //x=10.485 //y=0.37 //x2=11.215 //y2=0.755
cc_79 ( N_GND_c_79_p N_noxref_5_c_614_n ) capacitor c=0.0118602f //x=11.505 \
 //y=0.535 //x2=11.37 //y2=0.91
cc_80 ( N_GND_M6_noxref_s N_noxref_5_c_614_n ) capacitor c=0.0143355f \
 //x=10.485 //y=0.37 //x2=11.37 //y2=0.91
cc_81 ( N_GND_M6_noxref_s N_noxref_5_c_616_n ) capacitor c=0.0074042f \
 //x=10.485 //y=0.37 //x2=11.37 //y2=1.255
cc_82 ( N_GND_c_62_p N_noxref_5_c_617_n ) capacitor c=2.1838e-19 //x=11.02 \
 //y=0.535 //x2=10.73 //y2=2.085
cc_83 ( N_GND_c_4_p N_noxref_5_c_617_n ) capacitor c=0.0108179f //x=9.99 //y=0 \
 //x2=10.73 //y2=2.085
cc_84 ( N_GND_M6_noxref_s N_noxref_5_c_617_n ) capacitor c=0.00652238f \
 //x=10.485 //y=0.37 //x2=10.73 //y2=2.085
cc_85 ( N_GND_c_3_p N_noxref_5_M5_noxref_d ) capacitor c=8.58106e-19 //x=6.66 \
 //y=0 //x2=8.62 //y2=0.905
cc_86 ( N_GND_c_4_p N_noxref_5_M5_noxref_d ) capacitor c=0.00616547f //x=9.99 \
 //y=0 //x2=8.62 //y2=0.905
cc_87 ( N_GND_M4_noxref_d N_noxref_5_M5_noxref_d ) capacitor c=0.00143464f \
 //x=7.65 //y=0.865 //x2=8.62 //y2=0.905
cc_88 ( N_GND_M6_noxref_s N_noxref_5_M5_noxref_d ) capacitor c=2.09402e-19 \
 //x=10.485 //y=0.37 //x2=8.62 //y2=0.905
cc_89 ( N_GND_c_1_p N_A_c_723_n ) capacitor c=0.0180518f //x=0.74 //y=0 \
 //x2=1.11 //y2=2.08
cc_90 ( N_GND_c_90_p N_A_c_724_n ) capacitor c=0.00135046f //x=1.095 //y=0 \
 //x2=0.915 //y2=0.865
cc_91 ( N_GND_M0_noxref_d N_A_c_724_n ) capacitor c=0.00220047f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=0.865
cc_92 ( N_GND_M0_noxref_d N_A_c_726_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=1.21
cc_93 ( N_GND_c_1_p N_A_c_727_n ) capacitor c=0.00264481f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.52
cc_94 ( N_GND_c_1_p N_A_c_728_n ) capacitor c=0.0121947f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.915
cc_95 ( N_GND_M0_noxref_d N_A_c_729_n ) capacitor c=0.0131326f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=0.71
cc_96 ( N_GND_M0_noxref_d N_A_c_730_n ) capacitor c=0.00193127f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=1.365
cc_97 ( N_GND_c_97_p N_A_c_731_n ) capacitor c=0.00130622f //x=3.16 //y=0 \
 //x2=1.445 //y2=0.865
cc_98 ( N_GND_M0_noxref_d N_A_c_731_n ) capacitor c=0.00257848f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=0.865
cc_99 ( N_GND_M0_noxref_d N_A_c_733_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=1.21
cc_100 ( N_GND_c_1_p N_B_c_778_n ) capacitor c=9.2064e-19 //x=0.74 //y=0 \
 //x2=1.85 //y2=2.08
cc_101 ( N_GND_c_2_p N_B_c_778_n ) capacitor c=0.00110071f //x=3.33 //y=0 \
 //x2=1.85 //y2=2.08
cc_102 ( N_GND_c_14_p N_noxref_8_c_842_n ) capacitor c=0.00710948f //x=11.47 \
 //y=0 //x2=1.58 //y2=1.58
cc_103 ( N_GND_c_90_p N_noxref_8_c_842_n ) capacitor c=0.00111428f //x=1.095 \
 //y=0 //x2=1.58 //y2=1.58
cc_104 ( N_GND_c_97_p N_noxref_8_c_842_n ) capacitor c=0.00180846f //x=3.16 \
 //y=0 //x2=1.58 //y2=1.58
cc_105 ( N_GND_M0_noxref_d N_noxref_8_c_842_n ) capacitor c=0.0090983f \
 //x=0.99 //y=0.865 //x2=1.58 //y2=1.58
cc_106 ( N_GND_c_14_p N_noxref_8_c_846_n ) capacitor c=0.00723598f //x=11.47 \
 //y=0 //x2=1.665 //y2=0.615
cc_107 ( N_GND_c_97_p N_noxref_8_c_846_n ) capacitor c=0.0146208f //x=3.16 \
 //y=0 //x2=1.665 //y2=0.615
cc_108 ( N_GND_c_5_p N_noxref_8_c_846_n ) capacitor c=0.00145873f //x=11.59 \
 //y=0 //x2=1.665 //y2=0.615
cc_109 ( N_GND_M0_noxref_d N_noxref_8_c_846_n ) capacitor c=0.033812f //x=0.99 \
 //y=0.865 //x2=1.665 //y2=0.615
cc_110 ( N_GND_c_1_p N_noxref_8_c_850_n ) capacitor c=2.91423e-19 //x=0.74 \
 //y=0 //x2=1.665 //y2=1.495
cc_111 ( N_GND_c_14_p N_noxref_8_c_851_n ) capacitor c=0.0199727f //x=11.47 \
 //y=0 //x2=2.55 //y2=0.53
cc_112 ( N_GND_c_97_p N_noxref_8_c_851_n ) capacitor c=0.0371035f //x=3.16 \
 //y=0 //x2=2.55 //y2=0.53
cc_113 ( N_GND_c_5_p N_noxref_8_c_851_n ) capacitor c=0.00199095f //x=11.59 \
 //y=0 //x2=2.55 //y2=0.53
cc_114 ( N_GND_c_14_p N_noxref_8_c_854_n ) capacitor c=0.00719615f //x=11.47 \
 //y=0 //x2=2.635 //y2=0.615
cc_115 ( N_GND_c_97_p N_noxref_8_c_854_n ) capacitor c=0.0144264f //x=3.16 \
 //y=0 //x2=2.635 //y2=0.615
cc_116 ( N_GND_c_116_p N_noxref_8_c_854_n ) capacitor c=9.02073e-19 //x=4.025 \
 //y=0.445 //x2=2.635 //y2=0.615
cc_117 ( N_GND_c_2_p N_noxref_8_c_854_n ) capacitor c=0.0431718f //x=3.33 \
 //y=0 //x2=2.635 //y2=0.615
cc_118 ( N_GND_c_5_p N_noxref_8_c_854_n ) capacitor c=0.00145015f //x=11.59 \
 //y=0 //x2=2.635 //y2=0.615
cc_119 ( N_GND_c_14_p N_noxref_8_M0_noxref_s ) capacitor c=0.00723598f \
 //x=11.47 //y=0 //x2=0.56 //y2=0.365
cc_120 ( N_GND_c_90_p N_noxref_8_M0_noxref_s ) capacitor c=0.0146208f \
 //x=1.095 //y=0 //x2=0.56 //y2=0.365
cc_121 ( N_GND_c_1_p N_noxref_8_M0_noxref_s ) capacitor c=0.0594057f //x=0.74 \
 //y=0 //x2=0.56 //y2=0.365
cc_122 ( N_GND_c_2_p N_noxref_8_M0_noxref_s ) capacitor c=0.00198043f //x=3.33 \
 //y=0 //x2=0.56 //y2=0.365
cc_123 ( N_GND_c_5_p N_noxref_8_M0_noxref_s ) capacitor c=0.00145873f \
 //x=11.59 //y=0 //x2=0.56 //y2=0.365
cc_124 ( N_GND_M0_noxref_d N_noxref_8_M0_noxref_s ) capacitor c=0.0334197f \
 //x=0.99 //y=0.865 //x2=0.56 //y2=0.365
cc_125 ( N_GND_M2_noxref_s N_noxref_8_M0_noxref_s ) capacitor c=9.02073e-19 \
 //x=3.89 //y=0.365 //x2=0.56 //y2=0.365
cc_126 ( N_GND_c_2_p N_C_c_893_n ) capacitor c=0.00112835f //x=3.33 //y=0 \
 //x2=5.18 //y2=2.08
cc_127 ( N_GND_c_3_p N_C_c_893_n ) capacitor c=0.00110071f //x=6.66 //y=0 \
 //x2=5.18 //y2=2.08
cc_128 ( N_GND_c_34_p N_C_c_895_n ) capacitor c=0.0109802f //x=5.395 //y=0.53 \
 //x2=5.215 //y2=0.905
cc_129 ( N_GND_M2_noxref_s N_C_c_895_n ) capacitor c=0.00590563f //x=3.89 \
 //y=0.365 //x2=5.215 //y2=0.905
cc_130 ( N_GND_M2_noxref_s N_C_c_897_n ) capacitor c=0.00466751f //x=3.89 \
 //y=0.365 //x2=5.59 //y2=0.75
cc_131 ( N_GND_M2_noxref_s N_C_c_898_n ) capacitor c=0.00316186f //x=3.89 \
 //y=0.365 //x2=5.59 //y2=1.405
cc_132 ( N_GND_c_37_p N_C_c_899_n ) capacitor c=0.0112321f //x=5.88 //y=0.53 \
 //x2=5.745 //y2=0.905
cc_133 ( N_GND_M2_noxref_s N_C_c_899_n ) capacitor c=0.0142835f //x=3.89 \
 //y=0.365 //x2=5.745 //y2=0.905
cc_134 ( N_GND_c_3_p N_D_c_1007_n ) capacitor c=0.00112835f //x=6.66 //y=0 \
 //x2=8.51 //y2=2.08
cc_135 ( N_GND_c_4_p N_D_c_1007_n ) capacitor c=0.00110071f //x=9.99 //y=0 \
 //x2=8.51 //y2=2.08
cc_136 ( N_GND_c_14_p N_noxref_12_c_1073_n ) capacitor c=0.00708088f //x=11.47 \
 //y=0 //x2=8.24 //y2=1.58
cc_137 ( N_GND_c_43_p N_noxref_12_c_1073_n ) capacitor c=0.00111428f //x=7.755 \
 //y=0 //x2=8.24 //y2=1.58
cc_138 ( N_GND_c_50_p N_noxref_12_c_1073_n ) capacitor c=0.00180846f //x=9.82 \
 //y=0 //x2=8.24 //y2=1.58
cc_139 ( N_GND_M4_noxref_d N_noxref_12_c_1073_n ) capacitor c=0.00880942f \
 //x=7.65 //y=0.865 //x2=8.24 //y2=1.58
cc_140 ( N_GND_c_14_p N_noxref_12_c_1077_n ) capacitor c=0.00723598f //x=11.47 \
 //y=0 //x2=8.325 //y2=0.615
cc_141 ( N_GND_c_50_p N_noxref_12_c_1077_n ) capacitor c=0.0146208f //x=9.82 \
 //y=0 //x2=8.325 //y2=0.615
cc_142 ( N_GND_c_5_p N_noxref_12_c_1077_n ) capacitor c=0.00145873f //x=11.59 \
 //y=0 //x2=8.325 //y2=0.615
cc_143 ( N_GND_M4_noxref_d N_noxref_12_c_1077_n ) capacitor c=0.033812f \
 //x=7.65 //y=0.865 //x2=8.325 //y2=0.615
cc_144 ( N_GND_c_3_p N_noxref_12_c_1081_n ) capacitor c=2.91423e-19 //x=6.66 \
 //y=0 //x2=8.325 //y2=1.495
cc_145 ( N_GND_c_14_p N_noxref_12_c_1082_n ) capacitor c=0.0199727f //x=11.47 \
 //y=0 //x2=9.21 //y2=0.53
cc_146 ( N_GND_c_50_p N_noxref_12_c_1082_n ) capacitor c=0.0371035f //x=9.82 \
 //y=0 //x2=9.21 //y2=0.53
cc_147 ( N_GND_c_5_p N_noxref_12_c_1082_n ) capacitor c=0.00199095f //x=11.59 \
 //y=0 //x2=9.21 //y2=0.53
cc_148 ( N_GND_c_14_p N_noxref_12_c_1085_n ) capacitor c=0.00719615f //x=11.47 \
 //y=0 //x2=9.295 //y2=0.615
cc_149 ( N_GND_c_50_p N_noxref_12_c_1085_n ) capacitor c=0.0144264f //x=9.82 \
 //y=0 //x2=9.295 //y2=0.615
cc_150 ( N_GND_c_150_p N_noxref_12_c_1085_n ) capacitor c=9.77746e-19 \
 //x=10.62 //y=0.45 //x2=9.295 //y2=0.615
cc_151 ( N_GND_c_4_p N_noxref_12_c_1085_n ) capacitor c=0.0431718f //x=9.99 \
 //y=0 //x2=9.295 //y2=0.615
cc_152 ( N_GND_c_5_p N_noxref_12_c_1085_n ) capacitor c=0.00145015f //x=11.59 \
 //y=0 //x2=9.295 //y2=0.615
cc_153 ( N_GND_c_14_p N_noxref_12_M4_noxref_s ) capacitor c=0.00723598f \
 //x=11.47 //y=0 //x2=7.22 //y2=0.365
cc_154 ( N_GND_c_154_p N_noxref_12_M4_noxref_s ) capacitor c=0.00177507f \
 //x=5.965 //y=0.445 //x2=7.22 //y2=0.365
cc_155 ( N_GND_c_43_p N_noxref_12_M4_noxref_s ) capacitor c=0.0146208f \
 //x=7.755 //y=0 //x2=7.22 //y2=0.365
cc_156 ( N_GND_c_3_p N_noxref_12_M4_noxref_s ) capacitor c=0.058339f //x=6.66 \
 //y=0 //x2=7.22 //y2=0.365
cc_157 ( N_GND_c_4_p N_noxref_12_M4_noxref_s ) capacitor c=0.00198098f \
 //x=9.99 //y=0 //x2=7.22 //y2=0.365
cc_158 ( N_GND_c_5_p N_noxref_12_M4_noxref_s ) capacitor c=0.00145873f \
 //x=11.59 //y=0 //x2=7.22 //y2=0.365
cc_159 ( N_GND_M4_noxref_d N_noxref_12_M4_noxref_s ) capacitor c=0.0334197f \
 //x=7.65 //y=0.865 //x2=7.22 //y2=0.365
cc_160 ( N_GND_M6_noxref_s N_noxref_12_M4_noxref_s ) capacitor c=9.77746e-19 \
 //x=10.485 //y=0.37 //x2=7.22 //y2=0.365
cc_161 ( N_GND_c_4_p Y ) capacitor c=9.57726e-19 //x=9.99 //y=0 //x2=11.47 \
 //y2=2.22
cc_162 ( N_GND_c_14_p N_Y_c_1129_n ) capacitor c=0.0021242f //x=11.47 //y=0 \
 //x2=11.385 //y2=2.08
cc_163 ( N_GND_c_5_p N_Y_c_1129_n ) capacitor c=0.029556f //x=11.59 //y=0 \
 //x2=11.385 //y2=2.08
cc_164 ( N_GND_M6_noxref_s N_Y_c_1129_n ) capacitor c=0.00999304f //x=10.485 \
 //y=0.37 //x2=11.385 //y2=2.08
cc_165 ( N_GND_c_14_p N_Y_M6_noxref_d ) capacitor c=0.00194883f //x=11.47 \
 //y=0 //x2=10.915 //y2=0.91
cc_166 ( N_GND_c_62_p N_Y_M6_noxref_d ) capacitor c=0.0146043f //x=11.02 \
 //y=0.535 //x2=10.915 //y2=0.91
cc_167 ( N_GND_c_4_p N_Y_M6_noxref_d ) capacitor c=0.00924905f //x=9.99 //y=0 \
 //x2=10.915 //y2=0.91
cc_168 ( N_GND_c_5_p N_Y_M6_noxref_d ) capacitor c=0.00973758f //x=11.59 //y=0 \
 //x2=10.915 //y2=0.91
cc_169 ( N_GND_M6_noxref_s N_Y_M6_noxref_d ) capacitor c=0.076995f //x=10.485 \
 //y=0.37 //x2=10.915 //y2=0.91
cc_170 ( N_VDD_c_171_n N_noxref_3_c_311_n ) capacitor c=0.00382812f //x=3.33 \
 //y=7.4 //x2=4.325 //y2=2.59
cc_171 ( N_VDD_c_176_p N_noxref_3_c_334_n ) capacitor c=5.76712e-19 //x=1.585 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_172 ( N_VDD_c_177_p N_noxref_3_c_334_n ) capacitor c=5.76712e-19 //x=2.465 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_173 ( N_VDD_M8_noxref_d N_noxref_3_c_334_n ) capacitor c=0.0132775f \
 //x=1.525 //y=5.02 //x2=2.025 //y2=5.2
cc_174 ( N_VDD_c_170_n N_noxref_3_c_337_n ) capacitor c=0.00989999f //x=0.74 \
 //y=7.4 //x2=1.315 //y2=5.2
cc_175 ( N_VDD_M7_noxref_s N_noxref_3_c_337_n ) capacitor c=0.087833f \
 //x=0.655 //y=5.02 //x2=1.315 //y2=5.2
cc_176 ( N_VDD_c_177_p N_noxref_3_c_339_n ) capacitor c=8.71806e-19 //x=2.465 \
 //y=7.4 //x2=2.505 //y2=5.2
cc_177 ( N_VDD_M10_noxref_d N_noxref_3_c_339_n ) capacitor c=0.0167784f \
 //x=2.405 //y=5.02 //x2=2.505 //y2=5.2
cc_178 ( N_VDD_c_170_n N_noxref_3_c_317_n ) capacitor c=0.00159771f //x=0.74 \
 //y=7.4 //x2=2.59 //y2=2.59
cc_179 ( N_VDD_c_171_n N_noxref_3_c_317_n ) capacitor c=0.0462672f //x=3.33 \
 //y=7.4 //x2=2.59 //y2=2.59
cc_180 ( N_VDD_c_171_n N_noxref_3_c_319_n ) capacitor c=0.0103855f //x=3.33 \
 //y=7.4 //x2=4.44 //y2=2.08
cc_181 ( N_VDD_c_171_n N_noxref_3_c_344_n ) capacitor c=0.00860173f //x=3.33 \
 //y=7.4 //x2=4.285 //y2=4.705
cc_182 ( N_VDD_M11_noxref_d N_noxref_3_c_344_n ) capacitor c=2.85008e-19 \
 //x=4.415 //y=5.025 //x2=4.285 //y2=4.705
cc_183 ( N_VDD_c_188_p N_noxref_3_M11_noxref_g ) capacitor c=0.0067918f \
 //x=4.475 //y=7.4 //x2=4.34 //y2=6.025
cc_184 ( N_VDD_c_171_n N_noxref_3_M11_noxref_g ) capacitor c=0.0105272f \
 //x=3.33 //y=7.4 //x2=4.34 //y2=6.025
cc_185 ( N_VDD_M11_noxref_d N_noxref_3_M11_noxref_g ) capacitor c=0.0156786f \
 //x=4.415 //y=5.025 //x2=4.34 //y2=6.025
cc_186 ( N_VDD_c_191_p N_noxref_3_M12_noxref_g ) capacitor c=0.00678153f \
 //x=6.49 //y=7.4 //x2=4.78 //y2=6.025
cc_187 ( N_VDD_M11_noxref_d N_noxref_3_M12_noxref_g ) capacitor c=0.0183011f \
 //x=4.415 //y=5.025 //x2=4.78 //y2=6.025
cc_188 ( N_VDD_c_171_n N_noxref_3_c_351_n ) capacitor c=0.00890932f //x=3.33 \
 //y=7.4 //x2=4.285 //y2=4.705
cc_189 ( N_VDD_c_194_p N_noxref_3_M7_noxref_d ) capacitor c=0.00719513f \
 //x=11.47 //y=7.4 //x2=1.085 //y2=5.02
cc_190 ( N_VDD_c_176_p N_noxref_3_M7_noxref_d ) capacitor c=0.0138103f \
 //x=1.585 //y=7.4 //x2=1.085 //y2=5.02
cc_191 ( N_VDD_c_171_n N_noxref_3_M7_noxref_d ) capacitor c=6.94454e-19 \
 //x=3.33 //y=7.4 //x2=1.085 //y2=5.02
cc_192 ( N_VDD_c_174_n N_noxref_3_M7_noxref_d ) capacitor c=0.00135231f \
 //x=11.47 //y=7.4 //x2=1.085 //y2=5.02
cc_193 ( N_VDD_M8_noxref_d N_noxref_3_M7_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.085 //y2=5.02
cc_194 ( N_VDD_c_194_p N_noxref_3_M9_noxref_d ) capacitor c=0.00719513f \
 //x=11.47 //y=7.4 //x2=1.965 //y2=5.02
cc_195 ( N_VDD_c_177_p N_noxref_3_M9_noxref_d ) capacitor c=0.0138379f \
 //x=2.465 //y=7.4 //x2=1.965 //y2=5.02
cc_196 ( N_VDD_c_171_n N_noxref_3_M9_noxref_d ) capacitor c=0.0120541f \
 //x=3.33 //y=7.4 //x2=1.965 //y2=5.02
cc_197 ( N_VDD_c_174_n N_noxref_3_M9_noxref_d ) capacitor c=0.00135231f \
 //x=11.47 //y=7.4 //x2=1.965 //y2=5.02
cc_198 ( N_VDD_M7_noxref_s N_noxref_3_M9_noxref_d ) capacitor c=0.00111971f \
 //x=0.655 //y=5.02 //x2=1.965 //y2=5.02
cc_199 ( N_VDD_M8_noxref_d N_noxref_3_M9_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.965 //y2=5.02
cc_200 ( N_VDD_M10_noxref_d N_noxref_3_M9_noxref_d ) capacitor c=0.0664752f \
 //x=2.405 //y=5.02 //x2=1.965 //y2=5.02
cc_201 ( N_VDD_c_172_n N_noxref_4_c_455_n ) capacitor c=0.00382812f //x=6.66 \
 //y=7.4 //x2=7.655 //y2=2.59
cc_202 ( N_VDD_c_191_p N_noxref_4_c_490_n ) capacitor c=9.65117e-19 //x=6.49 \
 //y=7.4 //x2=5.835 //y2=5.21
cc_203 ( N_VDD_M15_noxref_s N_noxref_4_c_490_n ) capacitor c=2.47894e-19 \
 //x=7.315 //y=5.02 //x2=5.835 //y2=5.21
cc_204 ( N_VDD_c_171_n N_noxref_4_c_492_n ) capacitor c=8.9933e-19 //x=3.33 \
 //y=7.4 //x2=5.525 //y2=5.21
cc_205 ( N_VDD_c_171_n N_noxref_4_c_467_n ) capacitor c=0.00155409f //x=3.33 \
 //y=7.4 //x2=5.92 //y2=2.59
cc_206 ( N_VDD_c_172_n N_noxref_4_c_467_n ) capacitor c=0.0462858f //x=6.66 \
 //y=7.4 //x2=5.92 //y2=2.59
cc_207 ( N_VDD_c_212_p N_noxref_4_c_469_n ) capacitor c=3.97183e-19 //x=8.245 \
 //y=7.4 //x2=7.77 //y2=2.08
cc_208 ( N_VDD_c_172_n N_noxref_4_c_469_n ) capacitor c=0.0167437f //x=6.66 \
 //y=7.4 //x2=7.77 //y2=2.08
cc_209 ( N_VDD_c_212_p N_noxref_4_M15_noxref_g ) capacitor c=0.00726866f \
 //x=8.245 //y=7.4 //x2=7.67 //y2=6.02
cc_210 ( N_VDD_M15_noxref_s N_noxref_4_M15_noxref_g ) capacitor c=0.054195f \
 //x=7.315 //y=5.02 //x2=7.67 //y2=6.02
cc_211 ( N_VDD_c_212_p N_noxref_4_M16_noxref_g ) capacitor c=0.00672952f \
 //x=8.245 //y=7.4 //x2=8.11 //y2=6.02
cc_212 ( N_VDD_M16_noxref_d N_noxref_4_M16_noxref_g ) capacitor c=0.015318f \
 //x=8.185 //y=5.02 //x2=8.11 //y2=6.02
cc_213 ( N_VDD_c_172_n N_noxref_4_c_501_n ) capacitor c=0.0162221f //x=6.66 \
 //y=7.4 //x2=7.77 //y2=4.7
cc_214 ( N_VDD_c_172_n N_noxref_4_M13_noxref_d ) capacitor c=0.00966019f \
 //x=6.66 //y=7.4 //x2=5.295 //y2=5.025
cc_215 ( N_VDD_M11_noxref_d N_noxref_4_M13_noxref_d ) capacitor c=0.00561178f \
 //x=4.415 //y=5.025 //x2=5.295 //y2=5.025
cc_216 ( N_VDD_M15_noxref_s N_noxref_4_M13_noxref_d ) capacitor c=4.37644e-19 \
 //x=7.315 //y=5.02 //x2=5.295 //y2=5.025
cc_217 ( N_VDD_c_173_n N_noxref_5_c_597_n ) capacitor c=0.00382812f //x=9.99 \
 //y=7.4 //x2=10.615 //y2=2.59
cc_218 ( N_VDD_c_212_p N_noxref_5_c_625_n ) capacitor c=5.76712e-19 //x=8.245 \
 //y=7.4 //x2=8.685 //y2=5.2
cc_219 ( N_VDD_c_224_p N_noxref_5_c_625_n ) capacitor c=5.76712e-19 //x=9.125 \
 //y=7.4 //x2=8.685 //y2=5.2
cc_220 ( N_VDD_M16_noxref_d N_noxref_5_c_625_n ) capacitor c=0.0132775f \
 //x=8.185 //y=5.02 //x2=8.685 //y2=5.2
cc_221 ( N_VDD_c_172_n N_noxref_5_c_628_n ) capacitor c=0.00985474f //x=6.66 \
 //y=7.4 //x2=7.975 //y2=5.2
cc_222 ( N_VDD_M15_noxref_s N_noxref_5_c_628_n ) capacitor c=0.087833f \
 //x=7.315 //y=5.02 //x2=7.975 //y2=5.2
cc_223 ( N_VDD_c_224_p N_noxref_5_c_630_n ) capacitor c=8.71806e-19 //x=9.125 \
 //y=7.4 //x2=9.165 //y2=5.2
cc_224 ( N_VDD_M18_noxref_d N_noxref_5_c_630_n ) capacitor c=0.0167784f \
 //x=9.065 //y=5.02 //x2=9.165 //y2=5.2
cc_225 ( N_VDD_c_172_n N_noxref_5_c_603_n ) capacitor c=0.00151618f //x=6.66 \
 //y=7.4 //x2=9.25 //y2=2.59
cc_226 ( N_VDD_c_173_n N_noxref_5_c_603_n ) capacitor c=0.0461201f //x=9.99 \
 //y=7.4 //x2=9.25 //y2=2.59
cc_227 ( N_VDD_c_173_n N_noxref_5_c_605_n ) capacitor c=0.0272885f //x=9.99 \
 //y=7.4 //x2=10.73 //y2=2.085
cc_228 ( N_VDD_c_174_n N_noxref_5_c_605_n ) capacitor c=0.00144809f //x=11.47 \
 //y=7.4 //x2=10.73 //y2=2.085
cc_229 ( N_VDD_M19_noxref_s N_noxref_5_c_605_n ) capacitor c=0.00938034f \
 //x=10.53 //y=5.02 //x2=10.73 //y2=2.085
cc_230 ( N_VDD_c_235_p N_noxref_5_M19_noxref_g ) capacitor c=0.00748034f \
 //x=11.46 //y=7.4 //x2=10.885 //y2=6.02
cc_231 ( N_VDD_c_173_n N_noxref_5_M19_noxref_g ) capacitor c=0.00895557f \
 //x=9.99 //y=7.4 //x2=10.885 //y2=6.02
cc_232 ( N_VDD_M19_noxref_s N_noxref_5_M19_noxref_g ) capacitor c=0.0528676f \
 //x=10.53 //y=5.02 //x2=10.885 //y2=6.02
cc_233 ( N_VDD_c_235_p N_noxref_5_M20_noxref_g ) capacitor c=0.00697478f \
 //x=11.46 //y=7.4 //x2=11.325 //y2=6.02
cc_234 ( N_VDD_M20_noxref_d N_noxref_5_M20_noxref_g ) capacitor c=0.0528676f \
 //x=11.4 //y=5.02 //x2=11.325 //y2=6.02
cc_235 ( N_VDD_c_174_n N_noxref_5_c_642_n ) capacitor c=0.0287802f //x=11.47 \
 //y=7.4 //x2=11.25 //y2=4.79
cc_236 ( N_VDD_c_173_n N_noxref_5_c_643_n ) capacitor c=0.011132f //x=9.99 \
 //y=7.4 //x2=10.96 //y2=4.79
cc_237 ( N_VDD_M19_noxref_s N_noxref_5_c_643_n ) capacitor c=0.00665831f \
 //x=10.53 //y=5.02 //x2=10.96 //y2=4.79
cc_238 ( N_VDD_c_194_p N_noxref_5_M15_noxref_d ) capacitor c=0.00719513f \
 //x=11.47 //y=7.4 //x2=7.745 //y2=5.02
cc_239 ( N_VDD_c_212_p N_noxref_5_M15_noxref_d ) capacitor c=0.0138103f \
 //x=8.245 //y=7.4 //x2=7.745 //y2=5.02
cc_240 ( N_VDD_c_173_n N_noxref_5_M15_noxref_d ) capacitor c=6.94454e-19 \
 //x=9.99 //y=7.4 //x2=7.745 //y2=5.02
cc_241 ( N_VDD_c_174_n N_noxref_5_M15_noxref_d ) capacitor c=0.00135231f \
 //x=11.47 //y=7.4 //x2=7.745 //y2=5.02
cc_242 ( N_VDD_M16_noxref_d N_noxref_5_M15_noxref_d ) capacitor c=0.0664752f \
 //x=8.185 //y=5.02 //x2=7.745 //y2=5.02
cc_243 ( N_VDD_c_194_p N_noxref_5_M17_noxref_d ) capacitor c=0.00719513f \
 //x=11.47 //y=7.4 //x2=8.625 //y2=5.02
cc_244 ( N_VDD_c_224_p N_noxref_5_M17_noxref_d ) capacitor c=0.0138379f \
 //x=9.125 //y=7.4 //x2=8.625 //y2=5.02
cc_245 ( N_VDD_c_173_n N_noxref_5_M17_noxref_d ) capacitor c=0.0120541f \
 //x=9.99 //y=7.4 //x2=8.625 //y2=5.02
cc_246 ( N_VDD_c_174_n N_noxref_5_M17_noxref_d ) capacitor c=0.00135231f \
 //x=11.47 //y=7.4 //x2=8.625 //y2=5.02
cc_247 ( N_VDD_M15_noxref_s N_noxref_5_M17_noxref_d ) capacitor c=0.00111971f \
 //x=7.315 //y=5.02 //x2=8.625 //y2=5.02
cc_248 ( N_VDD_M16_noxref_d N_noxref_5_M17_noxref_d ) capacitor c=0.0664752f \
 //x=8.185 //y=5.02 //x2=8.625 //y2=5.02
cc_249 ( N_VDD_M18_noxref_d N_noxref_5_M17_noxref_d ) capacitor c=0.0664752f \
 //x=9.065 //y=5.02 //x2=8.625 //y2=5.02
cc_250 ( N_VDD_M19_noxref_s N_noxref_5_M17_noxref_d ) capacitor c=5.1407e-19 \
 //x=10.53 //y=5.02 //x2=8.625 //y2=5.02
cc_251 ( N_VDD_c_176_p N_A_c_723_n ) capacitor c=3.97183e-19 //x=1.585 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_252 ( N_VDD_c_170_n N_A_c_723_n ) capacitor c=0.016845f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_253 ( N_VDD_c_176_p N_A_M7_noxref_g ) capacitor c=0.00726866f //x=1.585 \
 //y=7.4 //x2=1.01 //y2=6.02
cc_254 ( N_VDD_M7_noxref_s N_A_M7_noxref_g ) capacitor c=0.054195f //x=0.655 \
 //y=5.02 //x2=1.01 //y2=6.02
cc_255 ( N_VDD_c_176_p N_A_M8_noxref_g ) capacitor c=0.00672952f //x=1.585 \
 //y=7.4 //x2=1.45 //y2=6.02
cc_256 ( N_VDD_M8_noxref_d N_A_M8_noxref_g ) capacitor c=0.015318f //x=1.525 \
 //y=5.02 //x2=1.45 //y2=6.02
cc_257 ( N_VDD_c_170_n N_A_c_740_n ) capacitor c=0.0292267f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=4.7
cc_258 ( N_VDD_c_170_n N_B_c_778_n ) capacitor c=6.61004e-19 //x=0.74 //y=7.4 \
 //x2=1.85 //y2=2.08
cc_259 ( N_VDD_c_171_n N_B_c_778_n ) capacitor c=6.09526e-19 //x=3.33 //y=7.4 \
 //x2=1.85 //y2=2.08
cc_260 ( N_VDD_c_177_p N_B_M9_noxref_g ) capacitor c=0.00673971f //x=2.465 \
 //y=7.4 //x2=1.89 //y2=6.02
cc_261 ( N_VDD_M8_noxref_d N_B_M9_noxref_g ) capacitor c=0.015318f //x=1.525 \
 //y=5.02 //x2=1.89 //y2=6.02
cc_262 ( N_VDD_c_177_p N_B_M10_noxref_g ) capacitor c=0.00672952f //x=2.465 \
 //y=7.4 //x2=2.33 //y2=6.02
cc_263 ( N_VDD_c_171_n N_B_M10_noxref_g ) capacitor c=0.00954586f //x=3.33 \
 //y=7.4 //x2=2.33 //y2=6.02
cc_264 ( N_VDD_M10_noxref_d N_B_M10_noxref_g ) capacitor c=0.0430452f \
 //x=2.405 //y=5.02 //x2=2.33 //y2=6.02
cc_265 ( N_VDD_c_171_n N_C_c_893_n ) capacitor c=7.02327e-19 //x=3.33 //y=7.4 \
 //x2=5.18 //y2=2.08
cc_266 ( N_VDD_c_172_n N_C_c_893_n ) capacitor c=6.16704e-19 //x=6.66 //y=7.4 \
 //x2=5.18 //y2=2.08
cc_267 ( N_VDD_c_191_p N_C_M13_noxref_g ) capacitor c=0.00513565f //x=6.49 \
 //y=7.4 //x2=5.22 //y2=6.025
cc_268 ( N_VDD_c_191_p N_C_M14_noxref_g ) capacitor c=0.00512552f //x=6.49 \
 //y=7.4 //x2=5.66 //y2=6.025
cc_269 ( N_VDD_c_172_n N_C_M14_noxref_g ) capacitor c=0.0116195f //x=6.66 \
 //y=7.4 //x2=5.66 //y2=6.025
cc_270 ( N_VDD_c_188_p N_noxref_10_c_964_n ) capacitor c=5.81484e-19 //x=4.475 \
 //y=7.4 //x2=4.915 //y2=5.21
cc_271 ( N_VDD_c_191_p N_noxref_10_c_964_n ) capacitor c=5.81484e-19 //x=6.49 \
 //y=7.4 //x2=4.915 //y2=5.21
cc_272 ( N_VDD_c_172_n N_noxref_10_c_964_n ) capacitor c=0.00289291f //x=6.66 \
 //y=7.4 //x2=4.915 //y2=5.21
cc_273 ( N_VDD_M11_noxref_d N_noxref_10_c_964_n ) capacitor c=0.0132432f \
 //x=4.415 //y=5.025 //x2=4.915 //y2=5.21
cc_274 ( N_VDD_c_171_n N_noxref_10_c_968_n ) capacitor c=0.0669114f //x=3.33 \
 //y=7.4 //x2=4.205 //y2=5.21
cc_275 ( N_VDD_c_174_n N_noxref_10_c_969_n ) capacitor c=0.00360102f //x=11.47 \
 //y=7.4 //x2=5.795 //y2=6.91
cc_276 ( N_VDD_c_194_p N_noxref_10_c_970_n ) capacitor c=0.0370274f //x=11.47 \
 //y=7.4 //x2=5.085 //y2=6.91
cc_277 ( N_VDD_c_191_p N_noxref_10_c_970_n ) capacitor c=0.0586694f //x=6.49 \
 //y=7.4 //x2=5.085 //y2=6.91
cc_278 ( N_VDD_c_174_n N_noxref_10_c_970_n ) capacitor c=0.00118659f //x=11.47 \
 //y=7.4 //x2=5.085 //y2=6.91
cc_279 ( N_VDD_c_194_p N_noxref_10_M11_noxref_s ) capacitor c=0.00726388f \
 //x=11.47 //y=7.4 //x2=3.985 //y2=5.025
cc_280 ( N_VDD_c_188_p N_noxref_10_M11_noxref_s ) capacitor c=0.0141117f \
 //x=4.475 //y=7.4 //x2=3.985 //y2=5.025
cc_281 ( N_VDD_c_174_n N_noxref_10_M11_noxref_s ) capacitor c=0.00138926f \
 //x=11.47 //y=7.4 //x2=3.985 //y2=5.025
cc_282 ( N_VDD_M10_noxref_d N_noxref_10_M11_noxref_s ) capacitor c=0.00196306f \
 //x=2.405 //y=5.02 //x2=3.985 //y2=5.025
cc_283 ( N_VDD_M11_noxref_d N_noxref_10_M11_noxref_s ) capacitor c=0.0667021f \
 //x=4.415 //y=5.025 //x2=3.985 //y2=5.025
cc_284 ( N_VDD_c_171_n N_noxref_10_M12_noxref_d ) capacitor c=8.88629e-19 \
 //x=3.33 //y=7.4 //x2=4.855 //y2=5.025
cc_285 ( N_VDD_M11_noxref_d N_noxref_10_M12_noxref_d ) capacitor c=0.0659925f \
 //x=4.415 //y=5.025 //x2=4.855 //y2=5.025
cc_286 ( N_VDD_c_172_n N_noxref_10_M14_noxref_d ) capacitor c=0.0520312f \
 //x=6.66 //y=7.4 //x2=5.735 //y2=5.025
cc_287 ( N_VDD_M11_noxref_d N_noxref_10_M14_noxref_d ) capacitor c=0.00107819f \
 //x=4.415 //y=5.025 //x2=5.735 //y2=5.025
cc_288 ( N_VDD_M15_noxref_s N_noxref_10_M14_noxref_d ) capacitor c=0.00195151f \
 //x=7.315 //y=5.02 //x2=5.735 //y2=5.025
cc_289 ( N_VDD_c_172_n N_D_c_1007_n ) capacitor c=6.61004e-19 //x=6.66 //y=7.4 \
 //x2=8.51 //y2=2.08
cc_290 ( N_VDD_c_173_n N_D_c_1007_n ) capacitor c=6.09526e-19 //x=9.99 //y=7.4 \
 //x2=8.51 //y2=2.08
cc_291 ( N_VDD_c_224_p N_D_M17_noxref_g ) capacitor c=0.00673971f //x=9.125 \
 //y=7.4 //x2=8.55 //y2=6.02
cc_292 ( N_VDD_M16_noxref_d N_D_M17_noxref_g ) capacitor c=0.015318f //x=8.185 \
 //y=5.02 //x2=8.55 //y2=6.02
cc_293 ( N_VDD_c_224_p N_D_M18_noxref_g ) capacitor c=0.00672952f //x=9.125 \
 //y=7.4 //x2=8.99 //y2=6.02
cc_294 ( N_VDD_c_173_n N_D_M18_noxref_g ) capacitor c=0.00904525f //x=9.99 \
 //y=7.4 //x2=8.99 //y2=6.02
cc_295 ( N_VDD_M18_noxref_d N_D_M18_noxref_g ) capacitor c=0.0430452f \
 //x=9.065 //y=5.02 //x2=8.99 //y2=6.02
cc_296 ( N_VDD_c_173_n Y ) capacitor c=4.80934e-19 //x=9.99 //y=7.4 //x2=11.47 \
 //y2=2.22
cc_297 ( N_VDD_c_174_n Y ) capacitor c=0.0232778f //x=11.47 //y=7.4 //x2=11.47 \
 //y2=2.22
cc_298 ( N_VDD_c_235_p N_Y_c_1139_n ) capacitor c=8.92854e-19 //x=11.46 \
 //y=7.4 //x2=11.385 //y2=4.58
cc_299 ( N_VDD_M20_noxref_d N_Y_c_1139_n ) capacitor c=0.00644908f //x=11.4 \
 //y=5.02 //x2=11.385 //y2=4.58
cc_300 ( N_VDD_c_173_n N_Y_c_1141_n ) capacitor c=0.017572f //x=9.99 //y=7.4 \
 //x2=11.19 //y2=4.58
cc_301 ( N_VDD_c_194_p N_Y_M19_noxref_d ) capacitor c=0.00722811f //x=11.47 \
 //y=7.4 //x2=10.96 //y2=5.02
cc_302 ( N_VDD_c_235_p N_Y_M19_noxref_d ) capacitor c=0.0139004f //x=11.46 \
 //y=7.4 //x2=10.96 //y2=5.02
cc_303 ( N_VDD_c_174_n N_Y_M19_noxref_d ) capacitor c=0.0219131f //x=11.47 \
 //y=7.4 //x2=10.96 //y2=5.02
cc_304 ( N_VDD_M19_noxref_s N_Y_M19_noxref_d ) capacitor c=0.0843065f \
 //x=10.53 //y=5.02 //x2=10.96 //y2=5.02
cc_305 ( N_VDD_M20_noxref_d N_Y_M19_noxref_d ) capacitor c=0.0832641f //x=11.4 \
 //y=5.02 //x2=10.96 //y2=5.02
cc_306 ( N_noxref_3_c_311_n N_noxref_4_c_457_n ) capacitor c=0.0114841f \
 //x=4.325 //y=2.59 //x2=6.035 //y2=2.59
cc_307 ( N_noxref_3_c_329_n N_noxref_4_c_459_n ) capacitor c=0.00431513f \
 //x=4.775 //y=1.25 //x2=5.395 //y2=1.655
cc_308 ( N_noxref_3_c_311_n N_noxref_4_c_507_n ) capacitor c=0.0018301f \
 //x=4.325 //y=2.59 //x2=4.595 //y2=1.655
cc_309 ( N_noxref_3_c_319_n N_noxref_4_c_507_n ) capacitor c=0.0107041f \
 //x=4.44 //y=2.08 //x2=4.595 //y2=1.655
cc_310 ( N_noxref_3_c_324_n N_noxref_4_c_507_n ) capacitor c=0.00524371f \
 //x=4.245 //y=1.915 //x2=4.595 //y2=1.655
cc_311 ( N_noxref_3_c_317_n N_noxref_4_c_467_n ) capacitor c=3.55699e-19 \
 //x=2.59 //y=2.59 //x2=5.92 //y2=2.59
cc_312 ( N_noxref_3_c_319_n N_noxref_4_c_467_n ) capacitor c=0.00354085f \
 //x=4.44 //y=2.08 //x2=5.92 //y2=2.59
cc_313 ( N_noxref_3_c_322_n N_noxref_4_M2_noxref_d ) capacitor c=0.0013184f \
 //x=4.245 //y=0.905 //x2=4.32 //y2=0.905
cc_314 ( N_noxref_3_c_372_p N_noxref_4_M2_noxref_d ) capacitor c=0.0034598f \
 //x=4.245 //y=1.25 //x2=4.32 //y2=0.905
cc_315 ( N_noxref_3_c_373_p N_noxref_4_M2_noxref_d ) capacitor c=0.00300148f \
 //x=4.245 //y=1.56 //x2=4.32 //y2=0.905
cc_316 ( N_noxref_3_c_324_n N_noxref_4_M2_noxref_d ) capacitor c=0.00273686f \
 //x=4.245 //y=1.915 //x2=4.32 //y2=0.905
cc_317 ( N_noxref_3_c_326_n N_noxref_4_M2_noxref_d ) capacitor c=0.00241102f \
 //x=4.62 //y=0.75 //x2=4.32 //y2=0.905
cc_318 ( N_noxref_3_c_376_p N_noxref_4_M2_noxref_d ) capacitor c=0.0123304f \
 //x=4.62 //y=1.405 //x2=4.32 //y2=0.905
cc_319 ( N_noxref_3_c_327_n N_noxref_4_M2_noxref_d ) capacitor c=0.00219619f \
 //x=4.775 //y=0.905 //x2=4.32 //y2=0.905
cc_320 ( N_noxref_3_c_329_n N_noxref_4_M2_noxref_d ) capacitor c=0.00603828f \
 //x=4.775 //y=1.25 //x2=4.32 //y2=0.905
cc_321 ( N_noxref_3_c_337_n N_A_c_723_n ) capacitor c=0.0055959f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=2.08
cc_322 ( N_noxref_3_c_317_n N_A_c_723_n ) capacitor c=0.00407922f //x=2.59 \
 //y=2.59 //x2=1.11 //y2=2.08
cc_323 ( N_noxref_3_c_337_n N_A_M7_noxref_g ) capacitor c=0.0177326f //x=1.315 \
 //y=5.2 //x2=1.01 //y2=6.02
cc_324 ( N_noxref_3_c_334_n N_A_M8_noxref_g ) capacitor c=0.0204115f //x=2.025 \
 //y=5.2 //x2=1.45 //y2=6.02
cc_325 ( N_noxref_3_M7_noxref_d N_A_M8_noxref_g ) capacitor c=0.0173476f \
 //x=1.085 //y=5.02 //x2=1.45 //y2=6.02
cc_326 ( N_noxref_3_c_337_n N_A_c_740_n ) capacitor c=0.00605692f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=4.7
cc_327 ( N_noxref_3_c_334_n N_B_c_787_n ) capacitor c=0.0127867f //x=2.025 \
 //y=5.2 //x2=1.85 //y2=4.535
cc_328 ( N_noxref_3_c_317_n N_B_c_787_n ) capacitor c=0.0101284f //x=2.59 \
 //y=2.59 //x2=1.85 //y2=4.535
cc_329 ( N_noxref_3_c_314_n N_B_c_778_n ) capacitor c=0.00732168f //x=2.705 \
 //y=2.59 //x2=1.85 //y2=2.08
cc_330 ( N_noxref_3_c_317_n N_B_c_778_n ) capacitor c=0.0813981f //x=2.59 \
 //y=2.59 //x2=1.85 //y2=2.08
cc_331 ( N_noxref_3_c_319_n N_B_c_778_n ) capacitor c=9.8819e-19 //x=4.44 \
 //y=2.08 //x2=1.85 //y2=2.08
cc_332 ( N_noxref_3_c_334_n N_B_M9_noxref_g ) capacitor c=0.0166699f //x=2.025 \
 //y=5.2 //x2=1.89 //y2=6.02
cc_333 ( N_noxref_3_M9_noxref_d N_B_M9_noxref_g ) capacitor c=0.0173477f \
 //x=1.965 //y=5.02 //x2=1.89 //y2=6.02
cc_334 ( N_noxref_3_c_339_n N_B_M10_noxref_g ) capacitor c=0.0223814f \
 //x=2.505 //y=5.2 //x2=2.33 //y2=6.02
cc_335 ( N_noxref_3_M9_noxref_d N_B_M10_noxref_g ) capacitor c=0.0179769f \
 //x=1.965 //y=5.02 //x2=2.33 //y2=6.02
cc_336 ( N_noxref_3_M1_noxref_d N_B_c_796_n ) capacitor c=0.00217566f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=0.905
cc_337 ( N_noxref_3_M1_noxref_d N_B_c_797_n ) capacitor c=0.0034598f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.25
cc_338 ( N_noxref_3_M1_noxref_d N_B_c_798_n ) capacitor c=0.0065582f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.56
cc_339 ( N_noxref_3_c_317_n N_B_c_799_n ) capacitor c=0.0142673f //x=2.59 \
 //y=2.59 //x2=2.255 //y2=4.79
cc_340 ( N_noxref_3_c_398_p N_B_c_799_n ) capacitor c=0.00421574f //x=2.11 \
 //y=5.2 //x2=2.255 //y2=4.79
cc_341 ( N_noxref_3_M1_noxref_d N_B_c_801_n ) capacitor c=0.00241102f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=0.75
cc_342 ( N_noxref_3_c_315_n N_B_c_802_n ) capacitor c=0.00359704f //x=2.505 \
 //y=1.655 //x2=2.26 //y2=1.405
cc_343 ( N_noxref_3_M1_noxref_d N_B_c_802_n ) capacitor c=0.0138845f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=1.405
cc_344 ( N_noxref_3_M1_noxref_d N_B_c_804_n ) capacitor c=0.00132245f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=0.905
cc_345 ( N_noxref_3_c_315_n N_B_c_805_n ) capacitor c=0.00457401f //x=2.505 \
 //y=1.655 //x2=2.415 //y2=1.25
cc_346 ( N_noxref_3_M1_noxref_d N_B_c_805_n ) capacitor c=0.00566463f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=1.25
cc_347 ( N_noxref_3_c_317_n N_B_c_807_n ) capacitor c=0.00877984f //x=2.59 \
 //y=2.59 //x2=1.85 //y2=2.08
cc_348 ( N_noxref_3_c_317_n N_B_c_808_n ) capacitor c=0.00306024f //x=2.59 \
 //y=2.59 //x2=1.85 //y2=1.915
cc_349 ( N_noxref_3_M1_noxref_d N_B_c_808_n ) capacitor c=0.00660593f //x=1.96 \
 //y=0.905 //x2=1.85 //y2=1.915
cc_350 ( N_noxref_3_c_334_n N_B_c_810_n ) capacitor c=0.00399417f //x=2.025 \
 //y=5.2 //x2=1.88 //y2=4.7
cc_351 ( N_noxref_3_c_317_n N_B_c_810_n ) capacitor c=0.00533692f //x=2.59 \
 //y=2.59 //x2=1.88 //y2=4.7
cc_352 ( N_noxref_3_c_410_p N_noxref_8_c_866_n ) capacitor c=3.15806e-19 \
 //x=2.235 //y=1.655 //x2=0.695 //y2=1.495
cc_353 ( N_noxref_3_c_410_p N_noxref_8_c_850_n ) capacitor c=0.0201674f \
 //x=2.235 //y=1.655 //x2=1.665 //y2=1.495
cc_354 ( N_noxref_3_c_315_n N_noxref_8_c_851_n ) capacitor c=0.00468333f \
 //x=2.505 //y=1.655 //x2=2.55 //y2=0.53
cc_355 ( N_noxref_3_M1_noxref_d N_noxref_8_c_851_n ) capacitor c=0.0118355f \
 //x=1.96 //y=0.905 //x2=2.55 //y2=0.53
cc_356 ( N_noxref_3_c_311_n N_noxref_8_M0_noxref_s ) capacitor c=3.03583e-19 \
 //x=4.325 //y=2.59 //x2=0.56 //y2=0.365
cc_357 ( N_noxref_3_c_314_n N_noxref_8_M0_noxref_s ) capacitor c=6.92363e-19 \
 //x=2.705 //y=2.59 //x2=0.56 //y2=0.365
cc_358 ( N_noxref_3_c_315_n N_noxref_8_M0_noxref_s ) capacitor c=0.0129465f \
 //x=2.505 //y=1.655 //x2=0.56 //y2=0.365
cc_359 ( N_noxref_3_M1_noxref_d N_noxref_8_M0_noxref_s ) capacitor \
 c=0.0437911f //x=1.96 //y=0.905 //x2=0.56 //y2=0.365
cc_360 ( N_noxref_3_c_344_n N_C_c_906_n ) capacitor c=0.0470738f //x=4.285 \
 //y=4.705 //x2=5.18 //y2=4.54
cc_361 ( N_noxref_3_c_419_p N_C_c_906_n ) capacitor c=0.00146509f //x=4.705 \
 //y=4.795 //x2=5.18 //y2=4.54
cc_362 ( N_noxref_3_c_351_n N_C_c_906_n ) capacitor c=0.00112871f //x=4.285 \
 //y=4.705 //x2=5.18 //y2=4.54
cc_363 ( N_noxref_3_c_311_n N_C_c_893_n ) capacitor c=0.00316948f //x=4.325 \
 //y=2.59 //x2=5.18 //y2=2.08
cc_364 ( N_noxref_3_c_317_n N_C_c_893_n ) capacitor c=9.8819e-19 //x=2.59 \
 //y=2.59 //x2=5.18 //y2=2.08
cc_365 ( N_noxref_3_c_319_n N_C_c_893_n ) capacitor c=0.0447305f //x=4.44 \
 //y=2.08 //x2=5.18 //y2=2.08
cc_366 ( N_noxref_3_c_324_n N_C_c_893_n ) capacitor c=0.00308814f //x=4.245 \
 //y=1.915 //x2=5.18 //y2=2.08
cc_367 ( N_noxref_3_M11_noxref_g N_C_M13_noxref_g ) capacitor c=0.0100243f \
 //x=4.34 //y=6.025 //x2=5.22 //y2=6.025
cc_368 ( N_noxref_3_M12_noxref_g N_C_M13_noxref_g ) capacitor c=0.107798f \
 //x=4.78 //y=6.025 //x2=5.22 //y2=6.025
cc_369 ( N_noxref_3_M12_noxref_g N_C_M14_noxref_g ) capacitor c=0.0094155f \
 //x=4.78 //y=6.025 //x2=5.66 //y2=6.025
cc_370 ( N_noxref_3_c_322_n N_C_c_895_n ) capacitor c=0.00125788f //x=4.245 \
 //y=0.905 //x2=5.215 //y2=0.905
cc_371 ( N_noxref_3_c_327_n N_C_c_895_n ) capacitor c=0.0126654f //x=4.775 \
 //y=0.905 //x2=5.215 //y2=0.905
cc_372 ( N_noxref_3_c_372_p N_C_c_918_n ) capacitor c=0.00148539f //x=4.245 \
 //y=1.25 //x2=5.215 //y2=1.255
cc_373 ( N_noxref_3_c_373_p N_C_c_918_n ) capacitor c=0.00105591f //x=4.245 \
 //y=1.56 //x2=5.215 //y2=1.255
cc_374 ( N_noxref_3_c_329_n N_C_c_918_n ) capacitor c=0.0126654f //x=4.775 \
 //y=1.25 //x2=5.215 //y2=1.255
cc_375 ( N_noxref_3_c_373_p N_C_c_921_n ) capacitor c=0.00109549f //x=4.245 \
 //y=1.56 //x2=5.215 //y2=1.56
cc_376 ( N_noxref_3_c_329_n N_C_c_921_n ) capacitor c=0.00886999f //x=4.775 \
 //y=1.25 //x2=5.215 //y2=1.56
cc_377 ( N_noxref_3_c_329_n N_C_c_898_n ) capacitor c=0.00123863f //x=4.775 \
 //y=1.25 //x2=5.59 //y2=1.405
cc_378 ( N_noxref_3_c_327_n N_C_c_899_n ) capacitor c=0.00132934f //x=4.775 \
 //y=0.905 //x2=5.745 //y2=0.905
cc_379 ( N_noxref_3_c_329_n N_C_c_925_n ) capacitor c=0.00150734f //x=4.775 \
 //y=1.25 //x2=5.745 //y2=1.255
cc_380 ( N_noxref_3_c_319_n N_C_c_926_n ) capacitor c=0.00307062f //x=4.44 \
 //y=2.08 //x2=5.18 //y2=2.08
cc_381 ( N_noxref_3_c_324_n N_C_c_926_n ) capacitor c=0.0179092f //x=4.245 \
 //y=1.915 //x2=5.18 //y2=2.08
cc_382 ( N_noxref_3_c_324_n N_C_c_928_n ) capacitor c=0.00577193f //x=4.245 \
 //y=1.915 //x2=5.18 //y2=1.915
cc_383 ( N_noxref_3_c_344_n N_C_c_929_n ) capacitor c=0.00336963f //x=4.285 \
 //y=4.705 //x2=5.215 //y2=4.705
cc_384 ( N_noxref_3_c_419_p N_C_c_929_n ) capacitor c=0.020271f //x=4.705 \
 //y=4.795 //x2=5.215 //y2=4.705
cc_385 ( N_noxref_3_c_351_n N_C_c_929_n ) capacitor c=0.00546725f //x=4.285 \
 //y=4.705 //x2=5.215 //y2=4.705
cc_386 ( N_noxref_3_c_344_n N_noxref_10_c_964_n ) capacitor c=0.00630079f \
 //x=4.285 //y=4.705 //x2=4.915 //y2=5.21
cc_387 ( N_noxref_3_M11_noxref_g N_noxref_10_c_964_n ) capacitor c=0.0182669f \
 //x=4.34 //y=6.025 //x2=4.915 //y2=5.21
cc_388 ( N_noxref_3_M12_noxref_g N_noxref_10_c_964_n ) capacitor c=0.0204082f \
 //x=4.78 //y=6.025 //x2=4.915 //y2=5.21
cc_389 ( N_noxref_3_c_419_p N_noxref_10_c_964_n ) capacitor c=0.00365818f \
 //x=4.705 //y=4.795 //x2=4.915 //y2=5.21
cc_390 ( N_noxref_3_c_351_n N_noxref_10_c_964_n ) capacitor c=0.0017421f \
 //x=4.285 //y=4.705 //x2=4.915 //y2=5.21
cc_391 ( N_noxref_3_c_339_n N_noxref_10_c_968_n ) capacitor c=2.87761e-19 \
 //x=2.505 //y=5.2 //x2=4.205 //y2=5.21
cc_392 ( N_noxref_3_c_344_n N_noxref_10_c_968_n ) capacitor c=0.0118415f \
 //x=4.285 //y=4.705 //x2=4.205 //y2=5.21
cc_393 ( N_noxref_3_c_351_n N_noxref_10_c_968_n ) capacitor c=0.00613395f \
 //x=4.285 //y=4.705 //x2=4.205 //y2=5.21
cc_394 ( N_noxref_3_M9_noxref_d N_noxref_10_c_968_n ) capacitor c=4.5543e-19 \
 //x=1.965 //y=5.02 //x2=4.205 //y2=5.21
cc_395 ( N_noxref_3_M11_noxref_g N_noxref_10_M11_noxref_s ) capacitor \
 c=0.0473218f //x=4.34 //y=6.025 //x2=3.985 //y2=5.025
cc_396 ( N_noxref_3_M12_noxref_g N_noxref_10_M12_noxref_d ) capacitor \
 c=0.0170604f //x=4.78 //y=6.025 //x2=4.855 //y2=5.025
cc_397 ( N_noxref_4_c_455_n N_noxref_5_c_600_n ) capacitor c=0.0114841f \
 //x=7.655 //y=2.59 //x2=9.365 //y2=2.59
cc_398 ( N_noxref_4_M16_noxref_g N_noxref_5_c_625_n ) capacitor c=0.0204115f \
 //x=8.11 //y=6.02 //x2=8.685 //y2=5.2
cc_399 ( N_noxref_4_c_469_n N_noxref_5_c_628_n ) capacitor c=0.0055959f \
 //x=7.77 //y=2.08 //x2=7.975 //y2=5.2
cc_400 ( N_noxref_4_M15_noxref_g N_noxref_5_c_628_n ) capacitor c=0.0177326f \
 //x=7.67 //y=6.02 //x2=7.975 //y2=5.2
cc_401 ( N_noxref_4_c_501_n N_noxref_5_c_628_n ) capacitor c=0.00605692f \
 //x=7.77 //y=4.7 //x2=7.975 //y2=5.2
cc_402 ( N_noxref_4_c_467_n N_noxref_5_c_603_n ) capacitor c=3.49822e-19 \
 //x=5.92 //y=2.59 //x2=9.25 //y2=2.59
cc_403 ( N_noxref_4_c_469_n N_noxref_5_c_603_n ) capacitor c=0.00369745f \
 //x=7.77 //y=2.08 //x2=9.25 //y2=2.59
cc_404 ( N_noxref_4_M16_noxref_g N_noxref_5_M15_noxref_d ) capacitor \
 c=0.0173476f //x=8.11 //y=6.02 //x2=7.745 //y2=5.02
cc_405 ( N_noxref_4_c_467_n N_C_c_906_n ) capacitor c=0.0102183f //x=5.92 \
 //y=2.59 //x2=5.18 //y2=4.54
cc_406 ( N_noxref_4_c_457_n N_C_c_893_n ) capacitor c=0.00316948f //x=6.035 \
 //y=2.59 //x2=5.18 //y2=2.08
cc_407 ( N_noxref_4_c_459_n N_C_c_893_n ) capacitor c=0.0162392f //x=5.395 \
 //y=1.655 //x2=5.18 //y2=2.08
cc_408 ( N_noxref_4_c_467_n N_C_c_893_n ) capacitor c=0.0822198f //x=5.92 \
 //y=2.59 //x2=5.18 //y2=2.08
cc_409 ( N_noxref_4_c_469_n N_C_c_893_n ) capacitor c=9.8819e-19 //x=7.77 \
 //y=2.08 //x2=5.18 //y2=2.08
cc_410 ( N_noxref_4_c_492_n N_C_M13_noxref_g ) capacitor c=0.0132788f \
 //x=5.525 //y=5.21 //x2=5.22 //y2=6.025
cc_411 ( N_noxref_4_c_490_n N_C_M14_noxref_g ) capacitor c=0.0217751f \
 //x=5.835 //y=5.21 //x2=5.66 //y2=6.025
cc_412 ( N_noxref_4_M13_noxref_d N_C_M14_noxref_g ) capacitor c=0.0136385f \
 //x=5.295 //y=5.025 //x2=5.66 //y2=6.025
cc_413 ( N_noxref_4_M3_noxref_d N_C_c_895_n ) capacitor c=0.00226395f //x=5.29 \
 //y=0.905 //x2=5.215 //y2=0.905
cc_414 ( N_noxref_4_M3_noxref_d N_C_c_918_n ) capacitor c=0.0035101f //x=5.29 \
 //y=0.905 //x2=5.215 //y2=1.255
cc_415 ( N_noxref_4_c_459_n N_C_c_921_n ) capacitor c=0.00218915f //x=5.395 \
 //y=1.655 //x2=5.215 //y2=1.56
cc_416 ( N_noxref_4_M2_noxref_d N_C_c_921_n ) capacitor c=0.00148728f //x=4.32 \
 //y=0.905 //x2=5.215 //y2=1.56
cc_417 ( N_noxref_4_M3_noxref_d N_C_c_921_n ) capacitor c=0.00546704f //x=5.29 \
 //y=0.905 //x2=5.215 //y2=1.56
cc_418 ( N_noxref_4_c_492_n N_C_c_945_n ) capacitor c=0.00417892f //x=5.525 \
 //y=5.21 //x2=5.585 //y2=4.795
cc_419 ( N_noxref_4_c_467_n N_C_c_945_n ) capacitor c=0.0144455f //x=5.92 \
 //y=2.59 //x2=5.585 //y2=4.795
cc_420 ( N_noxref_4_M3_noxref_d N_C_c_897_n ) capacitor c=0.00241102f //x=5.29 \
 //y=0.905 //x2=5.59 //y2=0.75
cc_421 ( N_noxref_4_c_463_n N_C_c_898_n ) capacitor c=0.00801563f //x=5.835 \
 //y=1.655 //x2=5.59 //y2=1.405
cc_422 ( N_noxref_4_M3_noxref_d N_C_c_898_n ) capacitor c=0.0158021f //x=5.29 \
 //y=0.905 //x2=5.59 //y2=1.405
cc_423 ( N_noxref_4_M3_noxref_d N_C_c_899_n ) capacitor c=0.00132831f //x=5.29 \
 //y=0.905 //x2=5.745 //y2=0.905
cc_424 ( N_noxref_4_M3_noxref_d N_C_c_925_n ) capacitor c=0.0035101f //x=5.29 \
 //y=0.905 //x2=5.745 //y2=1.255
cc_425 ( N_noxref_4_c_459_n N_C_c_926_n ) capacitor c=0.00633758f //x=5.395 \
 //y=1.655 //x2=5.18 //y2=2.08
cc_426 ( N_noxref_4_c_467_n N_C_c_926_n ) capacitor c=0.00877984f //x=5.92 \
 //y=2.59 //x2=5.18 //y2=2.08
cc_427 ( N_noxref_4_c_459_n N_C_c_928_n ) capacitor c=0.0189958f //x=5.395 \
 //y=1.655 //x2=5.18 //y2=1.915
cc_428 ( N_noxref_4_c_467_n N_C_c_928_n ) capacitor c=0.00306024f //x=5.92 \
 //y=2.59 //x2=5.18 //y2=1.915
cc_429 ( N_noxref_4_M3_noxref_d N_C_c_928_n ) capacitor c=3.4952e-19 //x=5.29 \
 //y=0.905 //x2=5.18 //y2=1.915
cc_430 ( N_noxref_4_c_467_n N_C_c_929_n ) capacitor c=0.00537091f //x=5.92 \
 //y=2.59 //x2=5.215 //y2=4.705
cc_431 ( N_noxref_4_c_492_n N_noxref_10_c_964_n ) capacitor c=0.0348754f \
 //x=5.525 //y=5.21 //x2=4.915 //y2=5.21
cc_432 ( N_noxref_4_c_490_n N_noxref_10_c_969_n ) capacitor c=0.00194034f \
 //x=5.835 //y=5.21 //x2=5.795 //y2=6.91
cc_433 ( N_noxref_4_M13_noxref_d N_noxref_10_c_969_n ) capacitor c=0.0118172f \
 //x=5.295 //y=5.025 //x2=5.795 //y2=6.91
cc_434 ( N_noxref_4_M13_noxref_d N_noxref_10_M11_noxref_s ) capacitor \
 c=0.00107541f //x=5.295 //y=5.025 //x2=3.985 //y2=5.025
cc_435 ( N_noxref_4_M13_noxref_d N_noxref_10_M12_noxref_d ) capacitor \
 c=0.0348754f //x=5.295 //y=5.025 //x2=4.855 //y2=5.025
cc_436 ( N_noxref_4_c_490_n N_noxref_10_M14_noxref_d ) capacitor c=0.0164221f \
 //x=5.835 //y=5.21 //x2=5.735 //y2=5.025
cc_437 ( N_noxref_4_M13_noxref_d N_noxref_10_M14_noxref_d ) capacitor \
 c=0.0458293f //x=5.295 //y=5.025 //x2=5.735 //y2=5.025
cc_438 ( N_noxref_4_c_469_n N_D_c_1016_n ) capacitor c=0.00400249f //x=7.77 \
 //y=2.08 //x2=8.51 //y2=4.535
cc_439 ( N_noxref_4_c_501_n N_D_c_1016_n ) capacitor c=0.00417994f //x=7.77 \
 //y=4.7 //x2=8.51 //y2=4.535
cc_440 ( N_noxref_4_c_455_n N_D_c_1007_n ) capacitor c=0.00316948f //x=7.655 \
 //y=2.59 //x2=8.51 //y2=2.08
cc_441 ( N_noxref_4_c_467_n N_D_c_1007_n ) capacitor c=9.8819e-19 //x=5.92 \
 //y=2.59 //x2=8.51 //y2=2.08
cc_442 ( N_noxref_4_c_469_n N_D_c_1007_n ) capacitor c=0.0872088f //x=7.77 \
 //y=2.08 //x2=8.51 //y2=2.08
cc_443 ( N_noxref_4_c_474_n N_D_c_1007_n ) capacitor c=0.00308814f //x=7.575 \
 //y=1.915 //x2=8.51 //y2=2.08
cc_444 ( N_noxref_4_M15_noxref_g N_D_M17_noxref_g ) capacitor c=0.0104611f \
 //x=7.67 //y=6.02 //x2=8.55 //y2=6.02
cc_445 ( N_noxref_4_M16_noxref_g N_D_M17_noxref_g ) capacitor c=0.106811f \
 //x=8.11 //y=6.02 //x2=8.55 //y2=6.02
cc_446 ( N_noxref_4_M16_noxref_g N_D_M18_noxref_g ) capacitor c=0.0100341f \
 //x=8.11 //y=6.02 //x2=8.99 //y2=6.02
cc_447 ( N_noxref_4_c_470_n N_D_c_1025_n ) capacitor c=4.86506e-19 //x=7.575 \
 //y=0.865 //x2=8.545 //y2=0.905
cc_448 ( N_noxref_4_c_472_n N_D_c_1025_n ) capacitor c=0.00152104f //x=7.575 \
 //y=1.21 //x2=8.545 //y2=0.905
cc_449 ( N_noxref_4_c_477_n N_D_c_1025_n ) capacitor c=0.0151475f //x=8.105 \
 //y=0.865 //x2=8.545 //y2=0.905
cc_450 ( N_noxref_4_c_473_n N_D_c_1028_n ) capacitor c=0.00109982f //x=7.575 \
 //y=1.52 //x2=8.545 //y2=1.25
cc_451 ( N_noxref_4_c_479_n N_D_c_1028_n ) capacitor c=0.0111064f //x=8.105 \
 //y=1.21 //x2=8.545 //y2=1.25
cc_452 ( N_noxref_4_c_473_n N_D_c_1030_n ) capacitor c=9.57794e-19 //x=7.575 \
 //y=1.52 //x2=8.545 //y2=1.56
cc_453 ( N_noxref_4_c_474_n N_D_c_1030_n ) capacitor c=0.00662747f //x=7.575 \
 //y=1.915 //x2=8.545 //y2=1.56
cc_454 ( N_noxref_4_c_479_n N_D_c_1030_n ) capacitor c=0.00862358f //x=8.105 \
 //y=1.21 //x2=8.545 //y2=1.56
cc_455 ( N_noxref_4_c_477_n N_D_c_1033_n ) capacitor c=0.00124821f //x=8.105 \
 //y=0.865 //x2=9.075 //y2=0.905
cc_456 ( N_noxref_4_c_479_n N_D_c_1034_n ) capacitor c=0.00200715f //x=8.105 \
 //y=1.21 //x2=9.075 //y2=1.25
cc_457 ( N_noxref_4_c_469_n N_D_c_1035_n ) capacitor c=0.00307062f //x=7.77 \
 //y=2.08 //x2=8.51 //y2=2.08
cc_458 ( N_noxref_4_c_474_n N_D_c_1035_n ) capacitor c=0.0179092f //x=7.575 \
 //y=1.915 //x2=8.51 //y2=2.08
cc_459 ( N_noxref_4_c_469_n N_D_c_1037_n ) capacitor c=0.00344981f //x=7.77 \
 //y=2.08 //x2=8.54 //y2=4.7
cc_460 ( N_noxref_4_c_501_n N_D_c_1037_n ) capacitor c=0.0293367f //x=7.77 \
 //y=4.7 //x2=8.54 //y2=4.7
cc_461 ( N_noxref_4_c_455_n N_noxref_12_c_1098_n ) capacitor c=0.00491973f \
 //x=7.655 //y=2.59 //x2=7.355 //y2=1.495
cc_462 ( N_noxref_4_c_463_n N_noxref_12_c_1098_n ) capacitor c=3.37788e-19 \
 //x=5.835 //y=1.655 //x2=7.355 //y2=1.495
cc_463 ( N_noxref_4_c_474_n N_noxref_12_c_1098_n ) capacitor c=0.0034165f \
 //x=7.575 //y=1.915 //x2=7.355 //y2=1.495
cc_464 ( N_noxref_4_c_455_n N_noxref_12_c_1073_n ) capacitor c=0.0108509f \
 //x=7.655 //y=2.59 //x2=8.24 //y2=1.58
cc_465 ( N_noxref_4_c_469_n N_noxref_12_c_1073_n ) capacitor c=0.0114076f \
 //x=7.77 //y=2.08 //x2=8.24 //y2=1.58
cc_466 ( N_noxref_4_c_473_n N_noxref_12_c_1073_n ) capacitor c=0.00700575f \
 //x=7.575 //y=1.52 //x2=8.24 //y2=1.58
cc_467 ( N_noxref_4_c_474_n N_noxref_12_c_1073_n ) capacitor c=0.018562f \
 //x=7.575 //y=1.915 //x2=8.24 //y2=1.58
cc_468 ( N_noxref_4_c_476_n N_noxref_12_c_1073_n ) capacitor c=0.00780629f \
 //x=7.95 //y=1.365 //x2=8.24 //y2=1.58
cc_469 ( N_noxref_4_c_479_n N_noxref_12_c_1073_n ) capacitor c=0.00339872f \
 //x=8.105 //y=1.21 //x2=8.24 //y2=1.58
cc_470 ( N_noxref_4_c_474_n N_noxref_12_c_1081_n ) capacitor c=6.71402e-19 \
 //x=7.575 //y=1.915 //x2=8.325 //y2=1.495
cc_471 ( N_noxref_4_c_470_n N_noxref_12_M4_noxref_s ) capacitor c=0.0326693f \
 //x=7.575 //y=0.865 //x2=7.22 //y2=0.365
cc_472 ( N_noxref_4_c_473_n N_noxref_12_M4_noxref_s ) capacitor c=3.48408e-19 \
 //x=7.575 //y=1.52 //x2=7.22 //y2=0.365
cc_473 ( N_noxref_4_c_477_n N_noxref_12_M4_noxref_s ) capacitor c=0.0120759f \
 //x=8.105 //y=0.865 //x2=7.22 //y2=0.365
cc_474 ( N_noxref_5_c_625_n N_D_c_1016_n ) capacitor c=0.0127867f //x=8.685 \
 //y=5.2 //x2=8.51 //y2=4.535
cc_475 ( N_noxref_5_c_603_n N_D_c_1016_n ) capacitor c=0.0101115f //x=9.25 \
 //y=2.59 //x2=8.51 //y2=4.535
cc_476 ( N_noxref_5_c_600_n N_D_c_1007_n ) capacitor c=0.00316373f //x=9.365 \
 //y=2.59 //x2=8.51 //y2=2.08
cc_477 ( N_noxref_5_c_603_n N_D_c_1007_n ) capacitor c=0.0820562f //x=9.25 \
 //y=2.59 //x2=8.51 //y2=2.08
cc_478 ( N_noxref_5_c_605_n N_D_c_1007_n ) capacitor c=0.00108914f //x=10.73 \
 //y=2.085 //x2=8.51 //y2=2.08
cc_479 ( N_noxref_5_c_625_n N_D_M17_noxref_g ) capacitor c=0.0166699f \
 //x=8.685 //y=5.2 //x2=8.55 //y2=6.02
cc_480 ( N_noxref_5_M17_noxref_d N_D_M17_noxref_g ) capacitor c=0.0173476f \
 //x=8.625 //y=5.02 //x2=8.55 //y2=6.02
cc_481 ( N_noxref_5_c_630_n N_D_M18_noxref_g ) capacitor c=0.0223814f \
 //x=9.165 //y=5.2 //x2=8.99 //y2=6.02
cc_482 ( N_noxref_5_M17_noxref_d N_D_M18_noxref_g ) capacitor c=0.0179769f \
 //x=8.625 //y=5.02 //x2=8.99 //y2=6.02
cc_483 ( N_noxref_5_M5_noxref_d N_D_c_1025_n ) capacitor c=0.00217566f \
 //x=8.62 //y=0.905 //x2=8.545 //y2=0.905
cc_484 ( N_noxref_5_M5_noxref_d N_D_c_1028_n ) capacitor c=0.0034598f //x=8.62 \
 //y=0.905 //x2=8.545 //y2=1.25
cc_485 ( N_noxref_5_M5_noxref_d N_D_c_1030_n ) capacitor c=0.0065582f //x=8.62 \
 //y=0.905 //x2=8.545 //y2=1.56
cc_486 ( N_noxref_5_c_603_n N_D_c_1051_n ) capacitor c=0.0142673f //x=9.25 \
 //y=2.59 //x2=8.915 //y2=4.79
cc_487 ( N_noxref_5_c_679_p N_D_c_1051_n ) capacitor c=0.00421574f //x=8.77 \
 //y=5.2 //x2=8.915 //y2=4.79
cc_488 ( N_noxref_5_M5_noxref_d N_D_c_1053_n ) capacitor c=0.00241102f \
 //x=8.62 //y=0.905 //x2=8.92 //y2=0.75
cc_489 ( N_noxref_5_c_601_n N_D_c_1054_n ) capacitor c=0.00359704f //x=9.165 \
 //y=1.655 //x2=8.92 //y2=1.405
cc_490 ( N_noxref_5_M5_noxref_d N_D_c_1054_n ) capacitor c=0.0138845f //x=8.62 \
 //y=0.905 //x2=8.92 //y2=1.405
cc_491 ( N_noxref_5_M5_noxref_d N_D_c_1033_n ) capacitor c=0.00132245f \
 //x=8.62 //y=0.905 //x2=9.075 //y2=0.905
cc_492 ( N_noxref_5_c_601_n N_D_c_1034_n ) capacitor c=0.00457401f //x=9.165 \
 //y=1.655 //x2=9.075 //y2=1.25
cc_493 ( N_noxref_5_M5_noxref_d N_D_c_1034_n ) capacitor c=0.00566463f \
 //x=8.62 //y=0.905 //x2=9.075 //y2=1.25
cc_494 ( N_noxref_5_c_603_n N_D_c_1035_n ) capacitor c=0.00877984f //x=9.25 \
 //y=2.59 //x2=8.51 //y2=2.08
cc_495 ( N_noxref_5_c_603_n N_D_c_1060_n ) capacitor c=0.00306024f //x=9.25 \
 //y=2.59 //x2=8.51 //y2=1.915
cc_496 ( N_noxref_5_M5_noxref_d N_D_c_1060_n ) capacitor c=0.00660593f \
 //x=8.62 //y=0.905 //x2=8.51 //y2=1.915
cc_497 ( N_noxref_5_c_625_n N_D_c_1037_n ) capacitor c=0.00399417f //x=8.685 \
 //y=5.2 //x2=8.54 //y2=4.7
cc_498 ( N_noxref_5_c_603_n N_D_c_1037_n ) capacitor c=0.00533692f //x=9.25 \
 //y=2.59 //x2=8.54 //y2=4.7
cc_499 ( N_noxref_5_c_691_p N_noxref_12_c_1098_n ) capacitor c=3.15806e-19 \
 //x=8.895 //y=1.655 //x2=7.355 //y2=1.495
cc_500 ( N_noxref_5_c_691_p N_noxref_12_c_1081_n ) capacitor c=0.0203424f \
 //x=8.895 //y=1.655 //x2=8.325 //y2=1.495
cc_501 ( N_noxref_5_c_601_n N_noxref_12_c_1082_n ) capacitor c=0.00468333f \
 //x=9.165 //y=1.655 //x2=9.21 //y2=0.53
cc_502 ( N_noxref_5_M5_noxref_d N_noxref_12_c_1082_n ) capacitor c=0.0118355f \
 //x=8.62 //y=0.905 //x2=9.21 //y2=0.53
cc_503 ( N_noxref_5_c_597_n N_noxref_12_M4_noxref_s ) capacitor c=3.03583e-19 \
 //x=10.615 //y=2.59 //x2=7.22 //y2=0.365
cc_504 ( N_noxref_5_c_600_n N_noxref_12_M4_noxref_s ) capacitor c=6.92363e-19 \
 //x=9.365 //y=2.59 //x2=7.22 //y2=0.365
cc_505 ( N_noxref_5_c_601_n N_noxref_12_M4_noxref_s ) capacitor c=0.0129465f \
 //x=9.165 //y=1.655 //x2=7.22 //y2=0.365
cc_506 ( N_noxref_5_M5_noxref_d N_noxref_12_M4_noxref_s ) capacitor \
 c=0.043966f //x=8.62 //y=0.905 //x2=7.22 //y2=0.365
cc_507 ( N_noxref_5_c_597_n Y ) capacitor c=0.00730959f //x=10.615 //y=2.59 \
 //x2=11.47 //y2=2.22
cc_508 ( N_noxref_5_c_603_n Y ) capacitor c=0.00108914f //x=9.25 //y=2.59 \
 //x2=11.47 //y2=2.22
cc_509 ( N_noxref_5_c_605_n Y ) capacitor c=0.0712221f //x=10.73 //y=2.085 \
 //x2=11.47 //y2=2.22
cc_510 ( N_noxref_5_c_617_n Y ) capacitor c=8.49451e-19 //x=10.73 //y=2.085 \
 //x2=11.47 //y2=2.22
cc_511 ( N_noxref_5_c_703_p N_Y_c_1129_n ) capacitor c=0.0023507f //x=11.215 \
 //y=1.41 //x2=11.385 //y2=2.08
cc_512 ( N_noxref_5_c_617_n N_Y_c_1152_n ) capacitor c=0.0167852f //x=10.73 \
 //y=2.085 //x2=11.185 //y2=2.08
cc_513 ( N_noxref_5_c_642_n N_Y_c_1139_n ) capacitor c=0.0107726f //x=11.25 \
 //y=4.79 //x2=11.385 //y2=4.58
cc_514 ( N_noxref_5_c_605_n N_Y_c_1141_n ) capacitor c=0.0250789f //x=10.73 \
 //y=2.085 //x2=11.19 //y2=4.58
cc_515 ( N_noxref_5_c_643_n N_Y_c_1141_n ) capacitor c=0.00962086f //x=10.96 \
 //y=4.79 //x2=11.19 //y2=4.58
cc_516 ( N_noxref_5_c_603_n N_Y_M6_noxref_d ) capacitor c=3.35192e-19 //x=9.25 \
 //y=2.59 //x2=10.915 //y2=0.91
cc_517 ( N_noxref_5_c_605_n N_Y_M6_noxref_d ) capacitor c=0.0175773f //x=10.73 \
 //y=2.085 //x2=10.915 //y2=0.91
cc_518 ( N_noxref_5_c_610_n N_Y_M6_noxref_d ) capacitor c=0.00218556f \
 //x=10.84 //y=0.91 //x2=10.915 //y2=0.91
cc_519 ( N_noxref_5_c_711_p N_Y_M6_noxref_d ) capacitor c=0.00347355f \
 //x=10.84 //y=1.255 //x2=10.915 //y2=0.91
cc_520 ( N_noxref_5_c_712_p N_Y_M6_noxref_d ) capacitor c=0.00742431f \
 //x=10.84 //y=1.565 //x2=10.915 //y2=0.91
cc_521 ( N_noxref_5_c_612_n N_Y_M6_noxref_d ) capacitor c=0.00957707f \
 //x=10.84 //y=1.92 //x2=10.915 //y2=0.91
cc_522 ( N_noxref_5_c_613_n N_Y_M6_noxref_d ) capacitor c=0.00220879f \
 //x=11.215 //y=0.755 //x2=10.915 //y2=0.91
cc_523 ( N_noxref_5_c_703_p N_Y_M6_noxref_d ) capacitor c=0.0138447f \
 //x=11.215 //y=1.41 //x2=10.915 //y2=0.91
cc_524 ( N_noxref_5_c_614_n N_Y_M6_noxref_d ) capacitor c=0.00218624f \
 //x=11.37 //y=0.91 //x2=10.915 //y2=0.91
cc_525 ( N_noxref_5_c_616_n N_Y_M6_noxref_d ) capacitor c=0.00601286f \
 //x=11.37 //y=1.255 //x2=10.915 //y2=0.91
cc_526 ( N_noxref_5_c_603_n N_Y_M19_noxref_d ) capacitor c=6.3502e-19 //x=9.25 \
 //y=2.59 //x2=10.96 //y2=5.02
cc_527 ( N_noxref_5_M19_noxref_g N_Y_M19_noxref_d ) capacitor c=0.0219309f \
 //x=10.885 //y=6.02 //x2=10.96 //y2=5.02
cc_528 ( N_noxref_5_M20_noxref_g N_Y_M19_noxref_d ) capacitor c=0.021902f \
 //x=11.325 //y=6.02 //x2=10.96 //y2=5.02
cc_529 ( N_noxref_5_c_642_n N_Y_M19_noxref_d ) capacitor c=0.0148755f \
 //x=11.25 //y=4.79 //x2=10.96 //y2=5.02
cc_530 ( N_noxref_5_c_643_n N_Y_M19_noxref_d ) capacitor c=0.00307344f \
 //x=10.96 //y=4.79 //x2=10.96 //y2=5.02
cc_531 ( N_A_c_723_n N_B_c_787_n ) capacitor c=0.00400249f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=4.535
cc_532 ( N_A_c_740_n N_B_c_787_n ) capacitor c=0.00417994f //x=1.11 //y=4.7 \
 //x2=1.85 //y2=4.535
cc_533 ( N_A_c_723_n N_B_c_778_n ) capacitor c=0.0887263f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_534 ( N_A_c_728_n N_B_c_778_n ) capacitor c=0.00308814f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_535 ( N_A_M7_noxref_g N_B_M9_noxref_g ) capacitor c=0.0104611f //x=1.01 \
 //y=6.02 //x2=1.89 //y2=6.02
cc_536 ( N_A_M8_noxref_g N_B_M9_noxref_g ) capacitor c=0.106811f //x=1.45 \
 //y=6.02 //x2=1.89 //y2=6.02
cc_537 ( N_A_M8_noxref_g N_B_M10_noxref_g ) capacitor c=0.0100341f //x=1.45 \
 //y=6.02 //x2=2.33 //y2=6.02
cc_538 ( N_A_c_724_n N_B_c_796_n ) capacitor c=4.86506e-19 //x=0.915 //y=0.865 \
 //x2=1.885 //y2=0.905
cc_539 ( N_A_c_726_n N_B_c_796_n ) capacitor c=0.00152104f //x=0.915 //y=1.21 \
 //x2=1.885 //y2=0.905
cc_540 ( N_A_c_731_n N_B_c_796_n ) capacitor c=0.0151475f //x=1.445 //y=0.865 \
 //x2=1.885 //y2=0.905
cc_541 ( N_A_c_727_n N_B_c_797_n ) capacitor c=0.00109982f //x=0.915 //y=1.52 \
 //x2=1.885 //y2=1.25
cc_542 ( N_A_c_733_n N_B_c_797_n ) capacitor c=0.0111064f //x=1.445 //y=1.21 \
 //x2=1.885 //y2=1.25
cc_543 ( N_A_c_727_n N_B_c_798_n ) capacitor c=9.57794e-19 //x=0.915 //y=1.52 \
 //x2=1.885 //y2=1.56
cc_544 ( N_A_c_728_n N_B_c_798_n ) capacitor c=0.00662747f //x=0.915 //y=1.915 \
 //x2=1.885 //y2=1.56
cc_545 ( N_A_c_733_n N_B_c_798_n ) capacitor c=0.00862358f //x=1.445 //y=1.21 \
 //x2=1.885 //y2=1.56
cc_546 ( N_A_c_731_n N_B_c_804_n ) capacitor c=0.00124821f //x=1.445 //y=0.865 \
 //x2=2.415 //y2=0.905
cc_547 ( N_A_c_733_n N_B_c_805_n ) capacitor c=0.00200715f //x=1.445 //y=1.21 \
 //x2=2.415 //y2=1.25
cc_548 ( N_A_c_723_n N_B_c_807_n ) capacitor c=0.00307062f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_549 ( N_A_c_728_n N_B_c_807_n ) capacitor c=0.0179092f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_550 ( N_A_c_723_n N_B_c_810_n ) capacitor c=0.00344981f //x=1.11 //y=2.08 \
 //x2=1.88 //y2=4.7
cc_551 ( N_A_c_740_n N_B_c_810_n ) capacitor c=0.0293367f //x=1.11 //y=4.7 \
 //x2=1.88 //y2=4.7
cc_552 ( N_A_c_728_n N_noxref_8_c_866_n ) capacitor c=0.0034165f //x=0.915 \
 //y=1.915 //x2=0.695 //y2=1.495
cc_553 ( N_A_c_723_n N_noxref_8_c_842_n ) capacitor c=0.0118986f //x=1.11 \
 //y=2.08 //x2=1.58 //y2=1.58
cc_554 ( N_A_c_727_n N_noxref_8_c_842_n ) capacitor c=0.00703567f //x=0.915 \
 //y=1.52 //x2=1.58 //y2=1.58
cc_555 ( N_A_c_728_n N_noxref_8_c_842_n ) capacitor c=0.0216532f //x=0.915 \
 //y=1.915 //x2=1.58 //y2=1.58
cc_556 ( N_A_c_730_n N_noxref_8_c_842_n ) capacitor c=0.00780629f //x=1.29 \
 //y=1.365 //x2=1.58 //y2=1.58
cc_557 ( N_A_c_733_n N_noxref_8_c_842_n ) capacitor c=0.00339872f //x=1.445 \
 //y=1.21 //x2=1.58 //y2=1.58
cc_558 ( N_A_c_728_n N_noxref_8_c_850_n ) capacitor c=6.71402e-19 //x=0.915 \
 //y=1.915 //x2=1.665 //y2=1.495
cc_559 ( N_A_c_724_n N_noxref_8_M0_noxref_s ) capacitor c=0.0326577f //x=0.915 \
 //y=0.865 //x2=0.56 //y2=0.365
cc_560 ( N_A_c_727_n N_noxref_8_M0_noxref_s ) capacitor c=3.48408e-19 \
 //x=0.915 //y=1.52 //x2=0.56 //y2=0.365
cc_561 ( N_A_c_731_n N_noxref_8_M0_noxref_s ) capacitor c=0.0120759f //x=1.445 \
 //y=0.865 //x2=0.56 //y2=0.365
cc_562 ( N_B_c_798_n N_noxref_8_c_850_n ) capacitor c=0.00623646f //x=1.885 \
 //y=1.56 //x2=1.665 //y2=1.495
cc_563 ( N_B_c_807_n N_noxref_8_c_850_n ) capacitor c=0.00172768f //x=1.85 \
 //y=2.08 //x2=1.665 //y2=1.495
cc_564 ( N_B_c_778_n N_noxref_8_c_851_n ) capacitor c=0.00161845f //x=1.85 \
 //y=2.08 //x2=2.55 //y2=0.53
cc_565 ( N_B_c_796_n N_noxref_8_c_851_n ) capacitor c=0.0186143f //x=1.885 \
 //y=0.905 //x2=2.55 //y2=0.53
cc_566 ( N_B_c_804_n N_noxref_8_c_851_n ) capacitor c=0.00656458f //x=2.415 \
 //y=0.905 //x2=2.55 //y2=0.53
cc_567 ( N_B_c_807_n N_noxref_8_c_851_n ) capacitor c=2.1838e-19 //x=1.85 \
 //y=2.08 //x2=2.55 //y2=0.53
cc_568 ( N_B_c_796_n N_noxref_8_M0_noxref_s ) capacitor c=0.00623646f \
 //x=1.885 //y=0.905 //x2=0.56 //y2=0.365
cc_569 ( N_B_c_804_n N_noxref_8_M0_noxref_s ) capacitor c=0.0143002f //x=2.415 \
 //y=0.905 //x2=0.56 //y2=0.365
cc_570 ( N_B_c_805_n N_noxref_8_M0_noxref_s ) capacitor c=0.00290153f \
 //x=2.415 //y=1.25 //x2=0.56 //y2=0.365
cc_571 ( N_C_M13_noxref_g N_noxref_10_c_964_n ) capacitor c=0.0170604f \
 //x=5.22 //y=6.025 //x2=4.915 //y2=5.21
cc_572 ( N_C_c_929_n N_noxref_10_c_964_n ) capacitor c=2.3112e-19 //x=5.215 \
 //y=4.705 //x2=4.915 //y2=5.21
cc_573 ( N_C_c_906_n N_noxref_10_c_969_n ) capacitor c=0.00109004f //x=5.18 \
 //y=4.54 //x2=5.795 //y2=6.91
cc_574 ( N_C_M13_noxref_g N_noxref_10_c_969_n ) capacitor c=0.0148484f \
 //x=5.22 //y=6.025 //x2=5.795 //y2=6.91
cc_575 ( N_C_M14_noxref_g N_noxref_10_c_969_n ) capacitor c=0.0163196f \
 //x=5.66 //y=6.025 //x2=5.795 //y2=6.91
cc_576 ( N_C_M14_noxref_g N_noxref_10_M14_noxref_d ) capacitor c=0.0351101f \
 //x=5.66 //y=6.025 //x2=5.735 //y2=5.025
cc_577 ( N_D_c_1030_n N_noxref_12_c_1081_n ) capacitor c=0.00623646f //x=8.545 \
 //y=1.56 //x2=8.325 //y2=1.495
cc_578 ( N_D_c_1035_n N_noxref_12_c_1081_n ) capacitor c=0.00172768f //x=8.51 \
 //y=2.08 //x2=8.325 //y2=1.495
cc_579 ( N_D_c_1007_n N_noxref_12_c_1082_n ) capacitor c=0.00161845f //x=8.51 \
 //y=2.08 //x2=9.21 //y2=0.53
cc_580 ( N_D_c_1025_n N_noxref_12_c_1082_n ) capacitor c=0.0186143f //x=8.545 \
 //y=0.905 //x2=9.21 //y2=0.53
cc_581 ( N_D_c_1033_n N_noxref_12_c_1082_n ) capacitor c=0.00656458f //x=9.075 \
 //y=0.905 //x2=9.21 //y2=0.53
cc_582 ( N_D_c_1035_n N_noxref_12_c_1082_n ) capacitor c=2.1838e-19 //x=8.51 \
 //y=2.08 //x2=9.21 //y2=0.53
cc_583 ( N_D_c_1025_n N_noxref_12_M4_noxref_s ) capacitor c=0.00623646f \
 //x=8.545 //y=0.905 //x2=7.22 //y2=0.365
cc_584 ( N_D_c_1033_n N_noxref_12_M4_noxref_s ) capacitor c=0.0143002f \
 //x=9.075 //y=0.905 //x2=7.22 //y2=0.365
cc_585 ( N_D_c_1034_n N_noxref_12_M4_noxref_s ) capacitor c=0.00290153f \
 //x=9.075 //y=1.25 //x2=7.22 //y2=0.365
