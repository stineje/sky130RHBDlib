VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AO3X1
  CLASS CORE ;
  FOREIGN AO3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.880 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 7.690 4.665 7.860 7.020 ;
        RECT 7.690 4.495 8.225 4.665 ;
        RECT 8.055 2.165 8.225 4.495 ;
        RECT 7.685 1.995 8.225 2.165 ;
        RECT 7.685 0.840 7.855 1.995 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.915 1.195 4.865 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.026450 ;
    PORT
      LAYER li1 ;
        RECT 5.130 4.710 5.300 4.870 ;
        RECT 5.095 4.540 5.300 4.710 ;
        RECT 5.095 1.915 5.265 4.540 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 9.315 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 9.050 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.475 5.555 4.645 7.230 ;
        RECT 6.490 4.110 6.830 7.230 ;
        RECT 7.250 5.185 7.420 7.230 ;
        RECT 8.130 5.185 8.300 7.230 ;
        RECT 8.710 4.110 9.050 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 9.050 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 9.050 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 3.940 0.615 4.110 1.745 ;
        RECT 4.910 0.615 5.080 1.390 ;
        RECT 5.880 0.615 6.050 1.390 ;
        RECT 3.940 0.445 6.050 0.615 ;
        RECT 3.940 0.170 4.110 0.445 ;
        RECT 4.425 0.170 4.595 0.445 ;
        RECT 4.910 0.170 5.080 0.445 ;
        RECT 5.395 0.170 5.565 0.445 ;
        RECT 5.880 0.170 6.050 0.445 ;
        RECT 6.490 0.170 6.830 2.720 ;
        RECT 7.205 0.620 7.375 1.750 ;
        RECT 8.175 0.620 8.345 1.750 ;
        RECT 7.205 0.450 8.345 0.620 ;
        RECT 7.205 0.170 7.375 0.450 ;
        RECT 7.690 0.170 7.860 0.450 ;
        RECT 8.175 0.170 8.345 0.450 ;
        RECT 8.710 0.170 9.050 2.720 ;
        RECT -0.170 -0.170 9.050 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 9.050 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 4.035 5.295 4.205 7.025 ;
        RECT 4.915 6.825 5.965 6.995 ;
        RECT 4.915 5.295 5.085 6.825 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 4.035 5.125 5.085 5.295 ;
        RECT 5.355 5.295 5.525 6.565 ;
        RECT 5.795 5.555 5.965 6.825 ;
        RECT 5.355 5.125 6.005 5.295 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.200 4.710 4.370 4.870 ;
        RECT 4.200 4.540 4.525 4.710 ;
        RECT 4.355 1.915 4.525 4.540 ;
        RECT 5.835 1.740 6.005 5.125 ;
        RECT 7.315 1.920 7.485 4.865 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 4.425 1.570 6.005 1.740 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 4.425 0.835 4.595 1.570 ;
        RECT 5.395 0.835 5.565 1.570 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 7.315 2.505 7.485 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 7.285 2.675 7.515 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 5.775 2.505 7.545 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 7.285 2.475 7.515 2.505 ;
  END
END AO3X1
END LIBRARY

