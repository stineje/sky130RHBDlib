* SPICE3 file created from TMRDFFQNX1.ext - technology: sky130A

.subckt TMRDFFQNX1 QN D CLK VDD GND
X0 GND dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 dffx1_pcell_0/m1_258_797# CLK dffx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X2 VDD dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/m1_258_797# VDD pshort w=2 l=0.15
X3 VDD CLK dffx1_pcell_0/m1_258_797# VDD pshort w=2 l=0.15
X4 GND dffx1_pcell_0/m1_833_723# dffx1_pcell_0/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X5 m1_3495_723# m1_3348_575# dffx1_pcell_0/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X6 VDD dffx1_pcell_0/m1_833_723# m1_3495_723# VDD pshort w=2 l=0.15
X7 VDD m1_3348_575# m1_3495_723# VDD pshort w=2 l=0.15
X8 GND m1_3495_723# dffx1_pcell_0/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X9 m1_3348_575# dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X10 VDD m1_3495_723# m1_3348_575# VDD pshort w=2 l=0.15
X11 VDD dffx1_pcell_0/m1_258_797# m1_3348_575# VDD pshort w=2 l=0.15
X12 GND dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X13 dffx1_pcell_0/m1_833_723# dffx1_pcell_0/m1_685_649# dffx1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X14 dffx1_pcell_0/nand3x1_pcell_0/li_393_182# CLK dffx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X15 VDD dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_833_723# VDD pshort w=2 l=0.15
X16 VDD CLK dffx1_pcell_0/m1_833_723# VDD pshort w=2 l=0.15
X17 VDD dffx1_pcell_0/m1_685_649# dffx1_pcell_0/m1_833_723# VDD pshort w=2 l=0.15
X18 GND dffx1_pcell_0/m1_833_723# dffx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X19 dffx1_pcell_0/m1_685_649# D dffx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X20 VDD dffx1_pcell_0/m1_833_723# dffx1_pcell_0/m1_685_649# VDD pshort w=2 l=0.15
X21 VDD D dffx1_pcell_0/m1_685_649# VDD pshort w=2 l=0.15
X22 GND dffx1_pcell_0/m1_685_649# dffx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X23 dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X24 VDD dffx1_pcell_0/m1_685_649# dffx1_pcell_0/m1_2165_649# VDD pshort w=2 l=0.15
X25 VDD dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_2165_649# VDD pshort w=2 l=0.15
X26 GND m1_11931_723# votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X27 GND m1_11931_723# votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X28 GND m1_3348_575# votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X29 votern3x1_pcell_0/a_805_1331# m1_11931_723# VDD VDD pshort w=2 l=0.15
X30 QN m1_3348_575# votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X31 votern3x1_pcell_0/a_805_1331# m1_7639_427# VDD VDD pshort w=2 l=0.15
X32 votern3x1_pcell_0/a_893_1059# m1_3348_575# votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X33 votern3x1_pcell_0/a_893_1059# m1_11931_723# votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X34 QN m1_3348_575# votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X35 QN m1_7639_427# votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X36 QN m1_7639_427# votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X37 QN m1_7639_427# votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X38 GND dffx1_pcell_1/m1_2165_649# dffx1_pcell_1/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X39 dffx1_pcell_1/m1_258_797# CLK dffx1_pcell_1/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X40 VDD dffx1_pcell_1/m1_2165_649# dffx1_pcell_1/m1_258_797# VDD pshort w=2 l=0.15
X41 VDD CLK dffx1_pcell_1/m1_258_797# VDD pshort w=2 l=0.15
X42 GND dffx1_pcell_1/m1_833_723# dffx1_pcell_1/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X43 m1_7741_723# m1_7639_427# dffx1_pcell_1/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X44 VDD dffx1_pcell_1/m1_833_723# m1_7741_723# VDD pshort w=2 l=0.15
X45 VDD m1_7639_427# m1_7741_723# VDD pshort w=2 l=0.15
X46 GND m1_7741_723# dffx1_pcell_1/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X47 m1_7639_427# dffx1_pcell_1/m1_258_797# dffx1_pcell_1/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X48 VDD m1_7741_723# m1_7639_427# VDD pshort w=2 l=0.15
X49 VDD dffx1_pcell_1/m1_258_797# m1_7639_427# VDD pshort w=2 l=0.15
X50 GND dffx1_pcell_1/m1_258_797# dffx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X51 dffx1_pcell_1/m1_833_723# dffx1_pcell_1/m1_685_649# dffx1_pcell_1/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X52 dffx1_pcell_1/nand3x1_pcell_0/li_393_182# CLK dffx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X53 VDD dffx1_pcell_1/m1_258_797# dffx1_pcell_1/m1_833_723# VDD pshort w=2 l=0.15
X54 VDD CLK dffx1_pcell_1/m1_833_723# VDD pshort w=2 l=0.15
X55 VDD dffx1_pcell_1/m1_685_649# dffx1_pcell_1/m1_833_723# VDD pshort w=2 l=0.15
X56 GND dffx1_pcell_1/m1_833_723# dffx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X57 dffx1_pcell_1/m1_685_649# D dffx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X58 VDD dffx1_pcell_1/m1_833_723# dffx1_pcell_1/m1_685_649# VDD pshort w=2 l=0.15
X59 VDD D dffx1_pcell_1/m1_685_649# VDD pshort w=2 l=0.15
X60 GND dffx1_pcell_1/m1_685_649# dffx1_pcell_1/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X61 dffx1_pcell_1/m1_2165_649# dffx1_pcell_1/m1_258_797# dffx1_pcell_1/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X62 VDD dffx1_pcell_1/m1_685_649# dffx1_pcell_1/m1_2165_649# VDD pshort w=2 l=0.15
X63 VDD dffx1_pcell_1/m1_258_797# dffx1_pcell_1/m1_2165_649# VDD pshort w=2 l=0.15
X64 GND dffx1_pcell_2/m1_2165_649# dffx1_pcell_2/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X65 dffx1_pcell_2/m1_258_797# CLK dffx1_pcell_2/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X66 VDD dffx1_pcell_2/m1_2165_649# dffx1_pcell_2/m1_258_797# VDD pshort w=2 l=0.15
X67 VDD CLK dffx1_pcell_2/m1_258_797# VDD pshort w=2 l=0.15
X68 GND dffx1_pcell_2/m1_833_723# dffx1_pcell_2/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X69 m1_12079_871# m1_11931_723# dffx1_pcell_2/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X70 VDD dffx1_pcell_2/m1_833_723# m1_12079_871# VDD pshort w=2 l=0.15
X71 VDD m1_11931_723# m1_12079_871# VDD pshort w=2 l=0.15
X72 GND m1_12079_871# dffx1_pcell_2/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X73 m1_11931_723# dffx1_pcell_2/m1_258_797# dffx1_pcell_2/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X74 VDD m1_12079_871# m1_11931_723# VDD pshort w=2 l=0.15
X75 VDD dffx1_pcell_2/m1_258_797# m1_11931_723# VDD pshort w=2 l=0.15
X76 GND dffx1_pcell_2/m1_258_797# dffx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X77 dffx1_pcell_2/m1_833_723# dffx1_pcell_2/m1_685_649# dffx1_pcell_2/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X78 dffx1_pcell_2/nand3x1_pcell_0/li_393_182# CLK dffx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X79 VDD dffx1_pcell_2/m1_258_797# dffx1_pcell_2/m1_833_723# VDD pshort w=2 l=0.15
X80 VDD CLK dffx1_pcell_2/m1_833_723# VDD pshort w=2 l=0.15
X81 VDD dffx1_pcell_2/m1_685_649# dffx1_pcell_2/m1_833_723# VDD pshort w=2 l=0.15
X82 GND dffx1_pcell_2/m1_833_723# dffx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X83 dffx1_pcell_2/m1_685_649# D dffx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X84 VDD dffx1_pcell_2/m1_833_723# dffx1_pcell_2/m1_685_649# VDD pshort w=2 l=0.15
X85 VDD D dffx1_pcell_2/m1_685_649# VDD pshort w=2 l=0.15
X86 GND dffx1_pcell_2/m1_685_649# dffx1_pcell_2/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X87 dffx1_pcell_2/m1_2165_649# dffx1_pcell_2/m1_258_797# dffx1_pcell_2/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X88 VDD dffx1_pcell_2/m1_685_649# dffx1_pcell_2/m1_2165_649# VDD pshort w=2 l=0.15
X89 VDD dffx1_pcell_2/m1_258_797# dffx1_pcell_2/m1_2165_649# VDD pshort w=2 l=0.15
C0 VDD dffx1_pcell_2/m1_258_797# 2.40fF
C1 VDD dffx1_pcell_1/m1_258_797# 2.41fF
C2 VDD dffx1_pcell_0/m1_258_797# 2.43fF
C3 VDD CLK 5.29fF
.ends
