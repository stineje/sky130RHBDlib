* SPICE3 file created from INVX1.ext - technology: sky130A

.subckt INVX1 Y A VDD VSS
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8p pd=4.58u as=1.1p ps=9.1u w=2u l=0.15u M=2
X1 Y A VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=1.1408p ps=8.1u w=3u l=0.15u
.ends
