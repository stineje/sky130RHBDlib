* SPICE3 file created from AND2X1.ext - technology: sky130A

.subckt AND2X1 Y A B VDD GND
X0 Y and2x1_pcell_0/m1_547_649# GND GND nshort w=3 l=0.15
X1 VDD and2x1_pcell_0/m1_547_649# Y VDD pshort w=2 l=0.15
X2 GND A and2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X3 and2x1_pcell_0/m1_547_649# B and2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X4 VDD A and2x1_pcell_0/m1_547_649# VDD pshort w=2 l=0.15
X5 VDD B and2x1_pcell_0/m1_547_649# VDD pshort w=2 l=0.15
C0 VDD GND 3.25fF
.ends
