magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 14 21 396 157
rect 29 -17 63 21
<< scnmos >>
rect 93 47 123 131
rect 165 47 195 131
rect 287 47 317 131
<< scpmoshvt >>
rect 93 413 123 497
rect 181 413 211 497
rect 335 369 365 497
<< ndiff >>
rect 40 106 93 131
rect 40 72 48 106
rect 82 72 93 106
rect 40 47 93 72
rect 123 47 165 131
rect 195 89 287 131
rect 195 55 219 89
rect 253 55 287 89
rect 195 47 287 55
rect 317 93 370 131
rect 317 59 328 93
rect 362 59 370 93
rect 317 47 370 59
<< pdiff >>
rect 40 485 93 497
rect 40 451 48 485
rect 82 451 93 485
rect 40 413 93 451
rect 123 477 181 497
rect 123 443 136 477
rect 170 443 181 477
rect 123 413 181 443
rect 211 485 335 497
rect 211 451 222 485
rect 256 451 290 485
rect 324 451 335 485
rect 211 417 335 451
rect 211 413 288 417
rect 237 383 288 413
rect 322 383 335 417
rect 237 369 335 383
rect 365 485 418 497
rect 365 451 376 485
rect 410 451 418 485
rect 365 417 418 451
rect 365 383 376 417
rect 410 383 418 417
rect 365 369 418 383
<< ndiffc >>
rect 48 72 82 106
rect 219 55 253 89
rect 328 59 362 93
<< pdiffc >>
rect 48 451 82 485
rect 136 443 170 477
rect 222 451 256 485
rect 290 451 324 485
rect 288 383 322 417
rect 376 451 410 485
rect 376 383 410 417
<< poly >>
rect 93 497 123 523
rect 181 497 211 523
rect 335 497 365 523
rect 93 376 123 413
rect 36 360 123 376
rect 36 326 52 360
rect 86 326 123 360
rect 181 342 211 413
rect 36 292 123 326
rect 36 258 52 292
rect 86 258 123 292
rect 36 242 123 258
rect 93 131 123 242
rect 165 321 254 342
rect 165 287 204 321
rect 238 287 254 321
rect 335 287 365 369
rect 165 253 254 287
rect 165 219 204 253
rect 238 219 254 253
rect 165 209 254 219
rect 296 271 365 287
rect 296 237 306 271
rect 340 237 365 271
rect 165 131 195 209
rect 296 203 365 237
rect 296 183 306 203
rect 287 169 306 183
rect 340 169 365 203
rect 287 153 365 169
rect 287 131 317 153
rect 93 21 123 47
rect 165 21 195 47
rect 287 21 317 47
<< polycont >>
rect 52 326 86 360
rect 52 258 86 292
rect 204 287 238 321
rect 204 219 238 253
rect 306 237 340 271
rect 306 169 340 203
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 32 485 86 527
rect 32 451 48 485
rect 82 451 86 485
rect 32 435 86 451
rect 120 477 173 493
rect 120 443 136 477
rect 170 443 173 477
rect 120 427 173 443
rect 222 485 324 527
rect 256 451 290 485
rect 17 360 86 391
rect 17 326 52 360
rect 17 292 86 326
rect 17 258 52 292
rect 17 237 86 258
rect 120 190 154 427
rect 222 417 324 451
rect 222 383 288 417
rect 322 383 324 417
rect 222 367 324 383
rect 358 485 443 493
rect 358 451 376 485
rect 410 451 443 485
rect 358 417 443 451
rect 358 383 376 417
rect 410 383 443 417
rect 358 367 443 383
rect 188 321 254 323
rect 188 287 204 321
rect 238 287 254 321
rect 188 253 254 287
rect 188 219 204 253
rect 238 219 254 253
rect 188 216 254 219
rect 290 271 356 287
rect 290 237 306 271
rect 340 237 356 271
rect 37 182 154 190
rect 290 203 356 237
rect 290 182 306 203
rect 37 169 306 182
rect 340 169 356 203
rect 37 139 356 169
rect 37 106 98 139
rect 37 72 48 106
rect 82 72 98 106
rect 390 105 443 367
rect 37 56 98 72
rect 190 89 278 105
rect 190 55 219 89
rect 253 55 278 89
rect 190 17 278 55
rect 312 93 443 105
rect 312 59 328 93
rect 362 59 443 93
rect 312 51 443 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 397 425 431 459 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 213 289 247 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 29 357 63 391 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
rlabel comment s 0 0 0 0 4 and2_0
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 3818138
string GDS_START 3813716
string path 0.000 0.000 11.500 0.000 
<< end >>
