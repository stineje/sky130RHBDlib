magic
tech sky130A
timestamp 1648060378
<< poly >>
rect -16 8 17 13
rect -16 -9 -8 8
rect 9 -9 17 8
rect -16 -14 17 -9
<< polycont >>
rect -8 -9 9 8
<< locali >>
rect -16 -9 -8 8
rect 9 -9 17 8
<< end >>
