* SPICE3 file created from TMRDFFQX1.ext - technology: sky130A

.subckt TMRDFFQX1 D CLK Q VDD GND
M1000 GND a_7469_1050.t5 a_8030_101.t0 nshort w=-1.605u l=1.765u
+  ad=4.9019p pd=41.07u as=0p ps=0u
M1001 a_599_989.t1 D.t0 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t43 a_10429_1050.t5 a_8731_187.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_13268_209.t5 a_7595_411.t5 a_13757_1051.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_10429_1050.t0 a_8731_187.t5 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD.t53 a_13268_209.t7 Q.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_7469_1050.t1 a_7595_411.t7 VDD.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t51 a_9183_989.t5 a_8861_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 GND a_1845_1050.t5 a_2406_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_4569_1050.t1 CLK.t0 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VDD.t2 a_4439_187.t5 a_6137_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1845_1050.t4 a_599_989.t5 VDD.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VDD.t29 a_8861_1050.t7 a_9183_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_8861_1050.t6 CLK.t1 VDD.t50 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 GND a_8861_1050.t8 a_9658_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_13093_1051.t1 a_11887_411.t5 VDD.t42 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VDD.t38 a_147_187.t6 a_1845_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_6137_1050.t1 a_4891_989.t5 VDD.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VDD.t32 a_4569_1050.t7 a_4891_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_13093_1051.t3 a_11887_411.t6 a_13757_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VDD.t21 a_4439_187.t6 a_7595_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t56 a_147_187.t7 a_277_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t15 a_6137_1050.t5 a_4439_187.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VDD.t69 a_8731_187.t8 a_8861_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 GND a_147_187.t8 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_3177_1050.t4 a_277_1050.t7 VDD.t77 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VDD.t66 a_1845_1050.t6 a_147_187.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_11887_411.t4 a_11761_1050.t5 VDD.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 VDD.t7 D.t2 a_9183_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 GND a_8861_1050.t9 a_11656_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1030 VDD.t4 D.t3 a_4891_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 GND a_10429_1050.t6 a_10990_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1032 GND a_4439_187.t8 a_4383_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1033 VDD.t39 a_7469_1050.t6 a_7595_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VDD.t60 CLK.t2 a_277_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_13757_1051.t4 a_7595_411.t8 a_13268_209.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_3177_1050.t1 a_3303_411.t7 VDD.t81 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VDD.t47 CLK.t5 a_147_187.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_11887_411.t2 a_8731_187.t10 VDD.t68 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 GND a_599_989.t8 a_1740_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1040 VDD.t41 a_11887_411.t7 a_11761_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 GND a_4569_1050.t9 a_5366_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1042 Q a_13268_209.t9 GND.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1043 VDD.t17 CLK.t6 a_4439_187.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 GND a_11887_411.t8 a_13654_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_9183_989.t0 D.t4 VDD.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_3303_411.t4 a_3177_1050.t5 VDD.t79 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 GND a_11887_411.t10 a_12988_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1048 VDD.t49 a_599_989.t7 a_277_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 VDD.t11 a_277_1050.t8 a_599_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_8731_187.t3 a_10429_1050.t7 VDD.t57 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_4569_1050.t6 a_4891_989.t7 VDD.t74 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 a_13757_1051.t2 a_3303_411.t8 a_13268_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 VDD.t61 a_9183_989.t6 a_10429_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 VDD.t37 a_147_187.t9 a_3303_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_7595_411.t4 a_7469_1050.t7 VDD.t54 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 Q.t0 a_13268_209.t8 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 VDD.t36 a_4569_1050.t8 a_7469_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_4439_187.t1 CLK.t7 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 a_1845_1050.t0 a_147_187.t10 VDD.t55 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 a_8861_1050.t1 a_9183_989.t7 VDD.t65 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 VDD.t33 a_4439_187.t10 a_4569_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_6137_1050.t2 a_4439_187.t11 VDD.t78 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 GND a_3177_1050.t6 a_3738_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1064 GND a_4569_1050.t10 a_7364_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1065 a_9183_989.t4 a_8861_1050.t10 VDD.t59 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 GND a_9183_989.t8 a_10324_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_13093_1051.t5 a_3303_411.t9 a_13757_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_11761_1050.t1 a_11887_411.t9 VDD.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_3303_411.t3 a_147_187.t11 VDD.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 VDD.t83 a_7595_411.t10 a_13093_1051.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 VDD.t9 D.t5 a_599_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_8731_187.t1 CLK.t9 VDD.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 a_13757_1051.t7 a_11887_411.t11 a_13093_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 VDD.t67 a_8731_187.t11 a_10429_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 a_277_1050.t2 a_147_187.t12 VDD.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 a_4439_187.t0 a_6137_1050.t6 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 VDD.t70 a_7595_411.t11 a_7469_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 GND a_277_1050.t9 a_1074_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1079 VDD.t35 CLK.t12 a_4569_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 VDD.t76 a_599_989.t9 a_1845_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 a_11761_1050.t4 a_8861_1050.t11 VDD.t48 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 VDD.t23 a_11887_411.t12 a_13093_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_4891_989.t1 D.t7 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 GND a_11761_1050.t7 a_12322_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_13757_1051.t1 a_3303_411.t10 a_13093_1051.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_277_1050.t0 CLK.t13 VDD.t64 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 VDD.t10 a_4891_989.t8 a_4569_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 VDD.t62 a_277_1050.t10 a_3177_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_147_187.t3 CLK.t15 VDD.t63 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 VDD.t19 a_11761_1050.t6 a_11887_411.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 GND a_6137_1050.t7 a_6698_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1092 GND a_277_1050.t12 a_3072_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_4891_989.t3 a_4569_1050.t11 VDD.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_7595_411.t3 a_4439_187.t12 VDD.t52 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 GND a_4891_989.t10 a_6032_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1096 a_277_1050.t4 a_599_989.t10 VDD.t46 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_599_989.t4 a_277_1050.t11 VDD.t44 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 GND a_3303_411.t5 a_14320_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1099 a_13268_209.t0 a_3303_411.t11 a_13757_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_8861_1050.t4 a_8731_187.t12 VDD.t82 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 VDD.t30 CLK.t16 a_8731_187.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_10429_1050.t1 a_9183_989.t10 VDD.t26 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_7469_1050.t3 a_4569_1050.t12 VDD.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_147_187.t1 a_1845_1050.t7 VDD.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 VDD.t80 a_3303_411.t12 a_3177_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VDD.t72 a_8731_187.t13 a_11887_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 VDD.t28 CLK.t17 a_8861_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 a_4569_1050.t4 a_4439_187.t13 VDD.t40 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 VDD.t16 a_4891_989.t9 a_6137_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 VDD.t58 a_8861_1050.t12 a_11761_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 GND a_8731_187.t7 a_8675_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1112 VDD.t13 a_3177_1050.t7 a_3303_411.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 a_13093_1051.t6 a_7595_411.t13 VDD.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD CLK 1.74fF
C1 VDD D 0.22fF
C2 VDD Q 0.76fF
C3 CLK D 0.45fF
R0 D.n5 D.t5 472.359
R1 D.n2 D.t3 472.359
R2 D.n0 D.t2 472.359
R3 D.n5 D.t0 384.527
R4 D.n2 D.t7 384.527
R5 D.n0 D.t4 384.527
R6 D.n6 D.n5 216.272
R7 D.n3 D.n2 216.272
R8 D.n1 D.n0 216.272
R9 D.n6 D.t1 141.114
R10 D.n3 D.t8 141.114
R11 D.n1 D.t6 141.114
R12 D.n4 D.n1 91.734
R13 D.n4 D.n3 76
R14 D.n7 D.n6 76
R15 D.n7 D.n4 15.734
R16 D.n7 D 0.046
R17 VDD.n799 VDD.n797 144.705
R18 VDD.n860 VDD.n858 144.705
R19 VDD.n921 VDD.n919 144.705
R20 VDD.n982 VDD.n980 144.705
R21 VDD.n1043 VDD.n1041 144.705
R22 VDD.n1104 VDD.n1102 144.705
R23 VDD.n1185 VDD.n1183 144.705
R24 VDD.n1246 VDD.n1244 144.705
R25 VDD.n1307 VDD.n1305 144.705
R26 VDD.n684 VDD.n682 144.705
R27 VDD.n1368 VDD.n1366 144.705
R28 VDD.n623 VDD.n621 144.705
R29 VDD.n542 VDD.n540 144.705
R30 VDD.n481 VDD.n479 144.705
R31 VDD.n420 VDD.n418 144.705
R32 VDD.n359 VDD.n357 144.705
R33 VDD.n298 VDD.n296 144.705
R34 VDD.n237 VDD.n235 144.705
R35 VDD.n176 VDD.n174 144.705
R36 VDD.n122 VDD.n120 144.705
R37 VDD.n68 VDD.n66 144.705
R38 VDD.n26 VDD.n25 77.792
R39 VDD.n35 VDD.n34 77.792
R40 VDD.n29 VDD.n23 76.145
R41 VDD.n29 VDD.n28 76
R42 VDD.n33 VDD.n32 76
R43 VDD.n39 VDD.n38 76
R44 VDD.n43 VDD.n42 76
R45 VDD.n70 VDD.n69 76
R46 VDD.n74 VDD.n73 76
R47 VDD.n78 VDD.n77 76
R48 VDD.n82 VDD.n81 76
R49 VDD.n86 VDD.n85 76
R50 VDD.n90 VDD.n89 76
R51 VDD.n94 VDD.n93 76
R52 VDD.n98 VDD.n97 76
R53 VDD.n124 VDD.n123 76
R54 VDD.n128 VDD.n127 76
R55 VDD.n132 VDD.n131 76
R56 VDD.n136 VDD.n135 76
R57 VDD.n140 VDD.n139 76
R58 VDD.n144 VDD.n143 76
R59 VDD.n148 VDD.n147 76
R60 VDD.n152 VDD.n151 76
R61 VDD.n178 VDD.n177 76
R62 VDD.n183 VDD.n182 76
R63 VDD.n188 VDD.n187 76
R64 VDD.n194 VDD.n193 76
R65 VDD.n199 VDD.n198 76
R66 VDD.n204 VDD.n203 76
R67 VDD.n209 VDD.n208 76
R68 VDD.n213 VDD.n212 76
R69 VDD.n239 VDD.n238 76
R70 VDD.n244 VDD.n243 76
R71 VDD.n249 VDD.n248 76
R72 VDD.n255 VDD.n254 76
R73 VDD.n260 VDD.n259 76
R74 VDD.n265 VDD.n264 76
R75 VDD.n270 VDD.n269 76
R76 VDD.n274 VDD.n273 76
R77 VDD.n300 VDD.n299 76
R78 VDD.n305 VDD.n304 76
R79 VDD.n310 VDD.n309 76
R80 VDD.n316 VDD.n315 76
R81 VDD.n321 VDD.n320 76
R82 VDD.n326 VDD.n325 76
R83 VDD.n331 VDD.n330 76
R84 VDD.n335 VDD.n334 76
R85 VDD.n361 VDD.n360 76
R86 VDD.n366 VDD.n365 76
R87 VDD.n371 VDD.n370 76
R88 VDD.n377 VDD.n376 76
R89 VDD.n382 VDD.n381 76
R90 VDD.n387 VDD.n386 76
R91 VDD.n392 VDD.n391 76
R92 VDD.n396 VDD.n395 76
R93 VDD.n422 VDD.n421 76
R94 VDD.n427 VDD.n426 76
R95 VDD.n432 VDD.n431 76
R96 VDD.n438 VDD.n437 76
R97 VDD.n443 VDD.n442 76
R98 VDD.n448 VDD.n447 76
R99 VDD.n453 VDD.n452 76
R100 VDD.n457 VDD.n456 76
R101 VDD.n483 VDD.n482 76
R102 VDD.n488 VDD.n487 76
R103 VDD.n493 VDD.n492 76
R104 VDD.n499 VDD.n498 76
R105 VDD.n504 VDD.n503 76
R106 VDD.n509 VDD.n508 76
R107 VDD.n514 VDD.n513 76
R108 VDD.n518 VDD.n517 76
R109 VDD.n544 VDD.n543 76
R110 VDD.n548 VDD.n547 76
R111 VDD.n552 VDD.n551 76
R112 VDD.n557 VDD.n556 76
R113 VDD.n564 VDD.n563 76
R114 VDD.n569 VDD.n568 76
R115 VDD.n574 VDD.n573 76
R116 VDD.n581 VDD.n580 76
R117 VDD.n586 VDD.n585 76
R118 VDD.n591 VDD.n590 76
R119 VDD.n595 VDD.n594 76
R120 VDD.n599 VDD.n598 76
R121 VDD.n625 VDD.n624 76
R122 VDD.n630 VDD.n629 76
R123 VDD.n635 VDD.n634 76
R124 VDD.n641 VDD.n640 76
R125 VDD.n646 VDD.n645 76
R126 VDD.n651 VDD.n650 76
R127 VDD.n656 VDD.n655 76
R128 VDD.n660 VDD.n659 76
R129 VDD.n686 VDD.n685 76
R130 VDD.n691 VDD.n690 76
R131 VDD.n696 VDD.n695 76
R132 VDD.n1391 VDD.n1390 76
R133 VDD.n1385 VDD.n1384 76
R134 VDD.n1380 VDD.n1379 76
R135 VDD.n1375 VDD.n1374 76
R136 VDD.n1370 VDD.n1369 76
R137 VDD.n1344 VDD.n1343 76
R138 VDD.n1340 VDD.n1339 76
R139 VDD.n1335 VDD.n1334 76
R140 VDD.n1330 VDD.n1329 76
R141 VDD.n1324 VDD.n1323 76
R142 VDD.n1319 VDD.n1318 76
R143 VDD.n1314 VDD.n1313 76
R144 VDD.n1309 VDD.n1308 76
R145 VDD.n1283 VDD.n1282 76
R146 VDD.n1279 VDD.n1278 76
R147 VDD.n1274 VDD.n1273 76
R148 VDD.n1269 VDD.n1268 76
R149 VDD.n1263 VDD.n1262 76
R150 VDD.n1258 VDD.n1257 76
R151 VDD.n1253 VDD.n1252 76
R152 VDD.n1248 VDD.n1247 76
R153 VDD.n1222 VDD.n1221 76
R154 VDD.n1218 VDD.n1217 76
R155 VDD.n1213 VDD.n1212 76
R156 VDD.n1208 VDD.n1207 76
R157 VDD.n1202 VDD.n1201 76
R158 VDD.n1197 VDD.n1196 76
R159 VDD.n1192 VDD.n1191 76
R160 VDD.n1187 VDD.n1186 76
R161 VDD.n1161 VDD.n1160 76
R162 VDD.n1157 VDD.n1156 76
R163 VDD.n1153 VDD.n1152 76
R164 VDD.n1149 VDD.n1148 76
R165 VDD.n1144 VDD.n1143 76
R166 VDD.n1137 VDD.n1136 76
R167 VDD.n1132 VDD.n1131 76
R168 VDD.n1127 VDD.n1126 76
R169 VDD.n1120 VDD.n1119 76
R170 VDD.n1115 VDD.n1114 76
R171 VDD.n1110 VDD.n1109 76
R172 VDD.n1106 VDD.n1105 76
R173 VDD.n1080 VDD.n1079 76
R174 VDD.n1076 VDD.n1075 76
R175 VDD.n1071 VDD.n1070 76
R176 VDD.n1066 VDD.n1065 76
R177 VDD.n1060 VDD.n1059 76
R178 VDD.n1055 VDD.n1054 76
R179 VDD.n1050 VDD.n1049 76
R180 VDD.n1045 VDD.n1044 76
R181 VDD.n1019 VDD.n1018 76
R182 VDD.n1015 VDD.n1014 76
R183 VDD.n1010 VDD.n1009 76
R184 VDD.n1005 VDD.n1004 76
R185 VDD.n999 VDD.n998 76
R186 VDD.n994 VDD.n993 76
R187 VDD.n989 VDD.n988 76
R188 VDD.n984 VDD.n983 76
R189 VDD.n958 VDD.n957 76
R190 VDD.n954 VDD.n953 76
R191 VDD.n949 VDD.n948 76
R192 VDD.n944 VDD.n943 76
R193 VDD.n938 VDD.n937 76
R194 VDD.n933 VDD.n932 76
R195 VDD.n928 VDD.n927 76
R196 VDD.n923 VDD.n922 76
R197 VDD.n897 VDD.n896 76
R198 VDD.n893 VDD.n892 76
R199 VDD.n888 VDD.n887 76
R200 VDD.n883 VDD.n882 76
R201 VDD.n877 VDD.n876 76
R202 VDD.n872 VDD.n871 76
R203 VDD.n867 VDD.n866 76
R204 VDD.n862 VDD.n861 76
R205 VDD.n836 VDD.n835 76
R206 VDD.n832 VDD.n831 76
R207 VDD.n827 VDD.n826 76
R208 VDD.n822 VDD.n821 76
R209 VDD.n816 VDD.n815 76
R210 VDD.n811 VDD.n810 76
R211 VDD.n806 VDD.n805 76
R212 VDD.n801 VDD.n800 76
R213 VDD.n774 VDD.n773 76
R214 VDD.n770 VDD.n769 76
R215 VDD.n766 VDD.n765 76
R216 VDD.n762 VDD.n761 76
R217 VDD.n757 VDD.n756 76
R218 VDD.n750 VDD.n749 76
R219 VDD.n745 VDD.n744 76
R220 VDD.n740 VDD.n739 76
R221 VDD.n733 VDD.n732 76
R222 VDD.n728 VDD.n727 76
R223 VDD.n723 VDD.n722 76
R224 VDD.n719 VDD.n718 76
R225 VDD.n554 VDD.n553 64.064
R226 VDD.n1146 VDD.n1145 64.064
R227 VDD.n759 VDD.n758 64.064
R228 VDD.n583 VDD.n582 59.488
R229 VDD.n1117 VDD.n1116 59.488
R230 VDD.n730 VDD.n729 59.488
R231 VDD.n205 VDD.t42 55.465
R232 VDD.n179 VDD.t83 55.465
R233 VDD.n724 VDD.t14 55.106
R234 VDD.n802 VDD.t44 55.106
R235 VDD.n863 VDD.t24 55.106
R236 VDD.n924 VDD.t31 55.106
R237 VDD.n985 VDD.t77 55.106
R238 VDD.n1046 VDD.t79 55.106
R239 VDD.n1111 VDD.t40 55.106
R240 VDD.n1188 VDD.t22 55.106
R241 VDD.n1249 VDD.t27 55.106
R242 VDD.n1310 VDD.t3 55.106
R243 VDD.n1371 VDD.t20 55.106
R244 VDD.n652 VDD.t54 55.106
R245 VDD.n587 VDD.t82 55.106
R246 VDD.n510 VDD.t59 55.106
R247 VDD.n449 VDD.t26 55.106
R248 VDD.n388 VDD.t57 55.106
R249 VDD.n327 VDD.t48 55.106
R250 VDD.n266 VDD.t73 55.106
R251 VDD.n37 VDD.t12 55.106
R252 VDD.n24 VDD.t53 55.106
R253 VDD.n765 VDD.t49 55.106
R254 VDD.n1152 VDD.t10 55.106
R255 VDD.n551 VDD.t51 55.106
R256 VDD.n828 VDD.t9 55.106
R257 VDD.n889 VDD.t38 55.106
R258 VDD.n950 VDD.t47 55.106
R259 VDD.n1011 VDD.t80 55.106
R260 VDD.n1072 VDD.t37 55.106
R261 VDD.n1214 VDD.t4 55.106
R262 VDD.n1275 VDD.t2 55.106
R263 VDD.n1336 VDD.t17 55.106
R264 VDD.n687 VDD.t70 55.106
R265 VDD.n626 VDD.t21 55.106
R266 VDD.n484 VDD.t7 55.106
R267 VDD.n423 VDD.t67 55.106
R268 VDD.n362 VDD.t30 55.106
R269 VDD.n301 VDD.t41 55.106
R270 VDD.n240 VDD.t72 55.106
R271 VDD.n190 VDD.n189 41.183
R272 VDD.n735 VDD.n734 40.824
R273 VDD.n755 VDD.n754 40.824
R274 VDD.n818 VDD.n817 40.824
R275 VDD.n879 VDD.n878 40.824
R276 VDD.n940 VDD.n939 40.824
R277 VDD.n1001 VDD.n1000 40.824
R278 VDD.n1062 VDD.n1061 40.824
R279 VDD.n1122 VDD.n1121 40.824
R280 VDD.n1142 VDD.n1141 40.824
R281 VDD.n1204 VDD.n1203 40.824
R282 VDD.n1265 VDD.n1264 40.824
R283 VDD.n1326 VDD.n1325 40.824
R284 VDD.n1387 VDD.n1386 40.824
R285 VDD.n637 VDD.n636 40.824
R286 VDD.n576 VDD.n575 40.824
R287 VDD.n562 VDD.n561 40.824
R288 VDD.n495 VDD.n494 40.824
R289 VDD.n434 VDD.n433 40.824
R290 VDD.n373 VDD.n372 40.824
R291 VDD.n312 VDD.n311 40.824
R292 VDD.n251 VDD.n250 40.824
R293 VDD.n841 VDD.n840 36.774
R294 VDD.n902 VDD.n901 36.774
R295 VDD.n963 VDD.n962 36.774
R296 VDD.n1024 VDD.n1023 36.774
R297 VDD.n1085 VDD.n1084 36.774
R298 VDD.n1166 VDD.n1165 36.774
R299 VDD.n1227 VDD.n1226 36.774
R300 VDD.n1288 VDD.n1287 36.774
R301 VDD.n1349 VDD.n1348 36.774
R302 VDD.n665 VDD.n664 36.774
R303 VDD.n604 VDD.n603 36.774
R304 VDD.n523 VDD.n522 36.774
R305 VDD.n462 VDD.n461 36.774
R306 VDD.n401 VDD.n400 36.774
R307 VDD.n340 VDD.n339 36.774
R308 VDD.n279 VDD.n278 36.774
R309 VDD.n218 VDD.n217 36.774
R310 VDD.n157 VDD.n156 36.774
R311 VDD.n103 VDD.n102 36.774
R312 VDD.n48 VDD.n47 36.774
R313 VDD.n790 VDD.n789 36.774
R314 VDD.n185 VDD.n184 36.608
R315 VDD.n246 VDD.n245 36.608
R316 VDD.n307 VDD.n306 36.608
R317 VDD.n368 VDD.n367 36.608
R318 VDD.n429 VDD.n428 36.608
R319 VDD.n490 VDD.n489 36.608
R320 VDD.n632 VDD.n631 36.608
R321 VDD.n693 VDD.n692 36.608
R322 VDD.n1332 VDD.n1331 36.608
R323 VDD.n1271 VDD.n1270 36.608
R324 VDD.n1210 VDD.n1209 36.608
R325 VDD.n1068 VDD.n1067 36.608
R326 VDD.n1007 VDD.n1006 36.608
R327 VDD.n946 VDD.n945 36.608
R328 VDD.n885 VDD.n884 36.608
R329 VDD.n824 VDD.n823 36.608
R330 VDD.n201 VDD.n200 32.032
R331 VDD.n262 VDD.n261 32.032
R332 VDD.n323 VDD.n322 32.032
R333 VDD.n384 VDD.n383 32.032
R334 VDD.n445 VDD.n444 32.032
R335 VDD.n506 VDD.n505 32.032
R336 VDD.n648 VDD.n647 32.032
R337 VDD.n1377 VDD.n1376 32.032
R338 VDD.n1316 VDD.n1315 32.032
R339 VDD.n1255 VDD.n1254 32.032
R340 VDD.n1194 VDD.n1193 32.032
R341 VDD.n1052 VDD.n1051 32.032
R342 VDD.n991 VDD.n990 32.032
R343 VDD.n930 VDD.n929 32.032
R344 VDD.n869 VDD.n868 32.032
R345 VDD.n808 VDD.n807 32.032
R346 VDD.n559 VDD.n558 27.456
R347 VDD.n1139 VDD.n1138 27.456
R348 VDD.n752 VDD.n751 27.456
R349 VDD.n578 VDD.n577 22.88
R350 VDD.n1124 VDD.n1123 22.88
R351 VDD.n737 VDD.n736 22.88
R352 VDD.n718 VDD.n715 21.841
R353 VDD.n23 VDD.n20 21.841
R354 VDD.n734 VDD.t64 14.282
R355 VDD.n734 VDD.t56 14.282
R356 VDD.n754 VDD.t46 14.282
R357 VDD.n754 VDD.t60 14.282
R358 VDD.n817 VDD.t8 14.282
R359 VDD.n817 VDD.t11 14.282
R360 VDD.n878 VDD.t55 14.282
R361 VDD.n878 VDD.t76 14.282
R362 VDD.n939 VDD.t63 14.282
R363 VDD.n939 VDD.t66 14.282
R364 VDD.n1000 VDD.t81 14.282
R365 VDD.n1000 VDD.t62 14.282
R366 VDD.n1061 VDD.t75 14.282
R367 VDD.n1061 VDD.t13 14.282
R368 VDD.n1121 VDD.t18 14.282
R369 VDD.n1121 VDD.t33 14.282
R370 VDD.n1141 VDD.t74 14.282
R371 VDD.n1141 VDD.t35 14.282
R372 VDD.n1203 VDD.t5 14.282
R373 VDD.n1203 VDD.t32 14.282
R374 VDD.n1264 VDD.t78 14.282
R375 VDD.n1264 VDD.t16 14.282
R376 VDD.n1325 VDD.t1 14.282
R377 VDD.n1325 VDD.t15 14.282
R378 VDD.n1386 VDD.t45 14.282
R379 VDD.n1386 VDD.t36 14.282
R380 VDD.n636 VDD.t52 14.282
R381 VDD.n636 VDD.t39 14.282
R382 VDD.n575 VDD.t50 14.282
R383 VDD.n575 VDD.t69 14.282
R384 VDD.n561 VDD.t65 14.282
R385 VDD.n561 VDD.t28 14.282
R386 VDD.n494 VDD.t6 14.282
R387 VDD.n494 VDD.t29 14.282
R388 VDD.n433 VDD.t0 14.282
R389 VDD.n433 VDD.t61 14.282
R390 VDD.n372 VDD.t25 14.282
R391 VDD.n372 VDD.t43 14.282
R392 VDD.n311 VDD.t34 14.282
R393 VDD.n311 VDD.t58 14.282
R394 VDD.n250 VDD.t68 14.282
R395 VDD.n250 VDD.t19 14.282
R396 VDD.n189 VDD.t71 14.282
R397 VDD.n189 VDD.t23 14.282
R398 VDD.n715 VDD.n698 14.167
R399 VDD.n698 VDD.n697 14.167
R400 VDD.n856 VDD.n838 14.167
R401 VDD.n838 VDD.n837 14.167
R402 VDD.n917 VDD.n899 14.167
R403 VDD.n899 VDD.n898 14.167
R404 VDD.n978 VDD.n960 14.167
R405 VDD.n960 VDD.n959 14.167
R406 VDD.n1039 VDD.n1021 14.167
R407 VDD.n1021 VDD.n1020 14.167
R408 VDD.n1100 VDD.n1082 14.167
R409 VDD.n1082 VDD.n1081 14.167
R410 VDD.n1181 VDD.n1163 14.167
R411 VDD.n1163 VDD.n1162 14.167
R412 VDD.n1242 VDD.n1224 14.167
R413 VDD.n1224 VDD.n1223 14.167
R414 VDD.n1303 VDD.n1285 14.167
R415 VDD.n1285 VDD.n1284 14.167
R416 VDD.n1364 VDD.n1346 14.167
R417 VDD.n1346 VDD.n1345 14.167
R418 VDD.n680 VDD.n662 14.167
R419 VDD.n662 VDD.n661 14.167
R420 VDD.n619 VDD.n601 14.167
R421 VDD.n601 VDD.n600 14.167
R422 VDD.n538 VDD.n520 14.167
R423 VDD.n520 VDD.n519 14.167
R424 VDD.n477 VDD.n459 14.167
R425 VDD.n459 VDD.n458 14.167
R426 VDD.n416 VDD.n398 14.167
R427 VDD.n398 VDD.n397 14.167
R428 VDD.n355 VDD.n337 14.167
R429 VDD.n337 VDD.n336 14.167
R430 VDD.n294 VDD.n276 14.167
R431 VDD.n276 VDD.n275 14.167
R432 VDD.n233 VDD.n215 14.167
R433 VDD.n215 VDD.n214 14.167
R434 VDD.n172 VDD.n154 14.167
R435 VDD.n154 VDD.n153 14.167
R436 VDD.n118 VDD.n100 14.167
R437 VDD.n100 VDD.n99 14.167
R438 VDD.n64 VDD.n45 14.167
R439 VDD.n45 VDD.n44 14.167
R440 VDD.n795 VDD.n776 14.167
R441 VDD.n776 VDD.n775 14.167
R442 VDD.n20 VDD.n19 14.167
R443 VDD.n19 VDD.n17 14.167
R444 VDD.n69 VDD.n65 14.167
R445 VDD.n123 VDD.n119 14.167
R446 VDD.n177 VDD.n173 14.167
R447 VDD.n238 VDD.n234 14.167
R448 VDD.n299 VDD.n295 14.167
R449 VDD.n360 VDD.n356 14.167
R450 VDD.n421 VDD.n417 14.167
R451 VDD.n482 VDD.n478 14.167
R452 VDD.n543 VDD.n539 14.167
R453 VDD.n624 VDD.n620 14.167
R454 VDD.n685 VDD.n681 14.167
R455 VDD.n1369 VDD.n1365 14.167
R456 VDD.n1308 VDD.n1304 14.167
R457 VDD.n1247 VDD.n1243 14.167
R458 VDD.n1186 VDD.n1182 14.167
R459 VDD.n1105 VDD.n1101 14.167
R460 VDD.n1044 VDD.n1040 14.167
R461 VDD.n983 VDD.n979 14.167
R462 VDD.n922 VDD.n918 14.167
R463 VDD.n861 VDD.n857 14.167
R464 VDD.n800 VDD.n796 14.167
R465 VDD.n571 VDD.n570 13.728
R466 VDD.n1129 VDD.n1128 13.728
R467 VDD.n742 VDD.n741 13.728
R468 VDD.n23 VDD.n22 13.653
R469 VDD.n22 VDD.n21 13.653
R470 VDD.n28 VDD.n27 13.653
R471 VDD.n27 VDD.n26 13.653
R472 VDD.n32 VDD.n31 13.653
R473 VDD.n31 VDD.n30 13.653
R474 VDD.n38 VDD.n36 13.653
R475 VDD.n36 VDD.n35 13.653
R476 VDD.n42 VDD.n41 13.653
R477 VDD.n41 VDD.n40 13.653
R478 VDD.n69 VDD.n68 13.653
R479 VDD.n68 VDD.n67 13.653
R480 VDD.n73 VDD.n72 13.653
R481 VDD.n72 VDD.n71 13.653
R482 VDD.n77 VDD.n76 13.653
R483 VDD.n76 VDD.n75 13.653
R484 VDD.n81 VDD.n80 13.653
R485 VDD.n80 VDD.n79 13.653
R486 VDD.n85 VDD.n84 13.653
R487 VDD.n84 VDD.n83 13.653
R488 VDD.n89 VDD.n88 13.653
R489 VDD.n88 VDD.n87 13.653
R490 VDD.n93 VDD.n92 13.653
R491 VDD.n92 VDD.n91 13.653
R492 VDD.n97 VDD.n96 13.653
R493 VDD.n96 VDD.n95 13.653
R494 VDD.n123 VDD.n122 13.653
R495 VDD.n122 VDD.n121 13.653
R496 VDD.n127 VDD.n126 13.653
R497 VDD.n126 VDD.n125 13.653
R498 VDD.n131 VDD.n130 13.653
R499 VDD.n130 VDD.n129 13.653
R500 VDD.n135 VDD.n134 13.653
R501 VDD.n134 VDD.n133 13.653
R502 VDD.n139 VDD.n138 13.653
R503 VDD.n138 VDD.n137 13.653
R504 VDD.n143 VDD.n142 13.653
R505 VDD.n142 VDD.n141 13.653
R506 VDD.n147 VDD.n146 13.653
R507 VDD.n146 VDD.n145 13.653
R508 VDD.n151 VDD.n150 13.653
R509 VDD.n150 VDD.n149 13.653
R510 VDD.n177 VDD.n176 13.653
R511 VDD.n176 VDD.n175 13.653
R512 VDD.n182 VDD.n181 13.653
R513 VDD.n181 VDD.n180 13.653
R514 VDD.n187 VDD.n186 13.653
R515 VDD.n186 VDD.n185 13.653
R516 VDD.n193 VDD.n192 13.653
R517 VDD.n192 VDD.n191 13.653
R518 VDD.n198 VDD.n197 13.653
R519 VDD.n197 VDD.n196 13.653
R520 VDD.n203 VDD.n202 13.653
R521 VDD.n202 VDD.n201 13.653
R522 VDD.n208 VDD.n207 13.653
R523 VDD.n207 VDD.n206 13.653
R524 VDD.n212 VDD.n211 13.653
R525 VDD.n211 VDD.n210 13.653
R526 VDD.n238 VDD.n237 13.653
R527 VDD.n237 VDD.n236 13.653
R528 VDD.n243 VDD.n242 13.653
R529 VDD.n242 VDD.n241 13.653
R530 VDD.n248 VDD.n247 13.653
R531 VDD.n247 VDD.n246 13.653
R532 VDD.n254 VDD.n253 13.653
R533 VDD.n253 VDD.n252 13.653
R534 VDD.n259 VDD.n258 13.653
R535 VDD.n258 VDD.n257 13.653
R536 VDD.n264 VDD.n263 13.653
R537 VDD.n263 VDD.n262 13.653
R538 VDD.n269 VDD.n268 13.653
R539 VDD.n268 VDD.n267 13.653
R540 VDD.n273 VDD.n272 13.653
R541 VDD.n272 VDD.n271 13.653
R542 VDD.n299 VDD.n298 13.653
R543 VDD.n298 VDD.n297 13.653
R544 VDD.n304 VDD.n303 13.653
R545 VDD.n303 VDD.n302 13.653
R546 VDD.n309 VDD.n308 13.653
R547 VDD.n308 VDD.n307 13.653
R548 VDD.n315 VDD.n314 13.653
R549 VDD.n314 VDD.n313 13.653
R550 VDD.n320 VDD.n319 13.653
R551 VDD.n319 VDD.n318 13.653
R552 VDD.n325 VDD.n324 13.653
R553 VDD.n324 VDD.n323 13.653
R554 VDD.n330 VDD.n329 13.653
R555 VDD.n329 VDD.n328 13.653
R556 VDD.n334 VDD.n333 13.653
R557 VDD.n333 VDD.n332 13.653
R558 VDD.n360 VDD.n359 13.653
R559 VDD.n359 VDD.n358 13.653
R560 VDD.n365 VDD.n364 13.653
R561 VDD.n364 VDD.n363 13.653
R562 VDD.n370 VDD.n369 13.653
R563 VDD.n369 VDD.n368 13.653
R564 VDD.n376 VDD.n375 13.653
R565 VDD.n375 VDD.n374 13.653
R566 VDD.n381 VDD.n380 13.653
R567 VDD.n380 VDD.n379 13.653
R568 VDD.n386 VDD.n385 13.653
R569 VDD.n385 VDD.n384 13.653
R570 VDD.n391 VDD.n390 13.653
R571 VDD.n390 VDD.n389 13.653
R572 VDD.n395 VDD.n394 13.653
R573 VDD.n394 VDD.n393 13.653
R574 VDD.n421 VDD.n420 13.653
R575 VDD.n420 VDD.n419 13.653
R576 VDD.n426 VDD.n425 13.653
R577 VDD.n425 VDD.n424 13.653
R578 VDD.n431 VDD.n430 13.653
R579 VDD.n430 VDD.n429 13.653
R580 VDD.n437 VDD.n436 13.653
R581 VDD.n436 VDD.n435 13.653
R582 VDD.n442 VDD.n441 13.653
R583 VDD.n441 VDD.n440 13.653
R584 VDD.n447 VDD.n446 13.653
R585 VDD.n446 VDD.n445 13.653
R586 VDD.n452 VDD.n451 13.653
R587 VDD.n451 VDD.n450 13.653
R588 VDD.n456 VDD.n455 13.653
R589 VDD.n455 VDD.n454 13.653
R590 VDD.n482 VDD.n481 13.653
R591 VDD.n481 VDD.n480 13.653
R592 VDD.n487 VDD.n486 13.653
R593 VDD.n486 VDD.n485 13.653
R594 VDD.n492 VDD.n491 13.653
R595 VDD.n491 VDD.n490 13.653
R596 VDD.n498 VDD.n497 13.653
R597 VDD.n497 VDD.n496 13.653
R598 VDD.n503 VDD.n502 13.653
R599 VDD.n502 VDD.n501 13.653
R600 VDD.n508 VDD.n507 13.653
R601 VDD.n507 VDD.n506 13.653
R602 VDD.n513 VDD.n512 13.653
R603 VDD.n512 VDD.n511 13.653
R604 VDD.n517 VDD.n516 13.653
R605 VDD.n516 VDD.n515 13.653
R606 VDD.n543 VDD.n542 13.653
R607 VDD.n542 VDD.n541 13.653
R608 VDD.n547 VDD.n546 13.653
R609 VDD.n546 VDD.n545 13.653
R610 VDD.n551 VDD.n550 13.653
R611 VDD.n550 VDD.n549 13.653
R612 VDD.n556 VDD.n555 13.653
R613 VDD.n555 VDD.n554 13.653
R614 VDD.n563 VDD.n560 13.653
R615 VDD.n560 VDD.n559 13.653
R616 VDD.n568 VDD.n567 13.653
R617 VDD.n567 VDD.n566 13.653
R618 VDD.n573 VDD.n572 13.653
R619 VDD.n572 VDD.n571 13.653
R620 VDD.n580 VDD.n579 13.653
R621 VDD.n579 VDD.n578 13.653
R622 VDD.n585 VDD.n584 13.653
R623 VDD.n584 VDD.n583 13.653
R624 VDD.n590 VDD.n589 13.653
R625 VDD.n589 VDD.n588 13.653
R626 VDD.n594 VDD.n593 13.653
R627 VDD.n593 VDD.n592 13.653
R628 VDD.n598 VDD.n597 13.653
R629 VDD.n597 VDD.n596 13.653
R630 VDD.n624 VDD.n623 13.653
R631 VDD.n623 VDD.n622 13.653
R632 VDD.n629 VDD.n628 13.653
R633 VDD.n628 VDD.n627 13.653
R634 VDD.n634 VDD.n633 13.653
R635 VDD.n633 VDD.n632 13.653
R636 VDD.n640 VDD.n639 13.653
R637 VDD.n639 VDD.n638 13.653
R638 VDD.n645 VDD.n644 13.653
R639 VDD.n644 VDD.n643 13.653
R640 VDD.n650 VDD.n649 13.653
R641 VDD.n649 VDD.n648 13.653
R642 VDD.n655 VDD.n654 13.653
R643 VDD.n654 VDD.n653 13.653
R644 VDD.n659 VDD.n658 13.653
R645 VDD.n658 VDD.n657 13.653
R646 VDD.n685 VDD.n684 13.653
R647 VDD.n684 VDD.n683 13.653
R648 VDD.n690 VDD.n689 13.653
R649 VDD.n689 VDD.n688 13.653
R650 VDD.n695 VDD.n694 13.653
R651 VDD.n694 VDD.n693 13.653
R652 VDD.n1390 VDD.n1389 13.653
R653 VDD.n1389 VDD.n1388 13.653
R654 VDD.n1384 VDD.n1383 13.653
R655 VDD.n1383 VDD.n1382 13.653
R656 VDD.n1379 VDD.n1378 13.653
R657 VDD.n1378 VDD.n1377 13.653
R658 VDD.n1374 VDD.n1373 13.653
R659 VDD.n1373 VDD.n1372 13.653
R660 VDD.n1369 VDD.n1368 13.653
R661 VDD.n1368 VDD.n1367 13.653
R662 VDD.n1343 VDD.n1342 13.653
R663 VDD.n1342 VDD.n1341 13.653
R664 VDD.n1339 VDD.n1338 13.653
R665 VDD.n1338 VDD.n1337 13.653
R666 VDD.n1334 VDD.n1333 13.653
R667 VDD.n1333 VDD.n1332 13.653
R668 VDD.n1329 VDD.n1328 13.653
R669 VDD.n1328 VDD.n1327 13.653
R670 VDD.n1323 VDD.n1322 13.653
R671 VDD.n1322 VDD.n1321 13.653
R672 VDD.n1318 VDD.n1317 13.653
R673 VDD.n1317 VDD.n1316 13.653
R674 VDD.n1313 VDD.n1312 13.653
R675 VDD.n1312 VDD.n1311 13.653
R676 VDD.n1308 VDD.n1307 13.653
R677 VDD.n1307 VDD.n1306 13.653
R678 VDD.n1282 VDD.n1281 13.653
R679 VDD.n1281 VDD.n1280 13.653
R680 VDD.n1278 VDD.n1277 13.653
R681 VDD.n1277 VDD.n1276 13.653
R682 VDD.n1273 VDD.n1272 13.653
R683 VDD.n1272 VDD.n1271 13.653
R684 VDD.n1268 VDD.n1267 13.653
R685 VDD.n1267 VDD.n1266 13.653
R686 VDD.n1262 VDD.n1261 13.653
R687 VDD.n1261 VDD.n1260 13.653
R688 VDD.n1257 VDD.n1256 13.653
R689 VDD.n1256 VDD.n1255 13.653
R690 VDD.n1252 VDD.n1251 13.653
R691 VDD.n1251 VDD.n1250 13.653
R692 VDD.n1247 VDD.n1246 13.653
R693 VDD.n1246 VDD.n1245 13.653
R694 VDD.n1221 VDD.n1220 13.653
R695 VDD.n1220 VDD.n1219 13.653
R696 VDD.n1217 VDD.n1216 13.653
R697 VDD.n1216 VDD.n1215 13.653
R698 VDD.n1212 VDD.n1211 13.653
R699 VDD.n1211 VDD.n1210 13.653
R700 VDD.n1207 VDD.n1206 13.653
R701 VDD.n1206 VDD.n1205 13.653
R702 VDD.n1201 VDD.n1200 13.653
R703 VDD.n1200 VDD.n1199 13.653
R704 VDD.n1196 VDD.n1195 13.653
R705 VDD.n1195 VDD.n1194 13.653
R706 VDD.n1191 VDD.n1190 13.653
R707 VDD.n1190 VDD.n1189 13.653
R708 VDD.n1186 VDD.n1185 13.653
R709 VDD.n1185 VDD.n1184 13.653
R710 VDD.n1160 VDD.n1159 13.653
R711 VDD.n1159 VDD.n1158 13.653
R712 VDD.n1156 VDD.n1155 13.653
R713 VDD.n1155 VDD.n1154 13.653
R714 VDD.n1152 VDD.n1151 13.653
R715 VDD.n1151 VDD.n1150 13.653
R716 VDD.n1148 VDD.n1147 13.653
R717 VDD.n1147 VDD.n1146 13.653
R718 VDD.n1143 VDD.n1140 13.653
R719 VDD.n1140 VDD.n1139 13.653
R720 VDD.n1136 VDD.n1135 13.653
R721 VDD.n1135 VDD.n1134 13.653
R722 VDD.n1131 VDD.n1130 13.653
R723 VDD.n1130 VDD.n1129 13.653
R724 VDD.n1126 VDD.n1125 13.653
R725 VDD.n1125 VDD.n1124 13.653
R726 VDD.n1119 VDD.n1118 13.653
R727 VDD.n1118 VDD.n1117 13.653
R728 VDD.n1114 VDD.n1113 13.653
R729 VDD.n1113 VDD.n1112 13.653
R730 VDD.n1109 VDD.n1108 13.653
R731 VDD.n1108 VDD.n1107 13.653
R732 VDD.n1105 VDD.n1104 13.653
R733 VDD.n1104 VDD.n1103 13.653
R734 VDD.n1079 VDD.n1078 13.653
R735 VDD.n1078 VDD.n1077 13.653
R736 VDD.n1075 VDD.n1074 13.653
R737 VDD.n1074 VDD.n1073 13.653
R738 VDD.n1070 VDD.n1069 13.653
R739 VDD.n1069 VDD.n1068 13.653
R740 VDD.n1065 VDD.n1064 13.653
R741 VDD.n1064 VDD.n1063 13.653
R742 VDD.n1059 VDD.n1058 13.653
R743 VDD.n1058 VDD.n1057 13.653
R744 VDD.n1054 VDD.n1053 13.653
R745 VDD.n1053 VDD.n1052 13.653
R746 VDD.n1049 VDD.n1048 13.653
R747 VDD.n1048 VDD.n1047 13.653
R748 VDD.n1044 VDD.n1043 13.653
R749 VDD.n1043 VDD.n1042 13.653
R750 VDD.n1018 VDD.n1017 13.653
R751 VDD.n1017 VDD.n1016 13.653
R752 VDD.n1014 VDD.n1013 13.653
R753 VDD.n1013 VDD.n1012 13.653
R754 VDD.n1009 VDD.n1008 13.653
R755 VDD.n1008 VDD.n1007 13.653
R756 VDD.n1004 VDD.n1003 13.653
R757 VDD.n1003 VDD.n1002 13.653
R758 VDD.n998 VDD.n997 13.653
R759 VDD.n997 VDD.n996 13.653
R760 VDD.n993 VDD.n992 13.653
R761 VDD.n992 VDD.n991 13.653
R762 VDD.n988 VDD.n987 13.653
R763 VDD.n987 VDD.n986 13.653
R764 VDD.n983 VDD.n982 13.653
R765 VDD.n982 VDD.n981 13.653
R766 VDD.n957 VDD.n956 13.653
R767 VDD.n956 VDD.n955 13.653
R768 VDD.n953 VDD.n952 13.653
R769 VDD.n952 VDD.n951 13.653
R770 VDD.n948 VDD.n947 13.653
R771 VDD.n947 VDD.n946 13.653
R772 VDD.n943 VDD.n942 13.653
R773 VDD.n942 VDD.n941 13.653
R774 VDD.n937 VDD.n936 13.653
R775 VDD.n936 VDD.n935 13.653
R776 VDD.n932 VDD.n931 13.653
R777 VDD.n931 VDD.n930 13.653
R778 VDD.n927 VDD.n926 13.653
R779 VDD.n926 VDD.n925 13.653
R780 VDD.n922 VDD.n921 13.653
R781 VDD.n921 VDD.n920 13.653
R782 VDD.n896 VDD.n895 13.653
R783 VDD.n895 VDD.n894 13.653
R784 VDD.n892 VDD.n891 13.653
R785 VDD.n891 VDD.n890 13.653
R786 VDD.n887 VDD.n886 13.653
R787 VDD.n886 VDD.n885 13.653
R788 VDD.n882 VDD.n881 13.653
R789 VDD.n881 VDD.n880 13.653
R790 VDD.n876 VDD.n875 13.653
R791 VDD.n875 VDD.n874 13.653
R792 VDD.n871 VDD.n870 13.653
R793 VDD.n870 VDD.n869 13.653
R794 VDD.n866 VDD.n865 13.653
R795 VDD.n865 VDD.n864 13.653
R796 VDD.n861 VDD.n860 13.653
R797 VDD.n860 VDD.n859 13.653
R798 VDD.n835 VDD.n834 13.653
R799 VDD.n834 VDD.n833 13.653
R800 VDD.n831 VDD.n830 13.653
R801 VDD.n830 VDD.n829 13.653
R802 VDD.n826 VDD.n825 13.653
R803 VDD.n825 VDD.n824 13.653
R804 VDD.n821 VDD.n820 13.653
R805 VDD.n820 VDD.n819 13.653
R806 VDD.n815 VDD.n814 13.653
R807 VDD.n814 VDD.n813 13.653
R808 VDD.n810 VDD.n809 13.653
R809 VDD.n809 VDD.n808 13.653
R810 VDD.n805 VDD.n804 13.653
R811 VDD.n804 VDD.n803 13.653
R812 VDD.n800 VDD.n799 13.653
R813 VDD.n799 VDD.n798 13.653
R814 VDD.n773 VDD.n772 13.653
R815 VDD.n772 VDD.n771 13.653
R816 VDD.n769 VDD.n768 13.653
R817 VDD.n768 VDD.n767 13.653
R818 VDD.n765 VDD.n764 13.653
R819 VDD.n764 VDD.n763 13.653
R820 VDD.n761 VDD.n760 13.653
R821 VDD.n760 VDD.n759 13.653
R822 VDD.n756 VDD.n753 13.653
R823 VDD.n753 VDD.n752 13.653
R824 VDD.n749 VDD.n748 13.653
R825 VDD.n748 VDD.n747 13.653
R826 VDD.n744 VDD.n743 13.653
R827 VDD.n743 VDD.n742 13.653
R828 VDD.n739 VDD.n738 13.653
R829 VDD.n738 VDD.n737 13.653
R830 VDD.n732 VDD.n731 13.653
R831 VDD.n731 VDD.n730 13.653
R832 VDD.n727 VDD.n726 13.653
R833 VDD.n726 VDD.n725 13.653
R834 VDD.n722 VDD.n721 13.653
R835 VDD.n721 VDD.n720 13.653
R836 VDD.n718 VDD.n717 13.653
R837 VDD.n717 VDD.n716 13.653
R838 VDD.n4 VDD.n2 12.915
R839 VDD.n4 VDD.n3 12.66
R840 VDD.n13 VDD.n12 12.343
R841 VDD.n11 VDD.n10 12.343
R842 VDD.n7 VDD.n6 12.343
R843 VDD.n566 VDD.n565 9.152
R844 VDD.n1134 VDD.n1133 9.152
R845 VDD.n747 VDD.n746 9.152
R846 VDD.n193 VDD.n190 8.658
R847 VDD.n254 VDD.n251 8.658
R848 VDD.n315 VDD.n312 8.658
R849 VDD.n376 VDD.n373 8.658
R850 VDD.n437 VDD.n434 8.658
R851 VDD.n498 VDD.n495 8.658
R852 VDD.n640 VDD.n637 8.658
R853 VDD.n1390 VDD.n1387 8.658
R854 VDD.n1329 VDD.n1326 8.658
R855 VDD.n1268 VDD.n1265 8.658
R856 VDD.n1207 VDD.n1204 8.658
R857 VDD.n1065 VDD.n1062 8.658
R858 VDD.n1004 VDD.n1001 8.658
R859 VDD.n943 VDD.n940 8.658
R860 VDD.n882 VDD.n879 8.658
R861 VDD.n821 VDD.n818 8.658
R862 VDD.n857 VDD.n856 7.674
R863 VDD.n918 VDD.n917 7.674
R864 VDD.n979 VDD.n978 7.674
R865 VDD.n1040 VDD.n1039 7.674
R866 VDD.n1101 VDD.n1100 7.674
R867 VDD.n1182 VDD.n1181 7.674
R868 VDD.n1243 VDD.n1242 7.674
R869 VDD.n1304 VDD.n1303 7.674
R870 VDD.n1365 VDD.n1364 7.674
R871 VDD.n681 VDD.n680 7.674
R872 VDD.n620 VDD.n619 7.674
R873 VDD.n539 VDD.n538 7.674
R874 VDD.n478 VDD.n477 7.674
R875 VDD.n417 VDD.n416 7.674
R876 VDD.n356 VDD.n355 7.674
R877 VDD.n295 VDD.n294 7.674
R878 VDD.n234 VDD.n233 7.674
R879 VDD.n173 VDD.n172 7.674
R880 VDD.n119 VDD.n118 7.674
R881 VDD.n65 VDD.n64 7.674
R882 VDD.n796 VDD.n795 7.674
R883 VDD.n59 VDD.n58 7.5
R884 VDD.n53 VDD.n52 7.5
R885 VDD.n55 VDD.n54 7.5
R886 VDD.n50 VDD.n49 7.5
R887 VDD.n64 VDD.n63 7.5
R888 VDD.n113 VDD.n112 7.5
R889 VDD.n107 VDD.n106 7.5
R890 VDD.n109 VDD.n108 7.5
R891 VDD.n115 VDD.n105 7.5
R892 VDD.n115 VDD.n103 7.5
R893 VDD.n118 VDD.n117 7.5
R894 VDD.n167 VDD.n166 7.5
R895 VDD.n161 VDD.n160 7.5
R896 VDD.n163 VDD.n162 7.5
R897 VDD.n169 VDD.n159 7.5
R898 VDD.n169 VDD.n157 7.5
R899 VDD.n172 VDD.n171 7.5
R900 VDD.n228 VDD.n227 7.5
R901 VDD.n222 VDD.n221 7.5
R902 VDD.n224 VDD.n223 7.5
R903 VDD.n230 VDD.n220 7.5
R904 VDD.n230 VDD.n218 7.5
R905 VDD.n233 VDD.n232 7.5
R906 VDD.n289 VDD.n288 7.5
R907 VDD.n283 VDD.n282 7.5
R908 VDD.n285 VDD.n284 7.5
R909 VDD.n291 VDD.n281 7.5
R910 VDD.n291 VDD.n279 7.5
R911 VDD.n294 VDD.n293 7.5
R912 VDD.n350 VDD.n349 7.5
R913 VDD.n344 VDD.n343 7.5
R914 VDD.n346 VDD.n345 7.5
R915 VDD.n352 VDD.n342 7.5
R916 VDD.n352 VDD.n340 7.5
R917 VDD.n355 VDD.n354 7.5
R918 VDD.n411 VDD.n410 7.5
R919 VDD.n405 VDD.n404 7.5
R920 VDD.n407 VDD.n406 7.5
R921 VDD.n413 VDD.n403 7.5
R922 VDD.n413 VDD.n401 7.5
R923 VDD.n416 VDD.n415 7.5
R924 VDD.n472 VDD.n471 7.5
R925 VDD.n466 VDD.n465 7.5
R926 VDD.n468 VDD.n467 7.5
R927 VDD.n474 VDD.n464 7.5
R928 VDD.n474 VDD.n462 7.5
R929 VDD.n477 VDD.n476 7.5
R930 VDD.n533 VDD.n532 7.5
R931 VDD.n527 VDD.n526 7.5
R932 VDD.n529 VDD.n528 7.5
R933 VDD.n535 VDD.n525 7.5
R934 VDD.n535 VDD.n523 7.5
R935 VDD.n538 VDD.n537 7.5
R936 VDD.n614 VDD.n613 7.5
R937 VDD.n608 VDD.n607 7.5
R938 VDD.n610 VDD.n609 7.5
R939 VDD.n616 VDD.n606 7.5
R940 VDD.n616 VDD.n604 7.5
R941 VDD.n619 VDD.n618 7.5
R942 VDD.n675 VDD.n674 7.5
R943 VDD.n669 VDD.n668 7.5
R944 VDD.n671 VDD.n670 7.5
R945 VDD.n677 VDD.n667 7.5
R946 VDD.n677 VDD.n665 7.5
R947 VDD.n680 VDD.n679 7.5
R948 VDD.n1359 VDD.n1358 7.5
R949 VDD.n1353 VDD.n1352 7.5
R950 VDD.n1355 VDD.n1354 7.5
R951 VDD.n1361 VDD.n1351 7.5
R952 VDD.n1361 VDD.n1349 7.5
R953 VDD.n1364 VDD.n1363 7.5
R954 VDD.n1298 VDD.n1297 7.5
R955 VDD.n1292 VDD.n1291 7.5
R956 VDD.n1294 VDD.n1293 7.5
R957 VDD.n1300 VDD.n1290 7.5
R958 VDD.n1300 VDD.n1288 7.5
R959 VDD.n1303 VDD.n1302 7.5
R960 VDD.n1237 VDD.n1236 7.5
R961 VDD.n1231 VDD.n1230 7.5
R962 VDD.n1233 VDD.n1232 7.5
R963 VDD.n1239 VDD.n1229 7.5
R964 VDD.n1239 VDD.n1227 7.5
R965 VDD.n1242 VDD.n1241 7.5
R966 VDD.n1176 VDD.n1175 7.5
R967 VDD.n1170 VDD.n1169 7.5
R968 VDD.n1172 VDD.n1171 7.5
R969 VDD.n1178 VDD.n1168 7.5
R970 VDD.n1178 VDD.n1166 7.5
R971 VDD.n1181 VDD.n1180 7.5
R972 VDD.n1095 VDD.n1094 7.5
R973 VDD.n1089 VDD.n1088 7.5
R974 VDD.n1091 VDD.n1090 7.5
R975 VDD.n1097 VDD.n1087 7.5
R976 VDD.n1097 VDD.n1085 7.5
R977 VDD.n1100 VDD.n1099 7.5
R978 VDD.n1034 VDD.n1033 7.5
R979 VDD.n1028 VDD.n1027 7.5
R980 VDD.n1030 VDD.n1029 7.5
R981 VDD.n1036 VDD.n1026 7.5
R982 VDD.n1036 VDD.n1024 7.5
R983 VDD.n1039 VDD.n1038 7.5
R984 VDD.n973 VDD.n972 7.5
R985 VDD.n967 VDD.n966 7.5
R986 VDD.n969 VDD.n968 7.5
R987 VDD.n975 VDD.n965 7.5
R988 VDD.n975 VDD.n963 7.5
R989 VDD.n978 VDD.n977 7.5
R990 VDD.n912 VDD.n911 7.5
R991 VDD.n906 VDD.n905 7.5
R992 VDD.n908 VDD.n907 7.5
R993 VDD.n914 VDD.n904 7.5
R994 VDD.n914 VDD.n902 7.5
R995 VDD.n917 VDD.n916 7.5
R996 VDD.n851 VDD.n850 7.5
R997 VDD.n845 VDD.n844 7.5
R998 VDD.n847 VDD.n846 7.5
R999 VDD.n853 VDD.n843 7.5
R1000 VDD.n853 VDD.n841 7.5
R1001 VDD.n856 VDD.n855 7.5
R1002 VDD.n780 VDD.n779 7.5
R1003 VDD.n783 VDD.n782 7.5
R1004 VDD.n785 VDD.n784 7.5
R1005 VDD.n788 VDD.n787 7.5
R1006 VDD.n795 VDD.n794 7.5
R1007 VDD.n710 VDD.n709 7.5
R1008 VDD.n704 VDD.n703 7.5
R1009 VDD.n706 VDD.n705 7.5
R1010 VDD.n712 VDD.n702 7.5
R1011 VDD.n712 VDD.n700 7.5
R1012 VDD.n715 VDD.n714 7.5
R1013 VDD.n20 VDD.n16 7.5
R1014 VDD.n2 VDD.n1 7.5
R1015 VDD.n6 VDD.n5 7.5
R1016 VDD.n10 VDD.n9 7.5
R1017 VDD.n19 VDD.n18 7.5
R1018 VDD.n14 VDD.n0 7.5
R1019 VDD.n51 VDD.n48 6.772
R1020 VDD.n62 VDD.n46 6.772
R1021 VDD.n60 VDD.n57 6.772
R1022 VDD.n56 VDD.n53 6.772
R1023 VDD.n116 VDD.n101 6.772
R1024 VDD.n114 VDD.n111 6.772
R1025 VDD.n110 VDD.n107 6.772
R1026 VDD.n170 VDD.n155 6.772
R1027 VDD.n168 VDD.n165 6.772
R1028 VDD.n164 VDD.n161 6.772
R1029 VDD.n231 VDD.n216 6.772
R1030 VDD.n229 VDD.n226 6.772
R1031 VDD.n225 VDD.n222 6.772
R1032 VDD.n292 VDD.n277 6.772
R1033 VDD.n290 VDD.n287 6.772
R1034 VDD.n286 VDD.n283 6.772
R1035 VDD.n353 VDD.n338 6.772
R1036 VDD.n351 VDD.n348 6.772
R1037 VDD.n347 VDD.n344 6.772
R1038 VDD.n414 VDD.n399 6.772
R1039 VDD.n412 VDD.n409 6.772
R1040 VDD.n408 VDD.n405 6.772
R1041 VDD.n475 VDD.n460 6.772
R1042 VDD.n473 VDD.n470 6.772
R1043 VDD.n469 VDD.n466 6.772
R1044 VDD.n536 VDD.n521 6.772
R1045 VDD.n534 VDD.n531 6.772
R1046 VDD.n530 VDD.n527 6.772
R1047 VDD.n617 VDD.n602 6.772
R1048 VDD.n615 VDD.n612 6.772
R1049 VDD.n611 VDD.n608 6.772
R1050 VDD.n678 VDD.n663 6.772
R1051 VDD.n676 VDD.n673 6.772
R1052 VDD.n672 VDD.n669 6.772
R1053 VDD.n1362 VDD.n1347 6.772
R1054 VDD.n1360 VDD.n1357 6.772
R1055 VDD.n1356 VDD.n1353 6.772
R1056 VDD.n1301 VDD.n1286 6.772
R1057 VDD.n1299 VDD.n1296 6.772
R1058 VDD.n1295 VDD.n1292 6.772
R1059 VDD.n1240 VDD.n1225 6.772
R1060 VDD.n1238 VDD.n1235 6.772
R1061 VDD.n1234 VDD.n1231 6.772
R1062 VDD.n1179 VDD.n1164 6.772
R1063 VDD.n1177 VDD.n1174 6.772
R1064 VDD.n1173 VDD.n1170 6.772
R1065 VDD.n1098 VDD.n1083 6.772
R1066 VDD.n1096 VDD.n1093 6.772
R1067 VDD.n1092 VDD.n1089 6.772
R1068 VDD.n1037 VDD.n1022 6.772
R1069 VDD.n1035 VDD.n1032 6.772
R1070 VDD.n1031 VDD.n1028 6.772
R1071 VDD.n976 VDD.n961 6.772
R1072 VDD.n974 VDD.n971 6.772
R1073 VDD.n970 VDD.n967 6.772
R1074 VDD.n915 VDD.n900 6.772
R1075 VDD.n913 VDD.n910 6.772
R1076 VDD.n909 VDD.n906 6.772
R1077 VDD.n854 VDD.n839 6.772
R1078 VDD.n852 VDD.n849 6.772
R1079 VDD.n848 VDD.n845 6.772
R1080 VDD.n713 VDD.n699 6.772
R1081 VDD.n711 VDD.n708 6.772
R1082 VDD.n707 VDD.n704 6.772
R1083 VDD.n51 VDD.n50 6.772
R1084 VDD.n56 VDD.n55 6.772
R1085 VDD.n60 VDD.n59 6.772
R1086 VDD.n63 VDD.n62 6.772
R1087 VDD.n110 VDD.n109 6.772
R1088 VDD.n114 VDD.n113 6.772
R1089 VDD.n117 VDD.n116 6.772
R1090 VDD.n164 VDD.n163 6.772
R1091 VDD.n168 VDD.n167 6.772
R1092 VDD.n171 VDD.n170 6.772
R1093 VDD.n225 VDD.n224 6.772
R1094 VDD.n229 VDD.n228 6.772
R1095 VDD.n232 VDD.n231 6.772
R1096 VDD.n286 VDD.n285 6.772
R1097 VDD.n290 VDD.n289 6.772
R1098 VDD.n293 VDD.n292 6.772
R1099 VDD.n347 VDD.n346 6.772
R1100 VDD.n351 VDD.n350 6.772
R1101 VDD.n354 VDD.n353 6.772
R1102 VDD.n408 VDD.n407 6.772
R1103 VDD.n412 VDD.n411 6.772
R1104 VDD.n415 VDD.n414 6.772
R1105 VDD.n469 VDD.n468 6.772
R1106 VDD.n473 VDD.n472 6.772
R1107 VDD.n476 VDD.n475 6.772
R1108 VDD.n530 VDD.n529 6.772
R1109 VDD.n534 VDD.n533 6.772
R1110 VDD.n537 VDD.n536 6.772
R1111 VDD.n611 VDD.n610 6.772
R1112 VDD.n615 VDD.n614 6.772
R1113 VDD.n618 VDD.n617 6.772
R1114 VDD.n672 VDD.n671 6.772
R1115 VDD.n676 VDD.n675 6.772
R1116 VDD.n679 VDD.n678 6.772
R1117 VDD.n1356 VDD.n1355 6.772
R1118 VDD.n1360 VDD.n1359 6.772
R1119 VDD.n1363 VDD.n1362 6.772
R1120 VDD.n1295 VDD.n1294 6.772
R1121 VDD.n1299 VDD.n1298 6.772
R1122 VDD.n1302 VDD.n1301 6.772
R1123 VDD.n1234 VDD.n1233 6.772
R1124 VDD.n1238 VDD.n1237 6.772
R1125 VDD.n1241 VDD.n1240 6.772
R1126 VDD.n1173 VDD.n1172 6.772
R1127 VDD.n1177 VDD.n1176 6.772
R1128 VDD.n1180 VDD.n1179 6.772
R1129 VDD.n1092 VDD.n1091 6.772
R1130 VDD.n1096 VDD.n1095 6.772
R1131 VDD.n1099 VDD.n1098 6.772
R1132 VDD.n1031 VDD.n1030 6.772
R1133 VDD.n1035 VDD.n1034 6.772
R1134 VDD.n1038 VDD.n1037 6.772
R1135 VDD.n970 VDD.n969 6.772
R1136 VDD.n974 VDD.n973 6.772
R1137 VDD.n977 VDD.n976 6.772
R1138 VDD.n909 VDD.n908 6.772
R1139 VDD.n913 VDD.n912 6.772
R1140 VDD.n916 VDD.n915 6.772
R1141 VDD.n848 VDD.n847 6.772
R1142 VDD.n852 VDD.n851 6.772
R1143 VDD.n855 VDD.n854 6.772
R1144 VDD.n707 VDD.n706 6.772
R1145 VDD.n711 VDD.n710 6.772
R1146 VDD.n714 VDD.n713 6.772
R1147 VDD.n794 VDD.n793 6.772
R1148 VDD.n781 VDD.n778 6.772
R1149 VDD.n786 VDD.n783 6.772
R1150 VDD.n791 VDD.n788 6.772
R1151 VDD.n791 VDD.n790 6.772
R1152 VDD.n786 VDD.n785 6.772
R1153 VDD.n781 VDD.n780 6.772
R1154 VDD.n793 VDD.n777 6.772
R1155 VDD.n580 VDD.n576 6.69
R1156 VDD.n1126 VDD.n1122 6.69
R1157 VDD.n739 VDD.n735 6.69
R1158 VDD.n16 VDD.n15 6.458
R1159 VDD.n563 VDD.n562 6.296
R1160 VDD.n1143 VDD.n1142 6.296
R1161 VDD.n756 VDD.n755 6.296
R1162 VDD.n105 VDD.n104 6.202
R1163 VDD.n159 VDD.n158 6.202
R1164 VDD.n220 VDD.n219 6.202
R1165 VDD.n281 VDD.n280 6.202
R1166 VDD.n342 VDD.n341 6.202
R1167 VDD.n403 VDD.n402 6.202
R1168 VDD.n464 VDD.n463 6.202
R1169 VDD.n525 VDD.n524 6.202
R1170 VDD.n606 VDD.n605 6.202
R1171 VDD.n667 VDD.n666 6.202
R1172 VDD.n1351 VDD.n1350 6.202
R1173 VDD.n1290 VDD.n1289 6.202
R1174 VDD.n1229 VDD.n1228 6.202
R1175 VDD.n1168 VDD.n1167 6.202
R1176 VDD.n1087 VDD.n1086 6.202
R1177 VDD.n1026 VDD.n1025 6.202
R1178 VDD.n965 VDD.n964 6.202
R1179 VDD.n904 VDD.n903 6.202
R1180 VDD.n843 VDD.n842 6.202
R1181 VDD.n702 VDD.n701 6.202
R1182 VDD.n196 VDD.n195 4.576
R1183 VDD.n257 VDD.n256 4.576
R1184 VDD.n318 VDD.n317 4.576
R1185 VDD.n379 VDD.n378 4.576
R1186 VDD.n440 VDD.n439 4.576
R1187 VDD.n501 VDD.n500 4.576
R1188 VDD.n643 VDD.n642 4.576
R1189 VDD.n1382 VDD.n1381 4.576
R1190 VDD.n1321 VDD.n1320 4.576
R1191 VDD.n1260 VDD.n1259 4.576
R1192 VDD.n1199 VDD.n1198 4.576
R1193 VDD.n1057 VDD.n1056 4.576
R1194 VDD.n996 VDD.n995 4.576
R1195 VDD.n935 VDD.n934 4.576
R1196 VDD.n874 VDD.n873 4.576
R1197 VDD.n813 VDD.n812 4.576
R1198 VDD.n208 VDD.n205 2.754
R1199 VDD.n269 VDD.n266 2.754
R1200 VDD.n330 VDD.n327 2.754
R1201 VDD.n391 VDD.n388 2.754
R1202 VDD.n452 VDD.n449 2.754
R1203 VDD.n513 VDD.n510 2.754
R1204 VDD.n655 VDD.n652 2.754
R1205 VDD.n1374 VDD.n1371 2.754
R1206 VDD.n1313 VDD.n1310 2.754
R1207 VDD.n1252 VDD.n1249 2.754
R1208 VDD.n1191 VDD.n1188 2.754
R1209 VDD.n1049 VDD.n1046 2.754
R1210 VDD.n988 VDD.n985 2.754
R1211 VDD.n927 VDD.n924 2.754
R1212 VDD.n866 VDD.n863 2.754
R1213 VDD.n805 VDD.n802 2.754
R1214 VDD.n182 VDD.n179 2.361
R1215 VDD.n243 VDD.n240 2.361
R1216 VDD.n304 VDD.n301 2.361
R1217 VDD.n365 VDD.n362 2.361
R1218 VDD.n426 VDD.n423 2.361
R1219 VDD.n487 VDD.n484 2.361
R1220 VDD.n629 VDD.n626 2.361
R1221 VDD.n690 VDD.n687 2.361
R1222 VDD.n1339 VDD.n1336 2.361
R1223 VDD.n1278 VDD.n1275 2.361
R1224 VDD.n1217 VDD.n1214 2.361
R1225 VDD.n1075 VDD.n1072 2.361
R1226 VDD.n1014 VDD.n1011 2.361
R1227 VDD.n953 VDD.n950 2.361
R1228 VDD.n892 VDD.n889 2.361
R1229 VDD.n831 VDD.n828 2.361
R1230 VDD.n28 VDD.n24 1.967
R1231 VDD.n38 VDD.n37 1.967
R1232 VDD.n14 VDD.n7 1.329
R1233 VDD.n14 VDD.n8 1.329
R1234 VDD.n14 VDD.n11 1.329
R1235 VDD.n14 VDD.n13 1.329
R1236 VDD.n15 VDD.n14 0.696
R1237 VDD.n14 VDD.n4 0.696
R1238 VDD.n590 VDD.n587 0.393
R1239 VDD.n1114 VDD.n1111 0.393
R1240 VDD.n727 VDD.n724 0.393
R1241 VDD.n61 VDD.n60 0.365
R1242 VDD.n61 VDD.n56 0.365
R1243 VDD.n61 VDD.n51 0.365
R1244 VDD.n62 VDD.n61 0.365
R1245 VDD.n115 VDD.n114 0.365
R1246 VDD.n115 VDD.n110 0.365
R1247 VDD.n116 VDD.n115 0.365
R1248 VDD.n169 VDD.n168 0.365
R1249 VDD.n169 VDD.n164 0.365
R1250 VDD.n170 VDD.n169 0.365
R1251 VDD.n230 VDD.n229 0.365
R1252 VDD.n230 VDD.n225 0.365
R1253 VDD.n231 VDD.n230 0.365
R1254 VDD.n291 VDD.n290 0.365
R1255 VDD.n291 VDD.n286 0.365
R1256 VDD.n292 VDD.n291 0.365
R1257 VDD.n352 VDD.n351 0.365
R1258 VDD.n352 VDD.n347 0.365
R1259 VDD.n353 VDD.n352 0.365
R1260 VDD.n413 VDD.n412 0.365
R1261 VDD.n413 VDD.n408 0.365
R1262 VDD.n414 VDD.n413 0.365
R1263 VDD.n474 VDD.n473 0.365
R1264 VDD.n474 VDD.n469 0.365
R1265 VDD.n475 VDD.n474 0.365
R1266 VDD.n535 VDD.n534 0.365
R1267 VDD.n535 VDD.n530 0.365
R1268 VDD.n536 VDD.n535 0.365
R1269 VDD.n616 VDD.n615 0.365
R1270 VDD.n616 VDD.n611 0.365
R1271 VDD.n617 VDD.n616 0.365
R1272 VDD.n677 VDD.n676 0.365
R1273 VDD.n677 VDD.n672 0.365
R1274 VDD.n678 VDD.n677 0.365
R1275 VDD.n1361 VDD.n1360 0.365
R1276 VDD.n1361 VDD.n1356 0.365
R1277 VDD.n1362 VDD.n1361 0.365
R1278 VDD.n1300 VDD.n1299 0.365
R1279 VDD.n1300 VDD.n1295 0.365
R1280 VDD.n1301 VDD.n1300 0.365
R1281 VDD.n1239 VDD.n1238 0.365
R1282 VDD.n1239 VDD.n1234 0.365
R1283 VDD.n1240 VDD.n1239 0.365
R1284 VDD.n1178 VDD.n1177 0.365
R1285 VDD.n1178 VDD.n1173 0.365
R1286 VDD.n1179 VDD.n1178 0.365
R1287 VDD.n1097 VDD.n1096 0.365
R1288 VDD.n1097 VDD.n1092 0.365
R1289 VDD.n1098 VDD.n1097 0.365
R1290 VDD.n1036 VDD.n1035 0.365
R1291 VDD.n1036 VDD.n1031 0.365
R1292 VDD.n1037 VDD.n1036 0.365
R1293 VDD.n975 VDD.n974 0.365
R1294 VDD.n975 VDD.n970 0.365
R1295 VDD.n976 VDD.n975 0.365
R1296 VDD.n914 VDD.n913 0.365
R1297 VDD.n914 VDD.n909 0.365
R1298 VDD.n915 VDD.n914 0.365
R1299 VDD.n853 VDD.n852 0.365
R1300 VDD.n853 VDD.n848 0.365
R1301 VDD.n854 VDD.n853 0.365
R1302 VDD.n712 VDD.n711 0.365
R1303 VDD.n712 VDD.n707 0.365
R1304 VDD.n713 VDD.n712 0.365
R1305 VDD.n792 VDD.n791 0.365
R1306 VDD.n792 VDD.n786 0.365
R1307 VDD.n792 VDD.n781 0.365
R1308 VDD.n793 VDD.n792 0.365
R1309 VDD.n70 VDD.n43 0.29
R1310 VDD.n124 VDD.n98 0.29
R1311 VDD.n178 VDD.n152 0.29
R1312 VDD.n239 VDD.n213 0.29
R1313 VDD.n300 VDD.n274 0.29
R1314 VDD.n361 VDD.n335 0.29
R1315 VDD.n422 VDD.n396 0.29
R1316 VDD.n483 VDD.n457 0.29
R1317 VDD.n544 VDD.n518 0.29
R1318 VDD.n625 VDD.n599 0.29
R1319 VDD.n686 VDD.n660 0.29
R1320 VDD.n1370 VDD.n1344 0.29
R1321 VDD.n1309 VDD.n1283 0.29
R1322 VDD.n1248 VDD.n1222 0.29
R1323 VDD.n1187 VDD.n1161 0.29
R1324 VDD.n1106 VDD.n1080 0.29
R1325 VDD.n1045 VDD.n1019 0.29
R1326 VDD.n984 VDD.n958 0.29
R1327 VDD.n923 VDD.n897 0.29
R1328 VDD.n862 VDD.n836 0.29
R1329 VDD.n801 VDD.n774 0.29
R1330 VDD.n719 VDD 0.207
R1331 VDD.n574 VDD.n569 0.197
R1332 VDD.n1137 VDD.n1132 0.197
R1333 VDD.n750 VDD.n745 0.197
R1334 VDD.n86 VDD.n82 0.181
R1335 VDD.n140 VDD.n136 0.181
R1336 VDD.n199 VDD.n194 0.181
R1337 VDD.n260 VDD.n255 0.181
R1338 VDD.n321 VDD.n316 0.181
R1339 VDD.n382 VDD.n377 0.181
R1340 VDD.n443 VDD.n438 0.181
R1341 VDD.n504 VDD.n499 0.181
R1342 VDD.n646 VDD.n641 0.181
R1343 VDD.n1391 VDD.n1385 0.181
R1344 VDD.n1330 VDD.n1324 0.181
R1345 VDD.n1269 VDD.n1263 0.181
R1346 VDD.n1208 VDD.n1202 0.181
R1347 VDD.n1066 VDD.n1060 0.181
R1348 VDD.n1005 VDD.n999 0.181
R1349 VDD.n944 VDD.n938 0.181
R1350 VDD.n883 VDD.n877 0.181
R1351 VDD.n822 VDD.n816 0.181
R1352 VDD.n33 VDD.n29 0.157
R1353 VDD.n39 VDD.n33 0.157
R1354 VDD.n43 VDD.n39 0.145
R1355 VDD.n74 VDD.n70 0.145
R1356 VDD.n78 VDD.n74 0.145
R1357 VDD.n82 VDD.n78 0.145
R1358 VDD.n90 VDD.n86 0.145
R1359 VDD.n94 VDD.n90 0.145
R1360 VDD.n98 VDD.n94 0.145
R1361 VDD.n128 VDD.n124 0.145
R1362 VDD.n132 VDD.n128 0.145
R1363 VDD.n136 VDD.n132 0.145
R1364 VDD.n144 VDD.n140 0.145
R1365 VDD.n148 VDD.n144 0.145
R1366 VDD.n152 VDD.n148 0.145
R1367 VDD.n183 VDD.n178 0.145
R1368 VDD.n188 VDD.n183 0.145
R1369 VDD.n194 VDD.n188 0.145
R1370 VDD.n204 VDD.n199 0.145
R1371 VDD.n209 VDD.n204 0.145
R1372 VDD.n213 VDD.n209 0.145
R1373 VDD.n244 VDD.n239 0.145
R1374 VDD.n249 VDD.n244 0.145
R1375 VDD.n255 VDD.n249 0.145
R1376 VDD.n265 VDD.n260 0.145
R1377 VDD.n270 VDD.n265 0.145
R1378 VDD.n274 VDD.n270 0.145
R1379 VDD.n305 VDD.n300 0.145
R1380 VDD.n310 VDD.n305 0.145
R1381 VDD.n316 VDD.n310 0.145
R1382 VDD.n326 VDD.n321 0.145
R1383 VDD.n331 VDD.n326 0.145
R1384 VDD.n335 VDD.n331 0.145
R1385 VDD.n366 VDD.n361 0.145
R1386 VDD.n371 VDD.n366 0.145
R1387 VDD.n377 VDD.n371 0.145
R1388 VDD.n387 VDD.n382 0.145
R1389 VDD.n392 VDD.n387 0.145
R1390 VDD.n396 VDD.n392 0.145
R1391 VDD.n427 VDD.n422 0.145
R1392 VDD.n432 VDD.n427 0.145
R1393 VDD.n438 VDD.n432 0.145
R1394 VDD.n448 VDD.n443 0.145
R1395 VDD.n453 VDD.n448 0.145
R1396 VDD.n457 VDD.n453 0.145
R1397 VDD.n488 VDD.n483 0.145
R1398 VDD.n493 VDD.n488 0.145
R1399 VDD.n499 VDD.n493 0.145
R1400 VDD.n509 VDD.n504 0.145
R1401 VDD.n514 VDD.n509 0.145
R1402 VDD.n518 VDD.n514 0.145
R1403 VDD.n548 VDD.n544 0.145
R1404 VDD.n552 VDD.n548 0.145
R1405 VDD.n557 VDD.n552 0.145
R1406 VDD.n564 VDD.n557 0.145
R1407 VDD.n569 VDD.n564 0.145
R1408 VDD.n581 VDD.n574 0.145
R1409 VDD.n586 VDD.n581 0.145
R1410 VDD.n591 VDD.n586 0.145
R1411 VDD.n595 VDD.n591 0.145
R1412 VDD.n599 VDD.n595 0.145
R1413 VDD.n630 VDD.n625 0.145
R1414 VDD.n635 VDD.n630 0.145
R1415 VDD.n641 VDD.n635 0.145
R1416 VDD.n651 VDD.n646 0.145
R1417 VDD.n656 VDD.n651 0.145
R1418 VDD.n660 VDD.n656 0.145
R1419 VDD.n691 VDD.n686 0.145
R1420 VDD.n696 VDD.n691 0.145
R1421 VDD.n1385 VDD.n1380 0.145
R1422 VDD.n1380 VDD.n1375 0.145
R1423 VDD.n1375 VDD.n1370 0.145
R1424 VDD.n1344 VDD.n1340 0.145
R1425 VDD.n1340 VDD.n1335 0.145
R1426 VDD.n1335 VDD.n1330 0.145
R1427 VDD.n1324 VDD.n1319 0.145
R1428 VDD.n1319 VDD.n1314 0.145
R1429 VDD.n1314 VDD.n1309 0.145
R1430 VDD.n1283 VDD.n1279 0.145
R1431 VDD.n1279 VDD.n1274 0.145
R1432 VDD.n1274 VDD.n1269 0.145
R1433 VDD.n1263 VDD.n1258 0.145
R1434 VDD.n1258 VDD.n1253 0.145
R1435 VDD.n1253 VDD.n1248 0.145
R1436 VDD.n1222 VDD.n1218 0.145
R1437 VDD.n1218 VDD.n1213 0.145
R1438 VDD.n1213 VDD.n1208 0.145
R1439 VDD.n1202 VDD.n1197 0.145
R1440 VDD.n1197 VDD.n1192 0.145
R1441 VDD.n1192 VDD.n1187 0.145
R1442 VDD.n1161 VDD.n1157 0.145
R1443 VDD.n1157 VDD.n1153 0.145
R1444 VDD.n1153 VDD.n1149 0.145
R1445 VDD.n1149 VDD.n1144 0.145
R1446 VDD.n1144 VDD.n1137 0.145
R1447 VDD.n1132 VDD.n1127 0.145
R1448 VDD.n1127 VDD.n1120 0.145
R1449 VDD.n1120 VDD.n1115 0.145
R1450 VDD.n1115 VDD.n1110 0.145
R1451 VDD.n1110 VDD.n1106 0.145
R1452 VDD.n1080 VDD.n1076 0.145
R1453 VDD.n1076 VDD.n1071 0.145
R1454 VDD.n1071 VDD.n1066 0.145
R1455 VDD.n1060 VDD.n1055 0.145
R1456 VDD.n1055 VDD.n1050 0.145
R1457 VDD.n1050 VDD.n1045 0.145
R1458 VDD.n1019 VDD.n1015 0.145
R1459 VDD.n1015 VDD.n1010 0.145
R1460 VDD.n1010 VDD.n1005 0.145
R1461 VDD.n999 VDD.n994 0.145
R1462 VDD.n994 VDD.n989 0.145
R1463 VDD.n989 VDD.n984 0.145
R1464 VDD.n958 VDD.n954 0.145
R1465 VDD.n954 VDD.n949 0.145
R1466 VDD.n949 VDD.n944 0.145
R1467 VDD.n938 VDD.n933 0.145
R1468 VDD.n933 VDD.n928 0.145
R1469 VDD.n928 VDD.n923 0.145
R1470 VDD.n897 VDD.n893 0.145
R1471 VDD.n893 VDD.n888 0.145
R1472 VDD.n888 VDD.n883 0.145
R1473 VDD.n877 VDD.n872 0.145
R1474 VDD.n872 VDD.n867 0.145
R1475 VDD.n867 VDD.n862 0.145
R1476 VDD.n836 VDD.n832 0.145
R1477 VDD.n832 VDD.n827 0.145
R1478 VDD.n827 VDD.n822 0.145
R1479 VDD.n816 VDD.n811 0.145
R1480 VDD.n811 VDD.n806 0.145
R1481 VDD.n806 VDD.n801 0.145
R1482 VDD.n774 VDD.n770 0.145
R1483 VDD.n770 VDD.n766 0.145
R1484 VDD.n766 VDD.n762 0.145
R1485 VDD.n762 VDD.n757 0.145
R1486 VDD.n757 VDD.n750 0.145
R1487 VDD.n745 VDD.n740 0.145
R1488 VDD.n740 VDD.n733 0.145
R1489 VDD.n733 VDD.n728 0.145
R1490 VDD.n728 VDD.n723 0.145
R1491 VDD.n723 VDD.n719 0.145
R1492 VDD VDD.n696 0.086
R1493 VDD VDD.n1391 0.058
R1494 a_599_989.n0 a_599_989.t9 480.392
R1495 a_599_989.n2 a_599_989.t10 454.685
R1496 a_599_989.n2 a_599_989.t7 428.979
R1497 a_599_989.n0 a_599_989.t5 403.272
R1498 a_599_989.n1 a_599_989.t8 283.48
R1499 a_599_989.n3 a_599_989.t6 237.959
R1500 a_599_989.n9 a_599_989.n8 210.592
R1501 a_599_989.n11 a_599_989.n9 152.499
R1502 a_599_989.n3 a_599_989.n2 98.447
R1503 a_599_989.n1 a_599_989.n0 98.447
R1504 a_599_989.n4 a_599_989.n3 78.947
R1505 a_599_989.n4 a_599_989.n1 77.315
R1506 a_599_989.n11 a_599_989.n10 76.002
R1507 a_599_989.n9 a_599_989.n4 76
R1508 a_599_989.n8 a_599_989.n7 30
R1509 a_599_989.n6 a_599_989.n5 24.383
R1510 a_599_989.n8 a_599_989.n6 23.684
R1511 a_599_989.n10 a_599_989.t3 14.282
R1512 a_599_989.n10 a_599_989.t4 14.282
R1513 a_599_989.n12 a_599_989.t0 14.282
R1514 a_599_989.t1 a_599_989.n12 14.282
R1515 a_599_989.n12 a_599_989.n11 12.848
R1516 a_3303_411.n4 a_3303_411.t8 512.525
R1517 a_3303_411.n3 a_3303_411.t10 512.525
R1518 a_3303_411.n8 a_3303_411.t12 472.359
R1519 a_3303_411.n8 a_3303_411.t7 384.527
R1520 a_3303_411.n4 a_3303_411.t11 371.139
R1521 a_3303_411.n3 a_3303_411.t9 371.139
R1522 a_3303_411.n5 a_3303_411.n4 265.439
R1523 a_3303_411.n9 a_3303_411.t6 214.619
R1524 a_3303_411.n13 a_3303_411.n11 190.561
R1525 a_3303_411.n7 a_3303_411.n3 185.78
R1526 a_3303_411.n11 a_3303_411.n2 179.052
R1527 a_3303_411.n5 a_3303_411.t5 176.995
R1528 a_3303_411.n6 a_3303_411.t13 170.569
R1529 a_3303_411.n6 a_3303_411.n5 153.043
R1530 a_3303_411.n9 a_3303_411.n8 136.613
R1531 a_3303_411.n10 a_3303_411.n7 112.41
R1532 a_3303_411.n7 a_3303_411.n6 79.658
R1533 a_3303_411.n10 a_3303_411.n9 78.947
R1534 a_3303_411.n2 a_3303_411.n1 76.002
R1535 a_3303_411.n11 a_3303_411.n10 76
R1536 a_3303_411.n13 a_3303_411.n12 15.218
R1537 a_3303_411.n0 a_3303_411.t2 14.282
R1538 a_3303_411.n0 a_3303_411.t3 14.282
R1539 a_3303_411.n1 a_3303_411.t0 14.282
R1540 a_3303_411.n1 a_3303_411.t4 14.282
R1541 a_3303_411.n2 a_3303_411.n0 12.85
R1542 a_3303_411.n14 a_3303_411.n13 12.014
R1543 a_14320_101.t0 a_14320_101.n1 93.333
R1544 a_14320_101.n4 a_14320_101.n2 55.07
R1545 a_14320_101.t0 a_14320_101.n0 8.137
R1546 a_14320_101.n4 a_14320_101.n3 4.619
R1547 a_14320_101.t0 a_14320_101.n4 0.071
R1548 GND.n30 GND.n29 219.745
R1549 GND.n60 GND.n58 219.745
R1550 GND.n90 GND.n88 219.745
R1551 GND.n400 GND.n399 219.745
R1552 GND.n433 GND.n431 219.745
R1553 GND.n466 GND.n464 219.745
R1554 GND.n496 GND.n494 219.745
R1555 GND.n526 GND.n524 219.745
R1556 GND.n559 GND.n557 219.745
R1557 GND.n601 GND.n599 219.745
R1558 GND.n631 GND.n629 219.745
R1559 GND.n661 GND.n659 219.745
R1560 GND.n691 GND.n689 219.745
R1561 GND.n348 GND.n346 219.745
R1562 GND.n318 GND.n316 219.745
R1563 GND.n276 GND.n274 219.745
R1564 GND.n246 GND.n244 219.745
R1565 GND.n213 GND.n211 219.745
R1566 GND.n183 GND.n181 219.745
R1567 GND.n153 GND.n151 219.745
R1568 GND.n120 GND.n119 219.745
R1569 GND.n307 GND.n306 85.559
R1570 GND.n568 GND.n567 85.559
R1571 GND.n367 GND.n366 85.559
R1572 GND.n30 GND.n28 85.529
R1573 GND.n60 GND.n59 85.529
R1574 GND.n90 GND.n89 85.529
R1575 GND.n400 GND.n398 85.529
R1576 GND.n433 GND.n432 85.529
R1577 GND.n466 GND.n465 85.529
R1578 GND.n496 GND.n495 85.529
R1579 GND.n526 GND.n525 85.529
R1580 GND.n559 GND.n558 85.529
R1581 GND.n601 GND.n600 85.529
R1582 GND.n631 GND.n630 85.529
R1583 GND.n661 GND.n660 85.529
R1584 GND.n691 GND.n690 85.529
R1585 GND.n348 GND.n347 85.529
R1586 GND.n318 GND.n317 85.529
R1587 GND.n276 GND.n275 85.529
R1588 GND.n246 GND.n245 85.529
R1589 GND.n213 GND.n212 85.529
R1590 GND.n183 GND.n182 85.529
R1591 GND.n153 GND.n152 85.529
R1592 GND.n120 GND.n118 85.529
R1593 GND.n78 GND.n77 84.842
R1594 GND.n108 GND.n107 84.842
R1595 GND.n171 GND.n170 84.842
R1596 GND.n201 GND.n200 84.842
R1597 GND.n264 GND.n263 84.842
R1598 GND.n336 GND.n335 84.842
R1599 GND.n669 GND.n668 84.842
R1600 GND.n639 GND.n638 84.842
R1601 GND.n609 GND.n608 84.842
R1602 GND.n504 GND.n503 84.842
R1603 GND.n474 GND.n473 84.842
R1604 GND.n48 GND.n47 84.842
R1605 GND.n9 GND.n1 76.145
R1606 GND.n361 GND.n360 76
R1607 GND.n73 GND.n72 76
R1608 GND.n76 GND.n75 76
R1609 GND.n81 GND.n80 76
R1610 GND.n84 GND.n83 76
R1611 GND.n87 GND.n86 76
R1612 GND.n94 GND.n93 76
R1613 GND.n97 GND.n96 76
R1614 GND.n100 GND.n99 76
R1615 GND.n103 GND.n102 76
R1616 GND.n106 GND.n105 76
R1617 GND.n111 GND.n110 76
R1618 GND.n114 GND.n113 76
R1619 GND.n117 GND.n116 76
R1620 GND.n124 GND.n123 76
R1621 GND.n127 GND.n126 76
R1622 GND.n130 GND.n129 76
R1623 GND.n133 GND.n132 76
R1624 GND.n136 GND.n135 76
R1625 GND.n144 GND.n143 76
R1626 GND.n147 GND.n146 76
R1627 GND.n150 GND.n149 76
R1628 GND.n157 GND.n156 76
R1629 GND.n160 GND.n159 76
R1630 GND.n163 GND.n162 76
R1631 GND.n166 GND.n165 76
R1632 GND.n169 GND.n168 76
R1633 GND.n174 GND.n173 76
R1634 GND.n177 GND.n176 76
R1635 GND.n180 GND.n179 76
R1636 GND.n187 GND.n186 76
R1637 GND.n190 GND.n189 76
R1638 GND.n193 GND.n192 76
R1639 GND.n196 GND.n195 76
R1640 GND.n199 GND.n198 76
R1641 GND.n204 GND.n203 76
R1642 GND.n207 GND.n206 76
R1643 GND.n210 GND.n209 76
R1644 GND.n217 GND.n216 76
R1645 GND.n220 GND.n219 76
R1646 GND.n223 GND.n222 76
R1647 GND.n226 GND.n225 76
R1648 GND.n229 GND.n228 76
R1649 GND.n237 GND.n236 76
R1650 GND.n240 GND.n239 76
R1651 GND.n243 GND.n242 76
R1652 GND.n250 GND.n249 76
R1653 GND.n253 GND.n252 76
R1654 GND.n256 GND.n255 76
R1655 GND.n259 GND.n258 76
R1656 GND.n262 GND.n261 76
R1657 GND.n267 GND.n266 76
R1658 GND.n270 GND.n269 76
R1659 GND.n273 GND.n272 76
R1660 GND.n280 GND.n279 76
R1661 GND.n283 GND.n282 76
R1662 GND.n286 GND.n285 76
R1663 GND.n289 GND.n288 76
R1664 GND.n292 GND.n291 76
R1665 GND.n295 GND.n294 76
R1666 GND.n298 GND.n297 76
R1667 GND.n301 GND.n300 76
R1668 GND.n304 GND.n303 76
R1669 GND.n309 GND.n308 76
R1670 GND.n312 GND.n311 76
R1671 GND.n315 GND.n314 76
R1672 GND.n322 GND.n321 76
R1673 GND.n325 GND.n324 76
R1674 GND.n328 GND.n327 76
R1675 GND.n331 GND.n330 76
R1676 GND.n334 GND.n333 76
R1677 GND.n339 GND.n338 76
R1678 GND.n342 GND.n341 76
R1679 GND.n345 GND.n344 76
R1680 GND.n352 GND.n351 76
R1681 GND.n355 GND.n354 76
R1682 GND.n358 GND.n357 76
R1683 GND.n711 GND.n710 76
R1684 GND.n708 GND.n707 76
R1685 GND.n705 GND.n704 76
R1686 GND.n697 GND.n696 76
R1687 GND.n694 GND.n693 76
R1688 GND.n687 GND.n686 76
R1689 GND.n684 GND.n683 76
R1690 GND.n681 GND.n680 76
R1691 GND.n678 GND.n677 76
R1692 GND.n675 GND.n674 76
R1693 GND.n672 GND.n671 76
R1694 GND.n667 GND.n666 76
R1695 GND.n664 GND.n663 76
R1696 GND.n657 GND.n656 76
R1697 GND.n654 GND.n653 76
R1698 GND.n651 GND.n650 76
R1699 GND.n648 GND.n647 76
R1700 GND.n645 GND.n644 76
R1701 GND.n642 GND.n641 76
R1702 GND.n637 GND.n636 76
R1703 GND.n634 GND.n633 76
R1704 GND.n627 GND.n626 76
R1705 GND.n624 GND.n623 76
R1706 GND.n621 GND.n620 76
R1707 GND.n618 GND.n617 76
R1708 GND.n615 GND.n614 76
R1709 GND.n612 GND.n611 76
R1710 GND.n607 GND.n606 76
R1711 GND.n604 GND.n603 76
R1712 GND.n597 GND.n596 76
R1713 GND.n594 GND.n593 76
R1714 GND.n591 GND.n590 76
R1715 GND.n588 GND.n587 76
R1716 GND.n585 GND.n584 76
R1717 GND.n582 GND.n581 76
R1718 GND.n579 GND.n578 76
R1719 GND.n576 GND.n575 76
R1720 GND.n573 GND.n572 76
R1721 GND.n570 GND.n569 76
R1722 GND.n565 GND.n564 76
R1723 GND.n562 GND.n561 76
R1724 GND.n555 GND.n554 76
R1725 GND.n552 GND.n551 76
R1726 GND.n549 GND.n548 76
R1727 GND.n546 GND.n545 76
R1728 GND.n543 GND.n542 76
R1729 GND.n540 GND.n539 76
R1730 GND.n532 GND.n531 76
R1731 GND.n529 GND.n528 76
R1732 GND.n522 GND.n521 76
R1733 GND.n519 GND.n518 76
R1734 GND.n516 GND.n515 76
R1735 GND.n513 GND.n512 76
R1736 GND.n510 GND.n509 76
R1737 GND.n507 GND.n506 76
R1738 GND.n502 GND.n501 76
R1739 GND.n499 GND.n498 76
R1740 GND.n492 GND.n491 76
R1741 GND.n489 GND.n488 76
R1742 GND.n486 GND.n485 76
R1743 GND.n483 GND.n482 76
R1744 GND.n480 GND.n479 76
R1745 GND.n477 GND.n476 76
R1746 GND.n472 GND.n471 76
R1747 GND.n469 GND.n468 76
R1748 GND.n462 GND.n461 76
R1749 GND.n459 GND.n458 76
R1750 GND.n456 GND.n455 76
R1751 GND.n453 GND.n452 76
R1752 GND.n450 GND.n449 76
R1753 GND.n447 GND.n446 76
R1754 GND.n439 GND.n438 76
R1755 GND.n436 GND.n435 76
R1756 GND.n429 GND.n428 76
R1757 GND.n426 GND.n425 76
R1758 GND.n423 GND.n422 76
R1759 GND.n420 GND.n419 76
R1760 GND.n417 GND.n416 76
R1761 GND.n414 GND.n413 76
R1762 GND.n406 GND.n405 76
R1763 GND.n403 GND.n402 76
R1764 GND.n396 GND.n395 76
R1765 GND.n393 GND.n392 76
R1766 GND.n390 GND.n389 76
R1767 GND.n387 GND.n386 76
R1768 GND.n384 GND.n383 76
R1769 GND.n381 GND.n380 76
R1770 GND.n378 GND.n377 76
R1771 GND.n375 GND.n374 76
R1772 GND.n372 GND.n371 76
R1773 GND.n369 GND.n368 76
R1774 GND.n364 GND.n363 76
R1775 GND.n9 GND.n8 76
R1776 GND.n17 GND.n16 76
R1777 GND.n24 GND.n23 76
R1778 GND.n27 GND.n26 76
R1779 GND.n34 GND.n33 76
R1780 GND.n37 GND.n36 76
R1781 GND.n40 GND.n39 76
R1782 GND.n43 GND.n42 76
R1783 GND.n46 GND.n45 76
R1784 GND.n51 GND.n50 76
R1785 GND.n54 GND.n53 76
R1786 GND.n57 GND.n56 76
R1787 GND.n64 GND.n63 76
R1788 GND.n67 GND.n66 76
R1789 GND.n70 GND.n69 76
R1790 GND.n141 GND.n140 63.835
R1791 GND.n234 GND.n233 63.835
R1792 GND.n702 GND.n701 63.835
R1793 GND.n537 GND.n536 63.835
R1794 GND.n444 GND.n443 63.835
R1795 GND.n411 GND.n410 63.835
R1796 GND.n5 GND.n4 35.01
R1797 GND.n3 GND.n2 29.127
R1798 GND.n140 GND.n139 28.421
R1799 GND.n233 GND.n232 28.421
R1800 GND.n701 GND.n700 28.421
R1801 GND.n536 GND.n535 28.421
R1802 GND.n443 GND.n442 28.421
R1803 GND.n410 GND.n409 28.421
R1804 GND.n140 GND.n138 25.263
R1805 GND.n233 GND.n231 25.263
R1806 GND.n701 GND.n699 25.263
R1807 GND.n536 GND.n534 25.263
R1808 GND.n443 GND.n441 25.263
R1809 GND.n410 GND.n408 25.263
R1810 GND.n138 GND.n137 24.383
R1811 GND.n231 GND.n230 24.383
R1812 GND.n699 GND.n698 24.383
R1813 GND.n534 GND.n533 24.383
R1814 GND.n441 GND.n440 24.383
R1815 GND.n408 GND.n407 24.383
R1816 GND.n12 GND.t1 20.794
R1817 GND.n6 GND.n5 19.735
R1818 GND.n14 GND.n13 19.735
R1819 GND.n21 GND.n20 19.735
R1820 GND.n5 GND.n3 19.017
R1821 GND.n33 GND.n31 14.167
R1822 GND.n63 GND.n61 14.167
R1823 GND.n93 GND.n91 14.167
R1824 GND.n123 GND.n121 14.167
R1825 GND.n156 GND.n154 14.167
R1826 GND.n186 GND.n184 14.167
R1827 GND.n216 GND.n214 14.167
R1828 GND.n249 GND.n247 14.167
R1829 GND.n279 GND.n277 14.167
R1830 GND.n321 GND.n319 14.167
R1831 GND.n351 GND.n349 14.167
R1832 GND.n693 GND.n692 14.167
R1833 GND.n663 GND.n662 14.167
R1834 GND.n633 GND.n632 14.167
R1835 GND.n603 GND.n602 14.167
R1836 GND.n561 GND.n560 14.167
R1837 GND.n528 GND.n527 14.167
R1838 GND.n498 GND.n497 14.167
R1839 GND.n468 GND.n467 14.167
R1840 GND.n435 GND.n434 14.167
R1841 GND.n402 GND.n401 14.167
R1842 GND.n363 GND.n362 13.653
R1843 GND.n368 GND.n365 13.653
R1844 GND.n371 GND.n370 13.653
R1845 GND.n374 GND.n373 13.653
R1846 GND.n377 GND.n376 13.653
R1847 GND.n380 GND.n379 13.653
R1848 GND.n383 GND.n382 13.653
R1849 GND.n386 GND.n385 13.653
R1850 GND.n389 GND.n388 13.653
R1851 GND.n392 GND.n391 13.653
R1852 GND.n395 GND.n394 13.653
R1853 GND.n402 GND.n397 13.653
R1854 GND.n405 GND.n404 13.653
R1855 GND.n413 GND.n412 13.653
R1856 GND.n416 GND.n415 13.653
R1857 GND.n419 GND.n418 13.653
R1858 GND.n422 GND.n421 13.653
R1859 GND.n425 GND.n424 13.653
R1860 GND.n428 GND.n427 13.653
R1861 GND.n435 GND.n430 13.653
R1862 GND.n438 GND.n437 13.653
R1863 GND.n446 GND.n445 13.653
R1864 GND.n449 GND.n448 13.653
R1865 GND.n452 GND.n451 13.653
R1866 GND.n455 GND.n454 13.653
R1867 GND.n458 GND.n457 13.653
R1868 GND.n461 GND.n460 13.653
R1869 GND.n468 GND.n463 13.653
R1870 GND.n471 GND.n470 13.653
R1871 GND.n476 GND.n475 13.653
R1872 GND.n479 GND.n478 13.653
R1873 GND.n482 GND.n481 13.653
R1874 GND.n485 GND.n484 13.653
R1875 GND.n488 GND.n487 13.653
R1876 GND.n491 GND.n490 13.653
R1877 GND.n498 GND.n493 13.653
R1878 GND.n501 GND.n500 13.653
R1879 GND.n506 GND.n505 13.653
R1880 GND.n509 GND.n508 13.653
R1881 GND.n512 GND.n511 13.653
R1882 GND.n515 GND.n514 13.653
R1883 GND.n518 GND.n517 13.653
R1884 GND.n521 GND.n520 13.653
R1885 GND.n528 GND.n523 13.653
R1886 GND.n531 GND.n530 13.653
R1887 GND.n539 GND.n538 13.653
R1888 GND.n542 GND.n541 13.653
R1889 GND.n545 GND.n544 13.653
R1890 GND.n548 GND.n547 13.653
R1891 GND.n551 GND.n550 13.653
R1892 GND.n554 GND.n553 13.653
R1893 GND.n561 GND.n556 13.653
R1894 GND.n564 GND.n563 13.653
R1895 GND.n569 GND.n566 13.653
R1896 GND.n572 GND.n571 13.653
R1897 GND.n575 GND.n574 13.653
R1898 GND.n578 GND.n577 13.653
R1899 GND.n581 GND.n580 13.653
R1900 GND.n584 GND.n583 13.653
R1901 GND.n587 GND.n586 13.653
R1902 GND.n590 GND.n589 13.653
R1903 GND.n593 GND.n592 13.653
R1904 GND.n596 GND.n595 13.653
R1905 GND.n603 GND.n598 13.653
R1906 GND.n606 GND.n605 13.653
R1907 GND.n611 GND.n610 13.653
R1908 GND.n614 GND.n613 13.653
R1909 GND.n617 GND.n616 13.653
R1910 GND.n620 GND.n619 13.653
R1911 GND.n623 GND.n622 13.653
R1912 GND.n626 GND.n625 13.653
R1913 GND.n633 GND.n628 13.653
R1914 GND.n636 GND.n635 13.653
R1915 GND.n641 GND.n640 13.653
R1916 GND.n644 GND.n643 13.653
R1917 GND.n647 GND.n646 13.653
R1918 GND.n650 GND.n649 13.653
R1919 GND.n653 GND.n652 13.653
R1920 GND.n656 GND.n655 13.653
R1921 GND.n663 GND.n658 13.653
R1922 GND.n666 GND.n665 13.653
R1923 GND.n671 GND.n670 13.653
R1924 GND.n674 GND.n673 13.653
R1925 GND.n677 GND.n676 13.653
R1926 GND.n680 GND.n679 13.653
R1927 GND.n683 GND.n682 13.653
R1928 GND.n686 GND.n685 13.653
R1929 GND.n693 GND.n688 13.653
R1930 GND.n696 GND.n695 13.653
R1931 GND.n704 GND.n703 13.653
R1932 GND.n707 GND.n706 13.653
R1933 GND.n710 GND.n709 13.653
R1934 GND.n357 GND.n356 13.653
R1935 GND.n354 GND.n353 13.653
R1936 GND.n351 GND.n350 13.653
R1937 GND.n344 GND.n343 13.653
R1938 GND.n341 GND.n340 13.653
R1939 GND.n338 GND.n337 13.653
R1940 GND.n333 GND.n332 13.653
R1941 GND.n330 GND.n329 13.653
R1942 GND.n327 GND.n326 13.653
R1943 GND.n324 GND.n323 13.653
R1944 GND.n321 GND.n320 13.653
R1945 GND.n314 GND.n313 13.653
R1946 GND.n311 GND.n310 13.653
R1947 GND.n308 GND.n305 13.653
R1948 GND.n303 GND.n302 13.653
R1949 GND.n300 GND.n299 13.653
R1950 GND.n297 GND.n296 13.653
R1951 GND.n294 GND.n293 13.653
R1952 GND.n291 GND.n290 13.653
R1953 GND.n288 GND.n287 13.653
R1954 GND.n285 GND.n284 13.653
R1955 GND.n282 GND.n281 13.653
R1956 GND.n279 GND.n278 13.653
R1957 GND.n272 GND.n271 13.653
R1958 GND.n269 GND.n268 13.653
R1959 GND.n266 GND.n265 13.653
R1960 GND.n261 GND.n260 13.653
R1961 GND.n258 GND.n257 13.653
R1962 GND.n255 GND.n254 13.653
R1963 GND.n252 GND.n251 13.653
R1964 GND.n249 GND.n248 13.653
R1965 GND.n242 GND.n241 13.653
R1966 GND.n239 GND.n238 13.653
R1967 GND.n236 GND.n235 13.653
R1968 GND.n228 GND.n227 13.653
R1969 GND.n225 GND.n224 13.653
R1970 GND.n222 GND.n221 13.653
R1971 GND.n219 GND.n218 13.653
R1972 GND.n216 GND.n215 13.653
R1973 GND.n209 GND.n208 13.653
R1974 GND.n206 GND.n205 13.653
R1975 GND.n203 GND.n202 13.653
R1976 GND.n198 GND.n197 13.653
R1977 GND.n195 GND.n194 13.653
R1978 GND.n192 GND.n191 13.653
R1979 GND.n189 GND.n188 13.653
R1980 GND.n186 GND.n185 13.653
R1981 GND.n179 GND.n178 13.653
R1982 GND.n176 GND.n175 13.653
R1983 GND.n173 GND.n172 13.653
R1984 GND.n168 GND.n167 13.653
R1985 GND.n165 GND.n164 13.653
R1986 GND.n162 GND.n161 13.653
R1987 GND.n159 GND.n158 13.653
R1988 GND.n156 GND.n155 13.653
R1989 GND.n149 GND.n148 13.653
R1990 GND.n146 GND.n145 13.653
R1991 GND.n143 GND.n142 13.653
R1992 GND.n135 GND.n134 13.653
R1993 GND.n132 GND.n131 13.653
R1994 GND.n129 GND.n128 13.653
R1995 GND.n126 GND.n125 13.653
R1996 GND.n123 GND.n122 13.653
R1997 GND.n116 GND.n115 13.653
R1998 GND.n113 GND.n112 13.653
R1999 GND.n110 GND.n109 13.653
R2000 GND.n105 GND.n104 13.653
R2001 GND.n102 GND.n101 13.653
R2002 GND.n99 GND.n98 13.653
R2003 GND.n96 GND.n95 13.653
R2004 GND.n93 GND.n92 13.653
R2005 GND.n86 GND.n85 13.653
R2006 GND.n83 GND.n82 13.653
R2007 GND.n80 GND.n79 13.653
R2008 GND.n75 GND.n74 13.653
R2009 GND.n72 GND.n71 13.653
R2010 GND.n8 GND.n7 13.653
R2011 GND.n16 GND.n15 13.653
R2012 GND.n23 GND.n22 13.653
R2013 GND.n26 GND.n25 13.653
R2014 GND.n33 GND.n32 13.653
R2015 GND.n36 GND.n35 13.653
R2016 GND.n39 GND.n38 13.653
R2017 GND.n42 GND.n41 13.653
R2018 GND.n45 GND.n44 13.653
R2019 GND.n50 GND.n49 13.653
R2020 GND.n53 GND.n52 13.653
R2021 GND.n56 GND.n55 13.653
R2022 GND.n63 GND.n62 13.653
R2023 GND.n66 GND.n65 13.653
R2024 GND.n69 GND.n68 13.653
R2025 GND.n20 GND.n19 12.837
R2026 GND.n19 GND.n18 7.566
R2027 GND.n31 GND.n30 7.312
R2028 GND.n61 GND.n60 7.312
R2029 GND.n91 GND.n90 7.312
R2030 GND.n401 GND.n400 7.312
R2031 GND.n434 GND.n433 7.312
R2032 GND.n467 GND.n466 7.312
R2033 GND.n497 GND.n496 7.312
R2034 GND.n527 GND.n526 7.312
R2035 GND.n560 GND.n559 7.312
R2036 GND.n602 GND.n601 7.312
R2037 GND.n632 GND.n631 7.312
R2038 GND.n662 GND.n661 7.312
R2039 GND.n692 GND.n691 7.312
R2040 GND.n349 GND.n348 7.312
R2041 GND.n319 GND.n318 7.312
R2042 GND.n277 GND.n276 7.312
R2043 GND.n247 GND.n246 7.312
R2044 GND.n214 GND.n213 7.312
R2045 GND.n184 GND.n183 7.312
R2046 GND.n154 GND.n153 7.312
R2047 GND.n121 GND.n120 7.312
R2048 GND.n11 GND.n10 4.551
R2049 GND.n8 GND.n6 3.935
R2050 GND.n50 GND.n48 3.935
R2051 GND.n80 GND.n78 3.935
R2052 GND.n110 GND.n108 3.935
R2053 GND.n143 GND.n141 3.935
R2054 GND.n173 GND.n171 3.935
R2055 GND.n203 GND.n201 3.935
R2056 GND.n236 GND.n234 3.935
R2057 GND.n266 GND.n264 3.935
R2058 GND.n338 GND.n336 3.935
R2059 GND.n704 GND.n702 3.935
R2060 GND.n671 GND.n669 3.935
R2061 GND.n641 GND.n639 3.935
R2062 GND.n611 GND.n609 3.935
R2063 GND.n539 GND.n537 3.935
R2064 GND.n506 GND.n504 3.935
R2065 GND.n476 GND.n474 3.935
R2066 GND.n446 GND.n444 3.935
R2067 GND.n413 GND.n411 3.935
R2068 GND.n23 GND.n21 3.541
R2069 GND.t1 GND.n11 2.238
R2070 GND.n360 GND.n359 0.596
R2071 GND.n1 GND.n0 0.596
R2072 GND.n13 GND.n12 0.358
R2073 GND.n34 GND.n27 0.29
R2074 GND.n64 GND.n57 0.29
R2075 GND.n94 GND.n87 0.29
R2076 GND.n124 GND.n117 0.29
R2077 GND.n157 GND.n150 0.29
R2078 GND.n187 GND.n180 0.29
R2079 GND.n217 GND.n210 0.29
R2080 GND.n250 GND.n243 0.29
R2081 GND.n280 GND.n273 0.29
R2082 GND.n322 GND.n315 0.29
R2083 GND.n352 GND.n345 0.29
R2084 GND.n694 GND.n687 0.29
R2085 GND.n664 GND.n657 0.29
R2086 GND.n634 GND.n627 0.29
R2087 GND.n604 GND.n597 0.29
R2088 GND.n562 GND.n555 0.29
R2089 GND.n529 GND.n522 0.29
R2090 GND.n499 GND.n492 0.29
R2091 GND.n469 GND.n462 0.29
R2092 GND.n436 GND.n429 0.29
R2093 GND.n403 GND.n396 0.29
R2094 GND.n361 GND 0.207
R2095 GND.n298 GND.n295 0.197
R2096 GND.n582 GND.n579 0.197
R2097 GND.n381 GND.n378 0.197
R2098 GND.n16 GND.n14 0.196
R2099 GND.n308 GND.n307 0.196
R2100 GND.n569 GND.n568 0.196
R2101 GND.n368 GND.n367 0.196
R2102 GND.n46 GND.n43 0.181
R2103 GND.n76 GND.n73 0.181
R2104 GND.n106 GND.n103 0.181
R2105 GND.n136 GND.n133 0.181
R2106 GND.n169 GND.n166 0.181
R2107 GND.n199 GND.n196 0.181
R2108 GND.n229 GND.n226 0.181
R2109 GND.n262 GND.n259 0.181
R2110 GND.n334 GND.n331 0.181
R2111 GND.n711 GND.n708 0.181
R2112 GND.n678 GND.n675 0.181
R2113 GND.n648 GND.n645 0.181
R2114 GND.n618 GND.n615 0.181
R2115 GND.n546 GND.n543 0.181
R2116 GND.n513 GND.n510 0.181
R2117 GND.n483 GND.n480 0.181
R2118 GND.n453 GND.n450 0.181
R2119 GND.n420 GND.n417 0.181
R2120 GND.n17 GND.n9 0.157
R2121 GND.n24 GND.n17 0.157
R2122 GND.n27 GND.n24 0.145
R2123 GND.n37 GND.n34 0.145
R2124 GND.n40 GND.n37 0.145
R2125 GND.n43 GND.n40 0.145
R2126 GND.n51 GND.n46 0.145
R2127 GND.n54 GND.n51 0.145
R2128 GND.n57 GND.n54 0.145
R2129 GND.n67 GND.n64 0.145
R2130 GND.n70 GND.n67 0.145
R2131 GND.n73 GND.n70 0.145
R2132 GND.n81 GND.n76 0.145
R2133 GND.n84 GND.n81 0.145
R2134 GND.n87 GND.n84 0.145
R2135 GND.n97 GND.n94 0.145
R2136 GND.n100 GND.n97 0.145
R2137 GND.n103 GND.n100 0.145
R2138 GND.n111 GND.n106 0.145
R2139 GND.n114 GND.n111 0.145
R2140 GND.n117 GND.n114 0.145
R2141 GND.n127 GND.n124 0.145
R2142 GND.n130 GND.n127 0.145
R2143 GND.n133 GND.n130 0.145
R2144 GND.n144 GND.n136 0.145
R2145 GND.n147 GND.n144 0.145
R2146 GND.n150 GND.n147 0.145
R2147 GND.n160 GND.n157 0.145
R2148 GND.n163 GND.n160 0.145
R2149 GND.n166 GND.n163 0.145
R2150 GND.n174 GND.n169 0.145
R2151 GND.n177 GND.n174 0.145
R2152 GND.n180 GND.n177 0.145
R2153 GND.n190 GND.n187 0.145
R2154 GND.n193 GND.n190 0.145
R2155 GND.n196 GND.n193 0.145
R2156 GND.n204 GND.n199 0.145
R2157 GND.n207 GND.n204 0.145
R2158 GND.n210 GND.n207 0.145
R2159 GND.n220 GND.n217 0.145
R2160 GND.n223 GND.n220 0.145
R2161 GND.n226 GND.n223 0.145
R2162 GND.n237 GND.n229 0.145
R2163 GND.n240 GND.n237 0.145
R2164 GND.n243 GND.n240 0.145
R2165 GND.n253 GND.n250 0.145
R2166 GND.n256 GND.n253 0.145
R2167 GND.n259 GND.n256 0.145
R2168 GND.n267 GND.n262 0.145
R2169 GND.n270 GND.n267 0.145
R2170 GND.n273 GND.n270 0.145
R2171 GND.n283 GND.n280 0.145
R2172 GND.n286 GND.n283 0.145
R2173 GND.n289 GND.n286 0.145
R2174 GND.n292 GND.n289 0.145
R2175 GND.n295 GND.n292 0.145
R2176 GND.n301 GND.n298 0.145
R2177 GND.n304 GND.n301 0.145
R2178 GND.n309 GND.n304 0.145
R2179 GND.n312 GND.n309 0.145
R2180 GND.n315 GND.n312 0.145
R2181 GND.n325 GND.n322 0.145
R2182 GND.n328 GND.n325 0.145
R2183 GND.n331 GND.n328 0.145
R2184 GND.n339 GND.n334 0.145
R2185 GND.n342 GND.n339 0.145
R2186 GND.n345 GND.n342 0.145
R2187 GND.n355 GND.n352 0.145
R2188 GND.n358 GND.n355 0.145
R2189 GND.n708 GND.n705 0.145
R2190 GND.n705 GND.n697 0.145
R2191 GND.n697 GND.n694 0.145
R2192 GND.n687 GND.n684 0.145
R2193 GND.n684 GND.n681 0.145
R2194 GND.n681 GND.n678 0.145
R2195 GND.n675 GND.n672 0.145
R2196 GND.n672 GND.n667 0.145
R2197 GND.n667 GND.n664 0.145
R2198 GND.n657 GND.n654 0.145
R2199 GND.n654 GND.n651 0.145
R2200 GND.n651 GND.n648 0.145
R2201 GND.n645 GND.n642 0.145
R2202 GND.n642 GND.n637 0.145
R2203 GND.n637 GND.n634 0.145
R2204 GND.n627 GND.n624 0.145
R2205 GND.n624 GND.n621 0.145
R2206 GND.n621 GND.n618 0.145
R2207 GND.n615 GND.n612 0.145
R2208 GND.n612 GND.n607 0.145
R2209 GND.n607 GND.n604 0.145
R2210 GND.n597 GND.n594 0.145
R2211 GND.n594 GND.n591 0.145
R2212 GND.n591 GND.n588 0.145
R2213 GND.n588 GND.n585 0.145
R2214 GND.n585 GND.n582 0.145
R2215 GND.n579 GND.n576 0.145
R2216 GND.n576 GND.n573 0.145
R2217 GND.n573 GND.n570 0.145
R2218 GND.n570 GND.n565 0.145
R2219 GND.n565 GND.n562 0.145
R2220 GND.n555 GND.n552 0.145
R2221 GND.n552 GND.n549 0.145
R2222 GND.n549 GND.n546 0.145
R2223 GND.n543 GND.n540 0.145
R2224 GND.n540 GND.n532 0.145
R2225 GND.n532 GND.n529 0.145
R2226 GND.n522 GND.n519 0.145
R2227 GND.n519 GND.n516 0.145
R2228 GND.n516 GND.n513 0.145
R2229 GND.n510 GND.n507 0.145
R2230 GND.n507 GND.n502 0.145
R2231 GND.n502 GND.n499 0.145
R2232 GND.n492 GND.n489 0.145
R2233 GND.n489 GND.n486 0.145
R2234 GND.n486 GND.n483 0.145
R2235 GND.n480 GND.n477 0.145
R2236 GND.n477 GND.n472 0.145
R2237 GND.n472 GND.n469 0.145
R2238 GND.n462 GND.n459 0.145
R2239 GND.n459 GND.n456 0.145
R2240 GND.n456 GND.n453 0.145
R2241 GND.n450 GND.n447 0.145
R2242 GND.n447 GND.n439 0.145
R2243 GND.n439 GND.n436 0.145
R2244 GND.n429 GND.n426 0.145
R2245 GND.n426 GND.n423 0.145
R2246 GND.n423 GND.n420 0.145
R2247 GND.n417 GND.n414 0.145
R2248 GND.n414 GND.n406 0.145
R2249 GND.n406 GND.n403 0.145
R2250 GND.n396 GND.n393 0.145
R2251 GND.n393 GND.n390 0.145
R2252 GND.n390 GND.n387 0.145
R2253 GND.n387 GND.n384 0.145
R2254 GND.n384 GND.n381 0.145
R2255 GND.n378 GND.n375 0.145
R2256 GND.n375 GND.n372 0.145
R2257 GND.n372 GND.n369 0.145
R2258 GND.n369 GND.n364 0.145
R2259 GND.n364 GND.n361 0.145
R2260 GND GND.n358 0.086
R2261 GND GND.n711 0.058
R2262 a_10429_1050.n3 a_10429_1050.t5 480.392
R2263 a_10429_1050.n3 a_10429_1050.t7 403.272
R2264 a_10429_1050.n4 a_10429_1050.t6 283.48
R2265 a_10429_1050.n7 a_10429_1050.n5 217.114
R2266 a_10429_1050.n5 a_10429_1050.n4 153.315
R2267 a_10429_1050.n5 a_10429_1050.n2 152.499
R2268 a_10429_1050.n4 a_10429_1050.n3 98.447
R2269 a_10429_1050.n2 a_10429_1050.n1 76.002
R2270 a_10429_1050.n7 a_10429_1050.n6 15.218
R2271 a_10429_1050.n0 a_10429_1050.t3 14.282
R2272 a_10429_1050.n0 a_10429_1050.t0 14.282
R2273 a_10429_1050.n1 a_10429_1050.t2 14.282
R2274 a_10429_1050.n1 a_10429_1050.t1 14.282
R2275 a_10429_1050.n2 a_10429_1050.n0 12.85
R2276 a_10429_1050.n8 a_10429_1050.n7 12.014
R2277 a_8731_187.n5 a_8731_187.t8 512.525
R2278 a_8731_187.n3 a_8731_187.t11 472.359
R2279 a_8731_187.n1 a_8731_187.t13 472.359
R2280 a_8731_187.n3 a_8731_187.t5 384.527
R2281 a_8731_187.n1 a_8731_187.t10 384.527
R2282 a_8731_187.n5 a_8731_187.t12 371.139
R2283 a_8731_187.n6 a_8731_187.t7 340.774
R2284 a_8731_187.n4 a_8731_187.t6 294.278
R2285 a_8731_187.n2 a_8731_187.t9 294.278
R2286 a_8731_187.n10 a_8731_187.n9 285.437
R2287 a_8731_187.n6 a_8731_187.n5 109.607
R2288 a_8731_187.n11 a_8731_187.n10 99.394
R2289 a_8731_187.n7 a_8731_187.n6 82.484
R2290 a_8731_187.n8 a_8731_187.n2 80.307
R2291 a_8731_187.n12 a_8731_187.n11 76.001
R2292 a_8731_187.n7 a_8731_187.n4 76
R2293 a_8731_187.n10 a_8731_187.n8 76
R2294 a_8731_187.n4 a_8731_187.n3 56.954
R2295 a_8731_187.n2 a_8731_187.n1 56.954
R2296 a_8731_187.n0 a_8731_187.t2 14.282
R2297 a_8731_187.n0 a_8731_187.t1 14.282
R2298 a_8731_187.t4 a_8731_187.n12 14.282
R2299 a_8731_187.n12 a_8731_187.t3 14.282
R2300 a_8731_187.n11 a_8731_187.n0 12.85
R2301 a_8731_187.n8 a_8731_187.n7 2.947
R2302 a_7595_411.n4 a_7595_411.t8 475.572
R2303 a_7595_411.n8 a_7595_411.t11 472.359
R2304 a_7595_411.n3 a_7595_411.t10 469.145
R2305 a_7595_411.n8 a_7595_411.t7 384.527
R2306 a_7595_411.n4 a_7595_411.t5 384.527
R2307 a_7595_411.n3 a_7595_411.t13 384.527
R2308 a_7595_411.n5 a_7595_411.t9 294.278
R2309 a_7595_411.n11 a_7595_411.n2 232.158
R2310 a_7595_411.n9 a_7595_411.n8 189.719
R2311 a_7595_411.n9 a_7595_411.t6 161.513
R2312 a_7595_411.n7 a_7595_411.t12 161.513
R2313 a_7595_411.n6 a_7595_411.n5 156.851
R2314 a_7595_411.n13 a_7595_411.n11 137.455
R2315 a_7595_411.n7 a_7595_411.n6 132.764
R2316 a_7595_411.n10 a_7595_411.n7 93.638
R2317 a_7595_411.n10 a_7595_411.n9 78.947
R2318 a_7595_411.n2 a_7595_411.n1 76.002
R2319 a_7595_411.n11 a_7595_411.n10 76
R2320 a_7595_411.n5 a_7595_411.n4 57.842
R2321 a_7595_411.n6 a_7595_411.n3 56.833
R2322 a_7595_411.n13 a_7595_411.n12 15.218
R2323 a_7595_411.n0 a_7595_411.t1 14.282
R2324 a_7595_411.n0 a_7595_411.t3 14.282
R2325 a_7595_411.n1 a_7595_411.t2 14.282
R2326 a_7595_411.n1 a_7595_411.t4 14.282
R2327 a_7595_411.n2 a_7595_411.n0 12.85
R2328 a_7595_411.n14 a_7595_411.n13 12.014
R2329 a_13757_1051.n4 a_13757_1051.n3 196.002
R2330 a_13757_1051.n2 a_13757_1051.t4 89.553
R2331 a_13757_1051.n4 a_13757_1051.n0 75.271
R2332 a_13757_1051.n3 a_13757_1051.n2 75.214
R2333 a_13757_1051.n5 a_13757_1051.n4 36.519
R2334 a_13757_1051.n3 a_13757_1051.t3 14.338
R2335 a_13757_1051.n1 a_13757_1051.t5 14.282
R2336 a_13757_1051.n1 a_13757_1051.t2 14.282
R2337 a_13757_1051.n0 a_13757_1051.t6 14.282
R2338 a_13757_1051.n0 a_13757_1051.t7 14.282
R2339 a_13757_1051.t0 a_13757_1051.n5 14.282
R2340 a_13757_1051.n5 a_13757_1051.t1 14.282
R2341 a_13757_1051.n2 a_13757_1051.n1 12.119
R2342 a_13268_209.n1 a_13268_209.t7 512.525
R2343 a_13268_209.n1 a_13268_209.t8 371.139
R2344 a_13268_209.n2 a_13268_209.t9 263.54
R2345 a_13268_209.n14 a_13268_209.n13 216.728
R2346 a_13268_209.n14 a_13268_209.n2 153.043
R2347 a_13268_209.n15 a_13268_209.n14 126.664
R2348 a_13268_209.n2 a_13268_209.n1 120.094
R2349 a_13268_209.n11 a_13268_209.n10 98.501
R2350 a_13268_209.n11 a_13268_209.n6 96.417
R2351 a_13268_209.n13 a_13268_209.n11 78.403
R2352 a_13268_209.n16 a_13268_209.n15 75.27
R2353 a_13268_209.n13 a_13268_209.n12 42.274
R2354 a_13268_209.n6 a_13268_209.n5 30
R2355 a_13268_209.n10 a_13268_209.n9 30
R2356 a_13268_209.n4 a_13268_209.n3 24.383
R2357 a_13268_209.n8 a_13268_209.n7 24.383
R2358 a_13268_209.n6 a_13268_209.n4 23.684
R2359 a_13268_209.n10 a_13268_209.n8 23.684
R2360 a_13268_209.n0 a_13268_209.t4 14.282
R2361 a_13268_209.n0 a_13268_209.t5 14.282
R2362 a_13268_209.t1 a_13268_209.n16 14.282
R2363 a_13268_209.n16 a_13268_209.t0 14.282
R2364 a_13268_209.n15 a_13268_209.n0 12.119
R2365 a_147_187.n7 a_147_187.t7 512.525
R2366 a_147_187.n5 a_147_187.t6 472.359
R2367 a_147_187.n3 a_147_187.t9 472.359
R2368 a_147_187.n5 a_147_187.t10 384.527
R2369 a_147_187.n3 a_147_187.t11 384.527
R2370 a_147_187.n7 a_147_187.t12 371.139
R2371 a_147_187.n8 a_147_187.t8 340.774
R2372 a_147_187.n6 a_147_187.t13 294.278
R2373 a_147_187.n4 a_147_187.t5 294.278
R2374 a_147_187.n13 a_147_187.n11 270.22
R2375 a_147_187.n8 a_147_187.n7 109.607
R2376 a_147_187.n11 a_147_187.n2 99.394
R2377 a_147_187.n9 a_147_187.n8 82.484
R2378 a_147_187.n10 a_147_187.n4 80.307
R2379 a_147_187.n2 a_147_187.n1 76.002
R2380 a_147_187.n9 a_147_187.n6 76
R2381 a_147_187.n11 a_147_187.n10 76
R2382 a_147_187.n6 a_147_187.n5 56.954
R2383 a_147_187.n4 a_147_187.n3 56.954
R2384 a_147_187.n13 a_147_187.n12 15.218
R2385 a_147_187.n0 a_147_187.t2 14.282
R2386 a_147_187.n0 a_147_187.t3 14.282
R2387 a_147_187.n1 a_147_187.t4 14.282
R2388 a_147_187.n1 a_147_187.t1 14.282
R2389 a_147_187.n2 a_147_187.n0 12.85
R2390 a_147_187.n14 a_147_187.n13 12.014
R2391 a_147_187.n10 a_147_187.n9 2.947
R2392 a_3738_101.n12 a_3738_101.n11 26.811
R2393 a_3738_101.n6 a_3738_101.n5 24.977
R2394 a_3738_101.n2 a_3738_101.n1 24.877
R2395 a_3738_101.t0 a_3738_101.n2 12.677
R2396 a_3738_101.t0 a_3738_101.n3 11.595
R2397 a_3738_101.t1 a_3738_101.n8 8.137
R2398 a_3738_101.t0 a_3738_101.n4 7.273
R2399 a_3738_101.t0 a_3738_101.n0 6.109
R2400 a_3738_101.t1 a_3738_101.n7 4.864
R2401 a_3738_101.t0 a_3738_101.n12 2.074
R2402 a_3738_101.n7 a_3738_101.n6 1.13
R2403 a_3738_101.n12 a_3738_101.t1 0.937
R2404 a_3738_101.t1 a_3738_101.n10 0.804
R2405 a_3738_101.n10 a_3738_101.n9 0.136
R2406 a_7364_101.t0 a_7364_101.n1 34.62
R2407 a_7364_101.t0 a_7364_101.n0 8.137
R2408 a_7364_101.t0 a_7364_101.n2 4.69
R2409 a_7469_1050.n0 a_7469_1050.t6 480.392
R2410 a_7469_1050.n0 a_7469_1050.t7 403.272
R2411 a_7469_1050.n1 a_7469_1050.t5 310.033
R2412 a_7469_1050.n3 a_7469_1050.n2 258.884
R2413 a_7469_1050.n3 a_7469_1050.n1 153.315
R2414 a_7469_1050.n5 a_7469_1050.n3 125.947
R2415 a_7469_1050.n5 a_7469_1050.n4 76.002
R2416 a_7469_1050.n1 a_7469_1050.n0 71.894
R2417 a_7469_1050.n4 a_7469_1050.t4 14.282
R2418 a_7469_1050.n4 a_7469_1050.t3 14.282
R2419 a_7469_1050.n6 a_7469_1050.t0 14.282
R2420 a_7469_1050.t1 a_7469_1050.n6 14.282
R2421 a_7469_1050.n6 a_7469_1050.n5 12.848
R2422 Q.n2 Q.n1 253.86
R2423 Q.n2 Q.n0 130.901
R2424 Q.n3 Q.n2 76
R2425 Q.n0 Q.t1 14.282
R2426 Q.n0 Q.t0 14.282
R2427 Q.n3 Q 0.046
R2428 a_10324_101.t0 a_10324_101.n1 34.62
R2429 a_10324_101.t0 a_10324_101.n0 8.137
R2430 a_10324_101.t0 a_10324_101.n2 4.69
R2431 a_9183_989.n0 a_9183_989.t6 480.392
R2432 a_9183_989.n2 a_9183_989.t7 454.685
R2433 a_9183_989.n2 a_9183_989.t5 428.979
R2434 a_9183_989.n0 a_9183_989.t10 403.272
R2435 a_9183_989.n1 a_9183_989.t8 283.48
R2436 a_9183_989.n3 a_9183_989.t9 237.959
R2437 a_9183_989.n9 a_9183_989.n8 210.592
R2438 a_9183_989.n11 a_9183_989.n9 152.499
R2439 a_9183_989.n3 a_9183_989.n2 98.447
R2440 a_9183_989.n1 a_9183_989.n0 98.447
R2441 a_9183_989.n4 a_9183_989.n3 78.947
R2442 a_9183_989.n4 a_9183_989.n1 77.315
R2443 a_9183_989.n11 a_9183_989.n10 76.002
R2444 a_9183_989.n9 a_9183_989.n4 76
R2445 a_9183_989.n8 a_9183_989.n7 30
R2446 a_9183_989.n6 a_9183_989.n5 24.383
R2447 a_9183_989.n8 a_9183_989.n6 23.684
R2448 a_9183_989.n10 a_9183_989.t3 14.282
R2449 a_9183_989.n10 a_9183_989.t4 14.282
R2450 a_9183_989.t1 a_9183_989.n12 14.282
R2451 a_9183_989.n12 a_9183_989.t0 14.282
R2452 a_9183_989.n12 a_9183_989.n11 12.848
R2453 a_8861_1050.n2 a_8861_1050.t7 480.392
R2454 a_8861_1050.n0 a_8861_1050.t12 480.392
R2455 a_8861_1050.n2 a_8861_1050.t10 403.272
R2456 a_8861_1050.n0 a_8861_1050.t11 403.272
R2457 a_8861_1050.n3 a_8861_1050.t8 310.033
R2458 a_8861_1050.n1 a_8861_1050.t9 310.033
R2459 a_8861_1050.n9 a_8861_1050.n8 239.657
R2460 a_8861_1050.n13 a_8861_1050.n9 144.246
R2461 a_8861_1050.n4 a_8861_1050.n1 83.3
R2462 a_8861_1050.n12 a_8861_1050.n11 79.232
R2463 a_8861_1050.n9 a_8861_1050.n4 77.315
R2464 a_8861_1050.n4 a_8861_1050.n3 76
R2465 a_8861_1050.n3 a_8861_1050.n2 71.894
R2466 a_8861_1050.n1 a_8861_1050.n0 71.894
R2467 a_8861_1050.n13 a_8861_1050.n12 63.152
R2468 a_8861_1050.n8 a_8861_1050.n7 30
R2469 a_8861_1050.n6 a_8861_1050.n5 24.383
R2470 a_8861_1050.n8 a_8861_1050.n6 23.684
R2471 a_8861_1050.n12 a_8861_1050.n10 16.08
R2472 a_8861_1050.n14 a_8861_1050.n13 16.078
R2473 a_8861_1050.n10 a_8861_1050.t0 14.282
R2474 a_8861_1050.n10 a_8861_1050.t6 14.282
R2475 a_8861_1050.n11 a_8861_1050.t5 14.282
R2476 a_8861_1050.n11 a_8861_1050.t4 14.282
R2477 a_8861_1050.t2 a_8861_1050.n14 14.282
R2478 a_8861_1050.n14 a_8861_1050.t1 14.282
R2479 CLK.n15 CLK.t5 472.359
R2480 CLK.n6 CLK.t6 472.359
R2481 CLK.n0 CLK.t16 472.359
R2482 CLK.n20 CLK.t2 459.505
R2483 CLK.n11 CLK.t12 459.505
R2484 CLK.n2 CLK.t17 459.505
R2485 CLK.n20 CLK.t13 384.527
R2486 CLK.n15 CLK.t15 384.527
R2487 CLK.n11 CLK.t0 384.527
R2488 CLK.n6 CLK.t7 384.527
R2489 CLK.n2 CLK.t1 384.527
R2490 CLK.n0 CLK.t9 384.527
R2491 CLK.n21 CLK.t8 322.152
R2492 CLK.n12 CLK.t11 322.151
R2493 CLK.n3 CLK.t4 322.151
R2494 CLK.n1 CLK.t14 321.724
R2495 CLK.n17 CLK.t10 319.581
R2496 CLK.n8 CLK.t3 319.581
R2497 CLK.n9 CLK.n8 75.621
R2498 CLK.n18 CLK.n17 75.621
R2499 CLK.n22 CLK.n21 49.342
R2500 CLK.n4 CLK.n3 49.342
R2501 CLK.n13 CLK.n12 49.342
R2502 CLK.n4 CLK.n1 44.933
R2503 CLK.n21 CLK.n20 27.599
R2504 CLK.n3 CLK.n2 27.599
R2505 CLK.n12 CLK.n11 27.599
R2506 CLK.n1 CLK.n0 23.329
R2507 CLK.n16 CLK.n15 21.176
R2508 CLK.n7 CLK.n6 21.176
R2509 CLK.n13 CLK.n10 8.078
R2510 CLK.n22 CLK.n19 8.078
R2511 CLK.n14 CLK.n13 7.797
R2512 CLK.n5 CLK.n4 7.564
R2513 CLK.n17 CLK.n16 4.419
R2514 CLK.n8 CLK.n7 4.419
R2515 CLK.n22 CLK 0.046
R2516 CLK.n10 CLK.n9 0.038
R2517 CLK.n19 CLK.n18 0.038
R2518 CLK.n9 CLK.n5 0.008
R2519 CLK.n18 CLK.n14 0.008
R2520 a_4569_1050.n3 a_4569_1050.t7 480.392
R2521 a_4569_1050.n1 a_4569_1050.t8 480.392
R2522 a_4569_1050.n3 a_4569_1050.t11 403.272
R2523 a_4569_1050.n1 a_4569_1050.t12 403.272
R2524 a_4569_1050.n4 a_4569_1050.t9 310.033
R2525 a_4569_1050.n2 a_4569_1050.t10 310.033
R2526 a_4569_1050.n7 a_4569_1050.n6 261.396
R2527 a_4569_1050.n8 a_4569_1050.n7 144.246
R2528 a_4569_1050.n5 a_4569_1050.n2 83.3
R2529 a_4569_1050.n10 a_4569_1050.n9 79.232
R2530 a_4569_1050.n7 a_4569_1050.n5 77.315
R2531 a_4569_1050.n5 a_4569_1050.n4 76
R2532 a_4569_1050.n4 a_4569_1050.n3 71.894
R2533 a_4569_1050.n2 a_4569_1050.n1 71.894
R2534 a_4569_1050.n10 a_4569_1050.n8 63.152
R2535 a_4569_1050.n8 a_4569_1050.n0 16.08
R2536 a_4569_1050.n11 a_4569_1050.n10 16.078
R2537 a_4569_1050.n0 a_4569_1050.t2 14.282
R2538 a_4569_1050.n0 a_4569_1050.t6 14.282
R2539 a_4569_1050.n9 a_4569_1050.t3 14.282
R2540 a_4569_1050.n9 a_4569_1050.t4 14.282
R2541 a_4569_1050.n11 a_4569_1050.t0 14.282
R2542 a_4569_1050.t1 a_4569_1050.n11 14.282
R2543 a_4439_187.n4 a_4439_187.t10 512.525
R2544 a_4439_187.n2 a_4439_187.t5 472.359
R2545 a_4439_187.n0 a_4439_187.t6 472.359
R2546 a_4439_187.n2 a_4439_187.t11 384.527
R2547 a_4439_187.n0 a_4439_187.t12 384.527
R2548 a_4439_187.n4 a_4439_187.t13 371.139
R2549 a_4439_187.n5 a_4439_187.t8 340.774
R2550 a_4439_187.n3 a_4439_187.t7 294.278
R2551 a_4439_187.n1 a_4439_187.t9 294.278
R2552 a_4439_187.n12 a_4439_187.n11 263.698
R2553 a_4439_187.n5 a_4439_187.n4 109.607
R2554 a_4439_187.n14 a_4439_187.n12 99.394
R2555 a_4439_187.n6 a_4439_187.n5 82.484
R2556 a_4439_187.n7 a_4439_187.n1 80.307
R2557 a_4439_187.n14 a_4439_187.n13 76.002
R2558 a_4439_187.n6 a_4439_187.n3 76
R2559 a_4439_187.n12 a_4439_187.n7 76
R2560 a_4439_187.n3 a_4439_187.n2 56.954
R2561 a_4439_187.n1 a_4439_187.n0 56.954
R2562 a_4439_187.n11 a_4439_187.n10 30
R2563 a_4439_187.n9 a_4439_187.n8 24.383
R2564 a_4439_187.n11 a_4439_187.n9 23.684
R2565 a_4439_187.n13 a_4439_187.t4 14.282
R2566 a_4439_187.n13 a_4439_187.t0 14.282
R2567 a_4439_187.t2 a_4439_187.n15 14.282
R2568 a_4439_187.n15 a_4439_187.t1 14.282
R2569 a_4439_187.n15 a_4439_187.n14 12.848
R2570 a_4439_187.n7 a_4439_187.n6 2.947
R2571 a_6137_1050.n0 a_6137_1050.t5 480.392
R2572 a_6137_1050.n0 a_6137_1050.t6 403.272
R2573 a_6137_1050.n1 a_6137_1050.t7 283.48
R2574 a_6137_1050.n6 a_6137_1050.n5 210.592
R2575 a_6137_1050.n6 a_6137_1050.n1 153.315
R2576 a_6137_1050.n8 a_6137_1050.n6 152.499
R2577 a_6137_1050.n1 a_6137_1050.n0 98.447
R2578 a_6137_1050.n8 a_6137_1050.n7 76.002
R2579 a_6137_1050.n5 a_6137_1050.n4 30
R2580 a_6137_1050.n3 a_6137_1050.n2 24.383
R2581 a_6137_1050.n5 a_6137_1050.n3 23.684
R2582 a_6137_1050.n7 a_6137_1050.t0 14.282
R2583 a_6137_1050.n7 a_6137_1050.t1 14.282
R2584 a_6137_1050.t3 a_6137_1050.n9 14.282
R2585 a_6137_1050.n9 a_6137_1050.t2 14.282
R2586 a_6137_1050.n9 a_6137_1050.n8 12.848
R2587 a_1845_1050.n0 a_1845_1050.t6 480.392
R2588 a_1845_1050.n0 a_1845_1050.t7 403.272
R2589 a_1845_1050.n1 a_1845_1050.t5 283.48
R2590 a_1845_1050.n6 a_1845_1050.n5 210.592
R2591 a_1845_1050.n6 a_1845_1050.n1 153.315
R2592 a_1845_1050.n8 a_1845_1050.n6 152.499
R2593 a_1845_1050.n1 a_1845_1050.n0 98.447
R2594 a_1845_1050.n8 a_1845_1050.n7 76.002
R2595 a_1845_1050.n5 a_1845_1050.n4 30
R2596 a_1845_1050.n3 a_1845_1050.n2 24.383
R2597 a_1845_1050.n5 a_1845_1050.n3 23.684
R2598 a_1845_1050.n7 a_1845_1050.t3 14.282
R2599 a_1845_1050.n7 a_1845_1050.t4 14.282
R2600 a_1845_1050.t1 a_1845_1050.n9 14.282
R2601 a_1845_1050.n9 a_1845_1050.t0 14.282
R2602 a_1845_1050.n9 a_1845_1050.n8 12.848
R2603 a_8675_103.n1 a_8675_103.n0 25.576
R2604 a_8675_103.n3 a_8675_103.n2 9.111
R2605 a_8675_103.n7 a_8675_103.n5 7.859
R2606 a_8675_103.t0 a_8675_103.n7 3.034
R2607 a_8675_103.n5 a_8675_103.n3 1.964
R2608 a_8675_103.n5 a_8675_103.n4 1.964
R2609 a_8675_103.t0 a_8675_103.n1 1.871
R2610 a_8675_103.n7 a_8675_103.n6 0.443
R2611 a_11887_411.n2 a_11887_411.t12 512.525
R2612 a_11887_411.n0 a_11887_411.t6 477.179
R2613 a_11887_411.n5 a_11887_411.t7 472.359
R2614 a_11887_411.n0 a_11887_411.t11 406.485
R2615 a_11887_411.n5 a_11887_411.t9 384.527
R2616 a_11887_411.n2 a_11887_411.t5 371.139
R2617 a_11887_411.n1 a_11887_411.t8 363.924
R2618 a_11887_411.n4 a_11887_411.t10 303.606
R2619 a_11887_411.n6 a_11887_411.t13 267.725
R2620 a_11887_411.n12 a_11887_411.n11 237.145
R2621 a_11887_411.n14 a_11887_411.n12 125.947
R2622 a_11887_411.n3 a_11887_411.n1 101.359
R2623 a_11887_411.n6 a_11887_411.n5 83.507
R2624 a_11887_411.n7 a_11887_411.n6 78.947
R2625 a_11887_411.n7 a_11887_411.n4 77.043
R2626 a_11887_411.n14 a_11887_411.n13 76.002
R2627 a_11887_411.n12 a_11887_411.n7 76
R2628 a_11887_411.n3 a_11887_411.n2 71.88
R2629 a_11887_411.n4 a_11887_411.n3 53.891
R2630 a_11887_411.n11 a_11887_411.n10 30
R2631 a_11887_411.n9 a_11887_411.n8 24.383
R2632 a_11887_411.n11 a_11887_411.n9 23.684
R2633 a_11887_411.n1 a_11887_411.n0 15.776
R2634 a_11887_411.n13 a_11887_411.t0 14.282
R2635 a_11887_411.n13 a_11887_411.t4 14.282
R2636 a_11887_411.n15 a_11887_411.t1 14.282
R2637 a_11887_411.t2 a_11887_411.n15 14.282
R2638 a_11887_411.n15 a_11887_411.n14 12.848
R2639 a_13093_1051.n4 a_13093_1051.n3 195.987
R2640 a_13093_1051.n2 a_13093_1051.t5 89.553
R2641 a_13093_1051.n5 a_13093_1051.n4 75.27
R2642 a_13093_1051.n3 a_13093_1051.n2 75.214
R2643 a_13093_1051.n4 a_13093_1051.n0 36.519
R2644 a_13093_1051.n3 a_13093_1051.t2 14.338
R2645 a_13093_1051.n0 a_13093_1051.t7 14.282
R2646 a_13093_1051.n0 a_13093_1051.t6 14.282
R2647 a_13093_1051.n1 a_13093_1051.t4 14.282
R2648 a_13093_1051.n1 a_13093_1051.t3 14.282
R2649 a_13093_1051.n5 a_13093_1051.t0 14.282
R2650 a_13093_1051.t1 a_13093_1051.n5 14.282
R2651 a_13093_1051.n2 a_13093_1051.n1 12.119
R2652 a_4891_989.n0 a_4891_989.t9 480.392
R2653 a_4891_989.n2 a_4891_989.t7 454.685
R2654 a_4891_989.n2 a_4891_989.t8 428.979
R2655 a_4891_989.n0 a_4891_989.t5 403.272
R2656 a_4891_989.n1 a_4891_989.t10 283.48
R2657 a_4891_989.n3 a_4891_989.t6 237.959
R2658 a_4891_989.n9 a_4891_989.n8 210.592
R2659 a_4891_989.n11 a_4891_989.n9 152.499
R2660 a_4891_989.n3 a_4891_989.n2 98.447
R2661 a_4891_989.n1 a_4891_989.n0 98.447
R2662 a_4891_989.n4 a_4891_989.n3 78.947
R2663 a_4891_989.n4 a_4891_989.n1 77.315
R2664 a_4891_989.n11 a_4891_989.n10 76.002
R2665 a_4891_989.n9 a_4891_989.n4 76
R2666 a_4891_989.n8 a_4891_989.n7 30
R2667 a_4891_989.n6 a_4891_989.n5 24.383
R2668 a_4891_989.n8 a_4891_989.n6 23.684
R2669 a_4891_989.n10 a_4891_989.t4 14.282
R2670 a_4891_989.n10 a_4891_989.t3 14.282
R2671 a_4891_989.t2 a_4891_989.n12 14.282
R2672 a_4891_989.n12 a_4891_989.t1 14.282
R2673 a_4891_989.n12 a_4891_989.n11 12.848
R2674 a_8030_101.n12 a_8030_101.n11 26.811
R2675 a_8030_101.n6 a_8030_101.n5 24.977
R2676 a_8030_101.n2 a_8030_101.n1 24.877
R2677 a_8030_101.t0 a_8030_101.n2 12.677
R2678 a_8030_101.t0 a_8030_101.n3 11.595
R2679 a_8030_101.t1 a_8030_101.n8 8.137
R2680 a_8030_101.t0 a_8030_101.n4 7.273
R2681 a_8030_101.t0 a_8030_101.n0 6.109
R2682 a_8030_101.t1 a_8030_101.n7 4.864
R2683 a_8030_101.t0 a_8030_101.n12 2.074
R2684 a_8030_101.n7 a_8030_101.n6 1.13
R2685 a_8030_101.n12 a_8030_101.t1 0.937
R2686 a_8030_101.t1 a_8030_101.n10 0.804
R2687 a_8030_101.n10 a_8030_101.n9 0.136
R2688 a_1074_101.t0 a_1074_101.n1 34.62
R2689 a_1074_101.t0 a_1074_101.n0 8.137
R2690 a_1074_101.t0 a_1074_101.n2 4.69
R2691 a_277_1050.n3 a_277_1050.t8 480.392
R2692 a_277_1050.n1 a_277_1050.t10 480.392
R2693 a_277_1050.n3 a_277_1050.t11 403.272
R2694 a_277_1050.n1 a_277_1050.t7 403.272
R2695 a_277_1050.n4 a_277_1050.t9 310.033
R2696 a_277_1050.n2 a_277_1050.t12 310.033
R2697 a_277_1050.n10 a_277_1050.n9 239.657
R2698 a_277_1050.n11 a_277_1050.n10 144.246
R2699 a_277_1050.n5 a_277_1050.n2 83.3
R2700 a_277_1050.n13 a_277_1050.n12 79.232
R2701 a_277_1050.n10 a_277_1050.n5 77.315
R2702 a_277_1050.n5 a_277_1050.n4 76
R2703 a_277_1050.n4 a_277_1050.n3 71.894
R2704 a_277_1050.n2 a_277_1050.n1 71.894
R2705 a_277_1050.n13 a_277_1050.n11 63.152
R2706 a_277_1050.n9 a_277_1050.n8 30
R2707 a_277_1050.n7 a_277_1050.n6 24.383
R2708 a_277_1050.n9 a_277_1050.n7 23.684
R2709 a_277_1050.n11 a_277_1050.n0 16.08
R2710 a_277_1050.n14 a_277_1050.n13 16.078
R2711 a_277_1050.n0 a_277_1050.t5 14.282
R2712 a_277_1050.n0 a_277_1050.t4 14.282
R2713 a_277_1050.n12 a_277_1050.t3 14.282
R2714 a_277_1050.n12 a_277_1050.t2 14.282
R2715 a_277_1050.t1 a_277_1050.n14 14.282
R2716 a_277_1050.n14 a_277_1050.t0 14.282
R2717 a_3177_1050.n0 a_3177_1050.t7 480.392
R2718 a_3177_1050.n0 a_3177_1050.t5 403.272
R2719 a_3177_1050.n1 a_3177_1050.t6 310.033
R2720 a_3177_1050.n6 a_3177_1050.n5 237.145
R2721 a_3177_1050.n6 a_3177_1050.n1 153.315
R2722 a_3177_1050.n8 a_3177_1050.n6 125.947
R2723 a_3177_1050.n8 a_3177_1050.n7 76.002
R2724 a_3177_1050.n1 a_3177_1050.n0 71.894
R2725 a_3177_1050.n5 a_3177_1050.n4 30
R2726 a_3177_1050.n3 a_3177_1050.n2 24.383
R2727 a_3177_1050.n5 a_3177_1050.n3 23.684
R2728 a_3177_1050.n7 a_3177_1050.t3 14.282
R2729 a_3177_1050.n7 a_3177_1050.t4 14.282
R2730 a_3177_1050.n9 a_3177_1050.t0 14.282
R2731 a_3177_1050.t1 a_3177_1050.n9 14.282
R2732 a_3177_1050.n9 a_3177_1050.n8 12.848
R2733 a_12322_101.t0 a_12322_101.n1 34.62
R2734 a_12322_101.t0 a_12322_101.n0 8.137
R2735 a_12322_101.t0 a_12322_101.n2 4.69
R2736 a_2406_101.n12 a_2406_101.n11 26.811
R2737 a_2406_101.n6 a_2406_101.n5 24.977
R2738 a_2406_101.n2 a_2406_101.n1 24.877
R2739 a_2406_101.t0 a_2406_101.n2 12.677
R2740 a_2406_101.t0 a_2406_101.n3 11.595
R2741 a_2406_101.t1 a_2406_101.n8 8.137
R2742 a_2406_101.t0 a_2406_101.n4 7.273
R2743 a_2406_101.t0 a_2406_101.n0 6.109
R2744 a_2406_101.t1 a_2406_101.n7 4.864
R2745 a_2406_101.t0 a_2406_101.n12 2.074
R2746 a_2406_101.n7 a_2406_101.n6 1.13
R2747 a_2406_101.n12 a_2406_101.t1 0.937
R2748 a_2406_101.t1 a_2406_101.n10 0.804
R2749 a_2406_101.n10 a_2406_101.n9 0.136
R2750 a_372_210.n10 a_372_210.n8 82.852
R2751 a_372_210.n7 a_372_210.n6 32.833
R2752 a_372_210.n8 a_372_210.t1 32.416
R2753 a_372_210.n10 a_372_210.n9 27.2
R2754 a_372_210.n11 a_372_210.n0 23.498
R2755 a_372_210.n3 a_372_210.n2 23.284
R2756 a_372_210.n11 a_372_210.n10 22.4
R2757 a_372_210.n7 a_372_210.n4 19.017
R2758 a_372_210.n6 a_372_210.n5 13.494
R2759 a_372_210.t1 a_372_210.n1 7.04
R2760 a_372_210.t1 a_372_210.n3 5.727
R2761 a_372_210.n8 a_372_210.n7 1.435
R2762 a_11761_1050.n0 a_11761_1050.t6 480.392
R2763 a_11761_1050.n0 a_11761_1050.t5 403.272
R2764 a_11761_1050.n1 a_11761_1050.t7 363.924
R2765 a_11761_1050.n6 a_11761_1050.n5 290.251
R2766 a_11761_1050.n6 a_11761_1050.n1 126.657
R2767 a_11761_1050.n8 a_11761_1050.n7 76.002
R2768 a_11761_1050.n8 a_11761_1050.n6 72.841
R2769 a_11761_1050.n5 a_11761_1050.n4 30
R2770 a_11761_1050.n3 a_11761_1050.n2 24.383
R2771 a_11761_1050.n5 a_11761_1050.n3 23.684
R2772 a_11761_1050.n1 a_11761_1050.n0 15.545
R2773 a_11761_1050.n7 a_11761_1050.t3 14.282
R2774 a_11761_1050.n7 a_11761_1050.t4 14.282
R2775 a_11761_1050.t2 a_11761_1050.n9 14.282
R2776 a_11761_1050.n9 a_11761_1050.t1 14.282
R2777 a_11761_1050.n9 a_11761_1050.n8 12.848
R2778 a_9658_101.n12 a_9658_101.n11 26.811
R2779 a_9658_101.n6 a_9658_101.n5 24.977
R2780 a_9658_101.n2 a_9658_101.n1 24.877
R2781 a_9658_101.t0 a_9658_101.n2 12.677
R2782 a_9658_101.t0 a_9658_101.n3 11.595
R2783 a_9658_101.t1 a_9658_101.n8 8.137
R2784 a_9658_101.t0 a_9658_101.n4 7.273
R2785 a_9658_101.t0 a_9658_101.n0 6.109
R2786 a_9658_101.t1 a_9658_101.n7 4.864
R2787 a_9658_101.t0 a_9658_101.n12 2.074
R2788 a_9658_101.n7 a_9658_101.n6 1.13
R2789 a_9658_101.n12 a_9658_101.t1 0.937
R2790 a_9658_101.t1 a_9658_101.n10 0.804
R2791 a_9658_101.n10 a_9658_101.n9 0.136
R2792 a_4664_210.n10 a_4664_210.n8 82.852
R2793 a_4664_210.n7 a_4664_210.n6 32.833
R2794 a_4664_210.n8 a_4664_210.t1 32.416
R2795 a_4664_210.n10 a_4664_210.n9 27.2
R2796 a_4664_210.n11 a_4664_210.n0 23.498
R2797 a_4664_210.n3 a_4664_210.n2 23.284
R2798 a_4664_210.n11 a_4664_210.n10 22.4
R2799 a_4664_210.n7 a_4664_210.n4 19.017
R2800 a_4664_210.n6 a_4664_210.n5 13.494
R2801 a_4664_210.t1 a_4664_210.n1 7.04
R2802 a_4664_210.t1 a_4664_210.n3 5.727
R2803 a_4664_210.n8 a_4664_210.n7 1.435
R2804 a_3072_101.t0 a_3072_101.n1 34.62
R2805 a_3072_101.t0 a_3072_101.n0 8.137
R2806 a_3072_101.t0 a_3072_101.n2 4.69
R2807 a_6698_101.n12 a_6698_101.n11 26.811
R2808 a_6698_101.n6 a_6698_101.n5 24.977
R2809 a_6698_101.n2 a_6698_101.n1 24.877
R2810 a_6698_101.t0 a_6698_101.n2 12.677
R2811 a_6698_101.t0 a_6698_101.n3 11.595
R2812 a_6698_101.t1 a_6698_101.n8 8.137
R2813 a_6698_101.t0 a_6698_101.n4 7.273
R2814 a_6698_101.t0 a_6698_101.n0 6.109
R2815 a_6698_101.t1 a_6698_101.n7 4.864
R2816 a_6698_101.t0 a_6698_101.n12 2.074
R2817 a_6698_101.n7 a_6698_101.n6 1.13
R2818 a_6698_101.n12 a_6698_101.t1 0.937
R2819 a_6698_101.t1 a_6698_101.n10 0.804
R2820 a_6698_101.n10 a_6698_101.n9 0.136
R2821 a_6032_101.t0 a_6032_101.n1 34.62
R2822 a_6032_101.t0 a_6032_101.n0 8.137
R2823 a_6032_101.t0 a_6032_101.n2 4.69
R2824 a_91_103.n1 a_91_103.n0 25.576
R2825 a_91_103.n3 a_91_103.n2 9.111
R2826 a_91_103.n7 a_91_103.n6 2.455
R2827 a_91_103.n5 a_91_103.n3 1.964
R2828 a_91_103.n5 a_91_103.n4 1.964
R2829 a_91_103.t0 a_91_103.n1 1.871
R2830 a_91_103.n7 a_91_103.n5 0.636
R2831 a_91_103.t0 a_91_103.n7 0.246
R2832 a_8956_210.n10 a_8956_210.n8 82.852
R2833 a_8956_210.n11 a_8956_210.n0 49.6
R2834 a_8956_210.n7 a_8956_210.n6 32.833
R2835 a_8956_210.n8 a_8956_210.t1 32.416
R2836 a_8956_210.n10 a_8956_210.n9 27.2
R2837 a_8956_210.n3 a_8956_210.n2 23.284
R2838 a_8956_210.n11 a_8956_210.n10 22.4
R2839 a_8956_210.n7 a_8956_210.n4 19.017
R2840 a_8956_210.n6 a_8956_210.n5 13.494
R2841 a_8956_210.t1 a_8956_210.n1 7.04
R2842 a_8956_210.t1 a_8956_210.n3 5.727
R2843 a_8956_210.n8 a_8956_210.n7 1.435
R2844 a_11656_101.t0 a_11656_101.n1 34.62
R2845 a_11656_101.t0 a_11656_101.n0 8.137
R2846 a_11656_101.t0 a_11656_101.n2 4.69
R2847 a_10990_101.t0 a_10990_101.n1 34.62
R2848 a_10990_101.t0 a_10990_101.n0 8.137
R2849 a_10990_101.t0 a_10990_101.n2 4.69
R2850 a_4383_103.n1 a_4383_103.n0 25.576
R2851 a_4383_103.n3 a_4383_103.n2 9.111
R2852 a_4383_103.n7 a_4383_103.n6 2.455
R2853 a_4383_103.n5 a_4383_103.n3 1.964
R2854 a_4383_103.n5 a_4383_103.n4 1.964
R2855 a_4383_103.t0 a_4383_103.n1 1.871
R2856 a_4383_103.n7 a_4383_103.n5 0.636
R2857 a_4383_103.t0 a_4383_103.n7 0.246
R2858 a_5366_101.t0 a_5366_101.n1 34.62
R2859 a_5366_101.t0 a_5366_101.n0 8.137
R2860 a_5366_101.t0 a_5366_101.n2 4.69
R2861 a_1740_101.t0 a_1740_101.n1 34.62
R2862 a_1740_101.t0 a_1740_101.n0 8.137
R2863 a_1740_101.t0 a_1740_101.n2 4.69
R2864 a_13654_101.t0 a_13654_101.n0 34.602
R2865 a_13654_101.t0 a_13654_101.n1 2.138
R2866 a_12988_101.n13 a_12988_101.n12 26.811
R2867 a_12988_101.n6 a_12988_101.n5 24.977
R2868 a_12988_101.n2 a_12988_101.n1 24.877
R2869 a_12988_101.t0 a_12988_101.n2 12.677
R2870 a_12988_101.t0 a_12988_101.n3 11.595
R2871 a_12988_101.n11 a_12988_101.n10 8.561
R2872 a_12988_101.t0 a_12988_101.n4 7.273
R2873 a_12988_101.n9 a_12988_101.n8 7.066
R2874 a_12988_101.t0 a_12988_101.n0 6.109
R2875 a_12988_101.t1 a_12988_101.n7 4.864
R2876 a_12988_101.t0 a_12988_101.n13 2.074
R2877 a_12988_101.n7 a_12988_101.n6 1.13
R2878 a_12988_101.t1 a_12988_101.n11 0.958
R2879 a_12988_101.n13 a_12988_101.t1 0.937
R2880 a_12988_101.t1 a_12988_101.n9 0.86
C4 VDD GND 56.51fF
C5 a_12988_101.n0 GND 0.02fF
C6 a_12988_101.n1 GND 0.09fF
C7 a_12988_101.n2 GND 0.05fF
C8 a_12988_101.n3 GND 0.06fF
C9 a_12988_101.n4 GND 0.00fF
C10 a_12988_101.n5 GND 0.04fF
C11 a_12988_101.n6 GND 0.05fF
C12 a_12988_101.n7 GND 0.02fF
C13 a_12988_101.n8 GND 0.05fF
C14 a_12988_101.n9 GND 0.09fF
C15 a_12988_101.n10 GND 0.21fF
C16 a_12988_101.n11 GND 0.07fF
C17 a_12988_101.t1 GND 0.14fF
C18 a_12988_101.n12 GND 0.04fF
C19 a_12988_101.n13 GND 0.00fF
C20 a_13654_101.n0 GND 0.13fF
C21 a_13654_101.n1 GND 0.13fF
C22 a_1740_101.n0 GND 0.05fF
C23 a_1740_101.n1 GND 0.12fF
C24 a_1740_101.n2 GND 0.04fF
C25 a_5366_101.n0 GND 0.05fF
C26 a_5366_101.n1 GND 0.12fF
C27 a_5366_101.n2 GND 0.04fF
C28 a_4383_103.n0 GND 0.09fF
C29 a_4383_103.n1 GND 0.10fF
C30 a_4383_103.n2 GND 0.05fF
C31 a_4383_103.n3 GND 0.03fF
C32 a_4383_103.n4 GND 0.04fF
C33 a_4383_103.n5 GND 0.03fF
C34 a_4383_103.n6 GND 0.04fF
C35 a_10990_101.n0 GND 0.05fF
C36 a_10990_101.n1 GND 0.12fF
C37 a_10990_101.n2 GND 0.04fF
C38 a_11656_101.n0 GND 0.05fF
C39 a_11656_101.n1 GND 0.12fF
C40 a_11656_101.n2 GND 0.04fF
C41 a_8956_210.n0 GND 0.02fF
C42 a_8956_210.n1 GND 0.09fF
C43 a_8956_210.n2 GND 0.13fF
C44 a_8956_210.n3 GND 0.11fF
C45 a_8956_210.t1 GND 0.30fF
C46 a_8956_210.n4 GND 0.09fF
C47 a_8956_210.n5 GND 0.06fF
C48 a_8956_210.n6 GND 0.01fF
C49 a_8956_210.n7 GND 0.03fF
C50 a_8956_210.n8 GND 0.11fF
C51 a_8956_210.n9 GND 0.02fF
C52 a_8956_210.n10 GND 0.05fF
C53 a_8956_210.n11 GND 0.02fF
C54 a_91_103.n0 GND 0.09fF
C55 a_91_103.n1 GND 0.09fF
C56 a_91_103.n2 GND 0.04fF
C57 a_91_103.n3 GND 0.03fF
C58 a_91_103.n4 GND 0.04fF
C59 a_91_103.n5 GND 0.03fF
C60 a_91_103.n6 GND 0.04fF
C61 a_6032_101.n0 GND 0.05fF
C62 a_6032_101.n1 GND 0.12fF
C63 a_6032_101.n2 GND 0.04fF
C64 a_6698_101.n0 GND 0.02fF
C65 a_6698_101.n1 GND 0.10fF
C66 a_6698_101.n2 GND 0.06fF
C67 a_6698_101.n3 GND 0.06fF
C68 a_6698_101.n4 GND 0.00fF
C69 a_6698_101.n5 GND 0.04fF
C70 a_6698_101.n6 GND 0.05fF
C71 a_6698_101.n7 GND 0.02fF
C72 a_6698_101.n8 GND 0.05fF
C73 a_6698_101.n9 GND 0.08fF
C74 a_6698_101.n10 GND 0.17fF
C75 a_6698_101.t1 GND 0.23fF
C76 a_6698_101.n11 GND 0.09fF
C77 a_6698_101.n12 GND 0.00fF
C78 a_3072_101.n0 GND 0.05fF
C79 a_3072_101.n1 GND 0.12fF
C80 a_3072_101.n2 GND 0.04fF
C81 a_4664_210.n0 GND 0.02fF
C82 a_4664_210.n1 GND 0.09fF
C83 a_4664_210.n2 GND 0.13fF
C84 a_4664_210.n3 GND 0.11fF
C85 a_4664_210.t1 GND 0.30fF
C86 a_4664_210.n4 GND 0.09fF
C87 a_4664_210.n5 GND 0.06fF
C88 a_4664_210.n6 GND 0.01fF
C89 a_4664_210.n7 GND 0.03fF
C90 a_4664_210.n8 GND 0.11fF
C91 a_4664_210.n9 GND 0.02fF
C92 a_4664_210.n10 GND 0.05fF
C93 a_4664_210.n11 GND 0.03fF
C94 a_9658_101.n0 GND 0.02fF
C95 a_9658_101.n1 GND 0.10fF
C96 a_9658_101.n2 GND 0.06fF
C97 a_9658_101.n3 GND 0.06fF
C98 a_9658_101.n4 GND 0.00fF
C99 a_9658_101.n5 GND 0.04fF
C100 a_9658_101.n6 GND 0.05fF
C101 a_9658_101.n7 GND 0.02fF
C102 a_9658_101.n8 GND 0.05fF
C103 a_9658_101.n9 GND 0.08fF
C104 a_9658_101.n10 GND 0.17fF
C105 a_9658_101.t1 GND 0.23fF
C106 a_9658_101.n11 GND 0.09fF
C107 a_9658_101.n12 GND 0.00fF
C108 a_11761_1050.n0 GND 0.27fF
C109 a_11761_1050.n1 GND 0.62fF
C110 a_11761_1050.n2 GND 0.04fF
C111 a_11761_1050.n3 GND 0.05fF
C112 a_11761_1050.n4 GND 0.03fF
C113 a_11761_1050.n5 GND 0.39fF
C114 a_11761_1050.n6 GND 0.56fF
C115 a_11761_1050.n7 GND 0.62fF
C116 a_11761_1050.n8 GND 0.21fF
C117 a_11761_1050.n9 GND 0.53fF
C118 a_372_210.n0 GND 0.02fF
C119 a_372_210.n1 GND 0.09fF
C120 a_372_210.n2 GND 0.13fF
C121 a_372_210.n3 GND 0.11fF
C122 a_372_210.t1 GND 0.30fF
C123 a_372_210.n4 GND 0.09fF
C124 a_372_210.n5 GND 0.06fF
C125 a_372_210.n6 GND 0.01fF
C126 a_372_210.n7 GND 0.03fF
C127 a_372_210.n8 GND 0.11fF
C128 a_372_210.n9 GND 0.02fF
C129 a_372_210.n10 GND 0.05fF
C130 a_372_210.n11 GND 0.03fF
C131 a_2406_101.n0 GND 0.02fF
C132 a_2406_101.n1 GND 0.10fF
C133 a_2406_101.n2 GND 0.06fF
C134 a_2406_101.n3 GND 0.06fF
C135 a_2406_101.n4 GND 0.00fF
C136 a_2406_101.n5 GND 0.04fF
C137 a_2406_101.n6 GND 0.05fF
C138 a_2406_101.n7 GND 0.02fF
C139 a_2406_101.n8 GND 0.05fF
C140 a_2406_101.n9 GND 0.08fF
C141 a_2406_101.n10 GND 0.17fF
C142 a_2406_101.t1 GND 0.23fF
C143 a_2406_101.n11 GND 0.09fF
C144 a_2406_101.n12 GND 0.00fF
C145 a_12322_101.n0 GND 0.05fF
C146 a_12322_101.n1 GND 0.12fF
C147 a_12322_101.n2 GND 0.04fF
C148 a_3177_1050.n0 GND 0.36fF
C149 a_3177_1050.n1 GND 0.60fF
C150 a_3177_1050.n2 GND 0.04fF
C151 a_3177_1050.n3 GND 0.06fF
C152 a_3177_1050.n4 GND 0.04fF
C153 a_3177_1050.n5 GND 0.34fF
C154 a_3177_1050.n6 GND 0.62fF
C155 a_3177_1050.n7 GND 0.65fF
C156 a_3177_1050.n8 GND 0.29fF
C157 a_3177_1050.n9 GND 0.55fF
C158 a_277_1050.n0 GND 0.72fF
C159 a_277_1050.n1 GND 0.46fF
C160 a_277_1050.n2 GND 0.64fF
C161 a_277_1050.n3 GND 0.46fF
C162 a_277_1050.n4 GND 0.54fF
C163 a_277_1050.n5 GND 2.59fF
C164 a_277_1050.n6 GND 0.05fF
C165 a_277_1050.n7 GND 0.07fF
C166 a_277_1050.n8 GND 0.05fF
C167 a_277_1050.n9 GND 0.45fF
C168 a_277_1050.n10 GND 0.61fF
C169 a_277_1050.n11 GND 0.37fF
C170 a_277_1050.n12 GND 0.85fF
C171 a_277_1050.n13 GND 0.27fF
C172 a_277_1050.n14 GND 0.72fF
C173 a_1074_101.n0 GND 0.05fF
C174 a_1074_101.n1 GND 0.12fF
C175 a_1074_101.n2 GND 0.04fF
C176 a_8030_101.n0 GND 0.02fF
C177 a_8030_101.n1 GND 0.10fF
C178 a_8030_101.n2 GND 0.06fF
C179 a_8030_101.n3 GND 0.06fF
C180 a_8030_101.n4 GND 0.00fF
C181 a_8030_101.n5 GND 0.04fF
C182 a_8030_101.n6 GND 0.05fF
C183 a_8030_101.n7 GND 0.02fF
C184 a_8030_101.n8 GND 0.05fF
C185 a_8030_101.n9 GND 0.08fF
C186 a_8030_101.n10 GND 0.17fF
C187 a_8030_101.t1 GND 0.23fF
C188 a_8030_101.n11 GND 0.09fF
C189 a_8030_101.n12 GND 0.00fF
C190 a_4891_989.n0 GND 0.49fF
C191 a_4891_989.n1 GND 0.52fF
C192 a_4891_989.n2 GND 0.49fF
C193 a_4891_989.t6 GND 0.69fF
C194 a_4891_989.n3 GND 0.50fF
C195 a_4891_989.n4 GND 1.33fF
C196 a_4891_989.n5 GND 0.05fF
C197 a_4891_989.n6 GND 0.07fF
C198 a_4891_989.n7 GND 0.04fF
C199 a_4891_989.n8 GND 0.39fF
C200 a_4891_989.n9 GND 0.56fF
C201 a_4891_989.n10 GND 0.82fF
C202 a_4891_989.n11 GND 0.40fF
C203 a_4891_989.n12 GND 0.69fF
C204 a_13093_1051.n0 GND 0.37fF
C205 a_13093_1051.n1 GND 0.33fF
C206 a_13093_1051.n2 GND 0.24fF
C207 a_13093_1051.n3 GND 0.63fF
C208 a_13093_1051.n4 GND 0.28fF
C209 a_13093_1051.n5 GND 0.41fF
C210 a_11887_411.n0 GND 0.28fF
C211 a_11887_411.n1 GND 0.74fF
C212 a_11887_411.n2 GND 0.25fF
C213 a_11887_411.n3 GND 0.50fF
C214 a_11887_411.n4 GND 0.37fF
C215 a_11887_411.n5 GND 0.31fF
C216 a_11887_411.t13 GND 0.56fF
C217 a_11887_411.n6 GND 0.40fF
C218 a_11887_411.n7 GND 0.96fF
C219 a_11887_411.n8 GND 0.04fF
C220 a_11887_411.n9 GND 0.05fF
C221 a_11887_411.n10 GND 0.03fF
C222 a_11887_411.n11 GND 0.33fF
C223 a_11887_411.n12 GND 0.43fF
C224 a_11887_411.n13 GND 0.63fF
C225 a_11887_411.n14 GND 0.28fF
C226 a_11887_411.n15 GND 0.53fF
C227 a_8675_103.n0 GND 0.09fF
C228 a_8675_103.n1 GND 0.10fF
C229 a_8675_103.n2 GND 0.05fF
C230 a_8675_103.n3 GND 0.03fF
C231 a_8675_103.n4 GND 0.04fF
C232 a_8675_103.n5 GND 0.11fF
C233 a_8675_103.n6 GND 0.04fF
C234 a_1845_1050.n0 GND 0.39fF
C235 a_1845_1050.n1 GND 0.59fF
C236 a_1845_1050.n2 GND 0.04fF
C237 a_1845_1050.n3 GND 0.06fF
C238 a_1845_1050.n4 GND 0.04fF
C239 a_1845_1050.n5 GND 0.31fF
C240 a_1845_1050.n6 GND 0.62fF
C241 a_1845_1050.n7 GND 0.64fF
C242 a_1845_1050.n8 GND 0.31fF
C243 a_1845_1050.n9 GND 0.54fF
C244 a_6137_1050.n0 GND 0.43fF
C245 a_6137_1050.n1 GND 0.65fF
C246 a_6137_1050.n2 GND 0.05fF
C247 a_6137_1050.n3 GND 0.06fF
C248 a_6137_1050.n4 GND 0.04fF
C249 a_6137_1050.n5 GND 0.34fF
C250 a_6137_1050.n6 GND 0.69fF
C251 a_6137_1050.n7 GND 0.71fF
C252 a_6137_1050.n8 GND 0.35fF
C253 a_6137_1050.n9 GND 0.60fF
C254 a_4439_187.n0 GND 0.45fF
C255 a_4439_187.t9 GND 0.96fF
C256 a_4439_187.n1 GND 0.66fF
C257 a_4439_187.n2 GND 0.45fF
C258 a_4439_187.t7 GND 0.96fF
C259 a_4439_187.n3 GND 0.62fF
C260 a_4439_187.n4 GND 0.44fF
C261 a_4439_187.n5 GND 0.88fF
C262 a_4439_187.n6 GND 2.85fF
C263 a_4439_187.n7 GND 2.12fF
C264 a_4439_187.n8 GND 0.07fF
C265 a_4439_187.n9 GND 0.09fF
C266 a_4439_187.n10 GND 0.06fF
C267 a_4439_187.n11 GND 0.58fF
C268 a_4439_187.n12 GND 0.69fF
C269 a_4439_187.n13 GND 1.01fF
C270 a_4439_187.n14 GND 0.40fF
C271 a_4439_187.n15 GND 0.86fF
C272 a_4569_1050.n0 GND 0.79fF
C273 a_4569_1050.n1 GND 0.51fF
C274 a_4569_1050.n2 GND 0.70fF
C275 a_4569_1050.n3 GND 0.51fF
C276 a_4569_1050.n4 GND 0.59fF
C277 a_4569_1050.n5 GND 2.84fF
C278 a_4569_1050.n6 GND 0.64fF
C279 a_4569_1050.n7 GND 0.71fF
C280 a_4569_1050.n8 GND 0.41fF
C281 a_4569_1050.n9 GND 0.93fF
C282 a_4569_1050.n10 GND 0.29fF
C283 a_4569_1050.n11 GND 0.79fF
C284 a_8861_1050.n0 GND 0.51fF
C285 a_8861_1050.n1 GND 0.69fF
C286 a_8861_1050.n2 GND 0.51fF
C287 a_8861_1050.n3 GND 0.59fF
C288 a_8861_1050.n4 GND 2.83fF
C289 a_8861_1050.n5 GND 0.06fF
C290 a_8861_1050.n6 GND 0.08fF
C291 a_8861_1050.n7 GND 0.05fF
C292 a_8861_1050.n8 GND 0.49fF
C293 a_8861_1050.n9 GND 0.67fF
C294 a_8861_1050.n10 GND 0.79fF
C295 a_8861_1050.n11 GND 0.93fF
C296 a_8861_1050.n12 GND 0.29fF
C297 a_8861_1050.n13 GND 0.41fF
C298 a_8861_1050.n14 GND 0.79fF
C299 a_9183_989.n0 GND 0.50fF
C300 a_9183_989.n1 GND 0.53fF
C301 a_9183_989.n2 GND 0.50fF
C302 a_9183_989.t9 GND 0.71fF
C303 a_9183_989.n3 GND 0.51fF
C304 a_9183_989.n4 GND 1.36fF
C305 a_9183_989.n5 GND 0.05fF
C306 a_9183_989.n6 GND 0.07fF
C307 a_9183_989.n7 GND 0.05fF
C308 a_9183_989.n8 GND 0.40fF
C309 a_9183_989.n9 GND 0.57fF
C310 a_9183_989.n10 GND 0.84fF
C311 a_9183_989.n11 GND 0.41fF
C312 a_9183_989.n12 GND 0.71fF
C313 a_10324_101.n0 GND 0.05fF
C314 a_10324_101.n1 GND 0.12fF
C315 a_10324_101.n2 GND 0.04fF
C316 Q.n0 GND 0.75fF
C317 Q.n1 GND 0.45fF
C318 Q.n2 GND 0.51fF
C319 Q.n3 GND 0.01fF
C320 a_7469_1050.n0 GND 0.37fF
C321 a_7469_1050.n1 GND 0.61fF
C322 a_7469_1050.n2 GND 0.46fF
C323 a_7469_1050.n3 GND 0.67fF
C324 a_7469_1050.n4 GND 0.67fF
C325 a_7469_1050.n5 GND 0.29fF
C326 a_7469_1050.n6 GND 0.56fF
C327 a_7364_101.n0 GND 0.05fF
C328 a_7364_101.n1 GND 0.12fF
C329 a_7364_101.n2 GND 0.04fF
C330 a_3738_101.n0 GND 0.02fF
C331 a_3738_101.n1 GND 0.10fF
C332 a_3738_101.n2 GND 0.06fF
C333 a_3738_101.n3 GND 0.06fF
C334 a_3738_101.n4 GND 0.00fF
C335 a_3738_101.n5 GND 0.04fF
C336 a_3738_101.n6 GND 0.05fF
C337 a_3738_101.n7 GND 0.02fF
C338 a_3738_101.n8 GND 0.05fF
C339 a_3738_101.n9 GND 0.08fF
C340 a_3738_101.n10 GND 0.17fF
C341 a_3738_101.t1 GND 0.23fF
C342 a_3738_101.n11 GND 0.09fF
C343 a_3738_101.n12 GND 0.00fF
C344 a_147_187.n0 GND 0.79fF
C345 a_147_187.n1 GND 0.93fF
C346 a_147_187.n2 GND 0.36fF
C347 a_147_187.n3 GND 0.41fF
C348 a_147_187.t5 GND 0.88fF
C349 a_147_187.n4 GND 0.61fF
C350 a_147_187.n5 GND 0.41fF
C351 a_147_187.t13 GND 0.88fF
C352 a_147_187.n6 GND 0.57fF
C353 a_147_187.n7 GND 0.41fF
C354 a_147_187.n8 GND 0.81fF
C355 a_147_187.n9 GND 2.62fF
C356 a_147_187.n10 GND 1.95fF
C357 a_147_187.n11 GND 0.64fF
C358 a_147_187.n12 GND 0.12fF
C359 a_147_187.n13 GND 0.52fF
C360 a_147_187.n14 GND 0.07fF
C361 a_13268_209.n0 GND 0.37fF
C362 a_13268_209.n1 GND 0.26fF
C363 a_13268_209.n2 GND 0.48fF
C364 a_13268_209.n3 GND 0.03fF
C365 a_13268_209.n4 GND 0.04fF
C366 a_13268_209.n5 GND 0.03fF
C367 a_13268_209.n6 GND 0.08fF
C368 a_13268_209.n7 GND 0.03fF
C369 a_13268_209.n8 GND 0.04fF
C370 a_13268_209.n9 GND 0.03fF
C371 a_13268_209.n10 GND 0.09fF
C372 a_13268_209.n11 GND 0.96fF
C373 a_13268_209.n12 GND 0.12fF
C374 a_13268_209.n13 GND 0.29fF
C375 a_13268_209.n14 GND 0.45fF
C376 a_13268_209.n15 GND 0.23fF
C377 a_13268_209.n16 GND 0.45fF
C378 a_13757_1051.n0 GND 0.36fF
C379 a_13757_1051.n1 GND 0.29fF
C380 a_13757_1051.n2 GND 0.20fF
C381 a_13757_1051.n3 GND 0.57fF
C382 a_13757_1051.n4 GND 0.25fF
C383 a_13757_1051.n5 GND 0.28fF
C384 a_7595_411.n0 GND 0.69fF
C385 a_7595_411.n1 GND 0.81fF
C386 a_7595_411.n2 GND 0.52fF
C387 a_7595_411.n3 GND 0.36fF
C388 a_7595_411.n4 GND 0.40fF
C389 a_7595_411.t9 GND 0.76fF
C390 a_7595_411.n5 GND 1.26fF
C391 a_7595_411.n6 GND 1.02fF
C392 a_7595_411.t12 GND 0.59fF
C393 a_7595_411.n7 GND 0.88fF
C394 a_7595_411.n8 GND 0.55fF
C395 a_7595_411.t6 GND 0.59fF
C396 a_7595_411.n9 GND 0.50fF
C397 a_7595_411.n10 GND 5.53fF
C398 a_7595_411.n11 GND 0.57fF
C399 a_7595_411.n12 GND 0.11fF
C400 a_7595_411.n13 GND 0.25fF
C401 a_7595_411.n14 GND 0.06fF
C402 a_8731_187.n0 GND 0.84fF
C403 a_8731_187.n1 GND 0.44fF
C404 a_8731_187.t9 GND 0.94fF
C405 a_8731_187.n2 GND 0.65fF
C406 a_8731_187.n3 GND 0.44fF
C407 a_8731_187.t6 GND 0.94fF
C408 a_8731_187.n4 GND 0.61fF
C409 a_8731_187.n5 GND 0.43fF
C410 a_8731_187.n6 GND 0.86fF
C411 a_8731_187.n7 GND 2.79fF
C412 a_8731_187.n8 GND 2.08fF
C413 a_8731_187.n9 GND 0.73fF
C414 a_8731_187.n10 GND 0.72fF
C415 a_8731_187.n11 GND 0.39fF
C416 a_8731_187.n12 GND 0.99fF
C417 a_10429_1050.n0 GND 0.60fF
C418 a_10429_1050.n1 GND 0.71fF
C419 a_10429_1050.n2 GND 0.35fF
C420 a_10429_1050.n3 GND 0.43fF
C421 a_10429_1050.n4 GND 0.65fF
C422 a_10429_1050.n5 GND 0.69fF
C423 a_10429_1050.n6 GND 0.09fF
C424 a_10429_1050.n7 GND 0.33fF
C425 a_10429_1050.n8 GND 0.05fF
C426 a_14320_101.n0 GND 0.06fF
C427 a_14320_101.n1 GND 0.03fF
C428 a_14320_101.n2 GND 0.14fF
C429 a_14320_101.n3 GND 0.04fF
C430 a_14320_101.n4 GND 0.18fF
C431 a_3303_411.n0 GND 0.81fF
C432 a_3303_411.n1 GND 0.96fF
C433 a_3303_411.n2 GND 0.52fF
C434 a_3303_411.n3 GND 0.58fF
C435 a_3303_411.n4 GND 0.73fF
C436 a_3303_411.n5 GND 0.89fF
C437 a_3303_411.t13 GND 0.67fF
C438 a_3303_411.n6 GND 0.56fF
C439 a_3303_411.n7 GND 2.50fF
C440 a_3303_411.n8 GND 0.56fF
C441 a_3303_411.t6 GND 0.78fF
C442 a_3303_411.n9 GND 0.60fF
C443 a_3303_411.n10 GND 11.50fF
C444 a_3303_411.n11 GND 0.67fF
C445 a_3303_411.n12 GND 0.13fF
C446 a_3303_411.n13 GND 0.40fF
C447 a_3303_411.n14 GND 0.07fF
C448 a_599_989.n0 GND 0.40fF
C449 a_599_989.n1 GND 0.43fF
C450 a_599_989.n2 GND 0.40fF
C451 a_599_989.t6 GND 0.57fF
C452 a_599_989.n3 GND 0.41fF
C453 a_599_989.n4 GND 1.09fF
C454 a_599_989.n5 GND 0.04fF
C455 a_599_989.n6 GND 0.06fF
C456 a_599_989.n7 GND 0.04fF
C457 a_599_989.n8 GND 0.32fF
C458 a_599_989.n9 GND 0.46fF
C459 a_599_989.n10 GND 0.67fF
C460 a_599_989.n11 GND 0.33fF
C461 a_599_989.n12 GND 0.57fF
C462 VDD.n0 GND 0.12fF
C463 VDD.n1 GND 0.03fF
C464 VDD.n2 GND 0.02fF
C465 VDD.n3 GND 0.05fF
C466 VDD.n4 GND 0.01fF
C467 VDD.n5 GND 0.02fF
C468 VDD.n6 GND 0.02fF
C469 VDD.n9 GND 0.02fF
C470 VDD.n10 GND 0.02fF
C471 VDD.n12 GND 0.02fF
C472 VDD.n14 GND 0.47fF
C473 VDD.n16 GND 0.03fF
C474 VDD.n17 GND 0.02fF
C475 VDD.n18 GND 0.02fF
C476 VDD.n19 GND 0.02fF
C477 VDD.n20 GND 0.04fF
C478 VDD.n21 GND 0.28fF
C479 VDD.n22 GND 0.02fF
C480 VDD.n23 GND 0.03fF
C481 VDD.n24 GND 0.06fF
C482 VDD.n25 GND 0.15fF
C483 VDD.n26 GND 0.21fF
C484 VDD.n27 GND 0.01fF
C485 VDD.n28 GND 0.01fF
C486 VDD.n29 GND 0.07fF
C487 VDD.n30 GND 0.17fF
C488 VDD.n31 GND 0.01fF
C489 VDD.n32 GND 0.03fF
C490 VDD.n33 GND 0.03fF
C491 VDD.n34 GND 0.15fF
C492 VDD.n35 GND 0.21fF
C493 VDD.n36 GND 0.01fF
C494 VDD.n37 GND 0.06fF
C495 VDD.n38 GND 0.01fF
C496 VDD.n39 GND 0.02fF
C497 VDD.n40 GND 0.28fF
C498 VDD.n41 GND 0.01fF
C499 VDD.n42 GND 0.02fF
C500 VDD.n43 GND 0.03fF
C501 VDD.n44 GND 0.02fF
C502 VDD.n45 GND 0.02fF
C503 VDD.n46 GND 0.02fF
C504 VDD.n47 GND 0.19fF
C505 VDD.n48 GND 0.04fF
C506 VDD.n49 GND 0.04fF
C507 VDD.n50 GND 0.02fF
C508 VDD.n52 GND 0.02fF
C509 VDD.n53 GND 0.02fF
C510 VDD.n54 GND 0.02fF
C511 VDD.n55 GND 0.02fF
C512 VDD.n57 GND 0.02fF
C513 VDD.n58 GND 0.02fF
C514 VDD.n59 GND 0.02fF
C515 VDD.n61 GND 0.28fF
C516 VDD.n63 GND 0.02fF
C517 VDD.n64 GND 0.02fF
C518 VDD.n65 GND 0.03fF
C519 VDD.n66 GND 0.02fF
C520 VDD.n67 GND 0.28fF
C521 VDD.n68 GND 0.01fF
C522 VDD.n69 GND 0.02fF
C523 VDD.n70 GND 0.03fF
C524 VDD.n71 GND 0.28fF
C525 VDD.n72 GND 0.01fF
C526 VDD.n73 GND 0.02fF
C527 VDD.n74 GND 0.02fF
C528 VDD.n75 GND 0.28fF
C529 VDD.n76 GND 0.01fF
C530 VDD.n77 GND 0.02fF
C531 VDD.n78 GND 0.02fF
C532 VDD.n79 GND 0.31fF
C533 VDD.n80 GND 0.01fF
C534 VDD.n81 GND 0.03fF
C535 VDD.n82 GND 0.03fF
C536 VDD.n83 GND 0.31fF
C537 VDD.n84 GND 0.01fF
C538 VDD.n85 GND 0.03fF
C539 VDD.n86 GND 0.03fF
C540 VDD.n87 GND 0.28fF
C541 VDD.n88 GND 0.01fF
C542 VDD.n89 GND 0.02fF
C543 VDD.n90 GND 0.02fF
C544 VDD.n91 GND 0.28fF
C545 VDD.n92 GND 0.01fF
C546 VDD.n93 GND 0.02fF
C547 VDD.n94 GND 0.02fF
C548 VDD.n95 GND 0.28fF
C549 VDD.n96 GND 0.01fF
C550 VDD.n97 GND 0.02fF
C551 VDD.n98 GND 0.03fF
C552 VDD.n99 GND 0.02fF
C553 VDD.n100 GND 0.02fF
C554 VDD.n101 GND 0.02fF
C555 VDD.n102 GND 0.22fF
C556 VDD.n103 GND 0.04fF
C557 VDD.n104 GND 0.03fF
C558 VDD.n105 GND 0.02fF
C559 VDD.n106 GND 0.02fF
C560 VDD.n107 GND 0.02fF
C561 VDD.n108 GND 0.03fF
C562 VDD.n109 GND 0.02fF
C563 VDD.n111 GND 0.02fF
C564 VDD.n112 GND 0.02fF
C565 VDD.n113 GND 0.02fF
C566 VDD.n115 GND 0.28fF
C567 VDD.n117 GND 0.02fF
C568 VDD.n118 GND 0.02fF
C569 VDD.n119 GND 0.03fF
C570 VDD.n120 GND 0.02fF
C571 VDD.n121 GND 0.28fF
C572 VDD.n122 GND 0.01fF
C573 VDD.n123 GND 0.02fF
C574 VDD.n124 GND 0.03fF
C575 VDD.n125 GND 0.28fF
C576 VDD.n126 GND 0.01fF
C577 VDD.n127 GND 0.02fF
C578 VDD.n128 GND 0.02fF
C579 VDD.n129 GND 0.28fF
C580 VDD.n130 GND 0.01fF
C581 VDD.n131 GND 0.02fF
C582 VDD.n132 GND 0.02fF
C583 VDD.n133 GND 0.31fF
C584 VDD.n134 GND 0.01fF
C585 VDD.n135 GND 0.03fF
C586 VDD.n136 GND 0.03fF
C587 VDD.n137 GND 0.31fF
C588 VDD.n138 GND 0.01fF
C589 VDD.n139 GND 0.03fF
C590 VDD.n140 GND 0.03fF
C591 VDD.n141 GND 0.28fF
C592 VDD.n142 GND 0.01fF
C593 VDD.n143 GND 0.02fF
C594 VDD.n144 GND 0.02fF
C595 VDD.n145 GND 0.28fF
C596 VDD.n146 GND 0.01fF
C597 VDD.n147 GND 0.02fF
C598 VDD.n148 GND 0.02fF
C599 VDD.n149 GND 0.28fF
C600 VDD.n150 GND 0.01fF
C601 VDD.n151 GND 0.02fF
C602 VDD.n152 GND 0.03fF
C603 VDD.n153 GND 0.02fF
C604 VDD.n154 GND 0.02fF
C605 VDD.n155 GND 0.02fF
C606 VDD.n156 GND 0.22fF
C607 VDD.n157 GND 0.04fF
C608 VDD.n158 GND 0.03fF
C609 VDD.n159 GND 0.02fF
C610 VDD.n160 GND 0.02fF
C611 VDD.n161 GND 0.02fF
C612 VDD.n162 GND 0.03fF
C613 VDD.n163 GND 0.02fF
C614 VDD.n165 GND 0.02fF
C615 VDD.n166 GND 0.02fF
C616 VDD.n167 GND 0.02fF
C617 VDD.n169 GND 0.28fF
C618 VDD.n171 GND 0.02fF
C619 VDD.n172 GND 0.02fF
C620 VDD.n173 GND 0.03fF
C621 VDD.n174 GND 0.02fF
C622 VDD.n175 GND 0.28fF
C623 VDD.n176 GND 0.01fF
C624 VDD.n177 GND 0.02fF
C625 VDD.n178 GND 0.03fF
C626 VDD.n179 GND 0.06fF
C627 VDD.n180 GND 0.25fF
C628 VDD.n181 GND 0.01fF
C629 VDD.n182 GND 0.01fF
C630 VDD.n183 GND 0.02fF
C631 VDD.n184 GND 0.14fF
C632 VDD.n185 GND 0.17fF
C633 VDD.n186 GND 0.01fF
C634 VDD.n187 GND 0.02fF
C635 VDD.n188 GND 0.02fF
C636 VDD.n189 GND 0.11fF
C637 VDD.n190 GND 0.03fF
C638 VDD.n191 GND 0.31fF
C639 VDD.n192 GND 0.01fF
C640 VDD.n193 GND 0.02fF
C641 VDD.n194 GND 0.03fF
C642 VDD.n195 GND 0.17fF
C643 VDD.n196 GND 0.14fF
C644 VDD.n197 GND 0.01fF
C645 VDD.n198 GND 0.02fF
C646 VDD.n199 GND 0.03fF
C647 VDD.n200 GND 0.14fF
C648 VDD.n201 GND 0.17fF
C649 VDD.n202 GND 0.01fF
C650 VDD.n203 GND 0.02fF
C651 VDD.n204 GND 0.02fF
C652 VDD.n205 GND 0.06fF
C653 VDD.n206 GND 0.25fF
C654 VDD.n207 GND 0.01fF
C655 VDD.n208 GND 0.01fF
C656 VDD.n209 GND 0.02fF
C657 VDD.n210 GND 0.28fF
C658 VDD.n211 GND 0.01fF
C659 VDD.n212 GND 0.02fF
C660 VDD.n213 GND 0.03fF
C661 VDD.n214 GND 0.02fF
C662 VDD.n215 GND 0.02fF
C663 VDD.n216 GND 0.02fF
C664 VDD.n217 GND 0.22fF
C665 VDD.n218 GND 0.04fF
C666 VDD.n219 GND 0.03fF
C667 VDD.n220 GND 0.02fF
C668 VDD.n221 GND 0.02fF
C669 VDD.n222 GND 0.02fF
C670 VDD.n223 GND 0.03fF
C671 VDD.n224 GND 0.02fF
C672 VDD.n226 GND 0.02fF
C673 VDD.n227 GND 0.02fF
C674 VDD.n228 GND 0.02fF
C675 VDD.n230 GND 0.28fF
C676 VDD.n232 GND 0.02fF
C677 VDD.n233 GND 0.02fF
C678 VDD.n234 GND 0.03fF
C679 VDD.n235 GND 0.02fF
C680 VDD.n236 GND 0.28fF
C681 VDD.n237 GND 0.01fF
C682 VDD.n238 GND 0.02fF
C683 VDD.n239 GND 0.03fF
C684 VDD.n240 GND 0.06fF
C685 VDD.n241 GND 0.25fF
C686 VDD.n242 GND 0.01fF
C687 VDD.n243 GND 0.01fF
C688 VDD.n244 GND 0.02fF
C689 VDD.n245 GND 0.14fF
C690 VDD.n246 GND 0.17fF
C691 VDD.n247 GND 0.01fF
C692 VDD.n248 GND 0.02fF
C693 VDD.n249 GND 0.02fF
C694 VDD.n250 GND 0.11fF
C695 VDD.n251 GND 0.03fF
C696 VDD.n252 GND 0.31fF
C697 VDD.n253 GND 0.01fF
C698 VDD.n254 GND 0.02fF
C699 VDD.n255 GND 0.03fF
C700 VDD.n256 GND 0.17fF
C701 VDD.n257 GND 0.14fF
C702 VDD.n258 GND 0.01fF
C703 VDD.n259 GND 0.02fF
C704 VDD.n260 GND 0.03fF
C705 VDD.n261 GND 0.14fF
C706 VDD.n262 GND 0.17fF
C707 VDD.n263 GND 0.01fF
C708 VDD.n264 GND 0.02fF
C709 VDD.n265 GND 0.02fF
C710 VDD.n266 GND 0.06fF
C711 VDD.n267 GND 0.25fF
C712 VDD.n268 GND 0.01fF
C713 VDD.n269 GND 0.01fF
C714 VDD.n270 GND 0.02fF
C715 VDD.n271 GND 0.28fF
C716 VDD.n272 GND 0.01fF
C717 VDD.n273 GND 0.02fF
C718 VDD.n274 GND 0.03fF
C719 VDD.n275 GND 0.02fF
C720 VDD.n276 GND 0.02fF
C721 VDD.n277 GND 0.02fF
C722 VDD.n278 GND 0.22fF
C723 VDD.n279 GND 0.04fF
C724 VDD.n280 GND 0.03fF
C725 VDD.n281 GND 0.02fF
C726 VDD.n282 GND 0.02fF
C727 VDD.n283 GND 0.02fF
C728 VDD.n284 GND 0.03fF
C729 VDD.n285 GND 0.02fF
C730 VDD.n287 GND 0.02fF
C731 VDD.n288 GND 0.02fF
C732 VDD.n289 GND 0.02fF
C733 VDD.n291 GND 0.28fF
C734 VDD.n293 GND 0.02fF
C735 VDD.n294 GND 0.02fF
C736 VDD.n295 GND 0.03fF
C737 VDD.n296 GND 0.02fF
C738 VDD.n297 GND 0.28fF
C739 VDD.n298 GND 0.01fF
C740 VDD.n299 GND 0.02fF
C741 VDD.n300 GND 0.03fF
C742 VDD.n301 GND 0.06fF
C743 VDD.n302 GND 0.25fF
C744 VDD.n303 GND 0.01fF
C745 VDD.n304 GND 0.01fF
C746 VDD.n305 GND 0.02fF
C747 VDD.n306 GND 0.14fF
C748 VDD.n307 GND 0.17fF
C749 VDD.n308 GND 0.01fF
C750 VDD.n309 GND 0.02fF
C751 VDD.n310 GND 0.02fF
C752 VDD.n311 GND 0.11fF
C753 VDD.n312 GND 0.03fF
C754 VDD.n313 GND 0.31fF
C755 VDD.n314 GND 0.01fF
C756 VDD.n315 GND 0.02fF
C757 VDD.n316 GND 0.03fF
C758 VDD.n317 GND 0.17fF
C759 VDD.n318 GND 0.14fF
C760 VDD.n319 GND 0.01fF
C761 VDD.n320 GND 0.02fF
C762 VDD.n321 GND 0.03fF
C763 VDD.n322 GND 0.14fF
C764 VDD.n323 GND 0.17fF
C765 VDD.n324 GND 0.01fF
C766 VDD.n325 GND 0.02fF
C767 VDD.n326 GND 0.02fF
C768 VDD.n327 GND 0.06fF
C769 VDD.n328 GND 0.25fF
C770 VDD.n329 GND 0.01fF
C771 VDD.n330 GND 0.01fF
C772 VDD.n331 GND 0.02fF
C773 VDD.n332 GND 0.28fF
C774 VDD.n333 GND 0.01fF
C775 VDD.n334 GND 0.02fF
C776 VDD.n335 GND 0.03fF
C777 VDD.n336 GND 0.02fF
C778 VDD.n337 GND 0.02fF
C779 VDD.n338 GND 0.02fF
C780 VDD.n339 GND 0.22fF
C781 VDD.n340 GND 0.04fF
C782 VDD.n341 GND 0.03fF
C783 VDD.n342 GND 0.02fF
C784 VDD.n343 GND 0.02fF
C785 VDD.n344 GND 0.02fF
C786 VDD.n345 GND 0.03fF
C787 VDD.n346 GND 0.02fF
C788 VDD.n348 GND 0.02fF
C789 VDD.n349 GND 0.02fF
C790 VDD.n350 GND 0.02fF
C791 VDD.n352 GND 0.28fF
C792 VDD.n354 GND 0.02fF
C793 VDD.n355 GND 0.02fF
C794 VDD.n356 GND 0.03fF
C795 VDD.n357 GND 0.02fF
C796 VDD.n358 GND 0.28fF
C797 VDD.n359 GND 0.01fF
C798 VDD.n360 GND 0.02fF
C799 VDD.n361 GND 0.03fF
C800 VDD.n362 GND 0.06fF
C801 VDD.n363 GND 0.25fF
C802 VDD.n364 GND 0.01fF
C803 VDD.n365 GND 0.01fF
C804 VDD.n366 GND 0.02fF
C805 VDD.n367 GND 0.14fF
C806 VDD.n368 GND 0.17fF
C807 VDD.n369 GND 0.01fF
C808 VDD.n370 GND 0.02fF
C809 VDD.n371 GND 0.02fF
C810 VDD.n372 GND 0.11fF
C811 VDD.n373 GND 0.03fF
C812 VDD.n374 GND 0.31fF
C813 VDD.n375 GND 0.01fF
C814 VDD.n376 GND 0.02fF
C815 VDD.n377 GND 0.03fF
C816 VDD.n378 GND 0.17fF
C817 VDD.n379 GND 0.14fF
C818 VDD.n380 GND 0.01fF
C819 VDD.n381 GND 0.02fF
C820 VDD.n382 GND 0.03fF
C821 VDD.n383 GND 0.14fF
C822 VDD.n384 GND 0.17fF
C823 VDD.n385 GND 0.01fF
C824 VDD.n386 GND 0.02fF
C825 VDD.n387 GND 0.02fF
C826 VDD.n388 GND 0.06fF
C827 VDD.n389 GND 0.25fF
C828 VDD.n390 GND 0.01fF
C829 VDD.n391 GND 0.01fF
C830 VDD.n392 GND 0.02fF
C831 VDD.n393 GND 0.28fF
C832 VDD.n394 GND 0.01fF
C833 VDD.n395 GND 0.02fF
C834 VDD.n396 GND 0.03fF
C835 VDD.n397 GND 0.02fF
C836 VDD.n398 GND 0.02fF
C837 VDD.n399 GND 0.02fF
C838 VDD.n400 GND 0.22fF
C839 VDD.n401 GND 0.04fF
C840 VDD.n402 GND 0.03fF
C841 VDD.n403 GND 0.02fF
C842 VDD.n404 GND 0.02fF
C843 VDD.n405 GND 0.02fF
C844 VDD.n406 GND 0.03fF
C845 VDD.n407 GND 0.02fF
C846 VDD.n409 GND 0.02fF
C847 VDD.n410 GND 0.02fF
C848 VDD.n411 GND 0.02fF
C849 VDD.n413 GND 0.28fF
C850 VDD.n415 GND 0.02fF
C851 VDD.n416 GND 0.02fF
C852 VDD.n417 GND 0.03fF
C853 VDD.n418 GND 0.02fF
C854 VDD.n419 GND 0.28fF
C855 VDD.n420 GND 0.01fF
C856 VDD.n421 GND 0.02fF
C857 VDD.n422 GND 0.03fF
C858 VDD.n423 GND 0.06fF
C859 VDD.n424 GND 0.25fF
C860 VDD.n425 GND 0.01fF
C861 VDD.n426 GND 0.01fF
C862 VDD.n427 GND 0.02fF
C863 VDD.n428 GND 0.14fF
C864 VDD.n429 GND 0.17fF
C865 VDD.n430 GND 0.01fF
C866 VDD.n431 GND 0.02fF
C867 VDD.n432 GND 0.02fF
C868 VDD.n433 GND 0.11fF
C869 VDD.n434 GND 0.03fF
C870 VDD.n435 GND 0.31fF
C871 VDD.n436 GND 0.01fF
C872 VDD.n437 GND 0.02fF
C873 VDD.n438 GND 0.03fF
C874 VDD.n439 GND 0.17fF
C875 VDD.n440 GND 0.14fF
C876 VDD.n441 GND 0.01fF
C877 VDD.n442 GND 0.02fF
C878 VDD.n443 GND 0.03fF
C879 VDD.n444 GND 0.14fF
C880 VDD.n445 GND 0.17fF
C881 VDD.n446 GND 0.01fF
C882 VDD.n447 GND 0.02fF
C883 VDD.n448 GND 0.02fF
C884 VDD.n449 GND 0.06fF
C885 VDD.n450 GND 0.25fF
C886 VDD.n451 GND 0.01fF
C887 VDD.n452 GND 0.01fF
C888 VDD.n453 GND 0.02fF
C889 VDD.n454 GND 0.28fF
C890 VDD.n455 GND 0.01fF
C891 VDD.n456 GND 0.02fF
C892 VDD.n457 GND 0.03fF
C893 VDD.n458 GND 0.02fF
C894 VDD.n459 GND 0.02fF
C895 VDD.n460 GND 0.02fF
C896 VDD.n461 GND 0.22fF
C897 VDD.n462 GND 0.04fF
C898 VDD.n463 GND 0.03fF
C899 VDD.n464 GND 0.02fF
C900 VDD.n465 GND 0.02fF
C901 VDD.n466 GND 0.02fF
C902 VDD.n467 GND 0.03fF
C903 VDD.n468 GND 0.02fF
C904 VDD.n470 GND 0.02fF
C905 VDD.n471 GND 0.02fF
C906 VDD.n472 GND 0.02fF
C907 VDD.n474 GND 0.28fF
C908 VDD.n476 GND 0.02fF
C909 VDD.n477 GND 0.02fF
C910 VDD.n478 GND 0.03fF
C911 VDD.n479 GND 0.02fF
C912 VDD.n480 GND 0.28fF
C913 VDD.n481 GND 0.01fF
C914 VDD.n482 GND 0.02fF
C915 VDD.n483 GND 0.03fF
C916 VDD.n484 GND 0.06fF
C917 VDD.n485 GND 0.25fF
C918 VDD.n486 GND 0.01fF
C919 VDD.n487 GND 0.01fF
C920 VDD.n488 GND 0.02fF
C921 VDD.n489 GND 0.14fF
C922 VDD.n490 GND 0.17fF
C923 VDD.n491 GND 0.01fF
C924 VDD.n492 GND 0.02fF
C925 VDD.n493 GND 0.02fF
C926 VDD.n494 GND 0.11fF
C927 VDD.n495 GND 0.03fF
C928 VDD.n496 GND 0.31fF
C929 VDD.n497 GND 0.01fF
C930 VDD.n498 GND 0.02fF
C931 VDD.n499 GND 0.03fF
C932 VDD.n500 GND 0.17fF
C933 VDD.n501 GND 0.14fF
C934 VDD.n502 GND 0.01fF
C935 VDD.n503 GND 0.02fF
C936 VDD.n504 GND 0.03fF
C937 VDD.n505 GND 0.14fF
C938 VDD.n506 GND 0.17fF
C939 VDD.n507 GND 0.01fF
C940 VDD.n508 GND 0.02fF
C941 VDD.n509 GND 0.02fF
C942 VDD.n510 GND 0.06fF
C943 VDD.n511 GND 0.25fF
C944 VDD.n512 GND 0.01fF
C945 VDD.n513 GND 0.01fF
C946 VDD.n514 GND 0.02fF
C947 VDD.n515 GND 0.28fF
C948 VDD.n516 GND 0.01fF
C949 VDD.n517 GND 0.02fF
C950 VDD.n518 GND 0.03fF
C951 VDD.n519 GND 0.02fF
C952 VDD.n520 GND 0.02fF
C953 VDD.n521 GND 0.02fF
C954 VDD.n522 GND 0.27fF
C955 VDD.n523 GND 0.04fF
C956 VDD.n524 GND 0.03fF
C957 VDD.n525 GND 0.02fF
C958 VDD.n526 GND 0.02fF
C959 VDD.n527 GND 0.02fF
C960 VDD.n528 GND 0.03fF
C961 VDD.n529 GND 0.02fF
C962 VDD.n531 GND 0.02fF
C963 VDD.n532 GND 0.02fF
C964 VDD.n533 GND 0.02fF
C965 VDD.n535 GND 0.28fF
C966 VDD.n537 GND 0.02fF
C967 VDD.n538 GND 0.02fF
C968 VDD.n539 GND 0.03fF
C969 VDD.n540 GND 0.02fF
C970 VDD.n541 GND 0.28fF
C971 VDD.n542 GND 0.01fF
C972 VDD.n543 GND 0.02fF
C973 VDD.n544 GND 0.03fF
C974 VDD.n545 GND 0.28fF
C975 VDD.n546 GND 0.01fF
C976 VDD.n547 GND 0.02fF
C977 VDD.n548 GND 0.02fF
C978 VDD.n549 GND 0.23fF
C979 VDD.n550 GND 0.01fF
C980 VDD.n551 GND 0.07fF
C981 VDD.n552 GND 0.02fF
C982 VDD.n553 GND 0.14fF
C983 VDD.n554 GND 0.17fF
C984 VDD.n555 GND 0.01fF
C985 VDD.n556 GND 0.02fF
C986 VDD.n557 GND 0.02fF
C987 VDD.n558 GND 0.14fF
C988 VDD.n559 GND 0.16fF
C989 VDD.n560 GND 0.01fF
C990 VDD.n561 GND 0.11fF
C991 VDD.n562 GND 0.02fF
C992 VDD.n563 GND 0.02fF
C993 VDD.n564 GND 0.02fF
C994 VDD.n565 GND 0.18fF
C995 VDD.n566 GND 0.15fF
C996 VDD.n567 GND 0.02fF
C997 VDD.n568 GND 0.02fF
C998 VDD.n569 GND 0.03fF
C999 VDD.n570 GND 0.18fF
C1000 VDD.n571 GND 0.15fF
C1001 VDD.n572 GND 0.02fF
C1002 VDD.n573 GND 0.02fF
C1003 VDD.n574 GND 0.03fF
C1004 VDD.n575 GND 0.11fF
C1005 VDD.n576 GND 0.02fF
C1006 VDD.n577 GND 0.14fF
C1007 VDD.n578 GND 0.16fF
C1008 VDD.n579 GND 0.01fF
C1009 VDD.n580 GND 0.02fF
C1010 VDD.n581 GND 0.02fF
C1011 VDD.n582 GND 0.14fF
C1012 VDD.n583 GND 0.17fF
C1013 VDD.n584 GND 0.01fF
C1014 VDD.n585 GND 0.02fF
C1015 VDD.n586 GND 0.02fF
C1016 VDD.n587 GND 0.06fF
C1017 VDD.n588 GND 0.23fF
C1018 VDD.n589 GND 0.01fF
C1019 VDD.n590 GND 0.01fF
C1020 VDD.n591 GND 0.02fF
C1021 VDD.n592 GND 0.28fF
C1022 VDD.n593 GND 0.01fF
C1023 VDD.n594 GND 0.02fF
C1024 VDD.n595 GND 0.02fF
C1025 VDD.n596 GND 0.28fF
C1026 VDD.n597 GND 0.01fF
C1027 VDD.n598 GND 0.02fF
C1028 VDD.n599 GND 0.03fF
C1029 VDD.n600 GND 0.02fF
C1030 VDD.n601 GND 0.02fF
C1031 VDD.n602 GND 0.02fF
C1032 VDD.n603 GND 0.27fF
C1033 VDD.n604 GND 0.04fF
C1034 VDD.n605 GND 0.03fF
C1035 VDD.n606 GND 0.02fF
C1036 VDD.n607 GND 0.02fF
C1037 VDD.n608 GND 0.02fF
C1038 VDD.n609 GND 0.03fF
C1039 VDD.n610 GND 0.02fF
C1040 VDD.n612 GND 0.02fF
C1041 VDD.n613 GND 0.02fF
C1042 VDD.n614 GND 0.02fF
C1043 VDD.n616 GND 0.28fF
C1044 VDD.n618 GND 0.02fF
C1045 VDD.n619 GND 0.02fF
C1046 VDD.n620 GND 0.03fF
C1047 VDD.n621 GND 0.02fF
C1048 VDD.n622 GND 0.28fF
C1049 VDD.n623 GND 0.01fF
C1050 VDD.n624 GND 0.02fF
C1051 VDD.n625 GND 0.03fF
C1052 VDD.n626 GND 0.06fF
C1053 VDD.n627 GND 0.25fF
C1054 VDD.n628 GND 0.01fF
C1055 VDD.n629 GND 0.01fF
C1056 VDD.n630 GND 0.02fF
C1057 VDD.n631 GND 0.14fF
C1058 VDD.n632 GND 0.17fF
C1059 VDD.n633 GND 0.01fF
C1060 VDD.n634 GND 0.02fF
C1061 VDD.n635 GND 0.02fF
C1062 VDD.n636 GND 0.11fF
C1063 VDD.n637 GND 0.03fF
C1064 VDD.n638 GND 0.31fF
C1065 VDD.n639 GND 0.01fF
C1066 VDD.n640 GND 0.02fF
C1067 VDD.n641 GND 0.03fF
C1068 VDD.n642 GND 0.17fF
C1069 VDD.n643 GND 0.14fF
C1070 VDD.n644 GND 0.01fF
C1071 VDD.n645 GND 0.02fF
C1072 VDD.n646 GND 0.03fF
C1073 VDD.n647 GND 0.14fF
C1074 VDD.n648 GND 0.17fF
C1075 VDD.n649 GND 0.01fF
C1076 VDD.n650 GND 0.02fF
C1077 VDD.n651 GND 0.02fF
C1078 VDD.n652 GND 0.06fF
C1079 VDD.n653 GND 0.25fF
C1080 VDD.n654 GND 0.01fF
C1081 VDD.n655 GND 0.01fF
C1082 VDD.n656 GND 0.02fF
C1083 VDD.n657 GND 0.28fF
C1084 VDD.n658 GND 0.01fF
C1085 VDD.n659 GND 0.02fF
C1086 VDD.n660 GND 0.03fF
C1087 VDD.n661 GND 0.02fF
C1088 VDD.n662 GND 0.02fF
C1089 VDD.n663 GND 0.02fF
C1090 VDD.n664 GND 0.22fF
C1091 VDD.n665 GND 0.04fF
C1092 VDD.n666 GND 0.03fF
C1093 VDD.n667 GND 0.02fF
C1094 VDD.n668 GND 0.02fF
C1095 VDD.n669 GND 0.02fF
C1096 VDD.n670 GND 0.03fF
C1097 VDD.n671 GND 0.02fF
C1098 VDD.n673 GND 0.02fF
C1099 VDD.n674 GND 0.02fF
C1100 VDD.n675 GND 0.02fF
C1101 VDD.n677 GND 0.28fF
C1102 VDD.n679 GND 0.02fF
C1103 VDD.n680 GND 0.02fF
C1104 VDD.n681 GND 0.03fF
C1105 VDD.n682 GND 0.02fF
C1106 VDD.n683 GND 0.28fF
C1107 VDD.n684 GND 0.01fF
C1108 VDD.n685 GND 0.02fF
C1109 VDD.n686 GND 0.03fF
C1110 VDD.n687 GND 0.06fF
C1111 VDD.n688 GND 0.25fF
C1112 VDD.n689 GND 0.01fF
C1113 VDD.n690 GND 0.01fF
C1114 VDD.n691 GND 0.02fF
C1115 VDD.n692 GND 0.14fF
C1116 VDD.n693 GND 0.17fF
C1117 VDD.n694 GND 0.01fF
C1118 VDD.n695 GND 0.02fF
C1119 VDD.n696 GND 0.02fF
C1120 VDD.n697 GND 0.02fF
C1121 VDD.n698 GND 0.02fF
C1122 VDD.n699 GND 0.02fF
C1123 VDD.n700 GND 0.21fF
C1124 VDD.n701 GND 0.03fF
C1125 VDD.n702 GND 0.02fF
C1126 VDD.n703 GND 0.02fF
C1127 VDD.n704 GND 0.02fF
C1128 VDD.n705 GND 0.03fF
C1129 VDD.n706 GND 0.02fF
C1130 VDD.n708 GND 0.02fF
C1131 VDD.n709 GND 0.02fF
C1132 VDD.n710 GND 0.02fF
C1133 VDD.n712 GND 0.47fF
C1134 VDD.n714 GND 0.03fF
C1135 VDD.n715 GND 0.04fF
C1136 VDD.n716 GND 0.28fF
C1137 VDD.n717 GND 0.02fF
C1138 VDD.n718 GND 0.03fF
C1139 VDD.n719 GND 0.03fF
C1140 VDD.n720 GND 0.28fF
C1141 VDD.n721 GND 0.01fF
C1142 VDD.n722 GND 0.02fF
C1143 VDD.n723 GND 0.02fF
C1144 VDD.n724 GND 0.06fF
C1145 VDD.n725 GND 0.23fF
C1146 VDD.n726 GND 0.01fF
C1147 VDD.n727 GND 0.01fF
C1148 VDD.n728 GND 0.02fF
C1149 VDD.n729 GND 0.14fF
C1150 VDD.n730 GND 0.17fF
C1151 VDD.n731 GND 0.01fF
C1152 VDD.n732 GND 0.02fF
C1153 VDD.n733 GND 0.02fF
C1154 VDD.n734 GND 0.11fF
C1155 VDD.n735 GND 0.02fF
C1156 VDD.n736 GND 0.14fF
C1157 VDD.n737 GND 0.16fF
C1158 VDD.n738 GND 0.01fF
C1159 VDD.n739 GND 0.02fF
C1160 VDD.n740 GND 0.02fF
C1161 VDD.n741 GND 0.18fF
C1162 VDD.n742 GND 0.15fF
C1163 VDD.n743 GND 0.02fF
C1164 VDD.n744 GND 0.02fF
C1165 VDD.n745 GND 0.03fF
C1166 VDD.n746 GND 0.18fF
C1167 VDD.n747 GND 0.15fF
C1168 VDD.n748 GND 0.02fF
C1169 VDD.n749 GND 0.02fF
C1170 VDD.n750 GND 0.03fF
C1171 VDD.n751 GND 0.14fF
C1172 VDD.n752 GND 0.16fF
C1173 VDD.n753 GND 0.01fF
C1174 VDD.n754 GND 0.11fF
C1175 VDD.n755 GND 0.02fF
C1176 VDD.n756 GND 0.02fF
C1177 VDD.n757 GND 0.02fF
C1178 VDD.n758 GND 0.14fF
C1179 VDD.n759 GND 0.17fF
C1180 VDD.n760 GND 0.01fF
C1181 VDD.n761 GND 0.02fF
C1182 VDD.n762 GND 0.02fF
C1183 VDD.n763 GND 0.23fF
C1184 VDD.n764 GND 0.01fF
C1185 VDD.n765 GND 0.07fF
C1186 VDD.n766 GND 0.02fF
C1187 VDD.n767 GND 0.28fF
C1188 VDD.n768 GND 0.01fF
C1189 VDD.n769 GND 0.02fF
C1190 VDD.n770 GND 0.02fF
C1191 VDD.n771 GND 0.28fF
C1192 VDD.n772 GND 0.01fF
C1193 VDD.n773 GND 0.02fF
C1194 VDD.n774 GND 0.03fF
C1195 VDD.n775 GND 0.02fF
C1196 VDD.n776 GND 0.02fF
C1197 VDD.n777 GND 0.02fF
C1198 VDD.n778 GND 0.02fF
C1199 VDD.n779 GND 0.02fF
C1200 VDD.n780 GND 0.02fF
C1201 VDD.n782 GND 0.02fF
C1202 VDD.n783 GND 0.02fF
C1203 VDD.n784 GND 0.02fF
C1204 VDD.n785 GND 0.02fF
C1205 VDD.n787 GND 0.04fF
C1206 VDD.n788 GND 0.02fF
C1207 VDD.n789 GND 0.27fF
C1208 VDD.n790 GND 0.04fF
C1209 VDD.n792 GND 0.28fF
C1210 VDD.n794 GND 0.02fF
C1211 VDD.n795 GND 0.02fF
C1212 VDD.n796 GND 0.03fF
C1213 VDD.n797 GND 0.02fF
C1214 VDD.n798 GND 0.28fF
C1215 VDD.n799 GND 0.01fF
C1216 VDD.n800 GND 0.02fF
C1217 VDD.n801 GND 0.03fF
C1218 VDD.n802 GND 0.06fF
C1219 VDD.n803 GND 0.25fF
C1220 VDD.n804 GND 0.01fF
C1221 VDD.n805 GND 0.01fF
C1222 VDD.n806 GND 0.02fF
C1223 VDD.n807 GND 0.14fF
C1224 VDD.n808 GND 0.17fF
C1225 VDD.n809 GND 0.01fF
C1226 VDD.n810 GND 0.02fF
C1227 VDD.n811 GND 0.02fF
C1228 VDD.n812 GND 0.17fF
C1229 VDD.n813 GND 0.14fF
C1230 VDD.n814 GND 0.01fF
C1231 VDD.n815 GND 0.02fF
C1232 VDD.n816 GND 0.03fF
C1233 VDD.n817 GND 0.11fF
C1234 VDD.n818 GND 0.03fF
C1235 VDD.n819 GND 0.31fF
C1236 VDD.n820 GND 0.01fF
C1237 VDD.n821 GND 0.02fF
C1238 VDD.n822 GND 0.03fF
C1239 VDD.n823 GND 0.14fF
C1240 VDD.n824 GND 0.17fF
C1241 VDD.n825 GND 0.01fF
C1242 VDD.n826 GND 0.02fF
C1243 VDD.n827 GND 0.02fF
C1244 VDD.n828 GND 0.06fF
C1245 VDD.n829 GND 0.25fF
C1246 VDD.n830 GND 0.01fF
C1247 VDD.n831 GND 0.01fF
C1248 VDD.n832 GND 0.02fF
C1249 VDD.n833 GND 0.28fF
C1250 VDD.n834 GND 0.01fF
C1251 VDD.n835 GND 0.02fF
C1252 VDD.n836 GND 0.03fF
C1253 VDD.n837 GND 0.02fF
C1254 VDD.n838 GND 0.02fF
C1255 VDD.n839 GND 0.02fF
C1256 VDD.n840 GND 0.22fF
C1257 VDD.n841 GND 0.04fF
C1258 VDD.n842 GND 0.03fF
C1259 VDD.n843 GND 0.02fF
C1260 VDD.n844 GND 0.02fF
C1261 VDD.n845 GND 0.02fF
C1262 VDD.n846 GND 0.03fF
C1263 VDD.n847 GND 0.02fF
C1264 VDD.n849 GND 0.02fF
C1265 VDD.n850 GND 0.02fF
C1266 VDD.n851 GND 0.02fF
C1267 VDD.n853 GND 0.28fF
C1268 VDD.n855 GND 0.02fF
C1269 VDD.n856 GND 0.02fF
C1270 VDD.n857 GND 0.03fF
C1271 VDD.n858 GND 0.02fF
C1272 VDD.n859 GND 0.28fF
C1273 VDD.n860 GND 0.01fF
C1274 VDD.n861 GND 0.02fF
C1275 VDD.n862 GND 0.03fF
C1276 VDD.n863 GND 0.06fF
C1277 VDD.n864 GND 0.25fF
C1278 VDD.n865 GND 0.01fF
C1279 VDD.n866 GND 0.01fF
C1280 VDD.n867 GND 0.02fF
C1281 VDD.n868 GND 0.14fF
C1282 VDD.n869 GND 0.17fF
C1283 VDD.n870 GND 0.01fF
C1284 VDD.n871 GND 0.02fF
C1285 VDD.n872 GND 0.02fF
C1286 VDD.n873 GND 0.17fF
C1287 VDD.n874 GND 0.14fF
C1288 VDD.n875 GND 0.01fF
C1289 VDD.n876 GND 0.02fF
C1290 VDD.n877 GND 0.03fF
C1291 VDD.n878 GND 0.11fF
C1292 VDD.n879 GND 0.03fF
C1293 VDD.n880 GND 0.31fF
C1294 VDD.n881 GND 0.01fF
C1295 VDD.n882 GND 0.02fF
C1296 VDD.n883 GND 0.03fF
C1297 VDD.n884 GND 0.14fF
C1298 VDD.n885 GND 0.17fF
C1299 VDD.n886 GND 0.01fF
C1300 VDD.n887 GND 0.02fF
C1301 VDD.n888 GND 0.02fF
C1302 VDD.n889 GND 0.06fF
C1303 VDD.n890 GND 0.25fF
C1304 VDD.n891 GND 0.01fF
C1305 VDD.n892 GND 0.01fF
C1306 VDD.n893 GND 0.02fF
C1307 VDD.n894 GND 0.28fF
C1308 VDD.n895 GND 0.01fF
C1309 VDD.n896 GND 0.02fF
C1310 VDD.n897 GND 0.03fF
C1311 VDD.n898 GND 0.02fF
C1312 VDD.n899 GND 0.02fF
C1313 VDD.n900 GND 0.02fF
C1314 VDD.n901 GND 0.22fF
C1315 VDD.n902 GND 0.04fF
C1316 VDD.n903 GND 0.03fF
C1317 VDD.n904 GND 0.02fF
C1318 VDD.n905 GND 0.02fF
C1319 VDD.n906 GND 0.02fF
C1320 VDD.n907 GND 0.03fF
C1321 VDD.n908 GND 0.02fF
C1322 VDD.n910 GND 0.02fF
C1323 VDD.n911 GND 0.02fF
C1324 VDD.n912 GND 0.02fF
C1325 VDD.n914 GND 0.28fF
C1326 VDD.n916 GND 0.02fF
C1327 VDD.n917 GND 0.02fF
C1328 VDD.n918 GND 0.03fF
C1329 VDD.n919 GND 0.02fF
C1330 VDD.n920 GND 0.28fF
C1331 VDD.n921 GND 0.01fF
C1332 VDD.n922 GND 0.02fF
C1333 VDD.n923 GND 0.03fF
C1334 VDD.n924 GND 0.06fF
C1335 VDD.n925 GND 0.25fF
C1336 VDD.n926 GND 0.01fF
C1337 VDD.n927 GND 0.01fF
C1338 VDD.n928 GND 0.02fF
C1339 VDD.n929 GND 0.14fF
C1340 VDD.n930 GND 0.17fF
C1341 VDD.n931 GND 0.01fF
C1342 VDD.n932 GND 0.02fF
C1343 VDD.n933 GND 0.02fF
C1344 VDD.n934 GND 0.17fF
C1345 VDD.n935 GND 0.14fF
C1346 VDD.n936 GND 0.01fF
C1347 VDD.n937 GND 0.02fF
C1348 VDD.n938 GND 0.03fF
C1349 VDD.n939 GND 0.11fF
C1350 VDD.n940 GND 0.03fF
C1351 VDD.n941 GND 0.31fF
C1352 VDD.n942 GND 0.01fF
C1353 VDD.n943 GND 0.02fF
C1354 VDD.n944 GND 0.03fF
C1355 VDD.n945 GND 0.14fF
C1356 VDD.n946 GND 0.17fF
C1357 VDD.n947 GND 0.01fF
C1358 VDD.n948 GND 0.02fF
C1359 VDD.n949 GND 0.02fF
C1360 VDD.n950 GND 0.06fF
C1361 VDD.n951 GND 0.25fF
C1362 VDD.n952 GND 0.01fF
C1363 VDD.n953 GND 0.01fF
C1364 VDD.n954 GND 0.02fF
C1365 VDD.n955 GND 0.28fF
C1366 VDD.n956 GND 0.01fF
C1367 VDD.n957 GND 0.02fF
C1368 VDD.n958 GND 0.03fF
C1369 VDD.n959 GND 0.02fF
C1370 VDD.n960 GND 0.02fF
C1371 VDD.n961 GND 0.02fF
C1372 VDD.n962 GND 0.22fF
C1373 VDD.n963 GND 0.04fF
C1374 VDD.n964 GND 0.03fF
C1375 VDD.n965 GND 0.02fF
C1376 VDD.n966 GND 0.02fF
C1377 VDD.n967 GND 0.02fF
C1378 VDD.n968 GND 0.03fF
C1379 VDD.n969 GND 0.02fF
C1380 VDD.n971 GND 0.02fF
C1381 VDD.n972 GND 0.02fF
C1382 VDD.n973 GND 0.02fF
C1383 VDD.n975 GND 0.28fF
C1384 VDD.n977 GND 0.02fF
C1385 VDD.n978 GND 0.02fF
C1386 VDD.n979 GND 0.03fF
C1387 VDD.n980 GND 0.02fF
C1388 VDD.n981 GND 0.28fF
C1389 VDD.n982 GND 0.01fF
C1390 VDD.n983 GND 0.02fF
C1391 VDD.n984 GND 0.03fF
C1392 VDD.n985 GND 0.06fF
C1393 VDD.n986 GND 0.25fF
C1394 VDD.n987 GND 0.01fF
C1395 VDD.n988 GND 0.01fF
C1396 VDD.n989 GND 0.02fF
C1397 VDD.n990 GND 0.14fF
C1398 VDD.n991 GND 0.17fF
C1399 VDD.n992 GND 0.01fF
C1400 VDD.n993 GND 0.02fF
C1401 VDD.n994 GND 0.02fF
C1402 VDD.n995 GND 0.17fF
C1403 VDD.n996 GND 0.14fF
C1404 VDD.n997 GND 0.01fF
C1405 VDD.n998 GND 0.02fF
C1406 VDD.n999 GND 0.03fF
C1407 VDD.n1000 GND 0.11fF
C1408 VDD.n1001 GND 0.03fF
C1409 VDD.n1002 GND 0.31fF
C1410 VDD.n1003 GND 0.01fF
C1411 VDD.n1004 GND 0.02fF
C1412 VDD.n1005 GND 0.03fF
C1413 VDD.n1006 GND 0.14fF
C1414 VDD.n1007 GND 0.17fF
C1415 VDD.n1008 GND 0.01fF
C1416 VDD.n1009 GND 0.02fF
C1417 VDD.n1010 GND 0.02fF
C1418 VDD.n1011 GND 0.06fF
C1419 VDD.n1012 GND 0.25fF
C1420 VDD.n1013 GND 0.01fF
C1421 VDD.n1014 GND 0.01fF
C1422 VDD.n1015 GND 0.02fF
C1423 VDD.n1016 GND 0.28fF
C1424 VDD.n1017 GND 0.01fF
C1425 VDD.n1018 GND 0.02fF
C1426 VDD.n1019 GND 0.03fF
C1427 VDD.n1020 GND 0.02fF
C1428 VDD.n1021 GND 0.02fF
C1429 VDD.n1022 GND 0.02fF
C1430 VDD.n1023 GND 0.22fF
C1431 VDD.n1024 GND 0.04fF
C1432 VDD.n1025 GND 0.03fF
C1433 VDD.n1026 GND 0.02fF
C1434 VDD.n1027 GND 0.02fF
C1435 VDD.n1028 GND 0.02fF
C1436 VDD.n1029 GND 0.03fF
C1437 VDD.n1030 GND 0.02fF
C1438 VDD.n1032 GND 0.02fF
C1439 VDD.n1033 GND 0.02fF
C1440 VDD.n1034 GND 0.02fF
C1441 VDD.n1036 GND 0.28fF
C1442 VDD.n1038 GND 0.02fF
C1443 VDD.n1039 GND 0.02fF
C1444 VDD.n1040 GND 0.03fF
C1445 VDD.n1041 GND 0.02fF
C1446 VDD.n1042 GND 0.28fF
C1447 VDD.n1043 GND 0.01fF
C1448 VDD.n1044 GND 0.02fF
C1449 VDD.n1045 GND 0.03fF
C1450 VDD.n1046 GND 0.06fF
C1451 VDD.n1047 GND 0.25fF
C1452 VDD.n1048 GND 0.01fF
C1453 VDD.n1049 GND 0.01fF
C1454 VDD.n1050 GND 0.02fF
C1455 VDD.n1051 GND 0.14fF
C1456 VDD.n1052 GND 0.17fF
C1457 VDD.n1053 GND 0.01fF
C1458 VDD.n1054 GND 0.02fF
C1459 VDD.n1055 GND 0.02fF
C1460 VDD.n1056 GND 0.17fF
C1461 VDD.n1057 GND 0.14fF
C1462 VDD.n1058 GND 0.01fF
C1463 VDD.n1059 GND 0.02fF
C1464 VDD.n1060 GND 0.03fF
C1465 VDD.n1061 GND 0.11fF
C1466 VDD.n1062 GND 0.03fF
C1467 VDD.n1063 GND 0.31fF
C1468 VDD.n1064 GND 0.01fF
C1469 VDD.n1065 GND 0.02fF
C1470 VDD.n1066 GND 0.03fF
C1471 VDD.n1067 GND 0.14fF
C1472 VDD.n1068 GND 0.17fF
C1473 VDD.n1069 GND 0.01fF
C1474 VDD.n1070 GND 0.02fF
C1475 VDD.n1071 GND 0.02fF
C1476 VDD.n1072 GND 0.06fF
C1477 VDD.n1073 GND 0.25fF
C1478 VDD.n1074 GND 0.01fF
C1479 VDD.n1075 GND 0.01fF
C1480 VDD.n1076 GND 0.02fF
C1481 VDD.n1077 GND 0.28fF
C1482 VDD.n1078 GND 0.01fF
C1483 VDD.n1079 GND 0.02fF
C1484 VDD.n1080 GND 0.03fF
C1485 VDD.n1081 GND 0.02fF
C1486 VDD.n1082 GND 0.02fF
C1487 VDD.n1083 GND 0.02fF
C1488 VDD.n1084 GND 0.27fF
C1489 VDD.n1085 GND 0.04fF
C1490 VDD.n1086 GND 0.03fF
C1491 VDD.n1087 GND 0.02fF
C1492 VDD.n1088 GND 0.02fF
C1493 VDD.n1089 GND 0.02fF
C1494 VDD.n1090 GND 0.03fF
C1495 VDD.n1091 GND 0.02fF
C1496 VDD.n1093 GND 0.02fF
C1497 VDD.n1094 GND 0.02fF
C1498 VDD.n1095 GND 0.02fF
C1499 VDD.n1097 GND 0.28fF
C1500 VDD.n1099 GND 0.02fF
C1501 VDD.n1100 GND 0.02fF
C1502 VDD.n1101 GND 0.03fF
C1503 VDD.n1102 GND 0.02fF
C1504 VDD.n1103 GND 0.28fF
C1505 VDD.n1104 GND 0.01fF
C1506 VDD.n1105 GND 0.02fF
C1507 VDD.n1106 GND 0.03fF
C1508 VDD.n1107 GND 0.28fF
C1509 VDD.n1108 GND 0.01fF
C1510 VDD.n1109 GND 0.02fF
C1511 VDD.n1110 GND 0.02fF
C1512 VDD.n1111 GND 0.06fF
C1513 VDD.n1112 GND 0.23fF
C1514 VDD.n1113 GND 0.01fF
C1515 VDD.n1114 GND 0.01fF
C1516 VDD.n1115 GND 0.02fF
C1517 VDD.n1116 GND 0.14fF
C1518 VDD.n1117 GND 0.17fF
C1519 VDD.n1118 GND 0.01fF
C1520 VDD.n1119 GND 0.02fF
C1521 VDD.n1120 GND 0.02fF
C1522 VDD.n1121 GND 0.11fF
C1523 VDD.n1122 GND 0.02fF
C1524 VDD.n1123 GND 0.14fF
C1525 VDD.n1124 GND 0.16fF
C1526 VDD.n1125 GND 0.01fF
C1527 VDD.n1126 GND 0.02fF
C1528 VDD.n1127 GND 0.02fF
C1529 VDD.n1128 GND 0.18fF
C1530 VDD.n1129 GND 0.15fF
C1531 VDD.n1130 GND 0.02fF
C1532 VDD.n1131 GND 0.02fF
C1533 VDD.n1132 GND 0.03fF
C1534 VDD.n1133 GND 0.18fF
C1535 VDD.n1134 GND 0.15fF
C1536 VDD.n1135 GND 0.02fF
C1537 VDD.n1136 GND 0.02fF
C1538 VDD.n1137 GND 0.03fF
C1539 VDD.n1138 GND 0.14fF
C1540 VDD.n1139 GND 0.16fF
C1541 VDD.n1140 GND 0.01fF
C1542 VDD.n1141 GND 0.11fF
C1543 VDD.n1142 GND 0.02fF
C1544 VDD.n1143 GND 0.02fF
C1545 VDD.n1144 GND 0.02fF
C1546 VDD.n1145 GND 0.14fF
C1547 VDD.n1146 GND 0.17fF
C1548 VDD.n1147 GND 0.01fF
C1549 VDD.n1148 GND 0.02fF
C1550 VDD.n1149 GND 0.02fF
C1551 VDD.n1150 GND 0.23fF
C1552 VDD.n1151 GND 0.01fF
C1553 VDD.n1152 GND 0.07fF
C1554 VDD.n1153 GND 0.02fF
C1555 VDD.n1154 GND 0.28fF
C1556 VDD.n1155 GND 0.01fF
C1557 VDD.n1156 GND 0.02fF
C1558 VDD.n1157 GND 0.02fF
C1559 VDD.n1158 GND 0.28fF
C1560 VDD.n1159 GND 0.01fF
C1561 VDD.n1160 GND 0.02fF
C1562 VDD.n1161 GND 0.03fF
C1563 VDD.n1162 GND 0.02fF
C1564 VDD.n1163 GND 0.02fF
C1565 VDD.n1164 GND 0.02fF
C1566 VDD.n1165 GND 0.27fF
C1567 VDD.n1166 GND 0.04fF
C1568 VDD.n1167 GND 0.03fF
C1569 VDD.n1168 GND 0.02fF
C1570 VDD.n1169 GND 0.02fF
C1571 VDD.n1170 GND 0.02fF
C1572 VDD.n1171 GND 0.03fF
C1573 VDD.n1172 GND 0.02fF
C1574 VDD.n1174 GND 0.02fF
C1575 VDD.n1175 GND 0.02fF
C1576 VDD.n1176 GND 0.02fF
C1577 VDD.n1178 GND 0.28fF
C1578 VDD.n1180 GND 0.02fF
C1579 VDD.n1181 GND 0.02fF
C1580 VDD.n1182 GND 0.03fF
C1581 VDD.n1183 GND 0.02fF
C1582 VDD.n1184 GND 0.28fF
C1583 VDD.n1185 GND 0.01fF
C1584 VDD.n1186 GND 0.02fF
C1585 VDD.n1187 GND 0.03fF
C1586 VDD.n1188 GND 0.06fF
C1587 VDD.n1189 GND 0.25fF
C1588 VDD.n1190 GND 0.01fF
C1589 VDD.n1191 GND 0.01fF
C1590 VDD.n1192 GND 0.02fF
C1591 VDD.n1193 GND 0.14fF
C1592 VDD.n1194 GND 0.17fF
C1593 VDD.n1195 GND 0.01fF
C1594 VDD.n1196 GND 0.02fF
C1595 VDD.n1197 GND 0.02fF
C1596 VDD.n1198 GND 0.17fF
C1597 VDD.n1199 GND 0.14fF
C1598 VDD.n1200 GND 0.01fF
C1599 VDD.n1201 GND 0.02fF
C1600 VDD.n1202 GND 0.03fF
C1601 VDD.n1203 GND 0.11fF
C1602 VDD.n1204 GND 0.03fF
C1603 VDD.n1205 GND 0.31fF
C1604 VDD.n1206 GND 0.01fF
C1605 VDD.n1207 GND 0.02fF
C1606 VDD.n1208 GND 0.03fF
C1607 VDD.n1209 GND 0.14fF
C1608 VDD.n1210 GND 0.17fF
C1609 VDD.n1211 GND 0.01fF
C1610 VDD.n1212 GND 0.02fF
C1611 VDD.n1213 GND 0.02fF
C1612 VDD.n1214 GND 0.06fF
C1613 VDD.n1215 GND 0.25fF
C1614 VDD.n1216 GND 0.01fF
C1615 VDD.n1217 GND 0.01fF
C1616 VDD.n1218 GND 0.02fF
C1617 VDD.n1219 GND 0.28fF
C1618 VDD.n1220 GND 0.01fF
C1619 VDD.n1221 GND 0.02fF
C1620 VDD.n1222 GND 0.03fF
C1621 VDD.n1223 GND 0.02fF
C1622 VDD.n1224 GND 0.02fF
C1623 VDD.n1225 GND 0.02fF
C1624 VDD.n1226 GND 0.22fF
C1625 VDD.n1227 GND 0.04fF
C1626 VDD.n1228 GND 0.03fF
C1627 VDD.n1229 GND 0.02fF
C1628 VDD.n1230 GND 0.02fF
C1629 VDD.n1231 GND 0.02fF
C1630 VDD.n1232 GND 0.03fF
C1631 VDD.n1233 GND 0.02fF
C1632 VDD.n1235 GND 0.02fF
C1633 VDD.n1236 GND 0.02fF
C1634 VDD.n1237 GND 0.02fF
C1635 VDD.n1239 GND 0.28fF
C1636 VDD.n1241 GND 0.02fF
C1637 VDD.n1242 GND 0.02fF
C1638 VDD.n1243 GND 0.03fF
C1639 VDD.n1244 GND 0.02fF
C1640 VDD.n1245 GND 0.28fF
C1641 VDD.n1246 GND 0.01fF
C1642 VDD.n1247 GND 0.02fF
C1643 VDD.n1248 GND 0.03fF
C1644 VDD.n1249 GND 0.06fF
C1645 VDD.n1250 GND 0.25fF
C1646 VDD.n1251 GND 0.01fF
C1647 VDD.n1252 GND 0.01fF
C1648 VDD.n1253 GND 0.02fF
C1649 VDD.n1254 GND 0.14fF
C1650 VDD.n1255 GND 0.17fF
C1651 VDD.n1256 GND 0.01fF
C1652 VDD.n1257 GND 0.02fF
C1653 VDD.n1258 GND 0.02fF
C1654 VDD.n1259 GND 0.17fF
C1655 VDD.n1260 GND 0.14fF
C1656 VDD.n1261 GND 0.01fF
C1657 VDD.n1262 GND 0.02fF
C1658 VDD.n1263 GND 0.03fF
C1659 VDD.n1264 GND 0.11fF
C1660 VDD.n1265 GND 0.03fF
C1661 VDD.n1266 GND 0.31fF
C1662 VDD.n1267 GND 0.01fF
C1663 VDD.n1268 GND 0.02fF
C1664 VDD.n1269 GND 0.03fF
C1665 VDD.n1270 GND 0.14fF
C1666 VDD.n1271 GND 0.17fF
C1667 VDD.n1272 GND 0.01fF
C1668 VDD.n1273 GND 0.02fF
C1669 VDD.n1274 GND 0.02fF
C1670 VDD.n1275 GND 0.06fF
C1671 VDD.n1276 GND 0.25fF
C1672 VDD.n1277 GND 0.01fF
C1673 VDD.n1278 GND 0.01fF
C1674 VDD.n1279 GND 0.02fF
C1675 VDD.n1280 GND 0.28fF
C1676 VDD.n1281 GND 0.01fF
C1677 VDD.n1282 GND 0.02fF
C1678 VDD.n1283 GND 0.03fF
C1679 VDD.n1284 GND 0.02fF
C1680 VDD.n1285 GND 0.02fF
C1681 VDD.n1286 GND 0.02fF
C1682 VDD.n1287 GND 0.22fF
C1683 VDD.n1288 GND 0.04fF
C1684 VDD.n1289 GND 0.03fF
C1685 VDD.n1290 GND 0.02fF
C1686 VDD.n1291 GND 0.02fF
C1687 VDD.n1292 GND 0.02fF
C1688 VDD.n1293 GND 0.03fF
C1689 VDD.n1294 GND 0.02fF
C1690 VDD.n1296 GND 0.02fF
C1691 VDD.n1297 GND 0.02fF
C1692 VDD.n1298 GND 0.02fF
C1693 VDD.n1300 GND 0.28fF
C1694 VDD.n1302 GND 0.02fF
C1695 VDD.n1303 GND 0.02fF
C1696 VDD.n1304 GND 0.03fF
C1697 VDD.n1305 GND 0.02fF
C1698 VDD.n1306 GND 0.28fF
C1699 VDD.n1307 GND 0.01fF
C1700 VDD.n1308 GND 0.02fF
C1701 VDD.n1309 GND 0.03fF
C1702 VDD.n1310 GND 0.06fF
C1703 VDD.n1311 GND 0.25fF
C1704 VDD.n1312 GND 0.01fF
C1705 VDD.n1313 GND 0.01fF
C1706 VDD.n1314 GND 0.02fF
C1707 VDD.n1315 GND 0.14fF
C1708 VDD.n1316 GND 0.17fF
C1709 VDD.n1317 GND 0.01fF
C1710 VDD.n1318 GND 0.02fF
C1711 VDD.n1319 GND 0.02fF
C1712 VDD.n1320 GND 0.17fF
C1713 VDD.n1321 GND 0.14fF
C1714 VDD.n1322 GND 0.01fF
C1715 VDD.n1323 GND 0.02fF
C1716 VDD.n1324 GND 0.03fF
C1717 VDD.n1325 GND 0.11fF
C1718 VDD.n1326 GND 0.03fF
C1719 VDD.n1327 GND 0.31fF
C1720 VDD.n1328 GND 0.01fF
C1721 VDD.n1329 GND 0.02fF
C1722 VDD.n1330 GND 0.03fF
C1723 VDD.n1331 GND 0.14fF
C1724 VDD.n1332 GND 0.17fF
C1725 VDD.n1333 GND 0.01fF
C1726 VDD.n1334 GND 0.02fF
C1727 VDD.n1335 GND 0.02fF
C1728 VDD.n1336 GND 0.06fF
C1729 VDD.n1337 GND 0.25fF
C1730 VDD.n1338 GND 0.01fF
C1731 VDD.n1339 GND 0.01fF
C1732 VDD.n1340 GND 0.02fF
C1733 VDD.n1341 GND 0.28fF
C1734 VDD.n1342 GND 0.01fF
C1735 VDD.n1343 GND 0.02fF
C1736 VDD.n1344 GND 0.03fF
C1737 VDD.n1345 GND 0.02fF
C1738 VDD.n1346 GND 0.02fF
C1739 VDD.n1347 GND 0.02fF
C1740 VDD.n1348 GND 0.22fF
C1741 VDD.n1349 GND 0.04fF
C1742 VDD.n1350 GND 0.03fF
C1743 VDD.n1351 GND 0.02fF
C1744 VDD.n1352 GND 0.02fF
C1745 VDD.n1353 GND 0.02fF
C1746 VDD.n1354 GND 0.03fF
C1747 VDD.n1355 GND 0.02fF
C1748 VDD.n1357 GND 0.02fF
C1749 VDD.n1358 GND 0.02fF
C1750 VDD.n1359 GND 0.02fF
C1751 VDD.n1361 GND 0.28fF
C1752 VDD.n1363 GND 0.02fF
C1753 VDD.n1364 GND 0.02fF
C1754 VDD.n1365 GND 0.03fF
C1755 VDD.n1366 GND 0.02fF
C1756 VDD.n1367 GND 0.28fF
C1757 VDD.n1368 GND 0.01fF
C1758 VDD.n1369 GND 0.02fF
C1759 VDD.n1370 GND 0.03fF
C1760 VDD.n1371 GND 0.06fF
C1761 VDD.n1372 GND 0.25fF
C1762 VDD.n1373 GND 0.01fF
C1763 VDD.n1374 GND 0.01fF
C1764 VDD.n1375 GND 0.02fF
C1765 VDD.n1376 GND 0.14fF
C1766 VDD.n1377 GND 0.17fF
C1767 VDD.n1378 GND 0.01fF
C1768 VDD.n1379 GND 0.02fF
C1769 VDD.n1380 GND 0.02fF
C1770 VDD.n1381 GND 0.17fF
C1771 VDD.n1382 GND 0.14fF
C1772 VDD.n1383 GND 0.01fF
C1773 VDD.n1384 GND 0.02fF
C1774 VDD.n1385 GND 0.03fF
C1775 VDD.n1386 GND 0.11fF
C1776 VDD.n1387 GND 0.03fF
C1777 VDD.n1388 GND 0.31fF
C1778 VDD.n1389 GND 0.01fF
C1779 VDD.n1390 GND 0.02fF
C1780 VDD.n1391 GND 0.02fF
.ends
