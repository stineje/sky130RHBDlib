* SPICE3 file created from OR2X1.ext - technology: sky130A

.subckt OR2X1 Y A B VPB VNB
X0 a_198_181# a_164_908# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.0774e+12p ps=2.104e+07u w=3e+06u l=150000u
X1 a_851_182# a_198_181# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2 VPB a_198_181# a_851_182# VPB sky130_fd_pr__pfet_01v8 ad=1.68e+12p pd=1.368e+07u as=0p ps=0u w=2e+06u l=150000u M=2
X3 a_131_1005# a_164_908# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X4 a_131_1005# a_343_383# a_198_181# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X5 a_198_181# a_343_383# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
.ends
