* SPICE3 file created from INVX12.ext - technology: sky130A

.subckt INVX12 Y A VSS VDD
X0 Y A.t1 VSS.t0 VSS sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=0p ps=0u w=0u l=0u
X1 Y.t1 A.t0 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 Y A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.1408e+12p ps=8.1e+06u w=3e+06u l=150000u
X3 VDD.t1 A.t2 Y.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
R0 A.n0 A.t2 512.525
R1 A.n0 A.t0 371.139
R2 A.n1 A.t1 282.852
R3 A.n1 A.n0 247.347
R4 A.n2 A.n1 4.65
R5 A.n2 A 0.046
R6 VDD.n35 VDD.t3 135.17
R7 VDD.n24 VDD.t1 135.17
R8 VDD.n47 VDD.n46 92.5
R9 VDD.n45 VDD.n44 92.5
R10 VDD.n43 VDD.n42 92.5
R11 VDD.n41 VDD.n40 92.5
R12 VDD.n49 VDD.n48 92.5
R13 VDD.n14 VDD.n1 92.5
R14 VDD.n5 VDD.n4 92.5
R15 VDD.n7 VDD.n6 92.5
R16 VDD.n9 VDD.n8 92.5
R17 VDD.n11 VDD.n10 92.5
R18 VDD.n13 VDD.n12 92.5
R19 VDD.n21 VDD.n20 92.059
R20 VDD.n58 VDD.n57 92.059
R21 VDD.n20 VDD.n16 67.194
R22 VDD.n20 VDD.n17 67.194
R23 VDD.n20 VDD.n18 67.194
R24 VDD.n20 VDD.n19 67.194
R25 VDD.n5 VDD.n3 44.141
R26 VDD.n3 VDD.n2 44.107
R27 VDD.n25 VDD.t0 43.472
R28 VDD.n33 VDD.t2 43.472
R29 VDD.n20 VDD.n15 41.052
R30 VDD.n56 VDD.n54 39.742
R31 VDD.n56 VDD.n55 39.742
R32 VDD.n53 VDD.n52 39.742
R33 VDD.n1 VDD.n0 30.923
R34 VDD.n57 VDD.n56 26.38
R35 VDD.n57 VDD.n53 26.38
R36 VDD.n57 VDD.n51 26.38
R37 VDD.n57 VDD.n50 26.38
R38 VDD.n60 VDD.n49 22.915
R39 VDD.n23 VDD.n14 22.915
R40 VDD.n49 VDD.n47 14.864
R41 VDD.n47 VDD.n45 14.864
R42 VDD.n45 VDD.n43 14.864
R43 VDD.n43 VDD.n41 14.864
R44 VDD.n41 VDD.n39 14.864
R45 VDD.n39 VDD.n38 14.864
R46 VDD.n14 VDD.n13 14.864
R47 VDD.n13 VDD.n11 14.864
R48 VDD.n11 VDD.n9 14.864
R49 VDD.n9 VDD.n7 14.864
R50 VDD.n7 VDD.n5 14.864
R51 VDD.n23 VDD.n22 8.855
R52 VDD.n22 VDD.n21 8.855
R53 VDD.n27 VDD.n26 8.855
R54 VDD.n26 VDD.n25 8.855
R55 VDD.n31 VDD.n30 8.855
R56 VDD.n30 VDD.n29 8.855
R57 VDD.n36 VDD.n34 8.855
R58 VDD.n34 VDD.n33 8.855
R59 VDD.n60 VDD.n59 8.855
R60 VDD.n59 VDD.n58 8.855
R61 VDD.n28 VDD.n23 4.795
R62 VDD.n28 VDD.n27 4.65
R63 VDD.n32 VDD.n31 4.65
R64 VDD.n37 VDD.n36 4.65
R65 VDD.n61 VDD.n60 4.65
R66 VDD.n27 VDD.n24 2.064
R67 VDD.n36 VDD.n35 2.064
R68 VDD.n32 VDD.n28 0.157
R69 VDD.n37 VDD.n32 0.157
R70 VDD.n61 VDD.n37 0.145
R71 VDD.n61 VDD 0.034
R72 Y.n5 Y.n4 272.451
R73 Y.n5 Y.n0 271.281
R74 Y.n4 Y.n3 30
R75 Y.n2 Y.n1 24.383
R76 Y.n4 Y.n2 23.684
R77 Y.n0 Y.t0 14.282
R78 Y.n0 Y.t1 14.282
R79 Y.n6 Y.n5 4.65
R80 Y.n6 Y 0.046
R81 VSS.n21 VSS.n20 37.582
R82 VSS.t0 VSS.n18 32.601
R83 VSS.n18 VSS.n17 21.734
R84 VSS.n4 VSS.n3 20.705
R85 VSS.n10 VSS.n9 20.705
R86 VSS.n22 VSS.n21 20.705
R87 VSS.n3 VSS.n2 19.952
R88 VSS.n20 VSS.t0 15.644
R89 VSS.n20 VSS.n19 13.541
R90 VSS.n23 VSS.n14 9.154
R91 VSS.n12 VSS.n11 9.154
R92 VSS.n6 VSS.n5 9.154
R93 VSS.n7 VSS.n1 4.795
R94 VSS.n27 VSS.n26 4.65
R95 VSS.n7 VSS.n6 4.65
R96 VSS.n13 VSS.n12 4.65
R97 VSS.n24 VSS.n23 4.65
R98 VSS.n16 VSS.n15 4.504
R99 VSS.n6 VSS.n4 4.129
R100 VSS.n23 VSS.n22 3.716
R101 VSS.t0 VSS.n16 2.452
R102 VSS.n1 VSS.n0 0.474
R103 VSS.n26 VSS.n25 0.474
R104 VSS.n9 VSS.n8 0.376
R105 VSS.n12 VSS.n10 0.206
R106 VSS.n13 VSS.n7 0.157
R107 VSS.n24 VSS.n13 0.157
R108 VSS.n27 VSS.n24 0.145
R109 VSS.n27 VSS 0.034
.ends
