// File: nmos_bottom.spi.pex
// Created: Tue Oct 15 15:58:05 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
