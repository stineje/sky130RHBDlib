* SPICE3 file created from MUX2X1.ext - technology: sky130A

.subckt MUX2X1 Y A0 A1 S VDD GND
X0 a_661_1004 A0 VDD VDD pshort w=2 l=0.15 M=2
X1 VDD A1 a_1327_1004 VDD pshort w=2 l=0.15 M=2
X2 a_185_182 S GND GND nshort w=3 l=0.15
X3 a_661_1004 A0 a_556_73 GND nshort w=3 l=0.15
X4 a_661_1004 S VDD VDD pshort w=2 l=0.15 M=2
X5 VDD S a_185_182 VDD pshort w=2 l=0.15 M=2
X6 a_1327_1004 a_185_182 VDD VDD pshort w=2 l=0.15 M=2
X7 VDD a_1327_1004 Y VDD pshort w=2 l=0.15 M=2
X8 VDD a_661_1004 Y VDD pshort w=2 l=0.15 M=2
X9 GND a_661_1004 a_1888_73 GND nshort w=3 l=0.15
X10 GND a_185_182 a_1222_73 GND nshort w=3 l=0.15
X11 Y a_1327_1004 a_1888_73 GND nshort w=3 l=0.15
X12 GND S a_556_73 GND nshort w=3 l=0.15
X13 a_1327_1004 A1 a_1222_73 GND nshort w=3 l=0.15
C0 VDD GND 6.15fF
.ends
