* SPICE3 file created from TIEHI.ext - technology: sky130A

.subckt TIEHI Y VDD GND
X0 a_155_381# a_155_381# GND GND nshort w=3 l=0.15
X1 VDD a_155_381# Y VDD pshort w=2 l=0.15
.ends
