magic
tech sky130A
magscale 1 2
timestamp 1669564295
<< nwell >>
rect -87 786 7857 1550
<< pwell >>
rect -34 -34 7804 544
<< nmos >>
rect 155 297 185 350
tri 185 297 201 313 sw
rect 155 267 261 297
tri 261 267 291 297 sw
rect 155 166 185 267
tri 185 251 201 267 nw
tri 245 251 261 267 ne
tri 185 166 201 182 sw
tri 245 166 261 182 se
rect 261 166 291 267
tri 155 136 185 166 ne
rect 185 136 261 166
tri 261 136 291 166 nw
rect 612 289 642 350
tri 642 289 658 305 sw
rect 806 297 836 350
tri 836 297 852 313 sw
rect 612 259 718 289
tri 718 259 748 289 sw
rect 806 267 912 297
tri 912 267 942 297 sw
rect 612 158 642 259
tri 642 243 658 259 nw
tri 702 243 718 259 ne
tri 642 158 658 174 sw
tri 702 158 718 174 se
rect 718 158 748 259
rect 806 166 836 267
tri 836 251 852 267 nw
tri 896 251 912 267 ne
tri 836 166 852 182 sw
tri 896 166 912 182 se
rect 912 166 942 267
tri 612 128 642 158 ne
rect 642 128 718 158
tri 718 128 748 158 nw
tri 806 136 836 166 ne
rect 836 136 912 166
tri 912 136 942 166 nw
rect 1278 289 1308 350
tri 1308 289 1324 305 sw
rect 1472 297 1502 350
tri 1502 297 1518 313 sw
rect 1278 259 1384 289
tri 1384 259 1414 289 sw
rect 1472 267 1578 297
tri 1578 267 1608 297 sw
rect 1278 158 1308 259
tri 1308 243 1324 259 nw
tri 1368 243 1384 259 ne
tri 1308 158 1324 174 sw
tri 1368 158 1384 174 se
rect 1384 158 1414 259
rect 1472 166 1502 267
tri 1502 251 1518 267 nw
tri 1562 251 1578 267 ne
tri 1502 166 1518 182 sw
tri 1562 166 1578 182 se
rect 1578 166 1608 267
tri 1278 128 1308 158 ne
rect 1308 128 1384 158
tri 1384 128 1414 158 nw
tri 1472 136 1502 166 ne
rect 1502 136 1578 166
tri 1578 136 1608 166 nw
tri 2019 297 2035 313 se
rect 2035 297 2065 350
tri 1929 267 1959 297 se
rect 1959 267 2065 297
rect 1929 166 1959 267
tri 1959 251 1975 267 nw
tri 2019 251 2035 267 ne
tri 1959 166 1975 182 sw
tri 2019 166 2035 182 se
rect 2035 166 2065 267
tri 1929 136 1959 166 ne
rect 1959 136 2035 166
tri 2035 136 2065 166 nw
rect 2375 297 2405 350
tri 2405 297 2421 313 sw
rect 2375 267 2481 297
tri 2481 267 2511 297 sw
rect 2375 166 2405 267
tri 2405 251 2421 267 nw
tri 2465 251 2481 267 ne
tri 2405 166 2421 182 sw
tri 2465 166 2481 182 se
rect 2481 166 2511 267
tri 2375 136 2405 166 ne
rect 2405 136 2481 166
tri 2481 136 2511 166 nw
rect 2832 289 2862 350
tri 2862 289 2878 305 sw
rect 3026 297 3056 350
tri 3056 297 3072 313 sw
rect 2832 259 2938 289
tri 2938 259 2968 289 sw
rect 3026 267 3132 297
tri 3132 267 3162 297 sw
rect 2832 158 2862 259
tri 2862 243 2878 259 nw
tri 2922 243 2938 259 ne
tri 2862 158 2878 174 sw
tri 2922 158 2938 174 se
rect 2938 158 2968 259
rect 3026 166 3056 267
tri 3056 251 3072 267 nw
tri 3116 251 3132 267 ne
tri 3056 166 3072 182 sw
tri 3116 166 3132 182 se
rect 3132 166 3162 267
tri 2832 128 2862 158 ne
rect 2862 128 2938 158
tri 2938 128 2968 158 nw
tri 3026 136 3056 166 ne
rect 3056 136 3132 166
tri 3132 136 3162 166 nw
rect 3498 289 3528 350
tri 3528 289 3544 305 sw
rect 3692 297 3722 350
tri 3722 297 3738 313 sw
rect 3498 259 3604 289
tri 3604 259 3634 289 sw
rect 3692 267 3798 297
tri 3798 267 3828 297 sw
rect 3498 158 3528 259
tri 3528 243 3544 259 nw
tri 3588 243 3604 259 ne
tri 3528 158 3544 174 sw
tri 3588 158 3604 174 se
rect 3604 158 3634 259
rect 3692 166 3722 267
tri 3722 251 3738 267 nw
tri 3782 251 3798 267 ne
tri 3722 166 3738 182 sw
tri 3782 166 3798 182 se
rect 3798 166 3828 267
tri 3498 128 3528 158 ne
rect 3528 128 3604 158
tri 3604 128 3634 158 nw
tri 3692 136 3722 166 ne
rect 3722 136 3798 166
tri 3798 136 3828 166 nw
tri 4239 297 4255 313 se
rect 4255 297 4285 350
tri 4149 267 4179 297 se
rect 4179 267 4285 297
rect 4149 166 4179 267
tri 4179 251 4195 267 nw
tri 4239 251 4255 267 ne
tri 4179 166 4195 182 sw
tri 4239 166 4255 182 se
rect 4255 166 4285 267
tri 4149 136 4179 166 ne
rect 4179 136 4255 166
tri 4255 136 4285 166 nw
rect 4608 288 4638 349
tri 4638 288 4654 304 sw
rect 4802 296 4832 349
tri 4832 296 4848 312 sw
rect 4608 258 4714 288
tri 4714 258 4744 288 sw
rect 4802 266 4908 296
tri 4908 266 4938 296 sw
rect 4608 157 4638 258
tri 4638 242 4654 258 nw
tri 4698 242 4714 258 ne
tri 4638 157 4654 173 sw
tri 4698 157 4714 173 se
rect 4714 157 4744 258
rect 4802 165 4832 266
tri 4832 250 4848 266 nw
tri 4892 250 4908 266 ne
tri 4832 165 4848 181 sw
tri 4892 165 4908 181 se
rect 4908 165 4938 266
tri 4608 127 4638 157 ne
rect 4638 127 4714 157
tri 4714 127 4744 157 nw
tri 4802 135 4832 165 ne
rect 4832 135 4908 165
tri 4908 135 4938 165 nw
rect 5261 297 5291 350
tri 5291 297 5307 313 sw
rect 5261 267 5367 297
tri 5367 267 5397 297 sw
rect 5261 166 5291 267
tri 5291 251 5307 267 nw
tri 5351 251 5367 267 ne
tri 5291 166 5307 182 sw
tri 5351 166 5367 182 se
rect 5367 166 5397 267
tri 5261 136 5291 166 ne
rect 5291 136 5367 166
tri 5367 136 5397 166 nw
rect 5718 288 5748 349
tri 5748 288 5764 304 sw
rect 5912 296 5942 349
tri 5942 296 5958 312 sw
rect 5718 258 5824 288
tri 5824 258 5854 288 sw
rect 5912 266 6018 296
tri 6018 266 6048 296 sw
rect 5718 157 5748 258
tri 5748 242 5764 258 nw
tri 5808 242 5824 258 ne
tri 5748 157 5764 173 sw
tri 5808 157 5824 173 se
rect 5824 157 5854 258
rect 5912 165 5942 266
tri 5942 250 5958 266 nw
tri 6002 250 6018 266 ne
tri 5942 165 5958 181 sw
tri 6002 165 6018 181 se
rect 6018 165 6048 266
tri 5718 127 5748 157 ne
rect 5748 127 5824 157
tri 5824 127 5854 157 nw
tri 5912 135 5942 165 ne
rect 5942 135 6018 165
tri 6018 135 6048 165 nw
rect 6371 297 6401 350
tri 6401 297 6417 313 sw
rect 6371 267 6477 297
tri 6477 267 6507 297 sw
rect 6371 166 6401 267
tri 6401 251 6417 267 nw
tri 6461 251 6477 267 ne
tri 6401 166 6417 182 sw
tri 6461 166 6477 182 se
rect 6477 166 6507 267
tri 6371 136 6401 166 ne
rect 6401 136 6477 166
tri 6477 136 6507 166 nw
rect 6828 296 6858 349
tri 6858 296 6874 312 sw
rect 7022 296 7052 349
tri 7052 296 7068 312 sw
rect 6828 266 6934 296
tri 6934 266 6964 296 sw
rect 6828 165 6858 266
tri 6858 250 6874 266 nw
tri 6918 250 6934 266 ne
tri 6858 165 6874 181 sw
tri 6918 165 6934 181 se
rect 6934 165 6964 266
rect 7022 266 7128 296
tri 7128 266 7158 296 sw
rect 7022 251 7053 266
tri 7053 251 7068 266 nw
tri 7112 251 7127 266 ne
rect 7127 251 7158 266
tri 6828 135 6858 165 ne
rect 6858 135 6934 165
tri 6934 135 6964 165 nw
rect 7022 165 7052 251
tri 7052 165 7068 181 sw
tri 7112 165 7128 181 se
rect 7128 165 7158 251
tri 7022 135 7052 165 ne
rect 7052 135 7128 165
tri 7128 135 7158 165 nw
rect 7481 297 7511 350
tri 7511 297 7527 313 sw
rect 7481 267 7587 297
tri 7587 267 7617 297 sw
rect 7481 166 7511 267
tri 7511 251 7527 267 nw
tri 7571 251 7587 267 ne
tri 7511 166 7527 182 sw
tri 7571 166 7587 182 se
rect 7587 166 7617 267
tri 7481 136 7511 166 ne
rect 7511 136 7587 166
tri 7587 136 7617 166 nw
<< pmos >>
rect 164 1004 194 1404
rect 252 1004 282 1404
rect 631 1004 661 1404
rect 719 1004 749 1404
rect 807 1004 837 1404
rect 895 1004 925 1404
rect 1297 1004 1327 1404
rect 1385 1004 1415 1404
rect 1473 1004 1503 1404
rect 1561 1004 1591 1404
rect 1938 1004 1968 1404
rect 2026 1004 2056 1404
rect 2384 1004 2414 1404
rect 2472 1004 2502 1404
rect 2851 1004 2881 1404
rect 2939 1004 2969 1404
rect 3027 1004 3057 1404
rect 3115 1004 3145 1404
rect 3517 1004 3547 1404
rect 3605 1004 3635 1404
rect 3693 1004 3723 1404
rect 3781 1004 3811 1404
rect 4158 1004 4188 1404
rect 4246 1004 4276 1404
rect 4627 1004 4657 1404
rect 4715 1004 4745 1404
rect 4803 1004 4833 1404
rect 4891 1004 4921 1404
rect 5270 1004 5300 1404
rect 5358 1004 5388 1404
rect 5737 1004 5767 1404
rect 5825 1004 5855 1404
rect 5913 1004 5943 1404
rect 6001 1004 6031 1404
rect 6380 1004 6410 1404
rect 6468 1004 6498 1404
rect 6847 1005 6877 1405
rect 6935 1005 6965 1405
rect 7023 1005 7053 1405
rect 7111 1005 7141 1405
rect 7490 1004 7520 1404
rect 7578 1004 7608 1404
<< ndiff >>
rect 99 334 155 350
rect 99 300 109 334
rect 143 300 155 334
rect 99 262 155 300
rect 185 334 345 350
rect 185 313 303 334
tri 185 297 201 313 ne
rect 201 300 303 313
rect 337 300 345 334
rect 201 297 345 300
tri 261 267 291 297 ne
rect 99 228 109 262
rect 143 228 155 262
rect 99 194 155 228
rect 99 160 109 194
rect 143 160 155 194
tri 185 251 201 267 se
rect 201 251 245 267
tri 245 251 261 267 sw
rect 185 218 261 251
rect 185 184 205 218
rect 239 184 261 218
rect 185 182 261 184
tri 185 166 201 182 ne
rect 201 166 245 182
tri 245 166 261 182 nw
rect 291 262 345 297
rect 291 228 303 262
rect 337 228 345 262
rect 291 194 345 228
rect 99 136 155 160
tri 155 136 185 166 sw
tri 261 136 291 166 se
rect 291 160 303 194
rect 337 160 345 194
rect 291 136 345 160
rect 99 124 345 136
rect 99 90 109 124
rect 143 90 205 124
rect 239 90 303 124
rect 337 90 345 124
rect 99 74 345 90
rect 556 334 612 350
rect 556 300 566 334
rect 600 300 612 334
rect 556 262 612 300
rect 642 334 806 350
rect 642 305 663 334
tri 642 289 658 305 ne
rect 658 300 663 305
rect 697 300 760 334
rect 794 300 806 334
rect 658 289 806 300
rect 836 313 998 350
tri 836 297 852 313 ne
rect 852 297 998 313
rect 556 228 566 262
rect 600 228 612 262
tri 718 259 748 289 ne
rect 748 262 806 289
tri 912 267 942 297 ne
rect 556 194 612 228
rect 556 160 566 194
rect 600 160 612 194
rect 556 128 612 160
tri 642 243 658 259 se
rect 658 243 702 259
tri 702 243 718 259 sw
rect 642 209 718 243
rect 642 175 663 209
rect 697 175 718 209
rect 642 174 718 175
tri 642 158 658 174 ne
rect 658 158 702 174
tri 702 158 718 174 nw
rect 748 228 760 262
rect 794 228 806 262
rect 748 194 806 228
rect 748 160 760 194
rect 794 160 806 194
tri 836 251 852 267 se
rect 852 251 896 267
tri 896 251 912 267 sw
rect 836 218 912 251
rect 836 184 857 218
rect 891 184 912 218
rect 836 182 912 184
tri 836 166 852 182 ne
rect 852 166 896 182
tri 896 166 912 182 nw
rect 942 262 998 297
rect 942 228 954 262
rect 988 228 998 262
rect 942 194 998 228
tri 612 128 642 158 sw
tri 718 128 748 158 se
rect 748 136 806 160
tri 806 136 836 166 sw
tri 912 136 942 166 se
rect 942 160 954 194
rect 988 160 998 194
rect 942 136 998 160
rect 748 128 998 136
rect 556 124 998 128
rect 556 90 566 124
rect 600 90 760 124
rect 794 90 857 124
rect 891 90 954 124
rect 988 90 998 124
rect 556 74 998 90
rect 1222 334 1278 350
rect 1222 300 1232 334
rect 1266 300 1278 334
rect 1222 262 1278 300
rect 1308 334 1472 350
rect 1308 305 1329 334
tri 1308 289 1324 305 ne
rect 1324 300 1329 305
rect 1363 300 1426 334
rect 1460 300 1472 334
rect 1324 289 1472 300
rect 1502 313 1664 350
tri 1502 297 1518 313 ne
rect 1518 297 1664 313
rect 1222 228 1232 262
rect 1266 228 1278 262
tri 1384 259 1414 289 ne
rect 1414 262 1472 289
tri 1578 267 1608 297 ne
rect 1222 194 1278 228
rect 1222 160 1232 194
rect 1266 160 1278 194
rect 1222 128 1278 160
tri 1308 243 1324 259 se
rect 1324 243 1368 259
tri 1368 243 1384 259 sw
rect 1308 209 1384 243
rect 1308 175 1329 209
rect 1363 175 1384 209
rect 1308 174 1384 175
tri 1308 158 1324 174 ne
rect 1324 158 1368 174
tri 1368 158 1384 174 nw
rect 1414 228 1426 262
rect 1460 228 1472 262
rect 1414 194 1472 228
rect 1414 160 1426 194
rect 1460 160 1472 194
tri 1502 251 1518 267 se
rect 1518 251 1562 267
tri 1562 251 1578 267 sw
rect 1502 218 1578 251
rect 1502 184 1523 218
rect 1557 184 1578 218
rect 1502 182 1578 184
tri 1502 166 1518 182 ne
rect 1518 166 1562 182
tri 1562 166 1578 182 nw
rect 1608 262 1664 297
rect 1608 228 1620 262
rect 1654 228 1664 262
rect 1608 194 1664 228
tri 1278 128 1308 158 sw
tri 1384 128 1414 158 se
rect 1414 136 1472 160
tri 1472 136 1502 166 sw
tri 1578 136 1608 166 se
rect 1608 160 1620 194
rect 1654 160 1664 194
rect 1608 136 1664 160
rect 1414 128 1664 136
rect 1222 124 1664 128
rect 1222 90 1232 124
rect 1266 90 1426 124
rect 1460 90 1523 124
rect 1557 90 1620 124
rect 1654 90 1664 124
rect 1222 74 1664 90
rect 1875 334 2035 350
rect 1875 300 1883 334
rect 1917 313 2035 334
rect 1917 300 2019 313
rect 1875 297 2019 300
tri 2019 297 2035 313 nw
rect 2065 334 2121 350
rect 2065 300 2077 334
rect 2111 300 2121 334
rect 1875 262 1929 297
tri 1929 267 1959 297 nw
rect 1875 228 1883 262
rect 1917 228 1929 262
rect 1875 194 1929 228
rect 1875 160 1883 194
rect 1917 160 1929 194
tri 1959 251 1975 267 se
rect 1975 251 2019 267
tri 2019 251 2035 267 sw
rect 1959 218 2035 251
rect 1959 184 1981 218
rect 2015 184 2035 218
rect 1959 182 2035 184
tri 1959 166 1975 182 ne
rect 1975 166 2019 182
tri 2019 166 2035 182 nw
rect 2065 262 2121 300
rect 2065 228 2077 262
rect 2111 228 2121 262
rect 2065 194 2121 228
rect 1875 136 1929 160
tri 1929 136 1959 166 sw
tri 2035 136 2065 166 se
rect 2065 160 2077 194
rect 2111 160 2121 194
rect 2065 136 2121 160
rect 1875 124 2121 136
rect 1875 90 1883 124
rect 1917 90 1981 124
rect 2015 90 2077 124
rect 2111 90 2121 124
rect 1875 74 2121 90
rect 2319 334 2375 350
rect 2319 300 2329 334
rect 2363 300 2375 334
rect 2319 262 2375 300
rect 2405 334 2565 350
rect 2405 313 2523 334
tri 2405 297 2421 313 ne
rect 2421 300 2523 313
rect 2557 300 2565 334
rect 2421 297 2565 300
tri 2481 267 2511 297 ne
rect 2319 228 2329 262
rect 2363 228 2375 262
rect 2319 194 2375 228
rect 2319 160 2329 194
rect 2363 160 2375 194
tri 2405 251 2421 267 se
rect 2421 251 2465 267
tri 2465 251 2481 267 sw
rect 2405 218 2481 251
rect 2405 184 2425 218
rect 2459 184 2481 218
rect 2405 182 2481 184
tri 2405 166 2421 182 ne
rect 2421 166 2465 182
tri 2465 166 2481 182 nw
rect 2511 262 2565 297
rect 2511 228 2523 262
rect 2557 228 2565 262
rect 2511 194 2565 228
rect 2319 136 2375 160
tri 2375 136 2405 166 sw
tri 2481 136 2511 166 se
rect 2511 160 2523 194
rect 2557 160 2565 194
rect 2511 136 2565 160
rect 2319 124 2565 136
rect 2319 90 2329 124
rect 2363 90 2425 124
rect 2459 90 2523 124
rect 2557 90 2565 124
rect 2319 74 2565 90
rect 2776 334 2832 350
rect 2776 300 2786 334
rect 2820 300 2832 334
rect 2776 262 2832 300
rect 2862 334 3026 350
rect 2862 305 2883 334
tri 2862 289 2878 305 ne
rect 2878 300 2883 305
rect 2917 300 2980 334
rect 3014 300 3026 334
rect 2878 289 3026 300
rect 3056 313 3218 350
tri 3056 297 3072 313 ne
rect 3072 297 3218 313
rect 2776 228 2786 262
rect 2820 228 2832 262
tri 2938 259 2968 289 ne
rect 2968 262 3026 289
tri 3132 267 3162 297 ne
rect 2776 194 2832 228
rect 2776 160 2786 194
rect 2820 160 2832 194
rect 2776 128 2832 160
tri 2862 243 2878 259 se
rect 2878 243 2922 259
tri 2922 243 2938 259 sw
rect 2862 209 2938 243
rect 2862 175 2883 209
rect 2917 175 2938 209
rect 2862 174 2938 175
tri 2862 158 2878 174 ne
rect 2878 158 2922 174
tri 2922 158 2938 174 nw
rect 2968 228 2980 262
rect 3014 228 3026 262
rect 2968 194 3026 228
rect 2968 160 2980 194
rect 3014 160 3026 194
tri 3056 251 3072 267 se
rect 3072 251 3116 267
tri 3116 251 3132 267 sw
rect 3056 218 3132 251
rect 3056 184 3077 218
rect 3111 184 3132 218
rect 3056 182 3132 184
tri 3056 166 3072 182 ne
rect 3072 166 3116 182
tri 3116 166 3132 182 nw
rect 3162 262 3218 297
rect 3162 228 3174 262
rect 3208 228 3218 262
rect 3162 194 3218 228
tri 2832 128 2862 158 sw
tri 2938 128 2968 158 se
rect 2968 136 3026 160
tri 3026 136 3056 166 sw
tri 3132 136 3162 166 se
rect 3162 160 3174 194
rect 3208 160 3218 194
rect 3162 136 3218 160
rect 2968 128 3218 136
rect 2776 124 3218 128
rect 2776 90 2786 124
rect 2820 90 2980 124
rect 3014 90 3077 124
rect 3111 90 3174 124
rect 3208 90 3218 124
rect 2776 74 3218 90
rect 3442 334 3498 350
rect 3442 300 3452 334
rect 3486 300 3498 334
rect 3442 262 3498 300
rect 3528 334 3692 350
rect 3528 305 3549 334
tri 3528 289 3544 305 ne
rect 3544 300 3549 305
rect 3583 300 3646 334
rect 3680 300 3692 334
rect 3544 289 3692 300
rect 3722 313 3884 350
tri 3722 297 3738 313 ne
rect 3738 297 3884 313
rect 3442 228 3452 262
rect 3486 228 3498 262
tri 3604 259 3634 289 ne
rect 3634 262 3692 289
tri 3798 267 3828 297 ne
rect 3442 194 3498 228
rect 3442 160 3452 194
rect 3486 160 3498 194
rect 3442 128 3498 160
tri 3528 243 3544 259 se
rect 3544 243 3588 259
tri 3588 243 3604 259 sw
rect 3528 209 3604 243
rect 3528 175 3549 209
rect 3583 175 3604 209
rect 3528 174 3604 175
tri 3528 158 3544 174 ne
rect 3544 158 3588 174
tri 3588 158 3604 174 nw
rect 3634 228 3646 262
rect 3680 228 3692 262
rect 3634 194 3692 228
rect 3634 160 3646 194
rect 3680 160 3692 194
tri 3722 251 3738 267 se
rect 3738 251 3782 267
tri 3782 251 3798 267 sw
rect 3722 218 3798 251
rect 3722 184 3743 218
rect 3777 184 3798 218
rect 3722 182 3798 184
tri 3722 166 3738 182 ne
rect 3738 166 3782 182
tri 3782 166 3798 182 nw
rect 3828 262 3884 297
rect 3828 228 3840 262
rect 3874 228 3884 262
rect 3828 194 3884 228
tri 3498 128 3528 158 sw
tri 3604 128 3634 158 se
rect 3634 136 3692 160
tri 3692 136 3722 166 sw
tri 3798 136 3828 166 se
rect 3828 160 3840 194
rect 3874 160 3884 194
rect 3828 136 3884 160
rect 3634 128 3884 136
rect 3442 124 3884 128
rect 3442 90 3452 124
rect 3486 90 3646 124
rect 3680 90 3743 124
rect 3777 90 3840 124
rect 3874 90 3884 124
rect 3442 74 3884 90
rect 4095 334 4255 350
rect 4095 300 4103 334
rect 4137 313 4255 334
rect 4137 300 4239 313
rect 4095 297 4239 300
tri 4239 297 4255 313 nw
rect 4285 334 4341 350
rect 4285 300 4297 334
rect 4331 300 4341 334
rect 4095 262 4149 297
tri 4149 267 4179 297 nw
rect 4095 228 4103 262
rect 4137 228 4149 262
rect 4095 194 4149 228
rect 4095 160 4103 194
rect 4137 160 4149 194
tri 4179 251 4195 267 se
rect 4195 251 4239 267
tri 4239 251 4255 267 sw
rect 4179 218 4255 251
rect 4179 184 4201 218
rect 4235 184 4255 218
rect 4179 182 4255 184
tri 4179 166 4195 182 ne
rect 4195 166 4239 182
tri 4239 166 4255 182 nw
rect 4285 262 4341 300
rect 4285 228 4297 262
rect 4331 228 4341 262
rect 4285 194 4341 228
rect 4095 136 4149 160
tri 4149 136 4179 166 sw
tri 4255 136 4285 166 se
rect 4285 160 4297 194
rect 4331 160 4341 194
rect 4285 136 4341 160
rect 4095 124 4341 136
rect 4095 90 4103 124
rect 4137 90 4201 124
rect 4235 90 4297 124
rect 4331 90 4341 124
rect 4095 74 4341 90
rect 4552 333 4608 349
rect 4552 299 4562 333
rect 4596 299 4608 333
rect 4552 261 4608 299
rect 4638 333 4802 349
rect 4638 304 4659 333
tri 4638 288 4654 304 ne
rect 4654 299 4659 304
rect 4693 299 4756 333
rect 4790 299 4802 333
rect 4654 288 4802 299
rect 4832 312 4994 349
tri 4832 296 4848 312 ne
rect 4848 296 4994 312
rect 4552 227 4562 261
rect 4596 227 4608 261
tri 4714 258 4744 288 ne
rect 4744 261 4802 288
tri 4908 266 4938 296 ne
rect 4552 193 4608 227
rect 4552 159 4562 193
rect 4596 159 4608 193
rect 4552 127 4608 159
tri 4638 242 4654 258 se
rect 4654 242 4698 258
tri 4698 242 4714 258 sw
rect 4638 208 4714 242
rect 4638 174 4659 208
rect 4693 174 4714 208
rect 4638 173 4714 174
tri 4638 157 4654 173 ne
rect 4654 157 4698 173
tri 4698 157 4714 173 nw
rect 4744 227 4756 261
rect 4790 227 4802 261
rect 4744 193 4802 227
rect 4744 159 4756 193
rect 4790 159 4802 193
tri 4832 250 4848 266 se
rect 4848 250 4892 266
tri 4892 250 4908 266 sw
rect 4832 217 4908 250
rect 4832 183 4853 217
rect 4887 183 4908 217
rect 4832 181 4908 183
tri 4832 165 4848 181 ne
rect 4848 165 4892 181
tri 4892 165 4908 181 nw
rect 4938 261 4994 296
rect 4938 227 4950 261
rect 4984 227 4994 261
rect 4938 193 4994 227
tri 4608 127 4638 157 sw
tri 4714 127 4744 157 se
rect 4744 135 4802 159
tri 4802 135 4832 165 sw
tri 4908 135 4938 165 se
rect 4938 159 4950 193
rect 4984 159 4994 193
rect 4938 135 4994 159
rect 4744 127 4994 135
rect 4552 123 4994 127
rect 4552 89 4562 123
rect 4596 89 4756 123
rect 4790 89 4853 123
rect 4887 89 4950 123
rect 4984 89 4994 123
rect 4552 73 4994 89
rect 5205 334 5261 350
rect 5205 300 5215 334
rect 5249 300 5261 334
rect 5205 262 5261 300
rect 5291 334 5451 350
rect 5291 313 5409 334
tri 5291 297 5307 313 ne
rect 5307 300 5409 313
rect 5443 300 5451 334
rect 5307 297 5451 300
tri 5367 267 5397 297 ne
rect 5205 228 5215 262
rect 5249 228 5261 262
rect 5205 194 5261 228
rect 5205 160 5215 194
rect 5249 160 5261 194
tri 5291 251 5307 267 se
rect 5307 251 5351 267
tri 5351 251 5367 267 sw
rect 5291 218 5367 251
rect 5291 184 5311 218
rect 5345 184 5367 218
rect 5291 182 5367 184
tri 5291 166 5307 182 ne
rect 5307 166 5351 182
tri 5351 166 5367 182 nw
rect 5397 262 5451 297
rect 5397 228 5409 262
rect 5443 228 5451 262
rect 5397 194 5451 228
rect 5205 136 5261 160
tri 5261 136 5291 166 sw
tri 5367 136 5397 166 se
rect 5397 160 5409 194
rect 5443 160 5451 194
rect 5397 136 5451 160
rect 5205 124 5451 136
rect 5205 90 5215 124
rect 5249 90 5311 124
rect 5345 90 5409 124
rect 5443 90 5451 124
rect 5205 74 5451 90
rect 5662 333 5718 349
rect 5662 299 5672 333
rect 5706 299 5718 333
rect 5662 261 5718 299
rect 5748 333 5912 349
rect 5748 304 5769 333
tri 5748 288 5764 304 ne
rect 5764 299 5769 304
rect 5803 299 5866 333
rect 5900 299 5912 333
rect 5764 288 5912 299
rect 5942 312 6104 349
tri 5942 296 5958 312 ne
rect 5958 296 6104 312
rect 5662 227 5672 261
rect 5706 227 5718 261
tri 5824 258 5854 288 ne
rect 5854 261 5912 288
tri 6018 266 6048 296 ne
rect 5662 193 5718 227
rect 5662 159 5672 193
rect 5706 159 5718 193
rect 5662 127 5718 159
tri 5748 242 5764 258 se
rect 5764 242 5808 258
tri 5808 242 5824 258 sw
rect 5748 208 5824 242
rect 5748 174 5769 208
rect 5803 174 5824 208
rect 5748 173 5824 174
tri 5748 157 5764 173 ne
rect 5764 157 5808 173
tri 5808 157 5824 173 nw
rect 5854 227 5866 261
rect 5900 227 5912 261
rect 5854 193 5912 227
rect 5854 159 5866 193
rect 5900 159 5912 193
tri 5942 250 5958 266 se
rect 5958 250 6002 266
tri 6002 250 6018 266 sw
rect 5942 217 6018 250
rect 5942 183 5963 217
rect 5997 183 6018 217
rect 5942 181 6018 183
tri 5942 165 5958 181 ne
rect 5958 165 6002 181
tri 6002 165 6018 181 nw
rect 6048 261 6104 296
rect 6048 227 6060 261
rect 6094 227 6104 261
rect 6048 193 6104 227
tri 5718 127 5748 157 sw
tri 5824 127 5854 157 se
rect 5854 135 5912 159
tri 5912 135 5942 165 sw
tri 6018 135 6048 165 se
rect 6048 159 6060 193
rect 6094 159 6104 193
rect 6048 135 6104 159
rect 5854 127 6104 135
rect 5662 123 6104 127
rect 5662 89 5672 123
rect 5706 89 5866 123
rect 5900 89 5963 123
rect 5997 89 6060 123
rect 6094 89 6104 123
rect 5662 73 6104 89
rect 6315 334 6371 350
rect 6315 300 6325 334
rect 6359 300 6371 334
rect 6315 262 6371 300
rect 6401 334 6561 350
rect 6401 313 6519 334
tri 6401 297 6417 313 ne
rect 6417 300 6519 313
rect 6553 300 6561 334
rect 6417 297 6561 300
tri 6477 267 6507 297 ne
rect 6315 228 6325 262
rect 6359 228 6371 262
rect 6315 194 6371 228
rect 6315 160 6325 194
rect 6359 160 6371 194
tri 6401 251 6417 267 se
rect 6417 251 6461 267
tri 6461 251 6477 267 sw
rect 6401 218 6477 251
rect 6401 184 6421 218
rect 6455 184 6477 218
rect 6401 182 6477 184
tri 6401 166 6417 182 ne
rect 6417 166 6461 182
tri 6461 166 6477 182 nw
rect 6507 262 6561 297
rect 6507 228 6519 262
rect 6553 228 6561 262
rect 6507 194 6561 228
rect 6315 136 6371 160
tri 6371 136 6401 166 sw
tri 6477 136 6507 166 se
rect 6507 160 6519 194
rect 6553 160 6561 194
rect 6507 136 6561 160
rect 6315 124 6561 136
rect 6315 90 6325 124
rect 6359 90 6421 124
rect 6455 90 6519 124
rect 6553 90 6561 124
rect 6315 74 6561 90
rect 6772 333 6828 349
rect 6772 299 6782 333
rect 6816 299 6828 333
rect 6772 261 6828 299
rect 6858 312 7022 349
tri 6858 296 6874 312 ne
rect 6874 296 7022 312
rect 7052 312 7214 349
tri 7052 296 7068 312 ne
rect 7068 296 7214 312
tri 6934 266 6964 296 ne
rect 6772 227 6782 261
rect 6816 227 6828 261
rect 6772 193 6828 227
rect 6772 159 6782 193
rect 6816 159 6828 193
tri 6858 250 6874 266 se
rect 6874 250 6918 266
tri 6918 250 6934 266 sw
rect 6858 217 6934 250
rect 6858 183 6879 217
rect 6913 183 6934 217
rect 6858 181 6934 183
tri 6858 165 6874 181 ne
rect 6874 165 6918 181
tri 6918 165 6934 181 nw
rect 6964 261 7022 296
tri 7128 266 7158 296 ne
rect 6964 227 6976 261
rect 7010 227 7022 261
tri 7053 251 7068 266 se
rect 7068 251 7112 266
tri 7112 251 7127 266 sw
rect 7158 261 7214 296
rect 6964 193 7022 227
rect 6772 135 6828 159
tri 6828 135 6858 165 sw
tri 6934 135 6964 165 se
rect 6964 159 6976 193
rect 7010 159 7022 193
rect 7052 217 7128 251
rect 7052 183 7073 217
rect 7107 183 7128 217
rect 7052 181 7128 183
tri 7052 165 7068 181 ne
rect 7068 165 7112 181
tri 7112 165 7128 181 nw
rect 7158 227 7170 261
rect 7204 227 7214 261
rect 7158 193 7214 227
rect 6964 135 7022 159
tri 7022 135 7052 165 sw
tri 7128 135 7158 165 se
rect 7158 159 7170 193
rect 7204 159 7214 193
rect 7158 135 7214 159
rect 6772 123 7214 135
rect 6772 89 6782 123
rect 6816 89 6879 123
rect 6913 89 6976 123
rect 7010 89 7073 123
rect 7107 89 7170 123
rect 7204 89 7214 123
rect 6772 73 7214 89
rect 7425 334 7481 350
rect 7425 300 7435 334
rect 7469 300 7481 334
rect 7425 262 7481 300
rect 7511 334 7671 350
rect 7511 313 7629 334
tri 7511 297 7527 313 ne
rect 7527 300 7629 313
rect 7663 300 7671 334
rect 7527 297 7671 300
tri 7587 267 7617 297 ne
rect 7425 228 7435 262
rect 7469 228 7481 262
rect 7425 194 7481 228
rect 7425 160 7435 194
rect 7469 160 7481 194
tri 7511 251 7527 267 se
rect 7527 251 7571 267
tri 7571 251 7587 267 sw
rect 7511 218 7587 251
rect 7511 184 7531 218
rect 7565 184 7587 218
rect 7511 182 7587 184
tri 7511 166 7527 182 ne
rect 7527 166 7571 182
tri 7571 166 7587 182 nw
rect 7617 262 7671 297
rect 7617 228 7629 262
rect 7663 228 7671 262
rect 7617 194 7671 228
rect 7425 136 7481 160
tri 7481 136 7511 166 sw
tri 7587 136 7617 166 se
rect 7617 160 7629 194
rect 7663 160 7671 194
rect 7617 136 7671 160
rect 7425 124 7671 136
rect 7425 90 7435 124
rect 7469 90 7531 124
rect 7565 90 7629 124
rect 7663 90 7671 124
rect 7425 74 7671 90
<< pdiff >>
rect 108 1366 164 1404
rect 108 1332 118 1366
rect 152 1332 164 1366
rect 108 1298 164 1332
rect 108 1264 118 1298
rect 152 1264 164 1298
rect 108 1230 164 1264
rect 108 1196 118 1230
rect 152 1196 164 1230
rect 108 1162 164 1196
rect 108 1128 118 1162
rect 152 1128 164 1162
rect 108 1093 164 1128
rect 108 1059 118 1093
rect 152 1059 164 1093
rect 108 1004 164 1059
rect 194 1366 252 1404
rect 194 1332 206 1366
rect 240 1332 252 1366
rect 194 1298 252 1332
rect 194 1264 206 1298
rect 240 1264 252 1298
rect 194 1230 252 1264
rect 194 1196 206 1230
rect 240 1196 252 1230
rect 194 1162 252 1196
rect 194 1128 206 1162
rect 240 1128 252 1162
rect 194 1093 252 1128
rect 194 1059 206 1093
rect 240 1059 252 1093
rect 194 1004 252 1059
rect 282 1366 336 1404
rect 282 1332 294 1366
rect 328 1332 336 1366
rect 282 1298 336 1332
rect 282 1264 294 1298
rect 328 1264 336 1298
rect 282 1230 336 1264
rect 282 1196 294 1230
rect 328 1196 336 1230
rect 282 1162 336 1196
rect 282 1128 294 1162
rect 328 1128 336 1162
rect 282 1093 336 1128
rect 282 1059 294 1093
rect 328 1059 336 1093
rect 282 1004 336 1059
rect 575 1364 631 1404
rect 575 1330 585 1364
rect 619 1330 631 1364
rect 575 1296 631 1330
rect 575 1262 585 1296
rect 619 1262 631 1296
rect 575 1228 631 1262
rect 575 1194 585 1228
rect 619 1194 631 1228
rect 575 1160 631 1194
rect 575 1126 585 1160
rect 619 1126 631 1160
rect 575 1092 631 1126
rect 575 1058 585 1092
rect 619 1058 631 1092
rect 575 1004 631 1058
rect 661 1296 719 1404
rect 661 1262 673 1296
rect 707 1262 719 1296
rect 661 1228 719 1262
rect 661 1194 673 1228
rect 707 1194 719 1228
rect 661 1160 719 1194
rect 661 1126 673 1160
rect 707 1126 719 1160
rect 661 1004 719 1126
rect 749 1364 807 1404
rect 749 1330 761 1364
rect 795 1330 807 1364
rect 749 1296 807 1330
rect 749 1262 761 1296
rect 795 1262 807 1296
rect 749 1228 807 1262
rect 749 1194 761 1228
rect 795 1194 807 1228
rect 749 1160 807 1194
rect 749 1126 761 1160
rect 795 1126 807 1160
rect 749 1092 807 1126
rect 749 1058 761 1092
rect 795 1058 807 1092
rect 749 1004 807 1058
rect 837 1296 895 1404
rect 837 1262 849 1296
rect 883 1262 895 1296
rect 837 1228 895 1262
rect 837 1194 849 1228
rect 883 1194 895 1228
rect 837 1160 895 1194
rect 837 1126 849 1160
rect 883 1126 895 1160
rect 837 1092 895 1126
rect 837 1058 849 1092
rect 883 1058 895 1092
rect 837 1004 895 1058
rect 925 1364 979 1404
rect 925 1330 937 1364
rect 971 1330 979 1364
rect 925 1296 979 1330
rect 925 1262 937 1296
rect 971 1262 979 1296
rect 925 1228 979 1262
rect 925 1194 937 1228
rect 971 1194 979 1228
rect 925 1160 979 1194
rect 925 1126 937 1160
rect 971 1126 979 1160
rect 925 1004 979 1126
rect 1241 1364 1297 1404
rect 1241 1330 1251 1364
rect 1285 1330 1297 1364
rect 1241 1296 1297 1330
rect 1241 1262 1251 1296
rect 1285 1262 1297 1296
rect 1241 1228 1297 1262
rect 1241 1194 1251 1228
rect 1285 1194 1297 1228
rect 1241 1160 1297 1194
rect 1241 1126 1251 1160
rect 1285 1126 1297 1160
rect 1241 1092 1297 1126
rect 1241 1058 1251 1092
rect 1285 1058 1297 1092
rect 1241 1004 1297 1058
rect 1327 1296 1385 1404
rect 1327 1262 1339 1296
rect 1373 1262 1385 1296
rect 1327 1228 1385 1262
rect 1327 1194 1339 1228
rect 1373 1194 1385 1228
rect 1327 1160 1385 1194
rect 1327 1126 1339 1160
rect 1373 1126 1385 1160
rect 1327 1004 1385 1126
rect 1415 1364 1473 1404
rect 1415 1330 1427 1364
rect 1461 1330 1473 1364
rect 1415 1296 1473 1330
rect 1415 1262 1427 1296
rect 1461 1262 1473 1296
rect 1415 1228 1473 1262
rect 1415 1194 1427 1228
rect 1461 1194 1473 1228
rect 1415 1160 1473 1194
rect 1415 1126 1427 1160
rect 1461 1126 1473 1160
rect 1415 1092 1473 1126
rect 1415 1058 1427 1092
rect 1461 1058 1473 1092
rect 1415 1004 1473 1058
rect 1503 1296 1561 1404
rect 1503 1262 1515 1296
rect 1549 1262 1561 1296
rect 1503 1228 1561 1262
rect 1503 1194 1515 1228
rect 1549 1194 1561 1228
rect 1503 1160 1561 1194
rect 1503 1126 1515 1160
rect 1549 1126 1561 1160
rect 1503 1092 1561 1126
rect 1503 1058 1515 1092
rect 1549 1058 1561 1092
rect 1503 1004 1561 1058
rect 1591 1364 1645 1404
rect 1591 1330 1603 1364
rect 1637 1330 1645 1364
rect 1591 1296 1645 1330
rect 1591 1262 1603 1296
rect 1637 1262 1645 1296
rect 1591 1228 1645 1262
rect 1591 1194 1603 1228
rect 1637 1194 1645 1228
rect 1591 1160 1645 1194
rect 1591 1126 1603 1160
rect 1637 1126 1645 1160
rect 1591 1004 1645 1126
rect 1884 1366 1938 1404
rect 1884 1332 1892 1366
rect 1926 1332 1938 1366
rect 1884 1298 1938 1332
rect 1884 1264 1892 1298
rect 1926 1264 1938 1298
rect 1884 1230 1938 1264
rect 1884 1196 1892 1230
rect 1926 1196 1938 1230
rect 1884 1162 1938 1196
rect 1884 1128 1892 1162
rect 1926 1128 1938 1162
rect 1884 1093 1938 1128
rect 1884 1059 1892 1093
rect 1926 1059 1938 1093
rect 1884 1004 1938 1059
rect 1968 1366 2026 1404
rect 1968 1332 1980 1366
rect 2014 1332 2026 1366
rect 1968 1298 2026 1332
rect 1968 1264 1980 1298
rect 2014 1264 2026 1298
rect 1968 1230 2026 1264
rect 1968 1196 1980 1230
rect 2014 1196 2026 1230
rect 1968 1162 2026 1196
rect 1968 1128 1980 1162
rect 2014 1128 2026 1162
rect 1968 1093 2026 1128
rect 1968 1059 1980 1093
rect 2014 1059 2026 1093
rect 1968 1004 2026 1059
rect 2056 1366 2112 1404
rect 2056 1332 2068 1366
rect 2102 1332 2112 1366
rect 2056 1298 2112 1332
rect 2056 1264 2068 1298
rect 2102 1264 2112 1298
rect 2056 1230 2112 1264
rect 2056 1196 2068 1230
rect 2102 1196 2112 1230
rect 2056 1162 2112 1196
rect 2056 1128 2068 1162
rect 2102 1128 2112 1162
rect 2056 1093 2112 1128
rect 2056 1059 2068 1093
rect 2102 1059 2112 1093
rect 2056 1004 2112 1059
rect 2328 1366 2384 1404
rect 2328 1332 2338 1366
rect 2372 1332 2384 1366
rect 2328 1298 2384 1332
rect 2328 1264 2338 1298
rect 2372 1264 2384 1298
rect 2328 1230 2384 1264
rect 2328 1196 2338 1230
rect 2372 1196 2384 1230
rect 2328 1162 2384 1196
rect 2328 1128 2338 1162
rect 2372 1128 2384 1162
rect 2328 1093 2384 1128
rect 2328 1059 2338 1093
rect 2372 1059 2384 1093
rect 2328 1004 2384 1059
rect 2414 1366 2472 1404
rect 2414 1332 2426 1366
rect 2460 1332 2472 1366
rect 2414 1298 2472 1332
rect 2414 1264 2426 1298
rect 2460 1264 2472 1298
rect 2414 1230 2472 1264
rect 2414 1196 2426 1230
rect 2460 1196 2472 1230
rect 2414 1162 2472 1196
rect 2414 1128 2426 1162
rect 2460 1128 2472 1162
rect 2414 1093 2472 1128
rect 2414 1059 2426 1093
rect 2460 1059 2472 1093
rect 2414 1004 2472 1059
rect 2502 1366 2556 1404
rect 2502 1332 2514 1366
rect 2548 1332 2556 1366
rect 2502 1298 2556 1332
rect 2502 1264 2514 1298
rect 2548 1264 2556 1298
rect 2502 1230 2556 1264
rect 2502 1196 2514 1230
rect 2548 1196 2556 1230
rect 2502 1162 2556 1196
rect 2502 1128 2514 1162
rect 2548 1128 2556 1162
rect 2502 1093 2556 1128
rect 2502 1059 2514 1093
rect 2548 1059 2556 1093
rect 2502 1004 2556 1059
rect 2795 1364 2851 1404
rect 2795 1330 2805 1364
rect 2839 1330 2851 1364
rect 2795 1296 2851 1330
rect 2795 1262 2805 1296
rect 2839 1262 2851 1296
rect 2795 1228 2851 1262
rect 2795 1194 2805 1228
rect 2839 1194 2851 1228
rect 2795 1160 2851 1194
rect 2795 1126 2805 1160
rect 2839 1126 2851 1160
rect 2795 1092 2851 1126
rect 2795 1058 2805 1092
rect 2839 1058 2851 1092
rect 2795 1004 2851 1058
rect 2881 1296 2939 1404
rect 2881 1262 2893 1296
rect 2927 1262 2939 1296
rect 2881 1228 2939 1262
rect 2881 1194 2893 1228
rect 2927 1194 2939 1228
rect 2881 1160 2939 1194
rect 2881 1126 2893 1160
rect 2927 1126 2939 1160
rect 2881 1004 2939 1126
rect 2969 1364 3027 1404
rect 2969 1330 2981 1364
rect 3015 1330 3027 1364
rect 2969 1296 3027 1330
rect 2969 1262 2981 1296
rect 3015 1262 3027 1296
rect 2969 1228 3027 1262
rect 2969 1194 2981 1228
rect 3015 1194 3027 1228
rect 2969 1160 3027 1194
rect 2969 1126 2981 1160
rect 3015 1126 3027 1160
rect 2969 1092 3027 1126
rect 2969 1058 2981 1092
rect 3015 1058 3027 1092
rect 2969 1004 3027 1058
rect 3057 1296 3115 1404
rect 3057 1262 3069 1296
rect 3103 1262 3115 1296
rect 3057 1228 3115 1262
rect 3057 1194 3069 1228
rect 3103 1194 3115 1228
rect 3057 1160 3115 1194
rect 3057 1126 3069 1160
rect 3103 1126 3115 1160
rect 3057 1092 3115 1126
rect 3057 1058 3069 1092
rect 3103 1058 3115 1092
rect 3057 1004 3115 1058
rect 3145 1364 3199 1404
rect 3145 1330 3157 1364
rect 3191 1330 3199 1364
rect 3145 1296 3199 1330
rect 3145 1262 3157 1296
rect 3191 1262 3199 1296
rect 3145 1228 3199 1262
rect 3145 1194 3157 1228
rect 3191 1194 3199 1228
rect 3145 1160 3199 1194
rect 3145 1126 3157 1160
rect 3191 1126 3199 1160
rect 3145 1004 3199 1126
rect 3461 1364 3517 1404
rect 3461 1330 3471 1364
rect 3505 1330 3517 1364
rect 3461 1296 3517 1330
rect 3461 1262 3471 1296
rect 3505 1262 3517 1296
rect 3461 1228 3517 1262
rect 3461 1194 3471 1228
rect 3505 1194 3517 1228
rect 3461 1160 3517 1194
rect 3461 1126 3471 1160
rect 3505 1126 3517 1160
rect 3461 1092 3517 1126
rect 3461 1058 3471 1092
rect 3505 1058 3517 1092
rect 3461 1004 3517 1058
rect 3547 1296 3605 1404
rect 3547 1262 3559 1296
rect 3593 1262 3605 1296
rect 3547 1228 3605 1262
rect 3547 1194 3559 1228
rect 3593 1194 3605 1228
rect 3547 1160 3605 1194
rect 3547 1126 3559 1160
rect 3593 1126 3605 1160
rect 3547 1004 3605 1126
rect 3635 1364 3693 1404
rect 3635 1330 3647 1364
rect 3681 1330 3693 1364
rect 3635 1296 3693 1330
rect 3635 1262 3647 1296
rect 3681 1262 3693 1296
rect 3635 1228 3693 1262
rect 3635 1194 3647 1228
rect 3681 1194 3693 1228
rect 3635 1160 3693 1194
rect 3635 1126 3647 1160
rect 3681 1126 3693 1160
rect 3635 1092 3693 1126
rect 3635 1058 3647 1092
rect 3681 1058 3693 1092
rect 3635 1004 3693 1058
rect 3723 1296 3781 1404
rect 3723 1262 3735 1296
rect 3769 1262 3781 1296
rect 3723 1228 3781 1262
rect 3723 1194 3735 1228
rect 3769 1194 3781 1228
rect 3723 1160 3781 1194
rect 3723 1126 3735 1160
rect 3769 1126 3781 1160
rect 3723 1092 3781 1126
rect 3723 1058 3735 1092
rect 3769 1058 3781 1092
rect 3723 1004 3781 1058
rect 3811 1364 3865 1404
rect 3811 1330 3823 1364
rect 3857 1330 3865 1364
rect 3811 1296 3865 1330
rect 3811 1262 3823 1296
rect 3857 1262 3865 1296
rect 3811 1228 3865 1262
rect 3811 1194 3823 1228
rect 3857 1194 3865 1228
rect 3811 1160 3865 1194
rect 3811 1126 3823 1160
rect 3857 1126 3865 1160
rect 3811 1004 3865 1126
rect 4104 1366 4158 1404
rect 4104 1332 4112 1366
rect 4146 1332 4158 1366
rect 4104 1298 4158 1332
rect 4104 1264 4112 1298
rect 4146 1264 4158 1298
rect 4104 1230 4158 1264
rect 4104 1196 4112 1230
rect 4146 1196 4158 1230
rect 4104 1162 4158 1196
rect 4104 1128 4112 1162
rect 4146 1128 4158 1162
rect 4104 1093 4158 1128
rect 4104 1059 4112 1093
rect 4146 1059 4158 1093
rect 4104 1004 4158 1059
rect 4188 1366 4246 1404
rect 4188 1332 4200 1366
rect 4234 1332 4246 1366
rect 4188 1298 4246 1332
rect 4188 1264 4200 1298
rect 4234 1264 4246 1298
rect 4188 1230 4246 1264
rect 4188 1196 4200 1230
rect 4234 1196 4246 1230
rect 4188 1162 4246 1196
rect 4188 1128 4200 1162
rect 4234 1128 4246 1162
rect 4188 1093 4246 1128
rect 4188 1059 4200 1093
rect 4234 1059 4246 1093
rect 4188 1004 4246 1059
rect 4276 1366 4332 1404
rect 4276 1332 4288 1366
rect 4322 1332 4332 1366
rect 4276 1298 4332 1332
rect 4276 1264 4288 1298
rect 4322 1264 4332 1298
rect 4276 1230 4332 1264
rect 4276 1196 4288 1230
rect 4322 1196 4332 1230
rect 4276 1162 4332 1196
rect 4276 1128 4288 1162
rect 4322 1128 4332 1162
rect 4276 1093 4332 1128
rect 4276 1059 4288 1093
rect 4322 1059 4332 1093
rect 4276 1004 4332 1059
rect 4571 1366 4627 1404
rect 4571 1332 4581 1366
rect 4615 1332 4627 1366
rect 4571 1298 4627 1332
rect 4571 1264 4581 1298
rect 4615 1264 4627 1298
rect 4571 1230 4627 1264
rect 4571 1196 4581 1230
rect 4615 1196 4627 1230
rect 4571 1162 4627 1196
rect 4571 1128 4581 1162
rect 4615 1128 4627 1162
rect 4571 1093 4627 1128
rect 4571 1059 4581 1093
rect 4615 1059 4627 1093
rect 4571 1004 4627 1059
rect 4657 1366 4715 1404
rect 4657 1332 4669 1366
rect 4703 1332 4715 1366
rect 4657 1298 4715 1332
rect 4657 1264 4669 1298
rect 4703 1264 4715 1298
rect 4657 1230 4715 1264
rect 4657 1196 4669 1230
rect 4703 1196 4715 1230
rect 4657 1162 4715 1196
rect 4657 1128 4669 1162
rect 4703 1128 4715 1162
rect 4657 1093 4715 1128
rect 4657 1059 4669 1093
rect 4703 1059 4715 1093
rect 4657 1004 4715 1059
rect 4745 1366 4803 1404
rect 4745 1332 4757 1366
rect 4791 1332 4803 1366
rect 4745 1298 4803 1332
rect 4745 1264 4757 1298
rect 4791 1264 4803 1298
rect 4745 1230 4803 1264
rect 4745 1196 4757 1230
rect 4791 1196 4803 1230
rect 4745 1162 4803 1196
rect 4745 1128 4757 1162
rect 4791 1128 4803 1162
rect 4745 1004 4803 1128
rect 4833 1366 4891 1404
rect 4833 1332 4845 1366
rect 4879 1332 4891 1366
rect 4833 1298 4891 1332
rect 4833 1264 4845 1298
rect 4879 1264 4891 1298
rect 4833 1230 4891 1264
rect 4833 1196 4845 1230
rect 4879 1196 4891 1230
rect 4833 1162 4891 1196
rect 4833 1128 4845 1162
rect 4879 1128 4891 1162
rect 4833 1093 4891 1128
rect 4833 1059 4845 1093
rect 4879 1059 4891 1093
rect 4833 1004 4891 1059
rect 4921 1366 4975 1404
rect 4921 1332 4933 1366
rect 4967 1332 4975 1366
rect 4921 1298 4975 1332
rect 4921 1264 4933 1298
rect 4967 1264 4975 1298
rect 4921 1230 4975 1264
rect 4921 1196 4933 1230
rect 4967 1196 4975 1230
rect 4921 1162 4975 1196
rect 4921 1128 4933 1162
rect 4967 1128 4975 1162
rect 4921 1004 4975 1128
rect 5214 1366 5270 1404
rect 5214 1332 5224 1366
rect 5258 1332 5270 1366
rect 5214 1298 5270 1332
rect 5214 1264 5224 1298
rect 5258 1264 5270 1298
rect 5214 1230 5270 1264
rect 5214 1196 5224 1230
rect 5258 1196 5270 1230
rect 5214 1162 5270 1196
rect 5214 1128 5224 1162
rect 5258 1128 5270 1162
rect 5214 1093 5270 1128
rect 5214 1059 5224 1093
rect 5258 1059 5270 1093
rect 5214 1004 5270 1059
rect 5300 1366 5358 1404
rect 5300 1332 5312 1366
rect 5346 1332 5358 1366
rect 5300 1298 5358 1332
rect 5300 1264 5312 1298
rect 5346 1264 5358 1298
rect 5300 1230 5358 1264
rect 5300 1196 5312 1230
rect 5346 1196 5358 1230
rect 5300 1162 5358 1196
rect 5300 1128 5312 1162
rect 5346 1128 5358 1162
rect 5300 1093 5358 1128
rect 5300 1059 5312 1093
rect 5346 1059 5358 1093
rect 5300 1004 5358 1059
rect 5388 1366 5442 1404
rect 5388 1332 5400 1366
rect 5434 1332 5442 1366
rect 5388 1298 5442 1332
rect 5388 1264 5400 1298
rect 5434 1264 5442 1298
rect 5388 1230 5442 1264
rect 5388 1196 5400 1230
rect 5434 1196 5442 1230
rect 5388 1162 5442 1196
rect 5388 1128 5400 1162
rect 5434 1128 5442 1162
rect 5388 1093 5442 1128
rect 5388 1059 5400 1093
rect 5434 1059 5442 1093
rect 5388 1004 5442 1059
rect 5681 1366 5737 1404
rect 5681 1332 5691 1366
rect 5725 1332 5737 1366
rect 5681 1298 5737 1332
rect 5681 1264 5691 1298
rect 5725 1264 5737 1298
rect 5681 1230 5737 1264
rect 5681 1196 5691 1230
rect 5725 1196 5737 1230
rect 5681 1162 5737 1196
rect 5681 1128 5691 1162
rect 5725 1128 5737 1162
rect 5681 1093 5737 1128
rect 5681 1059 5691 1093
rect 5725 1059 5737 1093
rect 5681 1004 5737 1059
rect 5767 1366 5825 1404
rect 5767 1332 5779 1366
rect 5813 1332 5825 1366
rect 5767 1298 5825 1332
rect 5767 1264 5779 1298
rect 5813 1264 5825 1298
rect 5767 1230 5825 1264
rect 5767 1196 5779 1230
rect 5813 1196 5825 1230
rect 5767 1162 5825 1196
rect 5767 1128 5779 1162
rect 5813 1128 5825 1162
rect 5767 1093 5825 1128
rect 5767 1059 5779 1093
rect 5813 1059 5825 1093
rect 5767 1004 5825 1059
rect 5855 1366 5913 1404
rect 5855 1332 5867 1366
rect 5901 1332 5913 1366
rect 5855 1298 5913 1332
rect 5855 1264 5867 1298
rect 5901 1264 5913 1298
rect 5855 1230 5913 1264
rect 5855 1196 5867 1230
rect 5901 1196 5913 1230
rect 5855 1162 5913 1196
rect 5855 1128 5867 1162
rect 5901 1128 5913 1162
rect 5855 1004 5913 1128
rect 5943 1366 6001 1404
rect 5943 1332 5955 1366
rect 5989 1332 6001 1366
rect 5943 1298 6001 1332
rect 5943 1264 5955 1298
rect 5989 1264 6001 1298
rect 5943 1230 6001 1264
rect 5943 1196 5955 1230
rect 5989 1196 6001 1230
rect 5943 1162 6001 1196
rect 5943 1128 5955 1162
rect 5989 1128 6001 1162
rect 5943 1093 6001 1128
rect 5943 1059 5955 1093
rect 5989 1059 6001 1093
rect 5943 1004 6001 1059
rect 6031 1366 6085 1404
rect 6031 1332 6043 1366
rect 6077 1332 6085 1366
rect 6031 1298 6085 1332
rect 6031 1264 6043 1298
rect 6077 1264 6085 1298
rect 6031 1230 6085 1264
rect 6031 1196 6043 1230
rect 6077 1196 6085 1230
rect 6031 1162 6085 1196
rect 6031 1128 6043 1162
rect 6077 1128 6085 1162
rect 6031 1004 6085 1128
rect 6324 1366 6380 1404
rect 6324 1332 6334 1366
rect 6368 1332 6380 1366
rect 6324 1298 6380 1332
rect 6324 1264 6334 1298
rect 6368 1264 6380 1298
rect 6324 1230 6380 1264
rect 6324 1196 6334 1230
rect 6368 1196 6380 1230
rect 6324 1162 6380 1196
rect 6324 1128 6334 1162
rect 6368 1128 6380 1162
rect 6324 1093 6380 1128
rect 6324 1059 6334 1093
rect 6368 1059 6380 1093
rect 6324 1004 6380 1059
rect 6410 1366 6468 1404
rect 6410 1332 6422 1366
rect 6456 1332 6468 1366
rect 6410 1298 6468 1332
rect 6410 1264 6422 1298
rect 6456 1264 6468 1298
rect 6410 1230 6468 1264
rect 6410 1196 6422 1230
rect 6456 1196 6468 1230
rect 6410 1162 6468 1196
rect 6410 1128 6422 1162
rect 6456 1128 6468 1162
rect 6410 1093 6468 1128
rect 6410 1059 6422 1093
rect 6456 1059 6468 1093
rect 6410 1004 6468 1059
rect 6498 1366 6552 1404
rect 6498 1332 6510 1366
rect 6544 1332 6552 1366
rect 6498 1298 6552 1332
rect 6498 1264 6510 1298
rect 6544 1264 6552 1298
rect 6498 1230 6552 1264
rect 6498 1196 6510 1230
rect 6544 1196 6552 1230
rect 6498 1162 6552 1196
rect 6498 1128 6510 1162
rect 6544 1128 6552 1162
rect 6498 1093 6552 1128
rect 6498 1059 6510 1093
rect 6544 1059 6552 1093
rect 6498 1004 6552 1059
rect 6791 1365 6847 1405
rect 6791 1331 6801 1365
rect 6835 1331 6847 1365
rect 6791 1297 6847 1331
rect 6791 1263 6801 1297
rect 6835 1263 6847 1297
rect 6791 1229 6847 1263
rect 6791 1195 6801 1229
rect 6835 1195 6847 1229
rect 6791 1161 6847 1195
rect 6791 1127 6801 1161
rect 6835 1127 6847 1161
rect 6791 1093 6847 1127
rect 6791 1059 6801 1093
rect 6835 1059 6847 1093
rect 6791 1005 6847 1059
rect 6877 1365 6935 1405
rect 6877 1331 6889 1365
rect 6923 1331 6935 1365
rect 6877 1297 6935 1331
rect 6877 1263 6889 1297
rect 6923 1263 6935 1297
rect 6877 1229 6935 1263
rect 6877 1195 6889 1229
rect 6923 1195 6935 1229
rect 6877 1161 6935 1195
rect 6877 1127 6889 1161
rect 6923 1127 6935 1161
rect 6877 1005 6935 1127
rect 6965 1365 7023 1405
rect 6965 1331 6977 1365
rect 7011 1331 7023 1365
rect 6965 1297 7023 1331
rect 6965 1263 6977 1297
rect 7011 1263 7023 1297
rect 6965 1229 7023 1263
rect 6965 1195 6977 1229
rect 7011 1195 7023 1229
rect 6965 1161 7023 1195
rect 6965 1127 6977 1161
rect 7011 1127 7023 1161
rect 6965 1093 7023 1127
rect 6965 1059 6977 1093
rect 7011 1059 7023 1093
rect 6965 1005 7023 1059
rect 7053 1297 7111 1405
rect 7053 1263 7065 1297
rect 7099 1263 7111 1297
rect 7053 1229 7111 1263
rect 7053 1195 7065 1229
rect 7099 1195 7111 1229
rect 7053 1161 7111 1195
rect 7053 1127 7065 1161
rect 7099 1127 7111 1161
rect 7053 1093 7111 1127
rect 7053 1059 7065 1093
rect 7099 1059 7111 1093
rect 7053 1005 7111 1059
rect 7141 1365 7195 1405
rect 7141 1331 7153 1365
rect 7187 1331 7195 1365
rect 7141 1297 7195 1331
rect 7141 1263 7153 1297
rect 7187 1263 7195 1297
rect 7141 1229 7195 1263
rect 7141 1195 7153 1229
rect 7187 1195 7195 1229
rect 7141 1161 7195 1195
rect 7141 1127 7153 1161
rect 7187 1127 7195 1161
rect 7141 1005 7195 1127
rect 7434 1366 7490 1404
rect 7434 1332 7444 1366
rect 7478 1332 7490 1366
rect 7434 1298 7490 1332
rect 7434 1264 7444 1298
rect 7478 1264 7490 1298
rect 7434 1230 7490 1264
rect 7434 1196 7444 1230
rect 7478 1196 7490 1230
rect 7434 1162 7490 1196
rect 7434 1128 7444 1162
rect 7478 1128 7490 1162
rect 7434 1093 7490 1128
rect 7434 1059 7444 1093
rect 7478 1059 7490 1093
rect 7434 1004 7490 1059
rect 7520 1366 7578 1404
rect 7520 1332 7532 1366
rect 7566 1332 7578 1366
rect 7520 1298 7578 1332
rect 7520 1264 7532 1298
rect 7566 1264 7578 1298
rect 7520 1230 7578 1264
rect 7520 1196 7532 1230
rect 7566 1196 7578 1230
rect 7520 1162 7578 1196
rect 7520 1128 7532 1162
rect 7566 1128 7578 1162
rect 7520 1093 7578 1128
rect 7520 1059 7532 1093
rect 7566 1059 7578 1093
rect 7520 1004 7578 1059
rect 7608 1366 7662 1404
rect 7608 1332 7620 1366
rect 7654 1332 7662 1366
rect 7608 1298 7662 1332
rect 7608 1264 7620 1298
rect 7654 1264 7662 1298
rect 7608 1230 7662 1264
rect 7608 1196 7620 1230
rect 7654 1196 7662 1230
rect 7608 1162 7662 1196
rect 7608 1128 7620 1162
rect 7654 1128 7662 1162
rect 7608 1093 7662 1128
rect 7608 1059 7620 1093
rect 7654 1059 7662 1093
rect 7608 1004 7662 1059
<< ndiffc >>
rect 109 300 143 334
rect 303 300 337 334
rect 109 228 143 262
rect 109 160 143 194
rect 205 184 239 218
rect 303 228 337 262
rect 303 160 337 194
rect 109 90 143 124
rect 205 90 239 124
rect 303 90 337 124
rect 566 300 600 334
rect 663 300 697 334
rect 760 300 794 334
rect 566 228 600 262
rect 566 160 600 194
rect 663 175 697 209
rect 760 228 794 262
rect 760 160 794 194
rect 857 184 891 218
rect 954 228 988 262
rect 954 160 988 194
rect 566 90 600 124
rect 760 90 794 124
rect 857 90 891 124
rect 954 90 988 124
rect 1232 300 1266 334
rect 1329 300 1363 334
rect 1426 300 1460 334
rect 1232 228 1266 262
rect 1232 160 1266 194
rect 1329 175 1363 209
rect 1426 228 1460 262
rect 1426 160 1460 194
rect 1523 184 1557 218
rect 1620 228 1654 262
rect 1620 160 1654 194
rect 1232 90 1266 124
rect 1426 90 1460 124
rect 1523 90 1557 124
rect 1620 90 1654 124
rect 1883 300 1917 334
rect 2077 300 2111 334
rect 1883 228 1917 262
rect 1883 160 1917 194
rect 1981 184 2015 218
rect 2077 228 2111 262
rect 2077 160 2111 194
rect 1883 90 1917 124
rect 1981 90 2015 124
rect 2077 90 2111 124
rect 2329 300 2363 334
rect 2523 300 2557 334
rect 2329 228 2363 262
rect 2329 160 2363 194
rect 2425 184 2459 218
rect 2523 228 2557 262
rect 2523 160 2557 194
rect 2329 90 2363 124
rect 2425 90 2459 124
rect 2523 90 2557 124
rect 2786 300 2820 334
rect 2883 300 2917 334
rect 2980 300 3014 334
rect 2786 228 2820 262
rect 2786 160 2820 194
rect 2883 175 2917 209
rect 2980 228 3014 262
rect 2980 160 3014 194
rect 3077 184 3111 218
rect 3174 228 3208 262
rect 3174 160 3208 194
rect 2786 90 2820 124
rect 2980 90 3014 124
rect 3077 90 3111 124
rect 3174 90 3208 124
rect 3452 300 3486 334
rect 3549 300 3583 334
rect 3646 300 3680 334
rect 3452 228 3486 262
rect 3452 160 3486 194
rect 3549 175 3583 209
rect 3646 228 3680 262
rect 3646 160 3680 194
rect 3743 184 3777 218
rect 3840 228 3874 262
rect 3840 160 3874 194
rect 3452 90 3486 124
rect 3646 90 3680 124
rect 3743 90 3777 124
rect 3840 90 3874 124
rect 4103 300 4137 334
rect 4297 300 4331 334
rect 4103 228 4137 262
rect 4103 160 4137 194
rect 4201 184 4235 218
rect 4297 228 4331 262
rect 4297 160 4331 194
rect 4103 90 4137 124
rect 4201 90 4235 124
rect 4297 90 4331 124
rect 4562 299 4596 333
rect 4659 299 4693 333
rect 4756 299 4790 333
rect 4562 227 4596 261
rect 4562 159 4596 193
rect 4659 174 4693 208
rect 4756 227 4790 261
rect 4756 159 4790 193
rect 4853 183 4887 217
rect 4950 227 4984 261
rect 4950 159 4984 193
rect 4562 89 4596 123
rect 4756 89 4790 123
rect 4853 89 4887 123
rect 4950 89 4984 123
rect 5215 300 5249 334
rect 5409 300 5443 334
rect 5215 228 5249 262
rect 5215 160 5249 194
rect 5311 184 5345 218
rect 5409 228 5443 262
rect 5409 160 5443 194
rect 5215 90 5249 124
rect 5311 90 5345 124
rect 5409 90 5443 124
rect 5672 299 5706 333
rect 5769 299 5803 333
rect 5866 299 5900 333
rect 5672 227 5706 261
rect 5672 159 5706 193
rect 5769 174 5803 208
rect 5866 227 5900 261
rect 5866 159 5900 193
rect 5963 183 5997 217
rect 6060 227 6094 261
rect 6060 159 6094 193
rect 5672 89 5706 123
rect 5866 89 5900 123
rect 5963 89 5997 123
rect 6060 89 6094 123
rect 6325 300 6359 334
rect 6519 300 6553 334
rect 6325 228 6359 262
rect 6325 160 6359 194
rect 6421 184 6455 218
rect 6519 228 6553 262
rect 6519 160 6553 194
rect 6325 90 6359 124
rect 6421 90 6455 124
rect 6519 90 6553 124
rect 6782 299 6816 333
rect 6782 227 6816 261
rect 6782 159 6816 193
rect 6879 183 6913 217
rect 6976 227 7010 261
rect 6976 159 7010 193
rect 7073 183 7107 217
rect 7170 227 7204 261
rect 7170 159 7204 193
rect 6782 89 6816 123
rect 6879 89 6913 123
rect 6976 89 7010 123
rect 7073 89 7107 123
rect 7170 89 7204 123
rect 7435 300 7469 334
rect 7629 300 7663 334
rect 7435 228 7469 262
rect 7435 160 7469 194
rect 7531 184 7565 218
rect 7629 228 7663 262
rect 7629 160 7663 194
rect 7435 90 7469 124
rect 7531 90 7565 124
rect 7629 90 7663 124
<< pdiffc >>
rect 118 1332 152 1366
rect 118 1264 152 1298
rect 118 1196 152 1230
rect 118 1128 152 1162
rect 118 1059 152 1093
rect 206 1332 240 1366
rect 206 1264 240 1298
rect 206 1196 240 1230
rect 206 1128 240 1162
rect 206 1059 240 1093
rect 294 1332 328 1366
rect 294 1264 328 1298
rect 294 1196 328 1230
rect 294 1128 328 1162
rect 294 1059 328 1093
rect 585 1330 619 1364
rect 585 1262 619 1296
rect 585 1194 619 1228
rect 585 1126 619 1160
rect 585 1058 619 1092
rect 673 1262 707 1296
rect 673 1194 707 1228
rect 673 1126 707 1160
rect 761 1330 795 1364
rect 761 1262 795 1296
rect 761 1194 795 1228
rect 761 1126 795 1160
rect 761 1058 795 1092
rect 849 1262 883 1296
rect 849 1194 883 1228
rect 849 1126 883 1160
rect 849 1058 883 1092
rect 937 1330 971 1364
rect 937 1262 971 1296
rect 937 1194 971 1228
rect 937 1126 971 1160
rect 1251 1330 1285 1364
rect 1251 1262 1285 1296
rect 1251 1194 1285 1228
rect 1251 1126 1285 1160
rect 1251 1058 1285 1092
rect 1339 1262 1373 1296
rect 1339 1194 1373 1228
rect 1339 1126 1373 1160
rect 1427 1330 1461 1364
rect 1427 1262 1461 1296
rect 1427 1194 1461 1228
rect 1427 1126 1461 1160
rect 1427 1058 1461 1092
rect 1515 1262 1549 1296
rect 1515 1194 1549 1228
rect 1515 1126 1549 1160
rect 1515 1058 1549 1092
rect 1603 1330 1637 1364
rect 1603 1262 1637 1296
rect 1603 1194 1637 1228
rect 1603 1126 1637 1160
rect 1892 1332 1926 1366
rect 1892 1264 1926 1298
rect 1892 1196 1926 1230
rect 1892 1128 1926 1162
rect 1892 1059 1926 1093
rect 1980 1332 2014 1366
rect 1980 1264 2014 1298
rect 1980 1196 2014 1230
rect 1980 1128 2014 1162
rect 1980 1059 2014 1093
rect 2068 1332 2102 1366
rect 2068 1264 2102 1298
rect 2068 1196 2102 1230
rect 2068 1128 2102 1162
rect 2068 1059 2102 1093
rect 2338 1332 2372 1366
rect 2338 1264 2372 1298
rect 2338 1196 2372 1230
rect 2338 1128 2372 1162
rect 2338 1059 2372 1093
rect 2426 1332 2460 1366
rect 2426 1264 2460 1298
rect 2426 1196 2460 1230
rect 2426 1128 2460 1162
rect 2426 1059 2460 1093
rect 2514 1332 2548 1366
rect 2514 1264 2548 1298
rect 2514 1196 2548 1230
rect 2514 1128 2548 1162
rect 2514 1059 2548 1093
rect 2805 1330 2839 1364
rect 2805 1262 2839 1296
rect 2805 1194 2839 1228
rect 2805 1126 2839 1160
rect 2805 1058 2839 1092
rect 2893 1262 2927 1296
rect 2893 1194 2927 1228
rect 2893 1126 2927 1160
rect 2981 1330 3015 1364
rect 2981 1262 3015 1296
rect 2981 1194 3015 1228
rect 2981 1126 3015 1160
rect 2981 1058 3015 1092
rect 3069 1262 3103 1296
rect 3069 1194 3103 1228
rect 3069 1126 3103 1160
rect 3069 1058 3103 1092
rect 3157 1330 3191 1364
rect 3157 1262 3191 1296
rect 3157 1194 3191 1228
rect 3157 1126 3191 1160
rect 3471 1330 3505 1364
rect 3471 1262 3505 1296
rect 3471 1194 3505 1228
rect 3471 1126 3505 1160
rect 3471 1058 3505 1092
rect 3559 1262 3593 1296
rect 3559 1194 3593 1228
rect 3559 1126 3593 1160
rect 3647 1330 3681 1364
rect 3647 1262 3681 1296
rect 3647 1194 3681 1228
rect 3647 1126 3681 1160
rect 3647 1058 3681 1092
rect 3735 1262 3769 1296
rect 3735 1194 3769 1228
rect 3735 1126 3769 1160
rect 3735 1058 3769 1092
rect 3823 1330 3857 1364
rect 3823 1262 3857 1296
rect 3823 1194 3857 1228
rect 3823 1126 3857 1160
rect 4112 1332 4146 1366
rect 4112 1264 4146 1298
rect 4112 1196 4146 1230
rect 4112 1128 4146 1162
rect 4112 1059 4146 1093
rect 4200 1332 4234 1366
rect 4200 1264 4234 1298
rect 4200 1196 4234 1230
rect 4200 1128 4234 1162
rect 4200 1059 4234 1093
rect 4288 1332 4322 1366
rect 4288 1264 4322 1298
rect 4288 1196 4322 1230
rect 4288 1128 4322 1162
rect 4288 1059 4322 1093
rect 4581 1332 4615 1366
rect 4581 1264 4615 1298
rect 4581 1196 4615 1230
rect 4581 1128 4615 1162
rect 4581 1059 4615 1093
rect 4669 1332 4703 1366
rect 4669 1264 4703 1298
rect 4669 1196 4703 1230
rect 4669 1128 4703 1162
rect 4669 1059 4703 1093
rect 4757 1332 4791 1366
rect 4757 1264 4791 1298
rect 4757 1196 4791 1230
rect 4757 1128 4791 1162
rect 4845 1332 4879 1366
rect 4845 1264 4879 1298
rect 4845 1196 4879 1230
rect 4845 1128 4879 1162
rect 4845 1059 4879 1093
rect 4933 1332 4967 1366
rect 4933 1264 4967 1298
rect 4933 1196 4967 1230
rect 4933 1128 4967 1162
rect 5224 1332 5258 1366
rect 5224 1264 5258 1298
rect 5224 1196 5258 1230
rect 5224 1128 5258 1162
rect 5224 1059 5258 1093
rect 5312 1332 5346 1366
rect 5312 1264 5346 1298
rect 5312 1196 5346 1230
rect 5312 1128 5346 1162
rect 5312 1059 5346 1093
rect 5400 1332 5434 1366
rect 5400 1264 5434 1298
rect 5400 1196 5434 1230
rect 5400 1128 5434 1162
rect 5400 1059 5434 1093
rect 5691 1332 5725 1366
rect 5691 1264 5725 1298
rect 5691 1196 5725 1230
rect 5691 1128 5725 1162
rect 5691 1059 5725 1093
rect 5779 1332 5813 1366
rect 5779 1264 5813 1298
rect 5779 1196 5813 1230
rect 5779 1128 5813 1162
rect 5779 1059 5813 1093
rect 5867 1332 5901 1366
rect 5867 1264 5901 1298
rect 5867 1196 5901 1230
rect 5867 1128 5901 1162
rect 5955 1332 5989 1366
rect 5955 1264 5989 1298
rect 5955 1196 5989 1230
rect 5955 1128 5989 1162
rect 5955 1059 5989 1093
rect 6043 1332 6077 1366
rect 6043 1264 6077 1298
rect 6043 1196 6077 1230
rect 6043 1128 6077 1162
rect 6334 1332 6368 1366
rect 6334 1264 6368 1298
rect 6334 1196 6368 1230
rect 6334 1128 6368 1162
rect 6334 1059 6368 1093
rect 6422 1332 6456 1366
rect 6422 1264 6456 1298
rect 6422 1196 6456 1230
rect 6422 1128 6456 1162
rect 6422 1059 6456 1093
rect 6510 1332 6544 1366
rect 6510 1264 6544 1298
rect 6510 1196 6544 1230
rect 6510 1128 6544 1162
rect 6510 1059 6544 1093
rect 6801 1331 6835 1365
rect 6801 1263 6835 1297
rect 6801 1195 6835 1229
rect 6801 1127 6835 1161
rect 6801 1059 6835 1093
rect 6889 1331 6923 1365
rect 6889 1263 6923 1297
rect 6889 1195 6923 1229
rect 6889 1127 6923 1161
rect 6977 1331 7011 1365
rect 6977 1263 7011 1297
rect 6977 1195 7011 1229
rect 6977 1127 7011 1161
rect 6977 1059 7011 1093
rect 7065 1263 7099 1297
rect 7065 1195 7099 1229
rect 7065 1127 7099 1161
rect 7065 1059 7099 1093
rect 7153 1331 7187 1365
rect 7153 1263 7187 1297
rect 7153 1195 7187 1229
rect 7153 1127 7187 1161
rect 7444 1332 7478 1366
rect 7444 1264 7478 1298
rect 7444 1196 7478 1230
rect 7444 1128 7478 1162
rect 7444 1059 7478 1093
rect 7532 1332 7566 1366
rect 7532 1264 7566 1298
rect 7532 1196 7566 1230
rect 7532 1128 7566 1162
rect 7532 1059 7566 1093
rect 7620 1332 7654 1366
rect 7620 1264 7654 1298
rect 7620 1196 7654 1230
rect 7620 1128 7654 1162
rect 7620 1059 7654 1093
<< psubdiff >>
rect -34 482 7804 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 410 461 478 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 410 427 427 461
rect 461 427 478 461
rect 1076 461 1144 482
rect -34 313 34 353
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 410 313 478 353
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 1742 461 1810 482
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect -34 17 34 57
rect 410 57 427 91
rect 461 57 478 91
rect 1076 313 1144 353
rect 1742 427 1759 461
rect 1793 427 1810 461
rect 2186 461 2254 482
rect 1742 387 1810 427
rect 1742 353 1759 387
rect 1793 353 1810 387
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 410 17 478 57
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1742 313 1810 353
rect 2186 427 2203 461
rect 2237 427 2254 461
rect 2630 461 2698 482
rect 2186 387 2254 427
rect 2186 353 2203 387
rect 2237 353 2254 387
rect 2630 427 2647 461
rect 2681 427 2698 461
rect 3296 461 3364 482
rect 1742 279 1759 313
rect 1793 279 1810 313
rect 1742 239 1810 279
rect 1742 205 1759 239
rect 1793 205 1810 239
rect 1742 165 1810 205
rect 1742 131 1759 165
rect 1793 131 1810 165
rect 1742 91 1810 131
rect 1076 17 1144 57
rect 1742 57 1759 91
rect 1793 57 1810 91
rect 2186 313 2254 353
rect 2630 387 2698 427
rect 2630 353 2647 387
rect 2681 353 2698 387
rect 2186 279 2203 313
rect 2237 279 2254 313
rect 2186 239 2254 279
rect 2186 205 2203 239
rect 2237 205 2254 239
rect 2186 165 2254 205
rect 2186 131 2203 165
rect 2237 131 2254 165
rect 2186 91 2254 131
rect 1742 17 1810 57
rect 2186 57 2203 91
rect 2237 57 2254 91
rect 2630 313 2698 353
rect 3296 427 3313 461
rect 3347 427 3364 461
rect 3962 461 4030 482
rect 3296 387 3364 427
rect 3296 353 3313 387
rect 3347 353 3364 387
rect 2630 279 2647 313
rect 2681 279 2698 313
rect 2630 239 2698 279
rect 2630 205 2647 239
rect 2681 205 2698 239
rect 2630 165 2698 205
rect 2630 131 2647 165
rect 2681 131 2698 165
rect 2630 91 2698 131
rect 2186 17 2254 57
rect 2630 57 2647 91
rect 2681 57 2698 91
rect 3296 313 3364 353
rect 3962 427 3979 461
rect 4013 427 4030 461
rect 4406 461 4474 482
rect 3962 387 4030 427
rect 3962 353 3979 387
rect 4013 353 4030 387
rect 3296 279 3313 313
rect 3347 279 3364 313
rect 3296 239 3364 279
rect 3296 205 3313 239
rect 3347 205 3364 239
rect 3296 165 3364 205
rect 3296 131 3313 165
rect 3347 131 3364 165
rect 3296 91 3364 131
rect 2630 17 2698 57
rect 3296 57 3313 91
rect 3347 57 3364 91
rect 3962 313 4030 353
rect 4406 427 4423 461
rect 4457 427 4474 461
rect 5072 461 5140 482
rect 4406 387 4474 427
rect 4406 353 4423 387
rect 4457 353 4474 387
rect 3962 279 3979 313
rect 4013 279 4030 313
rect 3962 239 4030 279
rect 3962 205 3979 239
rect 4013 205 4030 239
rect 3962 165 4030 205
rect 3962 131 3979 165
rect 4013 131 4030 165
rect 3962 91 4030 131
rect 3296 17 3364 57
rect 3962 57 3979 91
rect 4013 57 4030 91
rect 4406 313 4474 353
rect 5072 427 5089 461
rect 5123 427 5140 461
rect 5516 461 5584 482
rect 5072 387 5140 427
rect 5072 353 5089 387
rect 5123 353 5140 387
rect 5516 427 5533 461
rect 5567 427 5584 461
rect 6182 461 6250 482
rect 4406 279 4423 313
rect 4457 279 4474 313
rect 4406 239 4474 279
rect 4406 205 4423 239
rect 4457 205 4474 239
rect 4406 165 4474 205
rect 4406 131 4423 165
rect 4457 131 4474 165
rect 4406 91 4474 131
rect 3962 17 4030 57
rect 4406 57 4423 91
rect 4457 57 4474 91
rect 5072 313 5140 353
rect 5516 387 5584 427
rect 5516 353 5533 387
rect 5567 353 5584 387
rect 5072 279 5089 313
rect 5123 279 5140 313
rect 5072 239 5140 279
rect 5072 205 5089 239
rect 5123 205 5140 239
rect 5072 165 5140 205
rect 5072 131 5089 165
rect 5123 131 5140 165
rect 5072 91 5140 131
rect 4406 17 4474 57
rect 5072 57 5089 91
rect 5123 57 5140 91
rect 5516 313 5584 353
rect 6182 427 6199 461
rect 6233 427 6250 461
rect 6626 461 6694 482
rect 6182 387 6250 427
rect 6182 353 6199 387
rect 6233 353 6250 387
rect 6626 427 6643 461
rect 6677 427 6694 461
rect 7292 461 7360 482
rect 5516 279 5533 313
rect 5567 279 5584 313
rect 5516 239 5584 279
rect 5516 205 5533 239
rect 5567 205 5584 239
rect 5516 165 5584 205
rect 5516 131 5533 165
rect 5567 131 5584 165
rect 5516 91 5584 131
rect 5072 17 5140 57
rect 5516 57 5533 91
rect 5567 57 5584 91
rect 6182 313 6250 353
rect 6626 387 6694 427
rect 6626 353 6643 387
rect 6677 353 6694 387
rect 6182 279 6199 313
rect 6233 279 6250 313
rect 6182 239 6250 279
rect 6182 205 6199 239
rect 6233 205 6250 239
rect 6182 165 6250 205
rect 6182 131 6199 165
rect 6233 131 6250 165
rect 6182 91 6250 131
rect 5516 17 5584 57
rect 6182 57 6199 91
rect 6233 57 6250 91
rect 6626 313 6694 353
rect 7292 427 7309 461
rect 7343 427 7360 461
rect 7736 461 7804 482
rect 7292 387 7360 427
rect 7292 353 7309 387
rect 7343 353 7360 387
rect 7736 427 7753 461
rect 7787 427 7804 461
rect 6626 279 6643 313
rect 6677 279 6694 313
rect 6626 239 6694 279
rect 6626 205 6643 239
rect 6677 205 6694 239
rect 6626 165 6694 205
rect 6626 131 6643 165
rect 6677 131 6694 165
rect 6626 91 6694 131
rect 6182 17 6250 57
rect 6626 57 6643 91
rect 6677 57 6694 91
rect 7292 313 7360 353
rect 7736 387 7804 427
rect 7736 353 7753 387
rect 7787 353 7804 387
rect 7292 279 7309 313
rect 7343 279 7360 313
rect 7292 239 7360 279
rect 7292 205 7309 239
rect 7343 205 7360 239
rect 7292 165 7360 205
rect 7292 131 7309 165
rect 7343 131 7360 165
rect 7292 91 7360 131
rect 6626 17 6694 57
rect 7292 57 7309 91
rect 7343 57 7360 91
rect 7736 313 7804 353
rect 7736 279 7753 313
rect 7787 279 7804 313
rect 7736 239 7804 279
rect 7736 205 7753 239
rect 7787 205 7804 239
rect 7736 165 7804 205
rect 7736 131 7753 165
rect 7787 131 7804 165
rect 7736 91 7804 131
rect 7292 17 7360 57
rect 7736 57 7753 91
rect 7787 57 7804 91
rect 7736 17 7804 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6569 17
rect 6603 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7804 17
rect -34 -34 7804 -17
<< nsubdiff >>
rect -34 1497 7804 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6569 1497
rect 6603 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7804 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 410 1423 478 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 1076 1423 1144 1463
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 410 979 478 1019
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1742 1423 1810 1463
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 410 945 427 979
rect 461 945 478 979
rect -34 871 -17 905
rect 17 884 34 905
rect 410 905 478 945
rect 1076 979 1144 1019
rect 1742 1389 1759 1423
rect 1793 1389 1810 1423
rect 2186 1423 2254 1463
rect 1742 1349 1810 1389
rect 1742 1315 1759 1349
rect 1793 1315 1810 1349
rect 1742 1275 1810 1315
rect 1742 1241 1759 1275
rect 1793 1241 1810 1275
rect 1742 1201 1810 1241
rect 1742 1167 1759 1201
rect 1793 1167 1810 1201
rect 1742 1127 1810 1167
rect 1742 1093 1759 1127
rect 1793 1093 1810 1127
rect 1742 1053 1810 1093
rect 1742 1019 1759 1053
rect 1793 1019 1810 1053
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 410 884 427 905
rect 17 871 427 884
rect 461 884 478 905
rect 1076 905 1144 945
rect 1742 979 1810 1019
rect 2186 1389 2203 1423
rect 2237 1389 2254 1423
rect 2630 1423 2698 1463
rect 2186 1349 2254 1389
rect 2186 1315 2203 1349
rect 2237 1315 2254 1349
rect 2186 1275 2254 1315
rect 2186 1241 2203 1275
rect 2237 1241 2254 1275
rect 2186 1201 2254 1241
rect 2186 1167 2203 1201
rect 2237 1167 2254 1201
rect 2186 1127 2254 1167
rect 2186 1093 2203 1127
rect 2237 1093 2254 1127
rect 2186 1053 2254 1093
rect 2186 1019 2203 1053
rect 2237 1019 2254 1053
rect 1742 945 1759 979
rect 1793 945 1810 979
rect 1076 884 1093 905
rect 461 871 1093 884
rect 1127 884 1144 905
rect 1742 905 1810 945
rect 2186 979 2254 1019
rect 2630 1389 2647 1423
rect 2681 1389 2698 1423
rect 3296 1423 3364 1463
rect 2630 1349 2698 1389
rect 2630 1315 2647 1349
rect 2681 1315 2698 1349
rect 2630 1275 2698 1315
rect 2630 1241 2647 1275
rect 2681 1241 2698 1275
rect 2630 1201 2698 1241
rect 2630 1167 2647 1201
rect 2681 1167 2698 1201
rect 2630 1127 2698 1167
rect 2630 1093 2647 1127
rect 2681 1093 2698 1127
rect 2630 1053 2698 1093
rect 2630 1019 2647 1053
rect 2681 1019 2698 1053
rect 2186 945 2203 979
rect 2237 945 2254 979
rect 1742 884 1759 905
rect 1127 871 1759 884
rect 1793 884 1810 905
rect 2186 905 2254 945
rect 2630 979 2698 1019
rect 3296 1389 3313 1423
rect 3347 1389 3364 1423
rect 3962 1423 4030 1463
rect 3296 1349 3364 1389
rect 3296 1315 3313 1349
rect 3347 1315 3364 1349
rect 3296 1275 3364 1315
rect 3296 1241 3313 1275
rect 3347 1241 3364 1275
rect 3296 1201 3364 1241
rect 3296 1167 3313 1201
rect 3347 1167 3364 1201
rect 3296 1127 3364 1167
rect 3296 1093 3313 1127
rect 3347 1093 3364 1127
rect 3296 1053 3364 1093
rect 3296 1019 3313 1053
rect 3347 1019 3364 1053
rect 2630 945 2647 979
rect 2681 945 2698 979
rect 2186 884 2203 905
rect 1793 871 2203 884
rect 2237 884 2254 905
rect 2630 905 2698 945
rect 3296 979 3364 1019
rect 3962 1389 3979 1423
rect 4013 1389 4030 1423
rect 4406 1423 4474 1463
rect 3962 1349 4030 1389
rect 3962 1315 3979 1349
rect 4013 1315 4030 1349
rect 3962 1275 4030 1315
rect 3962 1241 3979 1275
rect 4013 1241 4030 1275
rect 3962 1201 4030 1241
rect 3962 1167 3979 1201
rect 4013 1167 4030 1201
rect 3962 1127 4030 1167
rect 3962 1093 3979 1127
rect 4013 1093 4030 1127
rect 3962 1053 4030 1093
rect 3962 1019 3979 1053
rect 4013 1019 4030 1053
rect 3296 945 3313 979
rect 3347 945 3364 979
rect 2630 884 2647 905
rect 2237 871 2647 884
rect 2681 884 2698 905
rect 3296 905 3364 945
rect 3962 979 4030 1019
rect 4406 1389 4423 1423
rect 4457 1389 4474 1423
rect 5072 1423 5140 1463
rect 4406 1349 4474 1389
rect 4406 1315 4423 1349
rect 4457 1315 4474 1349
rect 4406 1275 4474 1315
rect 4406 1241 4423 1275
rect 4457 1241 4474 1275
rect 4406 1201 4474 1241
rect 4406 1167 4423 1201
rect 4457 1167 4474 1201
rect 4406 1127 4474 1167
rect 4406 1093 4423 1127
rect 4457 1093 4474 1127
rect 4406 1053 4474 1093
rect 4406 1019 4423 1053
rect 4457 1019 4474 1053
rect 3962 945 3979 979
rect 4013 945 4030 979
rect 3296 884 3313 905
rect 2681 871 3313 884
rect 3347 884 3364 905
rect 3962 905 4030 945
rect 4406 979 4474 1019
rect 5072 1389 5089 1423
rect 5123 1389 5140 1423
rect 5516 1423 5584 1463
rect 5072 1349 5140 1389
rect 5072 1315 5089 1349
rect 5123 1315 5140 1349
rect 5072 1275 5140 1315
rect 5072 1241 5089 1275
rect 5123 1241 5140 1275
rect 5072 1201 5140 1241
rect 5072 1167 5089 1201
rect 5123 1167 5140 1201
rect 5072 1127 5140 1167
rect 5072 1093 5089 1127
rect 5123 1093 5140 1127
rect 5072 1053 5140 1093
rect 5072 1019 5089 1053
rect 5123 1019 5140 1053
rect 4406 945 4423 979
rect 4457 945 4474 979
rect 3962 884 3979 905
rect 3347 871 3979 884
rect 4013 884 4030 905
rect 4406 905 4474 945
rect 5072 979 5140 1019
rect 5516 1389 5533 1423
rect 5567 1389 5584 1423
rect 6182 1423 6250 1463
rect 5516 1349 5584 1389
rect 5516 1315 5533 1349
rect 5567 1315 5584 1349
rect 5516 1275 5584 1315
rect 5516 1241 5533 1275
rect 5567 1241 5584 1275
rect 5516 1201 5584 1241
rect 5516 1167 5533 1201
rect 5567 1167 5584 1201
rect 5516 1127 5584 1167
rect 5516 1093 5533 1127
rect 5567 1093 5584 1127
rect 5516 1053 5584 1093
rect 5516 1019 5533 1053
rect 5567 1019 5584 1053
rect 5072 945 5089 979
rect 5123 945 5140 979
rect 4406 884 4423 905
rect 4013 871 4423 884
rect 4457 884 4474 905
rect 5072 905 5140 945
rect 5516 979 5584 1019
rect 6182 1389 6199 1423
rect 6233 1389 6250 1423
rect 6626 1423 6694 1463
rect 6182 1349 6250 1389
rect 6182 1315 6199 1349
rect 6233 1315 6250 1349
rect 6182 1275 6250 1315
rect 6182 1241 6199 1275
rect 6233 1241 6250 1275
rect 6182 1201 6250 1241
rect 6182 1167 6199 1201
rect 6233 1167 6250 1201
rect 6182 1127 6250 1167
rect 6182 1093 6199 1127
rect 6233 1093 6250 1127
rect 6182 1053 6250 1093
rect 6182 1019 6199 1053
rect 6233 1019 6250 1053
rect 5516 945 5533 979
rect 5567 945 5584 979
rect 5072 884 5089 905
rect 4457 871 5089 884
rect 5123 884 5140 905
rect 5516 905 5584 945
rect 6182 979 6250 1019
rect 6626 1389 6643 1423
rect 6677 1389 6694 1423
rect 7292 1423 7360 1463
rect 6626 1349 6694 1389
rect 6626 1315 6643 1349
rect 6677 1315 6694 1349
rect 6626 1275 6694 1315
rect 6626 1241 6643 1275
rect 6677 1241 6694 1275
rect 6626 1201 6694 1241
rect 6626 1167 6643 1201
rect 6677 1167 6694 1201
rect 6626 1127 6694 1167
rect 6626 1093 6643 1127
rect 6677 1093 6694 1127
rect 6626 1053 6694 1093
rect 6626 1019 6643 1053
rect 6677 1019 6694 1053
rect 6182 945 6199 979
rect 6233 945 6250 979
rect 5516 884 5533 905
rect 5123 871 5533 884
rect 5567 884 5584 905
rect 6182 905 6250 945
rect 6626 979 6694 1019
rect 7292 1389 7309 1423
rect 7343 1389 7360 1423
rect 7736 1423 7804 1463
rect 7292 1349 7360 1389
rect 7292 1315 7309 1349
rect 7343 1315 7360 1349
rect 7292 1275 7360 1315
rect 7292 1241 7309 1275
rect 7343 1241 7360 1275
rect 7292 1201 7360 1241
rect 7292 1167 7309 1201
rect 7343 1167 7360 1201
rect 7292 1127 7360 1167
rect 7292 1093 7309 1127
rect 7343 1093 7360 1127
rect 7292 1053 7360 1093
rect 7292 1019 7309 1053
rect 7343 1019 7360 1053
rect 6626 945 6643 979
rect 6677 945 6694 979
rect 6182 884 6199 905
rect 5567 871 6199 884
rect 6233 884 6250 905
rect 6626 905 6694 945
rect 7292 979 7360 1019
rect 7736 1389 7753 1423
rect 7787 1389 7804 1423
rect 7736 1349 7804 1389
rect 7736 1315 7753 1349
rect 7787 1315 7804 1349
rect 7736 1275 7804 1315
rect 7736 1241 7753 1275
rect 7787 1241 7804 1275
rect 7736 1201 7804 1241
rect 7736 1167 7753 1201
rect 7787 1167 7804 1201
rect 7736 1127 7804 1167
rect 7736 1093 7753 1127
rect 7787 1093 7804 1127
rect 7736 1053 7804 1093
rect 7736 1019 7753 1053
rect 7787 1019 7804 1053
rect 7292 945 7309 979
rect 7343 945 7360 979
rect 6626 884 6643 905
rect 6233 871 6643 884
rect 6677 884 6694 905
rect 7292 905 7360 945
rect 7736 979 7804 1019
rect 7736 945 7753 979
rect 7787 945 7804 979
rect 7292 884 7309 905
rect 6677 871 7309 884
rect 7343 884 7360 905
rect 7736 905 7804 945
rect 7736 884 7753 905
rect 7343 871 7753 884
rect 7787 871 7804 905
rect -34 822 7804 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 427 427 461 461
rect 427 353 461 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1093 427 1127 461
rect 1093 353 1127 387
rect 427 279 461 313
rect 427 205 461 239
rect 427 131 461 165
rect 427 57 461 91
rect 1759 427 1793 461
rect 1759 353 1793 387
rect 1093 279 1127 313
rect 1093 205 1127 239
rect 1093 131 1127 165
rect 1093 57 1127 91
rect 2203 427 2237 461
rect 2203 353 2237 387
rect 2647 427 2681 461
rect 1759 279 1793 313
rect 1759 205 1793 239
rect 1759 131 1793 165
rect 1759 57 1793 91
rect 2647 353 2681 387
rect 2203 279 2237 313
rect 2203 205 2237 239
rect 2203 131 2237 165
rect 2203 57 2237 91
rect 3313 427 3347 461
rect 3313 353 3347 387
rect 2647 279 2681 313
rect 2647 205 2681 239
rect 2647 131 2681 165
rect 2647 57 2681 91
rect 3979 427 4013 461
rect 3979 353 4013 387
rect 3313 279 3347 313
rect 3313 205 3347 239
rect 3313 131 3347 165
rect 3313 57 3347 91
rect 4423 427 4457 461
rect 4423 353 4457 387
rect 3979 279 4013 313
rect 3979 205 4013 239
rect 3979 131 4013 165
rect 3979 57 4013 91
rect 5089 427 5123 461
rect 5089 353 5123 387
rect 5533 427 5567 461
rect 4423 279 4457 313
rect 4423 205 4457 239
rect 4423 131 4457 165
rect 4423 57 4457 91
rect 5533 353 5567 387
rect 5089 279 5123 313
rect 5089 205 5123 239
rect 5089 131 5123 165
rect 5089 57 5123 91
rect 6199 427 6233 461
rect 6199 353 6233 387
rect 6643 427 6677 461
rect 5533 279 5567 313
rect 5533 205 5567 239
rect 5533 131 5567 165
rect 5533 57 5567 91
rect 6643 353 6677 387
rect 6199 279 6233 313
rect 6199 205 6233 239
rect 6199 131 6233 165
rect 6199 57 6233 91
rect 7309 427 7343 461
rect 7309 353 7343 387
rect 7753 427 7787 461
rect 6643 279 6677 313
rect 6643 205 6677 239
rect 6643 131 6677 165
rect 6643 57 6677 91
rect 7753 353 7787 387
rect 7309 279 7343 313
rect 7309 205 7343 239
rect 7309 131 7343 165
rect 7309 57 7343 91
rect 7753 279 7787 313
rect 7753 205 7787 239
rect 7753 131 7787 165
rect 7753 57 7787 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5163 -17 5197 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5755 -17 5789 17
rect 5829 -17 5863 17
rect 5903 -17 5937 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6125 -17 6159 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6495 -17 6529 17
rect 6569 -17 6603 17
rect 6717 -17 6751 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7087 -17 7121 17
rect 7161 -17 7195 17
rect 7235 -17 7269 17
rect 7383 -17 7417 17
rect 7457 -17 7491 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7679 -17 7713 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5163 1463 5197 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5755 1463 5789 1497
rect 5829 1463 5863 1497
rect 5903 1463 5937 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6125 1463 6159 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6495 1463 6529 1497
rect 6569 1463 6603 1497
rect 6717 1463 6751 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7087 1463 7121 1497
rect 7161 1463 7195 1497
rect 7235 1463 7269 1497
rect 7383 1463 7417 1497
rect 7457 1463 7491 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7679 1463 7713 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 427 1389 461 1423
rect 427 1315 461 1349
rect 427 1241 461 1275
rect 427 1167 461 1201
rect 427 1093 461 1127
rect 427 1019 461 1053
rect -17 945 17 979
rect 1093 1389 1127 1423
rect 1093 1315 1127 1349
rect 1093 1241 1127 1275
rect 1093 1167 1127 1201
rect 1093 1093 1127 1127
rect 1093 1019 1127 1053
rect 427 945 461 979
rect -17 871 17 905
rect 1759 1389 1793 1423
rect 1759 1315 1793 1349
rect 1759 1241 1793 1275
rect 1759 1167 1793 1201
rect 1759 1093 1793 1127
rect 1759 1019 1793 1053
rect 1093 945 1127 979
rect 427 871 461 905
rect 2203 1389 2237 1423
rect 2203 1315 2237 1349
rect 2203 1241 2237 1275
rect 2203 1167 2237 1201
rect 2203 1093 2237 1127
rect 2203 1019 2237 1053
rect 1759 945 1793 979
rect 1093 871 1127 905
rect 2647 1389 2681 1423
rect 2647 1315 2681 1349
rect 2647 1241 2681 1275
rect 2647 1167 2681 1201
rect 2647 1093 2681 1127
rect 2647 1019 2681 1053
rect 2203 945 2237 979
rect 1759 871 1793 905
rect 3313 1389 3347 1423
rect 3313 1315 3347 1349
rect 3313 1241 3347 1275
rect 3313 1167 3347 1201
rect 3313 1093 3347 1127
rect 3313 1019 3347 1053
rect 2647 945 2681 979
rect 2203 871 2237 905
rect 3979 1389 4013 1423
rect 3979 1315 4013 1349
rect 3979 1241 4013 1275
rect 3979 1167 4013 1201
rect 3979 1093 4013 1127
rect 3979 1019 4013 1053
rect 3313 945 3347 979
rect 2647 871 2681 905
rect 4423 1389 4457 1423
rect 4423 1315 4457 1349
rect 4423 1241 4457 1275
rect 4423 1167 4457 1201
rect 4423 1093 4457 1127
rect 4423 1019 4457 1053
rect 3979 945 4013 979
rect 3313 871 3347 905
rect 5089 1389 5123 1423
rect 5089 1315 5123 1349
rect 5089 1241 5123 1275
rect 5089 1167 5123 1201
rect 5089 1093 5123 1127
rect 5089 1019 5123 1053
rect 4423 945 4457 979
rect 3979 871 4013 905
rect 5533 1389 5567 1423
rect 5533 1315 5567 1349
rect 5533 1241 5567 1275
rect 5533 1167 5567 1201
rect 5533 1093 5567 1127
rect 5533 1019 5567 1053
rect 5089 945 5123 979
rect 4423 871 4457 905
rect 6199 1389 6233 1423
rect 6199 1315 6233 1349
rect 6199 1241 6233 1275
rect 6199 1167 6233 1201
rect 6199 1093 6233 1127
rect 6199 1019 6233 1053
rect 5533 945 5567 979
rect 5089 871 5123 905
rect 6643 1389 6677 1423
rect 6643 1315 6677 1349
rect 6643 1241 6677 1275
rect 6643 1167 6677 1201
rect 6643 1093 6677 1127
rect 6643 1019 6677 1053
rect 6199 945 6233 979
rect 5533 871 5567 905
rect 7309 1389 7343 1423
rect 7309 1315 7343 1349
rect 7309 1241 7343 1275
rect 7309 1167 7343 1201
rect 7309 1093 7343 1127
rect 7309 1019 7343 1053
rect 6643 945 6677 979
rect 6199 871 6233 905
rect 7753 1389 7787 1423
rect 7753 1315 7787 1349
rect 7753 1241 7787 1275
rect 7753 1167 7787 1201
rect 7753 1093 7787 1127
rect 7753 1019 7787 1053
rect 7309 945 7343 979
rect 6643 871 6677 905
rect 7753 945 7787 979
rect 7309 871 7343 905
rect 7753 871 7787 905
<< poly >>
rect 164 1404 194 1430
rect 252 1404 282 1430
rect 631 1404 661 1430
rect 719 1404 749 1430
rect 807 1404 837 1430
rect 895 1404 925 1430
rect 164 973 194 1004
rect 252 973 282 1004
rect 121 957 282 973
rect 121 923 131 957
rect 165 943 282 957
rect 1297 1404 1327 1430
rect 1385 1404 1415 1430
rect 1473 1404 1503 1430
rect 1561 1404 1591 1430
rect 165 923 175 943
rect 121 907 175 923
rect 631 973 661 1004
rect 719 973 749 1004
rect 631 957 749 973
rect 631 943 649 957
rect 639 923 649 943
rect 683 943 749 957
rect 807 973 837 1004
rect 895 973 925 1004
rect 807 957 925 973
rect 807 943 871 957
rect 683 923 693 943
rect 639 907 693 923
rect 861 923 871 943
rect 905 943 925 957
rect 1938 1404 1968 1430
rect 2026 1404 2056 1430
rect 905 923 915 943
rect 861 907 915 923
rect 1297 973 1327 1004
rect 1385 973 1415 1004
rect 1297 957 1415 973
rect 1297 943 1315 957
rect 1305 923 1315 943
rect 1349 943 1415 957
rect 1473 973 1503 1004
rect 1561 973 1591 1004
rect 1473 957 1591 973
rect 1473 943 1537 957
rect 1349 923 1359 943
rect 1305 907 1359 923
rect 1527 923 1537 943
rect 1571 943 1591 957
rect 2384 1404 2414 1430
rect 2472 1404 2502 1430
rect 1571 923 1581 943
rect 1527 907 1581 923
rect 1938 973 1968 1004
rect 2026 973 2056 1004
rect 2851 1404 2881 1430
rect 2939 1404 2969 1430
rect 3027 1404 3057 1430
rect 3115 1404 3145 1430
rect 1938 957 2099 973
rect 1938 943 2055 957
rect 2045 923 2055 943
rect 2089 923 2099 957
rect 2045 907 2099 923
rect 2384 973 2414 1004
rect 2472 973 2502 1004
rect 2341 957 2502 973
rect 2341 923 2351 957
rect 2385 943 2502 957
rect 3517 1404 3547 1430
rect 3605 1404 3635 1430
rect 3693 1404 3723 1430
rect 3781 1404 3811 1430
rect 2385 923 2395 943
rect 2341 907 2395 923
rect 2851 973 2881 1004
rect 2939 973 2969 1004
rect 2851 957 2969 973
rect 2851 943 2869 957
rect 2859 923 2869 943
rect 2903 943 2969 957
rect 3027 973 3057 1004
rect 3115 973 3145 1004
rect 3027 957 3145 973
rect 3027 943 3091 957
rect 2903 923 2913 943
rect 2859 907 2913 923
rect 3081 923 3091 943
rect 3125 943 3145 957
rect 4158 1404 4188 1430
rect 4246 1404 4276 1430
rect 3125 923 3135 943
rect 3081 907 3135 923
rect 3517 973 3547 1004
rect 3605 973 3635 1004
rect 3517 957 3635 973
rect 3517 943 3535 957
rect 3525 923 3535 943
rect 3569 943 3635 957
rect 3693 973 3723 1004
rect 3781 973 3811 1004
rect 3693 957 3811 973
rect 3693 943 3757 957
rect 3569 923 3579 943
rect 3525 907 3579 923
rect 3747 923 3757 943
rect 3791 943 3811 957
rect 4627 1404 4657 1430
rect 4715 1404 4745 1430
rect 4803 1404 4833 1430
rect 4891 1404 4921 1430
rect 3791 923 3801 943
rect 3747 907 3801 923
rect 4158 973 4188 1004
rect 4246 973 4276 1004
rect 5270 1404 5300 1430
rect 5358 1404 5388 1430
rect 4158 957 4319 973
rect 4158 943 4275 957
rect 4265 923 4275 943
rect 4309 923 4319 957
rect 4265 907 4319 923
rect 4627 973 4657 1004
rect 4715 973 4745 1004
rect 4803 973 4833 1004
rect 4891 973 4921 1004
rect 4627 957 4745 973
rect 4627 943 4645 957
rect 4635 923 4645 943
rect 4679 943 4745 957
rect 4789 957 4921 973
rect 4679 923 4689 943
rect 4635 907 4689 923
rect 4789 923 4799 957
rect 4833 943 4921 957
rect 5737 1404 5767 1430
rect 5825 1404 5855 1430
rect 5913 1404 5943 1430
rect 6001 1404 6031 1430
rect 5270 973 5300 1004
rect 5358 973 5388 1004
rect 4833 923 4843 943
rect 4789 907 4843 923
rect 5227 957 5388 973
rect 5227 923 5237 957
rect 5271 943 5388 957
rect 6380 1404 6410 1430
rect 6468 1404 6498 1430
rect 5271 923 5281 943
rect 5227 907 5281 923
rect 5737 973 5767 1004
rect 5825 973 5855 1004
rect 5913 973 5943 1004
rect 6001 973 6031 1004
rect 5737 957 5855 973
rect 5737 943 5755 957
rect 5745 923 5755 943
rect 5789 943 5855 957
rect 5899 957 6031 973
rect 5789 923 5799 943
rect 5745 907 5799 923
rect 5899 923 5909 957
rect 5943 943 6031 957
rect 6847 1405 6877 1431
rect 6935 1405 6965 1431
rect 7023 1405 7053 1431
rect 7111 1405 7141 1431
rect 6380 973 6410 1004
rect 6468 973 6498 1004
rect 5943 923 5953 943
rect 5899 907 5953 923
rect 6337 957 6498 973
rect 6337 923 6347 957
rect 6381 943 6498 957
rect 7490 1404 7520 1430
rect 7578 1404 7608 1430
rect 6847 974 6877 1005
rect 6935 974 6965 1005
rect 7023 974 7053 1005
rect 7111 974 7141 1005
rect 6381 923 6391 943
rect 6337 907 6391 923
rect 6824 958 6965 974
rect 6824 924 6834 958
rect 6868 944 6965 958
rect 7010 958 7141 974
rect 6868 924 6878 944
rect 6824 908 6878 924
rect 7010 924 7020 958
rect 7054 944 7141 958
rect 7490 973 7520 1004
rect 7578 973 7608 1004
rect 7054 924 7064 944
rect 7010 908 7064 924
rect 7447 957 7608 973
rect 7447 923 7457 957
rect 7491 943 7608 957
rect 7491 923 7501 943
rect 7447 907 7501 923
rect 121 434 175 450
rect 121 400 131 434
rect 165 413 175 434
rect 165 400 185 413
rect 121 384 185 400
rect 155 350 185 384
rect 639 434 693 450
rect 639 414 649 434
rect 612 400 649 414
rect 683 400 693 434
rect 861 434 915 450
rect 861 414 871 434
rect 612 384 693 400
rect 806 400 871 414
rect 905 400 915 434
rect 806 384 915 400
rect 1305 434 1359 450
rect 1305 414 1315 434
rect 612 350 642 384
rect 806 350 836 384
rect 1278 400 1315 414
rect 1349 400 1359 434
rect 1527 434 1581 450
rect 1527 414 1537 434
rect 1278 384 1359 400
rect 1472 400 1537 414
rect 1571 400 1581 434
rect 1472 384 1581 400
rect 2045 434 2099 450
rect 2045 413 2055 434
rect 1278 350 1308 384
rect 1472 350 1502 384
rect 2035 400 2055 413
rect 2089 400 2099 434
rect 2035 384 2099 400
rect 2035 350 2065 384
rect 2341 434 2395 450
rect 2341 400 2351 434
rect 2385 413 2395 434
rect 2385 400 2405 413
rect 2341 384 2405 400
rect 2375 350 2405 384
rect 2859 434 2913 450
rect 2859 414 2869 434
rect 2832 400 2869 414
rect 2903 400 2913 434
rect 3081 434 3135 450
rect 3081 414 3091 434
rect 2832 384 2913 400
rect 3026 400 3091 414
rect 3125 400 3135 434
rect 3026 384 3135 400
rect 3525 434 3579 450
rect 3525 414 3535 434
rect 2832 350 2862 384
rect 3026 350 3056 384
rect 3498 400 3535 414
rect 3569 400 3579 434
rect 3747 434 3801 450
rect 3747 414 3757 434
rect 3498 384 3579 400
rect 3692 400 3757 414
rect 3791 400 3801 434
rect 3692 384 3801 400
rect 4265 434 4319 450
rect 4265 413 4275 434
rect 3498 350 3528 384
rect 3692 350 3722 384
rect 4255 400 4275 413
rect 4309 400 4319 434
rect 4255 384 4319 400
rect 4635 433 4689 449
rect 4635 413 4645 433
rect 4255 350 4285 384
rect 4608 399 4645 413
rect 4679 399 4689 433
rect 4608 383 4689 399
rect 4783 433 4837 449
rect 4783 399 4793 433
rect 4827 399 4837 433
rect 4783 383 4837 399
rect 4608 349 4638 383
rect 4802 349 4832 383
rect 5227 434 5281 450
rect 5227 400 5237 434
rect 5271 413 5281 434
rect 5271 400 5291 413
rect 5227 384 5291 400
rect 5261 350 5291 384
rect 5745 433 5799 449
rect 5745 413 5755 433
rect 5718 399 5755 413
rect 5789 399 5799 433
rect 5718 383 5799 399
rect 5893 433 5947 449
rect 5893 399 5903 433
rect 5937 399 5947 433
rect 5893 383 5947 399
rect 5718 349 5748 383
rect 5912 349 5942 383
rect 6337 434 6391 450
rect 6337 400 6347 434
rect 6381 413 6391 434
rect 6381 400 6401 413
rect 6337 384 6401 400
rect 6371 350 6401 384
rect 6855 433 6909 449
rect 6855 413 6865 433
rect 6828 399 6865 413
rect 6899 399 6909 433
rect 6828 383 6909 399
rect 7003 433 7057 449
rect 7003 399 7013 433
rect 7047 399 7057 433
rect 7003 383 7057 399
rect 6828 349 6858 383
rect 7022 349 7052 383
rect 7447 434 7501 450
rect 7447 400 7457 434
rect 7491 413 7501 434
rect 7491 400 7511 413
rect 7447 384 7511 400
rect 7481 350 7511 384
<< polycont >>
rect 131 923 165 957
rect 649 923 683 957
rect 871 923 905 957
rect 1315 923 1349 957
rect 1537 923 1571 957
rect 2055 923 2089 957
rect 2351 923 2385 957
rect 2869 923 2903 957
rect 3091 923 3125 957
rect 3535 923 3569 957
rect 3757 923 3791 957
rect 4275 923 4309 957
rect 4645 923 4679 957
rect 4799 923 4833 957
rect 5237 923 5271 957
rect 5755 923 5789 957
rect 5909 923 5943 957
rect 6347 923 6381 957
rect 6834 924 6868 958
rect 7020 924 7054 958
rect 7457 923 7491 957
rect 131 400 165 434
rect 649 400 683 434
rect 871 400 905 434
rect 1315 400 1349 434
rect 1537 400 1571 434
rect 2055 400 2089 434
rect 2351 400 2385 434
rect 2869 400 2903 434
rect 3091 400 3125 434
rect 3535 400 3569 434
rect 3757 400 3791 434
rect 4275 400 4309 434
rect 4645 399 4679 433
rect 4793 399 4827 433
rect 5237 400 5271 434
rect 5755 399 5789 433
rect 5903 399 5937 433
rect 6347 400 6381 434
rect 6865 399 6899 433
rect 7013 399 7047 433
rect 7457 400 7491 434
<< locali >>
rect -34 1497 7804 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6569 1497
rect 6603 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7804 1497
rect -34 1446 7804 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 118 1366 152 1446
rect 118 1298 152 1332
rect 118 1230 152 1264
rect 118 1162 152 1196
rect 118 1093 152 1128
rect 118 1037 152 1059
rect 206 1366 240 1404
rect 206 1298 240 1332
rect 206 1230 240 1264
rect 206 1162 240 1196
rect 206 1093 240 1128
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 131 957 165 973
rect 131 831 165 923
rect 206 933 240 1059
rect 294 1366 328 1446
rect 294 1298 328 1332
rect 294 1230 328 1264
rect 294 1162 328 1196
rect 294 1093 328 1128
rect 294 1037 328 1059
rect 410 1423 478 1446
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect 585 1364 619 1380
rect 585 1296 619 1330
rect 585 1228 619 1262
rect 585 1160 619 1194
rect 585 1092 619 1126
rect 673 1296 707 1446
rect 1076 1423 1144 1446
rect 673 1228 707 1262
rect 673 1160 707 1194
rect 673 1110 707 1126
rect 761 1364 971 1398
rect 761 1296 795 1330
rect 761 1228 795 1262
rect 761 1160 795 1194
rect 761 1092 795 1126
rect 585 1024 795 1058
rect 849 1296 883 1312
rect 849 1228 883 1262
rect 849 1160 883 1194
rect 849 1092 883 1126
rect 937 1296 971 1330
rect 937 1228 971 1262
rect 937 1160 971 1194
rect 937 1110 971 1126
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 849 1024 979 1058
rect 410 979 478 1019
rect 410 945 427 979
rect 461 945 478 979
rect 206 899 313 933
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 131 434 165 797
rect 279 535 313 899
rect 410 905 478 945
rect 410 871 427 905
rect 461 871 478 905
rect 410 822 478 871
rect 649 957 683 973
rect 649 831 683 923
rect 279 433 313 501
rect 131 384 165 400
rect 205 399 313 433
rect 410 461 478 544
rect 649 461 683 797
rect 871 957 905 973
rect 871 831 905 923
rect 871 781 905 797
rect 945 757 979 1024
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 1251 1364 1285 1380
rect 1251 1296 1285 1330
rect 1251 1228 1285 1262
rect 1251 1160 1285 1194
rect 1251 1092 1285 1126
rect 1339 1296 1373 1446
rect 1742 1423 1810 1446
rect 1339 1228 1373 1262
rect 1339 1160 1373 1194
rect 1339 1110 1373 1126
rect 1427 1364 1637 1398
rect 1427 1296 1461 1330
rect 1427 1228 1461 1262
rect 1427 1160 1461 1194
rect 1427 1092 1461 1126
rect 1251 1024 1461 1058
rect 1515 1296 1549 1312
rect 1515 1228 1549 1262
rect 1515 1160 1549 1194
rect 1515 1092 1549 1126
rect 1603 1296 1637 1330
rect 1603 1228 1637 1262
rect 1603 1160 1637 1194
rect 1603 1110 1637 1126
rect 1742 1389 1759 1423
rect 1793 1389 1810 1423
rect 1742 1349 1810 1389
rect 1742 1315 1759 1349
rect 1793 1315 1810 1349
rect 1742 1275 1810 1315
rect 1742 1241 1759 1275
rect 1793 1241 1810 1275
rect 1742 1201 1810 1241
rect 1742 1167 1759 1201
rect 1793 1167 1810 1201
rect 1742 1127 1810 1167
rect 1742 1093 1759 1127
rect 1793 1093 1810 1127
rect 1515 1024 1645 1058
rect 1076 979 1144 1019
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 1076 905 1144 945
rect 1076 871 1093 905
rect 1127 871 1144 905
rect 1076 822 1144 871
rect 1315 957 1349 973
rect 1315 905 1349 923
rect 1315 855 1349 871
rect 1537 957 1571 973
rect 871 609 905 625
rect 410 427 427 461
rect 461 427 478 461
rect 633 427 649 461
rect 683 427 699 461
rect 871 434 905 575
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 109 334 143 350
rect 109 262 143 300
rect 109 194 143 228
rect 205 218 239 399
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect 649 384 683 400
rect 871 384 905 400
rect 205 168 239 184
rect 303 334 337 350
rect 303 262 337 300
rect 303 194 337 228
rect 109 124 143 160
rect 303 124 337 160
rect 143 90 205 124
rect 239 90 303 124
rect 109 34 143 90
rect 206 34 240 90
rect 303 34 337 90
rect 410 313 478 353
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect 410 57 427 91
rect 461 57 478 91
rect 566 334 600 350
rect 760 334 794 350
rect 945 348 979 723
rect 1315 683 1349 699
rect 600 300 663 334
rect 697 300 760 334
rect 566 262 600 300
rect 566 194 600 228
rect 760 262 794 300
rect 566 124 600 160
rect 566 74 600 90
rect 663 209 697 225
rect 410 34 478 57
rect 663 34 697 175
rect 760 194 794 228
rect 857 314 979 348
rect 1076 461 1144 544
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 1315 434 1349 649
rect 1315 384 1349 400
rect 1537 535 1571 923
rect 1537 434 1571 501
rect 1537 384 1571 400
rect 1611 757 1645 1024
rect 1742 1053 1810 1093
rect 1742 1019 1759 1053
rect 1793 1019 1810 1053
rect 1892 1366 1926 1446
rect 1892 1298 1926 1332
rect 1892 1230 1926 1264
rect 1892 1162 1926 1196
rect 1892 1093 1926 1128
rect 1892 1037 1926 1059
rect 1980 1366 2014 1404
rect 1980 1298 2014 1332
rect 1980 1230 2014 1264
rect 1980 1162 2014 1196
rect 1980 1093 2014 1128
rect 1742 979 1810 1019
rect 1742 945 1759 979
rect 1793 945 1810 979
rect 1742 905 1810 945
rect 1980 933 2014 1059
rect 2068 1366 2102 1446
rect 2068 1298 2102 1332
rect 2068 1230 2102 1264
rect 2068 1162 2102 1196
rect 2068 1093 2102 1128
rect 2068 1037 2102 1059
rect 2186 1423 2254 1446
rect 2186 1389 2203 1423
rect 2237 1389 2254 1423
rect 2186 1349 2254 1389
rect 2186 1315 2203 1349
rect 2237 1315 2254 1349
rect 2186 1275 2254 1315
rect 2186 1241 2203 1275
rect 2237 1241 2254 1275
rect 2186 1201 2254 1241
rect 2186 1167 2203 1201
rect 2237 1167 2254 1201
rect 2186 1127 2254 1167
rect 2186 1093 2203 1127
rect 2237 1093 2254 1127
rect 2186 1053 2254 1093
rect 2186 1019 2203 1053
rect 2237 1019 2254 1053
rect 2338 1366 2372 1446
rect 2338 1298 2372 1332
rect 2338 1230 2372 1264
rect 2338 1162 2372 1196
rect 2338 1093 2372 1128
rect 2338 1037 2372 1059
rect 2426 1366 2460 1404
rect 2426 1298 2460 1332
rect 2426 1230 2460 1264
rect 2426 1162 2460 1196
rect 2426 1093 2460 1128
rect 1742 871 1759 905
rect 1793 871 1810 905
rect 1742 822 1810 871
rect 1907 899 2014 933
rect 2055 979 2089 995
rect 2055 905 2089 923
rect 1907 831 1941 899
rect 857 218 891 314
rect 1076 313 1144 353
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 857 168 891 184
rect 954 262 988 278
rect 954 194 988 228
rect 760 124 794 160
rect 954 124 988 160
rect 794 90 857 124
rect 891 90 954 124
rect 760 74 794 90
rect 954 74 988 90
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1232 334 1266 350
rect 1426 334 1460 350
rect 1611 348 1645 723
rect 1907 683 1941 797
rect 1266 300 1329 334
rect 1363 300 1426 334
rect 1232 262 1266 300
rect 1232 194 1266 228
rect 1426 262 1460 300
rect 1232 124 1266 160
rect 1232 74 1266 90
rect 1329 209 1363 225
rect 1076 34 1144 57
rect 1329 34 1363 175
rect 1426 194 1460 228
rect 1523 314 1645 348
rect 1742 461 1810 544
rect 1742 427 1759 461
rect 1793 427 1810 461
rect 1742 387 1810 427
rect 1907 433 1941 649
rect 2055 609 2089 871
rect 2186 979 2254 1019
rect 2186 945 2203 979
rect 2237 945 2254 979
rect 2186 905 2254 945
rect 2186 871 2203 905
rect 2237 871 2254 905
rect 2186 822 2254 871
rect 2351 957 2385 973
rect 2351 831 2385 923
rect 2426 933 2460 1059
rect 2514 1366 2548 1446
rect 2514 1298 2548 1332
rect 2514 1230 2548 1264
rect 2514 1162 2548 1196
rect 2514 1093 2548 1128
rect 2514 1037 2548 1059
rect 2630 1423 2698 1446
rect 2630 1389 2647 1423
rect 2681 1389 2698 1423
rect 2630 1349 2698 1389
rect 2630 1315 2647 1349
rect 2681 1315 2698 1349
rect 2630 1275 2698 1315
rect 2630 1241 2647 1275
rect 2681 1241 2698 1275
rect 2630 1201 2698 1241
rect 2630 1167 2647 1201
rect 2681 1167 2698 1201
rect 2630 1127 2698 1167
rect 2630 1093 2647 1127
rect 2681 1093 2698 1127
rect 2630 1053 2698 1093
rect 2630 1019 2647 1053
rect 2681 1019 2698 1053
rect 2805 1364 2839 1380
rect 2805 1296 2839 1330
rect 2805 1228 2839 1262
rect 2805 1160 2839 1194
rect 2805 1092 2839 1126
rect 2893 1296 2927 1446
rect 3296 1423 3364 1446
rect 2893 1228 2927 1262
rect 2893 1160 2927 1194
rect 2893 1110 2927 1126
rect 2981 1364 3191 1398
rect 2981 1296 3015 1330
rect 2981 1228 3015 1262
rect 2981 1160 3015 1194
rect 2981 1092 3015 1126
rect 2805 1024 3015 1058
rect 3069 1296 3103 1312
rect 3069 1228 3103 1262
rect 3069 1160 3103 1194
rect 3069 1092 3103 1126
rect 3157 1296 3191 1330
rect 3157 1228 3191 1262
rect 3157 1160 3191 1194
rect 3157 1110 3191 1126
rect 3296 1389 3313 1423
rect 3347 1389 3364 1423
rect 3296 1349 3364 1389
rect 3296 1315 3313 1349
rect 3347 1315 3364 1349
rect 3296 1275 3364 1315
rect 3296 1241 3313 1275
rect 3347 1241 3364 1275
rect 3296 1201 3364 1241
rect 3296 1167 3313 1201
rect 3347 1167 3364 1201
rect 3296 1127 3364 1167
rect 3296 1093 3313 1127
rect 3347 1093 3364 1127
rect 3069 1024 3199 1058
rect 2630 979 2698 1019
rect 2630 945 2647 979
rect 2681 945 2698 979
rect 2426 899 2533 933
rect 2055 434 2089 575
rect 2351 757 2385 797
rect 1907 399 2015 433
rect 1742 353 1759 387
rect 1793 353 1810 387
rect 1523 218 1557 314
rect 1742 313 1810 353
rect 1742 279 1759 313
rect 1793 279 1810 313
rect 1523 168 1557 184
rect 1620 262 1654 278
rect 1620 194 1654 228
rect 1426 124 1460 160
rect 1620 124 1654 160
rect 1460 90 1523 124
rect 1557 90 1620 124
rect 1426 74 1460 90
rect 1620 74 1654 90
rect 1742 239 1810 279
rect 1742 205 1759 239
rect 1793 205 1810 239
rect 1742 165 1810 205
rect 1742 131 1759 165
rect 1793 131 1810 165
rect 1742 91 1810 131
rect 1742 57 1759 91
rect 1793 57 1810 91
rect 1742 34 1810 57
rect 1883 334 1917 350
rect 1883 262 1917 300
rect 1883 194 1917 228
rect 1981 218 2015 399
rect 2055 384 2089 400
rect 2186 461 2254 544
rect 2186 427 2203 461
rect 2237 427 2254 461
rect 2186 387 2254 427
rect 2186 353 2203 387
rect 2237 353 2254 387
rect 2351 461 2385 723
rect 2499 535 2533 899
rect 2630 905 2698 945
rect 2630 871 2647 905
rect 2681 871 2698 905
rect 2630 822 2698 871
rect 2869 957 2903 973
rect 2869 831 2903 923
rect 2499 433 2533 501
rect 2351 384 2385 400
rect 2425 399 2533 433
rect 2630 461 2698 544
rect 2630 427 2647 461
rect 2681 427 2698 461
rect 1981 168 2015 184
rect 2077 334 2111 350
rect 2077 262 2111 300
rect 2077 194 2111 228
rect 1883 124 1917 160
rect 2077 124 2111 160
rect 1917 90 1981 124
rect 2015 90 2077 124
rect 1883 34 1917 90
rect 1980 34 2014 90
rect 2077 34 2111 90
rect 2186 313 2254 353
rect 2186 279 2203 313
rect 2237 279 2254 313
rect 2186 239 2254 279
rect 2186 205 2203 239
rect 2237 205 2254 239
rect 2186 165 2254 205
rect 2186 131 2203 165
rect 2237 131 2254 165
rect 2186 91 2254 131
rect 2186 57 2203 91
rect 2237 57 2254 91
rect 2186 34 2254 57
rect 2329 334 2363 350
rect 2329 262 2363 300
rect 2329 194 2363 228
rect 2425 218 2459 399
rect 2630 387 2698 427
rect 2630 353 2647 387
rect 2681 353 2698 387
rect 2869 434 2903 797
rect 3091 957 3125 973
rect 3091 831 3125 923
rect 3091 781 3125 797
rect 3165 757 3199 1024
rect 3296 1053 3364 1093
rect 3296 1019 3313 1053
rect 3347 1019 3364 1053
rect 3471 1364 3505 1380
rect 3471 1296 3505 1330
rect 3471 1228 3505 1262
rect 3471 1160 3505 1194
rect 3471 1092 3505 1126
rect 3559 1296 3593 1446
rect 3962 1423 4030 1446
rect 3559 1228 3593 1262
rect 3559 1160 3593 1194
rect 3559 1110 3593 1126
rect 3647 1364 3857 1398
rect 3647 1296 3681 1330
rect 3647 1228 3681 1262
rect 3647 1160 3681 1194
rect 3647 1092 3681 1126
rect 3471 1024 3681 1058
rect 3735 1296 3769 1312
rect 3735 1228 3769 1262
rect 3735 1160 3769 1194
rect 3735 1092 3769 1126
rect 3823 1296 3857 1330
rect 3823 1228 3857 1262
rect 3823 1160 3857 1194
rect 3823 1110 3857 1126
rect 3962 1389 3979 1423
rect 4013 1389 4030 1423
rect 3962 1349 4030 1389
rect 3962 1315 3979 1349
rect 4013 1315 4030 1349
rect 3962 1275 4030 1315
rect 3962 1241 3979 1275
rect 4013 1241 4030 1275
rect 3962 1201 4030 1241
rect 3962 1167 3979 1201
rect 4013 1167 4030 1201
rect 3962 1127 4030 1167
rect 3962 1093 3979 1127
rect 4013 1093 4030 1127
rect 3735 1024 3865 1058
rect 3296 979 3364 1019
rect 3296 945 3313 979
rect 3347 945 3364 979
rect 3296 905 3364 945
rect 3296 871 3313 905
rect 3347 871 3364 905
rect 3296 822 3364 871
rect 3535 957 3569 973
rect 3535 905 3569 923
rect 3535 855 3569 871
rect 3757 957 3791 973
rect 2869 384 2903 400
rect 3091 609 3125 625
rect 3091 434 3125 575
rect 3091 384 3125 400
rect 2425 168 2459 184
rect 2523 334 2557 350
rect 2523 262 2557 300
rect 2523 194 2557 228
rect 2329 124 2363 160
rect 2523 124 2557 160
rect 2363 90 2425 124
rect 2459 90 2523 124
rect 2329 34 2363 90
rect 2426 34 2460 90
rect 2523 34 2557 90
rect 2630 313 2698 353
rect 2630 279 2647 313
rect 2681 279 2698 313
rect 2630 239 2698 279
rect 2630 205 2647 239
rect 2681 205 2698 239
rect 2630 165 2698 205
rect 2630 131 2647 165
rect 2681 131 2698 165
rect 2630 91 2698 131
rect 2630 57 2647 91
rect 2681 57 2698 91
rect 2786 334 2820 350
rect 2980 334 3014 350
rect 3165 348 3199 723
rect 3535 683 3569 699
rect 2820 300 2883 334
rect 2917 300 2980 334
rect 2786 262 2820 300
rect 2786 194 2820 228
rect 2980 262 3014 300
rect 2786 124 2820 160
rect 2786 74 2820 90
rect 2883 209 2917 225
rect 2630 34 2698 57
rect 2883 34 2917 175
rect 2980 194 3014 228
rect 3077 314 3199 348
rect 3296 461 3364 544
rect 3296 427 3313 461
rect 3347 427 3364 461
rect 3296 387 3364 427
rect 3296 353 3313 387
rect 3347 353 3364 387
rect 3535 434 3569 649
rect 3535 384 3569 400
rect 3757 535 3791 923
rect 3757 434 3791 501
rect 3757 384 3791 400
rect 3831 757 3865 1024
rect 3962 1053 4030 1093
rect 3962 1019 3979 1053
rect 4013 1019 4030 1053
rect 4112 1366 4146 1446
rect 4112 1298 4146 1332
rect 4112 1230 4146 1264
rect 4112 1162 4146 1196
rect 4112 1093 4146 1128
rect 4112 1037 4146 1059
rect 4200 1366 4234 1404
rect 4200 1298 4234 1332
rect 4200 1230 4234 1264
rect 4200 1162 4234 1196
rect 4200 1093 4234 1128
rect 3962 979 4030 1019
rect 3962 945 3979 979
rect 4013 945 4030 979
rect 3962 905 4030 945
rect 4200 933 4234 1059
rect 4288 1366 4322 1446
rect 4288 1298 4322 1332
rect 4288 1230 4322 1264
rect 4288 1162 4322 1196
rect 4288 1093 4322 1128
rect 4288 1037 4322 1059
rect 4406 1423 4474 1446
rect 4406 1389 4423 1423
rect 4457 1389 4474 1423
rect 4406 1349 4474 1389
rect 4406 1315 4423 1349
rect 4457 1315 4474 1349
rect 4406 1275 4474 1315
rect 4406 1241 4423 1275
rect 4457 1241 4474 1275
rect 4406 1201 4474 1241
rect 4406 1167 4423 1201
rect 4457 1167 4474 1201
rect 4406 1127 4474 1167
rect 4406 1093 4423 1127
rect 4457 1093 4474 1127
rect 4406 1053 4474 1093
rect 4406 1019 4423 1053
rect 4457 1019 4474 1053
rect 4581 1366 4615 1446
rect 4581 1298 4615 1332
rect 4581 1230 4615 1264
rect 4581 1162 4615 1196
rect 4581 1093 4615 1128
rect 4581 1027 4615 1059
rect 4669 1366 4703 1404
rect 4669 1298 4703 1332
rect 4669 1230 4703 1264
rect 4669 1162 4703 1196
rect 4669 1093 4703 1128
rect 4757 1366 4791 1446
rect 4757 1298 4791 1332
rect 4757 1230 4791 1264
rect 4757 1162 4791 1196
rect 4757 1111 4791 1128
rect 4845 1366 4879 1404
rect 4845 1298 4879 1332
rect 4845 1230 4879 1264
rect 4845 1162 4879 1196
rect 4669 1057 4703 1059
rect 4845 1093 4879 1128
rect 4933 1366 4967 1446
rect 4933 1298 4967 1332
rect 4933 1230 4967 1264
rect 4933 1162 4967 1196
rect 4933 1111 4967 1128
rect 5072 1423 5140 1446
rect 5072 1389 5089 1423
rect 5123 1389 5140 1423
rect 5072 1349 5140 1389
rect 5072 1315 5089 1349
rect 5123 1315 5140 1349
rect 5072 1275 5140 1315
rect 5072 1241 5089 1275
rect 5123 1241 5140 1275
rect 5072 1201 5140 1241
rect 5072 1167 5089 1201
rect 5123 1167 5140 1201
rect 5072 1127 5140 1167
rect 4845 1057 4879 1059
rect 5072 1093 5089 1127
rect 5123 1093 5140 1127
rect 4669 1023 4975 1057
rect 4406 979 4474 1019
rect 3962 871 3979 905
rect 4013 871 4030 905
rect 3962 822 4030 871
rect 4127 899 4234 933
rect 4275 957 4309 973
rect 4275 905 4309 923
rect 4127 831 4161 899
rect 3077 218 3111 314
rect 3296 313 3364 353
rect 3296 279 3313 313
rect 3347 279 3364 313
rect 3077 168 3111 184
rect 3174 262 3208 278
rect 3174 194 3208 228
rect 2980 124 3014 160
rect 3174 124 3208 160
rect 3014 90 3077 124
rect 3111 90 3174 124
rect 2980 74 3014 90
rect 3174 74 3208 90
rect 3296 239 3364 279
rect 3296 205 3313 239
rect 3347 205 3364 239
rect 3296 165 3364 205
rect 3296 131 3313 165
rect 3347 131 3364 165
rect 3296 91 3364 131
rect 3296 57 3313 91
rect 3347 57 3364 91
rect 3452 334 3486 350
rect 3646 334 3680 350
rect 3831 348 3865 723
rect 4127 683 4161 797
rect 3486 300 3549 334
rect 3583 300 3646 334
rect 3452 262 3486 300
rect 3452 194 3486 228
rect 3646 262 3680 300
rect 3452 124 3486 160
rect 3452 74 3486 90
rect 3549 209 3583 225
rect 3296 34 3364 57
rect 3549 34 3583 175
rect 3646 194 3680 228
rect 3743 314 3865 348
rect 3962 461 4030 544
rect 3962 427 3979 461
rect 4013 427 4030 461
rect 3962 387 4030 427
rect 4127 433 4161 649
rect 4275 609 4309 871
rect 4406 945 4423 979
rect 4457 945 4474 979
rect 4406 905 4474 945
rect 4406 871 4423 905
rect 4457 871 4474 905
rect 4406 822 4474 871
rect 4645 957 4679 973
rect 4799 957 4833 973
rect 4645 905 4679 923
rect 4275 434 4309 575
rect 4127 399 4235 433
rect 3962 353 3979 387
rect 4013 353 4030 387
rect 3743 218 3777 314
rect 3962 313 4030 353
rect 3962 279 3979 313
rect 4013 279 4030 313
rect 3743 168 3777 184
rect 3840 262 3874 278
rect 3840 194 3874 228
rect 3646 124 3680 160
rect 3840 124 3874 160
rect 3680 90 3743 124
rect 3777 90 3840 124
rect 3646 74 3680 90
rect 3840 74 3874 90
rect 3962 239 4030 279
rect 3962 205 3979 239
rect 4013 205 4030 239
rect 3962 165 4030 205
rect 3962 131 3979 165
rect 4013 131 4030 165
rect 3962 91 4030 131
rect 3962 57 3979 91
rect 4013 57 4030 91
rect 3962 34 4030 57
rect 4103 334 4137 350
rect 4103 262 4137 300
rect 4103 194 4137 228
rect 4201 218 4235 399
rect 4275 384 4309 400
rect 4406 461 4474 544
rect 4406 427 4423 461
rect 4457 427 4474 461
rect 4406 387 4474 427
rect 4406 353 4423 387
rect 4457 353 4474 387
rect 4645 433 4679 871
rect 4645 383 4679 399
rect 4793 923 4799 942
rect 4793 907 4833 923
rect 4793 461 4827 907
rect 4793 383 4827 399
rect 4941 683 4975 1023
rect 5072 1053 5140 1093
rect 5072 1019 5089 1053
rect 5123 1019 5140 1053
rect 5224 1366 5258 1446
rect 5224 1298 5258 1332
rect 5224 1230 5258 1264
rect 5224 1162 5258 1196
rect 5224 1093 5258 1128
rect 5224 1037 5258 1059
rect 5312 1366 5346 1404
rect 5312 1298 5346 1332
rect 5312 1230 5346 1264
rect 5312 1162 5346 1196
rect 5312 1093 5346 1128
rect 5072 979 5140 1019
rect 5072 945 5089 979
rect 5123 945 5140 979
rect 5072 905 5140 945
rect 5072 871 5089 905
rect 5123 871 5140 905
rect 5072 822 5140 871
rect 5237 957 5271 973
rect 4201 168 4235 184
rect 4297 334 4331 350
rect 4297 262 4331 300
rect 4297 194 4331 228
rect 4103 124 4137 160
rect 4297 124 4331 160
rect 4137 90 4201 124
rect 4235 90 4297 124
rect 4103 34 4137 90
rect 4200 34 4234 90
rect 4297 34 4331 90
rect 4406 313 4474 353
rect 4406 279 4423 313
rect 4457 279 4474 313
rect 4406 239 4474 279
rect 4406 205 4423 239
rect 4457 205 4474 239
rect 4406 165 4474 205
rect 4406 131 4423 165
rect 4457 131 4474 165
rect 4406 91 4474 131
rect 4406 57 4423 91
rect 4457 57 4474 91
rect 4562 333 4596 349
rect 4756 333 4790 349
rect 4941 348 4975 649
rect 5237 683 5271 923
rect 5312 933 5346 1059
rect 5400 1366 5434 1446
rect 5400 1298 5434 1332
rect 5400 1230 5434 1264
rect 5400 1162 5434 1196
rect 5400 1093 5434 1128
rect 5400 1037 5434 1059
rect 5516 1423 5584 1446
rect 5516 1389 5533 1423
rect 5567 1389 5584 1423
rect 5516 1349 5584 1389
rect 5516 1315 5533 1349
rect 5567 1315 5584 1349
rect 5516 1275 5584 1315
rect 5516 1241 5533 1275
rect 5567 1241 5584 1275
rect 5516 1201 5584 1241
rect 5516 1167 5533 1201
rect 5567 1167 5584 1201
rect 5516 1127 5584 1167
rect 5516 1093 5533 1127
rect 5567 1093 5584 1127
rect 5516 1053 5584 1093
rect 5516 1019 5533 1053
rect 5567 1019 5584 1053
rect 5691 1366 5725 1446
rect 5691 1298 5725 1332
rect 5691 1230 5725 1264
rect 5691 1162 5725 1196
rect 5691 1093 5725 1128
rect 5691 1027 5725 1059
rect 5779 1366 5813 1404
rect 5779 1298 5813 1332
rect 5779 1230 5813 1264
rect 5779 1162 5813 1196
rect 5779 1093 5813 1128
rect 5867 1366 5901 1446
rect 5867 1298 5901 1332
rect 5867 1230 5901 1264
rect 5867 1162 5901 1196
rect 5867 1111 5901 1128
rect 5955 1366 5989 1404
rect 5955 1298 5989 1332
rect 5955 1230 5989 1264
rect 5955 1162 5989 1196
rect 5779 1057 5813 1059
rect 5955 1093 5989 1128
rect 6043 1366 6077 1446
rect 6043 1298 6077 1332
rect 6043 1230 6077 1264
rect 6043 1162 6077 1196
rect 6043 1111 6077 1128
rect 6182 1423 6250 1446
rect 6182 1389 6199 1423
rect 6233 1389 6250 1423
rect 6182 1349 6250 1389
rect 6182 1315 6199 1349
rect 6233 1315 6250 1349
rect 6182 1275 6250 1315
rect 6182 1241 6199 1275
rect 6233 1241 6250 1275
rect 6182 1201 6250 1241
rect 6182 1167 6199 1201
rect 6233 1167 6250 1201
rect 6182 1127 6250 1167
rect 5955 1057 5989 1059
rect 6182 1093 6199 1127
rect 6233 1093 6250 1127
rect 5779 1023 6085 1057
rect 5516 979 5584 1019
rect 5516 945 5533 979
rect 5567 945 5584 979
rect 5312 899 5419 933
rect 4596 299 4659 333
rect 4693 299 4756 333
rect 4562 261 4596 299
rect 4562 193 4596 227
rect 4756 261 4790 299
rect 4562 123 4596 159
rect 4562 73 4596 89
rect 4659 208 4693 224
rect 4406 34 4474 57
rect 4659 34 4693 174
rect 4756 193 4790 227
rect 4853 314 4975 348
rect 5072 461 5140 544
rect 5072 427 5089 461
rect 5123 427 5140 461
rect 5072 387 5140 427
rect 5072 353 5089 387
rect 5123 353 5140 387
rect 5237 434 5271 649
rect 5385 609 5419 899
rect 5516 905 5584 945
rect 5755 957 5789 979
rect 5909 957 5943 973
rect 5739 909 5755 943
rect 5789 909 5805 943
rect 5903 923 5909 942
rect 5516 871 5533 905
rect 5567 871 5584 905
rect 5516 822 5584 871
rect 5385 433 5419 575
rect 5237 384 5271 400
rect 5311 399 5419 433
rect 5516 461 5584 544
rect 5516 427 5533 461
rect 5567 427 5584 461
rect 4853 217 4887 314
rect 5072 313 5140 353
rect 5072 279 5089 313
rect 5123 279 5140 313
rect 4853 167 4887 183
rect 4950 261 4984 277
rect 4950 193 4984 227
rect 4756 123 4790 159
rect 4950 123 4984 159
rect 4790 89 4853 123
rect 4887 89 4950 123
rect 4756 73 4790 89
rect 4950 73 4984 89
rect 5072 239 5140 279
rect 5072 205 5089 239
rect 5123 205 5140 239
rect 5072 165 5140 205
rect 5072 131 5089 165
rect 5123 131 5140 165
rect 5072 91 5140 131
rect 5072 57 5089 91
rect 5123 57 5140 91
rect 5072 34 5140 57
rect 5215 334 5249 350
rect 5215 262 5249 300
rect 5215 194 5249 228
rect 5311 218 5345 399
rect 5516 387 5584 427
rect 5516 353 5533 387
rect 5567 353 5584 387
rect 5755 433 5789 909
rect 5903 907 5943 923
rect 5903 461 5937 907
rect 6051 683 6085 1023
rect 6182 1053 6250 1093
rect 6182 1019 6199 1053
rect 6233 1019 6250 1053
rect 6334 1366 6368 1446
rect 6334 1298 6368 1332
rect 6334 1230 6368 1264
rect 6334 1162 6368 1196
rect 6334 1093 6368 1128
rect 6334 1037 6368 1059
rect 6422 1366 6456 1404
rect 6422 1298 6456 1332
rect 6422 1230 6456 1264
rect 6422 1162 6456 1196
rect 6422 1093 6456 1128
rect 6182 979 6250 1019
rect 6182 945 6199 979
rect 6233 945 6250 979
rect 6182 905 6250 945
rect 6182 871 6199 905
rect 6233 871 6250 905
rect 6182 822 6250 871
rect 6347 957 6381 973
rect 5887 427 5903 461
rect 5937 427 5953 461
rect 5755 383 5789 399
rect 5903 383 5937 399
rect 5311 168 5345 184
rect 5409 334 5443 350
rect 5409 262 5443 300
rect 5409 194 5443 228
rect 5215 124 5249 160
rect 5409 124 5443 160
rect 5249 90 5311 124
rect 5345 90 5409 124
rect 5215 34 5249 90
rect 5312 34 5346 90
rect 5409 34 5443 90
rect 5516 313 5584 353
rect 5516 279 5533 313
rect 5567 279 5584 313
rect 5516 239 5584 279
rect 5516 205 5533 239
rect 5567 205 5584 239
rect 5516 165 5584 205
rect 5516 131 5533 165
rect 5567 131 5584 165
rect 5516 91 5584 131
rect 5516 57 5533 91
rect 5567 57 5584 91
rect 5672 333 5706 349
rect 5866 333 5900 349
rect 6051 348 6085 649
rect 6347 683 6381 923
rect 6422 933 6456 1059
rect 6510 1366 6544 1446
rect 6510 1298 6544 1332
rect 6510 1230 6544 1264
rect 6510 1162 6544 1196
rect 6510 1093 6544 1128
rect 6510 1037 6544 1059
rect 6626 1423 6694 1446
rect 6626 1389 6643 1423
rect 6677 1389 6694 1423
rect 6626 1349 6694 1389
rect 6626 1315 6643 1349
rect 6677 1315 6694 1349
rect 6626 1275 6694 1315
rect 6626 1241 6643 1275
rect 6677 1241 6694 1275
rect 6626 1201 6694 1241
rect 6626 1167 6643 1201
rect 6677 1167 6694 1201
rect 6626 1127 6694 1167
rect 6626 1093 6643 1127
rect 6677 1093 6694 1127
rect 6626 1053 6694 1093
rect 6626 1019 6643 1053
rect 6677 1019 6694 1053
rect 6801 1365 6835 1405
rect 6801 1297 6835 1331
rect 6801 1229 6835 1263
rect 6801 1161 6835 1195
rect 6801 1093 6835 1127
rect 6889 1365 6923 1446
rect 7292 1423 7360 1446
rect 6889 1297 6923 1331
rect 6889 1229 6923 1263
rect 6889 1161 6923 1195
rect 6889 1111 6923 1127
rect 6977 1365 7187 1399
rect 6977 1297 7011 1331
rect 6977 1229 7011 1263
rect 6977 1161 7011 1195
rect 6977 1093 7011 1127
rect 6801 1025 7011 1059
rect 7065 1297 7099 1313
rect 7065 1229 7099 1263
rect 7065 1161 7099 1195
rect 7065 1093 7099 1127
rect 7153 1297 7187 1331
rect 7153 1229 7187 1263
rect 7153 1161 7187 1195
rect 7153 1111 7187 1127
rect 7292 1389 7309 1423
rect 7343 1389 7360 1423
rect 7292 1349 7360 1389
rect 7292 1315 7309 1349
rect 7343 1315 7360 1349
rect 7292 1275 7360 1315
rect 7292 1241 7309 1275
rect 7343 1241 7360 1275
rect 7292 1201 7360 1241
rect 7292 1167 7309 1201
rect 7343 1167 7360 1201
rect 7292 1127 7360 1167
rect 7292 1093 7309 1127
rect 7343 1093 7360 1127
rect 7065 1025 7195 1059
rect 6626 979 6694 1019
rect 6626 945 6643 979
rect 6677 945 6694 979
rect 6422 899 6529 933
rect 5706 299 5769 333
rect 5803 299 5866 333
rect 5672 261 5706 299
rect 5672 193 5706 227
rect 5866 261 5900 299
rect 5672 123 5706 159
rect 5672 73 5706 89
rect 5769 208 5803 224
rect 5516 34 5584 57
rect 5769 34 5803 174
rect 5866 193 5900 227
rect 5963 314 6085 348
rect 6182 461 6250 544
rect 6182 427 6199 461
rect 6233 427 6250 461
rect 6182 387 6250 427
rect 6182 353 6199 387
rect 6233 353 6250 387
rect 6347 434 6381 649
rect 6495 683 6529 899
rect 6626 905 6694 945
rect 6834 958 6868 974
rect 7020 958 7054 974
rect 6868 924 6899 942
rect 6834 908 6899 924
rect 6626 871 6643 905
rect 6677 871 6694 905
rect 6626 822 6694 871
rect 6495 433 6529 649
rect 6865 609 6899 908
rect 6347 384 6381 400
rect 6421 399 6529 433
rect 6626 461 6694 544
rect 6626 427 6643 461
rect 6677 427 6694 461
rect 5963 217 5997 314
rect 6182 313 6250 353
rect 6182 279 6199 313
rect 6233 279 6250 313
rect 5963 167 5997 183
rect 6060 261 6094 277
rect 6060 193 6094 227
rect 5866 123 5900 159
rect 6060 123 6094 159
rect 5900 89 5963 123
rect 5997 89 6060 123
rect 5866 73 5900 89
rect 6060 73 6094 89
rect 6182 239 6250 279
rect 6182 205 6199 239
rect 6233 205 6250 239
rect 6182 165 6250 205
rect 6182 131 6199 165
rect 6233 131 6250 165
rect 6182 91 6250 131
rect 6182 57 6199 91
rect 6233 57 6250 91
rect 6182 34 6250 57
rect 6325 334 6359 350
rect 6325 262 6359 300
rect 6325 194 6359 228
rect 6421 218 6455 399
rect 6626 387 6694 427
rect 6626 353 6643 387
rect 6677 353 6694 387
rect 6865 433 6899 575
rect 6865 383 6899 399
rect 7013 924 7020 942
rect 7013 908 7054 924
rect 7013 683 7047 908
rect 7013 433 7047 649
rect 7013 383 7047 399
rect 7161 683 7195 1025
rect 7292 1053 7360 1093
rect 7292 1019 7309 1053
rect 7343 1019 7360 1053
rect 7444 1366 7478 1446
rect 7444 1298 7478 1332
rect 7444 1230 7478 1264
rect 7444 1162 7478 1196
rect 7444 1093 7478 1128
rect 7444 1037 7478 1059
rect 7532 1366 7566 1404
rect 7532 1298 7566 1332
rect 7532 1230 7566 1264
rect 7532 1162 7566 1196
rect 7532 1093 7566 1128
rect 7292 979 7360 1019
rect 7292 945 7309 979
rect 7343 945 7360 979
rect 7292 905 7360 945
rect 7292 871 7309 905
rect 7343 871 7360 905
rect 7292 822 7360 871
rect 7457 957 7491 973
rect 6421 168 6455 184
rect 6519 334 6553 350
rect 6519 262 6553 300
rect 6519 194 6553 228
rect 6325 124 6359 160
rect 6519 124 6553 160
rect 6359 90 6421 124
rect 6455 90 6519 124
rect 6325 34 6359 90
rect 6422 34 6456 90
rect 6519 34 6553 90
rect 6626 313 6694 353
rect 6626 279 6643 313
rect 6677 279 6694 313
rect 6626 239 6694 279
rect 6626 205 6643 239
rect 6677 205 6694 239
rect 6626 165 6694 205
rect 6626 131 6643 165
rect 6677 131 6694 165
rect 6626 91 6694 131
rect 6626 57 6643 91
rect 6677 57 6694 91
rect 6626 34 6694 57
rect 6782 333 6816 349
rect 7161 348 7195 649
rect 7457 683 7491 923
rect 7532 933 7566 1059
rect 7620 1366 7654 1446
rect 7620 1298 7654 1332
rect 7620 1230 7654 1264
rect 7620 1162 7654 1196
rect 7620 1093 7654 1128
rect 7620 1037 7654 1059
rect 7736 1423 7804 1446
rect 7736 1389 7753 1423
rect 7787 1389 7804 1423
rect 7736 1349 7804 1389
rect 7736 1315 7753 1349
rect 7787 1315 7804 1349
rect 7736 1275 7804 1315
rect 7736 1241 7753 1275
rect 7787 1241 7804 1275
rect 7736 1201 7804 1241
rect 7736 1167 7753 1201
rect 7787 1167 7804 1201
rect 7736 1127 7804 1167
rect 7736 1093 7753 1127
rect 7787 1093 7804 1127
rect 7736 1053 7804 1093
rect 7736 1019 7753 1053
rect 7787 1019 7804 1053
rect 7736 979 7804 1019
rect 7736 945 7753 979
rect 7787 945 7804 979
rect 7532 899 7639 933
rect 6782 261 6816 299
rect 6782 193 6816 227
rect 6879 314 7195 348
rect 7292 461 7360 544
rect 7292 427 7309 461
rect 7343 427 7360 461
rect 7292 387 7360 427
rect 7292 353 7309 387
rect 7343 353 7360 387
rect 7457 434 7491 649
rect 7605 433 7639 899
rect 7736 905 7804 945
rect 7736 871 7753 905
rect 7787 871 7804 905
rect 7736 822 7804 871
rect 7457 384 7491 400
rect 7531 399 7639 433
rect 7736 461 7804 544
rect 7736 427 7753 461
rect 7787 427 7804 461
rect 6879 217 6913 314
rect 6879 167 6913 183
rect 6976 261 7010 278
rect 6976 193 7010 227
rect 6782 123 6816 159
rect 7073 217 7107 314
rect 7292 313 7360 353
rect 7292 279 7309 313
rect 7343 279 7360 313
rect 7073 167 7107 183
rect 7170 261 7204 278
rect 7170 193 7204 227
rect 6976 123 7010 159
rect 7170 123 7204 159
rect 6816 89 6879 123
rect 6913 89 6976 123
rect 7010 89 7073 123
rect 7107 89 7170 123
rect 6782 34 6816 89
rect 6879 34 6913 89
rect 6976 34 7010 89
rect 7073 34 7107 89
rect 7170 34 7204 89
rect 7292 239 7360 279
rect 7292 205 7309 239
rect 7343 205 7360 239
rect 7292 165 7360 205
rect 7292 131 7309 165
rect 7343 131 7360 165
rect 7292 91 7360 131
rect 7292 57 7309 91
rect 7343 57 7360 91
rect 7292 34 7360 57
rect 7435 334 7469 350
rect 7435 262 7469 300
rect 7435 194 7469 228
rect 7531 218 7565 399
rect 7736 387 7804 427
rect 7736 353 7753 387
rect 7787 353 7804 387
rect 7531 168 7565 184
rect 7629 334 7663 350
rect 7629 262 7663 300
rect 7629 194 7663 228
rect 7435 124 7469 160
rect 7629 124 7663 160
rect 7469 90 7531 124
rect 7565 90 7629 124
rect 7435 34 7469 90
rect 7532 34 7566 90
rect 7629 34 7663 90
rect 7736 313 7804 353
rect 7736 279 7753 313
rect 7787 279 7804 313
rect 7736 239 7804 279
rect 7736 205 7753 239
rect 7787 205 7804 239
rect 7736 165 7804 205
rect 7736 131 7753 165
rect 7787 131 7804 165
rect 7736 91 7804 131
rect 7736 57 7753 91
rect 7787 57 7804 91
rect 7736 34 7804 57
rect -34 17 7804 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6569 17
rect 6603 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7804 17
rect -34 -34 7804 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5163 1463 5197 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5755 1463 5789 1497
rect 5829 1463 5863 1497
rect 5903 1463 5937 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6125 1463 6159 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6495 1463 6529 1497
rect 6569 1463 6603 1497
rect 6717 1463 6751 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7087 1463 7121 1497
rect 7161 1463 7195 1497
rect 7235 1463 7269 1497
rect 7383 1463 7417 1497
rect 7457 1463 7491 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7679 1463 7713 1497
rect 131 797 165 831
rect 649 797 683 831
rect 279 501 313 535
rect 871 797 905 831
rect 1315 871 1349 905
rect 945 723 979 757
rect 871 575 905 609
rect 649 434 683 461
rect 649 427 683 434
rect 1315 649 1349 683
rect 1537 501 1571 535
rect 2055 957 2089 979
rect 2055 945 2089 957
rect 1611 723 1645 757
rect 1907 797 1941 831
rect 1907 649 1941 683
rect 2055 871 2089 905
rect 2055 575 2089 609
rect 2351 797 2385 831
rect 2351 723 2385 757
rect 2351 434 2385 461
rect 2351 427 2385 434
rect 2869 797 2903 831
rect 2499 501 2533 535
rect 3091 797 3125 831
rect 3535 871 3569 905
rect 3165 723 3199 757
rect 3091 575 3125 609
rect 3535 649 3569 683
rect 3757 501 3791 535
rect 3831 723 3865 757
rect 4127 797 4161 831
rect 4127 649 4161 683
rect 4275 871 4309 905
rect 4645 871 4679 905
rect 4275 575 4309 609
rect 4793 433 4827 461
rect 4793 427 4827 433
rect 4941 649 4975 683
rect 5237 649 5271 683
rect 5755 923 5789 943
rect 5755 909 5789 923
rect 5385 575 5419 609
rect 6051 649 6085 683
rect 5903 433 5937 461
rect 5903 427 5937 433
rect 6347 649 6381 683
rect 6495 649 6529 683
rect 6865 575 6899 609
rect 7013 649 7047 683
rect 7161 649 7195 683
rect 7457 649 7491 683
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5163 -17 5197 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5755 -17 5789 17
rect 5829 -17 5863 17
rect 5903 -17 5937 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6125 -17 6159 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6495 -17 6529 17
rect 6569 -17 6603 17
rect 6717 -17 6751 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7087 -17 7121 17
rect 7161 -17 7195 17
rect 7235 -17 7269 17
rect 7383 -17 7417 17
rect 7457 -17 7491 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7679 -17 7713 17
<< metal1 >>
rect -34 1497 7804 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6569 1497
rect 6603 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7804 1497
rect -34 1446 7804 1463
rect 2049 979 2095 985
rect 2043 945 2055 979
rect 2089 949 5789 979
rect 2089 945 5795 949
rect 2049 939 2095 945
rect 5749 943 5795 945
rect 1309 905 1355 911
rect 2049 905 2095 911
rect 3529 905 3575 911
rect 4269 905 4315 911
rect 4639 905 4685 911
rect 5749 909 5755 943
rect 5789 909 5795 943
rect 1303 871 1315 905
rect 1349 871 2055 905
rect 2089 871 2101 905
rect 3523 871 3535 905
rect 3569 871 4275 905
rect 4309 871 4645 905
rect 4679 871 4691 905
rect 5749 903 5795 909
rect 5755 897 5789 903
rect 1309 865 1355 871
rect 2049 865 2095 871
rect 3529 865 3575 871
rect 4269 865 4315 871
rect 4639 865 4685 871
rect 125 831 171 837
rect 643 831 689 837
rect 865 831 911 837
rect 1901 831 1947 837
rect 2345 831 2391 837
rect 2863 831 2909 837
rect 3085 831 3131 837
rect 4121 831 4167 837
rect 119 797 131 831
rect 165 797 649 831
rect 683 797 695 831
rect 859 797 871 831
rect 905 797 1907 831
rect 1941 797 1953 831
rect 2339 797 2351 831
rect 2385 797 2869 831
rect 2903 797 2915 831
rect 3079 797 3091 831
rect 3125 797 4127 831
rect 4161 797 4173 831
rect 125 791 171 797
rect 643 791 689 797
rect 865 791 911 797
rect 1901 791 1947 797
rect 2345 791 2391 797
rect 2863 791 2909 797
rect 3085 791 3131 797
rect 4121 791 4167 797
rect 939 757 985 763
rect 1605 757 1651 763
rect 2345 757 2391 763
rect 3159 757 3205 763
rect 3825 757 3871 763
rect 933 723 945 757
rect 979 723 1611 757
rect 1645 723 2351 757
rect 2385 723 2397 757
rect 3153 723 3165 757
rect 3199 723 3831 757
rect 3865 723 3877 757
rect 939 717 985 723
rect 1605 717 1651 723
rect 2345 717 2391 723
rect 3159 717 3205 723
rect 3825 717 3871 723
rect 1309 683 1355 689
rect 1901 683 1947 689
rect 3529 683 3575 689
rect 4121 683 4167 689
rect 4935 683 4981 689
rect 5231 683 5277 689
rect 6045 683 6091 689
rect 6341 683 6387 689
rect 6489 683 6535 689
rect 7007 683 7053 689
rect 7155 683 7201 689
rect 7451 683 7497 689
rect 1303 649 1315 683
rect 1349 649 1907 683
rect 1941 649 1953 683
rect 3523 649 3535 683
rect 3569 649 4127 683
rect 4161 649 4173 683
rect 4929 649 4941 683
rect 4975 649 5237 683
rect 5271 649 5283 683
rect 6039 649 6051 683
rect 6085 649 6347 683
rect 6381 649 6393 683
rect 6483 649 6495 683
rect 6529 649 7013 683
rect 7047 649 7059 683
rect 7149 649 7161 683
rect 7195 649 7457 683
rect 7491 649 7503 683
rect 1309 643 1355 649
rect 1901 643 1947 649
rect 3529 643 3575 649
rect 4121 643 4167 649
rect 4935 643 4981 649
rect 5231 643 5277 649
rect 6045 643 6091 649
rect 6341 643 6387 649
rect 6489 643 6535 649
rect 7007 643 7053 649
rect 7155 643 7201 649
rect 7451 643 7497 649
rect 865 609 911 615
rect 2049 609 2095 615
rect 3085 609 3131 615
rect 4269 609 4315 615
rect 5379 609 5425 615
rect 6859 609 6905 615
rect 859 575 871 609
rect 905 575 2055 609
rect 2089 575 2101 609
rect 3079 575 3091 609
rect 3125 575 4275 609
rect 4309 575 4321 609
rect 5373 575 5385 609
rect 5419 575 6865 609
rect 6899 575 6911 609
rect 865 569 911 575
rect 2049 569 2095 575
rect 3085 569 3131 575
rect 4269 569 4315 575
rect 5379 569 5425 575
rect 6859 569 6905 575
rect 273 535 319 541
rect 1531 535 1577 541
rect 2493 535 2539 541
rect 3751 535 3797 541
rect 267 501 279 535
rect 313 501 1537 535
rect 1571 501 1583 535
rect 2487 501 2499 535
rect 2533 501 3757 535
rect 3791 501 3803 535
rect 273 495 319 501
rect 1531 495 1577 501
rect 2493 495 2539 501
rect 3751 495 3797 501
rect 649 467 683 473
rect 5903 467 5937 473
rect 643 461 689 467
rect 2345 461 2391 467
rect 4787 461 4833 467
rect 5897 461 5943 467
rect 643 427 649 461
rect 683 427 689 461
rect 2339 427 2351 461
rect 2385 427 4793 461
rect 4827 427 4839 461
rect 5897 427 5903 461
rect 5937 427 5943 461
rect 643 421 689 427
rect 2345 421 2391 427
rect 4787 421 4833 427
rect 5897 421 5943 427
rect 649 387 683 421
rect 5903 387 5937 421
rect 649 353 5937 387
rect -34 17 7804 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6569 17
rect 6603 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7804 17
rect -34 -34 7804 -17
<< labels >>
rlabel metal1 3831 723 3865 757 1 SUM
port 1 n
rlabel metal1 3831 501 3865 535 1 SUM
port 2 n
rlabel metal1 3165 723 3199 757 1 SUM
port 3 n
rlabel metal1 3165 649 3199 683 1 SUM
port 4 n
rlabel metal1 3165 871 3199 905 1 SUM
port 5 n
rlabel metal1 7605 649 7639 683 1 COUT
port 6 n
rlabel metal1 7605 723 7639 757 1 COUT
port 7 n
rlabel metal1 7605 797 7639 831 1 COUT
port 8 n
rlabel metal1 7605 871 7639 905 1 COUT
port 9 n
rlabel metal1 7605 575 7639 609 1 COUT
port 10 n
rlabel metal1 7605 501 7639 535 1 COUT
port 11 n
rlabel metal1 7605 427 7639 461 1 COUT
port 12 n
rlabel metal1 131 871 165 905 1 A
port 13 n
rlabel metal1 131 723 165 757 1 A
port 14 n
rlabel metal1 131 649 165 683 1 A
port 15 n
rlabel metal1 131 575 165 609 1 A
port 16 n
rlabel metal1 131 501 165 535 1 A
port 17 n
rlabel metal1 649 871 683 905 1 A
port 18 n
rlabel metal1 649 797 683 831 1 A
port 19 n
rlabel metal1 649 723 683 757 1 A
port 20 n
rlabel metal1 649 649 683 683 1 A
port 21 n
rlabel metal1 649 575 683 609 1 A
port 22 n
rlabel metal1 649 427 683 461 1 A
port 23 n
rlabel metal1 5903 871 5937 905 1 A
port 24 n
rlabel metal1 5903 797 5937 831 1 A
port 25 n
rlabel metal1 5903 723 5937 757 1 A
port 26 n
rlabel metal1 5903 649 5937 683 1 A
port 27 n
rlabel metal1 5903 501 5937 535 1 A
port 28 n
rlabel metal1 5903 427 5937 461 1 A
port 29 n
rlabel metal1 131 797 165 831 1 A
port 30 n
rlabel metal1 1315 871 1349 905 1 B
port 31 n
rlabel metal1 2055 871 2089 905 1 B
port 32 n
rlabel metal1 2055 945 2089 979 1 B
port 33 n
rlabel metal1 2055 797 2089 831 1 B
port 34 n
rlabel metal1 2055 649 2089 683 1 B
port 35 n
rlabel metal1 2055 501 2089 535 1 B
port 36 n
rlabel metal1 2055 575 2089 609 1 B
port 37 n
rlabel metal1 871 575 905 609 1 B
port 38 n
rlabel metal1 871 427 905 461 1 B
port 39 n
rlabel metal1 5755 649 5789 683 1 B
port 40 n
rlabel metal1 5755 723 5789 757 1 B
port 41 n
rlabel metal1 5755 797 5789 831 1 B
port 42 n
rlabel metal1 5755 871 5789 905 1 B
port 43 n
rlabel metal1 5755 945 5789 979 1 B
port 44 n
rlabel metal1 5755 501 5789 535 1 B
port 45 n
rlabel metal1 4645 871 4679 905 1 CIN
port 46 n
rlabel metal1 4645 797 4679 831 1 CIN
port 47 n
rlabel metal1 4645 723 4679 757 1 CIN
port 48 n
rlabel metal1 4645 649 4679 683 1 CIN
port 49 n
rlabel metal1 4645 575 4679 609 1 CIN
port 50 n
rlabel metal1 4645 501 4679 535 1 CIN
port 51 n
rlabel metal1 4275 871 4309 905 1 CIN
port 52 n
rlabel metal1 4275 575 4309 609 1 CIN
port 53 n
rlabel metal1 4275 649 4309 683 1 CIN
port 54 n
rlabel metal1 4275 723 4309 757 1 CIN
port 55 n
rlabel metal1 4275 797 4309 831 1 CIN
port 56 n
rlabel metal1 4275 501 4309 535 1 CIN
port 57 n
rlabel metal1 3535 871 3569 905 1 CIN
port 58 n
rlabel metal1 3091 575 3125 609 1 CIN
port 59 n
rlabel metal1 -34 1446 7804 1514 1 VPWR
port 60 n
rlabel metal1 -34 -34 7804 34 1 VGND
port 61 n
rlabel nwell 57 1463 91 1497 1 VPB
port 62 n
rlabel pwell 57 -17 91 17 1 VNB
port 63 n
<< end >>
