magic
tech sky130A
magscale 1 2
timestamp 1669507589
<< nwell >>
rect -87 786 5267 1550
<< pwell >>
rect -34 -34 5214 544
<< nmos >>
rect 147 290 177 351
tri 177 290 193 306 sw
rect 447 290 477 351
rect 147 260 253 290
tri 253 260 283 290 sw
rect 147 159 177 260
tri 177 244 193 260 nw
tri 237 244 253 260 ne
tri 177 159 193 175 sw
tri 237 159 253 175 se
rect 253 159 283 260
tri 342 260 372 290 se
rect 372 260 477 290
rect 342 166 372 260
tri 372 244 388 260 nw
tri 431 244 447 260 ne
tri 372 166 388 182 sw
tri 431 166 447 182 se
rect 447 166 477 260
tri 147 129 177 159 ne
rect 177 129 253 159
tri 253 129 283 159 nw
tri 342 136 372 166 ne
rect 372 136 447 166
tri 447 136 477 166 nw
rect 649 298 679 351
tri 679 298 695 314 sw
rect 649 268 755 298
tri 755 268 785 298 sw
rect 649 167 679 268
tri 679 252 695 268 nw
tri 739 252 755 268 ne
tri 679 167 695 183 sw
tri 739 167 755 183 se
rect 755 167 785 268
tri 649 137 679 167 ne
rect 679 137 755 167
tri 755 137 785 167 nw
rect 1109 290 1139 351
tri 1139 290 1155 306 sw
rect 1409 290 1439 351
rect 1109 260 1215 290
tri 1215 260 1245 290 sw
rect 1109 159 1139 260
tri 1139 244 1155 260 nw
tri 1199 244 1215 260 ne
tri 1139 159 1155 175 sw
tri 1199 159 1215 175 se
rect 1215 159 1245 260
tri 1304 260 1334 290 se
rect 1334 260 1439 290
rect 1304 166 1334 260
tri 1334 244 1350 260 nw
tri 1393 244 1409 260 ne
tri 1334 166 1350 182 sw
tri 1393 166 1409 182 se
rect 1409 166 1439 260
tri 1109 129 1139 159 ne
rect 1139 129 1215 159
tri 1215 129 1245 159 nw
tri 1304 136 1334 166 ne
rect 1334 136 1409 166
tri 1409 136 1439 166 nw
rect 1611 298 1641 351
tri 1641 298 1657 314 sw
rect 1611 268 1717 298
tri 1717 268 1747 298 sw
rect 1611 167 1641 268
tri 1641 252 1657 268 nw
tri 1701 252 1717 268 ne
tri 1641 167 1657 183 sw
tri 1701 167 1717 183 se
rect 1717 167 1747 268
tri 1611 137 1641 167 ne
rect 1641 137 1717 167
tri 1717 137 1747 167 nw
rect 2092 288 2122 349
tri 2122 288 2138 304 sw
rect 2286 296 2316 349
tri 2316 296 2332 312 sw
rect 2092 258 2198 288
tri 2198 258 2228 288 sw
rect 2286 266 2392 296
tri 2392 266 2422 296 sw
rect 2092 157 2122 258
tri 2122 242 2138 258 nw
tri 2182 242 2198 258 ne
tri 2122 157 2138 173 sw
tri 2182 157 2198 173 se
rect 2198 157 2228 258
rect 2286 165 2316 266
tri 2316 250 2332 266 nw
tri 2376 250 2392 266 ne
tri 2316 165 2332 181 sw
tri 2376 165 2392 181 se
rect 2392 165 2422 266
tri 2092 127 2122 157 ne
rect 2122 127 2198 157
tri 2198 127 2228 157 nw
tri 2286 135 2316 165 ne
rect 2316 135 2392 165
tri 2392 135 2422 165 nw
rect 2737 290 2767 351
tri 2767 290 2783 306 sw
rect 3037 290 3067 351
rect 2737 260 2843 290
tri 2843 260 2873 290 sw
rect 2737 159 2767 260
tri 2767 244 2783 260 nw
tri 2827 244 2843 260 ne
tri 2767 159 2783 175 sw
tri 2827 159 2843 175 se
rect 2843 159 2873 260
tri 2932 260 2962 290 se
rect 2962 260 3067 290
rect 2932 166 2962 260
tri 2962 244 2978 260 nw
tri 3021 244 3037 260 ne
tri 2962 166 2978 182 sw
tri 3021 166 3037 182 se
rect 3037 166 3067 260
tri 2737 129 2767 159 ne
rect 2767 129 2843 159
tri 2843 129 2873 159 nw
tri 2932 136 2962 166 ne
rect 2962 136 3037 166
tri 3037 136 3067 166 nw
rect 3239 298 3269 351
tri 3269 298 3285 314 sw
rect 3239 268 3345 298
tri 3345 268 3375 298 sw
rect 3239 167 3269 268
tri 3269 252 3285 268 nw
tri 3329 252 3345 268 ne
tri 3269 167 3285 183 sw
tri 3329 167 3345 183 se
rect 3345 167 3375 268
tri 3239 137 3269 167 ne
rect 3269 137 3345 167
tri 3345 137 3375 167 nw
rect 3699 290 3729 351
tri 3729 290 3745 306 sw
rect 3999 290 4029 351
rect 3699 260 3805 290
tri 3805 260 3835 290 sw
rect 3699 159 3729 260
tri 3729 244 3745 260 nw
tri 3789 244 3805 260 ne
tri 3729 159 3745 175 sw
tri 3789 159 3805 175 se
rect 3805 159 3835 260
tri 3894 260 3924 290 se
rect 3924 260 4029 290
rect 3894 166 3924 260
tri 3924 244 3940 260 nw
tri 3983 244 3999 260 ne
tri 3924 166 3940 182 sw
tri 3983 166 3999 182 se
rect 3999 166 4029 260
tri 3699 129 3729 159 ne
rect 3729 129 3805 159
tri 3805 129 3835 159 nw
tri 3894 136 3924 166 ne
rect 3924 136 3999 166
tri 3999 136 4029 166 nw
rect 4201 298 4231 351
tri 4231 298 4247 314 sw
rect 4201 268 4307 298
tri 4307 268 4337 298 sw
rect 4201 167 4231 268
tri 4231 252 4247 268 nw
tri 4291 252 4307 268 ne
tri 4231 167 4247 183 sw
tri 4291 167 4307 183 se
rect 4307 167 4337 268
tri 4201 137 4231 167 ne
rect 4231 137 4307 167
tri 4307 137 4337 167 nw
rect 4682 288 4712 349
tri 4712 288 4728 304 sw
rect 4876 296 4906 349
tri 4906 296 4922 312 sw
rect 4682 258 4788 288
tri 4788 258 4818 288 sw
rect 4876 266 4982 296
tri 4982 266 5012 296 sw
rect 4682 157 4712 258
tri 4712 242 4728 258 nw
tri 4772 242 4788 258 ne
tri 4712 157 4728 173 sw
tri 4772 157 4788 173 se
rect 4788 157 4818 258
rect 4876 165 4906 266
tri 4906 250 4922 266 nw
tri 4966 250 4982 266 ne
tri 4906 165 4922 181 sw
tri 4966 165 4982 181 se
rect 4982 165 5012 266
tri 4682 127 4712 157 ne
rect 4712 127 4788 157
tri 4788 127 4818 157 nw
tri 4876 135 4906 165 ne
rect 4906 135 4982 165
tri 4982 135 5012 165 nw
<< pmos >>
rect 247 1004 277 1404
rect 335 1004 365 1404
rect 423 1004 453 1404
rect 511 1004 541 1404
rect 599 1004 629 1404
rect 687 1004 717 1404
rect 1209 1004 1239 1404
rect 1297 1004 1327 1404
rect 1385 1004 1415 1404
rect 1473 1004 1503 1404
rect 1561 1004 1591 1404
rect 1649 1004 1679 1404
rect 2111 1004 2141 1404
rect 2199 1004 2229 1404
rect 2287 1004 2317 1404
rect 2375 1004 2405 1404
rect 2837 1004 2867 1404
rect 2925 1004 2955 1404
rect 3013 1004 3043 1404
rect 3101 1004 3131 1404
rect 3189 1004 3219 1404
rect 3277 1004 3307 1404
rect 3799 1004 3829 1404
rect 3887 1004 3917 1404
rect 3975 1004 4005 1404
rect 4063 1004 4093 1404
rect 4151 1004 4181 1404
rect 4239 1004 4269 1404
rect 4701 1004 4731 1404
rect 4789 1004 4819 1404
rect 4877 1004 4907 1404
rect 4965 1004 4995 1404
<< ndiff >>
rect 91 335 147 351
rect 91 301 101 335
rect 135 301 147 335
rect 91 263 147 301
rect 177 335 447 351
rect 177 306 198 335
tri 177 290 193 306 ne
rect 193 301 198 306
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 447 335
rect 193 290 447 301
rect 477 335 533 351
rect 477 301 489 335
rect 523 301 533 335
rect 91 229 101 263
rect 135 229 147 263
tri 253 260 283 290 ne
rect 283 263 342 290
rect 91 195 147 229
rect 91 161 101 195
rect 135 161 147 195
rect 91 129 147 161
tri 177 244 193 260 se
rect 193 244 237 260
tri 237 244 253 260 sw
rect 177 210 253 244
rect 177 176 198 210
rect 232 176 253 210
rect 177 175 253 176
tri 177 159 193 175 ne
rect 193 159 237 175
tri 237 159 253 175 nw
rect 283 229 295 263
rect 329 229 342 263
tri 342 260 372 290 nw
rect 283 195 342 229
rect 283 161 295 195
rect 329 161 342 195
tri 372 244 388 260 se
rect 388 244 431 260
tri 431 244 447 260 sw
rect 372 216 447 244
rect 372 182 393 216
rect 427 182 447 216
tri 372 166 388 182 ne
rect 388 166 431 182
tri 431 166 447 182 nw
tri 147 129 177 159 sw
tri 253 129 283 159 se
rect 283 136 342 161
tri 342 136 372 166 sw
tri 447 136 477 166 se
rect 477 136 533 301
rect 283 129 533 136
rect 91 125 533 129
rect 91 91 101 125
rect 135 91 295 125
rect 329 91 392 125
rect 426 91 489 125
rect 523 91 533 125
rect 91 75 533 91
rect 593 335 649 351
rect 593 301 603 335
rect 637 301 649 335
rect 593 263 649 301
rect 679 314 841 351
tri 679 298 695 314 ne
rect 695 298 841 314
tri 755 268 785 298 ne
rect 593 229 603 263
rect 637 229 649 263
rect 593 195 649 229
rect 593 161 603 195
rect 637 161 649 195
tri 679 252 695 268 se
rect 695 252 739 268
tri 739 252 755 268 sw
rect 679 219 755 252
rect 679 185 700 219
rect 734 185 755 219
rect 679 183 755 185
tri 679 167 695 183 ne
rect 695 167 739 183
tri 739 167 755 183 nw
rect 785 263 841 298
rect 785 229 797 263
rect 831 229 841 263
rect 785 195 841 229
rect 593 137 649 161
tri 649 137 679 167 sw
tri 755 137 785 167 se
rect 785 161 797 195
rect 831 161 841 195
rect 785 137 841 161
rect 593 125 841 137
rect 593 91 603 125
rect 637 91 700 125
rect 734 91 797 125
rect 831 91 841 125
rect 593 75 841 91
rect 1053 335 1109 351
rect 1053 301 1063 335
rect 1097 301 1109 335
rect 1053 263 1109 301
rect 1139 335 1409 351
rect 1139 306 1160 335
tri 1139 290 1155 306 ne
rect 1155 301 1160 306
rect 1194 301 1257 335
rect 1291 301 1354 335
rect 1388 301 1409 335
rect 1155 290 1409 301
rect 1439 335 1495 351
rect 1439 301 1451 335
rect 1485 301 1495 335
rect 1053 229 1063 263
rect 1097 229 1109 263
tri 1215 260 1245 290 ne
rect 1245 263 1304 290
rect 1053 195 1109 229
rect 1053 161 1063 195
rect 1097 161 1109 195
rect 1053 129 1109 161
tri 1139 244 1155 260 se
rect 1155 244 1199 260
tri 1199 244 1215 260 sw
rect 1139 210 1215 244
rect 1139 176 1160 210
rect 1194 176 1215 210
rect 1139 175 1215 176
tri 1139 159 1155 175 ne
rect 1155 159 1199 175
tri 1199 159 1215 175 nw
rect 1245 229 1257 263
rect 1291 229 1304 263
tri 1304 260 1334 290 nw
rect 1245 195 1304 229
rect 1245 161 1257 195
rect 1291 161 1304 195
tri 1334 244 1350 260 se
rect 1350 244 1393 260
tri 1393 244 1409 260 sw
rect 1334 216 1409 244
rect 1334 182 1355 216
rect 1389 182 1409 216
tri 1334 166 1350 182 ne
rect 1350 166 1393 182
tri 1393 166 1409 182 nw
tri 1109 129 1139 159 sw
tri 1215 129 1245 159 se
rect 1245 136 1304 161
tri 1304 136 1334 166 sw
tri 1409 136 1439 166 se
rect 1439 136 1495 301
rect 1245 129 1495 136
rect 1053 125 1495 129
rect 1053 91 1063 125
rect 1097 91 1257 125
rect 1291 91 1354 125
rect 1388 91 1451 125
rect 1485 91 1495 125
rect 1053 75 1495 91
rect 1555 335 1611 351
rect 1555 301 1565 335
rect 1599 301 1611 335
rect 1555 263 1611 301
rect 1641 314 1803 351
tri 1641 298 1657 314 ne
rect 1657 298 1803 314
tri 1717 268 1747 298 ne
rect 1555 229 1565 263
rect 1599 229 1611 263
rect 1555 195 1611 229
rect 1555 161 1565 195
rect 1599 161 1611 195
tri 1641 252 1657 268 se
rect 1657 252 1701 268
tri 1701 252 1717 268 sw
rect 1641 219 1717 252
rect 1641 185 1662 219
rect 1696 185 1717 219
rect 1641 183 1717 185
tri 1641 167 1657 183 ne
rect 1657 167 1701 183
tri 1701 167 1717 183 nw
rect 1747 263 1803 298
rect 1747 229 1759 263
rect 1793 229 1803 263
rect 1747 195 1803 229
rect 1555 137 1611 161
tri 1611 137 1641 167 sw
tri 1717 137 1747 167 se
rect 1747 161 1759 195
rect 1793 161 1803 195
rect 1747 137 1803 161
rect 1555 125 1803 137
rect 1555 91 1565 125
rect 1599 91 1662 125
rect 1696 91 1759 125
rect 1793 91 1803 125
rect 1555 75 1803 91
rect 2036 333 2092 349
rect 2036 299 2046 333
rect 2080 299 2092 333
rect 2036 261 2092 299
rect 2122 333 2286 349
rect 2122 304 2143 333
tri 2122 288 2138 304 ne
rect 2138 299 2143 304
rect 2177 299 2240 333
rect 2274 299 2286 333
rect 2138 288 2286 299
rect 2316 312 2478 349
tri 2316 296 2332 312 ne
rect 2332 296 2478 312
rect 2036 227 2046 261
rect 2080 227 2092 261
tri 2198 258 2228 288 ne
rect 2228 261 2286 288
tri 2392 266 2422 296 ne
rect 2036 193 2092 227
rect 2036 159 2046 193
rect 2080 159 2092 193
rect 2036 127 2092 159
tri 2122 242 2138 258 se
rect 2138 242 2182 258
tri 2182 242 2198 258 sw
rect 2122 208 2198 242
rect 2122 174 2143 208
rect 2177 174 2198 208
rect 2122 173 2198 174
tri 2122 157 2138 173 ne
rect 2138 157 2182 173
tri 2182 157 2198 173 nw
rect 2228 227 2240 261
rect 2274 227 2286 261
rect 2228 193 2286 227
rect 2228 159 2240 193
rect 2274 159 2286 193
tri 2316 250 2332 266 se
rect 2332 250 2376 266
tri 2376 250 2392 266 sw
rect 2316 217 2392 250
rect 2316 183 2337 217
rect 2371 183 2392 217
rect 2316 181 2392 183
tri 2316 165 2332 181 ne
rect 2332 165 2376 181
tri 2376 165 2392 181 nw
rect 2422 261 2478 296
rect 2422 227 2434 261
rect 2468 227 2478 261
rect 2422 193 2478 227
tri 2092 127 2122 157 sw
tri 2198 127 2228 157 se
rect 2228 135 2286 159
tri 2286 135 2316 165 sw
tri 2392 135 2422 165 se
rect 2422 159 2434 193
rect 2468 159 2478 193
rect 2422 135 2478 159
rect 2228 127 2478 135
rect 2036 123 2478 127
rect 2036 89 2046 123
rect 2080 89 2240 123
rect 2274 89 2337 123
rect 2371 89 2434 123
rect 2468 89 2478 123
rect 2036 73 2478 89
rect 2681 335 2737 351
rect 2681 301 2691 335
rect 2725 301 2737 335
rect 2681 263 2737 301
rect 2767 335 3037 351
rect 2767 306 2788 335
tri 2767 290 2783 306 ne
rect 2783 301 2788 306
rect 2822 301 2885 335
rect 2919 301 2982 335
rect 3016 301 3037 335
rect 2783 290 3037 301
rect 3067 335 3123 351
rect 3067 301 3079 335
rect 3113 301 3123 335
rect 2681 229 2691 263
rect 2725 229 2737 263
tri 2843 260 2873 290 ne
rect 2873 263 2932 290
rect 2681 195 2737 229
rect 2681 161 2691 195
rect 2725 161 2737 195
rect 2681 129 2737 161
tri 2767 244 2783 260 se
rect 2783 244 2827 260
tri 2827 244 2843 260 sw
rect 2767 210 2843 244
rect 2767 176 2788 210
rect 2822 176 2843 210
rect 2767 175 2843 176
tri 2767 159 2783 175 ne
rect 2783 159 2827 175
tri 2827 159 2843 175 nw
rect 2873 229 2885 263
rect 2919 229 2932 263
tri 2932 260 2962 290 nw
rect 2873 195 2932 229
rect 2873 161 2885 195
rect 2919 161 2932 195
tri 2962 244 2978 260 se
rect 2978 244 3021 260
tri 3021 244 3037 260 sw
rect 2962 216 3037 244
rect 2962 182 2983 216
rect 3017 182 3037 216
tri 2962 166 2978 182 ne
rect 2978 166 3021 182
tri 3021 166 3037 182 nw
tri 2737 129 2767 159 sw
tri 2843 129 2873 159 se
rect 2873 136 2932 161
tri 2932 136 2962 166 sw
tri 3037 136 3067 166 se
rect 3067 136 3123 301
rect 2873 129 3123 136
rect 2681 125 3123 129
rect 2681 91 2691 125
rect 2725 91 2885 125
rect 2919 91 2982 125
rect 3016 91 3079 125
rect 3113 91 3123 125
rect 2681 75 3123 91
rect 3183 335 3239 351
rect 3183 301 3193 335
rect 3227 301 3239 335
rect 3183 263 3239 301
rect 3269 314 3431 351
tri 3269 298 3285 314 ne
rect 3285 298 3431 314
tri 3345 268 3375 298 ne
rect 3183 229 3193 263
rect 3227 229 3239 263
rect 3183 195 3239 229
rect 3183 161 3193 195
rect 3227 161 3239 195
tri 3269 252 3285 268 se
rect 3285 252 3329 268
tri 3329 252 3345 268 sw
rect 3269 219 3345 252
rect 3269 185 3290 219
rect 3324 185 3345 219
rect 3269 183 3345 185
tri 3269 167 3285 183 ne
rect 3285 167 3329 183
tri 3329 167 3345 183 nw
rect 3375 263 3431 298
rect 3375 229 3387 263
rect 3421 229 3431 263
rect 3375 195 3431 229
rect 3183 137 3239 161
tri 3239 137 3269 167 sw
tri 3345 137 3375 167 se
rect 3375 161 3387 195
rect 3421 161 3431 195
rect 3375 137 3431 161
rect 3183 125 3431 137
rect 3183 91 3193 125
rect 3227 91 3290 125
rect 3324 91 3387 125
rect 3421 91 3431 125
rect 3183 75 3431 91
rect 3643 335 3699 351
rect 3643 301 3653 335
rect 3687 301 3699 335
rect 3643 263 3699 301
rect 3729 335 3999 351
rect 3729 306 3750 335
tri 3729 290 3745 306 ne
rect 3745 301 3750 306
rect 3784 301 3847 335
rect 3881 301 3944 335
rect 3978 301 3999 335
rect 3745 290 3999 301
rect 4029 335 4085 351
rect 4029 301 4041 335
rect 4075 301 4085 335
rect 3643 229 3653 263
rect 3687 229 3699 263
tri 3805 260 3835 290 ne
rect 3835 263 3894 290
rect 3643 195 3699 229
rect 3643 161 3653 195
rect 3687 161 3699 195
rect 3643 129 3699 161
tri 3729 244 3745 260 se
rect 3745 244 3789 260
tri 3789 244 3805 260 sw
rect 3729 210 3805 244
rect 3729 176 3750 210
rect 3784 176 3805 210
rect 3729 175 3805 176
tri 3729 159 3745 175 ne
rect 3745 159 3789 175
tri 3789 159 3805 175 nw
rect 3835 229 3847 263
rect 3881 229 3894 263
tri 3894 260 3924 290 nw
rect 3835 195 3894 229
rect 3835 161 3847 195
rect 3881 161 3894 195
tri 3924 244 3940 260 se
rect 3940 244 3983 260
tri 3983 244 3999 260 sw
rect 3924 216 3999 244
rect 3924 182 3945 216
rect 3979 182 3999 216
tri 3924 166 3940 182 ne
rect 3940 166 3983 182
tri 3983 166 3999 182 nw
tri 3699 129 3729 159 sw
tri 3805 129 3835 159 se
rect 3835 136 3894 161
tri 3894 136 3924 166 sw
tri 3999 136 4029 166 se
rect 4029 136 4085 301
rect 3835 129 4085 136
rect 3643 125 4085 129
rect 3643 91 3653 125
rect 3687 91 3847 125
rect 3881 91 3944 125
rect 3978 91 4041 125
rect 4075 91 4085 125
rect 3643 75 4085 91
rect 4145 335 4201 351
rect 4145 301 4155 335
rect 4189 301 4201 335
rect 4145 263 4201 301
rect 4231 314 4393 351
tri 4231 298 4247 314 ne
rect 4247 298 4393 314
tri 4307 268 4337 298 ne
rect 4145 229 4155 263
rect 4189 229 4201 263
rect 4145 195 4201 229
rect 4145 161 4155 195
rect 4189 161 4201 195
tri 4231 252 4247 268 se
rect 4247 252 4291 268
tri 4291 252 4307 268 sw
rect 4231 219 4307 252
rect 4231 185 4252 219
rect 4286 185 4307 219
rect 4231 183 4307 185
tri 4231 167 4247 183 ne
rect 4247 167 4291 183
tri 4291 167 4307 183 nw
rect 4337 263 4393 298
rect 4337 229 4349 263
rect 4383 229 4393 263
rect 4337 195 4393 229
rect 4145 137 4201 161
tri 4201 137 4231 167 sw
tri 4307 137 4337 167 se
rect 4337 161 4349 195
rect 4383 161 4393 195
rect 4337 137 4393 161
rect 4145 125 4393 137
rect 4145 91 4155 125
rect 4189 91 4252 125
rect 4286 91 4349 125
rect 4383 91 4393 125
rect 4145 75 4393 91
rect 4626 333 4682 349
rect 4626 299 4636 333
rect 4670 299 4682 333
rect 4626 261 4682 299
rect 4712 333 4876 349
rect 4712 304 4733 333
tri 4712 288 4728 304 ne
rect 4728 299 4733 304
rect 4767 299 4830 333
rect 4864 299 4876 333
rect 4728 288 4876 299
rect 4906 312 5068 349
tri 4906 296 4922 312 ne
rect 4922 296 5068 312
rect 4626 227 4636 261
rect 4670 227 4682 261
tri 4788 258 4818 288 ne
rect 4818 261 4876 288
tri 4982 266 5012 296 ne
rect 4626 193 4682 227
rect 4626 159 4636 193
rect 4670 159 4682 193
rect 4626 127 4682 159
tri 4712 242 4728 258 se
rect 4728 242 4772 258
tri 4772 242 4788 258 sw
rect 4712 208 4788 242
rect 4712 174 4733 208
rect 4767 174 4788 208
rect 4712 173 4788 174
tri 4712 157 4728 173 ne
rect 4728 157 4772 173
tri 4772 157 4788 173 nw
rect 4818 227 4830 261
rect 4864 227 4876 261
rect 4818 193 4876 227
rect 4818 159 4830 193
rect 4864 159 4876 193
tri 4906 250 4922 266 se
rect 4922 250 4966 266
tri 4966 250 4982 266 sw
rect 4906 217 4982 250
rect 4906 183 4927 217
rect 4961 183 4982 217
rect 4906 181 4982 183
tri 4906 165 4922 181 ne
rect 4922 165 4966 181
tri 4966 165 4982 181 nw
rect 5012 261 5068 296
rect 5012 227 5024 261
rect 5058 227 5068 261
rect 5012 193 5068 227
tri 4682 127 4712 157 sw
tri 4788 127 4818 157 se
rect 4818 135 4876 159
tri 4876 135 4906 165 sw
tri 4982 135 5012 165 se
rect 5012 159 5024 193
rect 5058 159 5068 193
rect 5012 135 5068 159
rect 4818 127 5068 135
rect 4626 123 5068 127
rect 4626 89 4636 123
rect 4670 89 4830 123
rect 4864 89 4927 123
rect 4961 89 5024 123
rect 5058 89 5068 123
rect 4626 73 5068 89
<< pdiff >>
rect 191 1366 247 1404
rect 191 1332 201 1366
rect 235 1332 247 1366
rect 191 1298 247 1332
rect 191 1264 201 1298
rect 235 1264 247 1298
rect 191 1230 247 1264
rect 191 1196 201 1230
rect 235 1196 247 1230
rect 191 1162 247 1196
rect 191 1128 201 1162
rect 235 1128 247 1162
rect 191 1093 247 1128
rect 191 1059 201 1093
rect 235 1059 247 1093
rect 191 1004 247 1059
rect 277 1366 335 1404
rect 277 1332 289 1366
rect 323 1332 335 1366
rect 277 1298 335 1332
rect 277 1264 289 1298
rect 323 1264 335 1298
rect 277 1230 335 1264
rect 277 1196 289 1230
rect 323 1196 335 1230
rect 277 1162 335 1196
rect 277 1128 289 1162
rect 323 1128 335 1162
rect 277 1093 335 1128
rect 277 1059 289 1093
rect 323 1059 335 1093
rect 277 1004 335 1059
rect 365 1366 423 1404
rect 365 1332 377 1366
rect 411 1332 423 1366
rect 365 1298 423 1332
rect 365 1264 377 1298
rect 411 1264 423 1298
rect 365 1230 423 1264
rect 365 1196 377 1230
rect 411 1196 423 1230
rect 365 1162 423 1196
rect 365 1128 377 1162
rect 411 1128 423 1162
rect 365 1004 423 1128
rect 453 1366 511 1404
rect 453 1332 465 1366
rect 499 1332 511 1366
rect 453 1298 511 1332
rect 453 1264 465 1298
rect 499 1264 511 1298
rect 453 1230 511 1264
rect 453 1196 465 1230
rect 499 1196 511 1230
rect 453 1162 511 1196
rect 453 1128 465 1162
rect 499 1128 511 1162
rect 453 1093 511 1128
rect 453 1059 465 1093
rect 499 1059 511 1093
rect 453 1004 511 1059
rect 541 1366 599 1404
rect 541 1332 553 1366
rect 587 1332 599 1366
rect 541 1298 599 1332
rect 541 1264 553 1298
rect 587 1264 599 1298
rect 541 1230 599 1264
rect 541 1196 553 1230
rect 587 1196 599 1230
rect 541 1162 599 1196
rect 541 1128 553 1162
rect 587 1128 599 1162
rect 541 1004 599 1128
rect 629 1366 687 1404
rect 629 1332 641 1366
rect 675 1332 687 1366
rect 629 1298 687 1332
rect 629 1264 641 1298
rect 675 1264 687 1298
rect 629 1230 687 1264
rect 629 1196 641 1230
rect 675 1196 687 1230
rect 629 1162 687 1196
rect 629 1128 641 1162
rect 675 1128 687 1162
rect 629 1093 687 1128
rect 629 1059 641 1093
rect 675 1059 687 1093
rect 629 1004 687 1059
rect 717 1366 771 1404
rect 717 1332 729 1366
rect 763 1332 771 1366
rect 717 1298 771 1332
rect 717 1264 729 1298
rect 763 1264 771 1298
rect 717 1230 771 1264
rect 717 1196 729 1230
rect 763 1196 771 1230
rect 717 1162 771 1196
rect 717 1128 729 1162
rect 763 1128 771 1162
rect 717 1004 771 1128
rect 1153 1366 1209 1404
rect 1153 1332 1163 1366
rect 1197 1332 1209 1366
rect 1153 1298 1209 1332
rect 1153 1264 1163 1298
rect 1197 1264 1209 1298
rect 1153 1230 1209 1264
rect 1153 1196 1163 1230
rect 1197 1196 1209 1230
rect 1153 1162 1209 1196
rect 1153 1128 1163 1162
rect 1197 1128 1209 1162
rect 1153 1093 1209 1128
rect 1153 1059 1163 1093
rect 1197 1059 1209 1093
rect 1153 1004 1209 1059
rect 1239 1366 1297 1404
rect 1239 1332 1251 1366
rect 1285 1332 1297 1366
rect 1239 1298 1297 1332
rect 1239 1264 1251 1298
rect 1285 1264 1297 1298
rect 1239 1230 1297 1264
rect 1239 1196 1251 1230
rect 1285 1196 1297 1230
rect 1239 1162 1297 1196
rect 1239 1128 1251 1162
rect 1285 1128 1297 1162
rect 1239 1093 1297 1128
rect 1239 1059 1251 1093
rect 1285 1059 1297 1093
rect 1239 1004 1297 1059
rect 1327 1366 1385 1404
rect 1327 1332 1339 1366
rect 1373 1332 1385 1366
rect 1327 1298 1385 1332
rect 1327 1264 1339 1298
rect 1373 1264 1385 1298
rect 1327 1230 1385 1264
rect 1327 1196 1339 1230
rect 1373 1196 1385 1230
rect 1327 1162 1385 1196
rect 1327 1128 1339 1162
rect 1373 1128 1385 1162
rect 1327 1004 1385 1128
rect 1415 1366 1473 1404
rect 1415 1332 1427 1366
rect 1461 1332 1473 1366
rect 1415 1298 1473 1332
rect 1415 1264 1427 1298
rect 1461 1264 1473 1298
rect 1415 1230 1473 1264
rect 1415 1196 1427 1230
rect 1461 1196 1473 1230
rect 1415 1162 1473 1196
rect 1415 1128 1427 1162
rect 1461 1128 1473 1162
rect 1415 1093 1473 1128
rect 1415 1059 1427 1093
rect 1461 1059 1473 1093
rect 1415 1004 1473 1059
rect 1503 1366 1561 1404
rect 1503 1332 1515 1366
rect 1549 1332 1561 1366
rect 1503 1298 1561 1332
rect 1503 1264 1515 1298
rect 1549 1264 1561 1298
rect 1503 1230 1561 1264
rect 1503 1196 1515 1230
rect 1549 1196 1561 1230
rect 1503 1162 1561 1196
rect 1503 1128 1515 1162
rect 1549 1128 1561 1162
rect 1503 1004 1561 1128
rect 1591 1366 1649 1404
rect 1591 1332 1603 1366
rect 1637 1332 1649 1366
rect 1591 1298 1649 1332
rect 1591 1264 1603 1298
rect 1637 1264 1649 1298
rect 1591 1230 1649 1264
rect 1591 1196 1603 1230
rect 1637 1196 1649 1230
rect 1591 1162 1649 1196
rect 1591 1128 1603 1162
rect 1637 1128 1649 1162
rect 1591 1093 1649 1128
rect 1591 1059 1603 1093
rect 1637 1059 1649 1093
rect 1591 1004 1649 1059
rect 1679 1366 1733 1404
rect 1679 1332 1691 1366
rect 1725 1332 1733 1366
rect 1679 1298 1733 1332
rect 1679 1264 1691 1298
rect 1725 1264 1733 1298
rect 1679 1230 1733 1264
rect 1679 1196 1691 1230
rect 1725 1196 1733 1230
rect 1679 1162 1733 1196
rect 1679 1128 1691 1162
rect 1725 1128 1733 1162
rect 1679 1004 1733 1128
rect 2055 1366 2111 1404
rect 2055 1332 2065 1366
rect 2099 1332 2111 1366
rect 2055 1298 2111 1332
rect 2055 1264 2065 1298
rect 2099 1264 2111 1298
rect 2055 1230 2111 1264
rect 2055 1196 2065 1230
rect 2099 1196 2111 1230
rect 2055 1162 2111 1196
rect 2055 1128 2065 1162
rect 2099 1128 2111 1162
rect 2055 1093 2111 1128
rect 2055 1059 2065 1093
rect 2099 1059 2111 1093
rect 2055 1004 2111 1059
rect 2141 1366 2199 1404
rect 2141 1332 2153 1366
rect 2187 1332 2199 1366
rect 2141 1298 2199 1332
rect 2141 1264 2153 1298
rect 2187 1264 2199 1298
rect 2141 1230 2199 1264
rect 2141 1196 2153 1230
rect 2187 1196 2199 1230
rect 2141 1162 2199 1196
rect 2141 1128 2153 1162
rect 2187 1128 2199 1162
rect 2141 1093 2199 1128
rect 2141 1059 2153 1093
rect 2187 1059 2199 1093
rect 2141 1004 2199 1059
rect 2229 1366 2287 1404
rect 2229 1332 2241 1366
rect 2275 1332 2287 1366
rect 2229 1298 2287 1332
rect 2229 1264 2241 1298
rect 2275 1264 2287 1298
rect 2229 1230 2287 1264
rect 2229 1196 2241 1230
rect 2275 1196 2287 1230
rect 2229 1162 2287 1196
rect 2229 1128 2241 1162
rect 2275 1128 2287 1162
rect 2229 1004 2287 1128
rect 2317 1366 2375 1404
rect 2317 1332 2329 1366
rect 2363 1332 2375 1366
rect 2317 1298 2375 1332
rect 2317 1264 2329 1298
rect 2363 1264 2375 1298
rect 2317 1230 2375 1264
rect 2317 1196 2329 1230
rect 2363 1196 2375 1230
rect 2317 1162 2375 1196
rect 2317 1128 2329 1162
rect 2363 1128 2375 1162
rect 2317 1093 2375 1128
rect 2317 1059 2329 1093
rect 2363 1059 2375 1093
rect 2317 1004 2375 1059
rect 2405 1366 2459 1404
rect 2405 1332 2417 1366
rect 2451 1332 2459 1366
rect 2405 1298 2459 1332
rect 2405 1264 2417 1298
rect 2451 1264 2459 1298
rect 2405 1230 2459 1264
rect 2405 1196 2417 1230
rect 2451 1196 2459 1230
rect 2405 1162 2459 1196
rect 2405 1128 2417 1162
rect 2451 1128 2459 1162
rect 2405 1004 2459 1128
rect 2781 1366 2837 1404
rect 2781 1332 2791 1366
rect 2825 1332 2837 1366
rect 2781 1298 2837 1332
rect 2781 1264 2791 1298
rect 2825 1264 2837 1298
rect 2781 1230 2837 1264
rect 2781 1196 2791 1230
rect 2825 1196 2837 1230
rect 2781 1162 2837 1196
rect 2781 1128 2791 1162
rect 2825 1128 2837 1162
rect 2781 1093 2837 1128
rect 2781 1059 2791 1093
rect 2825 1059 2837 1093
rect 2781 1004 2837 1059
rect 2867 1366 2925 1404
rect 2867 1332 2879 1366
rect 2913 1332 2925 1366
rect 2867 1298 2925 1332
rect 2867 1264 2879 1298
rect 2913 1264 2925 1298
rect 2867 1230 2925 1264
rect 2867 1196 2879 1230
rect 2913 1196 2925 1230
rect 2867 1162 2925 1196
rect 2867 1128 2879 1162
rect 2913 1128 2925 1162
rect 2867 1093 2925 1128
rect 2867 1059 2879 1093
rect 2913 1059 2925 1093
rect 2867 1004 2925 1059
rect 2955 1366 3013 1404
rect 2955 1332 2967 1366
rect 3001 1332 3013 1366
rect 2955 1298 3013 1332
rect 2955 1264 2967 1298
rect 3001 1264 3013 1298
rect 2955 1230 3013 1264
rect 2955 1196 2967 1230
rect 3001 1196 3013 1230
rect 2955 1162 3013 1196
rect 2955 1128 2967 1162
rect 3001 1128 3013 1162
rect 2955 1004 3013 1128
rect 3043 1366 3101 1404
rect 3043 1332 3055 1366
rect 3089 1332 3101 1366
rect 3043 1298 3101 1332
rect 3043 1264 3055 1298
rect 3089 1264 3101 1298
rect 3043 1230 3101 1264
rect 3043 1196 3055 1230
rect 3089 1196 3101 1230
rect 3043 1162 3101 1196
rect 3043 1128 3055 1162
rect 3089 1128 3101 1162
rect 3043 1093 3101 1128
rect 3043 1059 3055 1093
rect 3089 1059 3101 1093
rect 3043 1004 3101 1059
rect 3131 1366 3189 1404
rect 3131 1332 3143 1366
rect 3177 1332 3189 1366
rect 3131 1298 3189 1332
rect 3131 1264 3143 1298
rect 3177 1264 3189 1298
rect 3131 1230 3189 1264
rect 3131 1196 3143 1230
rect 3177 1196 3189 1230
rect 3131 1162 3189 1196
rect 3131 1128 3143 1162
rect 3177 1128 3189 1162
rect 3131 1004 3189 1128
rect 3219 1366 3277 1404
rect 3219 1332 3231 1366
rect 3265 1332 3277 1366
rect 3219 1298 3277 1332
rect 3219 1264 3231 1298
rect 3265 1264 3277 1298
rect 3219 1230 3277 1264
rect 3219 1196 3231 1230
rect 3265 1196 3277 1230
rect 3219 1162 3277 1196
rect 3219 1128 3231 1162
rect 3265 1128 3277 1162
rect 3219 1093 3277 1128
rect 3219 1059 3231 1093
rect 3265 1059 3277 1093
rect 3219 1004 3277 1059
rect 3307 1366 3361 1404
rect 3307 1332 3319 1366
rect 3353 1332 3361 1366
rect 3307 1298 3361 1332
rect 3307 1264 3319 1298
rect 3353 1264 3361 1298
rect 3307 1230 3361 1264
rect 3307 1196 3319 1230
rect 3353 1196 3361 1230
rect 3307 1162 3361 1196
rect 3307 1128 3319 1162
rect 3353 1128 3361 1162
rect 3307 1004 3361 1128
rect 3743 1366 3799 1404
rect 3743 1332 3753 1366
rect 3787 1332 3799 1366
rect 3743 1298 3799 1332
rect 3743 1264 3753 1298
rect 3787 1264 3799 1298
rect 3743 1230 3799 1264
rect 3743 1196 3753 1230
rect 3787 1196 3799 1230
rect 3743 1162 3799 1196
rect 3743 1128 3753 1162
rect 3787 1128 3799 1162
rect 3743 1093 3799 1128
rect 3743 1059 3753 1093
rect 3787 1059 3799 1093
rect 3743 1004 3799 1059
rect 3829 1366 3887 1404
rect 3829 1332 3841 1366
rect 3875 1332 3887 1366
rect 3829 1298 3887 1332
rect 3829 1264 3841 1298
rect 3875 1264 3887 1298
rect 3829 1230 3887 1264
rect 3829 1196 3841 1230
rect 3875 1196 3887 1230
rect 3829 1162 3887 1196
rect 3829 1128 3841 1162
rect 3875 1128 3887 1162
rect 3829 1093 3887 1128
rect 3829 1059 3841 1093
rect 3875 1059 3887 1093
rect 3829 1004 3887 1059
rect 3917 1366 3975 1404
rect 3917 1332 3929 1366
rect 3963 1332 3975 1366
rect 3917 1298 3975 1332
rect 3917 1264 3929 1298
rect 3963 1264 3975 1298
rect 3917 1230 3975 1264
rect 3917 1196 3929 1230
rect 3963 1196 3975 1230
rect 3917 1162 3975 1196
rect 3917 1128 3929 1162
rect 3963 1128 3975 1162
rect 3917 1004 3975 1128
rect 4005 1366 4063 1404
rect 4005 1332 4017 1366
rect 4051 1332 4063 1366
rect 4005 1298 4063 1332
rect 4005 1264 4017 1298
rect 4051 1264 4063 1298
rect 4005 1230 4063 1264
rect 4005 1196 4017 1230
rect 4051 1196 4063 1230
rect 4005 1162 4063 1196
rect 4005 1128 4017 1162
rect 4051 1128 4063 1162
rect 4005 1093 4063 1128
rect 4005 1059 4017 1093
rect 4051 1059 4063 1093
rect 4005 1004 4063 1059
rect 4093 1366 4151 1404
rect 4093 1332 4105 1366
rect 4139 1332 4151 1366
rect 4093 1298 4151 1332
rect 4093 1264 4105 1298
rect 4139 1264 4151 1298
rect 4093 1230 4151 1264
rect 4093 1196 4105 1230
rect 4139 1196 4151 1230
rect 4093 1162 4151 1196
rect 4093 1128 4105 1162
rect 4139 1128 4151 1162
rect 4093 1004 4151 1128
rect 4181 1366 4239 1404
rect 4181 1332 4193 1366
rect 4227 1332 4239 1366
rect 4181 1298 4239 1332
rect 4181 1264 4193 1298
rect 4227 1264 4239 1298
rect 4181 1230 4239 1264
rect 4181 1196 4193 1230
rect 4227 1196 4239 1230
rect 4181 1162 4239 1196
rect 4181 1128 4193 1162
rect 4227 1128 4239 1162
rect 4181 1093 4239 1128
rect 4181 1059 4193 1093
rect 4227 1059 4239 1093
rect 4181 1004 4239 1059
rect 4269 1366 4323 1404
rect 4269 1332 4281 1366
rect 4315 1332 4323 1366
rect 4269 1298 4323 1332
rect 4269 1264 4281 1298
rect 4315 1264 4323 1298
rect 4269 1230 4323 1264
rect 4269 1196 4281 1230
rect 4315 1196 4323 1230
rect 4269 1162 4323 1196
rect 4269 1128 4281 1162
rect 4315 1128 4323 1162
rect 4269 1004 4323 1128
rect 4645 1366 4701 1404
rect 4645 1332 4655 1366
rect 4689 1332 4701 1366
rect 4645 1298 4701 1332
rect 4645 1264 4655 1298
rect 4689 1264 4701 1298
rect 4645 1230 4701 1264
rect 4645 1196 4655 1230
rect 4689 1196 4701 1230
rect 4645 1162 4701 1196
rect 4645 1128 4655 1162
rect 4689 1128 4701 1162
rect 4645 1093 4701 1128
rect 4645 1059 4655 1093
rect 4689 1059 4701 1093
rect 4645 1004 4701 1059
rect 4731 1366 4789 1404
rect 4731 1332 4743 1366
rect 4777 1332 4789 1366
rect 4731 1298 4789 1332
rect 4731 1264 4743 1298
rect 4777 1264 4789 1298
rect 4731 1230 4789 1264
rect 4731 1196 4743 1230
rect 4777 1196 4789 1230
rect 4731 1162 4789 1196
rect 4731 1128 4743 1162
rect 4777 1128 4789 1162
rect 4731 1093 4789 1128
rect 4731 1059 4743 1093
rect 4777 1059 4789 1093
rect 4731 1004 4789 1059
rect 4819 1366 4877 1404
rect 4819 1332 4831 1366
rect 4865 1332 4877 1366
rect 4819 1298 4877 1332
rect 4819 1264 4831 1298
rect 4865 1264 4877 1298
rect 4819 1230 4877 1264
rect 4819 1196 4831 1230
rect 4865 1196 4877 1230
rect 4819 1162 4877 1196
rect 4819 1128 4831 1162
rect 4865 1128 4877 1162
rect 4819 1004 4877 1128
rect 4907 1366 4965 1404
rect 4907 1332 4919 1366
rect 4953 1332 4965 1366
rect 4907 1298 4965 1332
rect 4907 1264 4919 1298
rect 4953 1264 4965 1298
rect 4907 1230 4965 1264
rect 4907 1196 4919 1230
rect 4953 1196 4965 1230
rect 4907 1162 4965 1196
rect 4907 1128 4919 1162
rect 4953 1128 4965 1162
rect 4907 1093 4965 1128
rect 4907 1059 4919 1093
rect 4953 1059 4965 1093
rect 4907 1004 4965 1059
rect 4995 1366 5049 1404
rect 4995 1332 5007 1366
rect 5041 1332 5049 1366
rect 4995 1298 5049 1332
rect 4995 1264 5007 1298
rect 5041 1264 5049 1298
rect 4995 1230 5049 1264
rect 4995 1196 5007 1230
rect 5041 1196 5049 1230
rect 4995 1162 5049 1196
rect 4995 1128 5007 1162
rect 5041 1128 5049 1162
rect 4995 1004 5049 1128
<< ndiffc >>
rect 101 301 135 335
rect 198 301 232 335
rect 295 301 329 335
rect 392 301 426 335
rect 489 301 523 335
rect 101 229 135 263
rect 101 161 135 195
rect 198 176 232 210
rect 295 229 329 263
rect 295 161 329 195
rect 393 182 427 216
rect 101 91 135 125
rect 295 91 329 125
rect 392 91 426 125
rect 489 91 523 125
rect 603 301 637 335
rect 603 229 637 263
rect 603 161 637 195
rect 700 185 734 219
rect 797 229 831 263
rect 797 161 831 195
rect 603 91 637 125
rect 700 91 734 125
rect 797 91 831 125
rect 1063 301 1097 335
rect 1160 301 1194 335
rect 1257 301 1291 335
rect 1354 301 1388 335
rect 1451 301 1485 335
rect 1063 229 1097 263
rect 1063 161 1097 195
rect 1160 176 1194 210
rect 1257 229 1291 263
rect 1257 161 1291 195
rect 1355 182 1389 216
rect 1063 91 1097 125
rect 1257 91 1291 125
rect 1354 91 1388 125
rect 1451 91 1485 125
rect 1565 301 1599 335
rect 1565 229 1599 263
rect 1565 161 1599 195
rect 1662 185 1696 219
rect 1759 229 1793 263
rect 1759 161 1793 195
rect 1565 91 1599 125
rect 1662 91 1696 125
rect 1759 91 1793 125
rect 2046 299 2080 333
rect 2143 299 2177 333
rect 2240 299 2274 333
rect 2046 227 2080 261
rect 2046 159 2080 193
rect 2143 174 2177 208
rect 2240 227 2274 261
rect 2240 159 2274 193
rect 2337 183 2371 217
rect 2434 227 2468 261
rect 2434 159 2468 193
rect 2046 89 2080 123
rect 2240 89 2274 123
rect 2337 89 2371 123
rect 2434 89 2468 123
rect 2691 301 2725 335
rect 2788 301 2822 335
rect 2885 301 2919 335
rect 2982 301 3016 335
rect 3079 301 3113 335
rect 2691 229 2725 263
rect 2691 161 2725 195
rect 2788 176 2822 210
rect 2885 229 2919 263
rect 2885 161 2919 195
rect 2983 182 3017 216
rect 2691 91 2725 125
rect 2885 91 2919 125
rect 2982 91 3016 125
rect 3079 91 3113 125
rect 3193 301 3227 335
rect 3193 229 3227 263
rect 3193 161 3227 195
rect 3290 185 3324 219
rect 3387 229 3421 263
rect 3387 161 3421 195
rect 3193 91 3227 125
rect 3290 91 3324 125
rect 3387 91 3421 125
rect 3653 301 3687 335
rect 3750 301 3784 335
rect 3847 301 3881 335
rect 3944 301 3978 335
rect 4041 301 4075 335
rect 3653 229 3687 263
rect 3653 161 3687 195
rect 3750 176 3784 210
rect 3847 229 3881 263
rect 3847 161 3881 195
rect 3945 182 3979 216
rect 3653 91 3687 125
rect 3847 91 3881 125
rect 3944 91 3978 125
rect 4041 91 4075 125
rect 4155 301 4189 335
rect 4155 229 4189 263
rect 4155 161 4189 195
rect 4252 185 4286 219
rect 4349 229 4383 263
rect 4349 161 4383 195
rect 4155 91 4189 125
rect 4252 91 4286 125
rect 4349 91 4383 125
rect 4636 299 4670 333
rect 4733 299 4767 333
rect 4830 299 4864 333
rect 4636 227 4670 261
rect 4636 159 4670 193
rect 4733 174 4767 208
rect 4830 227 4864 261
rect 4830 159 4864 193
rect 4927 183 4961 217
rect 5024 227 5058 261
rect 5024 159 5058 193
rect 4636 89 4670 123
rect 4830 89 4864 123
rect 4927 89 4961 123
rect 5024 89 5058 123
<< pdiffc >>
rect 201 1332 235 1366
rect 201 1264 235 1298
rect 201 1196 235 1230
rect 201 1128 235 1162
rect 201 1059 235 1093
rect 289 1332 323 1366
rect 289 1264 323 1298
rect 289 1196 323 1230
rect 289 1128 323 1162
rect 289 1059 323 1093
rect 377 1332 411 1366
rect 377 1264 411 1298
rect 377 1196 411 1230
rect 377 1128 411 1162
rect 465 1332 499 1366
rect 465 1264 499 1298
rect 465 1196 499 1230
rect 465 1128 499 1162
rect 465 1059 499 1093
rect 553 1332 587 1366
rect 553 1264 587 1298
rect 553 1196 587 1230
rect 553 1128 587 1162
rect 641 1332 675 1366
rect 641 1264 675 1298
rect 641 1196 675 1230
rect 641 1128 675 1162
rect 641 1059 675 1093
rect 729 1332 763 1366
rect 729 1264 763 1298
rect 729 1196 763 1230
rect 729 1128 763 1162
rect 1163 1332 1197 1366
rect 1163 1264 1197 1298
rect 1163 1196 1197 1230
rect 1163 1128 1197 1162
rect 1163 1059 1197 1093
rect 1251 1332 1285 1366
rect 1251 1264 1285 1298
rect 1251 1196 1285 1230
rect 1251 1128 1285 1162
rect 1251 1059 1285 1093
rect 1339 1332 1373 1366
rect 1339 1264 1373 1298
rect 1339 1196 1373 1230
rect 1339 1128 1373 1162
rect 1427 1332 1461 1366
rect 1427 1264 1461 1298
rect 1427 1196 1461 1230
rect 1427 1128 1461 1162
rect 1427 1059 1461 1093
rect 1515 1332 1549 1366
rect 1515 1264 1549 1298
rect 1515 1196 1549 1230
rect 1515 1128 1549 1162
rect 1603 1332 1637 1366
rect 1603 1264 1637 1298
rect 1603 1196 1637 1230
rect 1603 1128 1637 1162
rect 1603 1059 1637 1093
rect 1691 1332 1725 1366
rect 1691 1264 1725 1298
rect 1691 1196 1725 1230
rect 1691 1128 1725 1162
rect 2065 1332 2099 1366
rect 2065 1264 2099 1298
rect 2065 1196 2099 1230
rect 2065 1128 2099 1162
rect 2065 1059 2099 1093
rect 2153 1332 2187 1366
rect 2153 1264 2187 1298
rect 2153 1196 2187 1230
rect 2153 1128 2187 1162
rect 2153 1059 2187 1093
rect 2241 1332 2275 1366
rect 2241 1264 2275 1298
rect 2241 1196 2275 1230
rect 2241 1128 2275 1162
rect 2329 1332 2363 1366
rect 2329 1264 2363 1298
rect 2329 1196 2363 1230
rect 2329 1128 2363 1162
rect 2329 1059 2363 1093
rect 2417 1332 2451 1366
rect 2417 1264 2451 1298
rect 2417 1196 2451 1230
rect 2417 1128 2451 1162
rect 2791 1332 2825 1366
rect 2791 1264 2825 1298
rect 2791 1196 2825 1230
rect 2791 1128 2825 1162
rect 2791 1059 2825 1093
rect 2879 1332 2913 1366
rect 2879 1264 2913 1298
rect 2879 1196 2913 1230
rect 2879 1128 2913 1162
rect 2879 1059 2913 1093
rect 2967 1332 3001 1366
rect 2967 1264 3001 1298
rect 2967 1196 3001 1230
rect 2967 1128 3001 1162
rect 3055 1332 3089 1366
rect 3055 1264 3089 1298
rect 3055 1196 3089 1230
rect 3055 1128 3089 1162
rect 3055 1059 3089 1093
rect 3143 1332 3177 1366
rect 3143 1264 3177 1298
rect 3143 1196 3177 1230
rect 3143 1128 3177 1162
rect 3231 1332 3265 1366
rect 3231 1264 3265 1298
rect 3231 1196 3265 1230
rect 3231 1128 3265 1162
rect 3231 1059 3265 1093
rect 3319 1332 3353 1366
rect 3319 1264 3353 1298
rect 3319 1196 3353 1230
rect 3319 1128 3353 1162
rect 3753 1332 3787 1366
rect 3753 1264 3787 1298
rect 3753 1196 3787 1230
rect 3753 1128 3787 1162
rect 3753 1059 3787 1093
rect 3841 1332 3875 1366
rect 3841 1264 3875 1298
rect 3841 1196 3875 1230
rect 3841 1128 3875 1162
rect 3841 1059 3875 1093
rect 3929 1332 3963 1366
rect 3929 1264 3963 1298
rect 3929 1196 3963 1230
rect 3929 1128 3963 1162
rect 4017 1332 4051 1366
rect 4017 1264 4051 1298
rect 4017 1196 4051 1230
rect 4017 1128 4051 1162
rect 4017 1059 4051 1093
rect 4105 1332 4139 1366
rect 4105 1264 4139 1298
rect 4105 1196 4139 1230
rect 4105 1128 4139 1162
rect 4193 1332 4227 1366
rect 4193 1264 4227 1298
rect 4193 1196 4227 1230
rect 4193 1128 4227 1162
rect 4193 1059 4227 1093
rect 4281 1332 4315 1366
rect 4281 1264 4315 1298
rect 4281 1196 4315 1230
rect 4281 1128 4315 1162
rect 4655 1332 4689 1366
rect 4655 1264 4689 1298
rect 4655 1196 4689 1230
rect 4655 1128 4689 1162
rect 4655 1059 4689 1093
rect 4743 1332 4777 1366
rect 4743 1264 4777 1298
rect 4743 1196 4777 1230
rect 4743 1128 4777 1162
rect 4743 1059 4777 1093
rect 4831 1332 4865 1366
rect 4831 1264 4865 1298
rect 4831 1196 4865 1230
rect 4831 1128 4865 1162
rect 4919 1332 4953 1366
rect 4919 1264 4953 1298
rect 4919 1196 4953 1230
rect 4919 1128 4953 1162
rect 4919 1059 4953 1093
rect 5007 1332 5041 1366
rect 5007 1264 5041 1298
rect 5007 1196 5041 1230
rect 5007 1128 5041 1162
<< psubdiff >>
rect -34 482 5214 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 928 461 996 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 928 427 945 461
rect 979 427 996 461
rect 1890 461 1958 482
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 928 313 996 353
rect 1890 427 1907 461
rect 1941 427 1958 461
rect 2556 461 2624 482
rect 1890 387 1958 427
rect 1890 353 1907 387
rect 1941 353 1958 387
rect 928 279 945 313
rect 979 279 996 313
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect -34 17 34 57
rect 928 57 945 91
rect 979 57 996 91
rect 1890 313 1958 353
rect 2556 427 2573 461
rect 2607 427 2624 461
rect 3518 461 3586 482
rect 2556 387 2624 427
rect 2556 353 2573 387
rect 2607 353 2624 387
rect 1890 279 1907 313
rect 1941 279 1958 313
rect 1890 239 1958 279
rect 1890 205 1907 239
rect 1941 205 1958 239
rect 1890 165 1958 205
rect 1890 131 1907 165
rect 1941 131 1958 165
rect 1890 91 1958 131
rect 928 17 996 57
rect 1890 57 1907 91
rect 1941 57 1958 91
rect 2556 313 2624 353
rect 3518 427 3535 461
rect 3569 427 3586 461
rect 4480 461 4548 482
rect 3518 387 3586 427
rect 3518 353 3535 387
rect 3569 353 3586 387
rect 2556 279 2573 313
rect 2607 279 2624 313
rect 2556 239 2624 279
rect 2556 205 2573 239
rect 2607 205 2624 239
rect 2556 165 2624 205
rect 2556 131 2573 165
rect 2607 131 2624 165
rect 2556 91 2624 131
rect 1890 17 1958 57
rect 2556 57 2573 91
rect 2607 57 2624 91
rect 3518 313 3586 353
rect 4480 427 4497 461
rect 4531 427 4548 461
rect 5146 461 5214 482
rect 4480 387 4548 427
rect 4480 353 4497 387
rect 4531 353 4548 387
rect 3518 279 3535 313
rect 3569 279 3586 313
rect 3518 239 3586 279
rect 3518 205 3535 239
rect 3569 205 3586 239
rect 3518 165 3586 205
rect 3518 131 3535 165
rect 3569 131 3586 165
rect 3518 91 3586 131
rect 2556 17 2624 57
rect 3518 57 3535 91
rect 3569 57 3586 91
rect 4480 313 4548 353
rect 5146 427 5163 461
rect 5197 427 5214 461
rect 5146 387 5214 427
rect 5146 353 5163 387
rect 5197 353 5214 387
rect 4480 279 4497 313
rect 4531 279 4548 313
rect 4480 239 4548 279
rect 4480 205 4497 239
rect 4531 205 4548 239
rect 4480 165 4548 205
rect 4480 131 4497 165
rect 4531 131 4548 165
rect 4480 91 4548 131
rect 3518 17 3586 57
rect 4480 57 4497 91
rect 4531 57 4548 91
rect 5146 313 5214 353
rect 5146 279 5163 313
rect 5197 279 5214 313
rect 5146 239 5214 279
rect 5146 205 5163 239
rect 5197 205 5214 239
rect 5146 165 5214 205
rect 5146 131 5163 165
rect 5197 131 5214 165
rect 5146 91 5214 131
rect 4480 17 4548 57
rect 5146 57 5163 91
rect 5197 57 5214 91
rect 5146 17 5214 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5214 17
rect -34 -34 5214 -17
<< nsubdiff >>
rect -34 1497 5214 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5214 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 928 1423 996 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 1890 1423 1958 1463
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect 928 1019 945 1053
rect 979 1019 996 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 928 979 996 1019
rect 1890 1389 1907 1423
rect 1941 1389 1958 1423
rect 2556 1423 2624 1463
rect 1890 1349 1958 1389
rect 1890 1315 1907 1349
rect 1941 1315 1958 1349
rect 1890 1275 1958 1315
rect 1890 1241 1907 1275
rect 1941 1241 1958 1275
rect 1890 1201 1958 1241
rect 1890 1167 1907 1201
rect 1941 1167 1958 1201
rect 1890 1127 1958 1167
rect 1890 1093 1907 1127
rect 1941 1093 1958 1127
rect 1890 1053 1958 1093
rect 1890 1019 1907 1053
rect 1941 1019 1958 1053
rect 928 945 945 979
rect 979 945 996 979
rect -34 871 -17 905
rect 17 884 34 905
rect 928 905 996 945
rect 1890 979 1958 1019
rect 2556 1389 2573 1423
rect 2607 1389 2624 1423
rect 3518 1423 3586 1463
rect 2556 1349 2624 1389
rect 2556 1315 2573 1349
rect 2607 1315 2624 1349
rect 2556 1275 2624 1315
rect 2556 1241 2573 1275
rect 2607 1241 2624 1275
rect 2556 1201 2624 1241
rect 2556 1167 2573 1201
rect 2607 1167 2624 1201
rect 2556 1127 2624 1167
rect 2556 1093 2573 1127
rect 2607 1093 2624 1127
rect 2556 1053 2624 1093
rect 2556 1019 2573 1053
rect 2607 1019 2624 1053
rect 1890 945 1907 979
rect 1941 945 1958 979
rect 928 884 945 905
rect 17 871 945 884
rect 979 884 996 905
rect 1890 905 1958 945
rect 2556 979 2624 1019
rect 3518 1389 3535 1423
rect 3569 1389 3586 1423
rect 4480 1423 4548 1463
rect 3518 1349 3586 1389
rect 3518 1315 3535 1349
rect 3569 1315 3586 1349
rect 3518 1275 3586 1315
rect 3518 1241 3535 1275
rect 3569 1241 3586 1275
rect 3518 1201 3586 1241
rect 3518 1167 3535 1201
rect 3569 1167 3586 1201
rect 3518 1127 3586 1167
rect 3518 1093 3535 1127
rect 3569 1093 3586 1127
rect 3518 1053 3586 1093
rect 3518 1019 3535 1053
rect 3569 1019 3586 1053
rect 2556 945 2573 979
rect 2607 945 2624 979
rect 1890 884 1907 905
rect 979 871 1907 884
rect 1941 884 1958 905
rect 2556 905 2624 945
rect 3518 979 3586 1019
rect 4480 1389 4497 1423
rect 4531 1389 4548 1423
rect 5146 1423 5214 1463
rect 4480 1349 4548 1389
rect 4480 1315 4497 1349
rect 4531 1315 4548 1349
rect 4480 1275 4548 1315
rect 4480 1241 4497 1275
rect 4531 1241 4548 1275
rect 4480 1201 4548 1241
rect 4480 1167 4497 1201
rect 4531 1167 4548 1201
rect 4480 1127 4548 1167
rect 4480 1093 4497 1127
rect 4531 1093 4548 1127
rect 4480 1053 4548 1093
rect 4480 1019 4497 1053
rect 4531 1019 4548 1053
rect 3518 945 3535 979
rect 3569 945 3586 979
rect 2556 884 2573 905
rect 1941 871 2573 884
rect 2607 884 2624 905
rect 3518 905 3586 945
rect 4480 979 4548 1019
rect 5146 1389 5163 1423
rect 5197 1389 5214 1423
rect 5146 1349 5214 1389
rect 5146 1315 5163 1349
rect 5197 1315 5214 1349
rect 5146 1275 5214 1315
rect 5146 1241 5163 1275
rect 5197 1241 5214 1275
rect 5146 1201 5214 1241
rect 5146 1167 5163 1201
rect 5197 1167 5214 1201
rect 5146 1127 5214 1167
rect 5146 1093 5163 1127
rect 5197 1093 5214 1127
rect 5146 1053 5214 1093
rect 5146 1019 5163 1053
rect 5197 1019 5214 1053
rect 4480 945 4497 979
rect 4531 945 4548 979
rect 3518 884 3535 905
rect 2607 871 3535 884
rect 3569 884 3586 905
rect 4480 905 4548 945
rect 5146 979 5214 1019
rect 5146 945 5163 979
rect 5197 945 5214 979
rect 4480 884 4497 905
rect 3569 871 4497 884
rect 4531 884 4548 905
rect 5146 905 5214 945
rect 5146 884 5163 905
rect 4531 871 5163 884
rect 5197 871 5214 905
rect -34 822 5214 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 945 427 979 461
rect 945 353 979 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1907 427 1941 461
rect 1907 353 1941 387
rect 945 279 979 313
rect 945 205 979 239
rect 945 131 979 165
rect 945 57 979 91
rect 2573 427 2607 461
rect 2573 353 2607 387
rect 1907 279 1941 313
rect 1907 205 1941 239
rect 1907 131 1941 165
rect 1907 57 1941 91
rect 3535 427 3569 461
rect 3535 353 3569 387
rect 2573 279 2607 313
rect 2573 205 2607 239
rect 2573 131 2607 165
rect 2573 57 2607 91
rect 4497 427 4531 461
rect 4497 353 4531 387
rect 3535 279 3569 313
rect 3535 205 3569 239
rect 3535 131 3569 165
rect 3535 57 3569 91
rect 5163 427 5197 461
rect 5163 353 5197 387
rect 4497 279 4531 313
rect 4497 205 4531 239
rect 4497 131 4531 165
rect 4497 57 4531 91
rect 5163 279 5197 313
rect 5163 205 5197 239
rect 5163 131 5197 165
rect 5163 57 5197 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 945 1389 979 1423
rect 945 1315 979 1349
rect 945 1241 979 1275
rect 945 1167 979 1201
rect 945 1093 979 1127
rect 945 1019 979 1053
rect -17 945 17 979
rect 1907 1389 1941 1423
rect 1907 1315 1941 1349
rect 1907 1241 1941 1275
rect 1907 1167 1941 1201
rect 1907 1093 1941 1127
rect 1907 1019 1941 1053
rect 945 945 979 979
rect -17 871 17 905
rect 2573 1389 2607 1423
rect 2573 1315 2607 1349
rect 2573 1241 2607 1275
rect 2573 1167 2607 1201
rect 2573 1093 2607 1127
rect 2573 1019 2607 1053
rect 1907 945 1941 979
rect 945 871 979 905
rect 3535 1389 3569 1423
rect 3535 1315 3569 1349
rect 3535 1241 3569 1275
rect 3535 1167 3569 1201
rect 3535 1093 3569 1127
rect 3535 1019 3569 1053
rect 2573 945 2607 979
rect 1907 871 1941 905
rect 4497 1389 4531 1423
rect 4497 1315 4531 1349
rect 4497 1241 4531 1275
rect 4497 1167 4531 1201
rect 4497 1093 4531 1127
rect 4497 1019 4531 1053
rect 3535 945 3569 979
rect 2573 871 2607 905
rect 5163 1389 5197 1423
rect 5163 1315 5197 1349
rect 5163 1241 5197 1275
rect 5163 1167 5197 1201
rect 5163 1093 5197 1127
rect 5163 1019 5197 1053
rect 4497 945 4531 979
rect 3535 871 3569 905
rect 5163 945 5197 979
rect 4497 871 4531 905
rect 5163 871 5197 905
<< poly >>
rect 247 1404 277 1430
rect 335 1404 365 1430
rect 423 1404 453 1430
rect 511 1404 541 1430
rect 599 1404 629 1430
rect 687 1404 717 1430
rect 1209 1404 1239 1430
rect 1297 1404 1327 1430
rect 1385 1404 1415 1430
rect 1473 1404 1503 1430
rect 1561 1404 1591 1430
rect 1649 1404 1679 1430
rect 247 973 277 1004
rect 335 973 365 1004
rect 423 973 453 1004
rect 511 973 541 1004
rect 195 957 365 973
rect 195 923 205 957
rect 239 943 365 957
rect 417 957 541 973
rect 239 923 249 943
rect 195 907 249 923
rect 417 923 427 957
rect 461 943 541 957
rect 599 973 629 1004
rect 687 973 717 1004
rect 599 957 717 973
rect 599 943 649 957
rect 461 923 471 943
rect 417 907 471 923
rect 639 923 649 943
rect 683 943 717 957
rect 2111 1404 2141 1430
rect 2199 1404 2229 1430
rect 2287 1404 2317 1430
rect 2375 1404 2405 1430
rect 1209 973 1239 1004
rect 1297 973 1327 1004
rect 1385 973 1415 1004
rect 1473 973 1503 1004
rect 683 923 693 943
rect 639 907 693 923
rect 1157 957 1327 973
rect 1157 923 1167 957
rect 1201 943 1327 957
rect 1379 957 1503 973
rect 1201 923 1211 943
rect 1157 907 1211 923
rect 1379 923 1389 957
rect 1423 943 1503 957
rect 1561 973 1591 1004
rect 1649 973 1679 1004
rect 1561 957 1679 973
rect 1561 943 1611 957
rect 1423 923 1433 943
rect 1379 907 1433 923
rect 1601 923 1611 943
rect 1645 943 1679 957
rect 2837 1404 2867 1430
rect 2925 1404 2955 1430
rect 3013 1404 3043 1430
rect 3101 1404 3131 1430
rect 3189 1404 3219 1430
rect 3277 1404 3307 1430
rect 1645 923 1655 943
rect 1601 907 1655 923
rect 2111 973 2141 1004
rect 2199 973 2229 1004
rect 2287 973 2317 1004
rect 2375 973 2405 1004
rect 2111 957 2229 973
rect 2111 943 2129 957
rect 2119 923 2129 943
rect 2163 943 2229 957
rect 2273 957 2405 973
rect 2163 923 2173 943
rect 2119 907 2173 923
rect 2273 923 2283 957
rect 2317 943 2405 957
rect 3799 1404 3829 1430
rect 3887 1404 3917 1430
rect 3975 1404 4005 1430
rect 4063 1404 4093 1430
rect 4151 1404 4181 1430
rect 4239 1404 4269 1430
rect 2837 973 2867 1004
rect 2925 973 2955 1004
rect 3013 973 3043 1004
rect 3101 973 3131 1004
rect 2317 923 2327 943
rect 2273 907 2327 923
rect 2785 957 2955 973
rect 2785 923 2795 957
rect 2829 943 2955 957
rect 3007 957 3131 973
rect 2829 923 2839 943
rect 2785 907 2839 923
rect 3007 923 3017 957
rect 3051 943 3131 957
rect 3189 973 3219 1004
rect 3277 973 3307 1004
rect 3189 957 3307 973
rect 3189 943 3239 957
rect 3051 923 3061 943
rect 3007 907 3061 923
rect 3229 923 3239 943
rect 3273 943 3307 957
rect 4701 1404 4731 1430
rect 4789 1404 4819 1430
rect 4877 1404 4907 1430
rect 4965 1404 4995 1430
rect 3799 973 3829 1004
rect 3887 973 3917 1004
rect 3975 973 4005 1004
rect 4063 973 4093 1004
rect 3273 923 3283 943
rect 3229 907 3283 923
rect 3747 957 3917 973
rect 3747 923 3757 957
rect 3791 943 3917 957
rect 3969 957 4093 973
rect 3791 923 3801 943
rect 3747 907 3801 923
rect 3969 923 3979 957
rect 4013 943 4093 957
rect 4151 973 4181 1004
rect 4239 973 4269 1004
rect 4151 957 4269 973
rect 4151 943 4201 957
rect 4013 923 4023 943
rect 3969 907 4023 923
rect 4191 923 4201 943
rect 4235 943 4269 957
rect 4235 923 4245 943
rect 4191 907 4245 923
rect 4701 973 4731 1004
rect 4789 973 4819 1004
rect 4877 973 4907 1004
rect 4965 973 4995 1004
rect 4701 957 4819 973
rect 4701 943 4719 957
rect 4709 923 4719 943
rect 4753 943 4819 957
rect 4863 957 4995 973
rect 4753 923 4763 943
rect 4709 907 4763 923
rect 4863 923 4873 957
rect 4907 943 4995 957
rect 4907 923 4917 943
rect 4863 907 4917 923
rect 195 433 249 449
rect 195 413 205 433
rect 147 399 205 413
rect 239 399 249 433
rect 147 383 249 399
rect 417 433 471 449
rect 417 399 427 433
rect 461 413 471 433
rect 639 433 693 449
rect 461 399 477 413
rect 417 383 477 399
rect 639 399 649 433
rect 683 399 693 433
rect 639 383 693 399
rect 1157 433 1211 449
rect 1157 413 1167 433
rect 147 351 177 383
rect 447 351 477 383
rect 649 351 679 383
rect 1109 399 1167 413
rect 1201 399 1211 433
rect 1109 383 1211 399
rect 1379 433 1433 449
rect 1379 399 1389 433
rect 1423 413 1433 433
rect 1601 433 1655 449
rect 1423 399 1439 413
rect 1379 383 1439 399
rect 1601 399 1611 433
rect 1645 399 1655 433
rect 1601 383 1655 399
rect 2119 433 2173 449
rect 2119 413 2129 433
rect 1109 351 1139 383
rect 1409 351 1439 383
rect 1611 351 1641 383
rect 2092 399 2129 413
rect 2163 399 2173 433
rect 2092 383 2173 399
rect 2267 433 2321 449
rect 2267 399 2277 433
rect 2311 399 2321 433
rect 2267 383 2321 399
rect 2785 433 2839 449
rect 2785 413 2795 433
rect 2092 349 2122 383
rect 2286 349 2316 383
rect 2737 399 2795 413
rect 2829 399 2839 433
rect 2737 383 2839 399
rect 3007 433 3061 449
rect 3007 399 3017 433
rect 3051 413 3061 433
rect 3229 433 3283 449
rect 3051 399 3067 413
rect 3007 383 3067 399
rect 3229 399 3239 433
rect 3273 399 3283 433
rect 3229 383 3283 399
rect 3747 433 3801 449
rect 3747 413 3757 433
rect 2737 351 2767 383
rect 3037 351 3067 383
rect 3239 351 3269 383
rect 3699 399 3757 413
rect 3791 399 3801 433
rect 3699 383 3801 399
rect 3969 433 4023 449
rect 3969 399 3979 433
rect 4013 413 4023 433
rect 4191 433 4245 449
rect 4013 399 4029 413
rect 3969 383 4029 399
rect 4191 399 4201 433
rect 4235 399 4245 433
rect 4191 383 4245 399
rect 4709 433 4763 449
rect 4709 413 4719 433
rect 3699 351 3729 383
rect 3999 351 4029 383
rect 4201 351 4231 383
rect 4682 399 4719 413
rect 4753 399 4763 433
rect 4682 383 4763 399
rect 4857 433 4911 449
rect 4857 399 4867 433
rect 4901 399 4911 433
rect 4857 383 4911 399
rect 4682 349 4712 383
rect 4876 349 4906 383
<< polycont >>
rect 205 923 239 957
rect 427 923 461 957
rect 649 923 683 957
rect 1167 923 1201 957
rect 1389 923 1423 957
rect 1611 923 1645 957
rect 2129 923 2163 957
rect 2283 923 2317 957
rect 2795 923 2829 957
rect 3017 923 3051 957
rect 3239 923 3273 957
rect 3757 923 3791 957
rect 3979 923 4013 957
rect 4201 923 4235 957
rect 4719 923 4753 957
rect 4873 923 4907 957
rect 205 399 239 433
rect 427 399 461 433
rect 649 399 683 433
rect 1167 399 1201 433
rect 1389 399 1423 433
rect 1611 399 1645 433
rect 2129 399 2163 433
rect 2277 399 2311 433
rect 2795 399 2829 433
rect 3017 399 3051 433
rect 3239 399 3273 433
rect 3757 399 3791 433
rect 3979 399 4013 433
rect 4201 399 4235 433
rect 4719 399 4753 433
rect 4867 399 4901 433
<< locali >>
rect -34 1497 5214 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5214 1497
rect -34 1446 5214 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 201 1366 235 1446
rect 201 1298 235 1332
rect 201 1230 235 1264
rect 201 1162 235 1196
rect 201 1093 235 1128
rect 201 1043 235 1059
rect 289 1366 323 1404
rect 289 1298 323 1332
rect 289 1230 323 1264
rect 289 1162 323 1196
rect 289 1093 323 1128
rect 377 1366 411 1446
rect 377 1298 411 1332
rect 377 1230 411 1264
rect 377 1162 411 1196
rect 377 1111 411 1128
rect 465 1366 499 1404
rect 465 1298 499 1332
rect 465 1230 499 1264
rect 465 1162 499 1196
rect 289 1048 323 1059
rect 465 1093 499 1128
rect 553 1366 587 1446
rect 553 1298 587 1332
rect 553 1230 587 1264
rect 553 1162 587 1196
rect 553 1111 587 1128
rect 641 1366 675 1404
rect 641 1298 675 1332
rect 641 1230 675 1264
rect 641 1162 675 1196
rect 465 1048 499 1059
rect 641 1093 675 1128
rect 729 1366 763 1446
rect 729 1298 763 1332
rect 729 1230 763 1264
rect 729 1162 763 1196
rect 729 1111 763 1128
rect 928 1423 996 1446
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 641 1048 675 1059
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect -34 979 34 1019
rect 289 1014 831 1048
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 205 831 239 923
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 797
rect 205 383 239 399
rect 427 957 461 973
rect 427 905 461 923
rect 427 433 461 871
rect 427 383 461 399
rect 649 957 683 973
rect 649 683 683 923
rect 649 433 683 649
rect 649 383 683 399
rect 797 757 831 1014
rect 928 1019 945 1053
rect 979 1019 996 1053
rect 1163 1366 1197 1446
rect 1163 1298 1197 1332
rect 1163 1230 1197 1264
rect 1163 1162 1197 1196
rect 1163 1093 1197 1128
rect 1163 1043 1197 1059
rect 1251 1366 1285 1404
rect 1251 1298 1285 1332
rect 1251 1230 1285 1264
rect 1251 1162 1285 1196
rect 1251 1093 1285 1128
rect 1339 1366 1373 1446
rect 1339 1298 1373 1332
rect 1339 1230 1373 1264
rect 1339 1162 1373 1196
rect 1339 1111 1373 1128
rect 1427 1366 1461 1404
rect 1427 1298 1461 1332
rect 1427 1230 1461 1264
rect 1427 1162 1461 1196
rect 1251 1048 1285 1059
rect 1427 1093 1461 1128
rect 1515 1366 1549 1446
rect 1515 1298 1549 1332
rect 1515 1230 1549 1264
rect 1515 1162 1549 1196
rect 1515 1111 1549 1128
rect 1603 1366 1637 1404
rect 1603 1298 1637 1332
rect 1603 1230 1637 1264
rect 1603 1162 1637 1196
rect 1427 1048 1461 1059
rect 1603 1093 1637 1128
rect 1691 1366 1725 1446
rect 1691 1298 1725 1332
rect 1691 1230 1725 1264
rect 1691 1162 1725 1196
rect 1691 1111 1725 1128
rect 1890 1423 1958 1446
rect 1890 1389 1907 1423
rect 1941 1389 1958 1423
rect 1890 1349 1958 1389
rect 1890 1315 1907 1349
rect 1941 1315 1958 1349
rect 1890 1275 1958 1315
rect 1890 1241 1907 1275
rect 1941 1241 1958 1275
rect 1890 1201 1958 1241
rect 1890 1167 1907 1201
rect 1941 1167 1958 1201
rect 1890 1127 1958 1167
rect 1603 1048 1637 1059
rect 1890 1093 1907 1127
rect 1941 1093 1958 1127
rect 1890 1053 1958 1093
rect 928 979 996 1019
rect 1251 1014 1793 1048
rect 928 945 945 979
rect 979 945 996 979
rect 928 905 996 945
rect 928 871 945 905
rect 979 871 996 905
rect 928 822 996 871
rect 1167 957 1201 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 101 335 135 351
rect 295 335 329 351
rect 489 335 523 351
rect 135 301 198 335
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 489 335
rect 101 263 135 301
rect 101 195 135 229
rect 295 263 329 301
rect 489 285 523 301
rect 603 335 637 351
rect 797 350 831 723
rect 1167 757 1201 923
rect 603 263 637 301
rect 101 125 135 161
rect 101 75 135 91
rect 198 210 232 226
rect -34 34 34 57
rect 198 34 232 176
rect 295 195 329 229
rect 393 216 427 232
rect 603 216 637 229
rect 427 195 637 216
rect 427 182 603 195
rect 393 166 427 182
rect 295 125 329 161
rect 700 316 831 350
rect 928 461 996 544
rect 928 427 945 461
rect 979 427 996 461
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect 1167 433 1201 723
rect 1167 383 1201 399
rect 1389 957 1423 973
rect 1389 433 1423 923
rect 1389 383 1423 399
rect 1611 957 1645 973
rect 1611 461 1645 923
rect 1611 383 1645 399
rect 1759 683 1793 1014
rect 1890 1019 1907 1053
rect 1941 1019 1958 1053
rect 2065 1366 2099 1446
rect 2065 1298 2099 1332
rect 2065 1230 2099 1264
rect 2065 1162 2099 1196
rect 2065 1093 2099 1128
rect 2065 1027 2099 1059
rect 2153 1366 2187 1404
rect 2153 1298 2187 1332
rect 2153 1230 2187 1264
rect 2153 1162 2187 1196
rect 2153 1093 2187 1128
rect 2241 1366 2275 1446
rect 2241 1298 2275 1332
rect 2241 1230 2275 1264
rect 2241 1162 2275 1196
rect 2241 1111 2275 1128
rect 2329 1366 2363 1404
rect 2329 1298 2363 1332
rect 2329 1230 2363 1264
rect 2329 1162 2363 1196
rect 2153 1057 2187 1059
rect 2329 1093 2363 1128
rect 2417 1366 2451 1446
rect 2417 1298 2451 1332
rect 2417 1230 2451 1264
rect 2417 1162 2451 1196
rect 2417 1111 2451 1128
rect 2556 1423 2624 1446
rect 2556 1389 2573 1423
rect 2607 1389 2624 1423
rect 2556 1349 2624 1389
rect 2556 1315 2573 1349
rect 2607 1315 2624 1349
rect 2556 1275 2624 1315
rect 2556 1241 2573 1275
rect 2607 1241 2624 1275
rect 2556 1201 2624 1241
rect 2556 1167 2573 1201
rect 2607 1167 2624 1201
rect 2556 1127 2624 1167
rect 2329 1057 2363 1059
rect 2556 1093 2573 1127
rect 2607 1093 2624 1127
rect 2153 1023 2459 1057
rect 1890 979 1958 1019
rect 1890 945 1907 979
rect 1941 945 1958 979
rect 1890 905 1958 945
rect 1890 871 1907 905
rect 1941 871 1958 905
rect 1890 822 1958 871
rect 2129 957 2163 973
rect 2283 957 2317 973
rect 700 219 734 316
rect 928 313 996 353
rect 928 279 945 313
rect 979 279 996 313
rect 700 169 734 185
rect 797 263 831 279
rect 797 195 831 229
rect 489 125 523 141
rect 329 91 392 125
rect 426 91 489 125
rect 295 75 329 91
rect 489 75 523 91
rect 603 125 637 161
rect 797 125 831 161
rect 637 91 700 125
rect 734 91 797 125
rect 603 75 637 91
rect 797 75 831 91
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect 928 57 945 91
rect 979 57 996 91
rect 1063 335 1097 351
rect 1257 335 1291 351
rect 1451 335 1485 351
rect 1097 301 1160 335
rect 1194 301 1257 335
rect 1291 301 1354 335
rect 1388 301 1451 335
rect 1063 263 1097 301
rect 1063 195 1097 229
rect 1257 263 1291 301
rect 1451 285 1485 301
rect 1565 335 1599 351
rect 1759 350 1793 649
rect 2129 683 2163 923
rect 1565 263 1599 301
rect 1063 125 1097 161
rect 1063 75 1097 91
rect 1160 210 1194 226
rect 928 34 996 57
rect 1160 34 1194 176
rect 1257 195 1291 229
rect 1355 216 1389 232
rect 1565 216 1599 229
rect 1389 195 1599 216
rect 1389 182 1565 195
rect 1355 166 1389 182
rect 1257 125 1291 161
rect 1662 316 1793 350
rect 1890 461 1958 544
rect 1890 427 1907 461
rect 1941 427 1958 461
rect 1890 387 1958 427
rect 1890 353 1907 387
rect 1941 353 1958 387
rect 2129 433 2163 649
rect 2129 383 2163 399
rect 2277 923 2283 942
rect 2277 907 2317 923
rect 2277 831 2311 907
rect 2277 433 2311 797
rect 2277 383 2311 399
rect 2425 683 2459 1023
rect 2556 1053 2624 1093
rect 2556 1019 2573 1053
rect 2607 1019 2624 1053
rect 2791 1366 2825 1446
rect 2791 1298 2825 1332
rect 2791 1230 2825 1264
rect 2791 1162 2825 1196
rect 2791 1093 2825 1128
rect 2791 1043 2825 1059
rect 2879 1366 2913 1404
rect 2879 1298 2913 1332
rect 2879 1230 2913 1264
rect 2879 1162 2913 1196
rect 2879 1093 2913 1128
rect 2967 1366 3001 1446
rect 2967 1298 3001 1332
rect 2967 1230 3001 1264
rect 2967 1162 3001 1196
rect 2967 1111 3001 1128
rect 3055 1366 3089 1404
rect 3055 1298 3089 1332
rect 3055 1230 3089 1264
rect 3055 1162 3089 1196
rect 2879 1048 2913 1059
rect 3055 1093 3089 1128
rect 3143 1366 3177 1446
rect 3143 1298 3177 1332
rect 3143 1230 3177 1264
rect 3143 1162 3177 1196
rect 3143 1111 3177 1128
rect 3231 1366 3265 1404
rect 3231 1298 3265 1332
rect 3231 1230 3265 1264
rect 3231 1162 3265 1196
rect 3055 1048 3089 1059
rect 3231 1093 3265 1128
rect 3319 1366 3353 1446
rect 3319 1298 3353 1332
rect 3319 1230 3353 1264
rect 3319 1162 3353 1196
rect 3319 1111 3353 1128
rect 3518 1423 3586 1446
rect 3518 1389 3535 1423
rect 3569 1389 3586 1423
rect 3518 1349 3586 1389
rect 3518 1315 3535 1349
rect 3569 1315 3586 1349
rect 3518 1275 3586 1315
rect 3518 1241 3535 1275
rect 3569 1241 3586 1275
rect 3518 1201 3586 1241
rect 3518 1167 3535 1201
rect 3569 1167 3586 1201
rect 3518 1127 3586 1167
rect 3231 1048 3265 1059
rect 3518 1093 3535 1127
rect 3569 1093 3586 1127
rect 3518 1053 3586 1093
rect 2556 979 2624 1019
rect 2879 1014 3421 1048
rect 2556 945 2573 979
rect 2607 945 2624 979
rect 2556 905 2624 945
rect 2556 871 2573 905
rect 2607 871 2624 905
rect 2556 822 2624 871
rect 2795 957 2829 973
rect 1662 219 1696 316
rect 1890 313 1958 353
rect 1890 279 1907 313
rect 1941 279 1958 313
rect 1662 169 1696 185
rect 1759 263 1793 279
rect 1759 195 1793 229
rect 1451 125 1485 141
rect 1291 91 1354 125
rect 1388 91 1451 125
rect 1257 75 1291 91
rect 1451 75 1485 91
rect 1565 125 1599 161
rect 1759 125 1793 161
rect 1599 91 1662 125
rect 1696 91 1759 125
rect 1565 75 1599 91
rect 1759 75 1793 91
rect 1890 239 1958 279
rect 1890 205 1907 239
rect 1941 205 1958 239
rect 1890 165 1958 205
rect 1890 131 1907 165
rect 1941 131 1958 165
rect 1890 91 1958 131
rect 1890 57 1907 91
rect 1941 57 1958 91
rect 2046 333 2080 349
rect 2240 333 2274 349
rect 2425 348 2459 649
rect 2795 683 2829 923
rect 2080 299 2143 333
rect 2177 299 2240 333
rect 2046 261 2080 299
rect 2046 193 2080 227
rect 2240 261 2274 299
rect 2046 123 2080 159
rect 2046 73 2080 89
rect 2143 208 2177 224
rect 1890 34 1958 57
rect 2143 34 2177 174
rect 2240 193 2274 227
rect 2337 314 2459 348
rect 2556 461 2624 544
rect 2556 427 2573 461
rect 2607 427 2624 461
rect 2556 387 2624 427
rect 2556 353 2573 387
rect 2607 353 2624 387
rect 2795 433 2829 649
rect 2795 383 2829 399
rect 3017 957 3051 973
rect 3017 905 3051 923
rect 3017 433 3051 871
rect 3017 383 3051 399
rect 3239 957 3273 973
rect 3239 461 3273 923
rect 3239 383 3273 399
rect 3387 831 3421 1014
rect 3518 1019 3535 1053
rect 3569 1019 3586 1053
rect 3753 1366 3787 1446
rect 3753 1298 3787 1332
rect 3753 1230 3787 1264
rect 3753 1162 3787 1196
rect 3753 1093 3787 1128
rect 3753 1043 3787 1059
rect 3841 1366 3875 1404
rect 3841 1298 3875 1332
rect 3841 1230 3875 1264
rect 3841 1162 3875 1196
rect 3841 1093 3875 1128
rect 3929 1366 3963 1446
rect 3929 1298 3963 1332
rect 3929 1230 3963 1264
rect 3929 1162 3963 1196
rect 3929 1111 3963 1128
rect 4017 1366 4051 1404
rect 4017 1298 4051 1332
rect 4017 1230 4051 1264
rect 4017 1162 4051 1196
rect 3841 1048 3875 1059
rect 4017 1093 4051 1128
rect 4105 1366 4139 1446
rect 4105 1298 4139 1332
rect 4105 1230 4139 1264
rect 4105 1162 4139 1196
rect 4105 1111 4139 1128
rect 4193 1366 4227 1404
rect 4193 1298 4227 1332
rect 4193 1230 4227 1264
rect 4193 1162 4227 1196
rect 4017 1048 4051 1059
rect 4193 1093 4227 1128
rect 4281 1366 4315 1446
rect 4281 1298 4315 1332
rect 4281 1230 4315 1264
rect 4281 1162 4315 1196
rect 4281 1111 4315 1128
rect 4480 1423 4548 1446
rect 4480 1389 4497 1423
rect 4531 1389 4548 1423
rect 4480 1349 4548 1389
rect 4480 1315 4497 1349
rect 4531 1315 4548 1349
rect 4480 1275 4548 1315
rect 4480 1241 4497 1275
rect 4531 1241 4548 1275
rect 4480 1201 4548 1241
rect 4480 1167 4497 1201
rect 4531 1167 4548 1201
rect 4480 1127 4548 1167
rect 4193 1048 4227 1059
rect 4480 1093 4497 1127
rect 4531 1093 4548 1127
rect 4480 1053 4548 1093
rect 3518 979 3586 1019
rect 3841 1014 4383 1048
rect 3518 945 3535 979
rect 3569 945 3586 979
rect 3518 905 3586 945
rect 3518 871 3535 905
rect 3569 871 3586 905
rect 3518 822 3586 871
rect 3757 957 3791 973
rect 2337 217 2371 314
rect 2556 313 2624 353
rect 2556 279 2573 313
rect 2607 279 2624 313
rect 2337 167 2371 183
rect 2434 261 2468 277
rect 2434 193 2468 227
rect 2240 123 2274 159
rect 2434 123 2468 159
rect 2274 89 2337 123
rect 2371 89 2434 123
rect 2240 73 2274 89
rect 2434 73 2468 89
rect 2556 239 2624 279
rect 2556 205 2573 239
rect 2607 205 2624 239
rect 2556 165 2624 205
rect 2556 131 2573 165
rect 2607 131 2624 165
rect 2556 91 2624 131
rect 2556 57 2573 91
rect 2607 57 2624 91
rect 2691 335 2725 351
rect 2885 335 2919 351
rect 3079 335 3113 351
rect 2725 301 2788 335
rect 2822 301 2885 335
rect 2919 301 2982 335
rect 3016 301 3079 335
rect 2691 263 2725 301
rect 2691 195 2725 229
rect 2885 263 2919 301
rect 3079 285 3113 301
rect 3193 335 3227 351
rect 3387 350 3421 797
rect 3757 757 3791 923
rect 3193 263 3227 301
rect 2691 125 2725 161
rect 2691 75 2725 91
rect 2788 210 2822 226
rect 2556 34 2624 57
rect 2788 34 2822 176
rect 2885 195 2919 229
rect 2983 216 3017 232
rect 3193 216 3227 229
rect 3017 195 3227 216
rect 3017 182 3193 195
rect 2983 166 3017 182
rect 2885 125 2919 161
rect 3290 316 3421 350
rect 3518 461 3586 544
rect 3518 427 3535 461
rect 3569 427 3586 461
rect 3518 387 3586 427
rect 3518 353 3535 387
rect 3569 353 3586 387
rect 3757 433 3791 723
rect 3757 383 3791 399
rect 3979 957 4013 973
rect 3979 461 4013 923
rect 3979 383 4013 399
rect 4201 957 4235 973
rect 4201 757 4235 923
rect 4201 433 4235 723
rect 4201 383 4235 399
rect 4349 683 4383 1014
rect 4480 1019 4497 1053
rect 4531 1019 4548 1053
rect 4655 1366 4689 1446
rect 4655 1298 4689 1332
rect 4655 1230 4689 1264
rect 4655 1162 4689 1196
rect 4655 1093 4689 1128
rect 4655 1027 4689 1059
rect 4743 1366 4777 1404
rect 4743 1298 4777 1332
rect 4743 1230 4777 1264
rect 4743 1162 4777 1196
rect 4743 1093 4777 1128
rect 4831 1366 4865 1446
rect 4831 1298 4865 1332
rect 4831 1230 4865 1264
rect 4831 1162 4865 1196
rect 4831 1111 4865 1128
rect 4919 1366 4953 1404
rect 4919 1298 4953 1332
rect 4919 1230 4953 1264
rect 4919 1162 4953 1196
rect 4743 1057 4777 1059
rect 4919 1093 4953 1128
rect 5007 1366 5041 1446
rect 5007 1298 5041 1332
rect 5007 1230 5041 1264
rect 5007 1162 5041 1196
rect 5007 1111 5041 1128
rect 5146 1423 5214 1446
rect 5146 1389 5163 1423
rect 5197 1389 5214 1423
rect 5146 1349 5214 1389
rect 5146 1315 5163 1349
rect 5197 1315 5214 1349
rect 5146 1275 5214 1315
rect 5146 1241 5163 1275
rect 5197 1241 5214 1275
rect 5146 1201 5214 1241
rect 5146 1167 5163 1201
rect 5197 1167 5214 1201
rect 5146 1127 5214 1167
rect 4919 1057 4953 1059
rect 5146 1093 5163 1127
rect 5197 1093 5214 1127
rect 4743 1023 5049 1057
rect 4480 979 4548 1019
rect 4480 945 4497 979
rect 4531 945 4548 979
rect 4480 905 4548 945
rect 4480 871 4497 905
rect 4531 871 4548 905
rect 4480 822 4548 871
rect 4719 957 4753 973
rect 4873 957 4907 973
rect 3290 219 3324 316
rect 3518 313 3586 353
rect 3518 279 3535 313
rect 3569 279 3586 313
rect 3290 169 3324 185
rect 3387 263 3421 279
rect 3387 195 3421 229
rect 3079 125 3113 141
rect 2919 91 2982 125
rect 3016 91 3079 125
rect 2885 75 2919 91
rect 3079 75 3113 91
rect 3193 125 3227 161
rect 3387 125 3421 161
rect 3227 91 3290 125
rect 3324 91 3387 125
rect 3193 75 3227 91
rect 3387 75 3421 91
rect 3518 239 3586 279
rect 3518 205 3535 239
rect 3569 205 3586 239
rect 3518 165 3586 205
rect 3518 131 3535 165
rect 3569 131 3586 165
rect 3518 91 3586 131
rect 3518 57 3535 91
rect 3569 57 3586 91
rect 3653 335 3687 351
rect 3847 335 3881 351
rect 4041 335 4075 351
rect 3687 301 3750 335
rect 3784 301 3847 335
rect 3881 301 3944 335
rect 3978 301 4041 335
rect 3653 263 3687 301
rect 3653 195 3687 229
rect 3847 263 3881 301
rect 4041 285 4075 301
rect 4155 335 4189 351
rect 4349 350 4383 649
rect 4719 683 4753 923
rect 4155 263 4189 301
rect 3653 125 3687 161
rect 3653 75 3687 91
rect 3750 210 3784 226
rect 3518 34 3586 57
rect 3750 34 3784 176
rect 3847 195 3881 229
rect 3945 216 3979 232
rect 4155 216 4189 229
rect 3979 195 4189 216
rect 3979 182 4155 195
rect 3945 166 3979 182
rect 3847 125 3881 161
rect 4252 316 4383 350
rect 4480 461 4548 544
rect 4480 427 4497 461
rect 4531 427 4548 461
rect 4480 387 4548 427
rect 4480 353 4497 387
rect 4531 353 4548 387
rect 4719 433 4753 649
rect 4719 383 4753 399
rect 4867 923 4873 942
rect 4867 907 4907 923
rect 4867 831 4901 907
rect 4867 433 4901 797
rect 4867 383 4901 399
rect 5015 757 5049 1023
rect 5146 1053 5214 1093
rect 5146 1019 5163 1053
rect 5197 1019 5214 1053
rect 5146 979 5214 1019
rect 5146 945 5163 979
rect 5197 945 5214 979
rect 5146 905 5214 945
rect 5146 871 5163 905
rect 5197 871 5214 905
rect 5146 822 5214 871
rect 4252 219 4286 316
rect 4480 313 4548 353
rect 4480 279 4497 313
rect 4531 279 4548 313
rect 4252 169 4286 185
rect 4349 263 4383 279
rect 4349 195 4383 229
rect 4041 125 4075 141
rect 3881 91 3944 125
rect 3978 91 4041 125
rect 3847 75 3881 91
rect 4041 75 4075 91
rect 4155 125 4189 161
rect 4349 125 4383 161
rect 4189 91 4252 125
rect 4286 91 4349 125
rect 4155 75 4189 91
rect 4349 75 4383 91
rect 4480 239 4548 279
rect 4480 205 4497 239
rect 4531 205 4548 239
rect 4480 165 4548 205
rect 4480 131 4497 165
rect 4531 131 4548 165
rect 4480 91 4548 131
rect 4480 57 4497 91
rect 4531 57 4548 91
rect 4636 333 4670 349
rect 4830 333 4864 349
rect 5015 348 5049 723
rect 4670 299 4733 333
rect 4767 299 4830 333
rect 4636 261 4670 299
rect 4636 193 4670 227
rect 4830 261 4864 299
rect 4636 123 4670 159
rect 4636 73 4670 89
rect 4733 208 4767 224
rect 4480 34 4548 57
rect 4733 34 4767 174
rect 4830 193 4864 227
rect 4927 314 5049 348
rect 5146 461 5214 544
rect 5146 427 5163 461
rect 5197 427 5214 461
rect 5146 387 5214 427
rect 5146 353 5163 387
rect 5197 353 5214 387
rect 4927 217 4961 314
rect 5146 313 5214 353
rect 5146 279 5163 313
rect 5197 279 5214 313
rect 4927 167 4961 183
rect 5024 261 5058 277
rect 5024 193 5058 227
rect 4830 123 4864 159
rect 5024 123 5058 159
rect 4864 89 4927 123
rect 4961 89 5024 123
rect 4830 73 4864 89
rect 5024 73 5058 89
rect 5146 239 5214 279
rect 5146 205 5163 239
rect 5197 205 5214 239
rect 5146 165 5214 205
rect 5146 131 5163 165
rect 5197 131 5214 165
rect 5146 91 5214 131
rect 5146 57 5163 91
rect 5197 57 5214 91
rect 5146 34 5214 57
rect -34 17 5214 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5214 17
rect -34 -34 5214 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 205 797 239 831
rect 427 871 461 905
rect 649 649 683 683
rect 797 723 831 757
rect 1167 723 1201 757
rect 1611 433 1645 461
rect 1611 427 1645 433
rect 1759 649 1793 683
rect 2129 649 2163 683
rect 2277 797 2311 831
rect 2425 649 2459 683
rect 2795 649 2829 683
rect 3017 871 3051 905
rect 3239 433 3273 461
rect 3239 427 3273 433
rect 3387 797 3421 831
rect 3757 723 3791 757
rect 3979 433 4013 461
rect 3979 427 4013 433
rect 4201 723 4235 757
rect 4349 649 4383 683
rect 4719 649 4753 683
rect 4867 797 4901 831
rect 5015 723 5049 757
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
<< metal1 >>
rect -34 1497 5214 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5214 1497
rect -34 1446 5214 1463
rect 421 905 467 911
rect 3011 905 3057 911
rect 415 871 427 905
rect 461 871 3017 905
rect 3051 871 3063 905
rect 421 865 467 871
rect 3011 865 3057 871
rect 199 831 245 837
rect 2271 831 2317 837
rect 3381 831 3427 837
rect 4861 831 4907 837
rect 193 797 205 831
rect 239 797 2277 831
rect 2311 797 3387 831
rect 3421 797 4867 831
rect 4901 797 4913 831
rect 199 791 245 797
rect 2271 791 2317 797
rect 3381 791 3427 797
rect 4861 791 4907 797
rect 791 757 837 763
rect 1161 757 1207 763
rect 3751 757 3797 763
rect 4195 757 4241 763
rect 5009 757 5055 763
rect 785 723 797 757
rect 831 723 1167 757
rect 1201 723 3757 757
rect 3791 723 3803 757
rect 4189 723 4201 757
rect 4235 723 5015 757
rect 5049 723 5061 757
rect 791 717 837 723
rect 1161 717 1207 723
rect 3751 717 3797 723
rect 4195 717 4241 723
rect 5009 717 5055 723
rect 643 683 689 689
rect 1753 683 1799 689
rect 2123 683 2169 689
rect 2419 683 2465 689
rect 2789 683 2835 689
rect 4343 683 4389 689
rect 4713 683 4759 689
rect 637 649 649 683
rect 683 649 1759 683
rect 1793 649 2129 683
rect 2163 649 2175 683
rect 2413 649 2425 683
rect 2459 649 2795 683
rect 2829 649 2841 683
rect 4337 649 4349 683
rect 4383 649 4719 683
rect 4753 649 4765 683
rect 643 643 689 649
rect 1753 643 1799 649
rect 2123 643 2169 649
rect 2419 643 2465 649
rect 2789 643 2835 649
rect 4343 643 4389 649
rect 4713 643 4759 649
rect 1605 461 1651 467
rect 3233 461 3279 467
rect 3973 461 4019 467
rect 1599 427 1611 461
rect 1645 427 3239 461
rect 3273 427 3979 461
rect 4013 427 4025 461
rect 1605 421 1651 427
rect 3233 421 3279 427
rect 3973 421 4019 427
rect -34 17 5214 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5214 17
rect -34 -34 5214 -17
<< labels >>
rlabel metal1 4349 649 4383 683 1 QN
port 1 n
rlabel metal1 4349 871 4383 905 1 QN
port 2 n
rlabel metal1 4349 945 4383 979 1 QN
port 3 n
rlabel metal1 4349 575 4383 609 1 QN
port 4 n
rlabel metal1 4349 501 4383 535 1 QN
port 5 n
rlabel metal1 4349 427 4383 461 1 QN
port 6 n
rlabel metal1 4719 427 4753 461 1 QN
port 7 n
rlabel metal1 4719 501 4753 535 1 QN
port 8 n
rlabel metal1 4719 575 4753 609 1 QN
port 9 n
rlabel metal1 4719 649 4753 683 1 QN
port 10 n
rlabel metal1 4719 871 4753 905 1 QN
port 11 n
rlabel metal1 1389 501 1423 535 1 D
port 12 n
rlabel metal1 1389 575 1423 609 1 D
port 13 n
rlabel metal1 427 871 461 905 1 CLK
port 14 n
rlabel metal1 427 723 461 757 1 CLK
port 15 n
rlabel metal1 427 649 461 683 1 CLK
port 16 n
rlabel metal1 427 575 461 609 1 CLK
port 17 n
rlabel metal1 427 501 461 535 1 CLK
port 18 n
rlabel metal1 3017 649 3051 683 1 CLK
port 19 n
rlabel metal1 3017 575 3051 609 1 CLK
port 20 n
rlabel metal1 3017 501 3051 535 1 CLK
port 21 n
rlabel metal1 3017 871 3051 905 1 CLK
port 22 n
rlabel metal1 1611 427 1645 461 1 RN
port 23 n
rlabel metal1 1611 501 1645 535 1 RN
port 24 n
rlabel metal1 1611 575 1645 609 1 RN
port 25 n
rlabel metal1 3979 575 4013 609 1 RN
port 26 n
rlabel metal1 3979 501 4013 535 1 RN
port 27 n
rlabel metal1 3979 427 4013 461 1 RN
port 28 n
rlabel metal1 3979 649 4013 683 1 RN
port 29 n
rlabel metal1 3979 723 4013 757 1 RN
port 30 n
rlabel metal1 3239 427 3273 461 1 RN
port 31 n
rlabel metal1 3239 501 3273 535 1 RN
port 32 n
rlabel metal1 3239 575 3273 609 1 RN
port 33 n
rlabel metal1 3239 649 3273 683 1 RN
port 34 n
rlabel metal1 3979 871 4013 905 1 RN
port 35 n
rlabel metal1 3239 871 3273 905 1 RN
port 36 n
rlabel metal1 -34 1446 5214 1514 1 VPWR
port 37 n
rlabel metal1 -34 -34 5214 34 1 VGND
port 38 n
rlabel nwell 57 1463 91 1497 1 VPB
port 39 n
rlabel pwell 57 -17 91 17 1 VNB
port 40 n
<< end >>
