// File: pmos2_1.spi.PMOS2_1.pxi
// Created: Tue Oct 15 16:00:29 2024
// 
simulator lang=spectre
x_PM_PMOS2_1\%noxref_4 ( N_noxref_4_M0_noxref_g N_noxref_4_M1_noxref_g \
 N_noxref_4_c_18_n )  PM_PMOS2_1\%noxref_4
cc_1 ( noxref_1 noxref_2 ) capacitor c=0.0527767f //x=0.44 //y=-1.995 \
 //x2=0.87 //y2=-1.995
cc_2 ( noxref_1 noxref_3 ) capacitor c=0.00561178f //x=0.44 //y=-1.995 \
 //x2=1.31 //y2=-1.995
cc_3 ( noxref_1 N_noxref_4_M0_noxref_g ) capacitor c=0.0245018f //x=0.44 \
 //y=-1.995 //x2=0.795 //y2=-0.995
cc_4 ( noxref_2 noxref_3 ) capacitor c=0.0527767f //x=0.87 //y=-1.995 \
 //x2=1.31 //y2=-1.995
cc_5 ( noxref_2 N_noxref_4_M0_noxref_g ) capacitor c=0.00925495f //x=0.87 \
 //y=-1.995 //x2=0.795 //y2=-0.995
cc_6 ( noxref_2 N_noxref_4_M1_noxref_g ) capacitor c=0.00925495f //x=0.87 \
 //y=-1.995 //x2=1.235 //y2=-0.995
cc_7 ( noxref_2 N_noxref_4_c_18_n ) capacitor c=0.00280229f //x=0.87 \
 //y=-1.995 //x2=1.16 //y2=-2.225
cc_8 ( noxref_3 N_noxref_4_M1_noxref_g ) capacitor c=0.0245018f //x=1.31 \
 //y=-1.995 //x2=1.235 //y2=-0.995
