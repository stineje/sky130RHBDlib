// File: DFFSNQNX1.spi.DFFSNQNX1.pxi
// Created: Tue Oct 15 15:46:54 2024
// 
simulator lang=spectre
x_PM_DFFSNQNX1\%GND ( GND N_GND_c_8_p N_GND_c_134_p N_GND_c_2_p N_GND_c_9_p \
 N_GND_c_10_p N_GND_c_15_p N_GND_c_16_p N_GND_c_42_p N_GND_c_53_p N_GND_c_60_p \
 N_GND_c_74_p N_GND_c_81_p N_GND_c_89_p N_GND_c_1_p N_GND_c_3_p N_GND_c_4_p \
 N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p N_GND_M0_noxref_d N_GND_M2_noxref_d \
 N_GND_M5_noxref_d N_GND_M8_noxref_d N_GND_M10_noxref_d N_GND_M12_noxref_d )  \
 PM_DFFSNQNX1\%GND
x_PM_DFFSNQNX1\%VDD ( VDD N_VDD_c_295_p N_VDD_c_296_p N_VDD_c_297_p \
 N_VDD_c_399_p N_VDD_c_400_p N_VDD_c_312_p N_VDD_c_389_p N_VDD_c_426_p \
 N_VDD_c_374_p N_VDD_c_375_p N_VDD_c_316_p N_VDD_c_337_p N_VDD_c_343_p \
 N_VDD_c_347_p N_VDD_c_378_p N_VDD_c_351_p N_VDD_c_393_p N_VDD_c_407_p \
 N_VDD_c_408_p N_VDD_c_409_p N_VDD_c_465_p N_VDD_c_475_p N_VDD_c_500_p \
 N_VDD_c_531_p N_VDD_c_287_n N_VDD_c_288_n N_VDD_c_289_n N_VDD_c_290_n \
 N_VDD_c_291_n N_VDD_c_292_n N_VDD_c_293_n N_VDD_M15_noxref_s \
 N_VDD_M16_noxref_d N_VDD_M18_noxref_d N_VDD_M19_noxref_s N_VDD_M20_noxref_d \
 N_VDD_M22_noxref_d N_VDD_M24_noxref_d N_VDD_M25_noxref_s N_VDD_M26_noxref_d \
 N_VDD_M28_noxref_d N_VDD_M30_noxref_d N_VDD_M31_noxref_s N_VDD_M32_noxref_d \
 N_VDD_M34_noxref_d N_VDD_M35_noxref_s N_VDD_M36_noxref_d N_VDD_M38_noxref_d \
 N_VDD_M39_noxref_s N_VDD_M40_noxref_d N_VDD_M42_noxref_d N_VDD_M44_noxref_d ) \
 PM_DFFSNQNX1\%VDD
x_PM_DFFSNQNX1\%noxref_3 ( N_noxref_3_c_591_n N_noxref_3_c_595_n \
 N_noxref_3_c_597_n N_noxref_3_c_601_n N_noxref_3_c_632_n N_noxref_3_c_636_n \
 N_noxref_3_c_638_n N_noxref_3_c_603_n N_noxref_3_c_710_p N_noxref_3_c_604_n \
 N_noxref_3_c_606_n N_noxref_3_c_607_n N_noxref_3_c_740_p \
 N_noxref_3_M2_noxref_g N_noxref_3_M5_noxref_g N_noxref_3_M19_noxref_g \
 N_noxref_3_M20_noxref_g N_noxref_3_M25_noxref_g N_noxref_3_M26_noxref_g \
 N_noxref_3_c_608_n N_noxref_3_c_610_n N_noxref_3_c_611_n N_noxref_3_c_612_n \
 N_noxref_3_c_613_n N_noxref_3_c_614_n N_noxref_3_c_615_n N_noxref_3_c_617_n \
 N_noxref_3_c_687_p N_noxref_3_c_657_n N_noxref_3_c_618_n N_noxref_3_c_620_n \
 N_noxref_3_c_621_n N_noxref_3_c_622_n N_noxref_3_c_623_n N_noxref_3_c_624_n \
 N_noxref_3_c_625_n N_noxref_3_c_627_n N_noxref_3_c_675_p N_noxref_3_c_659_n \
 N_noxref_3_M1_noxref_d N_noxref_3_M15_noxref_d N_noxref_3_M17_noxref_d )  \
 PM_DFFSNQNX1\%noxref_3
x_PM_DFFSNQNX1\%noxref_4 ( N_noxref_4_c_831_n N_noxref_4_c_832_n \
 N_noxref_4_c_847_n N_noxref_4_c_851_n N_noxref_4_c_853_n N_noxref_4_c_857_n \
 N_noxref_4_c_833_n N_noxref_4_c_926_p N_noxref_4_c_834_n N_noxref_4_c_835_n \
 N_noxref_4_c_936_p N_noxref_4_c_946_p N_noxref_4_M8_noxref_g \
 N_noxref_4_M31_noxref_g N_noxref_4_M32_noxref_g N_noxref_4_c_836_n \
 N_noxref_4_c_838_n N_noxref_4_c_839_n N_noxref_4_c_840_n N_noxref_4_c_841_n \
 N_noxref_4_c_842_n N_noxref_4_c_843_n N_noxref_4_c_845_n N_noxref_4_c_869_n \
 N_noxref_4_M7_noxref_d N_noxref_4_M25_noxref_d N_noxref_4_M27_noxref_d \
 N_noxref_4_M29_noxref_d )  PM_DFFSNQNX1\%noxref_4
x_PM_DFFSNQNX1\%CLK ( N_CLK_c_994_n N_CLK_c_1005_n CLK CLK CLK CLK CLK CLK CLK \
 CLK N_CLK_c_991_n N_CLK_c_1054_n N_CLK_c_992_n N_CLK_M3_noxref_g \
 N_CLK_M9_noxref_g N_CLK_M21_noxref_g N_CLK_M22_noxref_g N_CLK_M33_noxref_g \
 N_CLK_M34_noxref_g N_CLK_c_1034_n N_CLK_c_1037_n N_CLK_c_1168_p \
 N_CLK_c_1175_p N_CLK_c_1039_n N_CLK_c_1040_n N_CLK_c_1041_n N_CLK_c_1042_n \
 N_CLK_c_1095_p N_CLK_c_1063_n N_CLK_c_1066_n N_CLK_c_1068_n N_CLK_c_1082_p \
 N_CLK_c_1153_p N_CLK_c_1101_p N_CLK_c_1071_n N_CLK_c_1072_n N_CLK_c_1045_n \
 N_CLK_c_1073_n N_CLK_c_1133_p N_CLK_c_1075_n )  PM_DFFSNQNX1\%CLK
x_PM_DFFSNQNX1\%noxref_6 ( N_noxref_6_c_1189_n N_noxref_6_c_1191_n \
 N_noxref_6_c_1215_n N_noxref_6_c_1224_n N_noxref_6_c_1284_n \
 N_noxref_6_c_1192_n N_noxref_6_c_1227_n N_noxref_6_c_1231_n \
 N_noxref_6_c_1233_n N_noxref_6_c_1237_n N_noxref_6_c_1194_n \
 N_noxref_6_c_1293_n N_noxref_6_c_1336_n N_noxref_6_c_1195_n \
 N_noxref_6_c_1339_n N_noxref_6_c_1375_p N_noxref_6_c_1244_n \
 N_noxref_6_c_1294_n N_noxref_6_M1_noxref_g N_noxref_6_M10_noxref_g \
 N_noxref_6_M17_noxref_g N_noxref_6_M18_noxref_g N_noxref_6_M35_noxref_g \
 N_noxref_6_M36_noxref_g N_noxref_6_c_1300_n N_noxref_6_c_1301_n \
 N_noxref_6_c_1302_n N_noxref_6_c_1303_n N_noxref_6_c_1305_n \
 N_noxref_6_c_1306_n N_noxref_6_c_1308_n N_noxref_6_c_1309_n \
 N_noxref_6_c_1196_n N_noxref_6_c_1198_n N_noxref_6_c_1199_n \
 N_noxref_6_c_1200_n N_noxref_6_c_1201_n N_noxref_6_c_1202_n \
 N_noxref_6_c_1203_n N_noxref_6_c_1205_n N_noxref_6_c_1311_n \
 N_noxref_6_c_1312_n N_noxref_6_c_1314_n N_noxref_6_c_1254_n \
 N_noxref_6_M4_noxref_d N_noxref_6_M19_noxref_d N_noxref_6_M21_noxref_d \
 N_noxref_6_M23_noxref_d )  PM_DFFSNQNX1\%noxref_6
x_PM_DFFSNQNX1\%QN ( N_QN_c_1475_n N_QN_c_1531_p QN QN QN QN QN QN QN QN QN \
 N_QN_c_1494_n N_QN_c_1498_n N_QN_c_1500_n N_QN_c_1477_n N_QN_c_1533_p \
 N_QN_c_1478_n N_QN_c_1589_p N_QN_M12_noxref_g N_QN_M39_noxref_g \
 N_QN_M40_noxref_g N_QN_c_1479_n N_QN_c_1481_n N_QN_c_1482_n N_QN_c_1483_n \
 N_QN_c_1484_n N_QN_c_1485_n N_QN_c_1486_n N_QN_c_1488_n N_QN_c_1540_p \
 N_QN_c_1510_n N_QN_M11_noxref_d N_QN_M35_noxref_d N_QN_M37_noxref_d )  \
 PM_DFFSNQNX1\%QN
x_PM_DFFSNQNX1\%SN ( N_SN_c_1620_n N_SN_c_1630_n SN SN SN SN SN SN SN SN SN \
 N_SN_c_1631_n N_SN_c_1632_n N_SN_M6_noxref_g N_SN_M13_noxref_g \
 N_SN_M27_noxref_g N_SN_M28_noxref_g N_SN_M41_noxref_g N_SN_M42_noxref_g \
 N_SN_c_1655_n N_SN_c_1658_n N_SN_c_1798_p N_SN_c_1806_p N_SN_c_1660_n \
 N_SN_c_1661_n N_SN_c_1662_n N_SN_c_1663_n N_SN_c_1680_n N_SN_c_1709_n \
 N_SN_c_1712_n N_SN_c_1834_p N_SN_c_1841_p N_SN_c_1714_n N_SN_c_1715_n \
 N_SN_c_1716_n N_SN_c_1717_n N_SN_c_1730_p N_SN_c_1665_n N_SN_c_1719_n )  \
 PM_DFFSNQNX1\%SN
x_PM_DFFSNQNX1\%noxref_9 ( N_noxref_9_c_1846_n N_noxref_9_c_1902_n \
 N_noxref_9_c_1848_n N_noxref_9_c_1912_n N_noxref_9_c_1849_n \
 N_noxref_9_c_1949_n N_noxref_9_c_1850_n N_noxref_9_c_1851_n \
 N_noxref_9_c_1864_n N_noxref_9_c_1868_n N_noxref_9_c_1870_n \
 N_noxref_9_c_1852_n N_noxref_9_c_2065_n N_noxref_9_c_1853_n \
 N_noxref_9_c_1854_n N_noxref_9_c_1972_n N_noxref_9_M4_noxref_g \
 N_noxref_9_M7_noxref_g N_noxref_9_M14_noxref_g N_noxref_9_M23_noxref_g \
 N_noxref_9_M24_noxref_g N_noxref_9_M29_noxref_g N_noxref_9_M30_noxref_g \
 N_noxref_9_M43_noxref_g N_noxref_9_M44_noxref_g N_noxref_9_c_1976_n \
 N_noxref_9_c_1977_n N_noxref_9_c_1978_n N_noxref_9_c_2028_n \
 N_noxref_9_c_2029_n N_noxref_9_c_2031_n N_noxref_9_c_2032_n \
 N_noxref_9_c_1927_n N_noxref_9_c_1928_n N_noxref_9_c_1929_n \
 N_noxref_9_c_1930_n N_noxref_9_c_1931_n N_noxref_9_c_1933_n \
 N_noxref_9_c_1934_n N_noxref_9_c_2081_n N_noxref_9_c_2082_n \
 N_noxref_9_c_2083_n N_noxref_9_c_2126_p N_noxref_9_c_2111_p \
 N_noxref_9_c_2128_p N_noxref_9_c_2112_p N_noxref_9_c_1907_n \
 N_noxref_9_c_1981_n N_noxref_9_c_1982_n N_noxref_9_c_1936_n \
 N_noxref_9_c_1937_n N_noxref_9_c_1939_n N_noxref_9_c_2092_n \
 N_noxref_9_c_2095_n N_noxref_9_c_2096_n N_noxref_9_M9_noxref_d \
 N_noxref_9_M31_noxref_d N_noxref_9_M33_noxref_d )  PM_DFFSNQNX1\%noxref_9
x_PM_DFFSNQNX1\%noxref_10 ( N_noxref_10_c_2170_n N_noxref_10_c_2213_n \
 N_noxref_10_c_2214_n N_noxref_10_c_2172_n N_noxref_10_c_2179_n \
 N_noxref_10_c_2183_n N_noxref_10_c_2185_n N_noxref_10_c_2189_n \
 N_noxref_10_c_2174_n N_noxref_10_c_2335_p N_noxref_10_c_2193_n \
 N_noxref_10_c_2280_n N_noxref_10_c_2304_n N_noxref_10_M11_noxref_g \
 N_noxref_10_M37_noxref_g N_noxref_10_M38_noxref_g N_noxref_10_c_2222_n \
 N_noxref_10_c_2225_n N_noxref_10_c_2227_n N_noxref_10_c_2257_n \
 N_noxref_10_c_2259_n N_noxref_10_c_2260_n N_noxref_10_c_2230_n \
 N_noxref_10_c_2231_n N_noxref_10_c_2232_n N_noxref_10_c_2266_n \
 N_noxref_10_c_2234_n N_noxref_10_M14_noxref_d N_noxref_10_M39_noxref_d \
 N_noxref_10_M41_noxref_d N_noxref_10_M43_noxref_d )  PM_DFFSNQNX1\%noxref_10
x_PM_DFFSNQNX1\%D ( D D D D D D D N_D_c_2340_n N_D_M0_noxref_g \
 N_D_M15_noxref_g N_D_M16_noxref_g N_D_c_2341_n N_D_c_2343_n N_D_c_2344_n \
 N_D_c_2345_n N_D_c_2346_n N_D_c_2347_n N_D_c_2348_n N_D_c_2350_n N_D_c_2358_n \
 )  PM_DFFSNQNX1\%D
x_PM_DFFSNQNX1\%noxref_12 ( N_noxref_12_c_2416_n N_noxref_12_c_2397_n \
 N_noxref_12_c_2401_n N_noxref_12_c_2404_n N_noxref_12_c_2405_n \
 N_noxref_12_c_2408_n N_noxref_12_M0_noxref_s )  PM_DFFSNQNX1\%noxref_12
x_PM_DFFSNQNX1\%noxref_13 ( N_noxref_13_c_2461_n N_noxref_13_c_2445_n \
 N_noxref_13_c_2449_n N_noxref_13_c_2452_n N_noxref_13_c_2472_n \
 N_noxref_13_M2_noxref_s )  PM_DFFSNQNX1\%noxref_13
x_PM_DFFSNQNX1\%noxref_14 ( N_noxref_14_c_2497_n N_noxref_14_c_2499_n \
 N_noxref_14_c_2502_n N_noxref_14_c_2505_n N_noxref_14_c_2528_n \
 N_noxref_14_M3_noxref_d N_noxref_14_M4_noxref_s )  PM_DFFSNQNX1\%noxref_14
x_PM_DFFSNQNX1\%noxref_15 ( N_noxref_15_c_2566_n N_noxref_15_c_2550_n \
 N_noxref_15_c_2554_n N_noxref_15_c_2557_n N_noxref_15_c_2583_n \
 N_noxref_15_M5_noxref_s )  PM_DFFSNQNX1\%noxref_15
x_PM_DFFSNQNX1\%noxref_16 ( N_noxref_16_c_2604_n N_noxref_16_c_2606_n \
 N_noxref_16_c_2609_n N_noxref_16_c_2612_n N_noxref_16_c_2620_n \
 N_noxref_16_M6_noxref_d N_noxref_16_M7_noxref_s )  PM_DFFSNQNX1\%noxref_16
x_PM_DFFSNQNX1\%noxref_17 ( N_noxref_17_c_2676_n N_noxref_17_c_2657_n \
 N_noxref_17_c_2661_n N_noxref_17_c_2664_n N_noxref_17_c_2665_n \
 N_noxref_17_c_2668_n N_noxref_17_M8_noxref_s )  PM_DFFSNQNX1\%noxref_17
x_PM_DFFSNQNX1\%noxref_18 ( N_noxref_18_c_2728_n N_noxref_18_c_2709_n \
 N_noxref_18_c_2713_n N_noxref_18_c_2716_n N_noxref_18_c_2717_n \
 N_noxref_18_c_2720_n N_noxref_18_M10_noxref_s )  PM_DFFSNQNX1\%noxref_18
x_PM_DFFSNQNX1\%noxref_19 ( N_noxref_19_c_2775_n N_noxref_19_c_2761_n \
 N_noxref_19_c_2765_n N_noxref_19_c_2768_n N_noxref_19_c_2791_n \
 N_noxref_19_M12_noxref_s )  PM_DFFSNQNX1\%noxref_19
x_PM_DFFSNQNX1\%noxref_20 ( N_noxref_20_c_2811_n N_noxref_20_c_2813_n \
 N_noxref_20_c_2816_n N_noxref_20_c_2818_n N_noxref_20_c_2839_n \
 N_noxref_20_M13_noxref_d N_noxref_20_M14_noxref_s )  PM_DFFSNQNX1\%noxref_20
cc_1 ( N_GND_c_1_p N_VDD_c_287_n ) capacitor c=0.00989031f //x=23.68 //y=0 \
 //x2=23.68 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_288_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_289_n ) capacitor c=0.00582097f //x=3.33 //y=0 \
 //x2=3.33 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_290_n ) capacitor c=0.0057235f //x=8.14 //y=0 \
 //x2=8.14 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_291_n ) capacitor c=0.0057235f //x=12.95 //y=0 \
 //x2=12.95 //y2=7.4
cc_6 ( N_GND_c_6_p N_VDD_c_292_n ) capacitor c=0.00524516f //x=16.28 //y=0 \
 //x2=16.28 //y2=7.4
cc_7 ( N_GND_c_7_p N_VDD_c_293_n ) capacitor c=0.00802221f //x=19.61 //y=0 \
 //x2=19.61 //y2=7.4
cc_8 ( N_GND_c_8_p N_noxref_3_c_591_n ) capacitor c=0.0139834f //x=23.68 //y=0 \
 //x2=4.295 //y2=2.59
cc_9 ( N_GND_c_9_p N_noxref_3_c_591_n ) capacitor c=0.00230866f //x=3.16 //y=0 \
 //x2=4.295 //y2=2.59
cc_10 ( N_GND_c_10_p N_noxref_3_c_591_n ) capacitor c=0.00221947f //x=4.32 \
 //y=0 //x2=4.295 //y2=2.59
cc_11 ( N_GND_c_3_p N_noxref_3_c_591_n ) capacitor c=0.038878f //x=3.33 //y=0 \
 //x2=4.295 //y2=2.59
cc_12 ( N_GND_c_8_p N_noxref_3_c_595_n ) capacitor c=0.00222479f //x=23.68 \
 //y=0 //x2=2.705 //y2=2.59
cc_13 ( N_GND_c_3_p N_noxref_3_c_595_n ) capacitor c=0.00111411f //x=3.33 \
 //y=0 //x2=2.705 //y2=2.59
cc_14 ( N_GND_c_8_p N_noxref_3_c_597_n ) capacitor c=0.0394349f //x=23.68 \
 //y=0 //x2=9.135 //y2=2.59
cc_15 ( N_GND_c_15_p N_noxref_3_c_597_n ) capacitor c=0.00344363f //x=7.97 \
 //y=0 //x2=9.135 //y2=2.59
cc_16 ( N_GND_c_16_p N_noxref_3_c_597_n ) capacitor c=0.00221947f //x=9.13 \
 //y=0 //x2=9.135 //y2=2.59
cc_17 ( N_GND_c_4_p N_noxref_3_c_597_n ) capacitor c=0.0392112f //x=8.14 //y=0 \
 //x2=9.135 //y2=2.59
cc_18 ( N_GND_c_8_p N_noxref_3_c_601_n ) capacitor c=0.0038075f //x=23.68 \
 //y=0 //x2=4.705 //y2=2.59
cc_19 ( N_GND_c_3_p N_noxref_3_c_601_n ) capacitor c=7.88768e-19 //x=3.33 \
 //y=0 //x2=4.705 //y2=2.59
cc_20 ( N_GND_c_3_p N_noxref_3_c_603_n ) capacitor c=0.0430571f //x=3.33 //y=0 \
 //x2=2.505 //y2=1.655
cc_21 ( N_GND_c_2_p N_noxref_3_c_604_n ) capacitor c=0.00101801f //x=0.74 \
 //y=0 //x2=2.59 //y2=2.59
cc_22 ( N_GND_c_3_p N_noxref_3_c_604_n ) capacitor c=5.56859e-19 //x=3.33 \
 //y=0 //x2=2.59 //y2=2.59
cc_23 ( N_GND_c_3_p N_noxref_3_c_606_n ) capacitor c=0.0150282f //x=3.33 //y=0 \
 //x2=4.44 //y2=2.08
cc_24 ( N_GND_c_4_p N_noxref_3_c_607_n ) capacitor c=0.0147449f //x=8.14 //y=0 \
 //x2=9.25 //y2=2.08
cc_25 ( N_GND_c_10_p N_noxref_3_c_608_n ) capacitor c=0.00132755f //x=4.32 \
 //y=0 //x2=4.14 //y2=0.875
cc_26 ( N_GND_M2_noxref_d N_noxref_3_c_608_n ) capacitor c=0.00211996f \
 //x=4.215 //y=0.875 //x2=4.14 //y2=0.875
cc_27 ( N_GND_M2_noxref_d N_noxref_3_c_610_n ) capacitor c=0.00255985f \
 //x=4.215 //y=0.875 //x2=4.14 //y2=1.22
cc_28 ( N_GND_c_3_p N_noxref_3_c_611_n ) capacitor c=0.00195164f //x=3.33 \
 //y=0 //x2=4.14 //y2=1.53
cc_29 ( N_GND_c_3_p N_noxref_3_c_612_n ) capacitor c=0.0126573f //x=3.33 //y=0 \
 //x2=4.14 //y2=1.915
cc_30 ( N_GND_M2_noxref_d N_noxref_3_c_613_n ) capacitor c=0.0131341f \
 //x=4.215 //y=0.875 //x2=4.515 //y2=0.72
cc_31 ( N_GND_M2_noxref_d N_noxref_3_c_614_n ) capacitor c=0.00193146f \
 //x=4.215 //y=0.875 //x2=4.515 //y2=1.375
cc_32 ( N_GND_c_15_p N_noxref_3_c_615_n ) capacitor c=0.00129018f //x=7.97 \
 //y=0 //x2=4.67 //y2=0.875
cc_33 ( N_GND_M2_noxref_d N_noxref_3_c_615_n ) capacitor c=0.00257848f \
 //x=4.215 //y=0.875 //x2=4.67 //y2=0.875
cc_34 ( N_GND_M2_noxref_d N_noxref_3_c_617_n ) capacitor c=0.00255985f \
 //x=4.215 //y=0.875 //x2=4.67 //y2=1.22
cc_35 ( N_GND_c_16_p N_noxref_3_c_618_n ) capacitor c=0.00132755f //x=9.13 \
 //y=0 //x2=8.95 //y2=0.875
cc_36 ( N_GND_M5_noxref_d N_noxref_3_c_618_n ) capacitor c=0.00211996f \
 //x=9.025 //y=0.875 //x2=8.95 //y2=0.875
cc_37 ( N_GND_M5_noxref_d N_noxref_3_c_620_n ) capacitor c=0.00255985f \
 //x=9.025 //y=0.875 //x2=8.95 //y2=1.22
cc_38 ( N_GND_c_4_p N_noxref_3_c_621_n ) capacitor c=0.00204716f //x=8.14 \
 //y=0 //x2=8.95 //y2=1.53
cc_39 ( N_GND_c_4_p N_noxref_3_c_622_n ) capacitor c=0.0118433f //x=8.14 //y=0 \
 //x2=8.95 //y2=1.915
cc_40 ( N_GND_M5_noxref_d N_noxref_3_c_623_n ) capacitor c=0.0131341f \
 //x=9.025 //y=0.875 //x2=9.325 //y2=0.72
cc_41 ( N_GND_M5_noxref_d N_noxref_3_c_624_n ) capacitor c=0.00193146f \
 //x=9.025 //y=0.875 //x2=9.325 //y2=1.375
cc_42 ( N_GND_c_42_p N_noxref_3_c_625_n ) capacitor c=0.00129018f //x=12.78 \
 //y=0 //x2=9.48 //y2=0.875
cc_43 ( N_GND_M5_noxref_d N_noxref_3_c_625_n ) capacitor c=0.00257848f \
 //x=9.025 //y=0.875 //x2=9.48 //y2=0.875
cc_44 ( N_GND_M5_noxref_d N_noxref_3_c_627_n ) capacitor c=0.00255985f \
 //x=9.025 //y=0.875 //x2=9.48 //y2=1.22
cc_45 ( N_GND_c_2_p N_noxref_3_M1_noxref_d ) capacitor c=8.58106e-19 //x=0.74 \
 //y=0 //x2=1.96 //y2=0.905
cc_46 ( N_GND_c_3_p N_noxref_3_M1_noxref_d ) capacitor c=0.00616547f //x=3.33 \
 //y=0 //x2=1.96 //y2=0.905
cc_47 ( N_GND_M0_noxref_d N_noxref_3_M1_noxref_d ) capacitor c=0.00143464f \
 //x=0.99 //y=0.865 //x2=1.96 //y2=0.905
cc_48 ( N_GND_c_5_p N_noxref_4_c_831_n ) capacitor c=0.026175f //x=12.95 //y=0 \
 //x2=13.945 //y2=2.59
cc_49 ( N_GND_c_5_p N_noxref_4_c_832_n ) capacitor c=0.00102529f //x=12.95 \
 //y=0 //x2=12.325 //y2=2.59
cc_50 ( N_GND_c_5_p N_noxref_4_c_833_n ) capacitor c=0.0401238f //x=12.95 \
 //y=0 //x2=12.125 //y2=1.665
cc_51 ( N_GND_c_5_p N_noxref_4_c_834_n ) capacitor c=5.56859e-19 //x=12.95 \
 //y=0 //x2=12.21 //y2=2.59
cc_52 ( N_GND_c_5_p N_noxref_4_c_835_n ) capacitor c=0.0128176f //x=12.95 \
 //y=0 //x2=14.06 //y2=2.08
cc_53 ( N_GND_c_53_p N_noxref_4_c_836_n ) capacitor c=0.00135046f //x=14.045 \
 //y=0 //x2=13.865 //y2=0.865
cc_54 ( N_GND_M8_noxref_d N_noxref_4_c_836_n ) capacitor c=0.00220047f \
 //x=13.94 //y=0.865 //x2=13.865 //y2=0.865
cc_55 ( N_GND_M8_noxref_d N_noxref_4_c_838_n ) capacitor c=0.00255985f \
 //x=13.94 //y=0.865 //x2=13.865 //y2=1.21
cc_56 ( N_GND_c_5_p N_noxref_4_c_839_n ) capacitor c=0.00189421f //x=12.95 \
 //y=0 //x2=13.865 //y2=1.52
cc_57 ( N_GND_c_5_p N_noxref_4_c_840_n ) capacitor c=0.00992619f //x=12.95 \
 //y=0 //x2=13.865 //y2=1.915
cc_58 ( N_GND_M8_noxref_d N_noxref_4_c_841_n ) capacitor c=0.0131326f \
 //x=13.94 //y=0.865 //x2=14.24 //y2=0.71
cc_59 ( N_GND_M8_noxref_d N_noxref_4_c_842_n ) capacitor c=0.00193127f \
 //x=13.94 //y=0.865 //x2=14.24 //y2=1.365
cc_60 ( N_GND_c_60_p N_noxref_4_c_843_n ) capacitor c=0.00130622f //x=16.11 \
 //y=0 //x2=14.395 //y2=0.865
cc_61 ( N_GND_M8_noxref_d N_noxref_4_c_843_n ) capacitor c=0.00257848f \
 //x=13.94 //y=0.865 //x2=14.395 //y2=0.865
cc_62 ( N_GND_M8_noxref_d N_noxref_4_c_845_n ) capacitor c=0.00255985f \
 //x=13.94 //y=0.865 //x2=14.395 //y2=1.21
cc_63 ( N_GND_c_5_p N_noxref_4_M7_noxref_d ) capacitor c=0.00591582f //x=12.95 \
 //y=0 //x2=11.535 //y2=0.915
cc_64 ( N_GND_c_3_p N_CLK_c_991_n ) capacitor c=7.5188e-19 //x=3.33 //y=0 \
 //x2=5.55 //y2=2.08
cc_65 ( N_GND_c_5_p N_CLK_c_992_n ) capacitor c=9.18594e-19 //x=12.95 //y=0 \
 //x2=14.8 //y2=2.08
cc_66 ( N_GND_c_6_p N_CLK_c_992_n ) capacitor c=0.00110048f //x=16.28 //y=0 \
 //x2=14.8 //y2=2.08
cc_67 ( N_GND_c_8_p N_noxref_6_c_1189_n ) capacitor c=0.00601678f //x=23.68 \
 //y=0 //x2=7.28 //y2=4.07
cc_68 ( N_GND_c_3_p N_noxref_6_c_1189_n ) capacitor c=0.00249386f //x=3.33 \
 //y=0 //x2=7.28 //y2=4.07
cc_69 ( N_GND_c_8_p N_noxref_6_c_1191_n ) capacitor c=0.00138452f //x=23.68 \
 //y=0 //x2=1.965 //y2=4.07
cc_70 ( N_GND_c_2_p N_noxref_6_c_1192_n ) capacitor c=0.00115206f //x=0.74 \
 //y=0 //x2=1.85 //y2=2.08
cc_71 ( N_GND_c_3_p N_noxref_6_c_1192_n ) capacitor c=0.00110672f //x=3.33 \
 //y=0 //x2=1.85 //y2=2.08
cc_72 ( N_GND_c_4_p N_noxref_6_c_1194_n ) capacitor c=0.0425027f //x=8.14 \
 //y=0 //x2=7.315 //y2=1.665
cc_73 ( N_GND_c_6_p N_noxref_6_c_1195_n ) capacitor c=0.0154414f //x=16.28 \
 //y=0 //x2=17.39 //y2=2.08
cc_74 ( N_GND_c_74_p N_noxref_6_c_1196_n ) capacitor c=0.00135046f //x=17.375 \
 //y=0 //x2=17.195 //y2=0.865
cc_75 ( N_GND_M10_noxref_d N_noxref_6_c_1196_n ) capacitor c=0.00220047f \
 //x=17.27 //y=0.865 //x2=17.195 //y2=0.865
cc_76 ( N_GND_M10_noxref_d N_noxref_6_c_1198_n ) capacitor c=0.00255985f \
 //x=17.27 //y=0.865 //x2=17.195 //y2=1.21
cc_77 ( N_GND_c_6_p N_noxref_6_c_1199_n ) capacitor c=0.0018059f //x=16.28 \
 //y=0 //x2=17.195 //y2=1.52
cc_78 ( N_GND_c_6_p N_noxref_6_c_1200_n ) capacitor c=0.0101006f //x=16.28 \
 //y=0 //x2=17.195 //y2=1.915
cc_79 ( N_GND_M10_noxref_d N_noxref_6_c_1201_n ) capacitor c=0.0131326f \
 //x=17.27 //y=0.865 //x2=17.57 //y2=0.71
cc_80 ( N_GND_M10_noxref_d N_noxref_6_c_1202_n ) capacitor c=0.00193127f \
 //x=17.27 //y=0.865 //x2=17.57 //y2=1.365
cc_81 ( N_GND_c_81_p N_noxref_6_c_1203_n ) capacitor c=0.00130622f //x=19.44 \
 //y=0 //x2=17.725 //y2=0.865
cc_82 ( N_GND_M10_noxref_d N_noxref_6_c_1203_n ) capacitor c=0.00257848f \
 //x=17.27 //y=0.865 //x2=17.725 //y2=0.865
cc_83 ( N_GND_M10_noxref_d N_noxref_6_c_1205_n ) capacitor c=0.00255985f \
 //x=17.27 //y=0.865 //x2=17.725 //y2=1.21
cc_84 ( N_GND_c_4_p N_noxref_6_M4_noxref_d ) capacitor c=0.00591582f //x=8.14 \
 //y=0 //x2=6.725 //y2=0.915
cc_85 ( N_GND_c_7_p N_QN_c_1475_n ) capacitor c=0.00949826f //x=19.61 //y=0 \
 //x2=20.605 //y2=2.96
cc_86 ( N_GND_c_6_p QN ) capacitor c=9.64732e-19 //x=16.28 //y=0 //x2=18.87 \
 //y2=2.59
cc_87 ( N_GND_c_7_p N_QN_c_1477_n ) capacitor c=0.0435299f //x=19.61 //y=0 \
 //x2=18.785 //y2=1.655
cc_88 ( N_GND_c_7_p N_QN_c_1478_n ) capacitor c=0.0156304f //x=19.61 //y=0 \
 //x2=20.72 //y2=2.08
cc_89 ( N_GND_c_89_p N_QN_c_1479_n ) capacitor c=0.00132755f //x=20.6 //y=0 \
 //x2=20.42 //y2=0.875
cc_90 ( N_GND_M12_noxref_d N_QN_c_1479_n ) capacitor c=0.00211996f //x=20.495 \
 //y=0.875 //x2=20.42 //y2=0.875
cc_91 ( N_GND_M12_noxref_d N_QN_c_1481_n ) capacitor c=0.00255985f //x=20.495 \
 //y=0.875 //x2=20.42 //y2=1.22
cc_92 ( N_GND_c_7_p N_QN_c_1482_n ) capacitor c=0.00195164f //x=19.61 //y=0 \
 //x2=20.42 //y2=1.53
cc_93 ( N_GND_c_7_p N_QN_c_1483_n ) capacitor c=0.0110952f //x=19.61 //y=0 \
 //x2=20.42 //y2=1.915
cc_94 ( N_GND_M12_noxref_d N_QN_c_1484_n ) capacitor c=0.0131341f //x=20.495 \
 //y=0.875 //x2=20.795 //y2=0.72
cc_95 ( N_GND_M12_noxref_d N_QN_c_1485_n ) capacitor c=0.00193146f //x=20.495 \
 //y=0.875 //x2=20.795 //y2=1.375
cc_96 ( N_GND_c_1_p N_QN_c_1486_n ) capacitor c=0.00129018f //x=23.68 //y=0 \
 //x2=20.95 //y2=0.875
cc_97 ( N_GND_M12_noxref_d N_QN_c_1486_n ) capacitor c=0.00257848f //x=20.495 \
 //y=0.875 //x2=20.95 //y2=0.875
cc_98 ( N_GND_M12_noxref_d N_QN_c_1488_n ) capacitor c=0.00255985f //x=20.495 \
 //y=0.875 //x2=20.95 //y2=1.22
cc_99 ( N_GND_c_6_p N_QN_M11_noxref_d ) capacitor c=8.58106e-19 //x=16.28 \
 //y=0 //x2=18.24 //y2=0.905
cc_100 ( N_GND_c_7_p N_QN_M11_noxref_d ) capacitor c=0.00616547f //x=19.61 \
 //y=0 //x2=18.24 //y2=0.905
cc_101 ( N_GND_M10_noxref_d N_QN_M11_noxref_d ) capacitor c=0.00143464f \
 //x=17.27 //y=0.865 //x2=18.24 //y2=0.905
cc_102 ( N_GND_c_8_p N_SN_c_1620_n ) capacitor c=0.108864f //x=23.68 //y=0 \
 //x2=21.715 //y2=2.22
cc_103 ( N_GND_c_42_p N_SN_c_1620_n ) capacitor c=0.00447829f //x=12.78 //y=0 \
 //x2=21.715 //y2=2.22
cc_104 ( N_GND_c_53_p N_SN_c_1620_n ) capacitor c=0.00347653f //x=14.045 //y=0 \
 //x2=21.715 //y2=2.22
cc_105 ( N_GND_c_60_p N_SN_c_1620_n ) capacitor c=0.00411932f //x=16.11 //y=0 \
 //x2=21.715 //y2=2.22
cc_106 ( N_GND_c_74_p N_SN_c_1620_n ) capacitor c=0.00347653f //x=17.375 //y=0 \
 //x2=21.715 //y2=2.22
cc_107 ( N_GND_c_81_p N_SN_c_1620_n ) capacitor c=0.00411932f //x=19.44 //y=0 \
 //x2=21.715 //y2=2.22
cc_108 ( N_GND_c_89_p N_SN_c_1620_n ) capacitor c=0.00274252f //x=20.6 //y=0 \
 //x2=21.715 //y2=2.22
cc_109 ( N_GND_c_5_p N_SN_c_1620_n ) capacitor c=0.0379964f //x=12.95 //y=0 \
 //x2=21.715 //y2=2.22
cc_110 ( N_GND_c_6_p N_SN_c_1620_n ) capacitor c=0.0430854f //x=16.28 //y=0 \
 //x2=21.715 //y2=2.22
cc_111 ( N_GND_c_7_p N_SN_c_1620_n ) capacitor c=0.0401775f //x=19.61 //y=0 \
 //x2=21.715 //y2=2.22
cc_112 ( N_GND_c_8_p N_SN_c_1630_n ) capacitor c=0.0019104f //x=23.68 //y=0 \
 //x2=10.475 //y2=2.22
cc_113 ( N_GND_c_4_p N_SN_c_1631_n ) capacitor c=9.83618e-19 //x=8.14 //y=0 \
 //x2=10.36 //y2=2.08
cc_114 ( N_GND_c_7_p N_SN_c_1632_n ) capacitor c=5.94159e-19 //x=19.61 //y=0 \
 //x2=21.83 //y2=2.08
cc_115 ( N_GND_c_8_p N_noxref_9_c_1846_n ) capacitor c=0.00925958f //x=23.68 \
 //y=0 //x2=11.355 //y2=3.7
cc_116 ( N_GND_c_4_p N_noxref_9_c_1846_n ) capacitor c=0.0034979f //x=8.14 \
 //y=0 //x2=11.355 //y2=3.7
cc_117 ( N_GND_c_5_p N_noxref_9_c_1848_n ) capacitor c=0.0034979f //x=12.95 \
 //y=0 //x2=15.425 //y2=3.7
cc_118 ( N_GND_c_6_p N_noxref_9_c_1849_n ) capacitor c=0.00390249f //x=16.28 \
 //y=0 //x2=22.825 //y2=3.7
cc_119 ( N_GND_c_4_p N_noxref_9_c_1850_n ) capacitor c=7.88616e-19 //x=8.14 \
 //y=0 //x2=6.66 //y2=2.08
cc_120 ( N_GND_c_5_p N_noxref_9_c_1851_n ) capacitor c=0.00101012f //x=12.95 \
 //y=0 //x2=11.47 //y2=2.08
cc_121 ( N_GND_c_6_p N_noxref_9_c_1852_n ) capacitor c=0.0432305f //x=16.28 \
 //y=0 //x2=15.455 //y2=1.655
cc_122 ( N_GND_c_5_p N_noxref_9_c_1853_n ) capacitor c=9.64732e-19 //x=12.95 \
 //y=0 //x2=15.54 //y2=3.7
cc_123 ( N_GND_c_1_p N_noxref_9_c_1854_n ) capacitor c=0.00128267f //x=23.68 \
 //y=0 //x2=22.94 //y2=2.08
cc_124 ( N_GND_c_5_p N_noxref_9_M9_noxref_d ) capacitor c=8.58106e-19 \
 //x=12.95 //y=0 //x2=14.91 //y2=0.905
cc_125 ( N_GND_c_6_p N_noxref_9_M9_noxref_d ) capacitor c=0.00616547f \
 //x=16.28 //y=0 //x2=14.91 //y2=0.905
cc_126 ( N_GND_M8_noxref_d N_noxref_9_M9_noxref_d ) capacitor c=0.00143464f \
 //x=13.94 //y=0.865 //x2=14.91 //y2=0.905
cc_127 ( N_GND_c_8_p N_noxref_10_c_2170_n ) capacitor c=0.0148039f //x=23.68 \
 //y=0 //x2=23.565 //y2=3.33
cc_128 ( N_GND_c_1_p N_noxref_10_c_2170_n ) capacitor c=8.39131e-19 //x=23.68 \
 //y=0 //x2=23.565 //y2=3.33
cc_129 ( N_GND_c_6_p N_noxref_10_c_2172_n ) capacitor c=7.1088e-19 //x=16.28 \
 //y=0 //x2=18.13 //y2=2.08
cc_130 ( N_GND_c_7_p N_noxref_10_c_2172_n ) capacitor c=7.76678e-19 //x=19.61 \
 //y=0 //x2=18.13 //y2=2.08
cc_131 ( N_GND_c_1_p N_noxref_10_c_2174_n ) capacitor c=0.0461865f //x=23.68 \
 //y=0 //x2=23.595 //y2=1.665
cc_132 ( N_GND_c_1_p N_noxref_10_M14_noxref_d ) capacitor c=0.00593061f \
 //x=23.68 //y=0 //x2=23.005 //y2=0.915
cc_133 ( N_GND_c_2_p N_D_c_2340_n ) capacitor c=0.0177675f //x=0.74 //y=0 \
 //x2=1.11 //y2=2.08
cc_134 ( N_GND_c_134_p N_D_c_2341_n ) capacitor c=0.00135046f //x=1.095 //y=0 \
 //x2=0.915 //y2=0.865
cc_135 ( N_GND_M0_noxref_d N_D_c_2341_n ) capacitor c=0.00220047f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=0.865
cc_136 ( N_GND_M0_noxref_d N_D_c_2343_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=1.21
cc_137 ( N_GND_c_2_p N_D_c_2344_n ) capacitor c=0.00264481f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.52
cc_138 ( N_GND_c_2_p N_D_c_2345_n ) capacitor c=0.0121947f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.915
cc_139 ( N_GND_M0_noxref_d N_D_c_2346_n ) capacitor c=0.0131326f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=0.71
cc_140 ( N_GND_M0_noxref_d N_D_c_2347_n ) capacitor c=0.00193127f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=1.365
cc_141 ( N_GND_c_9_p N_D_c_2348_n ) capacitor c=0.00130622f //x=3.16 //y=0 \
 //x2=1.445 //y2=0.865
cc_142 ( N_GND_M0_noxref_d N_D_c_2348_n ) capacitor c=0.00257848f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=0.865
cc_143 ( N_GND_M0_noxref_d N_D_c_2350_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=1.21
cc_144 ( N_GND_c_8_p N_noxref_12_c_2397_n ) capacitor c=0.00710948f //x=23.68 \
 //y=0 //x2=1.58 //y2=1.58
cc_145 ( N_GND_c_134_p N_noxref_12_c_2397_n ) capacitor c=0.00111428f \
 //x=1.095 //y=0 //x2=1.58 //y2=1.58
cc_146 ( N_GND_c_9_p N_noxref_12_c_2397_n ) capacitor c=0.00180846f //x=3.16 \
 //y=0 //x2=1.58 //y2=1.58
cc_147 ( N_GND_M0_noxref_d N_noxref_12_c_2397_n ) capacitor c=0.0090983f \
 //x=0.99 //y=0.865 //x2=1.58 //y2=1.58
cc_148 ( N_GND_c_8_p N_noxref_12_c_2401_n ) capacitor c=0.00686741f //x=23.68 \
 //y=0 //x2=1.665 //y2=0.615
cc_149 ( N_GND_c_9_p N_noxref_12_c_2401_n ) capacitor c=0.0146208f //x=3.16 \
 //y=0 //x2=1.665 //y2=0.615
cc_150 ( N_GND_M0_noxref_d N_noxref_12_c_2401_n ) capacitor c=0.033812f \
 //x=0.99 //y=0.865 //x2=1.665 //y2=0.615
cc_151 ( N_GND_c_2_p N_noxref_12_c_2404_n ) capacitor c=2.91423e-19 //x=0.74 \
 //y=0 //x2=1.665 //y2=1.495
cc_152 ( N_GND_c_8_p N_noxref_12_c_2405_n ) capacitor c=0.0134195f //x=23.68 \
 //y=0 //x2=2.55 //y2=0.53
cc_153 ( N_GND_c_9_p N_noxref_12_c_2405_n ) capacitor c=0.0372723f //x=3.16 \
 //y=0 //x2=2.55 //y2=0.53
cc_154 ( N_GND_c_1_p N_noxref_12_c_2405_n ) capacitor c=0.00198522f //x=23.68 \
 //y=0 //x2=2.55 //y2=0.53
cc_155 ( N_GND_c_8_p N_noxref_12_c_2408_n ) capacitor c=0.0027057f //x=23.68 \
 //y=0 //x2=2.635 //y2=0.615
cc_156 ( N_GND_c_9_p N_noxref_12_c_2408_n ) capacitor c=0.0147125f //x=3.16 \
 //y=0 //x2=2.635 //y2=0.615
cc_157 ( N_GND_c_3_p N_noxref_12_c_2408_n ) capacitor c=0.0431718f //x=3.33 \
 //y=0 //x2=2.635 //y2=0.615
cc_158 ( N_GND_c_8_p N_noxref_12_M0_noxref_s ) capacitor c=0.00723598f \
 //x=23.68 //y=0 //x2=0.56 //y2=0.365
cc_159 ( N_GND_c_134_p N_noxref_12_M0_noxref_s ) capacitor c=0.0146208f \
 //x=1.095 //y=0 //x2=0.56 //y2=0.365
cc_160 ( N_GND_c_2_p N_noxref_12_M0_noxref_s ) capacitor c=0.0594057f //x=0.74 \
 //y=0 //x2=0.56 //y2=0.365
cc_161 ( N_GND_c_3_p N_noxref_12_M0_noxref_s ) capacitor c=0.00198098f \
 //x=3.33 //y=0 //x2=0.56 //y2=0.365
cc_162 ( N_GND_M0_noxref_d N_noxref_12_M0_noxref_s ) capacitor c=0.0334197f \
 //x=0.99 //y=0.865 //x2=0.56 //y2=0.365
cc_163 ( N_GND_c_8_p N_noxref_13_c_2445_n ) capacitor c=0.00529429f //x=23.68 \
 //y=0 //x2=4.805 //y2=1.59
cc_164 ( N_GND_c_10_p N_noxref_13_c_2445_n ) capacitor c=0.00111496f //x=4.32 \
 //y=0 //x2=4.805 //y2=1.59
cc_165 ( N_GND_c_15_p N_noxref_13_c_2445_n ) capacitor c=0.0018066f //x=7.97 \
 //y=0 //x2=4.805 //y2=1.59
cc_166 ( N_GND_M2_noxref_d N_noxref_13_c_2445_n ) capacitor c=0.00868399f \
 //x=4.215 //y=0.875 //x2=4.805 //y2=1.59
cc_167 ( N_GND_c_8_p N_noxref_13_c_2449_n ) capacitor c=0.00266608f //x=23.68 \
 //y=0 //x2=4.89 //y2=0.625
cc_168 ( N_GND_c_15_p N_noxref_13_c_2449_n ) capacitor c=0.0141814f //x=7.97 \
 //y=0 //x2=4.89 //y2=0.625
cc_169 ( N_GND_M2_noxref_d N_noxref_13_c_2449_n ) capacitor c=0.033954f \
 //x=4.215 //y=0.875 //x2=4.89 //y2=0.625
cc_170 ( N_GND_c_8_p N_noxref_13_c_2452_n ) capacitor c=0.0109327f //x=23.68 \
 //y=0 //x2=5.775 //y2=0.54
cc_171 ( N_GND_c_15_p N_noxref_13_c_2452_n ) capacitor c=0.0361235f //x=7.97 \
 //y=0 //x2=5.775 //y2=0.54
cc_172 ( N_GND_c_1_p N_noxref_13_c_2452_n ) capacitor c=0.00177401f //x=23.68 \
 //y=0 //x2=5.775 //y2=0.54
cc_173 ( N_GND_c_8_p N_noxref_13_M2_noxref_s ) capacitor c=0.00532331f \
 //x=23.68 //y=0 //x2=3.785 //y2=0.375
cc_174 ( N_GND_c_10_p N_noxref_13_M2_noxref_s ) capacitor c=0.0141814f \
 //x=4.32 //y=0 //x2=3.785 //y2=0.375
cc_175 ( N_GND_c_15_p N_noxref_13_M2_noxref_s ) capacitor c=0.0132355f \
 //x=7.97 //y=0 //x2=3.785 //y2=0.375
cc_176 ( N_GND_c_3_p N_noxref_13_M2_noxref_s ) capacitor c=0.0696963f //x=3.33 \
 //y=0 //x2=3.785 //y2=0.375
cc_177 ( N_GND_c_4_p N_noxref_13_M2_noxref_s ) capacitor c=3.31601e-19 \
 //x=8.14 //y=0 //x2=3.785 //y2=0.375
cc_178 ( N_GND_M2_noxref_d N_noxref_13_M2_noxref_s ) capacitor c=0.033718f \
 //x=4.215 //y=0.875 //x2=3.785 //y2=0.375
cc_179 ( N_GND_c_8_p N_noxref_14_c_2497_n ) capacitor c=0.00364762f //x=23.68 \
 //y=0 //x2=6.345 //y2=0.995
cc_180 ( N_GND_c_15_p N_noxref_14_c_2497_n ) capacitor c=0.00940048f //x=7.97 \
 //y=0 //x2=6.345 //y2=0.995
cc_181 ( N_GND_c_8_p N_noxref_14_c_2499_n ) capacitor c=0.00266608f //x=23.68 \
 //y=0 //x2=6.43 //y2=0.625
cc_182 ( N_GND_c_15_p N_noxref_14_c_2499_n ) capacitor c=0.0141814f //x=7.97 \
 //y=0 //x2=6.43 //y2=0.625
cc_183 ( N_GND_M2_noxref_d N_noxref_14_c_2499_n ) capacitor c=6.21394e-19 \
 //x=4.215 //y=0.875 //x2=6.43 //y2=0.625
cc_184 ( N_GND_c_8_p N_noxref_14_c_2502_n ) capacitor c=0.0110095f //x=23.68 \
 //y=0 //x2=7.315 //y2=0.54
cc_185 ( N_GND_c_15_p N_noxref_14_c_2502_n ) capacitor c=0.0365163f //x=7.97 \
 //y=0 //x2=7.315 //y2=0.54
cc_186 ( N_GND_c_1_p N_noxref_14_c_2502_n ) capacitor c=0.00189501f //x=23.68 \
 //y=0 //x2=7.315 //y2=0.54
cc_187 ( N_GND_c_8_p N_noxref_14_c_2505_n ) capacitor c=0.00266421f //x=23.68 \
 //y=0 //x2=7.4 //y2=0.625
cc_188 ( N_GND_c_15_p N_noxref_14_c_2505_n ) capacitor c=0.0141195f //x=7.97 \
 //y=0 //x2=7.4 //y2=0.625
cc_189 ( N_GND_c_4_p N_noxref_14_c_2505_n ) capacitor c=0.0404137f //x=8.14 \
 //y=0 //x2=7.4 //y2=0.625
cc_190 ( N_GND_M2_noxref_d N_noxref_14_M3_noxref_d ) capacitor c=0.00162435f \
 //x=4.215 //y=0.875 //x2=5.19 //y2=0.91
cc_191 ( N_GND_c_3_p N_noxref_14_M4_noxref_s ) capacitor c=8.16352e-19 \
 //x=3.33 //y=0 //x2=6.295 //y2=0.375
cc_192 ( N_GND_c_4_p N_noxref_14_M4_noxref_s ) capacitor c=0.00180469f \
 //x=8.14 //y=0 //x2=6.295 //y2=0.375
cc_193 ( N_GND_c_8_p N_noxref_15_c_2550_n ) capacitor c=0.00537035f //x=23.68 \
 //y=0 //x2=9.615 //y2=1.59
cc_194 ( N_GND_c_16_p N_noxref_15_c_2550_n ) capacitor c=0.00111496f //x=9.13 \
 //y=0 //x2=9.615 //y2=1.59
cc_195 ( N_GND_c_42_p N_noxref_15_c_2550_n ) capacitor c=0.00179185f //x=12.78 \
 //y=0 //x2=9.615 //y2=1.59
cc_196 ( N_GND_M5_noxref_d N_noxref_15_c_2550_n ) capacitor c=0.00868586f \
 //x=9.025 //y=0.875 //x2=9.615 //y2=1.59
cc_197 ( N_GND_c_8_p N_noxref_15_c_2554_n ) capacitor c=0.00296961f //x=23.68 \
 //y=0 //x2=9.7 //y2=0.625
cc_198 ( N_GND_c_42_p N_noxref_15_c_2554_n ) capacitor c=0.0140218f //x=12.78 \
 //y=0 //x2=9.7 //y2=0.625
cc_199 ( N_GND_M5_noxref_d N_noxref_15_c_2554_n ) capacitor c=0.033954f \
 //x=9.025 //y=0.875 //x2=9.7 //y2=0.625
cc_200 ( N_GND_c_8_p N_noxref_15_c_2557_n ) capacitor c=0.0113461f //x=23.68 \
 //y=0 //x2=10.585 //y2=0.54
cc_201 ( N_GND_c_42_p N_noxref_15_c_2557_n ) capacitor c=0.0358309f //x=12.78 \
 //y=0 //x2=10.585 //y2=0.54
cc_202 ( N_GND_c_1_p N_noxref_15_c_2557_n ) capacitor c=0.00177401f //x=23.68 \
 //y=0 //x2=10.585 //y2=0.54
cc_203 ( N_GND_c_8_p N_noxref_15_M5_noxref_s ) capacitor c=0.00519789f \
 //x=23.68 //y=0 //x2=8.595 //y2=0.375
cc_204 ( N_GND_c_16_p N_noxref_15_M5_noxref_s ) capacitor c=0.0141814f \
 //x=9.13 //y=0 //x2=8.595 //y2=0.375
cc_205 ( N_GND_c_42_p N_noxref_15_M5_noxref_s ) capacitor c=0.0131437f \
 //x=12.78 //y=0 //x2=8.595 //y2=0.375
cc_206 ( N_GND_c_4_p N_noxref_15_M5_noxref_s ) capacitor c=0.0696963f //x=8.14 \
 //y=0 //x2=8.595 //y2=0.375
cc_207 ( N_GND_c_5_p N_noxref_15_M5_noxref_s ) capacitor c=3.31601e-19 \
 //x=12.95 //y=0 //x2=8.595 //y2=0.375
cc_208 ( N_GND_M5_noxref_d N_noxref_15_M5_noxref_s ) capacitor c=0.033718f \
 //x=9.025 //y=0.875 //x2=8.595 //y2=0.375
cc_209 ( N_GND_c_8_p N_noxref_16_c_2604_n ) capacitor c=0.00352952f //x=23.68 \
 //y=0 //x2=11.155 //y2=0.995
cc_210 ( N_GND_c_42_p N_noxref_16_c_2604_n ) capacitor c=0.00934524f //x=12.78 \
 //y=0 //x2=11.155 //y2=0.995
cc_211 ( N_GND_c_8_p N_noxref_16_c_2606_n ) capacitor c=0.00254475f //x=23.68 \
 //y=0 //x2=11.24 //y2=0.625
cc_212 ( N_GND_c_42_p N_noxref_16_c_2606_n ) capacitor c=0.0140928f //x=12.78 \
 //y=0 //x2=11.24 //y2=0.625
cc_213 ( N_GND_M5_noxref_d N_noxref_16_c_2606_n ) capacitor c=6.21394e-19 \
 //x=9.025 //y=0.875 //x2=11.24 //y2=0.625
cc_214 ( N_GND_c_8_p N_noxref_16_c_2609_n ) capacitor c=0.0105317f //x=23.68 \
 //y=0 //x2=12.125 //y2=0.54
cc_215 ( N_GND_c_42_p N_noxref_16_c_2609_n ) capacitor c=0.0364215f //x=12.78 \
 //y=0 //x2=12.125 //y2=0.54
cc_216 ( N_GND_c_1_p N_noxref_16_c_2609_n ) capacitor c=0.00189501f //x=23.68 \
 //y=0 //x2=12.125 //y2=0.54
cc_217 ( N_GND_c_8_p N_noxref_16_c_2612_n ) capacitor c=0.00254232f //x=23.68 \
 //y=0 //x2=12.21 //y2=0.625
cc_218 ( N_GND_c_42_p N_noxref_16_c_2612_n ) capacitor c=0.0140304f //x=12.78 \
 //y=0 //x2=12.21 //y2=0.625
cc_219 ( N_GND_c_5_p N_noxref_16_c_2612_n ) capacitor c=0.0404137f //x=12.95 \
 //y=0 //x2=12.21 //y2=0.625
cc_220 ( N_GND_M5_noxref_d N_noxref_16_M6_noxref_d ) capacitor c=0.00162435f \
 //x=9.025 //y=0.875 //x2=10 //y2=0.91
cc_221 ( N_GND_c_4_p N_noxref_16_M7_noxref_s ) capacitor c=8.16352e-19 \
 //x=8.14 //y=0 //x2=11.105 //y2=0.375
cc_222 ( N_GND_c_5_p N_noxref_16_M7_noxref_s ) capacitor c=0.00183576f \
 //x=12.95 //y=0 //x2=11.105 //y2=0.375
cc_223 ( N_GND_c_8_p N_noxref_17_c_2657_n ) capacitor c=0.00517234f //x=23.68 \
 //y=0 //x2=14.53 //y2=1.58
cc_224 ( N_GND_c_53_p N_noxref_17_c_2657_n ) capacitor c=0.00112872f \
 //x=14.045 //y=0 //x2=14.53 //y2=1.58
cc_225 ( N_GND_c_60_p N_noxref_17_c_2657_n ) capacitor c=0.0018229f //x=16.11 \
 //y=0 //x2=14.53 //y2=1.58
cc_226 ( N_GND_M8_noxref_d N_noxref_17_c_2657_n ) capacitor c=0.008625f \
 //x=13.94 //y=0.865 //x2=14.53 //y2=1.58
cc_227 ( N_GND_c_8_p N_noxref_17_c_2661_n ) capacitor c=0.00259029f //x=23.68 \
 //y=0 //x2=14.615 //y2=0.615
cc_228 ( N_GND_c_60_p N_noxref_17_c_2661_n ) capacitor c=0.0146901f //x=16.11 \
 //y=0 //x2=14.615 //y2=0.615
cc_229 ( N_GND_M8_noxref_d N_noxref_17_c_2661_n ) capacitor c=0.033812f \
 //x=13.94 //y=0.865 //x2=14.615 //y2=0.615
cc_230 ( N_GND_c_5_p N_noxref_17_c_2664_n ) capacitor c=2.91423e-19 //x=12.95 \
 //y=0 //x2=14.615 //y2=1.495
cc_231 ( N_GND_c_8_p N_noxref_17_c_2665_n ) capacitor c=0.0106919f //x=23.68 \
 //y=0 //x2=15.5 //y2=0.53
cc_232 ( N_GND_c_60_p N_noxref_17_c_2665_n ) capacitor c=0.0374253f //x=16.11 \
 //y=0 //x2=15.5 //y2=0.53
cc_233 ( N_GND_c_1_p N_noxref_17_c_2665_n ) capacitor c=0.00198522f //x=23.68 \
 //y=0 //x2=15.5 //y2=0.53
cc_234 ( N_GND_c_8_p N_noxref_17_c_2668_n ) capacitor c=0.00258845f //x=23.68 \
 //y=0 //x2=15.585 //y2=0.615
cc_235 ( N_GND_c_60_p N_noxref_17_c_2668_n ) capacitor c=0.0146256f //x=16.11 \
 //y=0 //x2=15.585 //y2=0.615
cc_236 ( N_GND_c_6_p N_noxref_17_c_2668_n ) capacitor c=0.0431718f //x=16.28 \
 //y=0 //x2=15.585 //y2=0.615
cc_237 ( N_GND_c_8_p N_noxref_17_M8_noxref_s ) capacitor c=0.00259029f \
 //x=23.68 //y=0 //x2=13.51 //y2=0.365
cc_238 ( N_GND_c_53_p N_noxref_17_M8_noxref_s ) capacitor c=0.0146901f \
 //x=14.045 //y=0 //x2=13.51 //y2=0.365
cc_239 ( N_GND_c_5_p N_noxref_17_M8_noxref_s ) capacitor c=0.0583534f \
 //x=12.95 //y=0 //x2=13.51 //y2=0.365
cc_240 ( N_GND_c_6_p N_noxref_17_M8_noxref_s ) capacitor c=0.00198043f \
 //x=16.28 //y=0 //x2=13.51 //y2=0.365
cc_241 ( N_GND_M8_noxref_d N_noxref_17_M8_noxref_s ) capacitor c=0.0334197f \
 //x=13.94 //y=0.865 //x2=13.51 //y2=0.365
cc_242 ( N_GND_c_8_p N_noxref_18_c_2709_n ) capacitor c=0.00517234f //x=23.68 \
 //y=0 //x2=17.86 //y2=1.58
cc_243 ( N_GND_c_74_p N_noxref_18_c_2709_n ) capacitor c=0.00112872f \
 //x=17.375 //y=0 //x2=17.86 //y2=1.58
cc_244 ( N_GND_c_81_p N_noxref_18_c_2709_n ) capacitor c=0.0018229f //x=19.44 \
 //y=0 //x2=17.86 //y2=1.58
cc_245 ( N_GND_M10_noxref_d N_noxref_18_c_2709_n ) capacitor c=0.008625f \
 //x=17.27 //y=0.865 //x2=17.86 //y2=1.58
cc_246 ( N_GND_c_8_p N_noxref_18_c_2713_n ) capacitor c=0.00259029f //x=23.68 \
 //y=0 //x2=17.945 //y2=0.615
cc_247 ( N_GND_c_81_p N_noxref_18_c_2713_n ) capacitor c=0.0143795f //x=19.44 \
 //y=0 //x2=17.945 //y2=0.615
cc_248 ( N_GND_M10_noxref_d N_noxref_18_c_2713_n ) capacitor c=0.033812f \
 //x=17.27 //y=0.865 //x2=17.945 //y2=0.615
cc_249 ( N_GND_c_6_p N_noxref_18_c_2716_n ) capacitor c=2.91423e-19 //x=16.28 \
 //y=0 //x2=17.945 //y2=1.495
cc_250 ( N_GND_c_8_p N_noxref_18_c_2717_n ) capacitor c=0.0106919f //x=23.68 \
 //y=0 //x2=18.83 //y2=0.53
cc_251 ( N_GND_c_81_p N_noxref_18_c_2717_n ) capacitor c=0.0374253f //x=19.44 \
 //y=0 //x2=18.83 //y2=0.53
cc_252 ( N_GND_c_1_p N_noxref_18_c_2717_n ) capacitor c=0.00198522f //x=23.68 \
 //y=0 //x2=18.83 //y2=0.53
cc_253 ( N_GND_c_8_p N_noxref_18_c_2720_n ) capacitor c=0.00258845f //x=23.68 \
 //y=0 //x2=18.915 //y2=0.615
cc_254 ( N_GND_c_81_p N_noxref_18_c_2720_n ) capacitor c=0.0146256f //x=19.44 \
 //y=0 //x2=18.915 //y2=0.615
cc_255 ( N_GND_c_7_p N_noxref_18_c_2720_n ) capacitor c=0.0431718f //x=19.61 \
 //y=0 //x2=18.915 //y2=0.615
cc_256 ( N_GND_c_8_p N_noxref_18_M10_noxref_s ) capacitor c=0.00259029f \
 //x=23.68 //y=0 //x2=16.84 //y2=0.365
cc_257 ( N_GND_c_74_p N_noxref_18_M10_noxref_s ) capacitor c=0.0146901f \
 //x=17.375 //y=0 //x2=16.84 //y2=0.365
cc_258 ( N_GND_c_6_p N_noxref_18_M10_noxref_s ) capacitor c=0.058339f \
 //x=16.28 //y=0 //x2=16.84 //y2=0.365
cc_259 ( N_GND_c_7_p N_noxref_18_M10_noxref_s ) capacitor c=0.00198098f \
 //x=19.61 //y=0 //x2=16.84 //y2=0.365
cc_260 ( N_GND_M10_noxref_d N_noxref_18_M10_noxref_s ) capacitor c=0.0334197f \
 //x=17.27 //y=0.865 //x2=16.84 //y2=0.365
cc_261 ( N_GND_c_8_p N_noxref_19_c_2761_n ) capacitor c=0.00517576f //x=23.68 \
 //y=0 //x2=21.085 //y2=1.59
cc_262 ( N_GND_c_89_p N_noxref_19_c_2761_n ) capacitor c=0.00111448f //x=20.6 \
 //y=0 //x2=21.085 //y2=1.59
cc_263 ( N_GND_c_1_p N_noxref_19_c_2761_n ) capacitor c=0.00180612f //x=23.68 \
 //y=0 //x2=21.085 //y2=1.59
cc_264 ( N_GND_M12_noxref_d N_noxref_19_c_2761_n ) capacitor c=0.00853078f \
 //x=20.495 //y=0.875 //x2=21.085 //y2=1.59
cc_265 ( N_GND_c_8_p N_noxref_19_c_2765_n ) capacitor c=0.00254475f //x=23.68 \
 //y=0 //x2=21.17 //y2=0.625
cc_266 ( N_GND_c_1_p N_noxref_19_c_2765_n ) capacitor c=0.0140928f //x=23.68 \
 //y=0 //x2=21.17 //y2=0.625
cc_267 ( N_GND_M12_noxref_d N_noxref_19_c_2765_n ) capacitor c=0.033954f \
 //x=20.495 //y=0.875 //x2=21.17 //y2=0.625
cc_268 ( N_GND_c_8_p N_noxref_19_c_2768_n ) capacitor c=0.0105704f //x=23.68 \
 //y=0 //x2=22.055 //y2=0.54
cc_269 ( N_GND_c_1_p N_noxref_19_c_2768_n ) capacitor c=0.0379112f //x=23.68 \
 //y=0 //x2=22.055 //y2=0.54
cc_270 ( N_GND_c_8_p N_noxref_19_M12_noxref_s ) capacitor c=0.00541939f \
 //x=23.68 //y=0 //x2=20.065 //y2=0.375
cc_271 ( N_GND_c_89_p N_noxref_19_M12_noxref_s ) capacitor c=0.0140928f \
 //x=20.6 //y=0 //x2=20.065 //y2=0.375
cc_272 ( N_GND_c_1_p N_noxref_19_M12_noxref_s ) capacitor c=0.013718f \
 //x=23.68 //y=0 //x2=20.065 //y2=0.375
cc_273 ( N_GND_c_7_p N_noxref_19_M12_noxref_s ) capacitor c=0.0696963f \
 //x=19.61 //y=0 //x2=20.065 //y2=0.375
cc_274 ( N_GND_M12_noxref_d N_noxref_19_M12_noxref_s ) capacitor c=0.033718f \
 //x=20.495 //y=0.875 //x2=20.065 //y2=0.375
cc_275 ( N_GND_c_8_p N_noxref_20_c_2811_n ) capacitor c=0.00385233f //x=23.68 \
 //y=0 //x2=22.625 //y2=0.995
cc_276 ( N_GND_c_1_p N_noxref_20_c_2811_n ) capacitor c=0.0096703f //x=23.68 \
 //y=0 //x2=22.625 //y2=0.995
cc_277 ( N_GND_c_8_p N_noxref_20_c_2813_n ) capacitor c=0.00287639f //x=23.68 \
 //y=0 //x2=22.71 //y2=0.625
cc_278 ( N_GND_c_1_p N_noxref_20_c_2813_n ) capacitor c=0.014327f //x=23.68 \
 //y=0 //x2=22.71 //y2=0.625
cc_279 ( N_GND_M12_noxref_d N_noxref_20_c_2813_n ) capacitor c=6.21394e-19 \
 //x=20.495 //y=0.875 //x2=22.71 //y2=0.625
cc_280 ( N_GND_c_8_p N_noxref_20_c_2816_n ) capacitor c=0.0118444f //x=23.68 \
 //y=0 //x2=23.595 //y2=0.54
cc_281 ( N_GND_c_1_p N_noxref_20_c_2816_n ) capacitor c=0.0384431f //x=23.68 \
 //y=0 //x2=23.595 //y2=0.54
cc_282 ( N_GND_c_8_p N_noxref_20_c_2818_n ) capacitor c=0.00286759f //x=23.68 \
 //y=0 //x2=23.68 //y2=0.625
cc_283 ( N_GND_c_1_p N_noxref_20_c_2818_n ) capacitor c=0.0553579f //x=23.68 \
 //y=0 //x2=23.68 //y2=0.625
cc_284 ( N_GND_M12_noxref_d N_noxref_20_M13_noxref_d ) capacitor c=0.00162435f \
 //x=20.495 //y=0.875 //x2=21.47 //y2=0.91
cc_285 ( N_GND_c_1_p N_noxref_20_M14_noxref_s ) capacitor c=0.00183576f \
 //x=23.68 //y=0 //x2=22.575 //y2=0.375
cc_286 ( N_GND_c_7_p N_noxref_20_M14_noxref_s ) capacitor c=8.16352e-19 \
 //x=19.61 //y=0 //x2=22.575 //y2=0.375
cc_287 ( N_VDD_c_289_n N_noxref_3_c_591_n ) capacitor c=0.00137387f //x=3.33 \
 //y=7.4 //x2=4.295 //y2=2.59
cc_288 ( N_VDD_c_295_p N_noxref_3_c_632_n ) capacitor c=0.00546694f //x=23.68 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_289 ( N_VDD_c_296_p N_noxref_3_c_632_n ) capacitor c=4.3394e-19 //x=1.585 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_290 ( N_VDD_c_297_p N_noxref_3_c_632_n ) capacitor c=4.48693e-19 //x=2.465 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_291 ( N_VDD_M16_noxref_d N_noxref_3_c_632_n ) capacitor c=0.0129678f \
 //x=1.525 //y=5.02 //x2=2.025 //y2=5.2
cc_292 ( N_VDD_c_288_n N_noxref_3_c_636_n ) capacitor c=0.00989999f //x=0.74 \
 //y=7.4 //x2=1.315 //y2=5.2
cc_293 ( N_VDD_M15_noxref_s N_noxref_3_c_636_n ) capacitor c=0.087833f \
 //x=0.655 //y=5.02 //x2=1.315 //y2=5.2
cc_294 ( N_VDD_c_295_p N_noxref_3_c_638_n ) capacitor c=0.00307195f //x=23.68 \
 //y=7.4 //x2=2.505 //y2=5.2
cc_295 ( N_VDD_c_297_p N_noxref_3_c_638_n ) capacitor c=7.73167e-19 //x=2.465 \
 //y=7.4 //x2=2.505 //y2=5.2
cc_296 ( N_VDD_M18_noxref_d N_noxref_3_c_638_n ) capacitor c=0.0161518f \
 //x=2.405 //y=5.02 //x2=2.505 //y2=5.2
cc_297 ( N_VDD_c_288_n N_noxref_3_c_604_n ) capacitor c=0.00159771f //x=0.74 \
 //y=7.4 //x2=2.59 //y2=2.59
cc_298 ( N_VDD_c_289_n N_noxref_3_c_604_n ) capacitor c=0.0452382f //x=3.33 \
 //y=7.4 //x2=2.59 //y2=2.59
cc_299 ( N_VDD_c_295_p N_noxref_3_c_606_n ) capacitor c=9.23542e-19 //x=23.68 \
 //y=7.4 //x2=4.44 //y2=2.08
cc_300 ( N_VDD_c_289_n N_noxref_3_c_606_n ) capacitor c=0.0157357f //x=3.33 \
 //y=7.4 //x2=4.44 //y2=2.08
cc_301 ( N_VDD_M19_noxref_s N_noxref_3_c_606_n ) capacitor c=0.0129925f \
 //x=4.285 //y=5.02 //x2=4.44 //y2=2.08
cc_302 ( N_VDD_c_295_p N_noxref_3_c_607_n ) capacitor c=9.10347e-19 //x=23.68 \
 //y=7.4 //x2=9.25 //y2=2.08
cc_303 ( N_VDD_c_290_n N_noxref_3_c_607_n ) capacitor c=0.013427f //x=8.14 \
 //y=7.4 //x2=9.25 //y2=2.08
cc_304 ( N_VDD_M25_noxref_s N_noxref_3_c_607_n ) capacitor c=0.0120327f \
 //x=9.095 //y=5.02 //x2=9.25 //y2=2.08
cc_305 ( N_VDD_c_312_p N_noxref_3_M19_noxref_g ) capacitor c=0.00749687f \
 //x=5.215 //y=7.4 //x2=4.64 //y2=6.02
cc_306 ( N_VDD_M19_noxref_s N_noxref_3_M19_noxref_g ) capacitor c=0.0477201f \
 //x=4.285 //y=5.02 //x2=4.64 //y2=6.02
cc_307 ( N_VDD_c_312_p N_noxref_3_M20_noxref_g ) capacitor c=0.00675175f \
 //x=5.215 //y=7.4 //x2=5.08 //y2=6.02
cc_308 ( N_VDD_M20_noxref_d N_noxref_3_M20_noxref_g ) capacitor c=0.015318f \
 //x=5.155 //y=5.02 //x2=5.08 //y2=6.02
cc_309 ( N_VDD_c_316_p N_noxref_3_M25_noxref_g ) capacitor c=0.00749687f \
 //x=10.025 //y=7.4 //x2=9.45 //y2=6.02
cc_310 ( N_VDD_M25_noxref_s N_noxref_3_M25_noxref_g ) capacitor c=0.0477201f \
 //x=9.095 //y=5.02 //x2=9.45 //y2=6.02
cc_311 ( N_VDD_c_316_p N_noxref_3_M26_noxref_g ) capacitor c=0.00675175f \
 //x=10.025 //y=7.4 //x2=9.89 //y2=6.02
cc_312 ( N_VDD_M26_noxref_d N_noxref_3_M26_noxref_g ) capacitor c=0.015318f \
 //x=9.965 //y=5.02 //x2=9.89 //y2=6.02
cc_313 ( N_VDD_c_289_n N_noxref_3_c_657_n ) capacitor c=0.00757682f //x=3.33 \
 //y=7.4 //x2=4.715 //y2=4.79
cc_314 ( N_VDD_M19_noxref_s N_noxref_3_c_657_n ) capacitor c=0.00445134f \
 //x=4.285 //y=5.02 //x2=4.715 //y2=4.79
cc_315 ( N_VDD_c_290_n N_noxref_3_c_659_n ) capacitor c=0.00757682f //x=8.14 \
 //y=7.4 //x2=9.525 //y2=4.79
cc_316 ( N_VDD_M25_noxref_s N_noxref_3_c_659_n ) capacitor c=0.00444914f \
 //x=9.095 //y=5.02 //x2=9.525 //y2=4.79
cc_317 ( N_VDD_c_295_p N_noxref_3_M15_noxref_d ) capacitor c=0.00706239f \
 //x=23.68 //y=7.4 //x2=1.085 //y2=5.02
cc_318 ( N_VDD_c_296_p N_noxref_3_M15_noxref_d ) capacitor c=0.0138103f \
 //x=1.585 //y=7.4 //x2=1.085 //y2=5.02
cc_319 ( N_VDD_c_289_n N_noxref_3_M15_noxref_d ) capacitor c=6.94454e-19 \
 //x=3.33 //y=7.4 //x2=1.085 //y2=5.02
cc_320 ( N_VDD_M16_noxref_d N_noxref_3_M15_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.085 //y2=5.02
cc_321 ( N_VDD_c_295_p N_noxref_3_M17_noxref_d ) capacitor c=0.00285083f \
 //x=23.68 //y=7.4 //x2=1.965 //y2=5.02
cc_322 ( N_VDD_c_297_p N_noxref_3_M17_noxref_d ) capacitor c=0.0140984f \
 //x=2.465 //y=7.4 //x2=1.965 //y2=5.02
cc_323 ( N_VDD_c_289_n N_noxref_3_M17_noxref_d ) capacitor c=0.0120541f \
 //x=3.33 //y=7.4 //x2=1.965 //y2=5.02
cc_324 ( N_VDD_M15_noxref_s N_noxref_3_M17_noxref_d ) capacitor c=0.00111971f \
 //x=0.655 //y=5.02 //x2=1.965 //y2=5.02
cc_325 ( N_VDD_M16_noxref_d N_noxref_3_M17_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.965 //y2=5.02
cc_326 ( N_VDD_M18_noxref_d N_noxref_3_M17_noxref_d ) capacitor c=0.0664752f \
 //x=2.405 //y=5.02 //x2=1.965 //y2=5.02
cc_327 ( N_VDD_M19_noxref_s N_noxref_3_M17_noxref_d ) capacitor c=3.73257e-19 \
 //x=4.285 //y=5.02 //x2=1.965 //y2=5.02
cc_328 ( N_VDD_c_295_p N_noxref_4_c_847_n ) capacitor c=0.00444892f //x=23.68 \
 //y=7.4 //x2=10.465 //y2=5.155
cc_329 ( N_VDD_c_316_p N_noxref_4_c_847_n ) capacitor c=4.31931e-19 //x=10.025 \
 //y=7.4 //x2=10.465 //y2=5.155
cc_330 ( N_VDD_c_337_p N_noxref_4_c_847_n ) capacitor c=4.31931e-19 //x=10.905 \
 //y=7.4 //x2=10.465 //y2=5.155
cc_331 ( N_VDD_M26_noxref_d N_noxref_4_c_847_n ) capacitor c=0.0112985f \
 //x=9.965 //y=5.02 //x2=10.465 //y2=5.155
cc_332 ( N_VDD_c_290_n N_noxref_4_c_851_n ) capacitor c=0.00863585f //x=8.14 \
 //y=7.4 //x2=9.755 //y2=5.155
cc_333 ( N_VDD_M25_noxref_s N_noxref_4_c_851_n ) capacitor c=0.0831083f \
 //x=9.095 //y=5.02 //x2=9.755 //y2=5.155
cc_334 ( N_VDD_c_295_p N_noxref_4_c_853_n ) capacitor c=0.0044221f //x=23.68 \
 //y=7.4 //x2=11.345 //y2=5.155
cc_335 ( N_VDD_c_337_p N_noxref_4_c_853_n ) capacitor c=4.31931e-19 //x=10.905 \
 //y=7.4 //x2=11.345 //y2=5.155
cc_336 ( N_VDD_c_343_p N_noxref_4_c_853_n ) capacitor c=4.31931e-19 //x=11.785 \
 //y=7.4 //x2=11.345 //y2=5.155
cc_337 ( N_VDD_M28_noxref_d N_noxref_4_c_853_n ) capacitor c=0.0112985f \
 //x=10.845 //y=5.02 //x2=11.345 //y2=5.155
cc_338 ( N_VDD_c_295_p N_noxref_4_c_857_n ) capacitor c=0.00434174f //x=23.68 \
 //y=7.4 //x2=12.125 //y2=5.155
cc_339 ( N_VDD_c_343_p N_noxref_4_c_857_n ) capacitor c=7.46626e-19 //x=11.785 \
 //y=7.4 //x2=12.125 //y2=5.155
cc_340 ( N_VDD_c_347_p N_noxref_4_c_857_n ) capacitor c=0.00198565f //x=12.78 \
 //y=7.4 //x2=12.125 //y2=5.155
cc_341 ( N_VDD_M30_noxref_d N_noxref_4_c_857_n ) capacitor c=0.0112985f \
 //x=11.725 //y=5.02 //x2=12.125 //y2=5.155
cc_342 ( N_VDD_c_291_n N_noxref_4_c_834_n ) capacitor c=0.042636f //x=12.95 \
 //y=7.4 //x2=12.21 //y2=2.59
cc_343 ( N_VDD_c_295_p N_noxref_4_c_835_n ) capacitor c=0.00125279f //x=23.68 \
 //y=7.4 //x2=14.06 //y2=2.08
cc_344 ( N_VDD_c_351_p N_noxref_4_c_835_n ) capacitor c=2.87256e-19 //x=14.535 \
 //y=7.4 //x2=14.06 //y2=2.08
cc_345 ( N_VDD_c_291_n N_noxref_4_c_835_n ) capacitor c=0.0133961f //x=12.95 \
 //y=7.4 //x2=14.06 //y2=2.08
cc_346 ( N_VDD_c_351_p N_noxref_4_M31_noxref_g ) capacitor c=0.00726866f \
 //x=14.535 //y=7.4 //x2=13.96 //y2=6.02
cc_347 ( N_VDD_M31_noxref_s N_noxref_4_M31_noxref_g ) capacitor c=0.054195f \
 //x=13.605 //y=5.02 //x2=13.96 //y2=6.02
cc_348 ( N_VDD_c_351_p N_noxref_4_M32_noxref_g ) capacitor c=0.00672952f \
 //x=14.535 //y=7.4 //x2=14.4 //y2=6.02
cc_349 ( N_VDD_M32_noxref_d N_noxref_4_M32_noxref_g ) capacitor c=0.015318f \
 //x=14.475 //y=5.02 //x2=14.4 //y2=6.02
cc_350 ( N_VDD_c_291_n N_noxref_4_c_869_n ) capacitor c=0.015293f //x=12.95 \
 //y=7.4 //x2=14.06 //y2=4.7
cc_351 ( N_VDD_c_295_p N_noxref_4_M25_noxref_d ) capacitor c=0.00275235f \
 //x=23.68 //y=7.4 //x2=9.525 //y2=5.02
cc_352 ( N_VDD_c_316_p N_noxref_4_M25_noxref_d ) capacitor c=0.014035f \
 //x=10.025 //y=7.4 //x2=9.525 //y2=5.02
cc_353 ( N_VDD_M26_noxref_d N_noxref_4_M25_noxref_d ) capacitor c=0.0664752f \
 //x=9.965 //y=5.02 //x2=9.525 //y2=5.02
cc_354 ( N_VDD_c_295_p N_noxref_4_M27_noxref_d ) capacitor c=0.00275235f \
 //x=23.68 //y=7.4 //x2=10.405 //y2=5.02
cc_355 ( N_VDD_c_337_p N_noxref_4_M27_noxref_d ) capacitor c=0.014035f \
 //x=10.905 //y=7.4 //x2=10.405 //y2=5.02
cc_356 ( N_VDD_c_291_n N_noxref_4_M27_noxref_d ) capacitor c=4.9285e-19 \
 //x=12.95 //y=7.4 //x2=10.405 //y2=5.02
cc_357 ( N_VDD_M25_noxref_s N_noxref_4_M27_noxref_d ) capacitor c=0.00130656f \
 //x=9.095 //y=5.02 //x2=10.405 //y2=5.02
cc_358 ( N_VDD_M26_noxref_d N_noxref_4_M27_noxref_d ) capacitor c=0.0664752f \
 //x=9.965 //y=5.02 //x2=10.405 //y2=5.02
cc_359 ( N_VDD_M28_noxref_d N_noxref_4_M27_noxref_d ) capacitor c=0.0664752f \
 //x=10.845 //y=5.02 //x2=10.405 //y2=5.02
cc_360 ( N_VDD_c_295_p N_noxref_4_M29_noxref_d ) capacitor c=0.00275235f \
 //x=23.68 //y=7.4 //x2=11.285 //y2=5.02
cc_361 ( N_VDD_c_343_p N_noxref_4_M29_noxref_d ) capacitor c=0.014035f \
 //x=11.785 //y=7.4 //x2=11.285 //y2=5.02
cc_362 ( N_VDD_c_291_n N_noxref_4_M29_noxref_d ) capacitor c=0.00939849f \
 //x=12.95 //y=7.4 //x2=11.285 //y2=5.02
cc_363 ( N_VDD_M28_noxref_d N_noxref_4_M29_noxref_d ) capacitor c=0.0664752f \
 //x=10.845 //y=5.02 //x2=11.285 //y2=5.02
cc_364 ( N_VDD_M30_noxref_d N_noxref_4_M29_noxref_d ) capacitor c=0.0664752f \
 //x=11.725 //y=5.02 //x2=11.285 //y2=5.02
cc_365 ( N_VDD_M31_noxref_s N_noxref_4_M29_noxref_d ) capacitor c=4.52683e-19 \
 //x=13.605 //y=5.02 //x2=11.285 //y2=5.02
cc_366 ( N_VDD_c_295_p N_CLK_c_994_n ) capacitor c=0.0693925f //x=23.68 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_367 ( N_VDD_c_374_p N_CLK_c_994_n ) capacitor c=0.00258496f //x=7.97 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_368 ( N_VDD_c_375_p N_CLK_c_994_n ) capacitor c=0.00328994f //x=9.145 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_369 ( N_VDD_c_316_p N_CLK_c_994_n ) capacitor c=0.00135925f //x=10.025 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_370 ( N_VDD_c_347_p N_CLK_c_994_n ) capacitor c=0.00258496f //x=12.78 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_371 ( N_VDD_c_378_p N_CLK_c_994_n ) capacitor c=0.00209689f //x=13.655 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_372 ( N_VDD_c_351_p N_CLK_c_994_n ) capacitor c=7.81728e-19 //x=14.535 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_373 ( N_VDD_c_290_n N_CLK_c_994_n ) capacitor c=0.0389825f //x=8.14 //y=7.4 \
 //x2=14.685 //y2=4.44
cc_374 ( N_VDD_c_291_n N_CLK_c_994_n ) capacitor c=0.0389825f //x=12.95 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_375 ( N_VDD_M25_noxref_s N_CLK_c_994_n ) capacitor c=0.00179496f //x=9.095 \
 //y=5.02 //x2=14.685 //y2=4.44
cc_376 ( N_VDD_M31_noxref_s N_CLK_c_994_n ) capacitor c=0.00541054f //x=13.605 \
 //y=5.02 //x2=14.685 //y2=4.44
cc_377 ( N_VDD_c_295_p N_CLK_c_1005_n ) capacitor c=0.00146064f //x=23.68 \
 //y=7.4 //x2=5.665 //y2=4.44
cc_378 ( N_VDD_c_295_p N_CLK_c_991_n ) capacitor c=2.03287e-19 //x=23.68 \
 //y=7.4 //x2=5.55 //y2=2.08
cc_379 ( N_VDD_c_289_n N_CLK_c_991_n ) capacitor c=8.47879e-19 //x=3.33 \
 //y=7.4 //x2=5.55 //y2=2.08
cc_380 ( N_VDD_c_291_n N_CLK_c_992_n ) capacitor c=4.60777e-19 //x=12.95 \
 //y=7.4 //x2=14.8 //y2=2.08
cc_381 ( N_VDD_c_292_n N_CLK_c_992_n ) capacitor c=7.28243e-19 //x=16.28 \
 //y=7.4 //x2=14.8 //y2=2.08
cc_382 ( N_VDD_c_389_p N_CLK_M21_noxref_g ) capacitor c=0.00676195f //x=6.095 \
 //y=7.4 //x2=5.52 //y2=6.02
cc_383 ( N_VDD_M20_noxref_d N_CLK_M21_noxref_g ) capacitor c=0.015318f \
 //x=5.155 //y=5.02 //x2=5.52 //y2=6.02
cc_384 ( N_VDD_c_389_p N_CLK_M22_noxref_g ) capacitor c=0.00675175f //x=6.095 \
 //y=7.4 //x2=5.96 //y2=6.02
cc_385 ( N_VDD_M22_noxref_d N_CLK_M22_noxref_g ) capacitor c=0.015318f \
 //x=6.035 //y=5.02 //x2=5.96 //y2=6.02
cc_386 ( N_VDD_c_393_p N_CLK_M33_noxref_g ) capacitor c=0.00673971f //x=15.415 \
 //y=7.4 //x2=14.84 //y2=6.02
cc_387 ( N_VDD_M32_noxref_d N_CLK_M33_noxref_g ) capacitor c=0.015318f \
 //x=14.475 //y=5.02 //x2=14.84 //y2=6.02
cc_388 ( N_VDD_c_393_p N_CLK_M34_noxref_g ) capacitor c=0.00672952f //x=15.415 \
 //y=7.4 //x2=15.28 //y2=6.02
cc_389 ( N_VDD_c_292_n N_CLK_M34_noxref_g ) capacitor c=0.00864163f //x=16.28 \
 //y=7.4 //x2=15.28 //y2=6.02
cc_390 ( N_VDD_M34_noxref_d N_CLK_M34_noxref_g ) capacitor c=0.0430452f \
 //x=15.355 //y=5.02 //x2=15.28 //y2=6.02
cc_391 ( N_VDD_c_295_p N_noxref_6_c_1189_n ) capacitor c=0.031669f //x=23.68 \
 //y=7.4 //x2=7.28 //y2=4.07
cc_392 ( N_VDD_c_399_p N_noxref_6_c_1189_n ) capacitor c=0.00168692f //x=3.16 \
 //y=7.4 //x2=7.28 //y2=4.07
cc_393 ( N_VDD_c_400_p N_noxref_6_c_1189_n ) capacitor c=0.0027159f //x=4.335 \
 //y=7.4 //x2=7.28 //y2=4.07
cc_394 ( N_VDD_c_312_p N_noxref_6_c_1189_n ) capacitor c=0.00113459f //x=5.215 \
 //y=7.4 //x2=7.28 //y2=4.07
cc_395 ( N_VDD_c_289_n N_noxref_6_c_1189_n ) capacitor c=0.0276227f //x=3.33 \
 //y=7.4 //x2=7.28 //y2=4.07
cc_396 ( N_VDD_M18_noxref_d N_noxref_6_c_1189_n ) capacitor c=5.05307e-19 \
 //x=2.405 //y=5.02 //x2=7.28 //y2=4.07
cc_397 ( N_VDD_M19_noxref_s N_noxref_6_c_1189_n ) capacitor c=0.00122826f \
 //x=4.285 //y=5.02 //x2=7.28 //y2=4.07
cc_398 ( N_VDD_c_295_p N_noxref_6_c_1191_n ) capacitor c=0.00181362f //x=23.68 \
 //y=7.4 //x2=1.965 //y2=4.07
cc_399 ( N_VDD_c_295_p N_noxref_6_c_1215_n ) capacitor c=0.046539f //x=23.68 \
 //y=7.4 //x2=17.275 //y2=4.07
cc_400 ( N_VDD_c_407_p N_noxref_6_c_1215_n ) capacitor c=0.00168692f //x=16.11 \
 //y=7.4 //x2=17.275 //y2=4.07
cc_401 ( N_VDD_c_408_p N_noxref_6_c_1215_n ) capacitor c=0.00172186f \
 //x=16.985 //y=7.4 //x2=17.275 //y2=4.07
cc_402 ( N_VDD_c_409_p N_noxref_6_c_1215_n ) capacitor c=6.62004e-19 \
 //x=17.865 //y=7.4 //x2=17.275 //y2=4.07
cc_403 ( N_VDD_c_290_n N_noxref_6_c_1215_n ) capacitor c=0.0140578f //x=8.14 \
 //y=7.4 //x2=17.275 //y2=4.07
cc_404 ( N_VDD_c_291_n N_noxref_6_c_1215_n ) capacitor c=0.0140578f //x=12.95 \
 //y=7.4 //x2=17.275 //y2=4.07
cc_405 ( N_VDD_c_292_n N_noxref_6_c_1215_n ) capacitor c=0.0277022f //x=16.28 \
 //y=7.4 //x2=17.275 //y2=4.07
cc_406 ( N_VDD_M34_noxref_d N_noxref_6_c_1215_n ) capacitor c=5.05307e-19 \
 //x=15.355 //y=5.02 //x2=17.275 //y2=4.07
cc_407 ( N_VDD_M35_noxref_s N_noxref_6_c_1215_n ) capacitor c=0.00363031f \
 //x=16.935 //y=5.02 //x2=17.275 //y2=4.07
cc_408 ( N_VDD_c_290_n N_noxref_6_c_1224_n ) capacitor c=0.00104411f //x=8.14 \
 //y=7.4 //x2=7.51 //y2=4.07
cc_409 ( N_VDD_c_288_n N_noxref_6_c_1192_n ) capacitor c=6.87732e-19 //x=0.74 \
 //y=7.4 //x2=1.85 //y2=2.08
cc_410 ( N_VDD_c_289_n N_noxref_6_c_1192_n ) capacitor c=5.66013e-19 //x=3.33 \
 //y=7.4 //x2=1.85 //y2=2.08
cc_411 ( N_VDD_c_295_p N_noxref_6_c_1227_n ) capacitor c=0.00449316f //x=23.68 \
 //y=7.4 //x2=5.655 //y2=5.155
cc_412 ( N_VDD_c_312_p N_noxref_6_c_1227_n ) capacitor c=4.32228e-19 //x=5.215 \
 //y=7.4 //x2=5.655 //y2=5.155
cc_413 ( N_VDD_c_389_p N_noxref_6_c_1227_n ) capacitor c=4.31906e-19 //x=6.095 \
 //y=7.4 //x2=5.655 //y2=5.155
cc_414 ( N_VDD_M20_noxref_d N_noxref_6_c_1227_n ) capacitor c=0.0115147f \
 //x=5.155 //y=5.02 //x2=5.655 //y2=5.155
cc_415 ( N_VDD_c_289_n N_noxref_6_c_1231_n ) capacitor c=0.00863585f //x=3.33 \
 //y=7.4 //x2=4.945 //y2=5.155
cc_416 ( N_VDD_M19_noxref_s N_noxref_6_c_1231_n ) capacitor c=0.0831083f \
 //x=4.285 //y=5.02 //x2=4.945 //y2=5.155
cc_417 ( N_VDD_c_295_p N_noxref_6_c_1233_n ) capacitor c=0.0044221f //x=23.68 \
 //y=7.4 //x2=6.535 //y2=5.155
cc_418 ( N_VDD_c_389_p N_noxref_6_c_1233_n ) capacitor c=4.31931e-19 //x=6.095 \
 //y=7.4 //x2=6.535 //y2=5.155
cc_419 ( N_VDD_c_426_p N_noxref_6_c_1233_n ) capacitor c=4.31931e-19 //x=6.975 \
 //y=7.4 //x2=6.535 //y2=5.155
cc_420 ( N_VDD_M22_noxref_d N_noxref_6_c_1233_n ) capacitor c=0.0112985f \
 //x=6.035 //y=5.02 //x2=6.535 //y2=5.155
cc_421 ( N_VDD_c_295_p N_noxref_6_c_1237_n ) capacitor c=0.00433242f //x=23.68 \
 //y=7.4 //x2=7.315 //y2=5.155
cc_422 ( N_VDD_c_426_p N_noxref_6_c_1237_n ) capacitor c=7.46626e-19 //x=6.975 \
 //y=7.4 //x2=7.315 //y2=5.155
cc_423 ( N_VDD_c_374_p N_noxref_6_c_1237_n ) capacitor c=0.00198565f //x=7.97 \
 //y=7.4 //x2=7.315 //y2=5.155
cc_424 ( N_VDD_M24_noxref_d N_noxref_6_c_1237_n ) capacitor c=0.0112985f \
 //x=6.915 //y=5.02 //x2=7.315 //y2=5.155
cc_425 ( N_VDD_c_295_p N_noxref_6_c_1195_n ) capacitor c=0.00126142f //x=23.68 \
 //y=7.4 //x2=17.39 //y2=2.08
cc_426 ( N_VDD_c_409_p N_noxref_6_c_1195_n ) capacitor c=2.8777e-19 //x=17.865 \
 //y=7.4 //x2=17.39 //y2=2.08
cc_427 ( N_VDD_c_292_n N_noxref_6_c_1195_n ) capacitor c=0.0156645f //x=16.28 \
 //y=7.4 //x2=17.39 //y2=2.08
cc_428 ( N_VDD_c_290_n N_noxref_6_c_1244_n ) capacitor c=0.0427201f //x=8.14 \
 //y=7.4 //x2=7.395 //y2=4.07
cc_429 ( N_VDD_c_297_p N_noxref_6_M17_noxref_g ) capacitor c=0.00673971f \
 //x=2.465 //y=7.4 //x2=1.89 //y2=6.02
cc_430 ( N_VDD_M16_noxref_d N_noxref_6_M17_noxref_g ) capacitor c=0.015318f \
 //x=1.525 //y=5.02 //x2=1.89 //y2=6.02
cc_431 ( N_VDD_c_297_p N_noxref_6_M18_noxref_g ) capacitor c=0.00672952f \
 //x=2.465 //y=7.4 //x2=2.33 //y2=6.02
cc_432 ( N_VDD_c_289_n N_noxref_6_M18_noxref_g ) capacitor c=0.00928743f \
 //x=3.33 //y=7.4 //x2=2.33 //y2=6.02
cc_433 ( N_VDD_M18_noxref_d N_noxref_6_M18_noxref_g ) capacitor c=0.0430452f \
 //x=2.405 //y=5.02 //x2=2.33 //y2=6.02
cc_434 ( N_VDD_c_409_p N_noxref_6_M35_noxref_g ) capacitor c=0.00726866f \
 //x=17.865 //y=7.4 //x2=17.29 //y2=6.02
cc_435 ( N_VDD_M35_noxref_s N_noxref_6_M35_noxref_g ) capacitor c=0.054195f \
 //x=16.935 //y=5.02 //x2=17.29 //y2=6.02
cc_436 ( N_VDD_c_409_p N_noxref_6_M36_noxref_g ) capacitor c=0.00672952f \
 //x=17.865 //y=7.4 //x2=17.73 //y2=6.02
cc_437 ( N_VDD_M36_noxref_d N_noxref_6_M36_noxref_g ) capacitor c=0.015318f \
 //x=17.805 //y=5.02 //x2=17.73 //y2=6.02
cc_438 ( N_VDD_c_292_n N_noxref_6_c_1254_n ) capacitor c=0.0149273f //x=16.28 \
 //y=7.4 //x2=17.39 //y2=4.7
cc_439 ( N_VDD_c_295_p N_noxref_6_M19_noxref_d ) capacitor c=0.00285091f \
 //x=23.68 //y=7.4 //x2=4.715 //y2=5.02
cc_440 ( N_VDD_c_312_p N_noxref_6_M19_noxref_d ) capacitor c=0.0141016f \
 //x=5.215 //y=7.4 //x2=4.715 //y2=5.02
cc_441 ( N_VDD_M20_noxref_d N_noxref_6_M19_noxref_d ) capacitor c=0.0664752f \
 //x=5.155 //y=5.02 //x2=4.715 //y2=5.02
cc_442 ( N_VDD_c_295_p N_noxref_6_M21_noxref_d ) capacitor c=0.00275186f \
 //x=23.68 //y=7.4 //x2=5.595 //y2=5.02
cc_443 ( N_VDD_c_389_p N_noxref_6_M21_noxref_d ) capacitor c=0.0140346f \
 //x=6.095 //y=7.4 //x2=5.595 //y2=5.02
cc_444 ( N_VDD_c_290_n N_noxref_6_M21_noxref_d ) capacitor c=4.9285e-19 \
 //x=8.14 //y=7.4 //x2=5.595 //y2=5.02
cc_445 ( N_VDD_M19_noxref_s N_noxref_6_M21_noxref_d ) capacitor c=0.00130656f \
 //x=4.285 //y=5.02 //x2=5.595 //y2=5.02
cc_446 ( N_VDD_M20_noxref_d N_noxref_6_M21_noxref_d ) capacitor c=0.0664752f \
 //x=5.155 //y=5.02 //x2=5.595 //y2=5.02
cc_447 ( N_VDD_M22_noxref_d N_noxref_6_M21_noxref_d ) capacitor c=0.0664752f \
 //x=6.035 //y=5.02 //x2=5.595 //y2=5.02
cc_448 ( N_VDD_c_295_p N_noxref_6_M23_noxref_d ) capacitor c=0.00275235f \
 //x=23.68 //y=7.4 //x2=6.475 //y2=5.02
cc_449 ( N_VDD_c_426_p N_noxref_6_M23_noxref_d ) capacitor c=0.014035f \
 //x=6.975 //y=7.4 //x2=6.475 //y2=5.02
cc_450 ( N_VDD_c_290_n N_noxref_6_M23_noxref_d ) capacitor c=0.00939849f \
 //x=8.14 //y=7.4 //x2=6.475 //y2=5.02
cc_451 ( N_VDD_M22_noxref_d N_noxref_6_M23_noxref_d ) capacitor c=0.0664752f \
 //x=6.035 //y=5.02 //x2=6.475 //y2=5.02
cc_452 ( N_VDD_M24_noxref_d N_noxref_6_M23_noxref_d ) capacitor c=0.0664752f \
 //x=6.915 //y=5.02 //x2=6.475 //y2=5.02
cc_453 ( N_VDD_M25_noxref_s N_noxref_6_M23_noxref_d ) capacitor c=3.57641e-19 \
 //x=9.095 //y=5.02 //x2=6.475 //y2=5.02
cc_454 ( N_VDD_c_292_n QN ) capacitor c=0.00151618f //x=16.28 //y=7.4 \
 //x2=18.87 //y2=2.59
cc_455 ( N_VDD_c_293_n QN ) capacitor c=0.0462279f //x=19.61 //y=7.4 \
 //x2=18.87 //y2=2.59
cc_456 ( N_VDD_c_295_p N_QN_c_1494_n ) capacitor c=0.0046595f //x=23.68 \
 //y=7.4 //x2=18.305 //y2=5.2
cc_457 ( N_VDD_c_409_p N_QN_c_1494_n ) capacitor c=4.3394e-19 //x=17.865 \
 //y=7.4 //x2=18.305 //y2=5.2
cc_458 ( N_VDD_c_465_p N_QN_c_1494_n ) capacitor c=4.3394e-19 //x=18.745 \
 //y=7.4 //x2=18.305 //y2=5.2
cc_459 ( N_VDD_M36_noxref_d N_QN_c_1494_n ) capacitor c=0.0128485f //x=17.805 \
 //y=5.02 //x2=18.305 //y2=5.2
cc_460 ( N_VDD_c_292_n N_QN_c_1498_n ) capacitor c=0.00985474f //x=16.28 \
 //y=7.4 //x2=17.595 //y2=5.2
cc_461 ( N_VDD_M35_noxref_s N_QN_c_1498_n ) capacitor c=0.087833f //x=16.935 \
 //y=5.02 //x2=17.595 //y2=5.2
cc_462 ( N_VDD_c_295_p N_QN_c_1500_n ) capacitor c=0.0031203f //x=23.68 \
 //y=7.4 //x2=18.785 //y2=5.2
cc_463 ( N_VDD_c_465_p N_QN_c_1500_n ) capacitor c=7.21492e-19 //x=18.745 \
 //y=7.4 //x2=18.785 //y2=5.2
cc_464 ( N_VDD_M38_noxref_d N_QN_c_1500_n ) capacitor c=0.0163486f //x=18.685 \
 //y=5.02 //x2=18.785 //y2=5.2
cc_465 ( N_VDD_c_295_p N_QN_c_1478_n ) capacitor c=9.35768e-19 //x=23.68 \
 //y=7.4 //x2=20.72 //y2=2.08
cc_466 ( N_VDD_c_293_n N_QN_c_1478_n ) capacitor c=0.0166656f //x=19.61 \
 //y=7.4 //x2=20.72 //y2=2.08
cc_467 ( N_VDD_M39_noxref_s N_QN_c_1478_n ) capacitor c=0.0125045f //x=20.565 \
 //y=5.02 //x2=20.72 //y2=2.08
cc_468 ( N_VDD_c_475_p N_QN_M39_noxref_g ) capacitor c=0.00749687f //x=21.495 \
 //y=7.4 //x2=20.92 //y2=6.02
cc_469 ( N_VDD_M39_noxref_s N_QN_M39_noxref_g ) capacitor c=0.0477201f \
 //x=20.565 //y=5.02 //x2=20.92 //y2=6.02
cc_470 ( N_VDD_c_475_p N_QN_M40_noxref_g ) capacitor c=0.00675175f //x=21.495 \
 //y=7.4 //x2=21.36 //y2=6.02
cc_471 ( N_VDD_M40_noxref_d N_QN_M40_noxref_g ) capacitor c=0.015318f \
 //x=21.435 //y=5.02 //x2=21.36 //y2=6.02
cc_472 ( N_VDD_c_293_n N_QN_c_1510_n ) capacitor c=0.0076931f //x=19.61 \
 //y=7.4 //x2=20.995 //y2=4.79
cc_473 ( N_VDD_M39_noxref_s N_QN_c_1510_n ) capacitor c=0.00446175f //x=20.565 \
 //y=5.02 //x2=20.995 //y2=4.79
cc_474 ( N_VDD_c_295_p N_QN_M35_noxref_d ) capacitor c=0.00287944f //x=23.68 \
 //y=7.4 //x2=17.365 //y2=5.02
cc_475 ( N_VDD_c_409_p N_QN_M35_noxref_d ) capacitor c=0.014004f //x=17.865 \
 //y=7.4 //x2=17.365 //y2=5.02
cc_476 ( N_VDD_c_293_n N_QN_M35_noxref_d ) capacitor c=6.94454e-19 //x=19.61 \
 //y=7.4 //x2=17.365 //y2=5.02
cc_477 ( N_VDD_M36_noxref_d N_QN_M35_noxref_d ) capacitor c=0.0664752f \
 //x=17.805 //y=5.02 //x2=17.365 //y2=5.02
cc_478 ( N_VDD_c_295_p N_QN_M37_noxref_d ) capacitor c=0.00294217f //x=23.68 \
 //y=7.4 //x2=18.245 //y2=5.02
cc_479 ( N_VDD_c_465_p N_QN_M37_noxref_d ) capacitor c=0.0138379f //x=18.745 \
 //y=7.4 //x2=18.245 //y2=5.02
cc_480 ( N_VDD_c_293_n N_QN_M37_noxref_d ) capacitor c=0.0120541f //x=19.61 \
 //y=7.4 //x2=18.245 //y2=5.02
cc_481 ( N_VDD_M35_noxref_s N_QN_M37_noxref_d ) capacitor c=0.00111971f \
 //x=16.935 //y=5.02 //x2=18.245 //y2=5.02
cc_482 ( N_VDD_M36_noxref_d N_QN_M37_noxref_d ) capacitor c=0.0664752f \
 //x=17.805 //y=5.02 //x2=18.245 //y2=5.02
cc_483 ( N_VDD_M38_noxref_d N_QN_M37_noxref_d ) capacitor c=0.0664752f \
 //x=18.685 //y=5.02 //x2=18.245 //y2=5.02
cc_484 ( N_VDD_M39_noxref_s N_QN_M37_noxref_d ) capacitor c=3.73257e-19 \
 //x=20.565 //y=5.02 //x2=18.245 //y2=5.02
cc_485 ( N_VDD_c_295_p N_SN_c_1631_n ) capacitor c=2.03486e-19 //x=23.68 \
 //y=7.4 //x2=10.36 //y2=2.08
cc_486 ( N_VDD_c_290_n N_SN_c_1631_n ) capacitor c=6.15069e-19 //x=8.14 \
 //y=7.4 //x2=10.36 //y2=2.08
cc_487 ( N_VDD_c_295_p N_SN_c_1632_n ) capacitor c=2.07998e-19 //x=23.68 \
 //y=7.4 //x2=21.83 //y2=2.08
cc_488 ( N_VDD_c_293_n N_SN_c_1632_n ) capacitor c=7.34553e-19 //x=19.61 \
 //y=7.4 //x2=21.83 //y2=2.08
cc_489 ( N_VDD_c_337_p N_SN_M27_noxref_g ) capacitor c=0.00676195f //x=10.905 \
 //y=7.4 //x2=10.33 //y2=6.02
cc_490 ( N_VDD_M26_noxref_d N_SN_M27_noxref_g ) capacitor c=0.015318f \
 //x=9.965 //y=5.02 //x2=10.33 //y2=6.02
cc_491 ( N_VDD_c_337_p N_SN_M28_noxref_g ) capacitor c=0.00675175f //x=10.905 \
 //y=7.4 //x2=10.77 //y2=6.02
cc_492 ( N_VDD_M28_noxref_d N_SN_M28_noxref_g ) capacitor c=0.015318f \
 //x=10.845 //y=5.02 //x2=10.77 //y2=6.02
cc_493 ( N_VDD_c_500_p N_SN_M41_noxref_g ) capacitor c=0.00676195f //x=22.375 \
 //y=7.4 //x2=21.8 //y2=6.02
cc_494 ( N_VDD_M40_noxref_d N_SN_M41_noxref_g ) capacitor c=0.015318f \
 //x=21.435 //y=5.02 //x2=21.8 //y2=6.02
cc_495 ( N_VDD_c_500_p N_SN_M42_noxref_g ) capacitor c=0.00675175f //x=22.375 \
 //y=7.4 //x2=22.24 //y2=6.02
cc_496 ( N_VDD_M42_noxref_d N_SN_M42_noxref_g ) capacitor c=0.015318f \
 //x=22.315 //y=5.02 //x2=22.24 //y2=6.02
cc_497 ( N_VDD_c_295_p N_noxref_9_c_1849_n ) capacitor c=0.040523f //x=23.68 \
 //y=7.4 //x2=22.825 //y2=3.7
cc_498 ( N_VDD_c_293_n N_noxref_9_c_1849_n ) capacitor c=0.0109524f //x=19.61 \
 //y=7.4 //x2=22.825 //y2=3.7
cc_499 ( N_VDD_M38_noxref_d N_noxref_9_c_1849_n ) capacitor c=4.00436e-19 \
 //x=18.685 //y=5.02 //x2=22.825 //y2=3.7
cc_500 ( N_VDD_M39_noxref_s N_noxref_9_c_1849_n ) capacitor c=9.16752e-19 \
 //x=20.565 //y=5.02 //x2=22.825 //y2=3.7
cc_501 ( N_VDD_c_290_n N_noxref_9_c_1850_n ) capacitor c=7.21808e-19 //x=8.14 \
 //y=7.4 //x2=6.66 //y2=2.08
cc_502 ( N_VDD_c_291_n N_noxref_9_c_1851_n ) capacitor c=6.21611e-19 //x=12.95 \
 //y=7.4 //x2=11.47 //y2=2.08
cc_503 ( N_VDD_c_295_p N_noxref_9_c_1864_n ) capacitor c=0.00453473f //x=23.68 \
 //y=7.4 //x2=14.975 //y2=5.2
cc_504 ( N_VDD_c_351_p N_noxref_9_c_1864_n ) capacitor c=4.48391e-19 \
 //x=14.535 //y=7.4 //x2=14.975 //y2=5.2
cc_505 ( N_VDD_c_393_p N_noxref_9_c_1864_n ) capacitor c=4.48377e-19 \
 //x=15.415 //y=7.4 //x2=14.975 //y2=5.2
cc_506 ( N_VDD_M32_noxref_d N_noxref_9_c_1864_n ) capacitor c=0.0124506f \
 //x=14.475 //y=5.02 //x2=14.975 //y2=5.2
cc_507 ( N_VDD_c_291_n N_noxref_9_c_1868_n ) capacitor c=0.00985474f //x=12.95 \
 //y=7.4 //x2=14.265 //y2=5.2
cc_508 ( N_VDD_M31_noxref_s N_noxref_9_c_1868_n ) capacitor c=0.087833f \
 //x=13.605 //y=5.02 //x2=14.265 //y2=5.2
cc_509 ( N_VDD_c_295_p N_noxref_9_c_1870_n ) capacitor c=0.00307195f //x=23.68 \
 //y=7.4 //x2=15.455 //y2=5.2
cc_510 ( N_VDD_c_393_p N_noxref_9_c_1870_n ) capacitor c=7.73167e-19 \
 //x=15.415 //y=7.4 //x2=15.455 //y2=5.2
cc_511 ( N_VDD_M34_noxref_d N_noxref_9_c_1870_n ) capacitor c=0.0161518f \
 //x=15.355 //y=5.02 //x2=15.455 //y2=5.2
cc_512 ( N_VDD_M35_noxref_s N_noxref_9_c_1870_n ) capacitor c=2.44532e-19 \
 //x=16.935 //y=5.02 //x2=15.455 //y2=5.2
cc_513 ( N_VDD_c_291_n N_noxref_9_c_1853_n ) capacitor c=0.00151618f //x=12.95 \
 //y=7.4 //x2=15.54 //y2=3.7
cc_514 ( N_VDD_c_292_n N_noxref_9_c_1853_n ) capacitor c=0.044931f //x=16.28 \
 //y=7.4 //x2=15.54 //y2=3.7
cc_515 ( N_VDD_c_287_n N_noxref_9_c_1854_n ) capacitor c=8.81482e-19 //x=23.68 \
 //y=7.4 //x2=22.94 //y2=2.08
cc_516 ( N_VDD_c_426_p N_noxref_9_M23_noxref_g ) capacitor c=0.00675175f \
 //x=6.975 //y=7.4 //x2=6.4 //y2=6.02
cc_517 ( N_VDD_M22_noxref_d N_noxref_9_M23_noxref_g ) capacitor c=0.015318f \
 //x=6.035 //y=5.02 //x2=6.4 //y2=6.02
cc_518 ( N_VDD_c_426_p N_noxref_9_M24_noxref_g ) capacitor c=0.00675379f \
 //x=6.975 //y=7.4 //x2=6.84 //y2=6.02
cc_519 ( N_VDD_M24_noxref_d N_noxref_9_M24_noxref_g ) capacitor c=0.0394719f \
 //x=6.915 //y=5.02 //x2=6.84 //y2=6.02
cc_520 ( N_VDD_c_343_p N_noxref_9_M29_noxref_g ) capacitor c=0.00675175f \
 //x=11.785 //y=7.4 //x2=11.21 //y2=6.02
cc_521 ( N_VDD_M28_noxref_d N_noxref_9_M29_noxref_g ) capacitor c=0.015318f \
 //x=10.845 //y=5.02 //x2=11.21 //y2=6.02
cc_522 ( N_VDD_c_343_p N_noxref_9_M30_noxref_g ) capacitor c=0.00675379f \
 //x=11.785 //y=7.4 //x2=11.65 //y2=6.02
cc_523 ( N_VDD_M30_noxref_d N_noxref_9_M30_noxref_g ) capacitor c=0.0394719f \
 //x=11.725 //y=5.02 //x2=11.65 //y2=6.02
cc_524 ( N_VDD_c_531_p N_noxref_9_M43_noxref_g ) capacitor c=0.00675175f \
 //x=23.255 //y=7.4 //x2=22.68 //y2=6.02
cc_525 ( N_VDD_M42_noxref_d N_noxref_9_M43_noxref_g ) capacitor c=0.015318f \
 //x=22.315 //y=5.02 //x2=22.68 //y2=6.02
cc_526 ( N_VDD_c_531_p N_noxref_9_M44_noxref_g ) capacitor c=0.00675379f \
 //x=23.255 //y=7.4 //x2=23.12 //y2=6.02
cc_527 ( N_VDD_M44_noxref_d N_noxref_9_M44_noxref_g ) capacitor c=0.0394719f \
 //x=23.195 //y=5.02 //x2=23.12 //y2=6.02
cc_528 ( N_VDD_c_295_p N_noxref_9_M31_noxref_d ) capacitor c=0.00275225f \
 //x=23.68 //y=7.4 //x2=14.035 //y2=5.02
cc_529 ( N_VDD_c_351_p N_noxref_9_M31_noxref_d ) capacitor c=0.0140317f \
 //x=14.535 //y=7.4 //x2=14.035 //y2=5.02
cc_530 ( N_VDD_c_292_n N_noxref_9_M31_noxref_d ) capacitor c=6.94454e-19 \
 //x=16.28 //y=7.4 //x2=14.035 //y2=5.02
cc_531 ( N_VDD_M32_noxref_d N_noxref_9_M31_noxref_d ) capacitor c=0.0664752f \
 //x=14.475 //y=5.02 //x2=14.035 //y2=5.02
cc_532 ( N_VDD_c_295_p N_noxref_9_M33_noxref_d ) capacitor c=0.00285083f \
 //x=23.68 //y=7.4 //x2=14.915 //y2=5.02
cc_533 ( N_VDD_c_393_p N_noxref_9_M33_noxref_d ) capacitor c=0.0140984f \
 //x=15.415 //y=7.4 //x2=14.915 //y2=5.02
cc_534 ( N_VDD_c_292_n N_noxref_9_M33_noxref_d ) capacitor c=0.0120541f \
 //x=16.28 //y=7.4 //x2=14.915 //y2=5.02
cc_535 ( N_VDD_M31_noxref_s N_noxref_9_M33_noxref_d ) capacitor c=0.00111971f \
 //x=13.605 //y=5.02 //x2=14.915 //y2=5.02
cc_536 ( N_VDD_M32_noxref_d N_noxref_9_M33_noxref_d ) capacitor c=0.0664752f \
 //x=14.475 //y=5.02 //x2=14.915 //y2=5.02
cc_537 ( N_VDD_M34_noxref_d N_noxref_9_M33_noxref_d ) capacitor c=0.0664752f \
 //x=15.355 //y=5.02 //x2=14.915 //y2=5.02
cc_538 ( N_VDD_M35_noxref_s N_noxref_9_M33_noxref_d ) capacitor c=4.54516e-19 \
 //x=16.935 //y=5.02 //x2=14.915 //y2=5.02
cc_539 ( N_VDD_c_295_p N_noxref_10_c_2170_n ) capacitor c=0.0215075f //x=23.68 \
 //y=7.4 //x2=23.565 //y2=3.33
cc_540 ( N_VDD_c_292_n N_noxref_10_c_2172_n ) capacitor c=9.96229e-19 \
 //x=16.28 //y=7.4 //x2=18.13 //y2=2.08
cc_541 ( N_VDD_c_293_n N_noxref_10_c_2172_n ) capacitor c=7.1514e-19 //x=19.61 \
 //y=7.4 //x2=18.13 //y2=2.08
cc_542 ( N_VDD_c_295_p N_noxref_10_c_2179_n ) capacitor c=0.00457327f \
 //x=23.68 //y=7.4 //x2=21.935 //y2=5.155
cc_543 ( N_VDD_c_475_p N_noxref_10_c_2179_n ) capacitor c=4.18223e-19 \
 //x=21.495 //y=7.4 //x2=21.935 //y2=5.155
cc_544 ( N_VDD_c_500_p N_noxref_10_c_2179_n ) capacitor c=4.18223e-19 \
 //x=22.375 //y=7.4 //x2=21.935 //y2=5.155
cc_545 ( N_VDD_M40_noxref_d N_noxref_10_c_2179_n ) capacitor c=0.0116565f \
 //x=21.435 //y=5.02 //x2=21.935 //y2=5.155
cc_546 ( N_VDD_c_293_n N_noxref_10_c_2183_n ) capacitor c=0.00863585f \
 //x=19.61 //y=7.4 //x2=21.225 //y2=5.155
cc_547 ( N_VDD_M39_noxref_s N_noxref_10_c_2183_n ) capacitor c=0.0831083f \
 //x=20.565 //y=5.02 //x2=21.225 //y2=5.155
cc_548 ( N_VDD_c_295_p N_noxref_10_c_2185_n ) capacitor c=0.00454915f \
 //x=23.68 //y=7.4 //x2=22.815 //y2=5.155
cc_549 ( N_VDD_c_500_p N_noxref_10_c_2185_n ) capacitor c=4.18223e-19 \
 //x=22.375 //y=7.4 //x2=22.815 //y2=5.155
cc_550 ( N_VDD_c_531_p N_noxref_10_c_2185_n ) capacitor c=4.18223e-19 \
 //x=23.255 //y=7.4 //x2=22.815 //y2=5.155
cc_551 ( N_VDD_M42_noxref_d N_noxref_10_c_2185_n ) capacitor c=0.0116565f \
 //x=22.315 //y=5.02 //x2=22.815 //y2=5.155
cc_552 ( N_VDD_c_295_p N_noxref_10_c_2189_n ) capacitor c=0.00455815f \
 //x=23.68 //y=7.4 //x2=23.595 //y2=5.155
cc_553 ( N_VDD_c_531_p N_noxref_10_c_2189_n ) capacitor c=6.98646e-19 \
 //x=23.255 //y=7.4 //x2=23.595 //y2=5.155
cc_554 ( N_VDD_c_287_n N_noxref_10_c_2189_n ) capacitor c=0.00179956f \
 //x=23.68 //y=7.4 //x2=23.595 //y2=5.155
cc_555 ( N_VDD_M44_noxref_d N_noxref_10_c_2189_n ) capacitor c=0.0117481f \
 //x=23.195 //y=5.02 //x2=23.595 //y2=5.155
cc_556 ( N_VDD_c_287_n N_noxref_10_c_2193_n ) capacitor c=0.046173f //x=23.68 \
 //y=7.4 //x2=23.68 //y2=3.33
cc_557 ( N_VDD_c_465_p N_noxref_10_M37_noxref_g ) capacitor c=0.00673971f \
 //x=18.745 //y=7.4 //x2=18.17 //y2=6.02
cc_558 ( N_VDD_M36_noxref_d N_noxref_10_M37_noxref_g ) capacitor c=0.015318f \
 //x=17.805 //y=5.02 //x2=18.17 //y2=6.02
cc_559 ( N_VDD_c_465_p N_noxref_10_M38_noxref_g ) capacitor c=0.00672952f \
 //x=18.745 //y=7.4 //x2=18.61 //y2=6.02
cc_560 ( N_VDD_c_293_n N_noxref_10_M38_noxref_g ) capacitor c=0.00928743f \
 //x=19.61 //y=7.4 //x2=18.61 //y2=6.02
cc_561 ( N_VDD_M38_noxref_d N_noxref_10_M38_noxref_g ) capacitor c=0.0430452f \
 //x=18.685 //y=5.02 //x2=18.61 //y2=6.02
cc_562 ( N_VDD_c_295_p N_noxref_10_M39_noxref_d ) capacitor c=0.00294223f \
 //x=23.68 //y=7.4 //x2=20.995 //y2=5.02
cc_563 ( N_VDD_c_475_p N_noxref_10_M39_noxref_d ) capacitor c=0.0138437f \
 //x=21.495 //y=7.4 //x2=20.995 //y2=5.02
cc_564 ( N_VDD_M40_noxref_d N_noxref_10_M39_noxref_d ) capacitor c=0.0664752f \
 //x=21.435 //y=5.02 //x2=20.995 //y2=5.02
cc_565 ( N_VDD_c_295_p N_noxref_10_M41_noxref_d ) capacitor c=0.00294223f \
 //x=23.68 //y=7.4 //x2=21.875 //y2=5.02
cc_566 ( N_VDD_c_500_p N_noxref_10_M41_noxref_d ) capacitor c=0.0138437f \
 //x=22.375 //y=7.4 //x2=21.875 //y2=5.02
cc_567 ( N_VDD_c_287_n N_noxref_10_M41_noxref_d ) capacitor c=4.9285e-19 \
 //x=23.68 //y=7.4 //x2=21.875 //y2=5.02
cc_568 ( N_VDD_M39_noxref_s N_noxref_10_M41_noxref_d ) capacitor c=0.00130656f \
 //x=20.565 //y=5.02 //x2=21.875 //y2=5.02
cc_569 ( N_VDD_M40_noxref_d N_noxref_10_M41_noxref_d ) capacitor c=0.0664752f \
 //x=21.435 //y=5.02 //x2=21.875 //y2=5.02
cc_570 ( N_VDD_M42_noxref_d N_noxref_10_M41_noxref_d ) capacitor c=0.0664752f \
 //x=22.315 //y=5.02 //x2=21.875 //y2=5.02
cc_571 ( N_VDD_c_295_p N_noxref_10_M43_noxref_d ) capacitor c=0.00293548f \
 //x=23.68 //y=7.4 //x2=22.755 //y2=5.02
cc_572 ( N_VDD_c_531_p N_noxref_10_M43_noxref_d ) capacitor c=0.0137718f \
 //x=23.255 //y=7.4 //x2=22.755 //y2=5.02
cc_573 ( N_VDD_c_287_n N_noxref_10_M43_noxref_d ) capacitor c=0.00963505f \
 //x=23.68 //y=7.4 //x2=22.755 //y2=5.02
cc_574 ( N_VDD_M42_noxref_d N_noxref_10_M43_noxref_d ) capacitor c=0.0664752f \
 //x=22.315 //y=5.02 //x2=22.755 //y2=5.02
cc_575 ( N_VDD_M44_noxref_d N_noxref_10_M43_noxref_d ) capacitor c=0.0664752f \
 //x=23.195 //y=5.02 //x2=22.755 //y2=5.02
cc_576 ( N_VDD_c_295_p N_D_c_2340_n ) capacitor c=0.00140404f //x=23.68 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_577 ( N_VDD_c_296_p N_D_c_2340_n ) capacitor c=2.63811e-19 //x=1.585 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_578 ( N_VDD_c_288_n N_D_c_2340_n ) capacitor c=0.01673f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_579 ( N_VDD_c_296_p N_D_M15_noxref_g ) capacitor c=0.00726866f //x=1.585 \
 //y=7.4 //x2=1.01 //y2=6.02
cc_580 ( N_VDD_M15_noxref_s N_D_M15_noxref_g ) capacitor c=0.054195f //x=0.655 \
 //y=5.02 //x2=1.01 //y2=6.02
cc_581 ( N_VDD_c_296_p N_D_M16_noxref_g ) capacitor c=0.00672952f //x=1.585 \
 //y=7.4 //x2=1.45 //y2=6.02
cc_582 ( N_VDD_M16_noxref_d N_D_M16_noxref_g ) capacitor c=0.015318f //x=1.525 \
 //y=5.02 //x2=1.45 //y2=6.02
cc_583 ( N_VDD_c_288_n N_D_c_2358_n ) capacitor c=0.0292267f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=4.7
cc_584 ( N_noxref_3_c_597_n N_noxref_4_c_832_n ) capacitor c=0.00564994f \
 //x=9.135 //y=2.59 //x2=12.325 //y2=2.59
cc_585 ( N_noxref_3_M26_noxref_g N_noxref_4_c_847_n ) capacitor c=0.0168349f \
 //x=9.89 //y=6.02 //x2=10.465 //y2=5.155
cc_586 ( N_noxref_3_M25_noxref_g N_noxref_4_c_851_n ) capacitor c=0.0213876f \
 //x=9.45 //y=6.02 //x2=9.755 //y2=5.155
cc_587 ( N_noxref_3_c_675_p N_noxref_4_c_851_n ) capacitor c=0.00428486f \
 //x=9.815 //y=4.79 //x2=9.755 //y2=5.155
cc_588 ( N_noxref_3_M26_noxref_g N_noxref_4_M25_noxref_d ) capacitor \
 c=0.0180032f //x=9.89 //y=6.02 //x2=9.525 //y2=5.02
cc_589 ( N_noxref_3_c_597_n N_CLK_c_994_n ) capacitor c=0.00559244f //x=9.135 \
 //y=2.59 //x2=14.685 //y2=4.44
cc_590 ( N_noxref_3_c_607_n N_CLK_c_994_n ) capacitor c=0.0208709f //x=9.25 \
 //y=2.08 //x2=14.685 //y2=4.44
cc_591 ( N_noxref_3_c_659_n N_CLK_c_994_n ) capacitor c=0.0166984f //x=9.525 \
 //y=4.79 //x2=14.685 //y2=4.44
cc_592 ( N_noxref_3_c_597_n N_CLK_c_1005_n ) capacitor c=6.22349e-19 //x=9.135 \
 //y=2.59 //x2=5.665 //y2=4.44
cc_593 ( N_noxref_3_c_606_n N_CLK_c_1005_n ) capacitor c=0.00551083f //x=4.44 \
 //y=2.08 //x2=5.665 //y2=4.44
cc_594 ( N_noxref_3_c_597_n N_CLK_c_991_n ) capacitor c=0.0273718f //x=9.135 \
 //y=2.59 //x2=5.55 //y2=2.08
cc_595 ( N_noxref_3_c_601_n N_CLK_c_991_n ) capacitor c=0.00103784f //x=4.705 \
 //y=2.59 //x2=5.55 //y2=2.08
cc_596 ( N_noxref_3_c_604_n N_CLK_c_991_n ) capacitor c=4.97515e-19 //x=2.59 \
 //y=2.59 //x2=5.55 //y2=2.08
cc_597 ( N_noxref_3_c_606_n N_CLK_c_991_n ) capacitor c=0.0511511f //x=4.44 \
 //y=2.08 //x2=5.55 //y2=2.08
cc_598 ( N_noxref_3_c_612_n N_CLK_c_991_n ) capacitor c=0.00238338f //x=4.14 \
 //y=1.915 //x2=5.55 //y2=2.08
cc_599 ( N_noxref_3_c_687_p N_CLK_c_991_n ) capacitor c=0.00147352f //x=5.005 \
 //y=4.79 //x2=5.55 //y2=2.08
cc_600 ( N_noxref_3_c_657_n N_CLK_c_991_n ) capacitor c=0.00141297f //x=4.715 \
 //y=4.79 //x2=5.55 //y2=2.08
cc_601 ( N_noxref_3_M19_noxref_g N_CLK_M21_noxref_g ) capacitor c=0.0105869f \
 //x=4.64 //y=6.02 //x2=5.52 //y2=6.02
cc_602 ( N_noxref_3_M20_noxref_g N_CLK_M21_noxref_g ) capacitor c=0.10632f \
 //x=5.08 //y=6.02 //x2=5.52 //y2=6.02
cc_603 ( N_noxref_3_M20_noxref_g N_CLK_M22_noxref_g ) capacitor c=0.0101598f \
 //x=5.08 //y=6.02 //x2=5.96 //y2=6.02
cc_604 ( N_noxref_3_c_608_n N_CLK_c_1034_n ) capacitor c=5.72482e-19 //x=4.14 \
 //y=0.875 //x2=5.115 //y2=0.91
cc_605 ( N_noxref_3_c_610_n N_CLK_c_1034_n ) capacitor c=0.00149976f //x=4.14 \
 //y=1.22 //x2=5.115 //y2=0.91
cc_606 ( N_noxref_3_c_615_n N_CLK_c_1034_n ) capacitor c=0.0160123f //x=4.67 \
 //y=0.875 //x2=5.115 //y2=0.91
cc_607 ( N_noxref_3_c_611_n N_CLK_c_1037_n ) capacitor c=0.00111227f //x=4.14 \
 //y=1.53 //x2=5.115 //y2=1.22
cc_608 ( N_noxref_3_c_617_n N_CLK_c_1037_n ) capacitor c=0.0124075f //x=4.67 \
 //y=1.22 //x2=5.115 //y2=1.22
cc_609 ( N_noxref_3_c_615_n N_CLK_c_1039_n ) capacitor c=0.00103227f //x=4.67 \
 //y=0.875 //x2=5.64 //y2=0.91
cc_610 ( N_noxref_3_c_617_n N_CLK_c_1040_n ) capacitor c=0.0010154f //x=4.67 \
 //y=1.22 //x2=5.64 //y2=1.22
cc_611 ( N_noxref_3_c_617_n N_CLK_c_1041_n ) capacitor c=9.23422e-19 //x=4.67 \
 //y=1.22 //x2=5.64 //y2=1.45
cc_612 ( N_noxref_3_c_597_n N_CLK_c_1042_n ) capacitor c=0.00233308f //x=9.135 \
 //y=2.59 //x2=5.64 //y2=1.915
cc_613 ( N_noxref_3_c_606_n N_CLK_c_1042_n ) capacitor c=0.00231304f //x=4.44 \
 //y=2.08 //x2=5.64 //y2=1.915
cc_614 ( N_noxref_3_c_612_n N_CLK_c_1042_n ) capacitor c=0.00964411f //x=4.14 \
 //y=1.915 //x2=5.64 //y2=1.915
cc_615 ( N_noxref_3_c_606_n N_CLK_c_1045_n ) capacitor c=0.00183762f //x=4.44 \
 //y=2.08 //x2=5.55 //y2=4.7
cc_616 ( N_noxref_3_c_687_p N_CLK_c_1045_n ) capacitor c=0.0168581f //x=5.005 \
 //y=4.79 //x2=5.55 //y2=4.7
cc_617 ( N_noxref_3_c_657_n N_CLK_c_1045_n ) capacitor c=0.00484466f //x=4.715 \
 //y=4.79 //x2=5.55 //y2=4.7
cc_618 ( N_noxref_3_c_591_n N_noxref_6_c_1189_n ) capacitor c=0.0375273f \
 //x=4.295 //y=2.59 //x2=7.28 //y2=4.07
cc_619 ( N_noxref_3_c_595_n N_noxref_6_c_1189_n ) capacitor c=0.0053071f \
 //x=2.705 //y=2.59 //x2=7.28 //y2=4.07
cc_620 ( N_noxref_3_c_601_n N_noxref_6_c_1189_n ) capacitor c=0.0491486f \
 //x=4.705 //y=2.59 //x2=7.28 //y2=4.07
cc_621 ( N_noxref_3_c_632_n N_noxref_6_c_1189_n ) capacitor c=0.0129784f \
 //x=2.025 //y=5.2 //x2=7.28 //y2=4.07
cc_622 ( N_noxref_3_c_710_p N_noxref_6_c_1189_n ) capacitor c=0.00308569f \
 //x=2.235 //y=1.655 //x2=7.28 //y2=4.07
cc_623 ( N_noxref_3_c_604_n N_noxref_6_c_1189_n ) capacitor c=0.0280719f \
 //x=2.59 //y=2.59 //x2=7.28 //y2=4.07
cc_624 ( N_noxref_3_c_606_n N_noxref_6_c_1189_n ) capacitor c=0.0283241f \
 //x=4.44 //y=2.08 //x2=7.28 //y2=4.07
cc_625 ( N_noxref_3_c_657_n N_noxref_6_c_1189_n ) capacitor c=0.0116469f \
 //x=4.715 //y=4.79 //x2=7.28 //y2=4.07
cc_626 ( N_noxref_3_c_632_n N_noxref_6_c_1191_n ) capacitor c=0.00198571f \
 //x=2.025 //y=5.2 //x2=1.965 //y2=4.07
cc_627 ( N_noxref_3_c_604_n N_noxref_6_c_1191_n ) capacitor c=0.00179385f \
 //x=2.59 //y=2.59 //x2=1.965 //y2=4.07
cc_628 ( N_noxref_3_c_597_n N_noxref_6_c_1215_n ) capacitor c=0.00635883f \
 //x=9.135 //y=2.59 //x2=17.275 //y2=4.07
cc_629 ( N_noxref_3_c_607_n N_noxref_6_c_1215_n ) capacitor c=0.0194977f \
 //x=9.25 //y=2.08 //x2=17.275 //y2=4.07
cc_630 ( N_noxref_3_c_597_n N_noxref_6_c_1224_n ) capacitor c=3.09116e-19 \
 //x=9.135 //y=2.59 //x2=7.51 //y2=4.07
cc_631 ( N_noxref_3_c_607_n N_noxref_6_c_1224_n ) capacitor c=3.49381e-19 \
 //x=9.25 //y=2.08 //x2=7.51 //y2=4.07
cc_632 ( N_noxref_3_c_632_n N_noxref_6_c_1284_n ) capacitor c=0.0129794f \
 //x=2.025 //y=5.2 //x2=1.85 //y2=4.535
cc_633 ( N_noxref_3_c_604_n N_noxref_6_c_1284_n ) capacitor c=0.0101115f \
 //x=2.59 //y=2.59 //x2=1.85 //y2=4.535
cc_634 ( N_noxref_3_c_595_n N_noxref_6_c_1192_n ) capacitor c=0.00691549f \
 //x=2.705 //y=2.59 //x2=1.85 //y2=2.08
cc_635 ( N_noxref_3_c_604_n N_noxref_6_c_1192_n ) capacitor c=0.0786485f \
 //x=2.59 //y=2.59 //x2=1.85 //y2=2.08
cc_636 ( N_noxref_3_c_606_n N_noxref_6_c_1192_n ) capacitor c=8.97258e-19 \
 //x=4.44 //y=2.08 //x2=1.85 //y2=2.08
cc_637 ( N_noxref_3_M20_noxref_g N_noxref_6_c_1227_n ) capacitor c=0.0178794f \
 //x=5.08 //y=6.02 //x2=5.655 //y2=5.155
cc_638 ( N_noxref_3_c_604_n N_noxref_6_c_1231_n ) capacitor c=2.97874e-19 \
 //x=2.59 //y=2.59 //x2=4.945 //y2=5.155
cc_639 ( N_noxref_3_M19_noxref_g N_noxref_6_c_1231_n ) capacitor c=0.0213876f \
 //x=4.64 //y=6.02 //x2=4.945 //y2=5.155
cc_640 ( N_noxref_3_c_687_p N_noxref_6_c_1231_n ) capacitor c=0.00429591f \
 //x=5.005 //y=4.79 //x2=4.945 //y2=5.155
cc_641 ( N_noxref_3_c_597_n N_noxref_6_c_1293_n ) capacitor c=0.011558f \
 //x=9.135 //y=2.59 //x2=7 //y2=1.665
cc_642 ( N_noxref_3_c_597_n N_noxref_6_c_1294_n ) capacitor c=0.024834f \
 //x=9.135 //y=2.59 //x2=7.397 //y2=3.905
cc_643 ( N_noxref_3_c_607_n N_noxref_6_c_1294_n ) capacitor c=0.0148121f \
 //x=9.25 //y=2.08 //x2=7.397 //y2=3.905
cc_644 ( N_noxref_3_c_632_n N_noxref_6_M17_noxref_g ) capacitor c=0.0166421f \
 //x=2.025 //y=5.2 //x2=1.89 //y2=6.02
cc_645 ( N_noxref_3_M17_noxref_d N_noxref_6_M17_noxref_g ) capacitor \
 c=0.0173476f //x=1.965 //y=5.02 //x2=1.89 //y2=6.02
cc_646 ( N_noxref_3_c_638_n N_noxref_6_M18_noxref_g ) capacitor c=0.0199348f \
 //x=2.505 //y=5.2 //x2=2.33 //y2=6.02
cc_647 ( N_noxref_3_M17_noxref_d N_noxref_6_M18_noxref_g ) capacitor \
 c=0.0179769f //x=1.965 //y=5.02 //x2=2.33 //y2=6.02
cc_648 ( N_noxref_3_M1_noxref_d N_noxref_6_c_1300_n ) capacitor c=0.00217566f \
 //x=1.96 //y=0.905 //x2=1.885 //y2=0.905
cc_649 ( N_noxref_3_M1_noxref_d N_noxref_6_c_1301_n ) capacitor c=0.0034598f \
 //x=1.96 //y=0.905 //x2=1.885 //y2=1.25
cc_650 ( N_noxref_3_M1_noxref_d N_noxref_6_c_1302_n ) capacitor c=0.0065582f \
 //x=1.96 //y=0.905 //x2=1.885 //y2=1.56
cc_651 ( N_noxref_3_c_604_n N_noxref_6_c_1303_n ) capacitor c=0.0142673f \
 //x=2.59 //y=2.59 //x2=2.255 //y2=4.79
cc_652 ( N_noxref_3_c_740_p N_noxref_6_c_1303_n ) capacitor c=0.00408717f \
 //x=2.11 //y=5.2 //x2=2.255 //y2=4.79
cc_653 ( N_noxref_3_M1_noxref_d N_noxref_6_c_1305_n ) capacitor c=0.00241102f \
 //x=1.96 //y=0.905 //x2=2.26 //y2=0.75
cc_654 ( N_noxref_3_c_603_n N_noxref_6_c_1306_n ) capacitor c=0.00359704f \
 //x=2.505 //y=1.655 //x2=2.26 //y2=1.405
cc_655 ( N_noxref_3_M1_noxref_d N_noxref_6_c_1306_n ) capacitor c=0.0138845f \
 //x=1.96 //y=0.905 //x2=2.26 //y2=1.405
cc_656 ( N_noxref_3_M1_noxref_d N_noxref_6_c_1308_n ) capacitor c=0.00132245f \
 //x=1.96 //y=0.905 //x2=2.415 //y2=0.905
cc_657 ( N_noxref_3_c_603_n N_noxref_6_c_1309_n ) capacitor c=0.00457401f \
 //x=2.505 //y=1.655 //x2=2.415 //y2=1.25
cc_658 ( N_noxref_3_M1_noxref_d N_noxref_6_c_1309_n ) capacitor c=0.00566463f \
 //x=1.96 //y=0.905 //x2=2.415 //y2=1.25
cc_659 ( N_noxref_3_c_604_n N_noxref_6_c_1311_n ) capacitor c=0.00877984f \
 //x=2.59 //y=2.59 //x2=1.85 //y2=2.08
cc_660 ( N_noxref_3_c_604_n N_noxref_6_c_1312_n ) capacitor c=0.00306024f \
 //x=2.59 //y=2.59 //x2=1.85 //y2=1.915
cc_661 ( N_noxref_3_M1_noxref_d N_noxref_6_c_1312_n ) capacitor c=0.00660593f \
 //x=1.96 //y=0.905 //x2=1.85 //y2=1.915
cc_662 ( N_noxref_3_c_632_n N_noxref_6_c_1314_n ) capacitor c=0.00346627f \
 //x=2.025 //y=5.2 //x2=1.88 //y2=4.7
cc_663 ( N_noxref_3_c_604_n N_noxref_6_c_1314_n ) capacitor c=0.00517969f \
 //x=2.59 //y=2.59 //x2=1.88 //y2=4.7
cc_664 ( N_noxref_3_M20_noxref_g N_noxref_6_M19_noxref_d ) capacitor \
 c=0.0180032f //x=5.08 //y=6.02 //x2=4.715 //y2=5.02
cc_665 ( N_noxref_3_c_607_n N_SN_c_1630_n ) capacitor c=0.00558344f //x=9.25 \
 //y=2.08 //x2=10.475 //y2=2.22
cc_666 ( N_noxref_3_c_622_n N_SN_c_1630_n ) capacitor c=0.00341397f //x=8.95 \
 //y=1.915 //x2=10.475 //y2=2.22
cc_667 ( N_noxref_3_c_597_n N_SN_c_1631_n ) capacitor c=0.00311593f //x=9.135 \
 //y=2.59 //x2=10.36 //y2=2.08
cc_668 ( N_noxref_3_c_607_n N_SN_c_1631_n ) capacitor c=0.0481863f //x=9.25 \
 //y=2.08 //x2=10.36 //y2=2.08
cc_669 ( N_noxref_3_c_622_n N_SN_c_1631_n ) capacitor c=0.00228225f //x=8.95 \
 //y=1.915 //x2=10.36 //y2=2.08
cc_670 ( N_noxref_3_c_675_p N_SN_c_1631_n ) capacitor c=0.00147352f //x=9.815 \
 //y=4.79 //x2=10.36 //y2=2.08
cc_671 ( N_noxref_3_c_659_n N_SN_c_1631_n ) capacitor c=0.00142741f //x=9.525 \
 //y=4.79 //x2=10.36 //y2=2.08
cc_672 ( N_noxref_3_M25_noxref_g N_SN_M27_noxref_g ) capacitor c=0.0105869f \
 //x=9.45 //y=6.02 //x2=10.33 //y2=6.02
cc_673 ( N_noxref_3_M26_noxref_g N_SN_M27_noxref_g ) capacitor c=0.10632f \
 //x=9.89 //y=6.02 //x2=10.33 //y2=6.02
cc_674 ( N_noxref_3_M26_noxref_g N_SN_M28_noxref_g ) capacitor c=0.0101598f \
 //x=9.89 //y=6.02 //x2=10.77 //y2=6.02
cc_675 ( N_noxref_3_c_618_n N_SN_c_1655_n ) capacitor c=5.72482e-19 //x=8.95 \
 //y=0.875 //x2=9.925 //y2=0.91
cc_676 ( N_noxref_3_c_620_n N_SN_c_1655_n ) capacitor c=0.00149976f //x=8.95 \
 //y=1.22 //x2=9.925 //y2=0.91
cc_677 ( N_noxref_3_c_625_n N_SN_c_1655_n ) capacitor c=0.0160123f //x=9.48 \
 //y=0.875 //x2=9.925 //y2=0.91
cc_678 ( N_noxref_3_c_621_n N_SN_c_1658_n ) capacitor c=0.00111227f //x=8.95 \
 //y=1.53 //x2=9.925 //y2=1.22
cc_679 ( N_noxref_3_c_627_n N_SN_c_1658_n ) capacitor c=0.0124075f //x=9.48 \
 //y=1.22 //x2=9.925 //y2=1.22
cc_680 ( N_noxref_3_c_625_n N_SN_c_1660_n ) capacitor c=0.00103227f //x=9.48 \
 //y=0.875 //x2=10.45 //y2=0.91
cc_681 ( N_noxref_3_c_627_n N_SN_c_1661_n ) capacitor c=0.0010154f //x=9.48 \
 //y=1.22 //x2=10.45 //y2=1.22
cc_682 ( N_noxref_3_c_627_n N_SN_c_1662_n ) capacitor c=9.23422e-19 //x=9.48 \
 //y=1.22 //x2=10.45 //y2=1.45
cc_683 ( N_noxref_3_c_607_n N_SN_c_1663_n ) capacitor c=0.00211714f //x=9.25 \
 //y=2.08 //x2=10.45 //y2=1.915
cc_684 ( N_noxref_3_c_622_n N_SN_c_1663_n ) capacitor c=0.00909574f //x=8.95 \
 //y=1.915 //x2=10.45 //y2=1.915
cc_685 ( N_noxref_3_c_607_n N_SN_c_1665_n ) capacitor c=0.00183762f //x=9.25 \
 //y=2.08 //x2=10.36 //y2=4.7
cc_686 ( N_noxref_3_c_675_p N_SN_c_1665_n ) capacitor c=0.0168581f //x=9.815 \
 //y=4.79 //x2=10.36 //y2=4.7
cc_687 ( N_noxref_3_c_659_n N_SN_c_1665_n ) capacitor c=0.00484466f //x=9.525 \
 //y=4.79 //x2=10.36 //y2=4.7
cc_688 ( N_noxref_3_c_597_n N_noxref_9_c_1846_n ) capacitor c=0.0761096f \
 //x=9.135 //y=2.59 //x2=11.355 //y2=3.7
cc_689 ( N_noxref_3_c_607_n N_noxref_9_c_1846_n ) capacitor c=0.0237114f \
 //x=9.25 //y=2.08 //x2=11.355 //y2=3.7
cc_690 ( N_noxref_3_c_597_n N_noxref_9_c_1902_n ) capacitor c=0.00777466f \
 //x=9.135 //y=2.59 //x2=6.775 //y2=3.7
cc_691 ( N_noxref_3_c_597_n N_noxref_9_c_1850_n ) capacitor c=0.025454f \
 //x=9.135 //y=2.59 //x2=6.66 //y2=2.08
cc_692 ( N_noxref_3_c_606_n N_noxref_9_c_1850_n ) capacitor c=0.00150385f \
 //x=4.44 //y=2.08 //x2=6.66 //y2=2.08
cc_693 ( N_noxref_3_c_607_n N_noxref_9_c_1850_n ) capacitor c=8.19041e-19 \
 //x=9.25 //y=2.08 //x2=6.66 //y2=2.08
cc_694 ( N_noxref_3_c_607_n N_noxref_9_c_1851_n ) capacitor c=0.00128526f \
 //x=9.25 //y=2.08 //x2=11.47 //y2=2.08
cc_695 ( N_noxref_3_c_597_n N_noxref_9_c_1907_n ) capacitor c=0.00232725f \
 //x=9.135 //y=2.59 //x2=6.66 //y2=2.08
cc_696 ( N_noxref_3_c_636_n N_D_c_2340_n ) capacitor c=0.00569255f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=2.08
cc_697 ( N_noxref_3_c_604_n N_D_c_2340_n ) capacitor c=0.0042593f //x=2.59 \
 //y=2.59 //x2=1.11 //y2=2.08
cc_698 ( N_noxref_3_c_636_n N_D_M15_noxref_g ) capacitor c=0.0177326f \
 //x=1.315 //y=5.2 //x2=1.01 //y2=6.02
cc_699 ( N_noxref_3_c_632_n N_D_M16_noxref_g ) capacitor c=0.0203837f \
 //x=2.025 //y=5.2 //x2=1.45 //y2=6.02
cc_700 ( N_noxref_3_M15_noxref_d N_D_M16_noxref_g ) capacitor c=0.0173476f \
 //x=1.085 //y=5.02 //x2=1.45 //y2=6.02
cc_701 ( N_noxref_3_c_636_n N_D_c_2358_n ) capacitor c=0.00571434f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=4.7
cc_702 ( N_noxref_3_c_710_p N_noxref_12_c_2416_n ) capacitor c=3.15806e-19 \
 //x=2.235 //y=1.655 //x2=0.695 //y2=1.495
cc_703 ( N_noxref_3_c_710_p N_noxref_12_c_2404_n ) capacitor c=0.0201674f \
 //x=2.235 //y=1.655 //x2=1.665 //y2=1.495
cc_704 ( N_noxref_3_c_603_n N_noxref_12_c_2405_n ) capacitor c=0.00467467f \
 //x=2.505 //y=1.655 //x2=2.55 //y2=0.53
cc_705 ( N_noxref_3_M1_noxref_d N_noxref_12_c_2405_n ) capacitor c=0.0118355f \
 //x=1.96 //y=0.905 //x2=2.55 //y2=0.53
cc_706 ( N_noxref_3_c_591_n N_noxref_12_M0_noxref_s ) capacitor c=2.68031e-19 \
 //x=4.295 //y=2.59 //x2=0.56 //y2=0.365
cc_707 ( N_noxref_3_c_595_n N_noxref_12_M0_noxref_s ) capacitor c=5.97427e-19 \
 //x=2.705 //y=2.59 //x2=0.56 //y2=0.365
cc_708 ( N_noxref_3_c_603_n N_noxref_12_M0_noxref_s ) capacitor c=0.0129465f \
 //x=2.505 //y=1.655 //x2=0.56 //y2=0.365
cc_709 ( N_noxref_3_M1_noxref_d N_noxref_12_M0_noxref_s ) capacitor \
 c=0.0437911f //x=1.96 //y=0.905 //x2=0.56 //y2=0.365
cc_710 ( N_noxref_3_c_591_n N_noxref_13_c_2461_n ) capacitor c=0.00448771f \
 //x=4.295 //y=2.59 //x2=3.92 //y2=1.505
cc_711 ( N_noxref_3_c_603_n N_noxref_13_c_2461_n ) capacitor c=4.08644e-19 \
 //x=2.505 //y=1.655 //x2=3.92 //y2=1.505
cc_712 ( N_noxref_3_c_612_n N_noxref_13_c_2461_n ) capacitor c=0.0034165f \
 //x=4.14 //y=1.915 //x2=3.92 //y2=1.505
cc_713 ( N_noxref_3_c_591_n N_noxref_13_c_2445_n ) capacitor c=0.00818794f \
 //x=4.295 //y=2.59 //x2=4.805 //y2=1.59
cc_714 ( N_noxref_3_c_597_n N_noxref_13_c_2445_n ) capacitor c=0.00225113f \
 //x=9.135 //y=2.59 //x2=4.805 //y2=1.59
cc_715 ( N_noxref_3_c_601_n N_noxref_13_c_2445_n ) capacitor c=0.00603529f \
 //x=4.705 //y=2.59 //x2=4.805 //y2=1.59
cc_716 ( N_noxref_3_c_606_n N_noxref_13_c_2445_n ) capacitor c=0.0117784f \
 //x=4.44 //y=2.08 //x2=4.805 //y2=1.59
cc_717 ( N_noxref_3_c_611_n N_noxref_13_c_2445_n ) capacitor c=0.00703864f \
 //x=4.14 //y=1.53 //x2=4.805 //y2=1.59
cc_718 ( N_noxref_3_c_612_n N_noxref_13_c_2445_n ) capacitor c=0.0215834f \
 //x=4.14 //y=1.915 //x2=4.805 //y2=1.59
cc_719 ( N_noxref_3_c_614_n N_noxref_13_c_2445_n ) capacitor c=0.00708583f \
 //x=4.515 //y=1.375 //x2=4.805 //y2=1.59
cc_720 ( N_noxref_3_c_617_n N_noxref_13_c_2445_n ) capacitor c=0.00698822f \
 //x=4.67 //y=1.22 //x2=4.805 //y2=1.59
cc_721 ( N_noxref_3_c_597_n N_noxref_13_c_2472_n ) capacitor c=0.0144126f \
 //x=9.135 //y=2.59 //x2=5.775 //y2=1.59
cc_722 ( N_noxref_3_c_597_n N_noxref_13_M2_noxref_s ) capacitor c=0.00867201f \
 //x=9.135 //y=2.59 //x2=3.785 //y2=0.375
cc_723 ( N_noxref_3_c_608_n N_noxref_13_M2_noxref_s ) capacitor c=0.0327271f \
 //x=4.14 //y=0.875 //x2=3.785 //y2=0.375
cc_724 ( N_noxref_3_c_611_n N_noxref_13_M2_noxref_s ) capacitor c=7.99997e-19 \
 //x=4.14 //y=1.53 //x2=3.785 //y2=0.375
cc_725 ( N_noxref_3_c_612_n N_noxref_13_M2_noxref_s ) capacitor c=0.00122123f \
 //x=4.14 //y=1.915 //x2=3.785 //y2=0.375
cc_726 ( N_noxref_3_c_615_n N_noxref_13_M2_noxref_s ) capacitor c=0.0121427f \
 //x=4.67 //y=0.875 //x2=3.785 //y2=0.375
cc_727 ( N_noxref_3_M1_noxref_d N_noxref_13_M2_noxref_s ) capacitor \
 c=2.53688e-19 //x=1.96 //y=0.905 //x2=3.785 //y2=0.375
cc_728 ( N_noxref_3_c_597_n N_noxref_14_c_2497_n ) capacitor c=0.00494691f \
 //x=9.135 //y=2.59 //x2=6.345 //y2=0.995
cc_729 ( N_noxref_3_c_597_n N_noxref_14_c_2502_n ) capacitor c=8.29806e-19 \
 //x=9.135 //y=2.59 //x2=7.315 //y2=0.54
cc_730 ( N_noxref_3_c_597_n N_noxref_14_M4_noxref_s ) capacitor c=0.00448771f \
 //x=9.135 //y=2.59 //x2=6.295 //y2=0.375
cc_731 ( N_noxref_3_c_597_n N_noxref_15_c_2566_n ) capacitor c=0.00448771f \
 //x=9.135 //y=2.59 //x2=8.73 //y2=1.505
cc_732 ( N_noxref_3_c_622_n N_noxref_15_c_2566_n ) capacitor c=0.0034165f \
 //x=8.95 //y=1.915 //x2=8.73 //y2=1.505
cc_733 ( N_noxref_3_c_597_n N_noxref_15_c_2550_n ) capacitor c=0.0116291f \
 //x=9.135 //y=2.59 //x2=9.615 //y2=1.59
cc_734 ( N_noxref_3_c_607_n N_noxref_15_c_2550_n ) capacitor c=0.0122435f \
 //x=9.25 //y=2.08 //x2=9.615 //y2=1.59
cc_735 ( N_noxref_3_c_621_n N_noxref_15_c_2550_n ) capacitor c=0.00703864f \
 //x=8.95 //y=1.53 //x2=9.615 //y2=1.59
cc_736 ( N_noxref_3_c_622_n N_noxref_15_c_2550_n ) capacitor c=0.0215834f \
 //x=8.95 //y=1.915 //x2=9.615 //y2=1.59
cc_737 ( N_noxref_3_c_624_n N_noxref_15_c_2550_n ) capacitor c=0.00708583f \
 //x=9.325 //y=1.375 //x2=9.615 //y2=1.59
cc_738 ( N_noxref_3_c_627_n N_noxref_15_c_2550_n ) capacitor c=0.00698822f \
 //x=9.48 //y=1.22 //x2=9.615 //y2=1.59
cc_739 ( N_noxref_3_c_618_n N_noxref_15_M5_noxref_s ) capacitor c=0.0327271f \
 //x=8.95 //y=0.875 //x2=8.595 //y2=0.375
cc_740 ( N_noxref_3_c_621_n N_noxref_15_M5_noxref_s ) capacitor c=7.99997e-19 \
 //x=8.95 //y=1.53 //x2=8.595 //y2=0.375
cc_741 ( N_noxref_3_c_622_n N_noxref_15_M5_noxref_s ) capacitor c=0.00122123f \
 //x=8.95 //y=1.915 //x2=8.595 //y2=0.375
cc_742 ( N_noxref_3_c_625_n N_noxref_15_M5_noxref_s ) capacitor c=0.0121427f \
 //x=9.48 //y=0.875 //x2=8.595 //y2=0.375
cc_743 ( N_noxref_4_c_847_n N_CLK_c_994_n ) capacitor c=0.032141f //x=10.465 \
 //y=5.155 //x2=14.685 //y2=4.44
cc_744 ( N_noxref_4_c_851_n N_CLK_c_994_n ) capacitor c=0.0230136f //x=9.755 \
 //y=5.155 //x2=14.685 //y2=4.44
cc_745 ( N_noxref_4_c_857_n N_CLK_c_994_n ) capacitor c=0.0183122f //x=12.125 \
 //y=5.155 //x2=14.685 //y2=4.44
cc_746 ( N_noxref_4_c_834_n N_CLK_c_994_n ) capacitor c=0.0210274f //x=12.21 \
 //y=2.59 //x2=14.685 //y2=4.44
cc_747 ( N_noxref_4_c_835_n N_CLK_c_994_n ) capacitor c=0.0215137f //x=14.06 \
 //y=2.08 //x2=14.685 //y2=4.44
cc_748 ( N_noxref_4_c_869_n N_CLK_c_994_n ) capacitor c=0.0109968f //x=14.06 \
 //y=4.7 //x2=14.685 //y2=4.44
cc_749 ( N_noxref_4_c_835_n N_CLK_c_1054_n ) capacitor c=0.00400249f //x=14.06 \
 //y=2.08 //x2=14.8 //y2=4.535
cc_750 ( N_noxref_4_c_869_n N_CLK_c_1054_n ) capacitor c=0.00415951f //x=14.06 \
 //y=4.7 //x2=14.8 //y2=4.535
cc_751 ( N_noxref_4_c_831_n N_CLK_c_992_n ) capacitor c=0.00720056f //x=13.945 \
 //y=2.59 //x2=14.8 //y2=2.08
cc_752 ( N_noxref_4_c_834_n N_CLK_c_992_n ) capacitor c=8.83058e-19 //x=12.21 \
 //y=2.59 //x2=14.8 //y2=2.08
cc_753 ( N_noxref_4_c_835_n N_CLK_c_992_n ) capacitor c=0.0762889f //x=14.06 \
 //y=2.08 //x2=14.8 //y2=2.08
cc_754 ( N_noxref_4_c_840_n N_CLK_c_992_n ) capacitor c=0.00284029f //x=13.865 \
 //y=1.915 //x2=14.8 //y2=2.08
cc_755 ( N_noxref_4_M31_noxref_g N_CLK_M33_noxref_g ) capacitor c=0.0104611f \
 //x=13.96 //y=6.02 //x2=14.84 //y2=6.02
cc_756 ( N_noxref_4_M32_noxref_g N_CLK_M33_noxref_g ) capacitor c=0.106811f \
 //x=14.4 //y=6.02 //x2=14.84 //y2=6.02
cc_757 ( N_noxref_4_M32_noxref_g N_CLK_M34_noxref_g ) capacitor c=0.0100341f \
 //x=14.4 //y=6.02 //x2=15.28 //y2=6.02
cc_758 ( N_noxref_4_c_836_n N_CLK_c_1063_n ) capacitor c=4.86506e-19 \
 //x=13.865 //y=0.865 //x2=14.835 //y2=0.905
cc_759 ( N_noxref_4_c_838_n N_CLK_c_1063_n ) capacitor c=0.00152104f \
 //x=13.865 //y=1.21 //x2=14.835 //y2=0.905
cc_760 ( N_noxref_4_c_843_n N_CLK_c_1063_n ) capacitor c=0.0151475f //x=14.395 \
 //y=0.865 //x2=14.835 //y2=0.905
cc_761 ( N_noxref_4_c_839_n N_CLK_c_1066_n ) capacitor c=0.00109982f \
 //x=13.865 //y=1.52 //x2=14.835 //y2=1.25
cc_762 ( N_noxref_4_c_845_n N_CLK_c_1066_n ) capacitor c=0.0111064f //x=14.395 \
 //y=1.21 //x2=14.835 //y2=1.25
cc_763 ( N_noxref_4_c_839_n N_CLK_c_1068_n ) capacitor c=9.57794e-19 \
 //x=13.865 //y=1.52 //x2=14.835 //y2=1.56
cc_764 ( N_noxref_4_c_840_n N_CLK_c_1068_n ) capacitor c=0.00662747f \
 //x=13.865 //y=1.915 //x2=14.835 //y2=1.56
cc_765 ( N_noxref_4_c_845_n N_CLK_c_1068_n ) capacitor c=0.00862358f \
 //x=14.395 //y=1.21 //x2=14.835 //y2=1.56
cc_766 ( N_noxref_4_c_843_n N_CLK_c_1071_n ) capacitor c=0.00124821f \
 //x=14.395 //y=0.865 //x2=15.365 //y2=0.905
cc_767 ( N_noxref_4_c_845_n N_CLK_c_1072_n ) capacitor c=0.00200715f \
 //x=14.395 //y=1.21 //x2=15.365 //y2=1.25
cc_768 ( N_noxref_4_c_835_n N_CLK_c_1073_n ) capacitor c=0.00282278f //x=14.06 \
 //y=2.08 //x2=14.8 //y2=2.08
cc_769 ( N_noxref_4_c_840_n N_CLK_c_1073_n ) capacitor c=0.0172771f //x=13.865 \
 //y=1.915 //x2=14.8 //y2=2.08
cc_770 ( N_noxref_4_c_835_n N_CLK_c_1075_n ) capacitor c=0.00342116f //x=14.06 \
 //y=2.08 //x2=14.83 //y2=4.7
cc_771 ( N_noxref_4_c_869_n N_CLK_c_1075_n ) capacitor c=0.0292158f //x=14.06 \
 //y=4.7 //x2=14.83 //y2=4.7
cc_772 ( N_noxref_4_c_831_n N_noxref_6_c_1215_n ) capacitor c=0.00628974f \
 //x=13.945 //y=2.59 //x2=17.275 //y2=4.07
cc_773 ( N_noxref_4_c_832_n N_noxref_6_c_1215_n ) capacitor c=5.0661e-19 \
 //x=12.325 //y=2.59 //x2=17.275 //y2=4.07
cc_774 ( N_noxref_4_c_834_n N_noxref_6_c_1215_n ) capacitor c=0.0181982f \
 //x=12.21 //y=2.59 //x2=17.275 //y2=4.07
cc_775 ( N_noxref_4_c_835_n N_noxref_6_c_1215_n ) capacitor c=0.0184765f \
 //x=14.06 //y=2.08 //x2=17.275 //y2=4.07
cc_776 ( N_noxref_4_c_851_n N_noxref_6_c_1237_n ) capacitor c=3.10026e-19 \
 //x=9.755 //y=5.155 //x2=7.315 //y2=5.155
cc_777 ( N_noxref_4_c_831_n N_SN_c_1620_n ) capacitor c=0.172308f //x=13.945 \
 //y=2.59 //x2=21.715 //y2=2.22
cc_778 ( N_noxref_4_c_832_n N_SN_c_1620_n ) capacitor c=0.0291301f //x=12.325 \
 //y=2.59 //x2=21.715 //y2=2.22
cc_779 ( N_noxref_4_c_926_p N_SN_c_1620_n ) capacitor c=0.016327f //x=11.81 \
 //y=1.665 //x2=21.715 //y2=2.22
cc_780 ( N_noxref_4_c_834_n N_SN_c_1620_n ) capacitor c=0.0215653f //x=12.21 \
 //y=2.59 //x2=21.715 //y2=2.22
cc_781 ( N_noxref_4_c_835_n N_SN_c_1620_n ) capacitor c=0.0203358f //x=14.06 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_782 ( N_noxref_4_c_840_n N_SN_c_1620_n ) capacitor c=0.00894156f //x=13.865 \
 //y=1.915 //x2=21.715 //y2=2.22
cc_783 ( N_noxref_4_c_847_n N_SN_c_1631_n ) capacitor c=0.0144268f //x=10.465 \
 //y=5.155 //x2=10.36 //y2=2.08
cc_784 ( N_noxref_4_c_834_n N_SN_c_1631_n ) capacitor c=0.00268713f //x=12.21 \
 //y=2.59 //x2=10.36 //y2=2.08
cc_785 ( N_noxref_4_c_847_n N_SN_M27_noxref_g ) capacitor c=0.0165266f \
 //x=10.465 //y=5.155 //x2=10.33 //y2=6.02
cc_786 ( N_noxref_4_M27_noxref_d N_SN_M27_noxref_g ) capacitor c=0.0180032f \
 //x=10.405 //y=5.02 //x2=10.33 //y2=6.02
cc_787 ( N_noxref_4_c_853_n N_SN_M28_noxref_g ) capacitor c=0.01736f \
 //x=11.345 //y=5.155 //x2=10.77 //y2=6.02
cc_788 ( N_noxref_4_M27_noxref_d N_SN_M28_noxref_g ) capacitor c=0.0180032f \
 //x=10.405 //y=5.02 //x2=10.77 //y2=6.02
cc_789 ( N_noxref_4_c_936_p N_SN_c_1680_n ) capacitor c=0.00426767f //x=10.55 \
 //y=5.155 //x2=10.695 //y2=4.79
cc_790 ( N_noxref_4_c_847_n N_SN_c_1665_n ) capacitor c=0.00322054f //x=10.465 \
 //y=5.155 //x2=10.36 //y2=4.7
cc_791 ( N_noxref_4_c_831_n N_noxref_9_c_1848_n ) capacitor c=0.0565623f \
 //x=13.945 //y=2.59 //x2=15.425 //y2=3.7
cc_792 ( N_noxref_4_c_832_n N_noxref_9_c_1848_n ) capacitor c=0.00783891f \
 //x=12.325 //y=2.59 //x2=15.425 //y2=3.7
cc_793 ( N_noxref_4_c_834_n N_noxref_9_c_1848_n ) capacitor c=0.0227211f \
 //x=12.21 //y=2.59 //x2=15.425 //y2=3.7
cc_794 ( N_noxref_4_c_835_n N_noxref_9_c_1848_n ) capacitor c=0.0226973f \
 //x=14.06 //y=2.08 //x2=15.425 //y2=3.7
cc_795 ( N_noxref_4_c_834_n N_noxref_9_c_1912_n ) capacitor c=0.00117715f \
 //x=12.21 //y=2.59 //x2=11.585 //y2=3.7
cc_796 ( N_noxref_4_c_832_n N_noxref_9_c_1851_n ) capacitor c=0.00456439f \
 //x=12.325 //y=2.59 //x2=11.47 //y2=2.08
cc_797 ( N_noxref_4_c_834_n N_noxref_9_c_1851_n ) capacitor c=0.081931f \
 //x=12.21 //y=2.59 //x2=11.47 //y2=2.08
cc_798 ( N_noxref_4_c_835_n N_noxref_9_c_1851_n ) capacitor c=7.74334e-19 \
 //x=14.06 //y=2.08 //x2=11.47 //y2=2.08
cc_799 ( N_noxref_4_c_946_p N_noxref_9_c_1851_n ) capacitor c=0.016476f \
 //x=11.43 //y=5.155 //x2=11.47 //y2=2.08
cc_800 ( N_noxref_4_M32_noxref_g N_noxref_9_c_1864_n ) capacitor c=0.0169521f \
 //x=14.4 //y=6.02 //x2=14.975 //y2=5.2
cc_801 ( N_noxref_4_c_835_n N_noxref_9_c_1868_n ) capacitor c=0.00539951f \
 //x=14.06 //y=2.08 //x2=14.265 //y2=5.2
cc_802 ( N_noxref_4_M31_noxref_g N_noxref_9_c_1868_n ) capacitor c=0.0177326f \
 //x=13.96 //y=6.02 //x2=14.265 //y2=5.2
cc_803 ( N_noxref_4_c_869_n N_noxref_9_c_1868_n ) capacitor c=0.00581252f \
 //x=14.06 //y=4.7 //x2=14.265 //y2=5.2
cc_804 ( N_noxref_4_c_834_n N_noxref_9_c_1853_n ) capacitor c=3.52729e-19 \
 //x=12.21 //y=2.59 //x2=15.54 //y2=3.7
cc_805 ( N_noxref_4_c_835_n N_noxref_9_c_1853_n ) capacitor c=0.00363124f \
 //x=14.06 //y=2.08 //x2=15.54 //y2=3.7
cc_806 ( N_noxref_4_c_853_n N_noxref_9_M29_noxref_g ) capacitor c=0.01736f \
 //x=11.345 //y=5.155 //x2=11.21 //y2=6.02
cc_807 ( N_noxref_4_M29_noxref_d N_noxref_9_M29_noxref_g ) capacitor \
 c=0.0180032f //x=11.285 //y=5.02 //x2=11.21 //y2=6.02
cc_808 ( N_noxref_4_c_857_n N_noxref_9_M30_noxref_g ) capacitor c=0.0194981f \
 //x=12.125 //y=5.155 //x2=11.65 //y2=6.02
cc_809 ( N_noxref_4_M29_noxref_d N_noxref_9_M30_noxref_g ) capacitor \
 c=0.0194246f //x=11.285 //y=5.02 //x2=11.65 //y2=6.02
cc_810 ( N_noxref_4_M7_noxref_d N_noxref_9_c_1927_n ) capacitor c=0.00217566f \
 //x=11.535 //y=0.915 //x2=11.46 //y2=0.915
cc_811 ( N_noxref_4_M7_noxref_d N_noxref_9_c_1928_n ) capacitor c=0.0034598f \
 //x=11.535 //y=0.915 //x2=11.46 //y2=1.26
cc_812 ( N_noxref_4_M7_noxref_d N_noxref_9_c_1929_n ) capacitor c=0.00546784f \
 //x=11.535 //y=0.915 //x2=11.46 //y2=1.57
cc_813 ( N_noxref_4_M7_noxref_d N_noxref_9_c_1930_n ) capacitor c=0.00241102f \
 //x=11.535 //y=0.915 //x2=11.835 //y2=0.76
cc_814 ( N_noxref_4_c_833_n N_noxref_9_c_1931_n ) capacitor c=0.00371277f \
 //x=12.125 //y=1.665 //x2=11.835 //y2=1.415
cc_815 ( N_noxref_4_M7_noxref_d N_noxref_9_c_1931_n ) capacitor c=0.0138621f \
 //x=11.535 //y=0.915 //x2=11.835 //y2=1.415
cc_816 ( N_noxref_4_M7_noxref_d N_noxref_9_c_1933_n ) capacitor c=0.00219619f \
 //x=11.535 //y=0.915 //x2=11.99 //y2=0.915
cc_817 ( N_noxref_4_c_833_n N_noxref_9_c_1934_n ) capacitor c=0.00457401f \
 //x=12.125 //y=1.665 //x2=11.99 //y2=1.26
cc_818 ( N_noxref_4_M7_noxref_d N_noxref_9_c_1934_n ) capacitor c=0.00603828f \
 //x=11.535 //y=0.915 //x2=11.99 //y2=1.26
cc_819 ( N_noxref_4_c_834_n N_noxref_9_c_1936_n ) capacitor c=0.00709342f \
 //x=12.21 //y=2.59 //x2=11.47 //y2=2.08
cc_820 ( N_noxref_4_c_834_n N_noxref_9_c_1937_n ) capacitor c=0.00283672f \
 //x=12.21 //y=2.59 //x2=11.47 //y2=1.915
cc_821 ( N_noxref_4_M7_noxref_d N_noxref_9_c_1937_n ) capacitor c=0.00661782f \
 //x=11.535 //y=0.915 //x2=11.47 //y2=1.915
cc_822 ( N_noxref_4_c_857_n N_noxref_9_c_1939_n ) capacitor c=0.00201851f \
 //x=12.125 //y=5.155 //x2=11.47 //y2=4.7
cc_823 ( N_noxref_4_c_834_n N_noxref_9_c_1939_n ) capacitor c=0.013693f \
 //x=12.21 //y=2.59 //x2=11.47 //y2=4.7
cc_824 ( N_noxref_4_c_946_p N_noxref_9_c_1939_n ) capacitor c=0.00475601f \
 //x=11.43 //y=5.155 //x2=11.47 //y2=4.7
cc_825 ( N_noxref_4_M32_noxref_g N_noxref_9_M31_noxref_d ) capacitor \
 c=0.0173476f //x=14.4 //y=6.02 //x2=14.035 //y2=5.02
cc_826 ( N_noxref_4_M7_noxref_d N_noxref_15_M5_noxref_s ) capacitor \
 c=0.00309936f //x=11.535 //y=0.915 //x2=8.595 //y2=0.375
cc_827 ( N_noxref_4_c_833_n N_noxref_16_c_2609_n ) capacitor c=0.00457167f \
 //x=12.125 //y=1.665 //x2=12.125 //y2=0.54
cc_828 ( N_noxref_4_M7_noxref_d N_noxref_16_c_2609_n ) capacitor c=0.0115903f \
 //x=11.535 //y=0.915 //x2=12.125 //y2=0.54
cc_829 ( N_noxref_4_c_926_p N_noxref_16_c_2620_n ) capacitor c=0.020048f \
 //x=11.81 //y=1.665 //x2=11.24 //y2=0.995
cc_830 ( N_noxref_4_M7_noxref_d N_noxref_16_M6_noxref_d ) capacitor \
 c=5.27807e-19 //x=11.535 //y=0.915 //x2=10 //y2=0.91
cc_831 ( N_noxref_4_c_833_n N_noxref_16_M7_noxref_s ) capacitor c=0.0184051f \
 //x=12.125 //y=1.665 //x2=11.105 //y2=0.375
cc_832 ( N_noxref_4_M7_noxref_d N_noxref_16_M7_noxref_s ) capacitor \
 c=0.0426444f //x=11.535 //y=0.915 //x2=11.105 //y2=0.375
cc_833 ( N_noxref_4_c_833_n N_noxref_17_c_2676_n ) capacitor c=3.04182e-19 \
 //x=12.125 //y=1.665 //x2=13.645 //y2=1.495
cc_834 ( N_noxref_4_c_840_n N_noxref_17_c_2676_n ) capacitor c=0.0034165f \
 //x=13.865 //y=1.915 //x2=13.645 //y2=1.495
cc_835 ( N_noxref_4_c_835_n N_noxref_17_c_2657_n ) capacitor c=0.011618f \
 //x=14.06 //y=2.08 //x2=14.53 //y2=1.58
cc_836 ( N_noxref_4_c_839_n N_noxref_17_c_2657_n ) capacitor c=0.00696403f \
 //x=13.865 //y=1.52 //x2=14.53 //y2=1.58
cc_837 ( N_noxref_4_c_840_n N_noxref_17_c_2657_n ) capacitor c=0.0174694f \
 //x=13.865 //y=1.915 //x2=14.53 //y2=1.58
cc_838 ( N_noxref_4_c_842_n N_noxref_17_c_2657_n ) capacitor c=0.00776811f \
 //x=14.24 //y=1.365 //x2=14.53 //y2=1.58
cc_839 ( N_noxref_4_c_845_n N_noxref_17_c_2657_n ) capacitor c=0.00339872f \
 //x=14.395 //y=1.21 //x2=14.53 //y2=1.58
cc_840 ( N_noxref_4_c_840_n N_noxref_17_c_2664_n ) capacitor c=6.71402e-19 \
 //x=13.865 //y=1.915 //x2=14.615 //y2=1.495
cc_841 ( N_noxref_4_c_836_n N_noxref_17_M8_noxref_s ) capacitor c=0.0327502f \
 //x=13.865 //y=0.865 //x2=13.51 //y2=0.365
cc_842 ( N_noxref_4_c_839_n N_noxref_17_M8_noxref_s ) capacitor c=3.48408e-19 \
 //x=13.865 //y=1.52 //x2=13.51 //y2=0.365
cc_843 ( N_noxref_4_c_843_n N_noxref_17_M8_noxref_s ) capacitor c=0.0120759f \
 //x=14.395 //y=0.865 //x2=13.51 //y2=0.365
cc_844 ( N_CLK_c_994_n N_noxref_6_c_1189_n ) capacitor c=0.139602f //x=14.685 \
 //y=4.44 //x2=7.28 //y2=4.07
cc_845 ( N_CLK_c_1005_n N_noxref_6_c_1189_n ) capacitor c=0.0291328f //x=5.665 \
 //y=4.44 //x2=7.28 //y2=4.07
cc_846 ( N_CLK_c_991_n N_noxref_6_c_1189_n ) capacitor c=0.0256971f //x=5.55 \
 //y=2.08 //x2=7.28 //y2=4.07
cc_847 ( N_CLK_c_994_n N_noxref_6_c_1215_n ) capacitor c=0.654862f //x=14.685 \
 //y=4.44 //x2=17.275 //y2=4.07
cc_848 ( N_CLK_c_992_n N_noxref_6_c_1215_n ) capacitor c=0.0187718f //x=14.8 \
 //y=2.08 //x2=17.275 //y2=4.07
cc_849 ( N_CLK_c_1082_p N_noxref_6_c_1215_n ) capacitor c=0.00756255f \
 //x=15.205 //y=4.79 //x2=17.275 //y2=4.07
cc_850 ( N_CLK_c_1075_n N_noxref_6_c_1215_n ) capacitor c=4.6185e-19 //x=14.83 \
 //y=4.7 //x2=17.275 //y2=4.07
cc_851 ( N_CLK_c_994_n N_noxref_6_c_1224_n ) capacitor c=0.0265302f //x=14.685 \
 //y=4.44 //x2=7.51 //y2=4.07
cc_852 ( N_CLK_c_1005_n N_noxref_6_c_1227_n ) capacitor c=0.00330099f \
 //x=5.665 //y=4.44 //x2=5.655 //y2=5.155
cc_853 ( N_CLK_c_991_n N_noxref_6_c_1227_n ) capacitor c=0.014564f //x=5.55 \
 //y=2.08 //x2=5.655 //y2=5.155
cc_854 ( N_CLK_M21_noxref_g N_noxref_6_c_1227_n ) capacitor c=0.016514f \
 //x=5.52 //y=6.02 //x2=5.655 //y2=5.155
cc_855 ( N_CLK_c_1045_n N_noxref_6_c_1227_n ) capacitor c=0.00322046f //x=5.55 \
 //y=4.7 //x2=5.655 //y2=5.155
cc_856 ( N_CLK_M22_noxref_g N_noxref_6_c_1233_n ) capacitor c=0.01736f \
 //x=5.96 //y=6.02 //x2=6.535 //y2=5.155
cc_857 ( N_CLK_c_994_n N_noxref_6_c_1237_n ) capacitor c=0.0182691f //x=14.685 \
 //y=4.44 //x2=7.315 //y2=5.155
cc_858 ( N_CLK_c_994_n N_noxref_6_c_1336_n ) capacitor c=0.0207896f //x=14.685 \
 //y=4.44 //x2=7.4 //y2=5.07
cc_859 ( N_CLK_c_991_n N_noxref_6_c_1336_n ) capacitor c=7.17254e-19 //x=5.55 \
 //y=2.08 //x2=7.4 //y2=5.07
cc_860 ( N_CLK_c_992_n N_noxref_6_c_1195_n ) capacitor c=0.00117524f //x=14.8 \
 //y=2.08 //x2=17.39 //y2=2.08
cc_861 ( N_CLK_c_994_n N_noxref_6_c_1339_n ) capacitor c=0.0311227f //x=14.685 \
 //y=4.44 //x2=5.74 //y2=5.155
cc_862 ( N_CLK_c_1095_p N_noxref_6_c_1339_n ) capacitor c=0.00426767f \
 //x=5.885 //y=4.79 //x2=5.74 //y2=5.155
cc_863 ( N_CLK_c_994_n N_noxref_6_c_1244_n ) capacitor c=0.00215288f \
 //x=14.685 //y=4.44 //x2=7.395 //y2=4.07
cc_864 ( N_CLK_c_991_n N_noxref_6_c_1294_n ) capacitor c=0.00212483f //x=5.55 \
 //y=2.08 //x2=7.397 //y2=3.905
cc_865 ( N_CLK_M21_noxref_g N_noxref_6_M21_noxref_d ) capacitor c=0.0180032f \
 //x=5.52 //y=6.02 //x2=5.595 //y2=5.02
cc_866 ( N_CLK_M22_noxref_g N_noxref_6_M21_noxref_d ) capacitor c=0.0180032f \
 //x=5.96 //y=6.02 //x2=5.595 //y2=5.02
cc_867 ( N_CLK_c_992_n N_SN_c_1620_n ) capacitor c=0.0226984f //x=14.8 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_868 ( N_CLK_c_1101_p N_SN_c_1620_n ) capacitor c=3.11115e-19 //x=15.21 \
 //y=1.405 //x2=21.715 //y2=2.22
cc_869 ( N_CLK_c_1073_n N_SN_c_1620_n ) capacitor c=0.00569088f //x=14.8 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_870 ( N_CLK_c_994_n N_SN_c_1631_n ) capacitor c=0.0210462f //x=14.685 \
 //y=4.44 //x2=10.36 //y2=2.08
cc_871 ( N_CLK_c_994_n N_SN_c_1680_n ) capacitor c=0.0085986f //x=14.685 \
 //y=4.44 //x2=10.695 //y2=4.79
cc_872 ( N_CLK_c_994_n N_SN_c_1665_n ) capacitor c=0.00293313f //x=14.685 \
 //y=4.44 //x2=10.36 //y2=4.7
cc_873 ( N_CLK_c_994_n N_noxref_9_c_1846_n ) capacitor c=0.0345106f //x=14.685 \
 //y=4.44 //x2=11.355 //y2=3.7
cc_874 ( N_CLK_c_994_n N_noxref_9_c_1902_n ) capacitor c=7.0371e-19 //x=14.685 \
 //y=4.44 //x2=6.775 //y2=3.7
cc_875 ( N_CLK_c_991_n N_noxref_9_c_1902_n ) capacitor c=0.00526349f //x=5.55 \
 //y=2.08 //x2=6.775 //y2=3.7
cc_876 ( N_CLK_c_994_n N_noxref_9_c_1848_n ) capacitor c=0.0218071f //x=14.685 \
 //y=4.44 //x2=15.425 //y2=3.7
cc_877 ( N_CLK_c_992_n N_noxref_9_c_1848_n ) capacitor c=0.0218063f //x=14.8 \
 //y=2.08 //x2=15.425 //y2=3.7
cc_878 ( N_CLK_c_994_n N_noxref_9_c_1912_n ) capacitor c=4.78625e-19 \
 //x=14.685 //y=4.44 //x2=11.585 //y2=3.7
cc_879 ( N_CLK_c_992_n N_noxref_9_c_1949_n ) capacitor c=0.00117715f //x=14.8 \
 //y=2.08 //x2=15.655 //y2=3.7
cc_880 ( N_CLK_c_994_n N_noxref_9_c_1850_n ) capacitor c=0.0200057f //x=14.685 \
 //y=4.44 //x2=6.66 //y2=2.08
cc_881 ( N_CLK_c_1005_n N_noxref_9_c_1850_n ) capacitor c=0.00153281f \
 //x=5.665 //y=4.44 //x2=6.66 //y2=2.08
cc_882 ( N_CLK_c_991_n N_noxref_9_c_1850_n ) capacitor c=0.0489927f //x=5.55 \
 //y=2.08 //x2=6.66 //y2=2.08
cc_883 ( N_CLK_c_1042_n N_noxref_9_c_1850_n ) capacitor c=0.0023343f //x=5.64 \
 //y=1.915 //x2=6.66 //y2=2.08
cc_884 ( N_CLK_c_1045_n N_noxref_9_c_1850_n ) capacitor c=0.00142741f //x=5.55 \
 //y=4.7 //x2=6.66 //y2=2.08
cc_885 ( N_CLK_c_994_n N_noxref_9_c_1851_n ) capacitor c=0.0200057f //x=14.685 \
 //y=4.44 //x2=11.47 //y2=2.08
cc_886 ( N_CLK_c_994_n N_noxref_9_c_1864_n ) capacitor c=0.00325337f \
 //x=14.685 //y=4.44 //x2=14.975 //y2=5.2
cc_887 ( N_CLK_c_1054_n N_noxref_9_c_1864_n ) capacitor c=0.0126974f //x=14.8 \
 //y=4.535 //x2=14.975 //y2=5.2
cc_888 ( N_CLK_c_992_n N_noxref_9_c_1864_n ) capacitor c=3.74769e-19 //x=14.8 \
 //y=2.08 //x2=14.975 //y2=5.2
cc_889 ( N_CLK_M33_noxref_g N_noxref_9_c_1864_n ) capacitor c=0.0166421f \
 //x=14.84 //y=6.02 //x2=14.975 //y2=5.2
cc_890 ( N_CLK_c_1075_n N_noxref_9_c_1864_n ) capacitor c=0.00346519f \
 //x=14.83 //y=4.7 //x2=14.975 //y2=5.2
cc_891 ( N_CLK_c_994_n N_noxref_9_c_1868_n ) capacitor c=0.0172877f //x=14.685 \
 //y=4.44 //x2=14.265 //y2=5.2
cc_892 ( N_CLK_M34_noxref_g N_noxref_9_c_1870_n ) capacitor c=0.0199348f \
 //x=15.28 //y=6.02 //x2=15.455 //y2=5.2
cc_893 ( N_CLK_c_1101_p N_noxref_9_c_1852_n ) capacitor c=0.00371277f \
 //x=15.21 //y=1.405 //x2=15.455 //y2=1.655
cc_894 ( N_CLK_c_1072_n N_noxref_9_c_1852_n ) capacitor c=0.00457401f \
 //x=15.365 //y=1.25 //x2=15.455 //y2=1.655
cc_895 ( N_CLK_c_994_n N_noxref_9_c_1853_n ) capacitor c=0.00707546f \
 //x=14.685 //y=4.44 //x2=15.54 //y2=3.7
cc_896 ( N_CLK_c_1054_n N_noxref_9_c_1853_n ) capacitor c=0.00923416f //x=14.8 \
 //y=4.535 //x2=15.54 //y2=3.7
cc_897 ( N_CLK_c_992_n N_noxref_9_c_1853_n ) capacitor c=0.0733345f //x=14.8 \
 //y=2.08 //x2=15.54 //y2=3.7
cc_898 ( N_CLK_c_1082_p N_noxref_9_c_1853_n ) capacitor c=0.0142673f \
 //x=15.205 //y=4.79 //x2=15.54 //y2=3.7
cc_899 ( N_CLK_c_1073_n N_noxref_9_c_1853_n ) capacitor c=0.00731987f //x=14.8 \
 //y=2.08 //x2=15.54 //y2=3.7
cc_900 ( N_CLK_c_1133_p N_noxref_9_c_1853_n ) capacitor c=0.00306024f //x=14.8 \
 //y=1.915 //x2=15.54 //y2=3.7
cc_901 ( N_CLK_c_1075_n N_noxref_9_c_1853_n ) capacitor c=0.00518077f \
 //x=14.83 //y=4.7 //x2=15.54 //y2=3.7
cc_902 ( N_CLK_c_1082_p N_noxref_9_c_1972_n ) capacitor c=0.00408717f \
 //x=15.205 //y=4.79 //x2=15.06 //y2=5.2
cc_903 ( N_CLK_M21_noxref_g N_noxref_9_M23_noxref_g ) capacitor c=0.0101598f \
 //x=5.52 //y=6.02 //x2=6.4 //y2=6.02
cc_904 ( N_CLK_M22_noxref_g N_noxref_9_M23_noxref_g ) capacitor c=0.0602553f \
 //x=5.96 //y=6.02 //x2=6.4 //y2=6.02
cc_905 ( N_CLK_M22_noxref_g N_noxref_9_M24_noxref_g ) capacitor c=0.0101598f \
 //x=5.96 //y=6.02 //x2=6.84 //y2=6.02
cc_906 ( N_CLK_c_1039_n N_noxref_9_c_1976_n ) capacitor c=0.00456962f //x=5.64 \
 //y=0.91 //x2=6.65 //y2=0.915
cc_907 ( N_CLK_c_1040_n N_noxref_9_c_1977_n ) capacitor c=0.00438372f //x=5.64 \
 //y=1.22 //x2=6.65 //y2=1.26
cc_908 ( N_CLK_c_1041_n N_noxref_9_c_1978_n ) capacitor c=0.00438372f //x=5.64 \
 //y=1.45 //x2=6.65 //y2=1.57
cc_909 ( N_CLK_c_991_n N_noxref_9_c_1907_n ) capacitor c=0.00228632f //x=5.55 \
 //y=2.08 //x2=6.66 //y2=2.08
cc_910 ( N_CLK_c_1042_n N_noxref_9_c_1907_n ) capacitor c=0.00933826f //x=5.64 \
 //y=1.915 //x2=6.66 //y2=2.08
cc_911 ( N_CLK_c_1042_n N_noxref_9_c_1981_n ) capacitor c=0.00438372f //x=5.64 \
 //y=1.915 //x2=6.66 //y2=1.915
cc_912 ( N_CLK_c_994_n N_noxref_9_c_1982_n ) capacitor c=0.0111881f //x=14.685 \
 //y=4.44 //x2=6.66 //y2=4.7
cc_913 ( N_CLK_c_991_n N_noxref_9_c_1982_n ) capacitor c=0.00218014f //x=5.55 \
 //y=2.08 //x2=6.66 //y2=4.7
cc_914 ( N_CLK_c_1095_p N_noxref_9_c_1982_n ) capacitor c=0.0611812f //x=5.885 \
 //y=4.79 //x2=6.66 //y2=4.7
cc_915 ( N_CLK_c_1045_n N_noxref_9_c_1982_n ) capacitor c=0.00487508f //x=5.55 \
 //y=4.7 //x2=6.66 //y2=4.7
cc_916 ( N_CLK_c_994_n N_noxref_9_c_1939_n ) capacitor c=0.0111881f //x=14.685 \
 //y=4.44 //x2=11.47 //y2=4.7
cc_917 ( N_CLK_c_1063_n N_noxref_9_M9_noxref_d ) capacitor c=0.00217566f \
 //x=14.835 //y=0.905 //x2=14.91 //y2=0.905
cc_918 ( N_CLK_c_1066_n N_noxref_9_M9_noxref_d ) capacitor c=0.0034598f \
 //x=14.835 //y=1.25 //x2=14.91 //y2=0.905
cc_919 ( N_CLK_c_1068_n N_noxref_9_M9_noxref_d ) capacitor c=0.00669531f \
 //x=14.835 //y=1.56 //x2=14.91 //y2=0.905
cc_920 ( N_CLK_c_1153_p N_noxref_9_M9_noxref_d ) capacitor c=0.00241102f \
 //x=15.21 //y=0.75 //x2=14.91 //y2=0.905
cc_921 ( N_CLK_c_1101_p N_noxref_9_M9_noxref_d ) capacitor c=0.0137169f \
 //x=15.21 //y=1.405 //x2=14.91 //y2=0.905
cc_922 ( N_CLK_c_1071_n N_noxref_9_M9_noxref_d ) capacitor c=0.00132245f \
 //x=15.365 //y=0.905 //x2=14.91 //y2=0.905
cc_923 ( N_CLK_c_1072_n N_noxref_9_M9_noxref_d ) capacitor c=0.00566463f \
 //x=15.365 //y=1.25 //x2=14.91 //y2=0.905
cc_924 ( N_CLK_c_1133_p N_noxref_9_M9_noxref_d ) capacitor c=0.00660593f \
 //x=14.8 //y=1.915 //x2=14.91 //y2=0.905
cc_925 ( N_CLK_M33_noxref_g N_noxref_9_M33_noxref_d ) capacitor c=0.0173476f \
 //x=14.84 //y=6.02 //x2=14.915 //y2=5.02
cc_926 ( N_CLK_M34_noxref_g N_noxref_9_M33_noxref_d ) capacitor c=0.0179769f \
 //x=15.28 //y=6.02 //x2=14.915 //y2=5.02
cc_927 ( N_CLK_c_1034_n N_noxref_13_c_2452_n ) capacitor c=0.0167228f \
 //x=5.115 //y=0.91 //x2=5.775 //y2=0.54
cc_928 ( N_CLK_c_1039_n N_noxref_13_c_2452_n ) capacitor c=0.00534519f \
 //x=5.64 //y=0.91 //x2=5.775 //y2=0.54
cc_929 ( N_CLK_c_991_n N_noxref_13_c_2472_n ) capacitor c=0.012334f //x=5.55 \
 //y=2.08 //x2=5.775 //y2=1.59
cc_930 ( N_CLK_c_1037_n N_noxref_13_c_2472_n ) capacitor c=0.0153476f \
 //x=5.115 //y=1.22 //x2=5.775 //y2=1.59
cc_931 ( N_CLK_c_1042_n N_noxref_13_c_2472_n ) capacitor c=0.0219329f //x=5.64 \
 //y=1.915 //x2=5.775 //y2=1.59
cc_932 ( N_CLK_c_1034_n N_noxref_13_M2_noxref_s ) capacitor c=0.00798959f \
 //x=5.115 //y=0.91 //x2=3.785 //y2=0.375
cc_933 ( N_CLK_c_1041_n N_noxref_13_M2_noxref_s ) capacitor c=0.00212176f \
 //x=5.64 //y=1.45 //x2=3.785 //y2=0.375
cc_934 ( N_CLK_c_1042_n N_noxref_13_M2_noxref_s ) capacitor c=0.00298115f \
 //x=5.64 //y=1.915 //x2=3.785 //y2=0.375
cc_935 ( N_CLK_c_1168_p N_noxref_14_c_2497_n ) capacitor c=2.14837e-19 \
 //x=5.485 //y=0.755 //x2=6.345 //y2=0.995
cc_936 ( N_CLK_c_1039_n N_noxref_14_c_2497_n ) capacitor c=0.00123426f \
 //x=5.64 //y=0.91 //x2=6.345 //y2=0.995
cc_937 ( N_CLK_c_1040_n N_noxref_14_c_2497_n ) capacitor c=0.0129288f //x=5.64 \
 //y=1.22 //x2=6.345 //y2=0.995
cc_938 ( N_CLK_c_1041_n N_noxref_14_c_2497_n ) capacitor c=0.00142359f \
 //x=5.64 //y=1.45 //x2=6.345 //y2=0.995
cc_939 ( N_CLK_c_1034_n N_noxref_14_M3_noxref_d ) capacitor c=0.00223875f \
 //x=5.115 //y=0.91 //x2=5.19 //y2=0.91
cc_940 ( N_CLK_c_1037_n N_noxref_14_M3_noxref_d ) capacitor c=0.00262485f \
 //x=5.115 //y=1.22 //x2=5.19 //y2=0.91
cc_941 ( N_CLK_c_1168_p N_noxref_14_M3_noxref_d ) capacitor c=0.00220746f \
 //x=5.485 //y=0.755 //x2=5.19 //y2=0.91
cc_942 ( N_CLK_c_1175_p N_noxref_14_M3_noxref_d ) capacitor c=0.00194798f \
 //x=5.485 //y=1.375 //x2=5.19 //y2=0.91
cc_943 ( N_CLK_c_1039_n N_noxref_14_M3_noxref_d ) capacitor c=0.00198465f \
 //x=5.64 //y=0.91 //x2=5.19 //y2=0.91
cc_944 ( N_CLK_c_1040_n N_noxref_14_M3_noxref_d ) capacitor c=0.00128384f \
 //x=5.64 //y=1.22 //x2=5.19 //y2=0.91
cc_945 ( N_CLK_c_1039_n N_noxref_14_M4_noxref_s ) capacitor c=7.21316e-19 \
 //x=5.64 //y=0.91 //x2=6.295 //y2=0.375
cc_946 ( N_CLK_c_1040_n N_noxref_14_M4_noxref_s ) capacitor c=0.00348171f \
 //x=5.64 //y=1.22 //x2=6.295 //y2=0.375
cc_947 ( N_CLK_c_1068_n N_noxref_17_c_2664_n ) capacitor c=0.00623646f \
 //x=14.835 //y=1.56 //x2=14.615 //y2=1.495
cc_948 ( N_CLK_c_1073_n N_noxref_17_c_2664_n ) capacitor c=0.00173579f \
 //x=14.8 //y=2.08 //x2=14.615 //y2=1.495
cc_949 ( N_CLK_c_992_n N_noxref_17_c_2665_n ) capacitor c=0.00156605f //x=14.8 \
 //y=2.08 //x2=15.5 //y2=0.53
cc_950 ( N_CLK_c_1063_n N_noxref_17_c_2665_n ) capacitor c=0.0188655f \
 //x=14.835 //y=0.905 //x2=15.5 //y2=0.53
cc_951 ( N_CLK_c_1071_n N_noxref_17_c_2665_n ) capacitor c=0.00656458f \
 //x=15.365 //y=0.905 //x2=15.5 //y2=0.53
cc_952 ( N_CLK_c_1073_n N_noxref_17_c_2665_n ) capacitor c=2.1838e-19 //x=14.8 \
 //y=2.08 //x2=15.5 //y2=0.53
cc_953 ( N_CLK_c_1063_n N_noxref_17_M8_noxref_s ) capacitor c=0.00623646f \
 //x=14.835 //y=0.905 //x2=13.51 //y2=0.365
cc_954 ( N_CLK_c_1071_n N_noxref_17_M8_noxref_s ) capacitor c=0.0143002f \
 //x=15.365 //y=0.905 //x2=13.51 //y2=0.365
cc_955 ( N_CLK_c_1072_n N_noxref_17_M8_noxref_s ) capacitor c=0.00290153f \
 //x=15.365 //y=1.25 //x2=13.51 //y2=0.365
cc_956 ( N_noxref_6_c_1195_n QN ) capacitor c=0.00396868f //x=17.39 //y=2.08 \
 //x2=18.87 //y2=2.59
cc_957 ( N_noxref_6_M36_noxref_g N_QN_c_1494_n ) capacitor c=0.0187084f \
 //x=17.73 //y=6.02 //x2=18.305 //y2=5.2
cc_958 ( N_noxref_6_c_1215_n N_QN_c_1498_n ) capacitor c=0.00144307f \
 //x=17.275 //y=4.07 //x2=17.595 //y2=5.2
cc_959 ( N_noxref_6_c_1195_n N_QN_c_1498_n ) capacitor c=0.00529872f //x=17.39 \
 //y=2.08 //x2=17.595 //y2=5.2
cc_960 ( N_noxref_6_M35_noxref_g N_QN_c_1498_n ) capacitor c=0.0177326f \
 //x=17.29 //y=6.02 //x2=17.595 //y2=5.2
cc_961 ( N_noxref_6_c_1254_n N_QN_c_1498_n ) capacitor c=0.00585724f //x=17.39 \
 //y=4.7 //x2=17.595 //y2=5.2
cc_962 ( N_noxref_6_M36_noxref_g N_QN_M35_noxref_d ) capacitor c=0.0173476f \
 //x=17.73 //y=6.02 //x2=17.365 //y2=5.02
cc_963 ( N_noxref_6_c_1215_n N_SN_c_1620_n ) capacitor c=0.0218224f //x=17.275 \
 //y=4.07 //x2=21.715 //y2=2.22
cc_964 ( N_noxref_6_c_1195_n N_SN_c_1620_n ) capacitor c=0.0233481f //x=17.39 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_965 ( N_noxref_6_c_1200_n N_SN_c_1620_n ) capacitor c=0.00814985f \
 //x=17.195 //y=1.915 //x2=21.715 //y2=2.22
cc_966 ( N_noxref_6_c_1215_n N_SN_c_1630_n ) capacitor c=5.95893e-19 \
 //x=17.275 //y=4.07 //x2=10.475 //y2=2.22
cc_967 ( N_noxref_6_c_1215_n N_SN_c_1631_n ) capacitor c=0.0190126f //x=17.275 \
 //y=4.07 //x2=10.36 //y2=2.08
cc_968 ( N_noxref_6_c_1294_n N_SN_c_1631_n ) capacitor c=4.52713e-19 //x=7.397 \
 //y=3.905 //x2=10.36 //y2=2.08
cc_969 ( N_noxref_6_c_1189_n N_noxref_9_c_1846_n ) capacitor c=0.044143f \
 //x=7.28 //y=4.07 //x2=11.355 //y2=3.7
cc_970 ( N_noxref_6_c_1215_n N_noxref_9_c_1846_n ) capacitor c=0.340271f \
 //x=17.275 //y=4.07 //x2=11.355 //y2=3.7
cc_971 ( N_noxref_6_c_1224_n N_noxref_9_c_1846_n ) capacitor c=0.0267581f \
 //x=7.51 //y=4.07 //x2=11.355 //y2=3.7
cc_972 ( N_noxref_6_c_1244_n N_noxref_9_c_1846_n ) capacitor c=0.00219785f \
 //x=7.395 //y=4.07 //x2=11.355 //y2=3.7
cc_973 ( N_noxref_6_c_1294_n N_noxref_9_c_1846_n ) capacitor c=0.0223643f \
 //x=7.397 //y=3.905 //x2=11.355 //y2=3.7
cc_974 ( N_noxref_6_c_1189_n N_noxref_9_c_1902_n ) capacitor c=0.0292842f \
 //x=7.28 //y=4.07 //x2=6.775 //y2=3.7
cc_975 ( N_noxref_6_c_1294_n N_noxref_9_c_1902_n ) capacitor c=0.00179385f \
 //x=7.397 //y=3.905 //x2=6.775 //y2=3.7
cc_976 ( N_noxref_6_c_1215_n N_noxref_9_c_1848_n ) capacitor c=0.339174f \
 //x=17.275 //y=4.07 //x2=15.425 //y2=3.7
cc_977 ( N_noxref_6_c_1215_n N_noxref_9_c_1912_n ) capacitor c=0.026596f \
 //x=17.275 //y=4.07 //x2=11.585 //y2=3.7
cc_978 ( N_noxref_6_c_1215_n N_noxref_9_c_1849_n ) capacitor c=0.17615f \
 //x=17.275 //y=4.07 //x2=22.825 //y2=3.7
cc_979 ( N_noxref_6_c_1195_n N_noxref_9_c_1849_n ) capacitor c=0.0253978f \
 //x=17.39 //y=2.08 //x2=22.825 //y2=3.7
cc_980 ( N_noxref_6_c_1254_n N_noxref_9_c_1849_n ) capacitor c=0.00463981f \
 //x=17.39 //y=4.7 //x2=22.825 //y2=3.7
cc_981 ( N_noxref_6_c_1215_n N_noxref_9_c_1949_n ) capacitor c=0.026743f \
 //x=17.275 //y=4.07 //x2=15.655 //y2=3.7
cc_982 ( N_noxref_6_c_1195_n N_noxref_9_c_1949_n ) capacitor c=7.01366e-19 \
 //x=17.39 //y=2.08 //x2=15.655 //y2=3.7
cc_983 ( N_noxref_6_c_1189_n N_noxref_9_c_1850_n ) capacitor c=0.0197867f \
 //x=7.28 //y=4.07 //x2=6.66 //y2=2.08
cc_984 ( N_noxref_6_c_1224_n N_noxref_9_c_1850_n ) capacitor c=0.00180189f \
 //x=7.51 //y=4.07 //x2=6.66 //y2=2.08
cc_985 ( N_noxref_6_c_1336_n N_noxref_9_c_1850_n ) capacitor c=0.0163236f \
 //x=7.4 //y=5.07 //x2=6.66 //y2=2.08
cc_986 ( N_noxref_6_c_1375_p N_noxref_9_c_1850_n ) capacitor c=0.016476f \
 //x=6.62 //y=5.155 //x2=6.66 //y2=2.08
cc_987 ( N_noxref_6_c_1244_n N_noxref_9_c_1850_n ) capacitor c=0.00966503f \
 //x=7.395 //y=4.07 //x2=6.66 //y2=2.08
cc_988 ( N_noxref_6_c_1294_n N_noxref_9_c_1850_n ) capacitor c=0.0580095f \
 //x=7.397 //y=3.905 //x2=6.66 //y2=2.08
cc_989 ( N_noxref_6_c_1215_n N_noxref_9_c_1851_n ) capacitor c=0.0198068f \
 //x=17.275 //y=4.07 //x2=11.47 //y2=2.08
cc_990 ( N_noxref_6_c_1215_n N_noxref_9_c_1864_n ) capacitor c=0.0126022f \
 //x=17.275 //y=4.07 //x2=14.975 //y2=5.2
cc_991 ( N_noxref_6_c_1215_n N_noxref_9_c_1853_n ) capacitor c=0.0253623f \
 //x=17.275 //y=4.07 //x2=15.54 //y2=3.7
cc_992 ( N_noxref_6_c_1195_n N_noxref_9_c_1853_n ) capacitor c=0.0145047f \
 //x=17.39 //y=2.08 //x2=15.54 //y2=3.7
cc_993 ( N_noxref_6_c_1233_n N_noxref_9_M23_noxref_g ) capacitor c=0.01736f \
 //x=6.535 //y=5.155 //x2=6.4 //y2=6.02
cc_994 ( N_noxref_6_M23_noxref_d N_noxref_9_M23_noxref_g ) capacitor \
 c=0.0180032f //x=6.475 //y=5.02 //x2=6.4 //y2=6.02
cc_995 ( N_noxref_6_c_1237_n N_noxref_9_M24_noxref_g ) capacitor c=0.0194981f \
 //x=7.315 //y=5.155 //x2=6.84 //y2=6.02
cc_996 ( N_noxref_6_M23_noxref_d N_noxref_9_M24_noxref_g ) capacitor \
 c=0.0194246f //x=6.475 //y=5.02 //x2=6.84 //y2=6.02
cc_997 ( N_noxref_6_M4_noxref_d N_noxref_9_c_1976_n ) capacitor c=0.00217566f \
 //x=6.725 //y=0.915 //x2=6.65 //y2=0.915
cc_998 ( N_noxref_6_M4_noxref_d N_noxref_9_c_1977_n ) capacitor c=0.0034598f \
 //x=6.725 //y=0.915 //x2=6.65 //y2=1.26
cc_999 ( N_noxref_6_M4_noxref_d N_noxref_9_c_1978_n ) capacitor c=0.00544291f \
 //x=6.725 //y=0.915 //x2=6.65 //y2=1.57
cc_1000 ( N_noxref_6_M4_noxref_d N_noxref_9_c_2028_n ) capacitor c=0.00241102f \
 //x=6.725 //y=0.915 //x2=7.025 //y2=0.76
cc_1001 ( N_noxref_6_c_1194_n N_noxref_9_c_2029_n ) capacitor c=0.00359704f \
 //x=7.315 //y=1.665 //x2=7.025 //y2=1.415
cc_1002 ( N_noxref_6_M4_noxref_d N_noxref_9_c_2029_n ) capacitor c=0.0140297f \
 //x=6.725 //y=0.915 //x2=7.025 //y2=1.415
cc_1003 ( N_noxref_6_M4_noxref_d N_noxref_9_c_2031_n ) capacitor c=0.00219619f \
 //x=6.725 //y=0.915 //x2=7.18 //y2=0.915
cc_1004 ( N_noxref_6_c_1194_n N_noxref_9_c_2032_n ) capacitor c=0.00457401f \
 //x=7.315 //y=1.665 //x2=7.18 //y2=1.26
cc_1005 ( N_noxref_6_M4_noxref_d N_noxref_9_c_2032_n ) capacitor c=0.00603828f \
 //x=6.725 //y=0.915 //x2=7.18 //y2=1.26
cc_1006 ( N_noxref_6_c_1294_n N_noxref_9_c_1907_n ) capacitor c=0.00772308f \
 //x=7.397 //y=3.905 //x2=6.66 //y2=2.08
cc_1007 ( N_noxref_6_c_1294_n N_noxref_9_c_1981_n ) capacitor c=0.00404774f \
 //x=7.397 //y=3.905 //x2=6.66 //y2=1.915
cc_1008 ( N_noxref_6_M4_noxref_d N_noxref_9_c_1981_n ) capacitor c=0.00661782f \
 //x=6.725 //y=0.915 //x2=6.66 //y2=1.915
cc_1009 ( N_noxref_6_c_1237_n N_noxref_9_c_1982_n ) capacitor c=0.00201851f \
 //x=7.315 //y=5.155 //x2=6.66 //y2=4.7
cc_1010 ( N_noxref_6_c_1336_n N_noxref_9_c_1982_n ) capacitor c=0.0151148f \
 //x=7.4 //y=5.07 //x2=6.66 //y2=4.7
cc_1011 ( N_noxref_6_c_1375_p N_noxref_9_c_1982_n ) capacitor c=0.00475601f \
 //x=6.62 //y=5.155 //x2=6.66 //y2=4.7
cc_1012 ( N_noxref_6_c_1195_n N_noxref_10_c_2213_n ) capacitor c=0.00735597f \
 //x=17.39 //y=2.08 //x2=18.245 //y2=3.33
cc_1013 ( N_noxref_6_c_1195_n N_noxref_10_c_2214_n ) capacitor c=0.00400249f \
 //x=17.39 //y=2.08 //x2=18.13 //y2=4.535
cc_1014 ( N_noxref_6_c_1254_n N_noxref_10_c_2214_n ) capacitor c=0.00417994f \
 //x=17.39 //y=4.7 //x2=18.13 //y2=4.535
cc_1015 ( N_noxref_6_c_1215_n N_noxref_10_c_2172_n ) capacitor c=0.00735597f \
 //x=17.275 //y=4.07 //x2=18.13 //y2=2.08
cc_1016 ( N_noxref_6_c_1195_n N_noxref_10_c_2172_n ) capacitor c=0.0788112f \
 //x=17.39 //y=2.08 //x2=18.13 //y2=2.08
cc_1017 ( N_noxref_6_c_1200_n N_noxref_10_c_2172_n ) capacitor c=0.00284029f \
 //x=17.195 //y=1.915 //x2=18.13 //y2=2.08
cc_1018 ( N_noxref_6_M35_noxref_g N_noxref_10_M37_noxref_g ) capacitor \
 c=0.0104611f //x=17.29 //y=6.02 //x2=18.17 //y2=6.02
cc_1019 ( N_noxref_6_M36_noxref_g N_noxref_10_M37_noxref_g ) capacitor \
 c=0.106811f //x=17.73 //y=6.02 //x2=18.17 //y2=6.02
cc_1020 ( N_noxref_6_M36_noxref_g N_noxref_10_M38_noxref_g ) capacitor \
 c=0.0100341f //x=17.73 //y=6.02 //x2=18.61 //y2=6.02
cc_1021 ( N_noxref_6_c_1196_n N_noxref_10_c_2222_n ) capacitor c=4.86506e-19 \
 //x=17.195 //y=0.865 //x2=18.165 //y2=0.905
cc_1022 ( N_noxref_6_c_1198_n N_noxref_10_c_2222_n ) capacitor c=0.00152104f \
 //x=17.195 //y=1.21 //x2=18.165 //y2=0.905
cc_1023 ( N_noxref_6_c_1203_n N_noxref_10_c_2222_n ) capacitor c=0.0151475f \
 //x=17.725 //y=0.865 //x2=18.165 //y2=0.905
cc_1024 ( N_noxref_6_c_1199_n N_noxref_10_c_2225_n ) capacitor c=0.00109982f \
 //x=17.195 //y=1.52 //x2=18.165 //y2=1.25
cc_1025 ( N_noxref_6_c_1205_n N_noxref_10_c_2225_n ) capacitor c=0.0111064f \
 //x=17.725 //y=1.21 //x2=18.165 //y2=1.25
cc_1026 ( N_noxref_6_c_1199_n N_noxref_10_c_2227_n ) capacitor c=9.57794e-19 \
 //x=17.195 //y=1.52 //x2=18.165 //y2=1.56
cc_1027 ( N_noxref_6_c_1200_n N_noxref_10_c_2227_n ) capacitor c=0.00662747f \
 //x=17.195 //y=1.915 //x2=18.165 //y2=1.56
cc_1028 ( N_noxref_6_c_1205_n N_noxref_10_c_2227_n ) capacitor c=0.00862358f \
 //x=17.725 //y=1.21 //x2=18.165 //y2=1.56
cc_1029 ( N_noxref_6_c_1203_n N_noxref_10_c_2230_n ) capacitor c=0.00124821f \
 //x=17.725 //y=0.865 //x2=18.695 //y2=0.905
cc_1030 ( N_noxref_6_c_1205_n N_noxref_10_c_2231_n ) capacitor c=0.00200715f \
 //x=17.725 //y=1.21 //x2=18.695 //y2=1.25
cc_1031 ( N_noxref_6_c_1195_n N_noxref_10_c_2232_n ) capacitor c=0.00282278f \
 //x=17.39 //y=2.08 //x2=18.13 //y2=2.08
cc_1032 ( N_noxref_6_c_1200_n N_noxref_10_c_2232_n ) capacitor c=0.0172771f \
 //x=17.195 //y=1.915 //x2=18.13 //y2=2.08
cc_1033 ( N_noxref_6_c_1195_n N_noxref_10_c_2234_n ) capacitor c=0.00344981f \
 //x=17.39 //y=2.08 //x2=18.16 //y2=4.7
cc_1034 ( N_noxref_6_c_1254_n N_noxref_10_c_2234_n ) capacitor c=0.0293367f \
 //x=17.39 //y=4.7 //x2=18.16 //y2=4.7
cc_1035 ( N_noxref_6_c_1191_n N_D_c_2340_n ) capacitor c=0.00642908f //x=1.965 \
 //y=4.07 //x2=1.11 //y2=2.08
cc_1036 ( N_noxref_6_c_1284_n N_D_c_2340_n ) capacitor c=0.00400249f //x=1.85 \
 //y=4.535 //x2=1.11 //y2=2.08
cc_1037 ( N_noxref_6_c_1192_n N_D_c_2340_n ) capacitor c=0.0865678f //x=1.85 \
 //y=2.08 //x2=1.11 //y2=2.08
cc_1038 ( N_noxref_6_c_1311_n N_D_c_2340_n ) capacitor c=0.00307062f //x=1.85 \
 //y=2.08 //x2=1.11 //y2=2.08
cc_1039 ( N_noxref_6_c_1314_n N_D_c_2340_n ) capacitor c=0.00344981f //x=1.88 \
 //y=4.7 //x2=1.11 //y2=2.08
cc_1040 ( N_noxref_6_M17_noxref_g N_D_M15_noxref_g ) capacitor c=0.0104611f \
 //x=1.89 //y=6.02 //x2=1.01 //y2=6.02
cc_1041 ( N_noxref_6_M17_noxref_g N_D_M16_noxref_g ) capacitor c=0.106811f \
 //x=1.89 //y=6.02 //x2=1.45 //y2=6.02
cc_1042 ( N_noxref_6_M18_noxref_g N_D_M16_noxref_g ) capacitor c=0.0100341f \
 //x=2.33 //y=6.02 //x2=1.45 //y2=6.02
cc_1043 ( N_noxref_6_c_1300_n N_D_c_2341_n ) capacitor c=4.86506e-19 //x=1.885 \
 //y=0.905 //x2=0.915 //y2=0.865
cc_1044 ( N_noxref_6_c_1300_n N_D_c_2343_n ) capacitor c=0.00152104f //x=1.885 \
 //y=0.905 //x2=0.915 //y2=1.21
cc_1045 ( N_noxref_6_c_1301_n N_D_c_2344_n ) capacitor c=0.00109982f //x=1.885 \
 //y=1.25 //x2=0.915 //y2=1.52
cc_1046 ( N_noxref_6_c_1302_n N_D_c_2344_n ) capacitor c=9.57794e-19 //x=1.885 \
 //y=1.56 //x2=0.915 //y2=1.52
cc_1047 ( N_noxref_6_c_1192_n N_D_c_2345_n ) capacitor c=0.00308814f //x=1.85 \
 //y=2.08 //x2=0.915 //y2=1.915
cc_1048 ( N_noxref_6_c_1302_n N_D_c_2345_n ) capacitor c=0.00662747f //x=1.885 \
 //y=1.56 //x2=0.915 //y2=1.915
cc_1049 ( N_noxref_6_c_1311_n N_D_c_2345_n ) capacitor c=0.0179092f //x=1.85 \
 //y=2.08 //x2=0.915 //y2=1.915
cc_1050 ( N_noxref_6_c_1300_n N_D_c_2348_n ) capacitor c=0.0151475f //x=1.885 \
 //y=0.905 //x2=1.445 //y2=0.865
cc_1051 ( N_noxref_6_c_1308_n N_D_c_2348_n ) capacitor c=0.00124821f //x=2.415 \
 //y=0.905 //x2=1.445 //y2=0.865
cc_1052 ( N_noxref_6_c_1301_n N_D_c_2350_n ) capacitor c=0.0111064f //x=1.885 \
 //y=1.25 //x2=1.445 //y2=1.21
cc_1053 ( N_noxref_6_c_1302_n N_D_c_2350_n ) capacitor c=0.00862358f //x=1.885 \
 //y=1.56 //x2=1.445 //y2=1.21
cc_1054 ( N_noxref_6_c_1309_n N_D_c_2350_n ) capacitor c=0.00200715f //x=2.415 \
 //y=1.25 //x2=1.445 //y2=1.21
cc_1055 ( N_noxref_6_c_1284_n N_D_c_2358_n ) capacitor c=0.00417994f //x=1.85 \
 //y=4.535 //x2=1.11 //y2=4.7
cc_1056 ( N_noxref_6_c_1314_n N_D_c_2358_n ) capacitor c=0.0293367f //x=1.88 \
 //y=4.7 //x2=1.11 //y2=4.7
cc_1057 ( N_noxref_6_c_1191_n N_noxref_12_c_2404_n ) capacitor c=3.32378e-19 \
 //x=1.965 //y=4.07 //x2=1.665 //y2=1.495
cc_1058 ( N_noxref_6_c_1302_n N_noxref_12_c_2404_n ) capacitor c=0.00623646f \
 //x=1.885 //y=1.56 //x2=1.665 //y2=1.495
cc_1059 ( N_noxref_6_c_1311_n N_noxref_12_c_2404_n ) capacitor c=0.00176439f \
 //x=1.85 //y=2.08 //x2=1.665 //y2=1.495
cc_1060 ( N_noxref_6_c_1192_n N_noxref_12_c_2405_n ) capacitor c=0.00161845f \
 //x=1.85 //y=2.08 //x2=2.55 //y2=0.53
cc_1061 ( N_noxref_6_c_1300_n N_noxref_12_c_2405_n ) capacitor c=0.0186143f \
 //x=1.885 //y=0.905 //x2=2.55 //y2=0.53
cc_1062 ( N_noxref_6_c_1308_n N_noxref_12_c_2405_n ) capacitor c=0.00656458f \
 //x=2.415 //y=0.905 //x2=2.55 //y2=0.53
cc_1063 ( N_noxref_6_c_1311_n N_noxref_12_c_2405_n ) capacitor c=2.1838e-19 \
 //x=1.85 //y=2.08 //x2=2.55 //y2=0.53
cc_1064 ( N_noxref_6_c_1300_n N_noxref_12_M0_noxref_s ) capacitor \
 c=0.00623646f //x=1.885 //y=0.905 //x2=0.56 //y2=0.365
cc_1065 ( N_noxref_6_c_1308_n N_noxref_12_M0_noxref_s ) capacitor c=0.0143002f \
 //x=2.415 //y=0.905 //x2=0.56 //y2=0.365
cc_1066 ( N_noxref_6_c_1309_n N_noxref_12_M0_noxref_s ) capacitor \
 c=0.00290153f //x=2.415 //y=1.25 //x2=0.56 //y2=0.365
cc_1067 ( N_noxref_6_M4_noxref_d N_noxref_13_M2_noxref_s ) capacitor \
 c=0.00309936f //x=6.725 //y=0.915 //x2=3.785 //y2=0.375
cc_1068 ( N_noxref_6_c_1194_n N_noxref_14_c_2502_n ) capacitor c=0.00461497f \
 //x=7.315 //y=1.665 //x2=7.315 //y2=0.54
cc_1069 ( N_noxref_6_M4_noxref_d N_noxref_14_c_2502_n ) capacitor c=0.0116817f \
 //x=6.725 //y=0.915 //x2=7.315 //y2=0.54
cc_1070 ( N_noxref_6_c_1293_n N_noxref_14_c_2528_n ) capacitor c=0.0200405f \
 //x=7 //y=1.665 //x2=6.43 //y2=0.995
cc_1071 ( N_noxref_6_M4_noxref_d N_noxref_14_M3_noxref_d ) capacitor \
 c=5.27807e-19 //x=6.725 //y=0.915 //x2=5.19 //y2=0.91
cc_1072 ( N_noxref_6_c_1194_n N_noxref_14_M4_noxref_s ) capacitor c=0.0201579f \
 //x=7.315 //y=1.665 //x2=6.295 //y2=0.375
cc_1073 ( N_noxref_6_M4_noxref_d N_noxref_14_M4_noxref_s ) capacitor \
 c=0.0426368f //x=6.725 //y=0.915 //x2=6.295 //y2=0.375
cc_1074 ( N_noxref_6_c_1194_n N_noxref_15_c_2566_n ) capacitor c=3.83325e-19 \
 //x=7.315 //y=1.665 //x2=8.73 //y2=1.505
cc_1075 ( N_noxref_6_M4_noxref_d N_noxref_15_M5_noxref_s ) capacitor \
 c=2.55333e-19 //x=6.725 //y=0.915 //x2=8.595 //y2=0.375
cc_1076 ( N_noxref_6_c_1200_n N_noxref_18_c_2728_n ) capacitor c=0.0034165f \
 //x=17.195 //y=1.915 //x2=16.975 //y2=1.495
cc_1077 ( N_noxref_6_c_1195_n N_noxref_18_c_2709_n ) capacitor c=0.0111916f \
 //x=17.39 //y=2.08 //x2=17.86 //y2=1.58
cc_1078 ( N_noxref_6_c_1199_n N_noxref_18_c_2709_n ) capacitor c=0.00696403f \
 //x=17.195 //y=1.52 //x2=17.86 //y2=1.58
cc_1079 ( N_noxref_6_c_1200_n N_noxref_18_c_2709_n ) capacitor c=0.0174694f \
 //x=17.195 //y=1.915 //x2=17.86 //y2=1.58
cc_1080 ( N_noxref_6_c_1202_n N_noxref_18_c_2709_n ) capacitor c=0.00776811f \
 //x=17.57 //y=1.365 //x2=17.86 //y2=1.58
cc_1081 ( N_noxref_6_c_1205_n N_noxref_18_c_2709_n ) capacitor c=0.00339872f \
 //x=17.725 //y=1.21 //x2=17.86 //y2=1.58
cc_1082 ( N_noxref_6_c_1200_n N_noxref_18_c_2716_n ) capacitor c=6.71402e-19 \
 //x=17.195 //y=1.915 //x2=17.945 //y2=1.495
cc_1083 ( N_noxref_6_c_1196_n N_noxref_18_M10_noxref_s ) capacitor \
 c=0.0326577f //x=17.195 //y=0.865 //x2=16.84 //y2=0.365
cc_1084 ( N_noxref_6_c_1199_n N_noxref_18_M10_noxref_s ) capacitor \
 c=3.48408e-19 //x=17.195 //y=1.52 //x2=16.84 //y2=0.365
cc_1085 ( N_noxref_6_c_1203_n N_noxref_18_M10_noxref_s ) capacitor \
 c=0.0120759f //x=17.725 //y=0.865 //x2=16.84 //y2=0.365
cc_1086 ( N_QN_c_1475_n N_SN_c_1620_n ) capacitor c=0.0838914f //x=20.605 \
 //y=2.96 //x2=21.715 //y2=2.22
cc_1087 ( N_QN_c_1531_p N_SN_c_1620_n ) capacitor c=0.0133375f //x=18.985 \
 //y=2.96 //x2=21.715 //y2=2.22
cc_1088 ( QN N_SN_c_1620_n ) capacitor c=0.0225629f //x=18.87 //y=2.59 \
 //x2=21.715 //y2=2.22
cc_1089 ( N_QN_c_1533_p N_SN_c_1620_n ) capacitor c=0.0146822f //x=18.515 \
 //y=1.655 //x2=21.715 //y2=2.22
cc_1090 ( N_QN_c_1478_n N_SN_c_1620_n ) capacitor c=0.0235839f //x=20.72 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_1091 ( N_QN_c_1483_n N_SN_c_1620_n ) capacitor c=0.0122202f //x=20.42 \
 //y=1.915 //x2=21.715 //y2=2.22
cc_1092 ( N_QN_c_1475_n N_SN_c_1632_n ) capacitor c=0.00520283f //x=20.605 \
 //y=2.96 //x2=21.83 //y2=2.08
cc_1093 ( QN N_SN_c_1632_n ) capacitor c=5.5948e-19 //x=18.87 //y=2.59 \
 //x2=21.83 //y2=2.08
cc_1094 ( N_QN_c_1478_n N_SN_c_1632_n ) capacitor c=0.0493665f //x=20.72 \
 //y=2.08 //x2=21.83 //y2=2.08
cc_1095 ( N_QN_c_1483_n N_SN_c_1632_n ) capacitor c=0.00208635f //x=20.42 \
 //y=1.915 //x2=21.83 //y2=2.08
cc_1096 ( N_QN_c_1540_p N_SN_c_1632_n ) capacitor c=0.00147352f //x=21.285 \
 //y=4.79 //x2=21.83 //y2=2.08
cc_1097 ( N_QN_c_1510_n N_SN_c_1632_n ) capacitor c=0.00142741f //x=20.995 \
 //y=4.79 //x2=21.83 //y2=2.08
cc_1098 ( N_QN_M39_noxref_g N_SN_M41_noxref_g ) capacitor c=0.0105869f \
 //x=20.92 //y=6.02 //x2=21.8 //y2=6.02
cc_1099 ( N_QN_M40_noxref_g N_SN_M41_noxref_g ) capacitor c=0.10632f //x=21.36 \
 //y=6.02 //x2=21.8 //y2=6.02
cc_1100 ( N_QN_M40_noxref_g N_SN_M42_noxref_g ) capacitor c=0.0101598f \
 //x=21.36 //y=6.02 //x2=22.24 //y2=6.02
cc_1101 ( N_QN_c_1479_n N_SN_c_1709_n ) capacitor c=5.72482e-19 //x=20.42 \
 //y=0.875 //x2=21.395 //y2=0.91
cc_1102 ( N_QN_c_1481_n N_SN_c_1709_n ) capacitor c=0.00149976f //x=20.42 \
 //y=1.22 //x2=21.395 //y2=0.91
cc_1103 ( N_QN_c_1486_n N_SN_c_1709_n ) capacitor c=0.0160123f //x=20.95 \
 //y=0.875 //x2=21.395 //y2=0.91
cc_1104 ( N_QN_c_1482_n N_SN_c_1712_n ) capacitor c=0.00111227f //x=20.42 \
 //y=1.53 //x2=21.395 //y2=1.22
cc_1105 ( N_QN_c_1488_n N_SN_c_1712_n ) capacitor c=0.0124075f //x=20.95 \
 //y=1.22 //x2=21.395 //y2=1.22
cc_1106 ( N_QN_c_1486_n N_SN_c_1714_n ) capacitor c=0.00103227f //x=20.95 \
 //y=0.875 //x2=21.92 //y2=0.91
cc_1107 ( N_QN_c_1488_n N_SN_c_1715_n ) capacitor c=0.0010154f //x=20.95 \
 //y=1.22 //x2=21.92 //y2=1.22
cc_1108 ( N_QN_c_1488_n N_SN_c_1716_n ) capacitor c=9.23422e-19 //x=20.95 \
 //y=1.22 //x2=21.92 //y2=1.45
cc_1109 ( N_QN_c_1478_n N_SN_c_1717_n ) capacitor c=0.00203769f //x=20.72 \
 //y=2.08 //x2=21.92 //y2=1.915
cc_1110 ( N_QN_c_1483_n N_SN_c_1717_n ) capacitor c=0.00834532f //x=20.42 \
 //y=1.915 //x2=21.92 //y2=1.915
cc_1111 ( N_QN_c_1478_n N_SN_c_1719_n ) capacitor c=0.00183762f //x=20.72 \
 //y=2.08 //x2=21.83 //y2=4.7
cc_1112 ( N_QN_c_1540_p N_SN_c_1719_n ) capacitor c=0.0168581f //x=21.285 \
 //y=4.79 //x2=21.83 //y2=4.7
cc_1113 ( N_QN_c_1510_n N_SN_c_1719_n ) capacitor c=0.00484466f //x=20.995 \
 //y=4.79 //x2=21.83 //y2=4.7
cc_1114 ( N_QN_c_1475_n N_noxref_9_c_1849_n ) capacitor c=0.0116974f \
 //x=20.605 //y=2.96 //x2=22.825 //y2=3.7
cc_1115 ( N_QN_c_1531_p N_noxref_9_c_1849_n ) capacitor c=8.88514e-19 \
 //x=18.985 //y=2.96 //x2=22.825 //y2=3.7
cc_1116 ( QN N_noxref_9_c_1849_n ) capacitor c=0.024198f //x=18.87 //y=2.59 \
 //x2=22.825 //y2=3.7
cc_1117 ( N_QN_c_1494_n N_noxref_9_c_1849_n ) capacitor c=0.0111288f \
 //x=18.305 //y=5.2 //x2=22.825 //y2=3.7
cc_1118 ( N_QN_c_1498_n N_noxref_9_c_1849_n ) capacitor c=0.0099085f \
 //x=17.595 //y=5.2 //x2=22.825 //y2=3.7
cc_1119 ( N_QN_c_1478_n N_noxref_9_c_1849_n ) capacitor c=0.0245091f //x=20.72 \
 //y=2.08 //x2=22.825 //y2=3.7
cc_1120 ( N_QN_c_1510_n N_noxref_9_c_1849_n ) capacitor c=0.0129605f \
 //x=20.995 //y=4.79 //x2=22.825 //y2=3.7
cc_1121 ( QN N_noxref_9_c_1853_n ) capacitor c=3.49822e-19 //x=18.87 //y=2.59 \
 //x2=15.54 //y2=3.7
cc_1122 ( N_QN_c_1478_n N_noxref_9_c_1854_n ) capacitor c=0.00143759f \
 //x=20.72 //y=2.08 //x2=22.94 //y2=2.08
cc_1123 ( N_QN_c_1475_n N_noxref_10_c_2170_n ) capacitor c=0.174207f \
 //x=20.605 //y=2.96 //x2=23.565 //y2=3.33
cc_1124 ( N_QN_c_1531_p N_noxref_10_c_2170_n ) capacitor c=0.0293964f \
 //x=18.985 //y=2.96 //x2=23.565 //y2=3.33
cc_1125 ( QN N_noxref_10_c_2170_n ) capacitor c=0.0206038f //x=18.87 //y=2.59 \
 //x2=23.565 //y2=3.33
cc_1126 ( N_QN_c_1478_n N_noxref_10_c_2170_n ) capacitor c=0.0216152f \
 //x=20.72 //y=2.08 //x2=23.565 //y2=3.33
cc_1127 ( QN N_noxref_10_c_2213_n ) capacitor c=0.00179385f //x=18.87 //y=2.59 \
 //x2=18.245 //y2=3.33
cc_1128 ( QN N_noxref_10_c_2214_n ) capacitor c=0.0101115f //x=18.87 //y=2.59 \
 //x2=18.13 //y2=4.535
cc_1129 ( N_QN_c_1494_n N_noxref_10_c_2214_n ) capacitor c=0.0131484f \
 //x=18.305 //y=5.2 //x2=18.13 //y2=4.535
cc_1130 ( N_QN_c_1531_p N_noxref_10_c_2172_n ) capacitor c=0.00720056f \
 //x=18.985 //y=2.96 //x2=18.13 //y2=2.08
cc_1131 ( QN N_noxref_10_c_2172_n ) capacitor c=0.0734318f //x=18.87 //y=2.59 \
 //x2=18.13 //y2=2.08
cc_1132 ( N_QN_c_1478_n N_noxref_10_c_2172_n ) capacitor c=0.00101891f \
 //x=20.72 //y=2.08 //x2=18.13 //y2=2.08
cc_1133 ( N_QN_M40_noxref_g N_noxref_10_c_2179_n ) capacitor c=0.0186539f \
 //x=21.36 //y=6.02 //x2=21.935 //y2=5.155
cc_1134 ( QN N_noxref_10_c_2183_n ) capacitor c=2.97874e-19 //x=18.87 //y=2.59 \
 //x2=21.225 //y2=5.155
cc_1135 ( N_QN_M39_noxref_g N_noxref_10_c_2183_n ) capacitor c=0.0213876f \
 //x=20.92 //y=6.02 //x2=21.225 //y2=5.155
cc_1136 ( N_QN_c_1540_p N_noxref_10_c_2183_n ) capacitor c=0.0044314f \
 //x=21.285 //y=4.79 //x2=21.225 //y2=5.155
cc_1137 ( N_QN_c_1494_n N_noxref_10_M37_noxref_g ) capacitor c=0.0166421f \
 //x=18.305 //y=5.2 //x2=18.17 //y2=6.02
cc_1138 ( N_QN_M37_noxref_d N_noxref_10_M37_noxref_g ) capacitor c=0.0173476f \
 //x=18.245 //y=5.02 //x2=18.17 //y2=6.02
cc_1139 ( N_QN_c_1500_n N_noxref_10_M38_noxref_g ) capacitor c=0.0206783f \
 //x=18.785 //y=5.2 //x2=18.61 //y2=6.02
cc_1140 ( N_QN_M37_noxref_d N_noxref_10_M38_noxref_g ) capacitor c=0.0179769f \
 //x=18.245 //y=5.02 //x2=18.61 //y2=6.02
cc_1141 ( N_QN_M11_noxref_d N_noxref_10_c_2222_n ) capacitor c=0.00217566f \
 //x=18.24 //y=0.905 //x2=18.165 //y2=0.905
cc_1142 ( N_QN_M11_noxref_d N_noxref_10_c_2225_n ) capacitor c=0.0034598f \
 //x=18.24 //y=0.905 //x2=18.165 //y2=1.25
cc_1143 ( N_QN_M11_noxref_d N_noxref_10_c_2227_n ) capacitor c=0.00669531f \
 //x=18.24 //y=0.905 //x2=18.165 //y2=1.56
cc_1144 ( QN N_noxref_10_c_2257_n ) capacitor c=0.0142673f //x=18.87 //y=2.59 \
 //x2=18.535 //y2=4.79
cc_1145 ( N_QN_c_1589_p N_noxref_10_c_2257_n ) capacitor c=0.00421574f \
 //x=18.39 //y=5.2 //x2=18.535 //y2=4.79
cc_1146 ( N_QN_M11_noxref_d N_noxref_10_c_2259_n ) capacitor c=0.00241102f \
 //x=18.24 //y=0.905 //x2=18.54 //y2=0.75
cc_1147 ( N_QN_c_1477_n N_noxref_10_c_2260_n ) capacitor c=0.00371277f \
 //x=18.785 //y=1.655 //x2=18.54 //y2=1.405
cc_1148 ( N_QN_M11_noxref_d N_noxref_10_c_2260_n ) capacitor c=0.0137169f \
 //x=18.24 //y=0.905 //x2=18.54 //y2=1.405
cc_1149 ( N_QN_M11_noxref_d N_noxref_10_c_2230_n ) capacitor c=0.00132245f \
 //x=18.24 //y=0.905 //x2=18.695 //y2=0.905
cc_1150 ( N_QN_c_1477_n N_noxref_10_c_2231_n ) capacitor c=0.00457401f \
 //x=18.785 //y=1.655 //x2=18.695 //y2=1.25
cc_1151 ( N_QN_M11_noxref_d N_noxref_10_c_2231_n ) capacitor c=0.00566463f \
 //x=18.24 //y=0.905 //x2=18.695 //y2=1.25
cc_1152 ( QN N_noxref_10_c_2232_n ) capacitor c=0.00709342f //x=18.87 //y=2.59 \
 //x2=18.13 //y2=2.08
cc_1153 ( QN N_noxref_10_c_2266_n ) capacitor c=0.00306024f //x=18.87 //y=2.59 \
 //x2=18.13 //y2=1.915
cc_1154 ( N_QN_M11_noxref_d N_noxref_10_c_2266_n ) capacitor c=0.00660593f \
 //x=18.24 //y=0.905 //x2=18.13 //y2=1.915
cc_1155 ( QN N_noxref_10_c_2234_n ) capacitor c=0.00533692f //x=18.87 //y=2.59 \
 //x2=18.16 //y2=4.7
cc_1156 ( N_QN_c_1494_n N_noxref_10_c_2234_n ) capacitor c=0.00345427f \
 //x=18.305 //y=5.2 //x2=18.16 //y2=4.7
cc_1157 ( N_QN_M40_noxref_g N_noxref_10_M39_noxref_d ) capacitor c=0.0180032f \
 //x=21.36 //y=6.02 //x2=20.995 //y2=5.02
cc_1158 ( N_QN_c_1533_p N_noxref_18_c_2728_n ) capacitor c=3.15806e-19 \
 //x=18.515 //y=1.655 //x2=16.975 //y2=1.495
cc_1159 ( N_QN_c_1533_p N_noxref_18_c_2716_n ) capacitor c=0.0203424f \
 //x=18.515 //y=1.655 //x2=17.945 //y2=1.495
cc_1160 ( N_QN_c_1477_n N_noxref_18_c_2717_n ) capacitor c=0.00457164f \
 //x=18.785 //y=1.655 //x2=18.83 //y2=0.53
cc_1161 ( N_QN_M11_noxref_d N_noxref_18_c_2717_n ) capacitor c=0.0115831f \
 //x=18.24 //y=0.905 //x2=18.83 //y2=0.53
cc_1162 ( N_QN_c_1477_n N_noxref_18_M10_noxref_s ) capacitor c=0.013435f \
 //x=18.785 //y=1.655 //x2=16.84 //y2=0.365
cc_1163 ( N_QN_M11_noxref_d N_noxref_18_M10_noxref_s ) capacitor c=0.043966f \
 //x=18.24 //y=0.905 //x2=16.84 //y2=0.365
cc_1164 ( N_QN_c_1477_n N_noxref_19_c_2775_n ) capacitor c=4.08644e-19 \
 //x=18.785 //y=1.655 //x2=20.2 //y2=1.505
cc_1165 ( N_QN_c_1483_n N_noxref_19_c_2775_n ) capacitor c=0.0034165f \
 //x=20.42 //y=1.915 //x2=20.2 //y2=1.505
cc_1166 ( N_QN_c_1478_n N_noxref_19_c_2761_n ) capacitor c=0.0115578f \
 //x=20.72 //y=2.08 //x2=21.085 //y2=1.59
cc_1167 ( N_QN_c_1482_n N_noxref_19_c_2761_n ) capacitor c=0.00697148f \
 //x=20.42 //y=1.53 //x2=21.085 //y2=1.59
cc_1168 ( N_QN_c_1483_n N_noxref_19_c_2761_n ) capacitor c=0.0204849f \
 //x=20.42 //y=1.915 //x2=21.085 //y2=1.59
cc_1169 ( N_QN_c_1485_n N_noxref_19_c_2761_n ) capacitor c=0.00610316f \
 //x=20.795 //y=1.375 //x2=21.085 //y2=1.59
cc_1170 ( N_QN_c_1488_n N_noxref_19_c_2761_n ) capacitor c=0.00698822f \
 //x=20.95 //y=1.22 //x2=21.085 //y2=1.59
cc_1171 ( N_QN_c_1479_n N_noxref_19_M12_noxref_s ) capacitor c=0.0327271f \
 //x=20.42 //y=0.875 //x2=20.065 //y2=0.375
cc_1172 ( N_QN_c_1482_n N_noxref_19_M12_noxref_s ) capacitor c=7.99997e-19 \
 //x=20.42 //y=1.53 //x2=20.065 //y2=0.375
cc_1173 ( N_QN_c_1483_n N_noxref_19_M12_noxref_s ) capacitor c=0.00122123f \
 //x=20.42 //y=1.915 //x2=20.065 //y2=0.375
cc_1174 ( N_QN_c_1486_n N_noxref_19_M12_noxref_s ) capacitor c=0.0121427f \
 //x=20.95 //y=0.875 //x2=20.065 //y2=0.375
cc_1175 ( N_QN_M11_noxref_d N_noxref_19_M12_noxref_s ) capacitor c=2.53688e-19 \
 //x=18.24 //y=0.905 //x2=20.065 //y2=0.375
cc_1176 ( N_SN_c_1620_n N_noxref_9_c_1846_n ) capacitor c=0.0185443f \
 //x=21.715 //y=2.22 //x2=11.355 //y2=3.7
cc_1177 ( N_SN_c_1630_n N_noxref_9_c_1846_n ) capacitor c=0.00502941f \
 //x=10.475 //y=2.22 //x2=11.355 //y2=3.7
cc_1178 ( N_SN_c_1631_n N_noxref_9_c_1846_n ) capacitor c=0.0239078f //x=10.36 \
 //y=2.08 //x2=11.355 //y2=3.7
cc_1179 ( N_SN_c_1620_n N_noxref_9_c_1848_n ) capacitor c=0.0402118f \
 //x=21.715 //y=2.22 //x2=15.425 //y2=3.7
cc_1180 ( N_SN_c_1620_n N_noxref_9_c_1912_n ) capacitor c=0.00450155f \
 //x=21.715 //y=2.22 //x2=11.585 //y2=3.7
cc_1181 ( N_SN_c_1631_n N_noxref_9_c_1912_n ) capacitor c=0.00128547f \
 //x=10.36 //y=2.08 //x2=11.585 //y2=3.7
cc_1182 ( N_SN_c_1620_n N_noxref_9_c_1849_n ) capacitor c=0.0604652f \
 //x=21.715 //y=2.22 //x2=22.825 //y2=3.7
cc_1183 ( N_SN_c_1632_n N_noxref_9_c_1849_n ) capacitor c=0.0250454f //x=21.83 \
 //y=2.08 //x2=22.825 //y2=3.7
cc_1184 ( N_SN_c_1730_p N_noxref_9_c_1849_n ) capacitor c=0.00535612f \
 //x=22.165 //y=4.79 //x2=22.825 //y2=3.7
cc_1185 ( N_SN_c_1719_n N_noxref_9_c_1849_n ) capacitor c=0.00138305f \
 //x=21.83 //y=4.7 //x2=22.825 //y2=3.7
cc_1186 ( N_SN_c_1620_n N_noxref_9_c_1949_n ) capacitor c=0.00445687f \
 //x=21.715 //y=2.22 //x2=15.655 //y2=3.7
cc_1187 ( N_SN_c_1620_n N_noxref_9_c_1851_n ) capacitor c=0.0234959f \
 //x=21.715 //y=2.22 //x2=11.47 //y2=2.08
cc_1188 ( N_SN_c_1630_n N_noxref_9_c_1851_n ) capacitor c=0.00165648f \
 //x=10.475 //y=2.22 //x2=11.47 //y2=2.08
cc_1189 ( N_SN_c_1631_n N_noxref_9_c_1851_n ) capacitor c=0.0480841f //x=10.36 \
 //y=2.08 //x2=11.47 //y2=2.08
cc_1190 ( N_SN_c_1663_n N_noxref_9_c_1851_n ) capacitor c=0.00205895f \
 //x=10.45 //y=1.915 //x2=11.47 //y2=2.08
cc_1191 ( N_SN_c_1665_n N_noxref_9_c_1851_n ) capacitor c=0.00142741f \
 //x=10.36 //y=4.7 //x2=11.47 //y2=2.08
cc_1192 ( N_SN_c_1620_n N_noxref_9_c_2065_n ) capacitor c=0.0146822f \
 //x=21.715 //y=2.22 //x2=15.185 //y2=1.655
cc_1193 ( N_SN_c_1620_n N_noxref_9_c_1853_n ) capacitor c=0.0247812f \
 //x=21.715 //y=2.22 //x2=15.54 //y2=3.7
cc_1194 ( N_SN_c_1620_n N_noxref_9_c_1854_n ) capacitor c=0.00558344f \
 //x=21.715 //y=2.22 //x2=22.94 //y2=2.08
cc_1195 ( N_SN_c_1632_n N_noxref_9_c_1854_n ) capacitor c=0.0512968f //x=21.83 \
 //y=2.08 //x2=22.94 //y2=2.08
cc_1196 ( N_SN_c_1717_n N_noxref_9_c_1854_n ) capacitor c=0.00213841f \
 //x=21.92 //y=1.915 //x2=22.94 //y2=2.08
cc_1197 ( N_SN_c_1719_n N_noxref_9_c_1854_n ) capacitor c=0.00142741f \
 //x=21.83 //y=4.7 //x2=22.94 //y2=2.08
cc_1198 ( N_SN_M27_noxref_g N_noxref_9_M29_noxref_g ) capacitor c=0.0101598f \
 //x=10.33 //y=6.02 //x2=11.21 //y2=6.02
cc_1199 ( N_SN_M28_noxref_g N_noxref_9_M29_noxref_g ) capacitor c=0.0602553f \
 //x=10.77 //y=6.02 //x2=11.21 //y2=6.02
cc_1200 ( N_SN_M28_noxref_g N_noxref_9_M30_noxref_g ) capacitor c=0.0101598f \
 //x=10.77 //y=6.02 //x2=11.65 //y2=6.02
cc_1201 ( N_SN_M41_noxref_g N_noxref_9_M43_noxref_g ) capacitor c=0.0101598f \
 //x=21.8 //y=6.02 //x2=22.68 //y2=6.02
cc_1202 ( N_SN_M42_noxref_g N_noxref_9_M43_noxref_g ) capacitor c=0.0602553f \
 //x=22.24 //y=6.02 //x2=22.68 //y2=6.02
cc_1203 ( N_SN_M42_noxref_g N_noxref_9_M44_noxref_g ) capacitor c=0.0101598f \
 //x=22.24 //y=6.02 //x2=23.12 //y2=6.02
cc_1204 ( N_SN_c_1660_n N_noxref_9_c_1927_n ) capacitor c=0.00456962f \
 //x=10.45 //y=0.91 //x2=11.46 //y2=0.915
cc_1205 ( N_SN_c_1661_n N_noxref_9_c_1928_n ) capacitor c=0.00438372f \
 //x=10.45 //y=1.22 //x2=11.46 //y2=1.26
cc_1206 ( N_SN_c_1662_n N_noxref_9_c_1929_n ) capacitor c=0.00438372f \
 //x=10.45 //y=1.45 //x2=11.46 //y2=1.57
cc_1207 ( N_SN_c_1620_n N_noxref_9_c_1931_n ) capacitor c=3.13485e-19 \
 //x=21.715 //y=2.22 //x2=11.835 //y2=1.415
cc_1208 ( N_SN_c_1714_n N_noxref_9_c_2081_n ) capacitor c=0.00456962f \
 //x=21.92 //y=0.91 //x2=22.93 //y2=0.915
cc_1209 ( N_SN_c_1715_n N_noxref_9_c_2082_n ) capacitor c=0.00438372f \
 //x=21.92 //y=1.22 //x2=22.93 //y2=1.26
cc_1210 ( N_SN_c_1716_n N_noxref_9_c_2083_n ) capacitor c=0.00438372f \
 //x=21.92 //y=1.45 //x2=22.93 //y2=1.57
cc_1211 ( N_SN_c_1620_n N_noxref_9_c_1936_n ) capacitor c=0.00581478f \
 //x=21.715 //y=2.22 //x2=11.47 //y2=2.08
cc_1212 ( N_SN_c_1630_n N_noxref_9_c_1936_n ) capacitor c=2.3323e-19 \
 //x=10.475 //y=2.22 //x2=11.47 //y2=2.08
cc_1213 ( N_SN_c_1631_n N_noxref_9_c_1936_n ) capacitor c=0.0019893f //x=10.36 \
 //y=2.08 //x2=11.47 //y2=2.08
cc_1214 ( N_SN_c_1663_n N_noxref_9_c_1936_n ) capacitor c=0.00828003f \
 //x=10.45 //y=1.915 //x2=11.47 //y2=2.08
cc_1215 ( N_SN_c_1663_n N_noxref_9_c_1937_n ) capacitor c=0.00438372f \
 //x=10.45 //y=1.915 //x2=11.47 //y2=1.915
cc_1216 ( N_SN_c_1631_n N_noxref_9_c_1939_n ) capacitor c=0.00219458f \
 //x=10.36 //y=2.08 //x2=11.47 //y2=4.7
cc_1217 ( N_SN_c_1680_n N_noxref_9_c_1939_n ) capacitor c=0.0611812f \
 //x=10.695 //y=4.79 //x2=11.47 //y2=4.7
cc_1218 ( N_SN_c_1665_n N_noxref_9_c_1939_n ) capacitor c=0.00487508f \
 //x=10.36 //y=4.7 //x2=11.47 //y2=4.7
cc_1219 ( N_SN_c_1620_n N_noxref_9_c_2092_n ) capacitor c=0.00341397f \
 //x=21.715 //y=2.22 //x2=22.94 //y2=2.08
cc_1220 ( N_SN_c_1632_n N_noxref_9_c_2092_n ) capacitor c=0.0021852f //x=21.83 \
 //y=2.08 //x2=22.94 //y2=2.08
cc_1221 ( N_SN_c_1717_n N_noxref_9_c_2092_n ) capacitor c=0.00896806f \
 //x=21.92 //y=1.915 //x2=22.94 //y2=2.08
cc_1222 ( N_SN_c_1717_n N_noxref_9_c_2095_n ) capacitor c=0.00438372f \
 //x=21.92 //y=1.915 //x2=22.94 //y2=1.915
cc_1223 ( N_SN_c_1632_n N_noxref_9_c_2096_n ) capacitor c=0.00219458f \
 //x=21.83 //y=2.08 //x2=22.94 //y2=4.7
cc_1224 ( N_SN_c_1730_p N_noxref_9_c_2096_n ) capacitor c=0.0611812f \
 //x=22.165 //y=4.79 //x2=22.94 //y2=4.7
cc_1225 ( N_SN_c_1719_n N_noxref_9_c_2096_n ) capacitor c=0.00487508f \
 //x=21.83 //y=4.7 //x2=22.94 //y2=4.7
cc_1226 ( N_SN_c_1620_n N_noxref_10_c_2170_n ) capacitor c=0.0553978f \
 //x=21.715 //y=2.22 //x2=23.565 //y2=3.33
cc_1227 ( N_SN_c_1632_n N_noxref_10_c_2170_n ) capacitor c=0.0229939f \
 //x=21.83 //y=2.08 //x2=23.565 //y2=3.33
cc_1228 ( N_SN_c_1620_n N_noxref_10_c_2213_n ) capacitor c=0.00751102f \
 //x=21.715 //y=2.22 //x2=18.245 //y2=3.33
cc_1229 ( N_SN_c_1620_n N_noxref_10_c_2172_n ) capacitor c=0.0218045f \
 //x=21.715 //y=2.22 //x2=18.13 //y2=2.08
cc_1230 ( N_SN_c_1632_n N_noxref_10_c_2179_n ) capacitor c=0.0149705f \
 //x=21.83 //y=2.08 //x2=21.935 //y2=5.155
cc_1231 ( N_SN_M41_noxref_g N_noxref_10_c_2179_n ) capacitor c=0.0167692f \
 //x=21.8 //y=6.02 //x2=21.935 //y2=5.155
cc_1232 ( N_SN_c_1719_n N_noxref_10_c_2179_n ) capacitor c=0.00325274f \
 //x=21.83 //y=4.7 //x2=21.935 //y2=5.155
cc_1233 ( N_SN_M42_noxref_g N_noxref_10_c_2185_n ) capacitor c=0.019179f \
 //x=22.24 //y=6.02 //x2=22.815 //y2=5.155
cc_1234 ( N_SN_c_1632_n N_noxref_10_c_2193_n ) capacitor c=0.00363599f \
 //x=21.83 //y=2.08 //x2=23.68 //y2=3.33
cc_1235 ( N_SN_c_1730_p N_noxref_10_c_2280_n ) capacitor c=0.00441288f \
 //x=22.165 //y=4.79 //x2=22.02 //y2=5.155
cc_1236 ( N_SN_c_1620_n N_noxref_10_c_2260_n ) capacitor c=3.11115e-19 \
 //x=21.715 //y=2.22 //x2=18.54 //y2=1.405
cc_1237 ( N_SN_c_1620_n N_noxref_10_c_2232_n ) capacitor c=0.00570196f \
 //x=21.715 //y=2.22 //x2=18.13 //y2=2.08
cc_1238 ( N_SN_M41_noxref_g N_noxref_10_M41_noxref_d ) capacitor c=0.0180032f \
 //x=21.8 //y=6.02 //x2=21.875 //y2=5.02
cc_1239 ( N_SN_M42_noxref_g N_noxref_10_M41_noxref_d ) capacitor c=0.0180032f \
 //x=22.24 //y=6.02 //x2=21.875 //y2=5.02
cc_1240 ( N_SN_c_1655_n N_noxref_15_c_2557_n ) capacitor c=0.0167228f \
 //x=9.925 //y=0.91 //x2=10.585 //y2=0.54
cc_1241 ( N_SN_c_1660_n N_noxref_15_c_2557_n ) capacitor c=0.00534519f \
 //x=10.45 //y=0.91 //x2=10.585 //y2=0.54
cc_1242 ( N_SN_c_1620_n N_noxref_15_c_2583_n ) capacitor c=0.00387656f \
 //x=21.715 //y=2.22 //x2=10.585 //y2=1.59
cc_1243 ( N_SN_c_1630_n N_noxref_15_c_2583_n ) capacitor c=0.00354473f \
 //x=10.475 //y=2.22 //x2=10.585 //y2=1.59
cc_1244 ( N_SN_c_1631_n N_noxref_15_c_2583_n ) capacitor c=0.0119919f \
 //x=10.36 //y=2.08 //x2=10.585 //y2=1.59
cc_1245 ( N_SN_c_1658_n N_noxref_15_c_2583_n ) capacitor c=0.0153695f \
 //x=9.925 //y=1.22 //x2=10.585 //y2=1.59
cc_1246 ( N_SN_c_1663_n N_noxref_15_c_2583_n ) capacitor c=0.0213278f \
 //x=10.45 //y=1.915 //x2=10.585 //y2=1.59
cc_1247 ( N_SN_c_1620_n N_noxref_15_M5_noxref_s ) capacitor c=0.00599513f \
 //x=21.715 //y=2.22 //x2=8.595 //y2=0.375
cc_1248 ( N_SN_c_1655_n N_noxref_15_M5_noxref_s ) capacitor c=0.00798959f \
 //x=9.925 //y=0.91 //x2=8.595 //y2=0.375
cc_1249 ( N_SN_c_1662_n N_noxref_15_M5_noxref_s ) capacitor c=0.00212176f \
 //x=10.45 //y=1.45 //x2=8.595 //y2=0.375
cc_1250 ( N_SN_c_1663_n N_noxref_15_M5_noxref_s ) capacitor c=0.00298115f \
 //x=10.45 //y=1.915 //x2=8.595 //y2=0.375
cc_1251 ( N_SN_c_1620_n N_noxref_16_c_2604_n ) capacitor c=0.00657782f \
 //x=21.715 //y=2.22 //x2=11.155 //y2=0.995
cc_1252 ( N_SN_c_1798_p N_noxref_16_c_2604_n ) capacitor c=2.14837e-19 \
 //x=10.295 //y=0.755 //x2=11.155 //y2=0.995
cc_1253 ( N_SN_c_1660_n N_noxref_16_c_2604_n ) capacitor c=0.00123426f \
 //x=10.45 //y=0.91 //x2=11.155 //y2=0.995
cc_1254 ( N_SN_c_1661_n N_noxref_16_c_2604_n ) capacitor c=0.0129288f \
 //x=10.45 //y=1.22 //x2=11.155 //y2=0.995
cc_1255 ( N_SN_c_1662_n N_noxref_16_c_2604_n ) capacitor c=0.00142359f \
 //x=10.45 //y=1.45 //x2=11.155 //y2=0.995
cc_1256 ( N_SN_c_1620_n N_noxref_16_c_2609_n ) capacitor c=0.00147946f \
 //x=21.715 //y=2.22 //x2=12.125 //y2=0.54
cc_1257 ( N_SN_c_1655_n N_noxref_16_M6_noxref_d ) capacitor c=0.00223875f \
 //x=9.925 //y=0.91 //x2=10 //y2=0.91
cc_1258 ( N_SN_c_1658_n N_noxref_16_M6_noxref_d ) capacitor c=0.00262485f \
 //x=9.925 //y=1.22 //x2=10 //y2=0.91
cc_1259 ( N_SN_c_1798_p N_noxref_16_M6_noxref_d ) capacitor c=0.00220746f \
 //x=10.295 //y=0.755 //x2=10 //y2=0.91
cc_1260 ( N_SN_c_1806_p N_noxref_16_M6_noxref_d ) capacitor c=0.00194798f \
 //x=10.295 //y=1.375 //x2=10 //y2=0.91
cc_1261 ( N_SN_c_1660_n N_noxref_16_M6_noxref_d ) capacitor c=0.00198465f \
 //x=10.45 //y=0.91 //x2=10 //y2=0.91
cc_1262 ( N_SN_c_1661_n N_noxref_16_M6_noxref_d ) capacitor c=0.00128384f \
 //x=10.45 //y=1.22 //x2=10 //y2=0.91
cc_1263 ( N_SN_c_1620_n N_noxref_16_M7_noxref_s ) capacitor c=0.00642985f \
 //x=21.715 //y=2.22 //x2=11.105 //y2=0.375
cc_1264 ( N_SN_c_1660_n N_noxref_16_M7_noxref_s ) capacitor c=7.21316e-19 \
 //x=10.45 //y=0.91 //x2=11.105 //y2=0.375
cc_1265 ( N_SN_c_1661_n N_noxref_16_M7_noxref_s ) capacitor c=0.00348171f \
 //x=10.45 //y=1.22 //x2=11.105 //y2=0.375
cc_1266 ( N_SN_c_1620_n N_noxref_17_c_2676_n ) capacitor c=0.00635755f \
 //x=21.715 //y=2.22 //x2=13.645 //y2=1.495
cc_1267 ( N_SN_c_1620_n N_noxref_17_c_2657_n ) capacitor c=0.0223494f \
 //x=21.715 //y=2.22 //x2=14.53 //y2=1.58
cc_1268 ( N_SN_c_1620_n N_noxref_17_c_2664_n ) capacitor c=0.00649228f \
 //x=21.715 //y=2.22 //x2=14.615 //y2=1.495
cc_1269 ( N_SN_c_1620_n N_noxref_17_c_2665_n ) capacitor c=0.00178534f \
 //x=21.715 //y=2.22 //x2=15.5 //y2=0.53
cc_1270 ( N_SN_c_1620_n N_noxref_17_M8_noxref_s ) capacitor c=0.00113237f \
 //x=21.715 //y=2.22 //x2=13.51 //y2=0.365
cc_1271 ( N_SN_c_1620_n N_noxref_18_c_2728_n ) capacitor c=0.00635755f \
 //x=21.715 //y=2.22 //x2=16.975 //y2=1.495
cc_1272 ( N_SN_c_1620_n N_noxref_18_c_2709_n ) capacitor c=0.0223494f \
 //x=21.715 //y=2.22 //x2=17.86 //y2=1.58
cc_1273 ( N_SN_c_1620_n N_noxref_18_c_2716_n ) capacitor c=0.00649228f \
 //x=21.715 //y=2.22 //x2=17.945 //y2=1.495
cc_1274 ( N_SN_c_1620_n N_noxref_18_c_2717_n ) capacitor c=0.00178534f \
 //x=21.715 //y=2.22 //x2=18.83 //y2=0.53
cc_1275 ( N_SN_c_1620_n N_noxref_18_M10_noxref_s ) capacitor c=0.00113237f \
 //x=21.715 //y=2.22 //x2=16.84 //y2=0.365
cc_1276 ( N_SN_c_1620_n N_noxref_19_c_2775_n ) capacitor c=0.00642985f \
 //x=21.715 //y=2.22 //x2=20.2 //y2=1.505
cc_1277 ( N_SN_c_1620_n N_noxref_19_c_2761_n ) capacitor c=0.0225733f \
 //x=21.715 //y=2.22 //x2=21.085 //y2=1.59
cc_1278 ( N_SN_c_1709_n N_noxref_19_c_2768_n ) capacitor c=0.0167228f \
 //x=21.395 //y=0.91 //x2=22.055 //y2=0.54
cc_1279 ( N_SN_c_1714_n N_noxref_19_c_2768_n ) capacitor c=0.00534519f \
 //x=21.92 //y=0.91 //x2=22.055 //y2=0.54
cc_1280 ( N_SN_c_1620_n N_noxref_19_c_2791_n ) capacitor c=0.0178105f \
 //x=21.715 //y=2.22 //x2=22.055 //y2=1.59
cc_1281 ( N_SN_c_1632_n N_noxref_19_c_2791_n ) capacitor c=0.0119919f \
 //x=21.83 //y=2.08 //x2=22.055 //y2=1.59
cc_1282 ( N_SN_c_1712_n N_noxref_19_c_2791_n ) capacitor c=0.0157358f \
 //x=21.395 //y=1.22 //x2=22.055 //y2=1.59
cc_1283 ( N_SN_c_1717_n N_noxref_19_c_2791_n ) capacitor c=0.0216647f \
 //x=21.92 //y=1.915 //x2=22.055 //y2=1.59
cc_1284 ( N_SN_c_1620_n N_noxref_19_M12_noxref_s ) capacitor c=0.00642985f \
 //x=21.715 //y=2.22 //x2=20.065 //y2=0.375
cc_1285 ( N_SN_c_1709_n N_noxref_19_M12_noxref_s ) capacitor c=0.00798959f \
 //x=21.395 //y=0.91 //x2=20.065 //y2=0.375
cc_1286 ( N_SN_c_1716_n N_noxref_19_M12_noxref_s ) capacitor c=0.00212176f \
 //x=21.92 //y=1.45 //x2=20.065 //y2=0.375
cc_1287 ( N_SN_c_1717_n N_noxref_19_M12_noxref_s ) capacitor c=0.00298115f \
 //x=21.92 //y=1.915 //x2=20.065 //y2=0.375
cc_1288 ( N_SN_c_1834_p N_noxref_20_c_2811_n ) capacitor c=2.14837e-19 \
 //x=21.765 //y=0.755 //x2=22.625 //y2=0.995
cc_1289 ( N_SN_c_1714_n N_noxref_20_c_2811_n ) capacitor c=0.00123426f \
 //x=21.92 //y=0.91 //x2=22.625 //y2=0.995
cc_1290 ( N_SN_c_1715_n N_noxref_20_c_2811_n ) capacitor c=0.0129288f \
 //x=21.92 //y=1.22 //x2=22.625 //y2=0.995
cc_1291 ( N_SN_c_1716_n N_noxref_20_c_2811_n ) capacitor c=0.00142359f \
 //x=21.92 //y=1.45 //x2=22.625 //y2=0.995
cc_1292 ( N_SN_c_1709_n N_noxref_20_M13_noxref_d ) capacitor c=0.00223875f \
 //x=21.395 //y=0.91 //x2=21.47 //y2=0.91
cc_1293 ( N_SN_c_1712_n N_noxref_20_M13_noxref_d ) capacitor c=0.00262485f \
 //x=21.395 //y=1.22 //x2=21.47 //y2=0.91
cc_1294 ( N_SN_c_1834_p N_noxref_20_M13_noxref_d ) capacitor c=0.00220746f \
 //x=21.765 //y=0.755 //x2=21.47 //y2=0.91
cc_1295 ( N_SN_c_1841_p N_noxref_20_M13_noxref_d ) capacitor c=0.00194798f \
 //x=21.765 //y=1.375 //x2=21.47 //y2=0.91
cc_1296 ( N_SN_c_1714_n N_noxref_20_M13_noxref_d ) capacitor c=0.00198465f \
 //x=21.92 //y=0.91 //x2=21.47 //y2=0.91
cc_1297 ( N_SN_c_1715_n N_noxref_20_M13_noxref_d ) capacitor c=0.00128384f \
 //x=21.92 //y=1.22 //x2=21.47 //y2=0.91
cc_1298 ( N_SN_c_1714_n N_noxref_20_M14_noxref_s ) capacitor c=7.21316e-19 \
 //x=21.92 //y=0.91 //x2=22.575 //y2=0.375
cc_1299 ( N_SN_c_1715_n N_noxref_20_M14_noxref_s ) capacitor c=0.00348171f \
 //x=21.92 //y=1.22 //x2=22.575 //y2=0.375
cc_1300 ( N_noxref_9_c_1849_n N_noxref_10_c_2170_n ) capacitor c=0.433921f \
 //x=22.825 //y=3.7 //x2=23.565 //y2=3.33
cc_1301 ( N_noxref_9_c_1854_n N_noxref_10_c_2170_n ) capacitor c=0.0269537f \
 //x=22.94 //y=2.08 //x2=23.565 //y2=3.33
cc_1302 ( N_noxref_9_c_1849_n N_noxref_10_c_2213_n ) capacitor c=0.0291821f \
 //x=22.825 //y=3.7 //x2=18.245 //y2=3.33
cc_1303 ( N_noxref_9_c_1849_n N_noxref_10_c_2214_n ) capacitor c=0.00113929f \
 //x=22.825 //y=3.7 //x2=18.13 //y2=4.535
cc_1304 ( N_noxref_9_c_1849_n N_noxref_10_c_2172_n ) capacitor c=0.0234812f \
 //x=22.825 //y=3.7 //x2=18.13 //y2=2.08
cc_1305 ( N_noxref_9_c_1853_n N_noxref_10_c_2172_n ) capacitor c=0.00118913f \
 //x=15.54 //y=3.7 //x2=18.13 //y2=2.08
cc_1306 ( N_noxref_9_c_1849_n N_noxref_10_c_2179_n ) capacitor c=0.0189263f \
 //x=22.825 //y=3.7 //x2=21.935 //y2=5.155
cc_1307 ( N_noxref_9_c_1849_n N_noxref_10_c_2183_n ) capacitor c=0.0135617f \
 //x=22.825 //y=3.7 //x2=21.225 //y2=5.155
cc_1308 ( N_noxref_9_M43_noxref_g N_noxref_10_c_2185_n ) capacitor c=0.019179f \
 //x=22.68 //y=6.02 //x2=22.815 //y2=5.155
cc_1309 ( N_noxref_9_c_1849_n N_noxref_10_c_2189_n ) capacitor c=0.00153992f \
 //x=22.825 //y=3.7 //x2=23.595 //y2=5.155
cc_1310 ( N_noxref_9_M44_noxref_g N_noxref_10_c_2189_n ) capacitor \
 c=0.0217141f //x=23.12 //y=6.02 //x2=23.595 //y2=5.155
cc_1311 ( N_noxref_9_c_2096_n N_noxref_10_c_2189_n ) capacitor c=0.00201851f \
 //x=22.94 //y=4.7 //x2=23.595 //y2=5.155
cc_1312 ( N_noxref_9_c_2111_p N_noxref_10_c_2174_n ) capacitor c=0.00359704f \
 //x=23.305 //y=1.415 //x2=23.595 //y2=1.665
cc_1313 ( N_noxref_9_c_2112_p N_noxref_10_c_2174_n ) capacitor c=0.00457401f \
 //x=23.46 //y=1.26 //x2=23.595 //y2=1.665
cc_1314 ( N_noxref_9_c_1849_n N_noxref_10_c_2193_n ) capacitor c=0.00599141f \
 //x=22.825 //y=3.7 //x2=23.68 //y2=3.33
cc_1315 ( N_noxref_9_c_1854_n N_noxref_10_c_2193_n ) capacitor c=0.0882467f \
 //x=22.94 //y=2.08 //x2=23.68 //y2=3.33
cc_1316 ( N_noxref_9_c_2092_n N_noxref_10_c_2193_n ) capacitor c=0.00772308f \
 //x=22.94 //y=2.08 //x2=23.68 //y2=3.33
cc_1317 ( N_noxref_9_c_2095_n N_noxref_10_c_2193_n ) capacitor c=0.00283672f \
 //x=22.94 //y=1.915 //x2=23.68 //y2=3.33
cc_1318 ( N_noxref_9_c_2096_n N_noxref_10_c_2193_n ) capacitor c=0.013844f \
 //x=22.94 //y=4.7 //x2=23.68 //y2=3.33
cc_1319 ( N_noxref_9_c_1849_n N_noxref_10_c_2304_n ) capacitor c=5.7529e-19 \
 //x=22.825 //y=3.7 //x2=22.9 //y2=5.155
cc_1320 ( N_noxref_9_c_1854_n N_noxref_10_c_2304_n ) capacitor c=0.017024f \
 //x=22.94 //y=2.08 //x2=22.9 //y2=5.155
cc_1321 ( N_noxref_9_c_2096_n N_noxref_10_c_2304_n ) capacitor c=0.00476349f \
 //x=22.94 //y=4.7 //x2=22.9 //y2=5.155
cc_1322 ( N_noxref_9_c_1849_n N_noxref_10_c_2257_n ) capacitor c=0.00624857f \
 //x=22.825 //y=3.7 //x2=18.535 //y2=4.79
cc_1323 ( N_noxref_9_c_1849_n N_noxref_10_c_2234_n ) capacitor c=9.84146e-19 \
 //x=22.825 //y=3.7 //x2=18.16 //y2=4.7
cc_1324 ( N_noxref_9_c_2081_n N_noxref_10_M14_noxref_d ) capacitor \
 c=0.00217566f //x=22.93 //y=0.915 //x2=23.005 //y2=0.915
cc_1325 ( N_noxref_9_c_2082_n N_noxref_10_M14_noxref_d ) capacitor \
 c=0.0034598f //x=22.93 //y=1.26 //x2=23.005 //y2=0.915
cc_1326 ( N_noxref_9_c_2083_n N_noxref_10_M14_noxref_d ) capacitor \
 c=0.00544291f //x=22.93 //y=1.57 //x2=23.005 //y2=0.915
cc_1327 ( N_noxref_9_c_2126_p N_noxref_10_M14_noxref_d ) capacitor \
 c=0.00241102f //x=23.305 //y=0.76 //x2=23.005 //y2=0.915
cc_1328 ( N_noxref_9_c_2111_p N_noxref_10_M14_noxref_d ) capacitor \
 c=0.0140297f //x=23.305 //y=1.415 //x2=23.005 //y2=0.915
cc_1329 ( N_noxref_9_c_2128_p N_noxref_10_M14_noxref_d ) capacitor \
 c=0.00219619f //x=23.46 //y=0.915 //x2=23.005 //y2=0.915
cc_1330 ( N_noxref_9_c_2112_p N_noxref_10_M14_noxref_d ) capacitor \
 c=0.00603828f //x=23.46 //y=1.26 //x2=23.005 //y2=0.915
cc_1331 ( N_noxref_9_c_2095_n N_noxref_10_M14_noxref_d ) capacitor \
 c=0.00661782f //x=22.94 //y=1.915 //x2=23.005 //y2=0.915
cc_1332 ( N_noxref_9_M43_noxref_g N_noxref_10_M43_noxref_d ) capacitor \
 c=0.0180032f //x=22.68 //y=6.02 //x2=22.755 //y2=5.02
cc_1333 ( N_noxref_9_M44_noxref_g N_noxref_10_M43_noxref_d ) capacitor \
 c=0.0194246f //x=23.12 //y=6.02 //x2=22.755 //y2=5.02
cc_1334 ( N_noxref_9_c_1850_n N_noxref_14_c_2502_n ) capacitor c=0.0020642f \
 //x=6.66 //y=2.08 //x2=7.315 //y2=0.54
cc_1335 ( N_noxref_9_c_1976_n N_noxref_14_c_2502_n ) capacitor c=0.0194423f \
 //x=6.65 //y=0.915 //x2=7.315 //y2=0.54
cc_1336 ( N_noxref_9_c_2031_n N_noxref_14_c_2502_n ) capacitor c=0.00656458f \
 //x=7.18 //y=0.915 //x2=7.315 //y2=0.54
cc_1337 ( N_noxref_9_c_1907_n N_noxref_14_c_2502_n ) capacitor c=2.20712e-19 \
 //x=6.66 //y=2.08 //x2=7.315 //y2=0.54
cc_1338 ( N_noxref_9_c_1977_n N_noxref_14_c_2528_n ) capacitor c=0.00538033f \
 //x=6.65 //y=1.26 //x2=6.43 //y2=0.995
cc_1339 ( N_noxref_9_c_1976_n N_noxref_14_M4_noxref_s ) capacitor \
 c=0.00538033f //x=6.65 //y=0.915 //x2=6.295 //y2=0.375
cc_1340 ( N_noxref_9_c_1978_n N_noxref_14_M4_noxref_s ) capacitor \
 c=0.00538033f //x=6.65 //y=1.57 //x2=6.295 //y2=0.375
cc_1341 ( N_noxref_9_c_2031_n N_noxref_14_M4_noxref_s ) capacitor c=0.0143002f \
 //x=7.18 //y=0.915 //x2=6.295 //y2=0.375
cc_1342 ( N_noxref_9_c_2032_n N_noxref_14_M4_noxref_s ) capacitor \
 c=0.00290153f //x=7.18 //y=1.26 //x2=6.295 //y2=0.375
cc_1343 ( N_noxref_9_c_1846_n N_noxref_15_c_2550_n ) capacitor c=0.00208074f \
 //x=11.355 //y=3.7 //x2=9.615 //y2=1.59
cc_1344 ( N_noxref_9_c_1846_n N_noxref_15_c_2583_n ) capacitor c=0.00393278f \
 //x=11.355 //y=3.7 //x2=10.585 //y2=1.59
cc_1345 ( N_noxref_9_c_1846_n N_noxref_15_M5_noxref_s ) capacitor \
 c=0.00188576f //x=11.355 //y=3.7 //x2=8.595 //y2=0.375
cc_1346 ( N_noxref_9_c_1851_n N_noxref_16_c_2609_n ) capacitor c=0.00204385f \
 //x=11.47 //y=2.08 //x2=12.125 //y2=0.54
cc_1347 ( N_noxref_9_c_1927_n N_noxref_16_c_2609_n ) capacitor c=0.0194423f \
 //x=11.46 //y=0.915 //x2=12.125 //y2=0.54
cc_1348 ( N_noxref_9_c_1933_n N_noxref_16_c_2609_n ) capacitor c=0.00656458f \
 //x=11.99 //y=0.915 //x2=12.125 //y2=0.54
cc_1349 ( N_noxref_9_c_1936_n N_noxref_16_c_2609_n ) capacitor c=2.20712e-19 \
 //x=11.47 //y=2.08 //x2=12.125 //y2=0.54
cc_1350 ( N_noxref_9_c_1928_n N_noxref_16_c_2620_n ) capacitor c=0.00538829f \
 //x=11.46 //y=1.26 //x2=11.24 //y2=0.995
cc_1351 ( N_noxref_9_c_1927_n N_noxref_16_M7_noxref_s ) capacitor \
 c=0.00538829f //x=11.46 //y=0.915 //x2=11.105 //y2=0.375
cc_1352 ( N_noxref_9_c_1929_n N_noxref_16_M7_noxref_s ) capacitor \
 c=0.00538829f //x=11.46 //y=1.57 //x2=11.105 //y2=0.375
cc_1353 ( N_noxref_9_c_1933_n N_noxref_16_M7_noxref_s ) capacitor c=0.0143002f \
 //x=11.99 //y=0.915 //x2=11.105 //y2=0.375
cc_1354 ( N_noxref_9_c_1934_n N_noxref_16_M7_noxref_s ) capacitor \
 c=0.00290153f //x=11.99 //y=1.26 //x2=11.105 //y2=0.375
cc_1355 ( N_noxref_9_c_2065_n N_noxref_17_c_2676_n ) capacitor c=3.15806e-19 \
 //x=15.185 //y=1.655 //x2=13.645 //y2=1.495
cc_1356 ( N_noxref_9_c_2065_n N_noxref_17_c_2664_n ) capacitor c=0.020324f \
 //x=15.185 //y=1.655 //x2=14.615 //y2=1.495
cc_1357 ( N_noxref_9_c_1852_n N_noxref_17_c_2665_n ) capacitor c=0.00457164f \
 //x=15.455 //y=1.655 //x2=15.5 //y2=0.53
cc_1358 ( N_noxref_9_M9_noxref_d N_noxref_17_c_2665_n ) capacitor c=0.0115831f \
 //x=14.91 //y=0.905 //x2=15.5 //y2=0.53
cc_1359 ( N_noxref_9_c_1852_n N_noxref_17_M8_noxref_s ) capacitor c=0.013435f \
 //x=15.455 //y=1.655 //x2=13.51 //y2=0.365
cc_1360 ( N_noxref_9_M9_noxref_d N_noxref_17_M8_noxref_s ) capacitor \
 c=0.0439476f //x=14.91 //y=0.905 //x2=13.51 //y2=0.365
cc_1361 ( N_noxref_9_c_1852_n N_noxref_18_c_2728_n ) capacitor c=3.22188e-19 \
 //x=15.455 //y=1.655 //x2=16.975 //y2=1.495
cc_1362 ( N_noxref_9_c_1854_n N_noxref_20_c_2816_n ) capacitor c=0.00208576f \
 //x=22.94 //y=2.08 //x2=23.595 //y2=0.54
cc_1363 ( N_noxref_9_c_2081_n N_noxref_20_c_2816_n ) capacitor c=0.0194423f \
 //x=22.93 //y=0.915 //x2=23.595 //y2=0.54
cc_1364 ( N_noxref_9_c_2128_p N_noxref_20_c_2816_n ) capacitor c=0.00656458f \
 //x=23.46 //y=0.915 //x2=23.595 //y2=0.54
cc_1365 ( N_noxref_9_c_2092_n N_noxref_20_c_2816_n ) capacitor c=2.20712e-19 \
 //x=22.94 //y=2.08 //x2=23.595 //y2=0.54
cc_1366 ( N_noxref_9_c_2082_n N_noxref_20_c_2839_n ) capacitor c=0.00538829f \
 //x=22.93 //y=1.26 //x2=22.71 //y2=0.995
cc_1367 ( N_noxref_9_c_2081_n N_noxref_20_M14_noxref_s ) capacitor \
 c=0.00538829f //x=22.93 //y=0.915 //x2=22.575 //y2=0.375
cc_1368 ( N_noxref_9_c_2083_n N_noxref_20_M14_noxref_s ) capacitor \
 c=0.00538829f //x=22.93 //y=1.57 //x2=22.575 //y2=0.375
cc_1369 ( N_noxref_9_c_2128_p N_noxref_20_M14_noxref_s ) capacitor \
 c=0.0143002f //x=23.46 //y=0.915 //x2=22.575 //y2=0.375
cc_1370 ( N_noxref_9_c_2112_p N_noxref_20_M14_noxref_s ) capacitor \
 c=0.00290153f //x=23.46 //y=1.26 //x2=22.575 //y2=0.375
cc_1371 ( N_noxref_10_c_2227_n N_noxref_18_c_2716_n ) capacitor c=0.00623646f \
 //x=18.165 //y=1.56 //x2=17.945 //y2=1.495
cc_1372 ( N_noxref_10_c_2232_n N_noxref_18_c_2716_n ) capacitor c=0.00173579f \
 //x=18.13 //y=2.08 //x2=17.945 //y2=1.495
cc_1373 ( N_noxref_10_c_2172_n N_noxref_18_c_2717_n ) capacitor c=0.00156605f \
 //x=18.13 //y=2.08 //x2=18.83 //y2=0.53
cc_1374 ( N_noxref_10_c_2222_n N_noxref_18_c_2717_n ) capacitor c=0.0188655f \
 //x=18.165 //y=0.905 //x2=18.83 //y2=0.53
cc_1375 ( N_noxref_10_c_2230_n N_noxref_18_c_2717_n ) capacitor c=0.00656458f \
 //x=18.695 //y=0.905 //x2=18.83 //y2=0.53
cc_1376 ( N_noxref_10_c_2232_n N_noxref_18_c_2717_n ) capacitor c=2.1838e-19 \
 //x=18.13 //y=2.08 //x2=18.83 //y2=0.53
cc_1377 ( N_noxref_10_c_2222_n N_noxref_18_M10_noxref_s ) capacitor \
 c=0.00623646f //x=18.165 //y=0.905 //x2=16.84 //y2=0.365
cc_1378 ( N_noxref_10_c_2230_n N_noxref_18_M10_noxref_s ) capacitor \
 c=0.0143002f //x=18.695 //y=0.905 //x2=16.84 //y2=0.365
cc_1379 ( N_noxref_10_c_2231_n N_noxref_18_M10_noxref_s ) capacitor \
 c=0.00290153f //x=18.695 //y=1.25 //x2=16.84 //y2=0.365
cc_1380 ( N_noxref_10_c_2170_n N_noxref_19_c_2791_n ) capacitor c=0.00124665f \
 //x=23.565 //y=3.33 //x2=22.055 //y2=1.59
cc_1381 ( N_noxref_10_c_2170_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00227057f //x=23.565 //y=3.33 //x2=20.065 //y2=0.375
cc_1382 ( N_noxref_10_M14_noxref_d N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00309936f //x=23.005 //y=0.915 //x2=20.065 //y2=0.375
cc_1383 ( N_noxref_10_c_2170_n N_noxref_20_c_2811_n ) capacitor c=0.00306157f \
 //x=23.565 //y=3.33 //x2=22.625 //y2=0.995
cc_1384 ( N_noxref_10_c_2170_n N_noxref_20_c_2816_n ) capacitor c=5.19687e-19 \
 //x=23.565 //y=3.33 //x2=23.595 //y2=0.54
cc_1385 ( N_noxref_10_c_2174_n N_noxref_20_c_2816_n ) capacitor c=0.00466084f \
 //x=23.595 //y=1.665 //x2=23.595 //y2=0.54
cc_1386 ( N_noxref_10_M14_noxref_d N_noxref_20_c_2816_n ) capacitor \
 c=0.0117786f //x=23.005 //y=0.915 //x2=23.595 //y2=0.54
cc_1387 ( N_noxref_10_c_2335_p N_noxref_20_c_2839_n ) capacitor c=0.0200405f \
 //x=23.28 //y=1.665 //x2=22.71 //y2=0.995
cc_1388 ( N_noxref_10_M14_noxref_d N_noxref_20_M13_noxref_d ) capacitor \
 c=5.27807e-19 //x=23.005 //y=0.915 //x2=21.47 //y2=0.91
cc_1389 ( N_noxref_10_c_2170_n N_noxref_20_M14_noxref_s ) capacitor \
 c=0.00243521f //x=23.565 //y=3.33 //x2=22.575 //y2=0.375
cc_1390 ( N_noxref_10_c_2174_n N_noxref_20_M14_noxref_s ) capacitor \
 c=0.020752f //x=23.595 //y=1.665 //x2=22.575 //y2=0.375
cc_1391 ( N_noxref_10_M14_noxref_d N_noxref_20_M14_noxref_s ) capacitor \
 c=0.0426368f //x=23.005 //y=0.915 //x2=22.575 //y2=0.375
cc_1392 ( N_D_c_2345_n N_noxref_12_c_2416_n ) capacitor c=0.0034165f //x=0.915 \
 //y=1.915 //x2=0.695 //y2=1.495
cc_1393 ( N_D_c_2340_n N_noxref_12_c_2397_n ) capacitor c=0.0118986f //x=1.11 \
 //y=2.08 //x2=1.58 //y2=1.58
cc_1394 ( N_D_c_2344_n N_noxref_12_c_2397_n ) capacitor c=0.00703567f \
 //x=0.915 //y=1.52 //x2=1.58 //y2=1.58
cc_1395 ( N_D_c_2345_n N_noxref_12_c_2397_n ) capacitor c=0.0216532f //x=0.915 \
 //y=1.915 //x2=1.58 //y2=1.58
cc_1396 ( N_D_c_2347_n N_noxref_12_c_2397_n ) capacitor c=0.00780629f //x=1.29 \
 //y=1.365 //x2=1.58 //y2=1.58
cc_1397 ( N_D_c_2350_n N_noxref_12_c_2397_n ) capacitor c=0.00339872f \
 //x=1.445 //y=1.21 //x2=1.58 //y2=1.58
cc_1398 ( N_D_c_2345_n N_noxref_12_c_2404_n ) capacitor c=6.71402e-19 \
 //x=0.915 //y=1.915 //x2=1.665 //y2=1.495
cc_1399 ( N_D_c_2341_n N_noxref_12_M0_noxref_s ) capacitor c=0.0326577f \
 //x=0.915 //y=0.865 //x2=0.56 //y2=0.365
cc_1400 ( N_D_c_2344_n N_noxref_12_M0_noxref_s ) capacitor c=3.48408e-19 \
 //x=0.915 //y=1.52 //x2=0.56 //y2=0.365
cc_1401 ( N_D_c_2348_n N_noxref_12_M0_noxref_s ) capacitor c=0.0120759f \
 //x=1.445 //y=0.865 //x2=0.56 //y2=0.365
cc_1402 ( N_noxref_12_c_2408_n N_noxref_13_M2_noxref_s ) capacitor \
 c=0.00199452f //x=2.635 //y=0.615 //x2=3.785 //y2=0.375
cc_1403 ( N_noxref_13_c_2452_n N_noxref_14_c_2497_n ) capacitor c=0.0133059f \
 //x=5.775 //y=0.54 //x2=6.345 //y2=0.995
cc_1404 ( N_noxref_13_c_2472_n N_noxref_14_c_2497_n ) capacitor c=0.0100097f \
 //x=5.775 //y=1.59 //x2=6.345 //y2=0.995
cc_1405 ( N_noxref_13_M2_noxref_s N_noxref_14_c_2497_n ) capacitor \
 c=0.0224457f //x=3.785 //y=0.375 //x2=6.345 //y2=0.995
cc_1406 ( N_noxref_13_M2_noxref_s N_noxref_14_c_2499_n ) capacitor \
 c=0.0180035f //x=3.785 //y=0.375 //x2=6.43 //y2=0.625
cc_1407 ( N_noxref_13_c_2452_n N_noxref_14_M3_noxref_d ) capacitor \
 c=0.0128027f //x=5.775 //y=0.54 //x2=5.19 //y2=0.91
cc_1408 ( N_noxref_13_c_2472_n N_noxref_14_M3_noxref_d ) capacitor \
 c=0.00879751f //x=5.775 //y=1.59 //x2=5.19 //y2=0.91
cc_1409 ( N_noxref_13_M2_noxref_s N_noxref_14_M3_noxref_d ) capacitor \
 c=0.0159202f //x=3.785 //y=0.375 //x2=5.19 //y2=0.91
cc_1410 ( N_noxref_13_M2_noxref_s N_noxref_14_M4_noxref_s ) capacitor \
 c=0.0213553f //x=3.785 //y=0.375 //x2=6.295 //y2=0.375
cc_1411 ( N_noxref_14_c_2505_n N_noxref_15_M5_noxref_s ) capacitor \
 c=0.00191848f //x=7.4 //y=0.625 //x2=8.595 //y2=0.375
cc_1412 ( N_noxref_15_c_2557_n N_noxref_16_c_2604_n ) capacitor c=0.0131801f \
 //x=10.585 //y=0.54 //x2=11.155 //y2=0.995
cc_1413 ( N_noxref_15_c_2583_n N_noxref_16_c_2604_n ) capacitor c=0.00980353f \
 //x=10.585 //y=1.59 //x2=11.155 //y2=0.995
cc_1414 ( N_noxref_15_M5_noxref_s N_noxref_16_c_2604_n ) capacitor \
 c=0.0221661f //x=8.595 //y=0.375 //x2=11.155 //y2=0.995
cc_1415 ( N_noxref_15_M5_noxref_s N_noxref_16_c_2606_n ) capacitor \
 c=0.0180035f //x=8.595 //y=0.375 //x2=11.24 //y2=0.625
cc_1416 ( N_noxref_15_c_2557_n N_noxref_16_M6_noxref_d ) capacitor \
 c=0.0128434f //x=10.585 //y=0.54 //x2=10 //y2=0.91
cc_1417 ( N_noxref_15_c_2583_n N_noxref_16_M6_noxref_d ) capacitor \
 c=0.00886823f //x=10.585 //y=1.59 //x2=10 //y2=0.91
cc_1418 ( N_noxref_15_M5_noxref_s N_noxref_16_M6_noxref_d ) capacitor \
 c=0.0159202f //x=8.595 //y=0.375 //x2=10 //y2=0.91
cc_1419 ( N_noxref_15_M5_noxref_s N_noxref_16_M7_noxref_s ) capacitor \
 c=0.0213553f //x=8.595 //y=0.375 //x2=11.105 //y2=0.375
cc_1420 ( N_noxref_16_c_2612_n N_noxref_17_M8_noxref_s ) capacitor \
 c=0.00164795f //x=12.21 //y=0.625 //x2=13.51 //y2=0.365
cc_1421 ( N_noxref_17_c_2668_n N_noxref_18_M10_noxref_s ) capacitor \
 c=0.00174327f //x=15.585 //y=0.615 //x2=16.84 //y2=0.365
cc_1422 ( N_noxref_18_c_2720_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00199452f //x=18.915 //y=0.615 //x2=20.065 //y2=0.375
cc_1423 ( N_noxref_19_c_2768_n N_noxref_20_c_2811_n ) capacitor c=0.0132461f \
 //x=22.055 //y=0.54 //x2=22.625 //y2=0.995
cc_1424 ( N_noxref_19_c_2791_n N_noxref_20_c_2811_n ) capacitor c=0.00990219f \
 //x=22.055 //y=1.59 //x2=22.625 //y2=0.995
cc_1425 ( N_noxref_19_M12_noxref_s N_noxref_20_c_2811_n ) capacitor \
 c=0.0227445f //x=20.065 //y=0.375 //x2=22.625 //y2=0.995
cc_1426 ( N_noxref_19_M12_noxref_s N_noxref_20_c_2813_n ) capacitor \
 c=0.0180035f //x=20.065 //y=0.375 //x2=22.71 //y2=0.625
cc_1427 ( N_noxref_19_c_2768_n N_noxref_20_M13_noxref_d ) capacitor \
 c=0.0127176f //x=22.055 //y=0.54 //x2=21.47 //y2=0.91
cc_1428 ( N_noxref_19_c_2791_n N_noxref_20_M13_noxref_d ) capacitor \
 c=0.0086073f //x=22.055 //y=1.59 //x2=21.47 //y2=0.91
cc_1429 ( N_noxref_19_M12_noxref_s N_noxref_20_M13_noxref_d ) capacitor \
 c=0.0159202f //x=20.065 //y=0.375 //x2=21.47 //y2=0.91
cc_1430 ( N_noxref_19_M12_noxref_s N_noxref_20_M14_noxref_s ) capacitor \
 c=0.0213553f //x=20.065 //y=0.375 //x2=22.575 //y2=0.375
