// File: TMRDFFSNRNQNX1.spi.pex
// Created: Tue Oct 15 15:53:00 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_TMRDFFSNRNQNX1\%GND ( 1 163 167 170 175 185 193 203 211 221 229 239 \
 247 257 265 275 283 293 301 311 319 329 337 347 355 365 373 383 391 401 409 \
 419 427 437 445 455 463 473 481 491 499 507 513 519 532 536 538 540 542 544 \
 546 548 550 552 554 556 558 560 562 564 566 568 570 572 575 577 578 579 580 \
 581 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 )
c1062 ( 597 0 ) capacitor c=0.0215012f //x=94.23 //y=0.865
c1063 ( 596 0 ) capacitor c=0.0215012f //x=90.9 //y=0.865
c1064 ( 595 0 ) capacitor c=0.0207058f //x=87.57 //y=0.865
c1065 ( 594 0 ) capacitor c=0.0225929f //x=82.655 //y=0.875
c1066 ( 593 0 ) capacitor c=0.0225954f //x=77.845 //y=0.875
c1067 ( 592 0 ) capacitor c=0.0225954f //x=73.035 //y=0.875
c1068 ( 591 0 ) capacitor c=0.0225954f //x=68.225 //y=0.875
c1069 ( 590 0 ) capacitor c=0.0225954f //x=63.415 //y=0.875
c1070 ( 589 0 ) capacitor c=0.0225954f //x=58.605 //y=0.875
c1071 ( 588 0 ) capacitor c=0.0225954f //x=53.795 //y=0.875
c1072 ( 587 0 ) capacitor c=0.0225954f //x=48.985 //y=0.875
c1073 ( 586 0 ) capacitor c=0.0225954f //x=44.175 //y=0.875
c1074 ( 585 0 ) capacitor c=0.0225954f //x=39.365 //y=0.875
c1075 ( 584 0 ) capacitor c=0.0225954f //x=34.555 //y=0.875
c1076 ( 583 0 ) capacitor c=0.0225954f //x=29.745 //y=0.875
c1077 ( 582 0 ) capacitor c=0.0225954f //x=24.935 //y=0.875
c1078 ( 581 0 ) capacitor c=0.0225954f //x=20.125 //y=0.875
c1079 ( 580 0 ) capacitor c=0.0225954f //x=15.315 //y=0.875
c1080 ( 579 0 ) capacitor c=0.0225954f //x=10.505 //y=0.875
c1081 ( 578 0 ) capacitor c=0.0225954f //x=5.695 //y=0.875
c1082 ( 577 0 ) capacitor c=0.022675f //x=0.885 //y=0.875
c1083 ( 576 0 ) capacitor c=0.00440095f //x=94.42 //y=0
c1084 ( 575 0 ) capacitor c=0.101195f //x=93.24 //y=0
c1085 ( 574 0 ) capacitor c=0.00440095f //x=91.02 //y=0
c1086 ( 572 0 ) capacitor c=0.116097f //x=89.91 //y=0
c1087 ( 571 0 ) capacitor c=0.00440095f //x=87.76 //y=0
c1088 ( 570 0 ) capacitor c=0.106684f //x=86.58 //y=0
c1089 ( 569 0 ) capacitor c=0.00440144f //x=82.845 //y=0
c1090 ( 568 0 ) capacitor c=0.107013f //x=81.77 //y=0
c1091 ( 567 0 ) capacitor c=0.00440144f //x=78.035 //y=0
c1092 ( 566 0 ) capacitor c=0.106777f //x=76.96 //y=0
c1093 ( 565 0 ) capacitor c=0.00440144f //x=73.225 //y=0
c1094 ( 564 0 ) capacitor c=0.107052f //x=72.15 //y=0
c1095 ( 563 0 ) capacitor c=0.00440144f //x=68.415 //y=0
c1096 ( 562 0 ) capacitor c=0.107294f //x=67.34 //y=0
c1097 ( 561 0 ) capacitor c=0.00440144f //x=63.605 //y=0
c1098 ( 560 0 ) capacitor c=0.10703f //x=62.53 //y=0
c1099 ( 559 0 ) capacitor c=0.00440144f //x=58.795 //y=0
c1100 ( 558 0 ) capacitor c=0.106176f //x=57.72 //y=0
c1101 ( 557 0 ) capacitor c=0.00440144f //x=53.985 //y=0
c1102 ( 556 0 ) capacitor c=0.107346f //x=52.91 //y=0
c1103 ( 555 0 ) capacitor c=0.00440144f //x=49.175 //y=0
c1104 ( 554 0 ) capacitor c=0.106777f //x=48.1 //y=0
c1105 ( 553 0 ) capacitor c=0.00440144f //x=44.365 //y=0
c1106 ( 552 0 ) capacitor c=0.107052f //x=43.29 //y=0
c1107 ( 551 0 ) capacitor c=0.00440144f //x=39.555 //y=0
c1108 ( 550 0 ) capacitor c=0.107294f //x=38.48 //y=0
c1109 ( 549 0 ) capacitor c=0.00440144f //x=34.745 //y=0
c1110 ( 548 0 ) capacitor c=0.10703f //x=33.67 //y=0
c1111 ( 547 0 ) capacitor c=0.00440144f //x=29.935 //y=0
c1112 ( 546 0 ) capacitor c=0.107024f //x=28.86 //y=0
c1113 ( 545 0 ) capacitor c=0.00440144f //x=25.125 //y=0
c1114 ( 544 0 ) capacitor c=0.10703f //x=24.05 //y=0
c1115 ( 543 0 ) capacitor c=0.00440144f //x=20.315 //y=0
c1116 ( 542 0 ) capacitor c=0.106903f //x=19.24 //y=0
c1117 ( 541 0 ) capacitor c=0.00440144f //x=15.505 //y=0
c1118 ( 540 0 ) capacitor c=0.107052f //x=14.43 //y=0
c1119 ( 539 0 ) capacitor c=0.00440144f //x=10.695 //y=0
c1120 ( 538 0 ) capacitor c=0.107294f //x=9.62 //y=0
c1121 ( 537 0 ) capacitor c=0.00440144f //x=5.885 //y=0
c1122 ( 536 0 ) capacitor c=0.10703f //x=4.81 //y=0
c1123 ( 535 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c1124 ( 532 0 ) capacitor c=0.258637f //x=95.83 //y=0
c1125 ( 519 0 ) capacitor c=0.0389876f //x=94.335 //y=0
c1126 ( 513 0 ) capacitor c=0.0716428f //x=93.07 //y=0
c1127 ( 507 0 ) capacitor c=0.0388276f //x=91.005 //y=0
c1128 ( 499 0 ) capacitor c=0.0717274f //x=89.74 //y=0
c1129 ( 491 0 ) capacitor c=0.039094f //x=87.675 //y=0
c1130 ( 481 0 ) capacitor c=0.133362f //x=86.41 //y=0
c1131 ( 473 0 ) capacitor c=0.0339325f //x=82.76 //y=0
c1132 ( 463 0 ) capacitor c=0.133705f //x=81.6 //y=0
c1133 ( 455 0 ) capacitor c=0.0339325f //x=77.95 //y=0
c1134 ( 445 0 ) capacitor c=0.133561f //x=76.79 //y=0
c1135 ( 437 0 ) capacitor c=0.0339325f //x=73.14 //y=0
c1136 ( 427 0 ) capacitor c=0.133362f //x=71.98 //y=0
c1137 ( 419 0 ) capacitor c=0.0339325f //x=68.33 //y=0
c1138 ( 409 0 ) capacitor c=0.133362f //x=67.17 //y=0
c1139 ( 401 0 ) capacitor c=0.0339325f //x=63.52 //y=0
c1140 ( 391 0 ) capacitor c=0.133362f //x=62.36 //y=0
c1141 ( 383 0 ) capacitor c=0.0339325f //x=58.71 //y=0
c1142 ( 373 0 ) capacitor c=0.133362f //x=57.55 //y=0
c1143 ( 365 0 ) capacitor c=0.0339325f //x=53.9 //y=0
c1144 ( 355 0 ) capacitor c=0.133362f //x=52.74 //y=0
c1145 ( 347 0 ) capacitor c=0.0339325f //x=49.09 //y=0
c1146 ( 337 0 ) capacitor c=0.133561f //x=47.93 //y=0
c1147 ( 329 0 ) capacitor c=0.0339325f //x=44.28 //y=0
c1148 ( 319 0 ) capacitor c=0.133362f //x=43.12 //y=0
c1149 ( 311 0 ) capacitor c=0.0339325f //x=39.47 //y=0
c1150 ( 301 0 ) capacitor c=0.133362f //x=38.31 //y=0
c1151 ( 293 0 ) capacitor c=0.0339325f //x=34.66 //y=0
c1152 ( 283 0 ) capacitor c=0.133362f //x=33.5 //y=0
c1153 ( 275 0 ) capacitor c=0.0339325f //x=29.85 //y=0
c1154 ( 265 0 ) capacitor c=0.133362f //x=28.69 //y=0
c1155 ( 257 0 ) capacitor c=0.0339325f //x=25.04 //y=0
c1156 ( 247 0 ) capacitor c=0.133362f //x=23.88 //y=0
c1157 ( 239 0 ) capacitor c=0.0339325f //x=20.23 //y=0
c1158 ( 229 0 ) capacitor c=0.133561f //x=19.07 //y=0
c1159 ( 221 0 ) capacitor c=0.0339325f //x=15.42 //y=0
c1160 ( 211 0 ) capacitor c=0.133362f //x=14.26 //y=0
c1161 ( 203 0 ) capacitor c=0.0339325f //x=10.61 //y=0
c1162 ( 193 0 ) capacitor c=0.133362f //x=9.45 //y=0
c1163 ( 185 0 ) capacitor c=0.0339325f //x=5.8 //y=0
c1164 ( 175 0 ) capacitor c=0.133402f //x=4.64 //y=0
c1165 ( 170 0 ) capacitor c=0.178058f //x=0.74 //y=0
c1166 ( 167 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c1167 ( 163 0 ) capacitor c=2.86297f //x=95.83 //y=0
r1168 (  530 532 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=94.72 //y=0 //x2=95.83 //y2=0
r1169 (  528 576 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.505 //y=0 //x2=94.42 //y2=0
r1170 (  528 530 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=94.505 //y=0 //x2=94.72 //y2=0
r1171 (  523 576 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=94.42 //y=0.17 //x2=94.42 //y2=0
r1172 (  523 597 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=94.42 //y=0.17 //x2=94.42 //y2=0.955
r1173 (  520 575 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=93.41 //y=0 //x2=93.24 //y2=0
r1174 (  520 522 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=93.41 //y=0 //x2=93.61 //y2=0
r1175 (  519 576 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.335 //y=0 //x2=94.42 //y2=0
r1176 (  519 522 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=94.335 //y=0 //x2=93.61 //y2=0
r1177 (  514 574 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.175 //y=0 //x2=91.09 //y2=0
r1178 (  514 516 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=91.175 //y=0 //x2=92.13 //y2=0
r1179 (  513 575 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=93.07 //y=0 //x2=93.24 //y2=0
r1180 (  513 516 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=93.07 //y=0 //x2=92.13 //y2=0
r1181 (  509 574 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=91.09 //y=0.17 //x2=91.09 //y2=0
r1182 (  509 596 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=91.09 //y=0.17 //x2=91.09 //y2=0.955
r1183 (  508 572 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=90.08 //y=0 //x2=89.91 //y2=0
r1184 (  507 574 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.005 //y=0 //x2=91.09 //y2=0
r1185 (  507 508 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=91.005 //y=0 //x2=90.08 //y2=0
r1186 (  502 504 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=88.43 //y=0 //x2=89.54 //y2=0
r1187 (  500 571 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=87.845 //y=0 //x2=87.76 //y2=0
r1188 (  500 502 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=87.845 //y=0 //x2=88.43 //y2=0
r1189 (  499 572 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=89.74 //y=0 //x2=89.91 //y2=0
r1190 (  499 504 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=89.74 //y=0 //x2=89.54 //y2=0
r1191 (  495 571 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=87.76 //y=0.17 //x2=87.76 //y2=0
r1192 (  495 595 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=87.76 //y=0.17 //x2=87.76 //y2=0.955
r1193 (  492 570 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=86.75 //y=0 //x2=86.58 //y2=0
r1194 (  492 494 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=86.75 //y=0 //x2=87.32 //y2=0
r1195 (  491 571 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=87.675 //y=0 //x2=87.76 //y2=0
r1196 (  491 494 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=87.675 //y=0 //x2=87.32 //y2=0
r1197 (  486 488 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=84.73 //y=0 //x2=85.84 //y2=0
r1198 (  484 486 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=83.62 //y=0 //x2=84.73 //y2=0
r1199 (  482 569 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.93 //y=0 //x2=82.845 //y2=0
r1200 (  482 484 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=82.93 //y=0 //x2=83.62 //y2=0
r1201 (  481 570 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=86.41 //y=0 //x2=86.58 //y2=0
r1202 (  481 488 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=86.41 //y=0 //x2=85.84 //y2=0
r1203 (  477 569 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=82.845 //y=0.17 //x2=82.845 //y2=0
r1204 (  477 594 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=82.845 //y=0.17 //x2=82.845 //y2=0.965
r1205 (  474 568 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.94 //y=0 //x2=81.77 //y2=0
r1206 (  474 476 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=81.94 //y=0 //x2=82.51 //y2=0
r1207 (  473 569 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.76 //y=0 //x2=82.845 //y2=0
r1208 (  473 476 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=82.76 //y=0 //x2=82.51 //y2=0
r1209 (  468 470 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=79.92 //y=0 //x2=81.03 //y2=0
r1210 (  466 468 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=78.81 //y=0 //x2=79.92 //y2=0
r1211 (  464 567 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.12 //y=0 //x2=78.035 //y2=0
r1212 (  464 466 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=78.12 //y=0 //x2=78.81 //y2=0
r1213 (  463 568 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.6 //y=0 //x2=81.77 //y2=0
r1214 (  463 470 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=81.6 //y=0 //x2=81.03 //y2=0
r1215 (  459 567 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=78.035 //y=0.17 //x2=78.035 //y2=0
r1216 (  459 593 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=78.035 //y=0.17 //x2=78.035 //y2=0.965
r1217 (  456 566 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.13 //y=0 //x2=76.96 //y2=0
r1218 (  456 458 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=77.13 //y=0 //x2=77.7 //y2=0
r1219 (  455 567 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.95 //y=0 //x2=78.035 //y2=0
r1220 (  455 458 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=77.95 //y=0 //x2=77.7 //y2=0
r1221 (  450 452 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=75.11 //y=0 //x2=76.22 //y2=0
r1222 (  448 450 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=74 //y=0 //x2=75.11 //y2=0
r1223 (  446 565 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.31 //y=0 //x2=73.225 //y2=0
r1224 (  446 448 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=73.31 //y=0 //x2=74 //y2=0
r1225 (  445 566 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.79 //y=0 //x2=76.96 //y2=0
r1226 (  445 452 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=76.79 //y=0 //x2=76.22 //y2=0
r1227 (  441 565 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.225 //y=0.17 //x2=73.225 //y2=0
r1228 (  441 592 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=73.225 //y=0.17 //x2=73.225 //y2=0.965
r1229 (  438 564 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=72.32 //y=0 //x2=72.15 //y2=0
r1230 (  438 440 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=72.32 //y=0 //x2=72.89 //y2=0
r1231 (  437 565 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.14 //y=0 //x2=73.225 //y2=0
r1232 (  437 440 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=73.14 //y=0 //x2=72.89 //y2=0
r1233 (  432 434 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=70.3 //y=0 //x2=71.41 //y2=0
r1234 (  430 432 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=69.19 //y=0 //x2=70.3 //y2=0
r1235 (  428 563 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.5 //y=0 //x2=68.415 //y2=0
r1236 (  428 430 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=68.5 //y=0 //x2=69.19 //y2=0
r1237 (  427 564 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.98 //y=0 //x2=72.15 //y2=0
r1238 (  427 434 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=71.98 //y=0 //x2=71.41 //y2=0
r1239 (  423 563 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.415 //y=0.17 //x2=68.415 //y2=0
r1240 (  423 591 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=68.415 //y=0.17 //x2=68.415 //y2=0.965
r1241 (  420 562 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.51 //y=0 //x2=67.34 //y2=0
r1242 (  420 422 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.51 //y=0 //x2=68.08 //y2=0
r1243 (  419 563 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.33 //y=0 //x2=68.415 //y2=0
r1244 (  419 422 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=68.33 //y=0 //x2=68.08 //y2=0
r1245 (  414 416 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=65.49 //y=0 //x2=66.6 //y2=0
r1246 (  412 414 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=64.38 //y=0 //x2=65.49 //y2=0
r1247 (  410 561 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.69 //y=0 //x2=63.605 //y2=0
r1248 (  410 412 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=63.69 //y=0 //x2=64.38 //y2=0
r1249 (  409 562 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.17 //y=0 //x2=67.34 //y2=0
r1250 (  409 416 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.17 //y=0 //x2=66.6 //y2=0
r1251 (  405 561 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=63.605 //y=0.17 //x2=63.605 //y2=0
r1252 (  405 590 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=63.605 //y=0.17 //x2=63.605 //y2=0.965
r1253 (  402 560 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.7 //y=0 //x2=62.53 //y2=0
r1254 (  402 404 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=62.7 //y=0 //x2=63.27 //y2=0
r1255 (  401 561 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.52 //y=0 //x2=63.605 //y2=0
r1256 (  401 404 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=63.52 //y=0 //x2=63.27 //y2=0
r1257 (  396 398 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=60.68 //y=0 //x2=61.79 //y2=0
r1258 (  394 396 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=59.57 //y=0 //x2=60.68 //y2=0
r1259 (  392 559 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.88 //y=0 //x2=58.795 //y2=0
r1260 (  392 394 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=58.88 //y=0 //x2=59.57 //y2=0
r1261 (  391 560 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.36 //y=0 //x2=62.53 //y2=0
r1262 (  391 398 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=62.36 //y=0 //x2=61.79 //y2=0
r1263 (  387 559 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.795 //y=0.17 //x2=58.795 //y2=0
r1264 (  387 589 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=58.795 //y=0.17 //x2=58.795 //y2=0.965
r1265 (  384 558 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.89 //y=0 //x2=57.72 //y2=0
r1266 (  384 386 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=57.89 //y=0 //x2=58.46 //y2=0
r1267 (  383 559 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.71 //y=0 //x2=58.795 //y2=0
r1268 (  383 386 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=58.71 //y=0 //x2=58.46 //y2=0
r1269 (  378 380 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=55.87 //y=0 //x2=56.98 //y2=0
r1270 (  376 378 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=54.76 //y=0 //x2=55.87 //y2=0
r1271 (  374 557 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.07 //y=0 //x2=53.985 //y2=0
r1272 (  374 376 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=54.07 //y=0 //x2=54.76 //y2=0
r1273 (  373 558 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.55 //y=0 //x2=57.72 //y2=0
r1274 (  373 380 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=57.55 //y=0 //x2=56.98 //y2=0
r1275 (  369 557 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.985 //y=0.17 //x2=53.985 //y2=0
r1276 (  369 588 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=53.985 //y=0.17 //x2=53.985 //y2=0.965
r1277 (  366 556 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.08 //y=0 //x2=52.91 //y2=0
r1278 (  366 368 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=53.08 //y=0 //x2=53.65 //y2=0
r1279 (  365 557 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.9 //y=0 //x2=53.985 //y2=0
r1280 (  365 368 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=53.9 //y=0 //x2=53.65 //y2=0
r1281 (  360 362 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=51.06 //y=0 //x2=52.17 //y2=0
r1282 (  358 360 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=49.95 //y=0 //x2=51.06 //y2=0
r1283 (  356 555 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.26 //y=0 //x2=49.175 //y2=0
r1284 (  356 358 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=49.26 //y=0 //x2=49.95 //y2=0
r1285 (  355 556 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.74 //y=0 //x2=52.91 //y2=0
r1286 (  355 362 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=52.74 //y=0 //x2=52.17 //y2=0
r1287 (  351 555 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.175 //y=0.17 //x2=49.175 //y2=0
r1288 (  351 587 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=49.175 //y=0.17 //x2=49.175 //y2=0.965
r1289 (  348 554 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.27 //y=0 //x2=48.1 //y2=0
r1290 (  348 350 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.27 //y=0 //x2=48.84 //y2=0
r1291 (  347 555 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.09 //y=0 //x2=49.175 //y2=0
r1292 (  347 350 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=49.09 //y=0 //x2=48.84 //y2=0
r1293 (  342 344 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=46.25 //y=0 //x2=47.36 //y2=0
r1294 (  340 342 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=45.14 //y=0 //x2=46.25 //y2=0
r1295 (  338 553 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.45 //y=0 //x2=44.365 //y2=0
r1296 (  338 340 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=44.45 //y=0 //x2=45.14 //y2=0
r1297 (  337 554 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.93 //y=0 //x2=48.1 //y2=0
r1298 (  337 344 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=47.93 //y=0 //x2=47.36 //y2=0
r1299 (  333 553 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.365 //y=0.17 //x2=44.365 //y2=0
r1300 (  333 586 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=44.365 //y=0.17 //x2=44.365 //y2=0.965
r1301 (  330 552 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.46 //y=0 //x2=43.29 //y2=0
r1302 (  330 332 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.46 //y=0 //x2=44.03 //y2=0
r1303 (  329 553 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.28 //y=0 //x2=44.365 //y2=0
r1304 (  329 332 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=44.28 //y=0 //x2=44.03 //y2=0
r1305 (  324 326 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=41.44 //y=0 //x2=42.55 //y2=0
r1306 (  322 324 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=40.33 //y=0 //x2=41.44 //y2=0
r1307 (  320 551 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.64 //y=0 //x2=39.555 //y2=0
r1308 (  320 322 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=39.64 //y=0 //x2=40.33 //y2=0
r1309 (  319 552 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.12 //y=0 //x2=43.29 //y2=0
r1310 (  319 326 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.12 //y=0 //x2=42.55 //y2=0
r1311 (  315 551 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.555 //y=0.17 //x2=39.555 //y2=0
r1312 (  315 585 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=39.555 //y=0.17 //x2=39.555 //y2=0.965
r1313 (  312 550 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.65 //y=0 //x2=38.48 //y2=0
r1314 (  312 314 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.65 //y=0 //x2=39.22 //y2=0
r1315 (  311 551 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.47 //y=0 //x2=39.555 //y2=0
r1316 (  311 314 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=39.47 //y=0 //x2=39.22 //y2=0
r1317 (  306 308 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=36.63 //y=0 //x2=37.74 //y2=0
r1318 (  304 306 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=35.52 //y=0 //x2=36.63 //y2=0
r1319 (  302 549 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.83 //y=0 //x2=34.745 //y2=0
r1320 (  302 304 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=34.83 //y=0 //x2=35.52 //y2=0
r1321 (  301 550 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.31 //y=0 //x2=38.48 //y2=0
r1322 (  301 308 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.31 //y=0 //x2=37.74 //y2=0
r1323 (  297 549 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.745 //y=0.17 //x2=34.745 //y2=0
r1324 (  297 584 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=34.745 //y=0.17 //x2=34.745 //y2=0.965
r1325 (  294 548 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.84 //y=0 //x2=33.67 //y2=0
r1326 (  294 296 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=33.84 //y=0 //x2=34.41 //y2=0
r1327 (  293 549 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.66 //y=0 //x2=34.745 //y2=0
r1328 (  293 296 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=34.66 //y=0 //x2=34.41 //y2=0
r1329 (  288 290 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=31.82 //y=0 //x2=32.93 //y2=0
r1330 (  286 288 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=30.71 //y=0 //x2=31.82 //y2=0
r1331 (  284 547 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.02 //y=0 //x2=29.935 //y2=0
r1332 (  284 286 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=30.02 //y=0 //x2=30.71 //y2=0
r1333 (  283 548 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.5 //y=0 //x2=33.67 //y2=0
r1334 (  283 290 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=33.5 //y=0 //x2=32.93 //y2=0
r1335 (  279 547 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.935 //y=0.17 //x2=29.935 //y2=0
r1336 (  279 583 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=29.935 //y=0.17 //x2=29.935 //y2=0.965
r1337 (  276 546 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.03 //y=0 //x2=28.86 //y2=0
r1338 (  276 278 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=29.03 //y=0 //x2=29.6 //y2=0
r1339 (  275 547 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.85 //y=0 //x2=29.935 //y2=0
r1340 (  275 278 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=29.85 //y=0 //x2=29.6 //y2=0
r1341 (  270 272 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=27.01 //y=0 //x2=28.12 //y2=0
r1342 (  268 270 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=25.9 //y=0 //x2=27.01 //y2=0
r1343 (  266 545 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.21 //y=0 //x2=25.125 //y2=0
r1344 (  266 268 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=25.21 //y=0 //x2=25.9 //y2=0
r1345 (  265 546 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.69 //y=0 //x2=28.86 //y2=0
r1346 (  265 272 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=28.69 //y=0 //x2=28.12 //y2=0
r1347 (  261 545 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.125 //y=0.17 //x2=25.125 //y2=0
r1348 (  261 582 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=25.125 //y=0.17 //x2=25.125 //y2=0.965
r1349 (  258 544 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.22 //y=0 //x2=24.05 //y2=0
r1350 (  258 260 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.22 //y=0 //x2=24.79 //y2=0
r1351 (  257 545 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.04 //y=0 //x2=25.125 //y2=0
r1352 (  257 260 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=25.04 //y=0 //x2=24.79 //y2=0
r1353 (  252 254 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=22.2 //y=0 //x2=23.31 //y2=0
r1354 (  250 252 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.09 //y=0 //x2=22.2 //y2=0
r1355 (  248 543 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.4 //y=0 //x2=20.315 //y2=0
r1356 (  248 250 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=20.4 //y=0 //x2=21.09 //y2=0
r1357 (  247 544 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.88 //y=0 //x2=24.05 //y2=0
r1358 (  247 254 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.88 //y=0 //x2=23.31 //y2=0
r1359 (  243 543 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.315 //y=0.17 //x2=20.315 //y2=0
r1360 (  243 581 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=20.315 //y=0.17 //x2=20.315 //y2=0.965
r1361 (  240 542 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.41 //y=0 //x2=19.24 //y2=0
r1362 (  240 242 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.41 //y=0 //x2=19.98 //y2=0
r1363 (  239 543 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.23 //y=0 //x2=20.315 //y2=0
r1364 (  239 242 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=20.23 //y=0 //x2=19.98 //y2=0
r1365 (  234 236 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.39 //y=0 //x2=18.5 //y2=0
r1366 (  232 234 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=16.28 //y=0 //x2=17.39 //y2=0
r1367 (  230 541 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.59 //y=0 //x2=15.505 //y2=0
r1368 (  230 232 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=15.59 //y=0 //x2=16.28 //y2=0
r1369 (  229 542 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.07 //y=0 //x2=19.24 //y2=0
r1370 (  229 236 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.07 //y=0 //x2=18.5 //y2=0
r1371 (  225 541 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.505 //y=0.17 //x2=15.505 //y2=0
r1372 (  225 580 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=15.505 //y=0.17 //x2=15.505 //y2=0.965
r1373 (  222 540 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=14.43 //y2=0
r1374 (  222 224 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=15.17 //y2=0
r1375 (  221 541 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.42 //y=0 //x2=15.505 //y2=0
r1376 (  221 224 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=15.42 //y=0 //x2=15.17 //y2=0
r1377 (  216 218 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=12.58 //y=0 //x2=13.69 //y2=0
r1378 (  214 216 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r1379 (  212 539 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.78 //y=0 //x2=10.695 //y2=0
r1380 (  212 214 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=10.78 //y=0 //x2=11.47 //y2=0
r1381 (  211 540 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=14.43 //y2=0
r1382 (  211 218 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=13.69 //y2=0
r1383 (  207 539 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.695 //y=0.17 //x2=10.695 //y2=0
r1384 (  207 579 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=10.695 //y=0.17 //x2=10.695 //y2=0.965
r1385 (  204 538 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=9.62 //y2=0
r1386 (  204 206 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=10.36 //y2=0
r1387 (  203 539 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.61 //y=0 //x2=10.695 //y2=0
r1388 (  203 206 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=10.61 //y=0 //x2=10.36 //y2=0
r1389 (  198 200 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.77 //y=0 //x2=8.88 //y2=0
r1390 (  196 198 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r1391 (  194 537 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=5.885 //y2=0
r1392 (  194 196 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=6.66 //y2=0
r1393 (  193 538 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=9.62 //y2=0
r1394 (  193 200 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=8.88 //y2=0
r1395 (  189 537 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0
r1396 (  189 578 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0.965
r1397 (  186 536 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=4.81 //y2=0
r1398 (  186 188 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=5.55 //y2=0
r1399 (  185 537 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.885 //y2=0
r1400 (  185 188 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.55 //y2=0
r1401 (  180 182 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r1402 (  178 180 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r1403 (  176 535 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r1404 (  176 178 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r1405 (  175 536 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.81 //y2=0
r1406 (  175 182 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r1407 (  171 535 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r1408 (  171 577 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r1409 (  167 535 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r1410 (  167 170 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r1411 (  163 532 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=95.83 //y=0 //x2=95.83 //y2=0
r1412 (  161 530 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=94.72 //y=0 //x2=94.72 //y2=0
r1413 (  161 163 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=94.72 //y=0 //x2=95.83 //y2=0
r1414 (  159 522 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=93.61 //y=0 //x2=93.61 //y2=0
r1415 (  159 161 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=93.61 //y=0 //x2=94.72 //y2=0
r1416 (  157 516 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=92.13 //y=0 //x2=92.13 //y2=0
r1417 (  157 159 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=92.13 //y=0 //x2=93.61 //y2=0
r1418 (  155 574 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=91.02 //y=0 //x2=91.02 //y2=0
r1419 (  155 157 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=91.02 //y=0 //x2=92.13 //y2=0
r1420 (  153 504 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=89.54 //y=0 //x2=89.54 //y2=0
r1421 (  153 155 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=89.54 //y=0 //x2=91.02 //y2=0
r1422 (  151 502 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=88.43 //y=0 //x2=88.43 //y2=0
r1423 (  151 153 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=88.43 //y=0 //x2=89.54 //y2=0
r1424 (  149 494 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=87.32 //y=0 //x2=87.32 //y2=0
r1425 (  149 151 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=87.32 //y=0 //x2=88.43 //y2=0
r1426 (  147 488 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=85.84 //y=0 //x2=85.84 //y2=0
r1427 (  147 149 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=85.84 //y=0 //x2=87.32 //y2=0
r1428 (  145 486 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=84.73 //y=0 //x2=84.73 //y2=0
r1429 (  145 147 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=84.73 //y=0 //x2=85.84 //y2=0
r1430 (  143 484 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=83.62 //y=0 //x2=83.62 //y2=0
r1431 (  143 145 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=83.62 //y=0 //x2=84.73 //y2=0
r1432 (  141 476 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.51 //y=0 //x2=82.51 //y2=0
r1433 (  141 143 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=82.51 //y=0 //x2=83.62 //y2=0
r1434 (  139 470 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=81.03 //y=0 //x2=81.03 //y2=0
r1435 (  139 141 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=81.03 //y=0 //x2=82.51 //y2=0
r1436 (  137 468 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=79.92 //y=0 //x2=79.92 //y2=0
r1437 (  137 139 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=79.92 //y=0 //x2=81.03 //y2=0
r1438 (  135 466 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.81 //y=0 //x2=78.81 //y2=0
r1439 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=78.81 //y=0 //x2=79.92 //y2=0
r1440 (  133 458 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=77.7 //y=0 //x2=77.7 //y2=0
r1441 (  133 135 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=77.7 //y=0 //x2=78.81 //y2=0
r1442 (  131 452 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.22 //y=0 //x2=76.22 //y2=0
r1443 (  131 133 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.22 //y=0 //x2=77.7 //y2=0
r1444 (  129 450 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.11 //y=0 //x2=75.11 //y2=0
r1445 (  129 131 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=0 //x2=76.22 //y2=0
r1446 (  127 448 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74 //y=0 //x2=74 //y2=0
r1447 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74 //y=0 //x2=75.11 //y2=0
r1448 (  125 440 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.89 //y=0 //x2=72.89 //y2=0
r1449 (  125 127 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=72.89 //y=0 //x2=74 //y2=0
r1450 (  123 434 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=0 //x2=71.41 //y2=0
r1451 (  123 125 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=0 //x2=72.89 //y2=0
r1452 (  121 432 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=70.3 //y=0 //x2=70.3 //y2=0
r1453 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=70.3 //y=0 //x2=71.41 //y2=0
r1454 (  119 430 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.19 //y=0 //x2=69.19 //y2=0
r1455 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.19 //y=0 //x2=70.3 //y2=0
r1456 (  117 422 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=68.08 //y=0 //x2=68.08 //y2=0
r1457 (  117 119 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=68.08 //y=0 //x2=69.19 //y2=0
r1458 (  115 416 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.6 //y=0 //x2=66.6 //y2=0
r1459 (  115 117 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=66.6 //y=0 //x2=68.08 //y2=0
r1460 (  113 414 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.49 //y=0 //x2=65.49 //y2=0
r1461 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.49 //y=0 //x2=66.6 //y2=0
r1462 (  111 412 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=64.38 //y=0 //x2=64.38 //y2=0
r1463 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=64.38 //y=0 //x2=65.49 //y2=0
r1464 (  109 404 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=63.27 //y=0 //x2=63.27 //y2=0
r1465 (  109 111 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=63.27 //y=0 //x2=64.38 //y2=0
r1466 (  107 398 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.79 //y=0 //x2=61.79 //y2=0
r1467 (  107 109 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.79 //y=0 //x2=63.27 //y2=0
r1468 (  105 396 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=60.68 //y=0 //x2=60.68 //y2=0
r1469 (  105 107 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=60.68 //y=0 //x2=61.79 //y2=0
r1470 (  103 394 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.57 //y=0 //x2=59.57 //y2=0
r1471 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.57 //y=0 //x2=60.68 //y2=0
r1472 (  101 386 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.46 //y=0 //x2=58.46 //y2=0
r1473 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.46 //y=0 //x2=59.57 //y2=0
r1474 (  99 380 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.98 //y=0 //x2=56.98 //y2=0
r1475 (  99 101 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.98 //y=0 //x2=58.46 //y2=0
r1476 (  97 378 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.87 //y=0 //x2=55.87 //y2=0
r1477 (  97 99 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.87 //y=0 //x2=56.98 //y2=0
r1478 (  95 376 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.76 //y=0 //x2=54.76 //y2=0
r1479 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.76 //y=0 //x2=55.87 //y2=0
r1480 (  93 368 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.65 //y=0 //x2=53.65 //y2=0
r1481 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=53.65 //y=0 //x2=54.76 //y2=0
r1482 (  91 362 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=52.17 //y=0 //x2=52.17 //y2=0
r1483 (  91 93 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=52.17 //y=0 //x2=53.65 //y2=0
r1484 (  89 360 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.06 //y=0 //x2=51.06 //y2=0
r1485 (  89 91 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=51.06 //y=0 //x2=52.17 //y2=0
r1486 (  87 358 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.95 //y=0 //x2=49.95 //y2=0
r1487 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.95 //y=0 //x2=51.06 //y2=0
r1488 (  85 350 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.84 //y=0 //x2=48.84 //y2=0
r1489 (  85 87 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=48.84 //y=0 //x2=49.95 //y2=0
r1490 (  82 344 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=47.36 //y=0 //x2=47.36 //y2=0
r1491 (  80 342 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.25 //y=0 //x2=46.25 //y2=0
r1492 (  80 82 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.25 //y=0 //x2=47.36 //y2=0
r1493 (  78 340 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.14 //y=0 //x2=45.14 //y2=0
r1494 (  78 80 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.14 //y=0 //x2=46.25 //y2=0
r1495 (  76 332 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.03 //y=0 //x2=44.03 //y2=0
r1496 (  76 78 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.03 //y=0 //x2=45.14 //y2=0
r1497 (  74 326 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.55 //y=0 //x2=42.55 //y2=0
r1498 (  74 76 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=42.55 //y=0 //x2=44.03 //y2=0
r1499 (  72 324 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.44 //y=0 //x2=41.44 //y2=0
r1500 (  72 74 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.44 //y=0 //x2=42.55 //y2=0
r1501 (  70 322 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=40.33 //y=0 //x2=40.33 //y2=0
r1502 (  70 72 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=40.33 //y=0 //x2=41.44 //y2=0
r1503 (  68 314 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.22 //y=0 //x2=39.22 //y2=0
r1504 (  68 70 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=39.22 //y=0 //x2=40.33 //y2=0
r1505 (  66 308 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37.74 //y=0 //x2=37.74 //y2=0
r1506 (  66 68 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=37.74 //y=0 //x2=39.22 //y2=0
r1507 (  64 306 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=36.63 //y=0 //x2=36.63 //y2=0
r1508 (  64 66 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=36.63 //y=0 //x2=37.74 //y2=0
r1509 (  62 304 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.52 //y=0 //x2=35.52 //y2=0
r1510 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.52 //y=0 //x2=36.63 //y2=0
r1511 (  60 296 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.41 //y=0 //x2=34.41 //y2=0
r1512 (  60 62 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.41 //y=0 //x2=35.52 //y2=0
r1513 (  58 290 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.93 //y=0 //x2=32.93 //y2=0
r1514 (  58 60 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.93 //y=0 //x2=34.41 //y2=0
r1515 (  56 288 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.82 //y=0 //x2=31.82 //y2=0
r1516 (  56 58 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.82 //y=0 //x2=32.93 //y2=0
r1517 (  54 286 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=30.71 //y=0 //x2=30.71 //y2=0
r1518 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=30.71 //y=0 //x2=31.82 //y2=0
r1519 (  52 278 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.6 //y=0 //x2=29.6 //y2=0
r1520 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=29.6 //y=0 //x2=30.71 //y2=0
r1521 (  50 272 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.12 //y=0 //x2=28.12 //y2=0
r1522 (  50 52 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=28.12 //y=0 //x2=29.6 //y2=0
r1523 (  48 270 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.01 //y=0 //x2=27.01 //y2=0
r1524 (  48 50 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.01 //y=0 //x2=28.12 //y2=0
r1525 (  46 268 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.9 //y=0 //x2=25.9 //y2=0
r1526 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.9 //y=0 //x2=27.01 //y2=0
r1527 (  44 260 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=0 //x2=24.79 //y2=0
r1528 (  44 46 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=0 //x2=25.9 //y2=0
r1529 (  42 254 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.31 //y=0 //x2=23.31 //y2=0
r1530 (  42 44 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.31 //y=0 //x2=24.79 //y2=0
r1531 (  40 252 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=0 //x2=22.2 //y2=0
r1532 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=0 //x2=23.31 //y2=0
r1533 (  38 250 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r1534 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=0 //x2=22.2 //y2=0
r1535 (  36 242 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=0 //x2=19.98 //y2=0
r1536 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=0 //x2=21.09 //y2=0
r1537 (  34 236 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=0 //x2=18.5 //y2=0
r1538 (  34 36 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=0 //x2=19.98 //y2=0
r1539 (  32 234 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=0 //x2=17.39 //y2=0
r1540 (  32 34 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=0 //x2=18.5 //y2=0
r1541 (  30 232 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=0 //x2=16.28 //y2=0
r1542 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=0 //x2=17.39 //y2=0
r1543 (  28 224 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r1544 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.28 //y2=0
r1545 (  26 218 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=0 //x2=13.69 //y2=0
r1546 (  26 28 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=0 //x2=15.17 //y2=0
r1547 (  24 216 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r1548 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=0 //x2=13.69 //y2=0
r1549 (  22 214 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r1550 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=0 //x2=12.58 //y2=0
r1551 (  20 206 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r1552 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r1553 (  18 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=0 //x2=8.88 //y2=0
r1554 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=0 //x2=10.36 //y2=0
r1555 (  16 198 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r1556 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=8.88 //y2=0
r1557 (  14 196 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r1558 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r1559 (  12 188 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r1560 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r1561 (  10 182 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r1562 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r1563 (  8 180 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r1564 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r1565 (  6 178 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r1566 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r1567 (  3 170 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r1568 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r1569 (  1 85 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=48.285 //y=0 //x2=48.84 //y2=0
r1570 (  1 82 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=48.285 //y=0 //x2=47.36 //y2=0
ends PM_TMRDFFSNRNQNX1\%GND

subckt PM_TMRDFFSNRNQNX1\%VDD ( 1 163 167 170 177 187 195 205 211 221 231 239 \
 249 255 265 275 283 293 299 309 319 327 337 343 353 363 371 381 387 397 407 \
 415 425 431 441 451 459 469 475 485 495 503 513 519 529 539 547 557 563 573 \
 583 591 601 607 617 627 635 645 651 661 671 679 689 695 705 715 723 733 739 \
 749 759 767 777 783 793 803 811 821 827 837 847 855 865 871 881 891 899 909 \
 915 925 935 943 953 959 967 975 985 991 1006 1013 1018 1023 1028 1033 1038 \
 1043 1048 1053 1058 1063 1068 1073 1078 1083 1088 1093 1098 1103 1104 1105 \
 1106 1107 1108 1109 1110 1111 1112 1113 1114 1115 1116 1117 1118 1119 1120 \
 1121 1122 1123 1124 1125 1126 1127 1128 1129 1130 1131 1132 1133 1134 1135 \
 1136 1137 1138 1139 1140 1141 1142 1143 1144 1145 1146 1147 1148 1149 1150 \
 1151 1152 1153 1154 1155 1156 1157 1158 1159 1160 1161 1162 1163 1164 1165 \
 1166 1167 1168 1169 1170 1171 1172 1173 1174 1175 1176 1177 1178 1179 )
c1158 ( 1179 0 ) capacitor c=0.0476806f //x=88.985 //y=5.025
c1159 ( 1178 0 ) capacitor c=0.0241714f //x=88.105 //y=5.025
c1160 ( 1177 0 ) capacitor c=0.0467094f //x=87.235 //y=5.025
c1161 ( 1176 0 ) capacitor c=0.0452179f //x=85.355 //y=5.02
c1162 ( 1175 0 ) capacitor c=0.024152f //x=84.475 //y=5.02
c1163 ( 1174 0 ) capacitor c=0.024152f //x=83.595 //y=5.02
c1164 ( 1173 0 ) capacitor c=0.053132f //x=82.725 //y=5.02
c1165 ( 1172 0 ) capacitor c=0.0452179f //x=80.545 //y=5.02
c1166 ( 1171 0 ) capacitor c=0.024152f //x=79.665 //y=5.02
c1167 ( 1170 0 ) capacitor c=0.024152f //x=78.785 //y=5.02
c1168 ( 1169 0 ) capacitor c=0.053132f //x=77.915 //y=5.02
c1169 ( 1168 0 ) capacitor c=0.0452179f //x=75.735 //y=5.02
c1170 ( 1167 0 ) capacitor c=0.0240372f //x=74.855 //y=5.02
c1171 ( 1166 0 ) capacitor c=0.0240372f //x=73.975 //y=5.02
c1172 ( 1165 0 ) capacitor c=0.0530795f //x=73.105 //y=5.02
c1173 ( 1164 0 ) capacitor c=0.0451031f //x=70.925 //y=5.02
c1174 ( 1163 0 ) capacitor c=0.0240372f //x=70.045 //y=5.02
c1175 ( 1162 0 ) capacitor c=0.0240372f //x=69.165 //y=5.02
c1176 ( 1161 0 ) capacitor c=0.0530795f //x=68.295 //y=5.02
c1177 ( 1160 0 ) capacitor c=0.0451031f //x=66.115 //y=5.02
c1178 ( 1159 0 ) capacitor c=0.0240372f //x=65.235 //y=5.02
c1179 ( 1158 0 ) capacitor c=0.0240372f //x=64.355 //y=5.02
c1180 ( 1157 0 ) capacitor c=0.0530795f //x=63.485 //y=5.02
c1181 ( 1156 0 ) capacitor c=0.0451031f //x=61.305 //y=5.02
c1182 ( 1155 0 ) capacitor c=0.0240372f //x=60.425 //y=5.02
c1183 ( 1154 0 ) capacitor c=0.0240372f //x=59.545 //y=5.02
c1184 ( 1153 0 ) capacitor c=0.0530795f //x=58.675 //y=5.02
c1185 ( 1152 0 ) capacitor c=0.0451031f //x=56.495 //y=5.02
c1186 ( 1151 0 ) capacitor c=0.0240372f //x=55.615 //y=5.02
c1187 ( 1150 0 ) capacitor c=0.0240372f //x=54.735 //y=5.02
c1188 ( 1149 0 ) capacitor c=0.0530795f //x=53.865 //y=5.02
c1189 ( 1148 0 ) capacitor c=0.0451031f //x=51.685 //y=5.02
c1190 ( 1147 0 ) capacitor c=0.0240372f //x=50.805 //y=5.02
c1191 ( 1146 0 ) capacitor c=0.0240372f //x=49.925 //y=5.02
c1192 ( 1145 0 ) capacitor c=0.0530795f //x=49.055 //y=5.02
c1193 ( 1144 0 ) capacitor c=0.0451031f //x=46.875 //y=5.02
c1194 ( 1143 0 ) capacitor c=0.0240372f //x=45.995 //y=5.02
c1195 ( 1142 0 ) capacitor c=0.0240372f //x=45.115 //y=5.02
c1196 ( 1141 0 ) capacitor c=0.0530795f //x=44.245 //y=5.02
c1197 ( 1140 0 ) capacitor c=0.0451031f //x=42.065 //y=5.02
c1198 ( 1139 0 ) capacitor c=0.0240372f //x=41.185 //y=5.02
c1199 ( 1138 0 ) capacitor c=0.0240372f //x=40.305 //y=5.02
c1200 ( 1137 0 ) capacitor c=0.0530795f //x=39.435 //y=5.02
c1201 ( 1136 0 ) capacitor c=0.0451031f //x=37.255 //y=5.02
c1202 ( 1135 0 ) capacitor c=0.0240372f //x=36.375 //y=5.02
c1203 ( 1134 0 ) capacitor c=0.0240372f //x=35.495 //y=5.02
c1204 ( 1133 0 ) capacitor c=0.0530795f //x=34.625 //y=5.02
c1205 ( 1132 0 ) capacitor c=0.0451031f //x=32.445 //y=5.02
c1206 ( 1131 0 ) capacitor c=0.0240372f //x=31.565 //y=5.02
c1207 ( 1130 0 ) capacitor c=0.0240372f //x=30.685 //y=5.02
c1208 ( 1129 0 ) capacitor c=0.0530795f //x=29.815 //y=5.02
c1209 ( 1128 0 ) capacitor c=0.0451031f //x=27.635 //y=5.02
c1210 ( 1127 0 ) capacitor c=0.0240372f //x=26.755 //y=5.02
c1211 ( 1126 0 ) capacitor c=0.0240372f //x=25.875 //y=5.02
c1212 ( 1125 0 ) capacitor c=0.0530795f //x=25.005 //y=5.02
c1213 ( 1124 0 ) capacitor c=0.0452179f //x=22.825 //y=5.02
c1214 ( 1123 0 ) capacitor c=0.024152f //x=21.945 //y=5.02
c1215 ( 1122 0 ) capacitor c=0.024152f //x=21.065 //y=5.02
c1216 ( 1121 0 ) capacitor c=0.053132f //x=20.195 //y=5.02
c1217 ( 1120 0 ) capacitor c=0.0452179f //x=18.015 //y=5.02
c1218 ( 1119 0 ) capacitor c=0.024152f //x=17.135 //y=5.02
c1219 ( 1118 0 ) capacitor c=0.024152f //x=16.255 //y=5.02
c1220 ( 1117 0 ) capacitor c=0.053132f //x=15.385 //y=5.02
c1221 ( 1116 0 ) capacitor c=0.0452179f //x=13.205 //y=5.02
c1222 ( 1115 0 ) capacitor c=0.024152f //x=12.325 //y=5.02
c1223 ( 1114 0 ) capacitor c=0.024152f //x=11.445 //y=5.02
c1224 ( 1113 0 ) capacitor c=0.053132f //x=10.575 //y=5.02
c1225 ( 1112 0 ) capacitor c=0.0452179f //x=8.395 //y=5.02
c1226 ( 1111 0 ) capacitor c=0.024152f //x=7.515 //y=5.02
c1227 ( 1110 0 ) capacitor c=0.02424f //x=6.635 //y=5.02
c1228 ( 1109 0 ) capacitor c=0.0531793f //x=5.765 //y=5.02
c1229 ( 1108 0 ) capacitor c=0.0453059f //x=3.585 //y=5.02
c1230 ( 1107 0 ) capacitor c=0.02424f //x=2.705 //y=5.02
c1231 ( 1106 0 ) capacitor c=0.02424f //x=1.825 //y=5.02
c1232 ( 1105 0 ) capacitor c=0.0531407f //x=0.955 //y=5.02
c1233 ( 1104 0 ) capacitor c=0.113329f //x=93.24 //y=7.4
c1234 ( 1103 0 ) capacitor c=0.121389f //x=89.91 //y=7.4
c1235 ( 1102 0 ) capacitor c=0.00591168f //x=89.13 //y=7.4
c1236 ( 1101 0 ) capacitor c=0.00591168f //x=88.25 //y=7.4
c1237 ( 1100 0 ) capacitor c=0.00591168f //x=87.32 //y=7.4
c1238 ( 1098 0 ) capacitor c=0.132974f //x=86.58 //y=7.4
c1239 ( 1097 0 ) capacitor c=0.00591168f //x=85.5 //y=7.4
c1240 ( 1096 0 ) capacitor c=0.00591168f //x=84.62 //y=7.4
c1241 ( 1095 0 ) capacitor c=0.00591168f //x=83.74 //y=7.4
c1242 ( 1094 0 ) capacitor c=0.00591168f //x=82.86 //y=7.4
c1243 ( 1093 0 ) capacitor c=0.155236f //x=81.77 //y=7.4
c1244 ( 1092 0 ) capacitor c=0.00591168f //x=80.69 //y=7.4
c1245 ( 1091 0 ) capacitor c=0.00591168f //x=79.81 //y=7.4
c1246 ( 1090 0 ) capacitor c=0.00591168f //x=78.93 //y=7.4
c1247 ( 1089 0 ) capacitor c=0.00591168f //x=78.05 //y=7.4
c1248 ( 1088 0 ) capacitor c=0.154686f //x=76.96 //y=7.4
c1249 ( 1087 0 ) capacitor c=0.00591168f //x=75.88 //y=7.4
c1250 ( 1086 0 ) capacitor c=0.00591168f //x=75 //y=7.4
c1251 ( 1085 0 ) capacitor c=0.00591168f //x=74.12 //y=7.4
c1252 ( 1084 0 ) capacitor c=0.00591168f //x=73.24 //y=7.4
c1253 ( 1083 0 ) capacitor c=0.153722f //x=72.15 //y=7.4
c1254 ( 1082 0 ) capacitor c=0.00591168f //x=71.07 //y=7.4
c1255 ( 1081 0 ) capacitor c=0.00591168f //x=70.19 //y=7.4
c1256 ( 1080 0 ) capacitor c=0.00591168f //x=69.31 //y=7.4
c1257 ( 1079 0 ) capacitor c=0.00591168f //x=68.43 //y=7.4
c1258 ( 1078 0 ) capacitor c=0.153803f //x=67.34 //y=7.4
c1259 ( 1077 0 ) capacitor c=0.00591168f //x=66.26 //y=7.4
c1260 ( 1076 0 ) capacitor c=0.00591168f //x=65.38 //y=7.4
c1261 ( 1075 0 ) capacitor c=0.00591168f //x=64.5 //y=7.4
c1262 ( 1074 0 ) capacitor c=0.00591168f //x=63.62 //y=7.4
c1263 ( 1073 0 ) capacitor c=0.158289f //x=62.53 //y=7.4
c1264 ( 1072 0 ) capacitor c=0.00591168f //x=61.45 //y=7.4
c1265 ( 1071 0 ) capacitor c=0.00591168f //x=60.57 //y=7.4
c1266 ( 1070 0 ) capacitor c=0.00591168f //x=59.69 //y=7.4
c1267 ( 1069 0 ) capacitor c=0.00591168f //x=58.81 //y=7.4
c1268 ( 1068 0 ) capacitor c=0.15374f //x=57.72 //y=7.4
c1269 ( 1067 0 ) capacitor c=0.00591168f //x=56.64 //y=7.4
c1270 ( 1066 0 ) capacitor c=0.00591168f //x=55.76 //y=7.4
c1271 ( 1065 0 ) capacitor c=0.00591168f //x=54.88 //y=7.4
c1272 ( 1064 0 ) capacitor c=0.00591168f //x=54 //y=7.4
c1273 ( 1063 0 ) capacitor c=0.15385f //x=52.91 //y=7.4
c1274 ( 1062 0 ) capacitor c=0.00591168f //x=51.83 //y=7.4
c1275 ( 1061 0 ) capacitor c=0.00591168f //x=50.95 //y=7.4
c1276 ( 1060 0 ) capacitor c=0.00591168f //x=50.07 //y=7.4
c1277 ( 1059 0 ) capacitor c=0.00591168f //x=49.19 //y=7.4
c1278 ( 1058 0 ) capacitor c=0.153803f //x=48.1 //y=7.4
c1279 ( 1057 0 ) capacitor c=0.00591168f //x=47.02 //y=7.4
c1280 ( 1056 0 ) capacitor c=0.00591168f //x=46.14 //y=7.4
c1281 ( 1055 0 ) capacitor c=0.00591168f //x=45.26 //y=7.4
c1282 ( 1054 0 ) capacitor c=0.00591168f //x=44.38 //y=7.4
c1283 ( 1053 0 ) capacitor c=0.153779f //x=43.29 //y=7.4
c1284 ( 1052 0 ) capacitor c=0.00591168f //x=42.21 //y=7.4
c1285 ( 1051 0 ) capacitor c=0.00591168f //x=41.33 //y=7.4
c1286 ( 1050 0 ) capacitor c=0.00591168f //x=40.45 //y=7.4
c1287 ( 1049 0 ) capacitor c=0.00591168f //x=39.57 //y=7.4
c1288 ( 1048 0 ) capacitor c=0.153803f //x=38.48 //y=7.4
c1289 ( 1047 0 ) capacitor c=0.00591168f //x=37.4 //y=7.4
c1290 ( 1046 0 ) capacitor c=0.00591168f //x=36.52 //y=7.4
c1291 ( 1045 0 ) capacitor c=0.00591168f //x=35.64 //y=7.4
c1292 ( 1044 0 ) capacitor c=0.00591168f //x=34.76 //y=7.4
c1293 ( 1043 0 ) capacitor c=0.153957f //x=33.67 //y=7.4
c1294 ( 1042 0 ) capacitor c=0.00591168f //x=32.59 //y=7.4
c1295 ( 1041 0 ) capacitor c=0.00591168f //x=31.71 //y=7.4
c1296 ( 1040 0 ) capacitor c=0.00591168f //x=30.83 //y=7.4
c1297 ( 1039 0 ) capacitor c=0.00591168f //x=29.95 //y=7.4
c1298 ( 1038 0 ) capacitor c=0.154054f //x=28.86 //y=7.4
c1299 ( 1037 0 ) capacitor c=0.00591168f //x=27.78 //y=7.4
c1300 ( 1036 0 ) capacitor c=0.00591168f //x=26.9 //y=7.4
c1301 ( 1035 0 ) capacitor c=0.00591168f //x=26.02 //y=7.4
c1302 ( 1034 0 ) capacitor c=0.00591168f //x=25.14 //y=7.4
c1303 ( 1033 0 ) capacitor c=0.153632f //x=24.05 //y=7.4
c1304 ( 1032 0 ) capacitor c=0.00591168f //x=22.97 //y=7.4
c1305 ( 1031 0 ) capacitor c=0.00591168f //x=22.09 //y=7.4
c1306 ( 1030 0 ) capacitor c=0.00591168f //x=21.21 //y=7.4
c1307 ( 1029 0 ) capacitor c=0.00591168f //x=20.33 //y=7.4
c1308 ( 1028 0 ) capacitor c=0.15519f //x=19.24 //y=7.4
c1309 ( 1027 0 ) capacitor c=0.00591168f //x=18.16 //y=7.4
c1310 ( 1026 0 ) capacitor c=0.00591168f //x=17.28 //y=7.4
c1311 ( 1025 0 ) capacitor c=0.00591168f //x=16.4 //y=7.4
c1312 ( 1024 0 ) capacitor c=0.00591168f //x=15.52 //y=7.4
c1313 ( 1023 0 ) capacitor c=0.155166f //x=14.43 //y=7.4
c1314 ( 1022 0 ) capacitor c=0.00591168f //x=13.35 //y=7.4
c1315 ( 1021 0 ) capacitor c=0.00591168f //x=12.47 //y=7.4
c1316 ( 1020 0 ) capacitor c=0.00591168f //x=11.59 //y=7.4
c1317 ( 1019 0 ) capacitor c=0.00591168f //x=10.71 //y=7.4
c1318 ( 1018 0 ) capacitor c=0.15519f //x=9.62 //y=7.4
c1319 ( 1017 0 ) capacitor c=0.00591168f //x=8.54 //y=7.4
c1320 ( 1016 0 ) capacitor c=0.00591168f //x=7.66 //y=7.4
c1321 ( 1015 0 ) capacitor c=0.00591168f //x=6.78 //y=7.4
c1322 ( 1014 0 ) capacitor c=0.00591168f //x=5.9 //y=7.4
c1323 ( 1013 0 ) capacitor c=0.157289f //x=4.81 //y=7.4
c1324 ( 1012 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c1325 ( 1011 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c1326 ( 1010 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c1327 ( 1009 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c1328 ( 1006 0 ) capacitor c=0.333243f //x=95.83 //y=7.4
c1329 ( 991 0 ) capacitor c=0.120978f //x=93.07 //y=7.4
c1330 ( 985 0 ) capacitor c=0.0236224f //x=89.74 //y=7.4
c1331 ( 975 0 ) capacitor c=0.028539f //x=89.045 //y=7.4
c1332 ( 967 0 ) capacitor c=0.0285075f //x=88.165 //y=7.4
c1333 ( 959 0 ) capacitor c=0.0240981f //x=87.285 //y=7.4
c1334 ( 953 0 ) capacitor c=0.0394667f //x=86.41 //y=7.4
c1335 ( 943 0 ) capacitor c=0.0288488f //x=85.415 //y=7.4
c1336 ( 935 0 ) capacitor c=0.0287514f //x=84.535 //y=7.4
c1337 ( 925 0 ) capacitor c=0.0284966f //x=83.655 //y=7.4
c1338 ( 915 0 ) capacitor c=0.0383672f //x=82.775 //y=7.4
c1339 ( 909 0 ) capacitor c=0.0394667f //x=81.6 //y=7.4
c1340 ( 899 0 ) capacitor c=0.0288488f //x=80.605 //y=7.4
c1341 ( 891 0 ) capacitor c=0.0287514f //x=79.725 //y=7.4
c1342 ( 881 0 ) capacitor c=0.0284966f //x=78.845 //y=7.4
c1343 ( 871 0 ) capacitor c=0.0383672f //x=77.965 //y=7.4
c1344 ( 865 0 ) capacitor c=0.0394667f //x=76.79 //y=7.4
c1345 ( 855 0 ) capacitor c=0.0288466f //x=75.795 //y=7.4
c1346 ( 847 0 ) capacitor c=0.028724f //x=74.915 //y=7.4
c1347 ( 837 0 ) capacitor c=0.0284804f //x=74.035 //y=7.4
c1348 ( 827 0 ) capacitor c=0.0383672f //x=73.155 //y=7.4
c1349 ( 821 0 ) capacitor c=0.0394025f //x=71.98 //y=7.4
c1350 ( 811 0 ) capacitor c=0.0288171f //x=70.985 //y=7.4
c1351 ( 803 0 ) capacitor c=0.028724f //x=70.105 //y=7.4
c1352 ( 793 0 ) capacitor c=0.0284804f //x=69.225 //y=7.4
c1353 ( 783 0 ) capacitor c=0.0383672f //x=68.345 //y=7.4
c1354 ( 777 0 ) capacitor c=0.0394025f //x=67.17 //y=7.4
c1355 ( 767 0 ) capacitor c=0.0288171f //x=66.175 //y=7.4
c1356 ( 759 0 ) capacitor c=0.028724f //x=65.295 //y=7.4
c1357 ( 749 0 ) capacitor c=0.0284804f //x=64.415 //y=7.4
c1358 ( 739 0 ) capacitor c=0.0383672f //x=63.535 //y=7.4
c1359 ( 733 0 ) capacitor c=0.0394025f //x=62.36 //y=7.4
c1360 ( 723 0 ) capacitor c=0.0288171f //x=61.365 //y=7.4
c1361 ( 715 0 ) capacitor c=0.028724f //x=60.485 //y=7.4
c1362 ( 705 0 ) capacitor c=0.0284804f //x=59.605 //y=7.4
c1363 ( 695 0 ) capacitor c=0.0383672f //x=58.725 //y=7.4
c1364 ( 689 0 ) capacitor c=0.0394025f //x=57.55 //y=7.4
c1365 ( 679 0 ) capacitor c=0.0288171f //x=56.555 //y=7.4
c1366 ( 671 0 ) capacitor c=0.028724f //x=55.675 //y=7.4
c1367 ( 661 0 ) capacitor c=0.0284804f //x=54.795 //y=7.4
c1368 ( 651 0 ) capacitor c=0.0383672f //x=53.915 //y=7.4
c1369 ( 645 0 ) capacitor c=0.0394025f //x=52.74 //y=7.4
c1370 ( 635 0 ) capacitor c=0.0288171f //x=51.745 //y=7.4
c1371 ( 627 0 ) capacitor c=0.028724f //x=50.865 //y=7.4
c1372 ( 617 0 ) capacitor c=0.0284804f //x=49.985 //y=7.4
c1373 ( 607 0 ) capacitor c=0.0383672f //x=49.105 //y=7.4
c1374 ( 601 0 ) capacitor c=0.0394025f //x=47.93 //y=7.4
c1375 ( 591 0 ) capacitor c=0.0288171f //x=46.935 //y=7.4
c1376 ( 583 0 ) capacitor c=0.028724f //x=46.055 //y=7.4
c1377 ( 573 0 ) capacitor c=0.0284804f //x=45.175 //y=7.4
c1378 ( 563 0 ) capacitor c=0.0383672f //x=44.295 //y=7.4
c1379 ( 557 0 ) capacitor c=0.0394025f //x=43.12 //y=7.4
c1380 ( 547 0 ) capacitor c=0.0288171f //x=42.125 //y=7.4
c1381 ( 539 0 ) capacitor c=0.028724f //x=41.245 //y=7.4
c1382 ( 529 0 ) capacitor c=0.0284804f //x=40.365 //y=7.4
c1383 ( 519 0 ) capacitor c=0.0383672f //x=39.485 //y=7.4
c1384 ( 513 0 ) capacitor c=0.0394025f //x=38.31 //y=7.4
c1385 ( 503 0 ) capacitor c=0.0288171f //x=37.315 //y=7.4
c1386 ( 495 0 ) capacitor c=0.028724f //x=36.435 //y=7.4
c1387 ( 485 0 ) capacitor c=0.0284804f //x=35.555 //y=7.4
c1388 ( 475 0 ) capacitor c=0.0383672f //x=34.675 //y=7.4
c1389 ( 469 0 ) capacitor c=0.0394025f //x=33.5 //y=7.4
c1390 ( 459 0 ) capacitor c=0.0288171f //x=32.505 //y=7.4
c1391 ( 451 0 ) capacitor c=0.028724f //x=31.625 //y=7.4
c1392 ( 441 0 ) capacitor c=0.0284804f //x=30.745 //y=7.4
c1393 ( 431 0 ) capacitor c=0.0383672f //x=29.865 //y=7.4
c1394 ( 425 0 ) capacitor c=0.0394025f //x=28.69 //y=7.4
c1395 ( 415 0 ) capacitor c=0.0288171f //x=27.695 //y=7.4
c1396 ( 407 0 ) capacitor c=0.028724f //x=26.815 //y=7.4
c1397 ( 397 0 ) capacitor c=0.0284804f //x=25.935 //y=7.4
c1398 ( 387 0 ) capacitor c=0.0383672f //x=25.055 //y=7.4
c1399 ( 381 0 ) capacitor c=0.0394119f //x=23.88 //y=7.4
c1400 ( 371 0 ) capacitor c=0.0288488f //x=22.885 //y=7.4
c1401 ( 363 0 ) capacitor c=0.0287514f //x=22.005 //y=7.4
c1402 ( 353 0 ) capacitor c=0.0284966f //x=21.125 //y=7.4
c1403 ( 343 0 ) capacitor c=0.0383672f //x=20.245 //y=7.4
c1404 ( 337 0 ) capacitor c=0.0394667f //x=19.07 //y=7.4
c1405 ( 327 0 ) capacitor c=0.0288488f //x=18.075 //y=7.4
c1406 ( 319 0 ) capacitor c=0.0287505f //x=17.195 //y=7.4
c1407 ( 309 0 ) capacitor c=0.0284966f //x=16.315 //y=7.4
c1408 ( 299 0 ) capacitor c=0.0383672f //x=15.435 //y=7.4
c1409 ( 293 0 ) capacitor c=0.0394667f //x=14.26 //y=7.4
c1410 ( 283 0 ) capacitor c=0.0288488f //x=13.265 //y=7.4
c1411 ( 275 0 ) capacitor c=0.0287514f //x=12.385 //y=7.4
c1412 ( 265 0 ) capacitor c=0.0284966f //x=11.505 //y=7.4
c1413 ( 255 0 ) capacitor c=0.0383672f //x=10.625 //y=7.4
c1414 ( 249 0 ) capacitor c=0.0394667f //x=9.45 //y=7.4
c1415 ( 239 0 ) capacitor c=0.0288488f //x=8.455 //y=7.4
c1416 ( 231 0 ) capacitor c=0.0287505f //x=7.575 //y=7.4
c1417 ( 221 0 ) capacitor c=0.028511f //x=6.695 //y=7.4
c1418 ( 211 0 ) capacitor c=0.0383672f //x=5.815 //y=7.4
c1419 ( 205 0 ) capacitor c=0.0395236f //x=4.64 //y=7.4
c1420 ( 195 0 ) capacitor c=0.0288769f //x=3.645 //y=7.4
c1421 ( 187 0 ) capacitor c=0.0287757f //x=2.765 //y=7.4
c1422 ( 177 0 ) capacitor c=0.028511f //x=1.885 //y=7.4
c1423 ( 170 0 ) capacitor c=0.234727f //x=0.74 //y=7.4
c1424 ( 167 0 ) capacitor c=0.0441843f //x=1.005 //y=7.4
c1425 ( 163 0 ) capacitor c=3.17938f //x=95.83 //y=7.4
r1426 (  1004 1006 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=94.72 //y=7.4 //x2=95.83 //y2=7.4
r1427 (  1002 1004 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=93.61 //y=7.4 //x2=94.72 //y2=7.4
r1428 (  1000 1104 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=93.41 //y=7.4 //x2=93.24 //y2=7.4
r1429 (  1000 1002 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=93.41 //y=7.4 //x2=93.61 //y2=7.4
r1430 (  994 996 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=91.02 //y=7.4 //x2=92.13 //y2=7.4
r1431 (  992 1103 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=90.08 //y=7.4 //x2=89.91 //y2=7.4
r1432 (  992 994 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=90.08 //y=7.4 //x2=91.02 //y2=7.4
r1433 (  991 1104 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=93.07 //y=7.4 //x2=93.24 //y2=7.4
r1434 (  991 996 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=93.07 //y=7.4 //x2=92.13 //y2=7.4
r1435 (  986 1102 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=89.215 //y=7.4 //x2=89.13 //y2=7.4
r1436 (  986 988 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=89.215 //y=7.4 //x2=89.54 //y2=7.4
r1437 (  985 1103 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=89.74 //y=7.4 //x2=89.91 //y2=7.4
r1438 (  985 988 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=89.74 //y=7.4 //x2=89.54 //y2=7.4
r1439 (  979 1102 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=89.13 //y=7.23 //x2=89.13 //y2=7.4
r1440 (  979 1179 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=89.13 //y=7.23 //x2=89.13 //y2=6.4
r1441 (  976 1101 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=88.335 //y=7.4 //x2=88.25 //y2=7.4
r1442 (  976 978 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=88.335 //y=7.4 //x2=88.43 //y2=7.4
r1443 (  975 1102 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=89.045 //y=7.4 //x2=89.13 //y2=7.4
r1444 (  975 978 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=89.045 //y=7.4 //x2=88.43 //y2=7.4
r1445 (  969 1101 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=88.25 //y=7.23 //x2=88.25 //y2=7.4
r1446 (  969 1178 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=88.25 //y=7.23 //x2=88.25 //y2=6.74
r1447 (  968 1100 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=87.455 //y=7.4 //x2=87.37 //y2=7.4
r1448 (  967 1101 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=88.165 //y=7.4 //x2=88.25 //y2=7.4
r1449 (  967 968 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=88.165 //y=7.4 //x2=87.455 //y2=7.4
r1450 (  961 1100 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=87.37 //y=7.23 //x2=87.37 //y2=7.4
r1451 (  961 1177 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=87.37 //y=7.23 //x2=87.37 //y2=6.4
r1452 (  960 1098 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=86.75 //y=7.4 //x2=86.58 //y2=7.4
r1453 (  959 1100 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=87.285 //y=7.4 //x2=87.37 //y2=7.4
r1454 (  959 960 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=87.285 //y=7.4 //x2=86.75 //y2=7.4
r1455 (  954 1097 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.585 //y=7.4 //x2=85.5 //y2=7.4
r1456 (  954 956 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=85.585 //y=7.4 //x2=85.84 //y2=7.4
r1457 (  953 1098 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=86.41 //y=7.4 //x2=86.58 //y2=7.4
r1458 (  953 956 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=86.41 //y=7.4 //x2=85.84 //y2=7.4
r1459 (  947 1097 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=85.5 //y=7.23 //x2=85.5 //y2=7.4
r1460 (  947 1176 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=85.5 //y=7.23 //x2=85.5 //y2=6.745
r1461 (  944 1096 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.705 //y=7.4 //x2=84.62 //y2=7.4
r1462 (  944 946 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=84.705 //y=7.4 //x2=84.73 //y2=7.4
r1463 (  943 1097 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.415 //y=7.4 //x2=85.5 //y2=7.4
r1464 (  943 946 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=85.415 //y=7.4 //x2=84.73 //y2=7.4
r1465 (  937 1096 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=84.62 //y=7.23 //x2=84.62 //y2=7.4
r1466 (  937 1175 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=84.62 //y=7.23 //x2=84.62 //y2=6.745
r1467 (  936 1095 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.825 //y=7.4 //x2=83.74 //y2=7.4
r1468 (  935 1096 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.535 //y=7.4 //x2=84.62 //y2=7.4
r1469 (  935 936 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=84.535 //y=7.4 //x2=83.825 //y2=7.4
r1470 (  929 1095 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=83.74 //y=7.23 //x2=83.74 //y2=7.4
r1471 (  929 1174 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=83.74 //y=7.23 //x2=83.74 //y2=6.745
r1472 (  926 1094 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.945 //y=7.4 //x2=82.86 //y2=7.4
r1473 (  926 928 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=82.945 //y=7.4 //x2=83.62 //y2=7.4
r1474 (  925 1095 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.655 //y=7.4 //x2=83.74 //y2=7.4
r1475 (  925 928 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=83.655 //y=7.4 //x2=83.62 //y2=7.4
r1476 (  919 1094 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=82.86 //y=7.23 //x2=82.86 //y2=7.4
r1477 (  919 1173 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=82.86 //y=7.23 //x2=82.86 //y2=6.405
r1478 (  916 1093 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.94 //y=7.4 //x2=81.77 //y2=7.4
r1479 (  916 918 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=81.94 //y=7.4 //x2=82.51 //y2=7.4
r1480 (  915 1094 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.775 //y=7.4 //x2=82.86 //y2=7.4
r1481 (  915 918 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=82.775 //y=7.4 //x2=82.51 //y2=7.4
r1482 (  910 1092 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.775 //y=7.4 //x2=80.69 //y2=7.4
r1483 (  910 912 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=80.775 //y=7.4 //x2=81.03 //y2=7.4
r1484 (  909 1093 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.6 //y=7.4 //x2=81.77 //y2=7.4
r1485 (  909 912 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=81.6 //y=7.4 //x2=81.03 //y2=7.4
r1486 (  903 1092 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=80.69 //y=7.23 //x2=80.69 //y2=7.4
r1487 (  903 1172 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=80.69 //y=7.23 //x2=80.69 //y2=6.745
r1488 (  900 1091 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.895 //y=7.4 //x2=79.81 //y2=7.4
r1489 (  900 902 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=79.895 //y=7.4 //x2=79.92 //y2=7.4
r1490 (  899 1092 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.605 //y=7.4 //x2=80.69 //y2=7.4
r1491 (  899 902 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=80.605 //y=7.4 //x2=79.92 //y2=7.4
r1492 (  893 1091 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=79.81 //y=7.23 //x2=79.81 //y2=7.4
r1493 (  893 1171 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=79.81 //y=7.23 //x2=79.81 //y2=6.745
r1494 (  892 1090 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.015 //y=7.4 //x2=78.93 //y2=7.4
r1495 (  891 1091 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.725 //y=7.4 //x2=79.81 //y2=7.4
r1496 (  891 892 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=79.725 //y=7.4 //x2=79.015 //y2=7.4
r1497 (  885 1090 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=78.93 //y=7.23 //x2=78.93 //y2=7.4
r1498 (  885 1170 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=78.93 //y=7.23 //x2=78.93 //y2=6.745
r1499 (  882 1089 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.135 //y=7.4 //x2=78.05 //y2=7.4
r1500 (  882 884 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=78.135 //y=7.4 //x2=78.81 //y2=7.4
r1501 (  881 1090 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.845 //y=7.4 //x2=78.93 //y2=7.4
r1502 (  881 884 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=78.845 //y=7.4 //x2=78.81 //y2=7.4
r1503 (  875 1089 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=78.05 //y=7.23 //x2=78.05 //y2=7.4
r1504 (  875 1169 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=78.05 //y=7.23 //x2=78.05 //y2=6.405
r1505 (  872 1088 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.13 //y=7.4 //x2=76.96 //y2=7.4
r1506 (  872 874 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=77.13 //y=7.4 //x2=77.7 //y2=7.4
r1507 (  871 1089 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.965 //y=7.4 //x2=78.05 //y2=7.4
r1508 (  871 874 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=77.965 //y=7.4 //x2=77.7 //y2=7.4
r1509 (  866 1087 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.965 //y=7.4 //x2=75.88 //y2=7.4
r1510 (  866 868 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=75.965 //y=7.4 //x2=76.22 //y2=7.4
r1511 (  865 1088 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.79 //y=7.4 //x2=76.96 //y2=7.4
r1512 (  865 868 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=76.79 //y=7.4 //x2=76.22 //y2=7.4
r1513 (  859 1087 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=75.88 //y=7.23 //x2=75.88 //y2=7.4
r1514 (  859 1168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=75.88 //y=7.23 //x2=75.88 //y2=6.745
r1515 (  856 1086 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.085 //y=7.4 //x2=75 //y2=7.4
r1516 (  856 858 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=75.085 //y=7.4 //x2=75.11 //y2=7.4
r1517 (  855 1087 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.795 //y=7.4 //x2=75.88 //y2=7.4
r1518 (  855 858 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=75.795 //y=7.4 //x2=75.11 //y2=7.4
r1519 (  849 1086 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=75 //y=7.23 //x2=75 //y2=7.4
r1520 (  849 1167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=75 //y=7.23 //x2=75 //y2=6.745
r1521 (  848 1085 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.205 //y=7.4 //x2=74.12 //y2=7.4
r1522 (  847 1086 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.915 //y=7.4 //x2=75 //y2=7.4
r1523 (  847 848 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=74.915 //y=7.4 //x2=74.205 //y2=7.4
r1524 (  841 1085 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.12 //y=7.23 //x2=74.12 //y2=7.4
r1525 (  841 1166 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=74.12 //y=7.23 //x2=74.12 //y2=6.745
r1526 (  838 1084 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.325 //y=7.4 //x2=73.24 //y2=7.4
r1527 (  838 840 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=73.325 //y=7.4 //x2=74 //y2=7.4
r1528 (  837 1085 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.035 //y=7.4 //x2=74.12 //y2=7.4
r1529 (  837 840 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=74.035 //y=7.4 //x2=74 //y2=7.4
r1530 (  831 1084 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.24 //y=7.23 //x2=73.24 //y2=7.4
r1531 (  831 1165 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=73.24 //y=7.23 //x2=73.24 //y2=6.405
r1532 (  828 1083 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=72.32 //y=7.4 //x2=72.15 //y2=7.4
r1533 (  828 830 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=72.32 //y=7.4 //x2=72.89 //y2=7.4
r1534 (  827 1084 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.155 //y=7.4 //x2=73.24 //y2=7.4
r1535 (  827 830 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=73.155 //y=7.4 //x2=72.89 //y2=7.4
r1536 (  822 1082 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.155 //y=7.4 //x2=71.07 //y2=7.4
r1537 (  822 824 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=71.155 //y=7.4 //x2=71.41 //y2=7.4
r1538 (  821 1083 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.98 //y=7.4 //x2=72.15 //y2=7.4
r1539 (  821 824 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=71.98 //y=7.4 //x2=71.41 //y2=7.4
r1540 (  815 1082 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.07 //y=7.23 //x2=71.07 //y2=7.4
r1541 (  815 1164 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=71.07 //y=7.23 //x2=71.07 //y2=6.745
r1542 (  812 1081 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.275 //y=7.4 //x2=70.19 //y2=7.4
r1543 (  812 814 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=70.275 //y=7.4 //x2=70.3 //y2=7.4
r1544 (  811 1082 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.985 //y=7.4 //x2=71.07 //y2=7.4
r1545 (  811 814 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=70.985 //y=7.4 //x2=70.3 //y2=7.4
r1546 (  805 1081 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=70.19 //y=7.23 //x2=70.19 //y2=7.4
r1547 (  805 1163 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=70.19 //y=7.23 //x2=70.19 //y2=6.745
r1548 (  804 1080 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.395 //y=7.4 //x2=69.31 //y2=7.4
r1549 (  803 1081 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.105 //y=7.4 //x2=70.19 //y2=7.4
r1550 (  803 804 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=70.105 //y=7.4 //x2=69.395 //y2=7.4
r1551 (  797 1080 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.31 //y=7.23 //x2=69.31 //y2=7.4
r1552 (  797 1162 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=69.31 //y=7.23 //x2=69.31 //y2=6.745
r1553 (  794 1079 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.515 //y=7.4 //x2=68.43 //y2=7.4
r1554 (  794 796 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=68.515 //y=7.4 //x2=69.19 //y2=7.4
r1555 (  793 1080 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.225 //y=7.4 //x2=69.31 //y2=7.4
r1556 (  793 796 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=69.225 //y=7.4 //x2=69.19 //y2=7.4
r1557 (  787 1079 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.43 //y=7.23 //x2=68.43 //y2=7.4
r1558 (  787 1161 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=68.43 //y=7.23 //x2=68.43 //y2=6.405
r1559 (  784 1078 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.51 //y=7.4 //x2=67.34 //y2=7.4
r1560 (  784 786 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.51 //y=7.4 //x2=68.08 //y2=7.4
r1561 (  783 1079 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.345 //y=7.4 //x2=68.43 //y2=7.4
r1562 (  783 786 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=68.345 //y=7.4 //x2=68.08 //y2=7.4
r1563 (  778 1077 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.345 //y=7.4 //x2=66.26 //y2=7.4
r1564 (  778 780 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=66.345 //y=7.4 //x2=66.6 //y2=7.4
r1565 (  777 1078 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.17 //y=7.4 //x2=67.34 //y2=7.4
r1566 (  777 780 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.17 //y=7.4 //x2=66.6 //y2=7.4
r1567 (  771 1077 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=66.26 //y=7.23 //x2=66.26 //y2=7.4
r1568 (  771 1160 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=66.26 //y=7.23 //x2=66.26 //y2=6.745
r1569 (  768 1076 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.465 //y=7.4 //x2=65.38 //y2=7.4
r1570 (  768 770 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=65.465 //y=7.4 //x2=65.49 //y2=7.4
r1571 (  767 1077 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.175 //y=7.4 //x2=66.26 //y2=7.4
r1572 (  767 770 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=66.175 //y=7.4 //x2=65.49 //y2=7.4
r1573 (  761 1076 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.38 //y=7.23 //x2=65.38 //y2=7.4
r1574 (  761 1159 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=65.38 //y=7.23 //x2=65.38 //y2=6.745
r1575 (  760 1075 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.585 //y=7.4 //x2=64.5 //y2=7.4
r1576 (  759 1076 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.295 //y=7.4 //x2=65.38 //y2=7.4
r1577 (  759 760 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=65.295 //y=7.4 //x2=64.585 //y2=7.4
r1578 (  753 1075 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.5 //y=7.23 //x2=64.5 //y2=7.4
r1579 (  753 1158 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=64.5 //y=7.23 //x2=64.5 //y2=6.745
r1580 (  750 1074 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.705 //y=7.4 //x2=63.62 //y2=7.4
r1581 (  750 752 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=63.705 //y=7.4 //x2=64.38 //y2=7.4
r1582 (  749 1075 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.415 //y=7.4 //x2=64.5 //y2=7.4
r1583 (  749 752 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=64.415 //y=7.4 //x2=64.38 //y2=7.4
r1584 (  743 1074 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=63.62 //y=7.23 //x2=63.62 //y2=7.4
r1585 (  743 1157 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=63.62 //y=7.23 //x2=63.62 //y2=6.405
r1586 (  740 1073 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.7 //y=7.4 //x2=62.53 //y2=7.4
r1587 (  740 742 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=62.7 //y=7.4 //x2=63.27 //y2=7.4
r1588 (  739 1074 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.535 //y=7.4 //x2=63.62 //y2=7.4
r1589 (  739 742 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=63.535 //y=7.4 //x2=63.27 //y2=7.4
r1590 (  734 1072 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.535 //y=7.4 //x2=61.45 //y2=7.4
r1591 (  734 736 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=61.535 //y=7.4 //x2=61.79 //y2=7.4
r1592 (  733 1073 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.36 //y=7.4 //x2=62.53 //y2=7.4
r1593 (  733 736 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=62.36 //y=7.4 //x2=61.79 //y2=7.4
r1594 (  727 1072 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.45 //y=7.23 //x2=61.45 //y2=7.4
r1595 (  727 1156 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=61.45 //y=7.23 //x2=61.45 //y2=6.745
r1596 (  724 1071 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.655 //y=7.4 //x2=60.57 //y2=7.4
r1597 (  724 726 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=60.655 //y=7.4 //x2=60.68 //y2=7.4
r1598 (  723 1072 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.365 //y=7.4 //x2=61.45 //y2=7.4
r1599 (  723 726 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=61.365 //y=7.4 //x2=60.68 //y2=7.4
r1600 (  717 1071 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=60.57 //y=7.23 //x2=60.57 //y2=7.4
r1601 (  717 1155 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.57 //y=7.23 //x2=60.57 //y2=6.745
r1602 (  716 1070 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.775 //y=7.4 //x2=59.69 //y2=7.4
r1603 (  715 1071 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.485 //y=7.4 //x2=60.57 //y2=7.4
r1604 (  715 716 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=60.485 //y=7.4 //x2=59.775 //y2=7.4
r1605 (  709 1070 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=59.69 //y=7.23 //x2=59.69 //y2=7.4
r1606 (  709 1154 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.69 //y=7.23 //x2=59.69 //y2=6.745
r1607 (  706 1069 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.895 //y=7.4 //x2=58.81 //y2=7.4
r1608 (  706 708 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=58.895 //y=7.4 //x2=59.57 //y2=7.4
r1609 (  705 1070 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.605 //y=7.4 //x2=59.69 //y2=7.4
r1610 (  705 708 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=59.605 //y=7.4 //x2=59.57 //y2=7.4
r1611 (  699 1069 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.81 //y=7.23 //x2=58.81 //y2=7.4
r1612 (  699 1153 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=58.81 //y=7.23 //x2=58.81 //y2=6.405
r1613 (  696 1068 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.89 //y=7.4 //x2=57.72 //y2=7.4
r1614 (  696 698 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=57.89 //y=7.4 //x2=58.46 //y2=7.4
r1615 (  695 1069 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.725 //y=7.4 //x2=58.81 //y2=7.4
r1616 (  695 698 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=58.725 //y=7.4 //x2=58.46 //y2=7.4
r1617 (  690 1067 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.725 //y=7.4 //x2=56.64 //y2=7.4
r1618 (  690 692 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=56.725 //y=7.4 //x2=56.98 //y2=7.4
r1619 (  689 1068 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.55 //y=7.4 //x2=57.72 //y2=7.4
r1620 (  689 692 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=57.55 //y=7.4 //x2=56.98 //y2=7.4
r1621 (  683 1067 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.64 //y=7.23 //x2=56.64 //y2=7.4
r1622 (  683 1152 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=56.64 //y=7.23 //x2=56.64 //y2=6.745
r1623 (  680 1066 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.845 //y=7.4 //x2=55.76 //y2=7.4
r1624 (  680 682 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=55.845 //y=7.4 //x2=55.87 //y2=7.4
r1625 (  679 1067 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.555 //y=7.4 //x2=56.64 //y2=7.4
r1626 (  679 682 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=56.555 //y=7.4 //x2=55.87 //y2=7.4
r1627 (  673 1066 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=55.76 //y=7.23 //x2=55.76 //y2=7.4
r1628 (  673 1151 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.76 //y=7.23 //x2=55.76 //y2=6.745
r1629 (  672 1065 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.965 //y=7.4 //x2=54.88 //y2=7.4
r1630 (  671 1066 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.675 //y=7.4 //x2=55.76 //y2=7.4
r1631 (  671 672 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=55.675 //y=7.4 //x2=54.965 //y2=7.4
r1632 (  665 1065 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=54.88 //y=7.23 //x2=54.88 //y2=7.4
r1633 (  665 1150 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.88 //y=7.23 //x2=54.88 //y2=6.745
r1634 (  662 1064 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.085 //y=7.4 //x2=54 //y2=7.4
r1635 (  662 664 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=54.085 //y=7.4 //x2=54.76 //y2=7.4
r1636 (  661 1065 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.795 //y=7.4 //x2=54.88 //y2=7.4
r1637 (  661 664 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=54.795 //y=7.4 //x2=54.76 //y2=7.4
r1638 (  655 1064 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=54 //y=7.23 //x2=54 //y2=7.4
r1639 (  655 1149 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=54 //y=7.23 //x2=54 //y2=6.405
r1640 (  652 1063 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.08 //y=7.4 //x2=52.91 //y2=7.4
r1641 (  652 654 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=53.08 //y=7.4 //x2=53.65 //y2=7.4
r1642 (  651 1064 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.915 //y=7.4 //x2=54 //y2=7.4
r1643 (  651 654 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=53.915 //y=7.4 //x2=53.65 //y2=7.4
r1644 (  646 1062 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.915 //y=7.4 //x2=51.83 //y2=7.4
r1645 (  646 648 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=51.915 //y=7.4 //x2=52.17 //y2=7.4
r1646 (  645 1063 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.74 //y=7.4 //x2=52.91 //y2=7.4
r1647 (  645 648 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=52.74 //y=7.4 //x2=52.17 //y2=7.4
r1648 (  639 1062 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.83 //y=7.23 //x2=51.83 //y2=7.4
r1649 (  639 1148 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=51.83 //y=7.23 //x2=51.83 //y2=6.745
r1650 (  636 1061 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.035 //y=7.4 //x2=50.95 //y2=7.4
r1651 (  636 638 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=51.035 //y=7.4 //x2=51.06 //y2=7.4
r1652 (  635 1062 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.745 //y=7.4 //x2=51.83 //y2=7.4
r1653 (  635 638 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=51.745 //y=7.4 //x2=51.06 //y2=7.4
r1654 (  629 1061 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.95 //y=7.23 //x2=50.95 //y2=7.4
r1655 (  629 1147 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.95 //y=7.23 //x2=50.95 //y2=6.745
r1656 (  628 1060 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.155 //y=7.4 //x2=50.07 //y2=7.4
r1657 (  627 1061 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.865 //y=7.4 //x2=50.95 //y2=7.4
r1658 (  627 628 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.865 //y=7.4 //x2=50.155 //y2=7.4
r1659 (  621 1060 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.07 //y=7.23 //x2=50.07 //y2=7.4
r1660 (  621 1146 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.07 //y=7.23 //x2=50.07 //y2=6.745
r1661 (  618 1059 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.275 //y=7.4 //x2=49.19 //y2=7.4
r1662 (  618 620 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=49.275 //y=7.4 //x2=49.95 //y2=7.4
r1663 (  617 1060 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.985 //y=7.4 //x2=50.07 //y2=7.4
r1664 (  617 620 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=49.985 //y=7.4 //x2=49.95 //y2=7.4
r1665 (  611 1059 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.19 //y=7.23 //x2=49.19 //y2=7.4
r1666 (  611 1145 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=49.19 //y=7.23 //x2=49.19 //y2=6.405
r1667 (  608 1058 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.27 //y=7.4 //x2=48.1 //y2=7.4
r1668 (  608 610 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.27 //y=7.4 //x2=48.84 //y2=7.4
r1669 (  607 1059 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.105 //y=7.4 //x2=49.19 //y2=7.4
r1670 (  607 610 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=49.105 //y=7.4 //x2=48.84 //y2=7.4
r1671 (  602 1057 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.105 //y=7.4 //x2=47.02 //y2=7.4
r1672 (  602 604 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=47.105 //y=7.4 //x2=47.36 //y2=7.4
r1673 (  601 1058 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.93 //y=7.4 //x2=48.1 //y2=7.4
r1674 (  601 604 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=47.93 //y=7.4 //x2=47.36 //y2=7.4
r1675 (  595 1057 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.02 //y=7.23 //x2=47.02 //y2=7.4
r1676 (  595 1144 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=47.02 //y=7.23 //x2=47.02 //y2=6.745
r1677 (  592 1056 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.225 //y=7.4 //x2=46.14 //y2=7.4
r1678 (  592 594 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=46.225 //y=7.4 //x2=46.25 //y2=7.4
r1679 (  591 1057 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.935 //y=7.4 //x2=47.02 //y2=7.4
r1680 (  591 594 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=46.935 //y=7.4 //x2=46.25 //y2=7.4
r1681 (  585 1056 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=46.14 //y=7.23 //x2=46.14 //y2=7.4
r1682 (  585 1143 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.14 //y=7.23 //x2=46.14 //y2=6.745
r1683 (  584 1055 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.345 //y=7.4 //x2=45.26 //y2=7.4
r1684 (  583 1056 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.055 //y=7.4 //x2=46.14 //y2=7.4
r1685 (  583 584 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.055 //y=7.4 //x2=45.345 //y2=7.4
r1686 (  577 1055 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=45.26 //y=7.23 //x2=45.26 //y2=7.4
r1687 (  577 1142 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.26 //y=7.23 //x2=45.26 //y2=6.745
r1688 (  574 1054 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.465 //y=7.4 //x2=44.38 //y2=7.4
r1689 (  574 576 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=44.465 //y=7.4 //x2=45.14 //y2=7.4
r1690 (  573 1055 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.175 //y=7.4 //x2=45.26 //y2=7.4
r1691 (  573 576 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=45.175 //y=7.4 //x2=45.14 //y2=7.4
r1692 (  567 1054 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.38 //y=7.23 //x2=44.38 //y2=7.4
r1693 (  567 1141 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=44.38 //y=7.23 //x2=44.38 //y2=6.405
r1694 (  564 1053 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.46 //y=7.4 //x2=43.29 //y2=7.4
r1695 (  564 566 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.46 //y=7.4 //x2=44.03 //y2=7.4
r1696 (  563 1054 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.295 //y=7.4 //x2=44.38 //y2=7.4
r1697 (  563 566 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=44.295 //y=7.4 //x2=44.03 //y2=7.4
r1698 (  558 1052 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.295 //y=7.4 //x2=42.21 //y2=7.4
r1699 (  558 560 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=42.295 //y=7.4 //x2=42.55 //y2=7.4
r1700 (  557 1053 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.12 //y=7.4 //x2=43.29 //y2=7.4
r1701 (  557 560 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.12 //y=7.4 //x2=42.55 //y2=7.4
r1702 (  551 1052 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=42.21 //y=7.23 //x2=42.21 //y2=7.4
r1703 (  551 1140 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=42.21 //y=7.23 //x2=42.21 //y2=6.745
r1704 (  548 1051 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.415 //y=7.4 //x2=41.33 //y2=7.4
r1705 (  548 550 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=41.415 //y=7.4 //x2=41.44 //y2=7.4
r1706 (  547 1052 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.125 //y=7.4 //x2=42.21 //y2=7.4
r1707 (  547 550 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=42.125 //y=7.4 //x2=41.44 //y2=7.4
r1708 (  541 1051 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=41.33 //y=7.23 //x2=41.33 //y2=7.4
r1709 (  541 1139 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=41.33 //y=7.23 //x2=41.33 //y2=6.745
r1710 (  540 1050 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.535 //y=7.4 //x2=40.45 //y2=7.4
r1711 (  539 1051 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.245 //y=7.4 //x2=41.33 //y2=7.4
r1712 (  539 540 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=41.245 //y=7.4 //x2=40.535 //y2=7.4
r1713 (  533 1050 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.45 //y=7.23 //x2=40.45 //y2=7.4
r1714 (  533 1138 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=40.45 //y=7.23 //x2=40.45 //y2=6.745
r1715 (  530 1049 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.655 //y=7.4 //x2=39.57 //y2=7.4
r1716 (  530 532 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=39.655 //y=7.4 //x2=40.33 //y2=7.4
r1717 (  529 1050 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.365 //y=7.4 //x2=40.45 //y2=7.4
r1718 (  529 532 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=40.365 //y=7.4 //x2=40.33 //y2=7.4
r1719 (  523 1049 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.57 //y=7.23 //x2=39.57 //y2=7.4
r1720 (  523 1137 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=39.57 //y=7.23 //x2=39.57 //y2=6.405
r1721 (  520 1048 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.65 //y=7.4 //x2=38.48 //y2=7.4
r1722 (  520 522 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.65 //y=7.4 //x2=39.22 //y2=7.4
r1723 (  519 1049 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.485 //y=7.4 //x2=39.57 //y2=7.4
r1724 (  519 522 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=39.485 //y=7.4 //x2=39.22 //y2=7.4
r1725 (  514 1047 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.485 //y=7.4 //x2=37.4 //y2=7.4
r1726 (  514 516 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=37.485 //y=7.4 //x2=37.74 //y2=7.4
r1727 (  513 1048 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.31 //y=7.4 //x2=38.48 //y2=7.4
r1728 (  513 516 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.31 //y=7.4 //x2=37.74 //y2=7.4
r1729 (  507 1047 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.4 //y=7.23 //x2=37.4 //y2=7.4
r1730 (  507 1136 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=37.4 //y=7.23 //x2=37.4 //y2=6.745
r1731 (  504 1046 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.605 //y=7.4 //x2=36.52 //y2=7.4
r1732 (  504 506 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=36.605 //y=7.4 //x2=36.63 //y2=7.4
r1733 (  503 1047 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.315 //y=7.4 //x2=37.4 //y2=7.4
r1734 (  503 506 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=37.315 //y=7.4 //x2=36.63 //y2=7.4
r1735 (  497 1046 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.52 //y=7.23 //x2=36.52 //y2=7.4
r1736 (  497 1135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=36.52 //y=7.23 //x2=36.52 //y2=6.745
r1737 (  496 1045 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.725 //y=7.4 //x2=35.64 //y2=7.4
r1738 (  495 1046 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.435 //y=7.4 //x2=36.52 //y2=7.4
r1739 (  495 496 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=36.435 //y=7.4 //x2=35.725 //y2=7.4
r1740 (  489 1045 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.64 //y=7.23 //x2=35.64 //y2=7.4
r1741 (  489 1134 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.64 //y=7.23 //x2=35.64 //y2=6.745
r1742 (  486 1044 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.845 //y=7.4 //x2=34.76 //y2=7.4
r1743 (  486 488 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=34.845 //y=7.4 //x2=35.52 //y2=7.4
r1744 (  485 1045 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.555 //y=7.4 //x2=35.64 //y2=7.4
r1745 (  485 488 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=35.555 //y=7.4 //x2=35.52 //y2=7.4
r1746 (  479 1044 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.76 //y=7.23 //x2=34.76 //y2=7.4
r1747 (  479 1133 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=34.76 //y=7.23 //x2=34.76 //y2=6.405
r1748 (  476 1043 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.84 //y=7.4 //x2=33.67 //y2=7.4
r1749 (  476 478 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=33.84 //y=7.4 //x2=34.41 //y2=7.4
r1750 (  475 1044 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.675 //y=7.4 //x2=34.76 //y2=7.4
r1751 (  475 478 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=34.675 //y=7.4 //x2=34.41 //y2=7.4
r1752 (  470 1042 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.675 //y=7.4 //x2=32.59 //y2=7.4
r1753 (  470 472 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=32.675 //y=7.4 //x2=32.93 //y2=7.4
r1754 (  469 1043 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.5 //y=7.4 //x2=33.67 //y2=7.4
r1755 (  469 472 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=33.5 //y=7.4 //x2=32.93 //y2=7.4
r1756 (  463 1042 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.59 //y=7.23 //x2=32.59 //y2=7.4
r1757 (  463 1132 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=32.59 //y=7.23 //x2=32.59 //y2=6.745
r1758 (  460 1041 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.795 //y=7.4 //x2=31.71 //y2=7.4
r1759 (  460 462 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=31.795 //y=7.4 //x2=31.82 //y2=7.4
r1760 (  459 1042 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.505 //y=7.4 //x2=32.59 //y2=7.4
r1761 (  459 462 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=32.505 //y=7.4 //x2=31.82 //y2=7.4
r1762 (  453 1041 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.71 //y=7.23 //x2=31.71 //y2=7.4
r1763 (  453 1131 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.71 //y=7.23 //x2=31.71 //y2=6.745
r1764 (  452 1040 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.915 //y=7.4 //x2=30.83 //y2=7.4
r1765 (  451 1041 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.625 //y=7.4 //x2=31.71 //y2=7.4
r1766 (  451 452 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=31.625 //y=7.4 //x2=30.915 //y2=7.4
r1767 (  445 1040 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.83 //y=7.23 //x2=30.83 //y2=7.4
r1768 (  445 1130 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=30.83 //y=7.23 //x2=30.83 //y2=6.745
r1769 (  442 1039 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.035 //y=7.4 //x2=29.95 //y2=7.4
r1770 (  442 444 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=30.035 //y=7.4 //x2=30.71 //y2=7.4
r1771 (  441 1040 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.745 //y=7.4 //x2=30.83 //y2=7.4
r1772 (  441 444 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=30.745 //y=7.4 //x2=30.71 //y2=7.4
r1773 (  435 1039 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.95 //y=7.23 //x2=29.95 //y2=7.4
r1774 (  435 1129 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=29.95 //y=7.23 //x2=29.95 //y2=6.405
r1775 (  432 1038 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.03 //y=7.4 //x2=28.86 //y2=7.4
r1776 (  432 434 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=29.03 //y=7.4 //x2=29.6 //y2=7.4
r1777 (  431 1039 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.865 //y=7.4 //x2=29.95 //y2=7.4
r1778 (  431 434 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=29.865 //y=7.4 //x2=29.6 //y2=7.4
r1779 (  426 1037 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.865 //y=7.4 //x2=27.78 //y2=7.4
r1780 (  426 428 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=27.865 //y=7.4 //x2=28.12 //y2=7.4
r1781 (  425 1038 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.69 //y=7.4 //x2=28.86 //y2=7.4
r1782 (  425 428 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=28.69 //y=7.4 //x2=28.12 //y2=7.4
r1783 (  419 1037 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.78 //y=7.23 //x2=27.78 //y2=7.4
r1784 (  419 1128 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.78 //y=7.23 //x2=27.78 //y2=6.745
r1785 (  416 1036 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.985 //y=7.4 //x2=26.9 //y2=7.4
r1786 (  416 418 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=26.985 //y=7.4 //x2=27.01 //y2=7.4
r1787 (  415 1037 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.695 //y=7.4 //x2=27.78 //y2=7.4
r1788 (  415 418 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=27.695 //y=7.4 //x2=27.01 //y2=7.4
r1789 (  409 1036 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.9 //y=7.23 //x2=26.9 //y2=7.4
r1790 (  409 1127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.9 //y=7.23 //x2=26.9 //y2=6.745
r1791 (  408 1035 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.105 //y=7.4 //x2=26.02 //y2=7.4
r1792 (  407 1036 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.815 //y=7.4 //x2=26.9 //y2=7.4
r1793 (  407 408 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.815 //y=7.4 //x2=26.105 //y2=7.4
r1794 (  401 1035 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.02 //y=7.23 //x2=26.02 //y2=7.4
r1795 (  401 1126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.02 //y=7.23 //x2=26.02 //y2=6.745
r1796 (  398 1034 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.225 //y=7.4 //x2=25.14 //y2=7.4
r1797 (  398 400 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=25.225 //y=7.4 //x2=25.9 //y2=7.4
r1798 (  397 1035 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.935 //y=7.4 //x2=26.02 //y2=7.4
r1799 (  397 400 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=25.935 //y=7.4 //x2=25.9 //y2=7.4
r1800 (  391 1034 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.14 //y=7.23 //x2=25.14 //y2=7.4
r1801 (  391 1125 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=25.14 //y=7.23 //x2=25.14 //y2=6.405
r1802 (  388 1033 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.22 //y=7.4 //x2=24.05 //y2=7.4
r1803 (  388 390 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.22 //y=7.4 //x2=24.79 //y2=7.4
r1804 (  387 1034 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.055 //y=7.4 //x2=25.14 //y2=7.4
r1805 (  387 390 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=25.055 //y=7.4 //x2=24.79 //y2=7.4
r1806 (  382 1032 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.055 //y=7.4 //x2=22.97 //y2=7.4
r1807 (  382 384 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=23.055 //y=7.4 //x2=23.31 //y2=7.4
r1808 (  381 1033 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.88 //y=7.4 //x2=24.05 //y2=7.4
r1809 (  381 384 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.88 //y=7.4 //x2=23.31 //y2=7.4
r1810 (  375 1032 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.97 //y=7.23 //x2=22.97 //y2=7.4
r1811 (  375 1124 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.97 //y=7.23 //x2=22.97 //y2=6.745
r1812 (  372 1031 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.175 //y=7.4 //x2=22.09 //y2=7.4
r1813 (  372 374 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=22.175 //y=7.4 //x2=22.2 //y2=7.4
r1814 (  371 1032 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.885 //y=7.4 //x2=22.97 //y2=7.4
r1815 (  371 374 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=22.885 //y=7.4 //x2=22.2 //y2=7.4
r1816 (  365 1031 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.09 //y=7.23 //x2=22.09 //y2=7.4
r1817 (  365 1123 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.09 //y=7.23 //x2=22.09 //y2=6.745
r1818 (  364 1030 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.295 //y=7.4 //x2=21.21 //y2=7.4
r1819 (  363 1031 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.005 //y=7.4 //x2=22.09 //y2=7.4
r1820 (  363 364 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.005 //y=7.4 //x2=21.295 //y2=7.4
r1821 (  357 1030 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.21 //y=7.23 //x2=21.21 //y2=7.4
r1822 (  357 1122 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.21 //y=7.23 //x2=21.21 //y2=6.745
r1823 (  354 1029 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.415 //y=7.4 //x2=20.33 //y2=7.4
r1824 (  354 356 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=20.415 //y=7.4 //x2=21.09 //y2=7.4
r1825 (  353 1030 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.125 //y=7.4 //x2=21.21 //y2=7.4
r1826 (  353 356 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=21.125 //y=7.4 //x2=21.09 //y2=7.4
r1827 (  347 1029 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.33 //y=7.23 //x2=20.33 //y2=7.4
r1828 (  347 1121 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=20.33 //y=7.23 //x2=20.33 //y2=6.405
r1829 (  344 1028 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.41 //y=7.4 //x2=19.24 //y2=7.4
r1830 (  344 346 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.41 //y=7.4 //x2=19.98 //y2=7.4
r1831 (  343 1029 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.245 //y=7.4 //x2=20.33 //y2=7.4
r1832 (  343 346 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.245 //y=7.4 //x2=19.98 //y2=7.4
r1833 (  338 1027 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.245 //y=7.4 //x2=18.16 //y2=7.4
r1834 (  338 340 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=18.245 //y=7.4 //x2=18.5 //y2=7.4
r1835 (  337 1028 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.07 //y=7.4 //x2=19.24 //y2=7.4
r1836 (  337 340 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.07 //y=7.4 //x2=18.5 //y2=7.4
r1837 (  331 1027 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.16 //y=7.23 //x2=18.16 //y2=7.4
r1838 (  331 1120 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=18.16 //y=7.23 //x2=18.16 //y2=6.745
r1839 (  328 1026 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.365 //y=7.4 //x2=17.28 //y2=7.4
r1840 (  328 330 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=17.365 //y=7.4 //x2=17.39 //y2=7.4
r1841 (  327 1027 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.075 //y=7.4 //x2=18.16 //y2=7.4
r1842 (  327 330 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=18.075 //y=7.4 //x2=17.39 //y2=7.4
r1843 (  321 1026 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.28 //y=7.23 //x2=17.28 //y2=7.4
r1844 (  321 1119 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.28 //y=7.23 //x2=17.28 //y2=6.745
r1845 (  320 1025 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.485 //y=7.4 //x2=16.4 //y2=7.4
r1846 (  319 1026 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.195 //y=7.4 //x2=17.28 //y2=7.4
r1847 (  319 320 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=17.195 //y=7.4 //x2=16.485 //y2=7.4
r1848 (  313 1025 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.4 //y=7.23 //x2=16.4 //y2=7.4
r1849 (  313 1118 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.4 //y=7.23 //x2=16.4 //y2=6.745
r1850 (  310 1024 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.605 //y=7.4 //x2=15.52 //y2=7.4
r1851 (  310 312 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=15.605 //y=7.4 //x2=16.28 //y2=7.4
r1852 (  309 1025 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.315 //y=7.4 //x2=16.4 //y2=7.4
r1853 (  309 312 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=16.315 //y=7.4 //x2=16.28 //y2=7.4
r1854 (  303 1024 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.52 //y=7.23 //x2=15.52 //y2=7.4
r1855 (  303 1117 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=15.52 //y=7.23 //x2=15.52 //y2=6.405
r1856 (  300 1023 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=14.43 //y2=7.4
r1857 (  300 302 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=15.17 //y2=7.4
r1858 (  299 1024 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.435 //y=7.4 //x2=15.52 //y2=7.4
r1859 (  299 302 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.435 //y=7.4 //x2=15.17 //y2=7.4
r1860 (  294 1022 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.435 //y=7.4 //x2=13.35 //y2=7.4
r1861 (  294 296 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=13.435 //y=7.4 //x2=13.69 //y2=7.4
r1862 (  293 1023 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=14.43 //y2=7.4
r1863 (  293 296 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=13.69 //y2=7.4
r1864 (  287 1022 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.35 //y=7.23 //x2=13.35 //y2=7.4
r1865 (  287 1116 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=13.35 //y=7.23 //x2=13.35 //y2=6.745
r1866 (  284 1021 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.555 //y=7.4 //x2=12.47 //y2=7.4
r1867 (  284 286 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=12.555 //y=7.4 //x2=12.58 //y2=7.4
r1868 (  283 1022 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.265 //y=7.4 //x2=13.35 //y2=7.4
r1869 (  283 286 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=13.265 //y=7.4 //x2=12.58 //y2=7.4
r1870 (  277 1021 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.47 //y=7.23 //x2=12.47 //y2=7.4
r1871 (  277 1115 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.47 //y=7.23 //x2=12.47 //y2=6.745
r1872 (  276 1020 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.675 //y=7.4 //x2=11.59 //y2=7.4
r1873 (  275 1021 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.385 //y=7.4 //x2=12.47 //y2=7.4
r1874 (  275 276 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=12.385 //y=7.4 //x2=11.675 //y2=7.4
r1875 (  269 1020 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.59 //y=7.23 //x2=11.59 //y2=7.4
r1876 (  269 1114 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.59 //y=7.23 //x2=11.59 //y2=6.745
r1877 (  266 1019 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.795 //y=7.4 //x2=10.71 //y2=7.4
r1878 (  266 268 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=10.795 //y=7.4 //x2=11.47 //y2=7.4
r1879 (  265 1020 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.505 //y=7.4 //x2=11.59 //y2=7.4
r1880 (  265 268 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=11.505 //y=7.4 //x2=11.47 //y2=7.4
r1881 (  259 1019 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.71 //y=7.23 //x2=10.71 //y2=7.4
r1882 (  259 1113 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.71 //y=7.23 //x2=10.71 //y2=6.405
r1883 (  256 1018 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=9.62 //y2=7.4
r1884 (  256 258 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=10.36 //y2=7.4
r1885 (  255 1019 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.625 //y=7.4 //x2=10.71 //y2=7.4
r1886 (  255 258 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=10.625 //y=7.4 //x2=10.36 //y2=7.4
r1887 (  250 1017 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.54 //y2=7.4
r1888 (  250 252 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.88 //y2=7.4
r1889 (  249 1018 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=9.62 //y2=7.4
r1890 (  249 252 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=8.88 //y2=7.4
r1891 (  243 1017 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=7.4
r1892 (  243 1112 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=6.745
r1893 (  240 1016 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.66 //y2=7.4
r1894 (  240 242 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.77 //y2=7.4
r1895 (  239 1017 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=8.54 //y2=7.4
r1896 (  239 242 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=7.77 //y2=7.4
r1897 (  233 1016 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=7.4
r1898 (  233 1111 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=6.745
r1899 (  232 1015 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=6.78 //y2=7.4
r1900 (  231 1016 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=7.66 //y2=7.4
r1901 (  231 232 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=6.865 //y2=7.4
r1902 (  225 1015 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=7.4
r1903 (  225 1110 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=6.745
r1904 (  222 1014 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=5.9 //y2=7.4
r1905 (  222 224 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=6.66 //y2=7.4
r1906 (  221 1015 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.78 //y2=7.4
r1907 (  221 224 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.66 //y2=7.4
r1908 (  215 1014 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=7.4
r1909 (  215 1109 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=6.405
r1910 (  212 1013 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r1911 (  212 214 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=5.55 //y2=7.4
r1912 (  211 1014 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.9 //y2=7.4
r1913 (  211 214 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.55 //y2=7.4
r1914 (  206 1012 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r1915 (  206 208 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r1916 (  205 1013 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r1917 (  205 208 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r1918 (  199 1012 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r1919 (  199 1108 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r1920 (  196 1011 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r1921 (  196 198 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r1922 (  195 1012 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r1923 (  195 198 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r1924 (  189 1011 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r1925 (  189 1107 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r1926 (  188 1010 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r1927 (  187 1011 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r1928 (  187 188 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r1929 (  181 1010 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r1930 (  181 1106 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r1931 (  178 1009 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r1932 (  178 180 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r1933 (  177 1010 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r1934 (  177 180 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r1935 (  171 1009 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r1936 (  171 1105 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r1937 (  167 1009 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r1938 (  167 170 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r1939 (  163 1006 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=95.83 //y=7.4 //x2=95.83 //y2=7.4
r1940 (  161 1004 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=94.72 //y=7.4 //x2=94.72 //y2=7.4
r1941 (  161 163 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=94.72 //y=7.4 //x2=95.83 //y2=7.4
r1942 (  159 1002 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=93.61 //y=7.4 //x2=93.61 //y2=7.4
r1943 (  159 161 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=93.61 //y=7.4 //x2=94.72 //y2=7.4
r1944 (  157 996 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=92.13 //y=7.4 //x2=92.13 //y2=7.4
r1945 (  157 159 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=92.13 //y=7.4 //x2=93.61 //y2=7.4
r1946 (  155 994 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=91.02 //y=7.4 //x2=91.02 //y2=7.4
r1947 (  155 157 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=91.02 //y=7.4 //x2=92.13 //y2=7.4
r1948 (  153 988 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=89.54 //y=7.4 //x2=89.54 //y2=7.4
r1949 (  153 155 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=89.54 //y=7.4 //x2=91.02 //y2=7.4
r1950 (  151 978 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=88.43 //y=7.4 //x2=88.43 //y2=7.4
r1951 (  151 153 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=88.43 //y=7.4 //x2=89.54 //y2=7.4
r1952 (  149 1100 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=87.32 //y=7.4 //x2=87.32 //y2=7.4
r1953 (  149 151 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=87.32 //y=7.4 //x2=88.43 //y2=7.4
r1954 (  147 956 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=85.84 //y=7.4 //x2=85.84 //y2=7.4
r1955 (  147 149 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=85.84 //y=7.4 //x2=87.32 //y2=7.4
r1956 (  145 946 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=84.73 //y=7.4 //x2=84.73 //y2=7.4
r1957 (  145 147 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=84.73 //y=7.4 //x2=85.84 //y2=7.4
r1958 (  143 928 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=83.62 //y=7.4 //x2=83.62 //y2=7.4
r1959 (  143 145 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=83.62 //y=7.4 //x2=84.73 //y2=7.4
r1960 (  141 918 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.51 //y=7.4 //x2=82.51 //y2=7.4
r1961 (  141 143 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=82.51 //y=7.4 //x2=83.62 //y2=7.4
r1962 (  139 912 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=81.03 //y=7.4 //x2=81.03 //y2=7.4
r1963 (  139 141 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=81.03 //y=7.4 //x2=82.51 //y2=7.4
r1964 (  137 902 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=79.92 //y=7.4 //x2=79.92 //y2=7.4
r1965 (  137 139 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=79.92 //y=7.4 //x2=81.03 //y2=7.4
r1966 (  135 884 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.81 //y=7.4 //x2=78.81 //y2=7.4
r1967 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=78.81 //y=7.4 //x2=79.92 //y2=7.4
r1968 (  133 874 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=77.7 //y=7.4 //x2=77.7 //y2=7.4
r1969 (  133 135 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=77.7 //y=7.4 //x2=78.81 //y2=7.4
r1970 (  131 868 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.22 //y=7.4 //x2=76.22 //y2=7.4
r1971 (  131 133 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.22 //y=7.4 //x2=77.7 //y2=7.4
r1972 (  129 858 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.11 //y=7.4 //x2=75.11 //y2=7.4
r1973 (  129 131 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=7.4 //x2=76.22 //y2=7.4
r1974 (  127 840 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74 //y=7.4 //x2=74 //y2=7.4
r1975 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74 //y=7.4 //x2=75.11 //y2=7.4
r1976 (  125 830 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.89 //y=7.4 //x2=72.89 //y2=7.4
r1977 (  125 127 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=72.89 //y=7.4 //x2=74 //y2=7.4
r1978 (  123 824 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=7.4 //x2=71.41 //y2=7.4
r1979 (  123 125 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=7.4 //x2=72.89 //y2=7.4
r1980 (  121 814 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=70.3 //y=7.4 //x2=70.3 //y2=7.4
r1981 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=70.3 //y=7.4 //x2=71.41 //y2=7.4
r1982 (  119 796 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.19 //y=7.4 //x2=69.19 //y2=7.4
r1983 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.19 //y=7.4 //x2=70.3 //y2=7.4
r1984 (  117 786 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=68.08 //y=7.4 //x2=68.08 //y2=7.4
r1985 (  117 119 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=68.08 //y=7.4 //x2=69.19 //y2=7.4
r1986 (  115 780 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.6 //y=7.4 //x2=66.6 //y2=7.4
r1987 (  115 117 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=66.6 //y=7.4 //x2=68.08 //y2=7.4
r1988 (  113 770 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.49 //y=7.4 //x2=65.49 //y2=7.4
r1989 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.49 //y=7.4 //x2=66.6 //y2=7.4
r1990 (  111 752 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=64.38 //y=7.4 //x2=64.38 //y2=7.4
r1991 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=64.38 //y=7.4 //x2=65.49 //y2=7.4
r1992 (  109 742 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=63.27 //y=7.4 //x2=63.27 //y2=7.4
r1993 (  109 111 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=63.27 //y=7.4 //x2=64.38 //y2=7.4
r1994 (  107 736 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.79 //y=7.4 //x2=61.79 //y2=7.4
r1995 (  107 109 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.79 //y=7.4 //x2=63.27 //y2=7.4
r1996 (  105 726 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=60.68 //y=7.4 //x2=60.68 //y2=7.4
r1997 (  105 107 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=60.68 //y=7.4 //x2=61.79 //y2=7.4
r1998 (  103 708 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.57 //y=7.4 //x2=59.57 //y2=7.4
r1999 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.57 //y=7.4 //x2=60.68 //y2=7.4
r2000 (  101 698 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.46 //y=7.4 //x2=58.46 //y2=7.4
r2001 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.46 //y=7.4 //x2=59.57 //y2=7.4
r2002 (  99 692 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.98 //y=7.4 //x2=56.98 //y2=7.4
r2003 (  99 101 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.98 //y=7.4 //x2=58.46 //y2=7.4
r2004 (  97 682 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.87 //y=7.4 //x2=55.87 //y2=7.4
r2005 (  97 99 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.87 //y=7.4 //x2=56.98 //y2=7.4
r2006 (  95 664 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.76 //y=7.4 //x2=54.76 //y2=7.4
r2007 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.76 //y=7.4 //x2=55.87 //y2=7.4
r2008 (  93 654 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.65 //y=7.4 //x2=53.65 //y2=7.4
r2009 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=53.65 //y=7.4 //x2=54.76 //y2=7.4
r2010 (  91 648 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=52.17 //y=7.4 //x2=52.17 //y2=7.4
r2011 (  91 93 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=52.17 //y=7.4 //x2=53.65 //y2=7.4
r2012 (  89 638 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.06 //y=7.4 //x2=51.06 //y2=7.4
r2013 (  89 91 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=51.06 //y=7.4 //x2=52.17 //y2=7.4
r2014 (  87 620 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.95 //y=7.4 //x2=49.95 //y2=7.4
r2015 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.95 //y=7.4 //x2=51.06 //y2=7.4
r2016 (  85 610 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.84 //y=7.4 //x2=48.84 //y2=7.4
r2017 (  85 87 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=48.84 //y=7.4 //x2=49.95 //y2=7.4
r2018 (  82 604 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=47.36 //y=7.4 //x2=47.36 //y2=7.4
r2019 (  80 594 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.25 //y=7.4 //x2=46.25 //y2=7.4
r2020 (  80 82 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.25 //y=7.4 //x2=47.36 //y2=7.4
r2021 (  78 576 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.14 //y=7.4 //x2=45.14 //y2=7.4
r2022 (  78 80 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.14 //y=7.4 //x2=46.25 //y2=7.4
r2023 (  76 566 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.03 //y=7.4 //x2=44.03 //y2=7.4
r2024 (  76 78 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.03 //y=7.4 //x2=45.14 //y2=7.4
r2025 (  74 560 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.55 //y=7.4 //x2=42.55 //y2=7.4
r2026 (  74 76 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=42.55 //y=7.4 //x2=44.03 //y2=7.4
r2027 (  72 550 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.44 //y=7.4 //x2=41.44 //y2=7.4
r2028 (  72 74 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.44 //y=7.4 //x2=42.55 //y2=7.4
r2029 (  70 532 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=40.33 //y=7.4 //x2=40.33 //y2=7.4
r2030 (  70 72 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=40.33 //y=7.4 //x2=41.44 //y2=7.4
r2031 (  68 522 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.22 //y=7.4 //x2=39.22 //y2=7.4
r2032 (  68 70 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=39.22 //y=7.4 //x2=40.33 //y2=7.4
r2033 (  66 516 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37.74 //y=7.4 //x2=37.74 //y2=7.4
r2034 (  66 68 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=37.74 //y=7.4 //x2=39.22 //y2=7.4
r2035 (  64 506 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=36.63 //y=7.4 //x2=36.63 //y2=7.4
r2036 (  64 66 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=36.63 //y=7.4 //x2=37.74 //y2=7.4
r2037 (  62 488 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.52 //y=7.4 //x2=35.52 //y2=7.4
r2038 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.52 //y=7.4 //x2=36.63 //y2=7.4
r2039 (  60 478 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.41 //y=7.4 //x2=34.41 //y2=7.4
r2040 (  60 62 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.41 //y=7.4 //x2=35.52 //y2=7.4
r2041 (  58 472 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.93 //y=7.4 //x2=32.93 //y2=7.4
r2042 (  58 60 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.93 //y=7.4 //x2=34.41 //y2=7.4
r2043 (  56 462 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.82 //y=7.4 //x2=31.82 //y2=7.4
r2044 (  56 58 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.82 //y=7.4 //x2=32.93 //y2=7.4
r2045 (  54 444 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=30.71 //y=7.4 //x2=30.71 //y2=7.4
r2046 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=30.71 //y=7.4 //x2=31.82 //y2=7.4
r2047 (  52 434 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.6 //y=7.4 //x2=29.6 //y2=7.4
r2048 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=29.6 //y=7.4 //x2=30.71 //y2=7.4
r2049 (  50 428 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.12 //y=7.4 //x2=28.12 //y2=7.4
r2050 (  50 52 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=28.12 //y=7.4 //x2=29.6 //y2=7.4
r2051 (  48 418 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.01 //y=7.4 //x2=27.01 //y2=7.4
r2052 (  48 50 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.01 //y=7.4 //x2=28.12 //y2=7.4
r2053 (  46 400 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.9 //y=7.4 //x2=25.9 //y2=7.4
r2054 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.9 //y=7.4 //x2=27.01 //y2=7.4
r2055 (  44 390 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=7.4 //x2=24.79 //y2=7.4
r2056 (  44 46 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=7.4 //x2=25.9 //y2=7.4
r2057 (  42 384 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.31 //y=7.4 //x2=23.31 //y2=7.4
r2058 (  42 44 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.31 //y=7.4 //x2=24.79 //y2=7.4
r2059 (  40 374 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=7.4 //x2=22.2 //y2=7.4
r2060 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=7.4 //x2=23.31 //y2=7.4
r2061 (  38 356 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=7.4 //x2=21.09 //y2=7.4
r2062 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=7.4 //x2=22.2 //y2=7.4
r2063 (  36 346 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=7.4 //x2=19.98 //y2=7.4
r2064 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=7.4 //x2=21.09 //y2=7.4
r2065 (  34 340 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=7.4 //x2=18.5 //y2=7.4
r2066 (  34 36 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=7.4 //x2=19.98 //y2=7.4
r2067 (  32 330 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r2068 (  32 34 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.4 //x2=18.5 //y2=7.4
r2069 (  30 312 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=7.4 //x2=16.28 //y2=7.4
r2070 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=7.4 //x2=17.39 //y2=7.4
r2071 (  28 302 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r2072 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.28 //y2=7.4
r2073 (  26 296 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=7.4 //x2=13.69 //y2=7.4
r2074 (  26 28 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=7.4 //x2=15.17 //y2=7.4
r2075 (  24 286 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r2076 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.4 //x2=13.69 //y2=7.4
r2077 (  22 268 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r2078 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=7.4 //x2=12.58 //y2=7.4
r2079 (  20 258 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r2080 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r2081 (  18 252 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=7.4 //x2=8.88 //y2=7.4
r2082 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=7.4 //x2=10.36 //y2=7.4
r2083 (  16 242 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r2084 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=8.88 //y2=7.4
r2085 (  14 224 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r2086 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r2087 (  12 214 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r2088 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r2089 (  10 208 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r2090 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.4 //x2=5.55 //y2=7.4
r2091 (  8 198 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r2092 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r2093 (  6 180 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r2094 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r2095 (  3 170 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r2096 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r2097 (  1 85 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=48.285 //y=7.4 //x2=48.84 //y2=7.4
r2098 (  1 82 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=48.285 //y=7.4 //x2=47.36 //y2=7.4
ends PM_TMRDFFSNRNQNX1\%VDD

subckt PM_TMRDFFSNRNQNX1\%noxref_3 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 \
 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c240 ( 127 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c241 ( 126 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c242 ( 125 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c243 ( 123 0 ) capacitor c=0.00853354f //x=3.395 //y=0.915
c244 ( 103 0 ) capacitor c=0.0556143f //x=11.005 //y=4.79
c245 ( 102 0 ) capacitor c=0.0293157f //x=11.295 //y=4.79
c246 ( 101 0 ) capacitor c=0.0347816f //x=10.96 //y=1.22
c247 ( 100 0 ) capacitor c=0.0187487f //x=10.96 //y=0.875
c248 ( 94 0 ) capacitor c=0.0137055f //x=10.805 //y=1.375
c249 ( 92 0 ) capacitor c=0.0149861f //x=10.805 //y=0.72
c250 ( 91 0 ) capacitor c=0.096037f //x=10.43 //y=1.915
c251 ( 90 0 ) capacitor c=0.0228993f //x=10.43 //y=1.53
c252 ( 89 0 ) capacitor c=0.0234352f //x=10.43 //y=1.22
c253 ( 88 0 ) capacitor c=0.0198724f //x=10.43 //y=0.875
c254 ( 84 0 ) capacitor c=0.055995f //x=6.195 //y=4.79
c255 ( 83 0 ) capacitor c=0.0298189f //x=6.485 //y=4.79
c256 ( 82 0 ) capacitor c=0.0347816f //x=6.15 //y=1.22
c257 ( 81 0 ) capacitor c=0.0187487f //x=6.15 //y=0.875
c258 ( 75 0 ) capacitor c=0.0137055f //x=5.995 //y=1.375
c259 ( 73 0 ) capacitor c=0.0149861f //x=5.995 //y=0.72
c260 ( 72 0 ) capacitor c=0.096037f //x=5.62 //y=1.915
c261 ( 71 0 ) capacitor c=0.0228993f //x=5.62 //y=1.53
c262 ( 70 0 ) capacitor c=0.0234352f //x=5.62 //y=1.22
c263 ( 69 0 ) capacitor c=0.0198724f //x=5.62 //y=0.875
c264 ( 68 0 ) capacitor c=0.110114f //x=11.37 //y=6.02
c265 ( 67 0 ) capacitor c=0.158956f //x=10.93 //y=6.02
c266 ( 66 0 ) capacitor c=0.110114f //x=6.56 //y=6.02
c267 ( 65 0 ) capacitor c=0.158956f //x=6.12 //y=6.02
c268 ( 62 0 ) capacitor c=0.00116729f //x=3.29 //y=5.155
c269 ( 61 0 ) capacitor c=0.00226015f //x=2.41 //y=5.155
c270 ( 54 0 ) capacitor c=0.0970684f //x=10.73 //y=2.08
c271 ( 46 0 ) capacitor c=0.102314f //x=5.92 //y=2.08
c272 ( 44 0 ) capacitor c=0.111586f //x=4.07 //y=2.59
c273 ( 40 0 ) capacitor c=0.00398962f //x=3.67 //y=1.665
c274 ( 39 0 ) capacitor c=0.0137288f //x=3.985 //y=1.665
c275 ( 33 0 ) capacitor c=0.0291119f //x=3.985 //y=5.155
c276 ( 25 0 ) capacitor c=0.0184197f //x=3.205 //y=5.155
c277 ( 18 0 ) capacitor c=0.00351598f //x=1.615 //y=5.155
c278 ( 17 0 ) capacitor c=0.0155255f //x=2.325 //y=5.155
c279 ( 4 0 ) capacitor c=0.00440131f //x=6.035 //y=2.59
c280 ( 3 0 ) capacitor c=0.0870935f //x=10.615 //y=2.59
c281 ( 2 0 ) capacitor c=0.0124623f //x=4.185 //y=2.59
c282 ( 1 0 ) capacitor c=0.0300768f //x=5.805 //y=2.59
r283 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.295 //y=4.79 //x2=11.37 //y2=4.865
r284 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=11.295 //y=4.79 //x2=11.005 //y2=4.79
r285 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.96 //y=1.22 //x2=10.92 //y2=1.375
r286 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.96 //y=0.875 //x2=10.92 //y2=0.72
r287 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.96 //y=0.875 //x2=10.96 //y2=1.22
r288 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.93 //y=4.865 //x2=11.005 //y2=4.79
r289 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=10.93 //y=4.865 //x2=10.73 //y2=4.7
r290 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.585 //y=1.375 //x2=10.47 //y2=1.375
r291 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.805 //y=1.375 //x2=10.92 //y2=1.375
r292 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.585 //y=0.72 //x2=10.47 //y2=0.72
r293 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.805 //y=0.72 //x2=10.92 //y2=0.72
r294 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.805 //y=0.72 //x2=10.585 //y2=0.72
r295 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.915 //x2=10.73 //y2=2.08
r296 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.53 //x2=10.47 //y2=1.375
r297 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.53 //x2=10.43 //y2=1.915
r298 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.22 //x2=10.47 //y2=1.375
r299 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=0.875 //x2=10.47 //y2=0.72
r300 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.43 //y=0.875 //x2=10.43 //y2=1.22
r301 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.56 //y2=4.865
r302 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.195 //y2=4.79
r303 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=1.22 //x2=6.11 //y2=1.375
r304 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.11 //y2=0.72
r305 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.15 //y2=1.22
r306 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=6.195 //y2=4.79
r307 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=5.92 //y2=4.7
r308 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=1.375 //x2=5.66 //y2=1.375
r309 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=1.375 //x2=6.11 //y2=1.375
r310 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=0.72 //x2=5.66 //y2=0.72
r311 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=6.11 //y2=0.72
r312 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=5.775 //y2=0.72
r313 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.915 //x2=5.92 //y2=2.08
r314 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.66 //y2=1.375
r315 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.62 //y2=1.915
r316 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.22 //x2=5.66 //y2=1.375
r317 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.66 //y2=0.72
r318 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.62 //y2=1.22
r319 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.37 //y=6.02 //x2=11.37 //y2=4.865
r320 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.93 //y=6.02 //x2=10.93 //y2=4.865
r321 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.56 //y=6.02 //x2=6.56 //y2=4.865
r322 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.12 //y=6.02 //x2=6.12 //y2=4.865
r323 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.695 //y=1.375 //x2=10.805 //y2=1.375
r324 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.695 //y=1.375 //x2=10.585 //y2=1.375
r325 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.995 //y2=1.375
r326 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.775 //y2=1.375
r327 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=4.7 //x2=10.73 //y2=4.7
r328 (  57 59 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.59 //x2=10.73 //y2=4.7
r329 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=2.08 //x2=10.73 //y2=2.08
r330 (  54 57 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.08 //x2=10.73 //y2=2.59
r331 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.7 //x2=5.92 //y2=4.7
r332 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.59 //x2=5.92 //y2=4.7
r333 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r334 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=2.59
r335 (  42 44 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=2.59
r336 (  41 44 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=2.59
r337 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r338 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r339 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r340 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r341 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r342 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r343 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r344 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r345 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r346 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r347 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r348 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r349 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r350 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r351 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r352 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r353 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r354 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r355 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=2.59 //x2=10.73 //y2=2.59
r356 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=2.59 //x2=5.92 //y2=2.59
r357 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=2.59 //x2=4.07 //y2=2.59
r358 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=2.59 //x2=5.92 //y2=2.59
r359 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.59 //x2=10.73 //y2=2.59
r360 (  3 4 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.59 //x2=6.035 //y2=2.59
r361 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=2.59 //x2=4.07 //y2=2.59
r362 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.805 //y=2.59 //x2=5.92 //y2=2.59
r363 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.805 //y=2.59 //x2=4.185 //y2=2.59
ends PM_TMRDFFSNRNQNX1\%noxref_3

subckt PM_TMRDFFSNRNQNX1\%noxref_4 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 \
 53 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c165 ( 85 0 ) capacitor c=0.023087f //x=12.765 //y=5.02
c166 ( 84 0 ) capacitor c=0.023519f //x=11.885 //y=5.02
c167 ( 83 0 ) capacitor c=0.0224735f //x=11.005 //y=5.02
c168 ( 81 0 ) capacitor c=0.00853354f //x=13.015 //y=0.915
c169 ( 69 0 ) capacitor c=0.0557698f //x=15.815 //y=4.79
c170 ( 68 0 ) capacitor c=0.0293157f //x=16.105 //y=4.79
c171 ( 67 0 ) capacitor c=0.0347816f //x=15.77 //y=1.22
c172 ( 66 0 ) capacitor c=0.0187487f //x=15.77 //y=0.875
c173 ( 60 0 ) capacitor c=0.0137055f //x=15.615 //y=1.375
c174 ( 58 0 ) capacitor c=0.0149861f //x=15.615 //y=0.72
c175 ( 57 0 ) capacitor c=0.096037f //x=15.24 //y=1.915
c176 ( 56 0 ) capacitor c=0.0228993f //x=15.24 //y=1.53
c177 ( 55 0 ) capacitor c=0.0234352f //x=15.24 //y=1.22
c178 ( 54 0 ) capacitor c=0.0198724f //x=15.24 //y=0.875
c179 ( 53 0 ) capacitor c=0.110114f //x=16.18 //y=6.02
c180 ( 52 0 ) capacitor c=0.158956f //x=15.74 //y=6.02
c181 ( 50 0 ) capacitor c=0.00106608f //x=12.91 //y=5.155
c182 ( 49 0 ) capacitor c=0.00207319f //x=12.03 //y=5.155
c183 ( 42 0 ) capacitor c=0.0939064f //x=15.54 //y=2.08
c184 ( 40 0 ) capacitor c=0.10406f //x=13.69 //y=2.59
c185 ( 36 0 ) capacitor c=0.00398962f //x=13.29 //y=1.665
c186 ( 35 0 ) capacitor c=0.0137288f //x=13.605 //y=1.665
c187 ( 29 0 ) capacitor c=0.0283082f //x=13.605 //y=5.155
c188 ( 21 0 ) capacitor c=0.0176454f //x=12.825 //y=5.155
c189 ( 14 0 ) capacitor c=0.00332903f //x=11.235 //y=5.155
c190 ( 13 0 ) capacitor c=0.0148427f //x=11.945 //y=5.155
c191 ( 2 0 ) capacitor c=0.00808366f //x=13.805 //y=2.59
c192 ( 1 0 ) capacitor c=0.0352679f //x=15.425 //y=2.59
r193 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=16.105 //y=4.79 //x2=16.18 //y2=4.865
r194 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=16.105 //y=4.79 //x2=15.815 //y2=4.79
r195 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.77 //y=1.22 //x2=15.73 //y2=1.375
r196 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.77 //y=0.875 //x2=15.73 //y2=0.72
r197 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.77 //y=0.875 //x2=15.77 //y2=1.22
r198 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.74 //y=4.865 //x2=15.815 //y2=4.79
r199 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=15.74 //y=4.865 //x2=15.54 //y2=4.7
r200 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.395 //y=1.375 //x2=15.28 //y2=1.375
r201 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.615 //y=1.375 //x2=15.73 //y2=1.375
r202 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.395 //y=0.72 //x2=15.28 //y2=0.72
r203 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.615 //y=0.72 //x2=15.73 //y2=0.72
r204 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.615 //y=0.72 //x2=15.395 //y2=0.72
r205 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.915 //x2=15.54 //y2=2.08
r206 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.53 //x2=15.28 //y2=1.375
r207 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.53 //x2=15.24 //y2=1.915
r208 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.22 //x2=15.28 //y2=1.375
r209 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=0.875 //x2=15.28 //y2=0.72
r210 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.24 //y=0.875 //x2=15.24 //y2=1.22
r211 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.18 //y=6.02 //x2=16.18 //y2=4.865
r212 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.74 //y=6.02 //x2=15.74 //y2=4.865
r213 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.505 //y=1.375 //x2=15.615 //y2=1.375
r214 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.505 //y=1.375 //x2=15.395 //y2=1.375
r215 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=4.7 //x2=15.54 //y2=4.7
r216 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=15.54 //y=2.59 //x2=15.54 //y2=4.7
r217 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=2.08 //x2=15.54 //y2=2.08
r218 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=15.54 //y=2.08 //x2=15.54 //y2=2.59
r219 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=13.69 //y=5.07 //x2=13.69 //y2=2.59
r220 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=13.69 //y=1.75 //x2=13.69 //y2=2.59
r221 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.665 //x2=13.69 //y2=1.75
r222 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.665 //x2=13.29 //y2=1.665
r223 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.205 //y=1.58 //x2=13.29 //y2=1.665
r224 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=13.205 //y=1.58 //x2=13.205 //y2=1.01
r225 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.995 //y=5.155 //x2=12.91 //y2=5.155
r226 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.155 //x2=13.69 //y2=5.07
r227 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.155 //x2=12.995 //y2=5.155
r228 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.91 //y=5.24 //x2=12.91 //y2=5.155
r229 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.91 //y=5.24 //x2=12.91 //y2=5.725
r230 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.115 //y=5.155 //x2=12.03 //y2=5.155
r231 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.825 //y=5.155 //x2=12.91 //y2=5.155
r232 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=12.825 //y=5.155 //x2=12.115 //y2=5.155
r233 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.03 //y=5.24 //x2=12.03 //y2=5.155
r234 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.03 //y=5.24 //x2=12.03 //y2=5.725
r235 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.945 //y=5.155 //x2=12.03 //y2=5.155
r236 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.945 //y=5.155 //x2=11.235 //y2=5.155
r237 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.15 //y=5.24 //x2=11.235 //y2=5.155
r238 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.15 //y=5.24 //x2=11.15 //y2=5.725
r239 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=2.59 //x2=15.54 //y2=2.59
r240 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=13.69 //y=2.59 //x2=13.69 //y2=2.59
r241 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.805 //y=2.59 //x2=13.69 //y2=2.59
r242 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=2.59 //x2=15.54 //y2=2.59
r243 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=15.425 //y=2.59 //x2=13.805 //y2=2.59
ends PM_TMRDFFSNRNQNX1\%noxref_4

subckt PM_TMRDFFSNRNQNX1\%noxref_5 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 \
 63 64 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 90 92 98 99 100 101 106 \
 107 112 123 125 126 127 )
c267 ( 127 0 ) capacitor c=0.023087f //x=7.955 //y=5.02
c268 ( 126 0 ) capacitor c=0.023519f //x=7.075 //y=5.02
c269 ( 125 0 ) capacitor c=0.0224735f //x=6.195 //y=5.02
c270 ( 123 0 ) capacitor c=0.00853354f //x=8.205 //y=0.915
c271 ( 112 0 ) capacitor c=0.059212f //x=3.33 //y=4.7
c272 ( 107 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c273 ( 106 0 ) capacitor c=0.045877f //x=3.33 //y=2.08
c274 ( 101 0 ) capacitor c=0.0556143f //x=20.625 //y=4.79
c275 ( 100 0 ) capacitor c=0.0293157f //x=20.915 //y=4.79
c276 ( 99 0 ) capacitor c=0.0347816f //x=20.58 //y=1.22
c277 ( 98 0 ) capacitor c=0.0187487f //x=20.58 //y=0.875
c278 ( 92 0 ) capacitor c=0.0137055f //x=20.425 //y=1.375
c279 ( 90 0 ) capacitor c=0.0149861f //x=20.425 //y=0.72
c280 ( 89 0 ) capacitor c=0.096037f //x=20.05 //y=1.915
c281 ( 88 0 ) capacitor c=0.0228993f //x=20.05 //y=1.53
c282 ( 87 0 ) capacitor c=0.0234352f //x=20.05 //y=1.22
c283 ( 86 0 ) capacitor c=0.0198724f //x=20.05 //y=0.875
c284 ( 85 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c285 ( 84 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c286 ( 81 0 ) capacitor c=0.0148873f //x=3.695 //y=1.415
c287 ( 79 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c288 ( 74 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c289 ( 73 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c290 ( 72 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c291 ( 68 0 ) capacitor c=0.110114f //x=20.99 //y=6.02
c292 ( 67 0 ) capacitor c=0.158956f //x=20.55 //y=6.02
c293 ( 66 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c294 ( 65 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c295 ( 62 0 ) capacitor c=0.00106608f //x=8.1 //y=5.155
c296 ( 61 0 ) capacitor c=0.00207162f //x=7.22 //y=5.155
c297 ( 54 0 ) capacitor c=0.0965808f //x=20.35 //y=2.08
c298 ( 52 0 ) capacitor c=0.10653f //x=8.88 //y=3.33
c299 ( 48 0 ) capacitor c=0.00398962f //x=8.48 //y=1.665
c300 ( 47 0 ) capacitor c=0.0137288f //x=8.795 //y=1.665
c301 ( 41 0 ) capacitor c=0.0283082f //x=8.795 //y=5.155
c302 ( 33 0 ) capacitor c=0.0176454f //x=8.015 //y=5.155
c303 ( 26 0 ) capacitor c=0.00351598f //x=6.425 //y=5.155
c304 ( 25 0 ) capacitor c=0.0154196f //x=7.135 //y=5.155
c305 ( 12 0 ) capacitor c=0.0883624f //x=3.33 //y=2.08
c306 ( 4 0 ) capacitor c=0.00578611f //x=8.995 //y=3.33
c307 ( 3 0 ) capacitor c=0.184375f //x=20.235 //y=3.33
c308 ( 2 0 ) capacitor c=0.0148738f //x=3.445 //y=3.33
c309 ( 1 0 ) capacitor c=0.107193f //x=8.765 //y=3.33
r310 (  106 107 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r311 (  100 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.915 //y=4.79 //x2=20.99 //y2=4.865
r312 (  100 101 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=20.915 //y=4.79 //x2=20.625 //y2=4.79
r313 (  99 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.58 //y=1.22 //x2=20.54 //y2=1.375
r314 (  98 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.58 //y=0.875 //x2=20.54 //y2=0.72
r315 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.58 //y=0.875 //x2=20.58 //y2=1.22
r316 (  95 101 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.55 //y=4.865 //x2=20.625 //y2=4.79
r317 (  95 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=20.55 //y=4.865 //x2=20.35 //y2=4.7
r318 (  93 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.205 //y=1.375 //x2=20.09 //y2=1.375
r319 (  92 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.425 //y=1.375 //x2=20.54 //y2=1.375
r320 (  91 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.205 //y=0.72 //x2=20.09 //y2=0.72
r321 (  90 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.425 //y=0.72 //x2=20.54 //y2=0.72
r322 (  90 91 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.425 //y=0.72 //x2=20.205 //y2=0.72
r323 (  89 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.915 //x2=20.35 //y2=2.08
r324 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.53 //x2=20.09 //y2=1.375
r325 (  88 89 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.53 //x2=20.05 //y2=1.915
r326 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.22 //x2=20.09 //y2=1.375
r327 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=0.875 //x2=20.09 //y2=0.72
r328 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.05 //y=0.875 //x2=20.05 //y2=1.22
r329 (  85 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r330 (  84 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r331 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r332 (  82 110 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r333 (  81 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r334 (  80 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r335 (  79 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r336 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r337 (  76 112 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r338 (  74 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r339 (  74 107 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r340 (  73 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r341 (  72 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r342 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r343 (  69 112 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r344 (  68 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.99 //y=6.02 //x2=20.99 //y2=4.865
r345 (  67 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.55 //y=6.02 //x2=20.55 //y2=4.865
r346 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r347 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r348 (  64 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.315 //y=1.375 //x2=20.425 //y2=1.375
r349 (  64 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.315 //y=1.375 //x2=20.205 //y2=1.375
r350 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r351 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r352 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.35 //y=4.7 //x2=20.35 //y2=4.7
r353 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=20.35 //y=3.33 //x2=20.35 //y2=4.7
r354 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.35 //y=2.08 //x2=20.35 //y2=2.08
r355 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=20.35 //y=2.08 //x2=20.35 //y2=3.33
r356 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=8.88 //y=5.07 //x2=8.88 //y2=3.33
r357 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=8.88 //y=1.75 //x2=8.88 //y2=3.33
r358 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.88 //y2=1.75
r359 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.48 //y2=1.665
r360 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.48 //y2=1.665
r361 (  43 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.395 //y2=1.01
r362 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.185 //y=5.155 //x2=8.1 //y2=5.155
r363 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.88 //y2=5.07
r364 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.185 //y2=5.155
r365 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.155
r366 (  35 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.725
r367 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.305 //y=5.155 //x2=7.22 //y2=5.155
r368 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=8.1 //y2=5.155
r369 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=7.305 //y2=5.155
r370 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.155
r371 (  27 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.725
r372 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=7.22 //y2=5.155
r373 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=6.425 //y2=5.155
r374 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.425 //y2=5.155
r375 (  19 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.34 //y2=5.725
r376 (  17 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r377 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.33 //x2=3.33 //y2=4.7
r378 (  12 106 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r379 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.33
r380 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.35 //y=3.33 //x2=20.35 //y2=3.33
r381 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.88 //y=3.33 //x2=8.88 //y2=3.33
r382 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.33 //x2=3.33 //y2=3.33
r383 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.995 //y=3.33 //x2=8.88 //y2=3.33
r384 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.235 //y=3.33 //x2=20.35 //y2=3.33
r385 (  3 4 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=20.235 //y=3.33 //x2=8.995 //y2=3.33
r386 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.445 //y=3.33 //x2=3.33 //y2=3.33
r387 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=8.88 //y2=3.33
r388 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=3.445 //y2=3.33
ends PM_TMRDFFSNRNQNX1\%noxref_5

subckt PM_TMRDFFSNRNQNX1\%noxref_6 ( 1 2 3 4 6 7 8 9 10 27 28 35 43 49 50 54 \
 58 66 74 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 98 104 105 106 107 \
 111 112 113 114 118 120 123 124 125 126 130 131 132 133 137 139 145 146 156 \
 169 172 174 175 176 )
c634 ( 176 0 ) capacitor c=0.023087f //x=22.385 //y=5.02
c635 ( 175 0 ) capacitor c=0.023519f //x=21.505 //y=5.02
c636 ( 174 0 ) capacitor c=0.0224735f //x=20.625 //y=5.02
c637 ( 172 0 ) capacitor c=0.00853354f //x=22.635 //y=0.915
c638 ( 169 0 ) capacitor c=0.0655948f //x=91.02 //y=4.705
c639 ( 156 0 ) capacitor c=0.054113f //x=87.32 //y=2.08
c640 ( 146 0 ) capacitor c=0.0342409f //x=91.355 //y=1.21
c641 ( 145 0 ) capacitor c=0.0187384f //x=91.355 //y=0.865
c642 ( 139 0 ) capacitor c=0.0141797f //x=91.2 //y=1.365
c643 ( 137 0 ) capacitor c=0.0149844f //x=91.2 //y=0.71
c644 ( 133 0 ) capacitor c=0.0954119f //x=90.825 //y=1.915
c645 ( 132 0 ) capacitor c=0.022465f //x=90.825 //y=1.52
c646 ( 131 0 ) capacitor c=0.0234376f //x=90.825 //y=1.21
c647 ( 130 0 ) capacitor c=0.0199343f //x=90.825 //y=0.865
c648 ( 126 0 ) capacitor c=0.0318948f //x=88.025 //y=1.21
c649 ( 125 0 ) capacitor c=0.0187384f //x=88.025 //y=0.865
c650 ( 124 0 ) capacitor c=0.0605713f //x=87.665 //y=4.795
c651 ( 123 0 ) capacitor c=0.0292043f //x=87.955 //y=4.795
c652 ( 120 0 ) capacitor c=0.0157913f //x=87.87 //y=1.365
c653 ( 118 0 ) capacitor c=0.0149844f //x=87.87 //y=0.71
c654 ( 114 0 ) capacitor c=0.0302441f //x=87.495 //y=1.915
c655 ( 113 0 ) capacitor c=0.0237559f //x=87.495 //y=1.52
c656 ( 112 0 ) capacitor c=0.0234352f //x=87.495 //y=1.21
c657 ( 111 0 ) capacitor c=0.0199931f //x=87.495 //y=0.865
c658 ( 107 0 ) capacitor c=0.0547611f //x=25.435 //y=4.79
c659 ( 106 0 ) capacitor c=0.0294456f //x=25.725 //y=4.79
c660 ( 105 0 ) capacitor c=0.0347816f //x=25.39 //y=1.22
c661 ( 104 0 ) capacitor c=0.0187487f //x=25.39 //y=0.875
c662 ( 98 0 ) capacitor c=0.0137055f //x=25.235 //y=1.375
c663 ( 96 0 ) capacitor c=0.0149861f //x=25.235 //y=0.72
c664 ( 95 0 ) capacitor c=0.096037f //x=24.86 //y=1.915
c665 ( 94 0 ) capacitor c=0.0228993f //x=24.86 //y=1.53
c666 ( 93 0 ) capacitor c=0.0234352f //x=24.86 //y=1.22
c667 ( 92 0 ) capacitor c=0.0198724f //x=24.86 //y=0.875
c668 ( 91 0 ) capacitor c=0.110336f //x=91.35 //y=6.025
c669 ( 90 0 ) capacitor c=0.154049f //x=90.91 //y=6.025
c670 ( 89 0 ) capacitor c=0.110003f //x=88.03 //y=6.025
c671 ( 88 0 ) capacitor c=0.15424f //x=87.59 //y=6.025
c672 ( 87 0 ) capacitor c=0.109949f //x=25.8 //y=6.02
c673 ( 86 0 ) capacitor c=0.158483f //x=25.36 //y=6.02
c674 ( 82 0 ) capacitor c=0.00106608f //x=22.53 //y=5.155
c675 ( 81 0 ) capacitor c=0.00207319f //x=21.65 //y=5.155
c676 ( 74 0 ) capacitor c=0.119551f //x=91.02 //y=2.08
c677 ( 66 0 ) capacitor c=0.0991032f //x=87.32 //y=2.08
c678 ( 58 0 ) capacitor c=0.0910382f //x=25.16 //y=2.08
c679 ( 54 0 ) capacitor c=0.102793f //x=23.31 //y=2.59
c680 ( 50 0 ) capacitor c=0.00398962f //x=22.91 //y=1.665
c681 ( 49 0 ) capacitor c=0.0137288f //x=23.225 //y=1.665
c682 ( 43 0 ) capacitor c=0.0282124f //x=23.225 //y=5.155
c683 ( 35 0 ) capacitor c=0.0176454f //x=22.445 //y=5.155
c684 ( 28 0 ) capacitor c=0.00332903f //x=20.855 //y=5.155
c685 ( 27 0 ) capacitor c=0.0148427f //x=21.565 //y=5.155
c686 ( 10 0 ) capacitor c=0.00638553f //x=87.435 //y=4.44
c687 ( 9 0 ) capacitor c=0.0799095f //x=90.905 //y=4.44
c688 ( 8 0 ) capacitor c=0.00309768f //x=75.195 //y=4.44
c689 ( 7 0 ) capacitor c=0.267484f //x=87.205 //y=4.44
c690 ( 6 0 ) capacitor c=0.00718365f //x=75.11 //y=4.725
c691 ( 4 0 ) capacitor c=0.0158574f //x=23.425 //y=4.81
c692 ( 3 0 ) capacitor c=0.939239f //x=75.025 //y=4.81
c693 ( 2 0 ) capacitor c=0.0116088f //x=23.425 //y=2.59
c694 ( 1 0 ) capacitor c=0.0351856f //x=25.045 //y=2.59
r695 (  167 169 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=90.91 //y=4.705 //x2=91.02 //y2=4.705
r696 (  146 171 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=91.355 //y=1.21 //x2=91.315 //y2=1.365
r697 (  145 170 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=91.355 //y=0.865 //x2=91.315 //y2=0.71
r698 (  145 146 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=91.355 //y=0.865 //x2=91.355 //y2=1.21
r699 (  142 169 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=91.35 //y=4.87 //x2=91.02 //y2=4.705
r700 (  140 166 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=90.98 //y=1.365 //x2=90.865 //y2=1.365
r701 (  139 171 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=91.2 //y=1.365 //x2=91.315 //y2=1.365
r702 (  138 165 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=90.98 //y=0.71 //x2=90.865 //y2=0.71
r703 (  137 170 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=91.2 //y=0.71 //x2=91.315 //y2=0.71
r704 (  137 138 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=91.2 //y=0.71 //x2=90.98 //y2=0.71
r705 (  134 167 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=90.91 //y=4.87 //x2=90.91 //y2=4.705
r706 (  133 164 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=90.825 //y=1.915 //x2=91.02 //y2=2.08
r707 (  132 166 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=90.825 //y=1.52 //x2=90.865 //y2=1.365
r708 (  132 133 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=90.825 //y=1.52 //x2=90.825 //y2=1.915
r709 (  131 166 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=90.825 //y=1.21 //x2=90.865 //y2=1.365
r710 (  130 165 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=90.825 //y=0.865 //x2=90.865 //y2=0.71
r711 (  130 131 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=90.825 //y=0.865 //x2=90.825 //y2=1.21
r712 (  126 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.025 //y=1.21 //x2=87.985 //y2=1.365
r713 (  125 161 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.025 //y=0.865 //x2=87.985 //y2=0.71
r714 (  125 126 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=88.025 //y=0.865 //x2=88.025 //y2=1.21
r715 (  123 127 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=87.955 //y=4.795 //x2=88.03 //y2=4.87
r716 (  123 124 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=87.955 //y=4.795 //x2=87.665 //y2=4.795
r717 (  121 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=87.65 //y=1.365 //x2=87.535 //y2=1.365
r718 (  120 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=87.87 //y=1.365 //x2=87.985 //y2=1.365
r719 (  119 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=87.65 //y=0.71 //x2=87.535 //y2=0.71
r720 (  118 161 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=87.87 //y=0.71 //x2=87.985 //y2=0.71
r721 (  118 119 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=87.87 //y=0.71 //x2=87.65 //y2=0.71
r722 (  115 124 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=87.59 //y=4.87 //x2=87.665 //y2=4.795
r723 (  115 158 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=87.59 //y=4.87 //x2=87.32 //y2=4.705
r724 (  114 156 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=87.495 //y=1.915 //x2=87.32 //y2=2.08
r725 (  113 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=87.495 //y=1.52 //x2=87.535 //y2=1.365
r726 (  113 114 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=87.495 //y=1.52 //x2=87.495 //y2=1.915
r727 (  112 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=87.495 //y=1.21 //x2=87.535 //y2=1.365
r728 (  111 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=87.495 //y=0.865 //x2=87.535 //y2=0.71
r729 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=87.495 //y=0.865 //x2=87.495 //y2=1.21
r730 (  106 108 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=25.725 //y=4.79 //x2=25.8 //y2=4.865
r731 (  106 107 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=25.725 //y=4.79 //x2=25.435 //y2=4.79
r732 (  105 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.39 //y=1.22 //x2=25.35 //y2=1.375
r733 (  104 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.39 //y=0.875 //x2=25.35 //y2=0.72
r734 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=25.39 //y=0.875 //x2=25.39 //y2=1.22
r735 (  101 107 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=25.36 //y=4.865 //x2=25.435 //y2=4.79
r736 (  101 152 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=25.36 //y=4.865 //x2=25.16 //y2=4.7
r737 (  99 148 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.015 //y=1.375 //x2=24.9 //y2=1.375
r738 (  98 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.235 //y=1.375 //x2=25.35 //y2=1.375
r739 (  97 147 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.015 //y=0.72 //x2=24.9 //y2=0.72
r740 (  96 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.235 //y=0.72 //x2=25.35 //y2=0.72
r741 (  96 97 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=25.235 //y=0.72 //x2=25.015 //y2=0.72
r742 (  95 150 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.915 //x2=25.16 //y2=2.08
r743 (  94 148 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.53 //x2=24.9 //y2=1.375
r744 (  94 95 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.53 //x2=24.86 //y2=1.915
r745 (  93 148 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.22 //x2=24.9 //y2=1.375
r746 (  92 147 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=0.875 //x2=24.9 //y2=0.72
r747 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.86 //y=0.875 //x2=24.86 //y2=1.22
r748 (  91 142 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=91.35 //y=6.025 //x2=91.35 //y2=4.87
r749 (  90 134 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=90.91 //y=6.025 //x2=90.91 //y2=4.87
r750 (  89 127 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=88.03 //y=6.025 //x2=88.03 //y2=4.87
r751 (  88 115 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=87.59 //y=6.025 //x2=87.59 //y2=4.87
r752 (  87 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.8 //y=6.02 //x2=25.8 //y2=4.865
r753 (  86 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.36 //y=6.02 //x2=25.36 //y2=4.865
r754 (  85 139 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=91.09 //y=1.365 //x2=91.2 //y2=1.365
r755 (  85 140 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=91.09 //y=1.365 //x2=90.98 //y2=1.365
r756 (  84 120 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=87.76 //y=1.365 //x2=87.87 //y2=1.365
r757 (  84 121 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=87.76 //y=1.365 //x2=87.65 //y2=1.365
r758 (  83 98 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.125 //y=1.375 //x2=25.235 //y2=1.375
r759 (  83 99 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.125 //y=1.375 //x2=25.015 //y2=1.375
r760 (  79 169 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=91.02 //y=4.705 //x2=91.02 //y2=4.705
r761 (  77 79 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=91.02 //y=4.44 //x2=91.02 //y2=4.705
r762 (  74 164 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=91.02 //y=2.08 //x2=91.02 //y2=2.08
r763 (  74 77 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=91.02 //y=2.08 //x2=91.02 //y2=4.44
r764 (  71 158 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=87.32 //y=4.705 //x2=87.32 //y2=4.705
r765 (  69 71 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=87.32 //y=4.44 //x2=87.32 //y2=4.705
r766 (  66 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=87.32 //y=2.08 //x2=87.32 //y2=2.08
r767 (  66 69 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=87.32 //y=2.08 //x2=87.32 //y2=4.44
r768 (  63 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.16 //y=4.7 //x2=25.16 //y2=4.7
r769 (  61 63 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.59 //x2=25.16 //y2=4.7
r770 (  58 150 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.16 //y=2.08 //x2=25.16 //y2=2.08
r771 (  58 61 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.08 //x2=25.16 //y2=2.59
r772 (  54 56 ) resistor r=151.957 //w=0.187 //l=2.22 //layer=li \
 //thickness=0.1 //x=23.31 //y=2.59 //x2=23.31 //y2=4.81
r773 (  52 56 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=23.31 //y=5.07 //x2=23.31 //y2=4.81
r774 (  51 54 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=23.31 //y=1.75 //x2=23.31 //y2=2.59
r775 (  49 51 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.225 //y=1.665 //x2=23.31 //y2=1.75
r776 (  49 50 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=23.225 //y=1.665 //x2=22.91 //y2=1.665
r777 (  45 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=22.825 //y=1.58 //x2=22.91 //y2=1.665
r778 (  45 172 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=22.825 //y=1.58 //x2=22.825 //y2=1.01
r779 (  44 82 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.615 //y=5.155 //x2=22.53 //y2=5.155
r780 (  43 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.225 //y=5.155 //x2=23.31 //y2=5.07
r781 (  43 44 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=23.225 //y=5.155 //x2=22.615 //y2=5.155
r782 (  37 82 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.53 //y=5.24 //x2=22.53 //y2=5.155
r783 (  37 176 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.53 //y=5.24 //x2=22.53 //y2=5.725
r784 (  36 81 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.735 //y=5.155 //x2=21.65 //y2=5.155
r785 (  35 82 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.445 //y=5.155 //x2=22.53 //y2=5.155
r786 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.445 //y=5.155 //x2=21.735 //y2=5.155
r787 (  29 81 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.65 //y=5.24 //x2=21.65 //y2=5.155
r788 (  29 175 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.65 //y=5.24 //x2=21.65 //y2=5.725
r789 (  27 81 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.565 //y=5.155 //x2=21.65 //y2=5.155
r790 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=21.565 //y=5.155 //x2=20.855 //y2=5.155
r791 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.77 //y=5.24 //x2=20.855 //y2=5.155
r792 (  21 174 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.77 //y=5.24 //x2=20.77 //y2=5.725
r793 (  20 77 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=91.02 //y=4.44 //x2=91.02 //y2=4.44
r794 (  18 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=87.32 //y=4.44 //x2=87.32 //y2=4.44
r795 (  16 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.16 //y=2.59 //x2=25.16 //y2=2.59
r796 (  14 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.31 //y=4.81 //x2=23.31 //y2=4.81
r797 (  12 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.31 //y=2.59 //x2=23.31 //y2=2.59
r798 (  10 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=87.435 //y=4.44 //x2=87.32 //y2=4.44
r799 (  9 20 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=90.905 //y=4.44 //x2=91.02 //y2=4.44
r800 (  9 10 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=90.905 //y=4.44 //x2=87.435 //y2=4.44
r801 (  7 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=87.205 //y=4.44 //x2=87.32 //y2=4.44
r802 (  7 8 ) resistor r=11.4599 //w=0.131 //l=12.01 //layer=m1 \
 //thickness=0.36 //x=87.205 //y=4.44 //x2=75.195 //y2=4.44
r803 (  5 8 ) resistor r=0.0718295 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=4.525 //x2=75.195 //y2=4.44
r804 (  5 6 ) resistor r=0.19084 //w=0.131 //l=0.2 //layer=m1 //thickness=0.36 \
 //x=75.11 //y=4.525 //x2=75.11 //y2=4.725
r805 (  4 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.425 //y=4.81 //x2=23.31 //y2=4.81
r806 (  3 6 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=75.025 //y=4.81 //x2=75.11 //y2=4.725
r807 (  3 4 ) resistor r=49.2366 //w=0.131 //l=51.6 //layer=m1 \
 //thickness=0.36 //x=75.025 //y=4.81 //x2=23.425 //y2=4.81
r808 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.425 //y=2.59 //x2=23.31 //y2=2.59
r809 (  1 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.045 //y=2.59 //x2=25.16 //y2=2.59
r810 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=25.045 //y=2.59 //x2=23.425 //y2=2.59
ends PM_TMRDFFSNRNQNX1\%noxref_6

subckt PM_TMRDFFSNRNQNX1\%noxref_7 ( 1 2 3 4 5 6 16 24 37 38 45 53 59 60 64 66 \
 73 74 75 76 77 78 79 80 81 82 83 87 88 89 94 96 99 100 104 105 106 111 113 \
 116 117 121 122 123 128 130 133 134 136 137 142 146 147 152 156 157 162 165 \
 167 168 169 )
c339 ( 169 0 ) capacitor c=0.023087f //x=17.575 //y=5.02
c340 ( 168 0 ) capacitor c=0.023519f //x=16.695 //y=5.02
c341 ( 167 0 ) capacitor c=0.0224735f //x=15.815 //y=5.02
c342 ( 165 0 ) capacitor c=0.00853354f //x=17.825 //y=0.915
c343 ( 162 0 ) capacitor c=0.0588394f //x=27.38 //y=4.7
c344 ( 157 0 ) capacitor c=0.0273931f //x=27.38 //y=1.915
c345 ( 156 0 ) capacitor c=0.0456313f //x=27.38 //y=2.08
c346 ( 152 0 ) capacitor c=0.0587755f //x=12.95 //y=4.7
c347 ( 147 0 ) capacitor c=0.0273931f //x=12.95 //y=1.915
c348 ( 146 0 ) capacitor c=0.0456313f //x=12.95 //y=2.08
c349 ( 142 0 ) capacitor c=0.058931f //x=8.14 //y=4.7
c350 ( 137 0 ) capacitor c=0.0273931f //x=8.14 //y=1.915
c351 ( 136 0 ) capacitor c=0.0456313f //x=8.14 //y=2.08
c352 ( 134 0 ) capacitor c=0.0432517f //x=27.9 //y=1.26
c353 ( 133 0 ) capacitor c=0.0200379f //x=27.9 //y=0.915
c354 ( 130 0 ) capacitor c=0.0148873f //x=27.745 //y=1.415
c355 ( 128 0 ) capacitor c=0.0157803f //x=27.745 //y=0.76
c356 ( 123 0 ) capacitor c=0.0218028f //x=27.37 //y=1.57
c357 ( 122 0 ) capacitor c=0.0207459f //x=27.37 //y=1.26
c358 ( 121 0 ) capacitor c=0.0194308f //x=27.37 //y=0.915
c359 ( 117 0 ) capacitor c=0.0432517f //x=13.47 //y=1.26
c360 ( 116 0 ) capacitor c=0.0200379f //x=13.47 //y=0.915
c361 ( 113 0 ) capacitor c=0.0148873f //x=13.315 //y=1.415
c362 ( 111 0 ) capacitor c=0.0157803f //x=13.315 //y=0.76
c363 ( 106 0 ) capacitor c=0.0218028f //x=12.94 //y=1.57
c364 ( 105 0 ) capacitor c=0.0207459f //x=12.94 //y=1.26
c365 ( 104 0 ) capacitor c=0.0194308f //x=12.94 //y=0.915
c366 ( 100 0 ) capacitor c=0.0432517f //x=8.66 //y=1.26
c367 ( 99 0 ) capacitor c=0.0200379f //x=8.66 //y=0.915
c368 ( 96 0 ) capacitor c=0.0148873f //x=8.505 //y=1.415
c369 ( 94 0 ) capacitor c=0.0157803f //x=8.505 //y=0.76
c370 ( 89 0 ) capacitor c=0.0218028f //x=8.13 //y=1.57
c371 ( 88 0 ) capacitor c=0.0207459f //x=8.13 //y=1.26
c372 ( 87 0 ) capacitor c=0.0194308f //x=8.13 //y=0.915
c373 ( 83 0 ) capacitor c=0.158754f //x=27.56 //y=6.02
c374 ( 82 0 ) capacitor c=0.109949f //x=27.12 //y=6.02
c375 ( 81 0 ) capacitor c=0.158794f //x=13.13 //y=6.02
c376 ( 80 0 ) capacitor c=0.110114f //x=12.69 //y=6.02
c377 ( 79 0 ) capacitor c=0.158794f //x=8.32 //y=6.02
c378 ( 78 0 ) capacitor c=0.110114f //x=7.88 //y=6.02
c379 ( 74 0 ) capacitor c=0.00106608f //x=17.72 //y=5.155
c380 ( 73 0 ) capacitor c=0.00207162f //x=16.84 //y=5.155
c381 ( 66 0 ) capacitor c=0.0796271f //x=27.38 //y=2.08
c382 ( 64 0 ) capacitor c=0.105458f //x=18.5 //y=3.7
c383 ( 60 0 ) capacitor c=0.00398962f //x=18.1 //y=1.665
c384 ( 59 0 ) capacitor c=0.0137288f //x=18.415 //y=1.665
c385 ( 53 0 ) capacitor c=0.0283082f //x=18.415 //y=5.155
c386 ( 45 0 ) capacitor c=0.0176454f //x=17.635 //y=5.155
c387 ( 38 0 ) capacitor c=0.00332903f //x=16.045 //y=5.155
c388 ( 37 0 ) capacitor c=0.014837f //x=16.755 //y=5.155
c389 ( 24 0 ) capacitor c=0.0810736f //x=12.95 //y=2.08
c390 ( 16 0 ) capacitor c=0.0819749f //x=8.14 //y=2.08
c391 ( 6 0 ) capacitor c=0.0055354f //x=18.615 //y=3.7
c392 ( 5 0 ) capacitor c=0.145577f //x=27.265 //y=3.7
c393 ( 4 0 ) capacitor c=0.00556898f //x=13.065 //y=3.7
c394 ( 3 0 ) capacitor c=0.0758356f //x=18.385 //y=3.7
c395 ( 2 0 ) capacitor c=0.0138772f //x=8.255 //y=3.7
c396 ( 1 0 ) capacitor c=0.067053f //x=12.835 //y=3.7
r397 (  156 157 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=27.38 //y=2.08 //x2=27.38 //y2=1.915
r398 (  146 147 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=12.95 //y=2.08 //x2=12.95 //y2=1.915
r399 (  136 137 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.14 //y=2.08 //x2=8.14 //y2=1.915
r400 (  134 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.9 //y=1.26 //x2=27.86 //y2=1.415
r401 (  133 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.9 //y=0.915 //x2=27.86 //y2=0.76
r402 (  133 134 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.9 //y=0.915 //x2=27.9 //y2=1.26
r403 (  131 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.525 //y=1.415 //x2=27.41 //y2=1.415
r404 (  130 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.745 //y=1.415 //x2=27.86 //y2=1.415
r405 (  129 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.525 //y=0.76 //x2=27.41 //y2=0.76
r406 (  128 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.745 //y=0.76 //x2=27.86 //y2=0.76
r407 (  128 129 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=27.745 //y=0.76 //x2=27.525 //y2=0.76
r408 (  125 162 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=27.56 //y=4.865 //x2=27.38 //y2=4.7
r409 (  123 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.57 //x2=27.41 //y2=1.415
r410 (  123 157 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.57 //x2=27.37 //y2=1.915
r411 (  122 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.26 //x2=27.41 //y2=1.415
r412 (  121 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=0.915 //x2=27.41 //y2=0.76
r413 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.37 //y=0.915 //x2=27.37 //y2=1.26
r414 (  118 162 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=27.12 //y=4.865 //x2=27.38 //y2=4.7
r415 (  117 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.47 //y=1.26 //x2=13.43 //y2=1.415
r416 (  116 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.47 //y=0.915 //x2=13.43 //y2=0.76
r417 (  116 117 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.47 //y=0.915 //x2=13.47 //y2=1.26
r418 (  114 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.095 //y=1.415 //x2=12.98 //y2=1.415
r419 (  113 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.315 //y=1.415 //x2=13.43 //y2=1.415
r420 (  112 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.095 //y=0.76 //x2=12.98 //y2=0.76
r421 (  111 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.315 //y=0.76 //x2=13.43 //y2=0.76
r422 (  111 112 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=13.315 //y=0.76 //x2=13.095 //y2=0.76
r423 (  108 152 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=13.13 //y=4.865 //x2=12.95 //y2=4.7
r424 (  106 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.57 //x2=12.98 //y2=1.415
r425 (  106 147 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.57 //x2=12.94 //y2=1.915
r426 (  105 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.26 //x2=12.98 //y2=1.415
r427 (  104 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=0.915 //x2=12.98 //y2=0.76
r428 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.94 //y=0.915 //x2=12.94 //y2=1.26
r429 (  101 152 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=12.69 //y=4.865 //x2=12.95 //y2=4.7
r430 (  100 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=1.26 //x2=8.62 //y2=1.415
r431 (  99 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.62 //y2=0.76
r432 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.66 //y2=1.26
r433 (  97 140 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=1.415 //x2=8.17 //y2=1.415
r434 (  96 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=1.415 //x2=8.62 //y2=1.415
r435 (  95 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=0.76 //x2=8.17 //y2=0.76
r436 (  94 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.62 //y2=0.76
r437 (  94 95 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.285 //y2=0.76
r438 (  91 142 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=8.32 //y=4.865 //x2=8.14 //y2=4.7
r439 (  89 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.17 //y2=1.415
r440 (  89 137 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.13 //y2=1.915
r441 (  88 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.26 //x2=8.17 //y2=1.415
r442 (  87 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.17 //y2=0.76
r443 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.13 //y2=1.26
r444 (  84 142 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=7.88 //y=4.865 //x2=8.14 //y2=4.7
r445 (  83 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.56 //y=6.02 //x2=27.56 //y2=4.865
r446 (  82 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.12 //y=6.02 //x2=27.12 //y2=4.865
r447 (  81 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.13 //y=6.02 //x2=13.13 //y2=4.865
r448 (  80 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.69 //y=6.02 //x2=12.69 //y2=4.865
r449 (  79 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.32 //y=6.02 //x2=8.32 //y2=4.865
r450 (  78 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.88 //y=6.02 //x2=7.88 //y2=4.865
r451 (  77 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.635 //y=1.415 //x2=27.745 //y2=1.415
r452 (  77 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.635 //y=1.415 //x2=27.525 //y2=1.415
r453 (  76 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.205 //y=1.415 //x2=13.315 //y2=1.415
r454 (  76 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.205 //y=1.415 //x2=13.095 //y2=1.415
r455 (  75 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.505 //y2=1.415
r456 (  75 97 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.285 //y2=1.415
r457 (  71 162 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=4.7 //x2=27.38 //y2=4.7
r458 (  69 71 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=27.38 //y=3.7 //x2=27.38 //y2=4.7
r459 (  66 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=2.08 //x2=27.38 //y2=2.08
r460 (  66 69 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=27.38 //y=2.08 //x2=27.38 //y2=3.7
r461 (  62 64 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=18.5 //y=5.07 //x2=18.5 //y2=3.7
r462 (  61 64 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=18.5 //y=1.75 //x2=18.5 //y2=3.7
r463 (  59 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.415 //y=1.665 //x2=18.5 //y2=1.75
r464 (  59 60 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=18.415 //y=1.665 //x2=18.1 //y2=1.665
r465 (  55 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.015 //y=1.58 //x2=18.1 //y2=1.665
r466 (  55 165 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=18.015 //y=1.58 //x2=18.015 //y2=1.01
r467 (  54 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.805 //y=5.155 //x2=17.72 //y2=5.155
r468 (  53 62 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.415 //y=5.155 //x2=18.5 //y2=5.07
r469 (  53 54 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=18.415 //y=5.155 //x2=17.805 //y2=5.155
r470 (  47 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.72 //y=5.24 //x2=17.72 //y2=5.155
r471 (  47 169 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.72 //y=5.24 //x2=17.72 //y2=5.725
r472 (  46 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.925 //y=5.155 //x2=16.84 //y2=5.155
r473 (  45 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.635 //y=5.155 //x2=17.72 //y2=5.155
r474 (  45 46 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=17.635 //y=5.155 //x2=16.925 //y2=5.155
r475 (  39 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.84 //y=5.24 //x2=16.84 //y2=5.155
r476 (  39 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.84 //y=5.24 //x2=16.84 //y2=5.725
r477 (  37 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.755 //y=5.155 //x2=16.84 //y2=5.155
r478 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.755 //y=5.155 //x2=16.045 //y2=5.155
r479 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.96 //y=5.24 //x2=16.045 //y2=5.155
r480 (  31 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.96 //y=5.24 //x2=15.96 //y2=5.725
r481 (  29 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.95 //y=4.7 //x2=12.95 //y2=4.7
r482 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=12.95 //y=3.7 //x2=12.95 //y2=4.7
r483 (  24 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.95 //y=2.08 //x2=12.95 //y2=2.08
r484 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=12.95 //y=2.08 //x2=12.95 //y2=3.7
r485 (  21 142 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=4.7 //x2=8.14 //y2=4.7
r486 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=8.14 //y=3.7 //x2=8.14 //y2=4.7
r487 (  16 136 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=2.08 //x2=8.14 //y2=2.08
r488 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.08 //x2=8.14 //y2=3.7
r489 (  14 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=27.38 //y=3.7 //x2=27.38 //y2=3.7
r490 (  12 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.5 //y=3.7 //x2=18.5 //y2=3.7
r491 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.95 //y=3.7 //x2=12.95 //y2=3.7
r492 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.14 //y=3.7 //x2=8.14 //y2=3.7
r493 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.615 //y=3.7 //x2=18.5 //y2=3.7
r494 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.265 //y=3.7 //x2=27.38 //y2=3.7
r495 (  5 6 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=27.265 //y=3.7 //x2=18.615 //y2=3.7
r496 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.065 //y=3.7 //x2=12.95 //y2=3.7
r497 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=3.7 //x2=18.5 //y2=3.7
r498 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=3.7 //x2=13.065 //y2=3.7
r499 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.255 //y=3.7 //x2=8.14 //y2=3.7
r500 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.835 //y=3.7 //x2=12.95 //y2=3.7
r501 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=12.835 //y=3.7 //x2=8.255 //y2=3.7
ends PM_TMRDFFSNRNQNX1\%noxref_7

subckt PM_TMRDFFSNRNQNX1\%noxref_8 ( 1 2 8 21 22 29 37 43 44 48 49 50 51 52 53 \
 57 58 59 64 66 69 70 72 73 78 81 83 84 85 )
c176 ( 85 0 ) capacitor c=0.023087f //x=27.195 //y=5.02
c177 ( 84 0 ) capacitor c=0.023519f //x=26.315 //y=5.02
c178 ( 83 0 ) capacitor c=0.0224735f //x=25.435 //y=5.02
c179 ( 81 0 ) capacitor c=0.00853354f //x=27.445 //y=0.915
c180 ( 78 0 ) capacitor c=0.0587755f //x=22.57 //y=4.7
c181 ( 73 0 ) capacitor c=0.0273931f //x=22.57 //y=1.915
c182 ( 72 0 ) capacitor c=0.0456313f //x=22.57 //y=2.08
c183 ( 70 0 ) capacitor c=0.0432517f //x=23.09 //y=1.26
c184 ( 69 0 ) capacitor c=0.0200379f //x=23.09 //y=0.915
c185 ( 66 0 ) capacitor c=0.0148873f //x=22.935 //y=1.415
c186 ( 64 0 ) capacitor c=0.0157803f //x=22.935 //y=0.76
c187 ( 59 0 ) capacitor c=0.0218028f //x=22.56 //y=1.57
c188 ( 58 0 ) capacitor c=0.0207459f //x=22.56 //y=1.26
c189 ( 57 0 ) capacitor c=0.0194308f //x=22.56 //y=0.915
c190 ( 53 0 ) capacitor c=0.158794f //x=22.75 //y=6.02
c191 ( 52 0 ) capacitor c=0.110114f //x=22.31 //y=6.02
c192 ( 50 0 ) capacitor c=9.74268e-19 //x=27.34 //y=5.155
c193 ( 49 0 ) capacitor c=0.00191414f //x=26.46 //y=5.155
c194 ( 48 0 ) capacitor c=0.107305f //x=28.12 //y=3.33
c195 ( 44 0 ) capacitor c=0.00398962f //x=27.72 //y=1.665
c196 ( 43 0 ) capacitor c=0.0137288f //x=28.035 //y=1.665
c197 ( 37 0 ) capacitor c=0.0276208f //x=28.035 //y=5.155
c198 ( 29 0 ) capacitor c=0.0169868f //x=27.255 //y=5.155
c199 ( 22 0 ) capacitor c=0.00316998f //x=25.665 //y=5.155
c200 ( 21 0 ) capacitor c=0.014258f //x=26.375 //y=5.155
c201 ( 8 0 ) capacitor c=0.0820026f //x=22.57 //y=2.08
c202 ( 2 0 ) capacitor c=0.00906635f //x=22.685 //y=3.33
c203 ( 1 0 ) capacitor c=0.0884963f //x=28.005 //y=3.33
r204 (  72 73 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=22.57 //y=2.08 //x2=22.57 //y2=1.915
r205 (  70 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.09 //y=1.26 //x2=23.05 //y2=1.415
r206 (  69 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.09 //y=0.915 //x2=23.05 //y2=0.76
r207 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.09 //y=0.915 //x2=23.09 //y2=1.26
r208 (  67 76 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.715 //y=1.415 //x2=22.6 //y2=1.415
r209 (  66 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.935 //y=1.415 //x2=23.05 //y2=1.415
r210 (  65 75 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.715 //y=0.76 //x2=22.6 //y2=0.76
r211 (  64 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.935 //y=0.76 //x2=23.05 //y2=0.76
r212 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=22.935 //y=0.76 //x2=22.715 //y2=0.76
r213 (  61 78 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=22.75 //y=4.865 //x2=22.57 //y2=4.7
r214 (  59 76 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.57 //x2=22.6 //y2=1.415
r215 (  59 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.57 //x2=22.56 //y2=1.915
r216 (  58 76 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.26 //x2=22.6 //y2=1.415
r217 (  57 75 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=0.915 //x2=22.6 //y2=0.76
r218 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.56 //y=0.915 //x2=22.56 //y2=1.26
r219 (  54 78 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=22.31 //y=4.865 //x2=22.57 //y2=4.7
r220 (  53 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.75 //y=6.02 //x2=22.75 //y2=4.865
r221 (  52 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.31 //y=6.02 //x2=22.31 //y2=4.865
r222 (  51 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.825 //y=1.415 //x2=22.935 //y2=1.415
r223 (  51 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.825 //y=1.415 //x2=22.715 //y2=1.415
r224 (  46 48 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=28.12 //y=5.07 //x2=28.12 //y2=3.33
r225 (  45 48 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=28.12 //y=1.75 //x2=28.12 //y2=3.33
r226 (  43 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.035 //y=1.665 //x2=28.12 //y2=1.75
r227 (  43 44 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=28.035 //y=1.665 //x2=27.72 //y2=1.665
r228 (  39 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=27.635 //y=1.58 //x2=27.72 //y2=1.665
r229 (  39 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=27.635 //y=1.58 //x2=27.635 //y2=1.01
r230 (  38 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.425 //y=5.155 //x2=27.34 //y2=5.155
r231 (  37 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.035 //y=5.155 //x2=28.12 //y2=5.07
r232 (  37 38 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=28.035 //y=5.155 //x2=27.425 //y2=5.155
r233 (  31 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.34 //y=5.24 //x2=27.34 //y2=5.155
r234 (  31 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.34 //y=5.24 //x2=27.34 //y2=5.725
r235 (  30 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.545 //y=5.155 //x2=26.46 //y2=5.155
r236 (  29 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.255 //y=5.155 //x2=27.34 //y2=5.155
r237 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=27.255 //y=5.155 //x2=26.545 //y2=5.155
r238 (  23 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.46 //y=5.24 //x2=26.46 //y2=5.155
r239 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.46 //y=5.24 //x2=26.46 //y2=5.725
r240 (  21 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.375 //y=5.155 //x2=26.46 //y2=5.155
r241 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.375 //y=5.155 //x2=25.665 //y2=5.155
r242 (  15 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.58 //y=5.24 //x2=25.665 //y2=5.155
r243 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=25.58 //y=5.24 //x2=25.58 //y2=5.725
r244 (  13 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=4.7 //x2=22.57 //y2=4.7
r245 (  11 13 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=22.57 //y=3.33 //x2=22.57 //y2=4.7
r246 (  8 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=2.08 //x2=22.57 //y2=2.08
r247 (  8 11 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=22.57 //y=2.08 //x2=22.57 //y2=3.33
r248 (  6 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.12 //y=3.33 //x2=28.12 //y2=3.33
r249 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=22.57 //y=3.33 //x2=22.57 //y2=3.33
r250 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=22.685 //y=3.33 //x2=22.57 //y2=3.33
r251 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=3.33 //x2=28.12 //y2=3.33
r252 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=3.33 //x2=22.685 //y2=3.33
ends PM_TMRDFFSNRNQNX1\%noxref_8

subckt PM_TMRDFFSNRNQNX1\%noxref_9 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 \
 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c253 ( 127 0 ) capacitor c=0.023087f //x=32.005 //y=5.02
c254 ( 126 0 ) capacitor c=0.023519f //x=31.125 //y=5.02
c255 ( 125 0 ) capacitor c=0.0224735f //x=30.245 //y=5.02
c256 ( 123 0 ) capacitor c=0.00853354f //x=32.255 //y=0.915
c257 ( 103 0 ) capacitor c=0.0547611f //x=39.865 //y=4.79
c258 ( 102 0 ) capacitor c=0.0294456f //x=40.155 //y=4.79
c259 ( 101 0 ) capacitor c=0.0347816f //x=39.82 //y=1.22
c260 ( 100 0 ) capacitor c=0.0187487f //x=39.82 //y=0.875
c261 ( 94 0 ) capacitor c=0.0137055f //x=39.665 //y=1.375
c262 ( 92 0 ) capacitor c=0.0149861f //x=39.665 //y=0.72
c263 ( 91 0 ) capacitor c=0.096037f //x=39.29 //y=1.915
c264 ( 90 0 ) capacitor c=0.0228993f //x=39.29 //y=1.53
c265 ( 89 0 ) capacitor c=0.0234352f //x=39.29 //y=1.22
c266 ( 88 0 ) capacitor c=0.0198724f //x=39.29 //y=0.875
c267 ( 84 0 ) capacitor c=0.0549166f //x=35.055 //y=4.79
c268 ( 83 0 ) capacitor c=0.0294456f //x=35.345 //y=4.79
c269 ( 82 0 ) capacitor c=0.0347816f //x=35.01 //y=1.22
c270 ( 81 0 ) capacitor c=0.0187487f //x=35.01 //y=0.875
c271 ( 75 0 ) capacitor c=0.0137055f //x=34.855 //y=1.375
c272 ( 73 0 ) capacitor c=0.0149861f //x=34.855 //y=0.72
c273 ( 72 0 ) capacitor c=0.096037f //x=34.48 //y=1.915
c274 ( 71 0 ) capacitor c=0.0228993f //x=34.48 //y=1.53
c275 ( 70 0 ) capacitor c=0.0234352f //x=34.48 //y=1.22
c276 ( 69 0 ) capacitor c=0.0198724f //x=34.48 //y=0.875
c277 ( 68 0 ) capacitor c=0.109949f //x=40.23 //y=6.02
c278 ( 67 0 ) capacitor c=0.158483f //x=39.79 //y=6.02
c279 ( 66 0 ) capacitor c=0.109949f //x=35.42 //y=6.02
c280 ( 65 0 ) capacitor c=0.158483f //x=34.98 //y=6.02
c281 ( 62 0 ) capacitor c=9.74268e-19 //x=32.15 //y=5.155
c282 ( 61 0 ) capacitor c=0.00191414f //x=31.27 //y=5.155
c283 ( 54 0 ) capacitor c=0.0914984f //x=39.59 //y=2.08
c284 ( 46 0 ) capacitor c=0.0942434f //x=34.78 //y=2.08
c285 ( 44 0 ) capacitor c=0.106133f //x=32.93 //y=2.59
c286 ( 40 0 ) capacitor c=0.00398962f //x=32.53 //y=1.665
c287 ( 39 0 ) capacitor c=0.0137288f //x=32.845 //y=1.665
c288 ( 33 0 ) capacitor c=0.0276208f //x=32.845 //y=5.155
c289 ( 25 0 ) capacitor c=0.0169868f //x=32.065 //y=5.155
c290 ( 18 0 ) capacitor c=0.00316998f //x=30.475 //y=5.155
c291 ( 17 0 ) capacitor c=0.014258f //x=31.185 //y=5.155
c292 ( 4 0 ) capacitor c=0.00401138f //x=34.895 //y=2.59
c293 ( 3 0 ) capacitor c=0.0706637f //x=39.475 //y=2.59
c294 ( 2 0 ) capacitor c=0.0120752f //x=33.045 //y=2.59
c295 ( 1 0 ) capacitor c=0.0233554f //x=34.665 //y=2.59
r296 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=40.155 //y=4.79 //x2=40.23 //y2=4.865
r297 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=40.155 //y=4.79 //x2=39.865 //y2=4.79
r298 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.82 //y=1.22 //x2=39.78 //y2=1.375
r299 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.82 //y=0.875 //x2=39.78 //y2=0.72
r300 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=39.82 //y=0.875 //x2=39.82 //y2=1.22
r301 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=39.79 //y=4.865 //x2=39.865 //y2=4.79
r302 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=39.79 //y=4.865 //x2=39.59 //y2=4.7
r303 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.445 //y=1.375 //x2=39.33 //y2=1.375
r304 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.665 //y=1.375 //x2=39.78 //y2=1.375
r305 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.445 //y=0.72 //x2=39.33 //y2=0.72
r306 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.665 //y=0.72 //x2=39.78 //y2=0.72
r307 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=39.665 //y=0.72 //x2=39.445 //y2=0.72
r308 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=39.29 //y=1.915 //x2=39.59 //y2=2.08
r309 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.29 //y=1.53 //x2=39.33 //y2=1.375
r310 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=39.29 //y=1.53 //x2=39.29 //y2=1.915
r311 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.29 //y=1.22 //x2=39.33 //y2=1.375
r312 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.29 //y=0.875 //x2=39.33 //y2=0.72
r313 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=39.29 //y=0.875 //x2=39.29 //y2=1.22
r314 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=35.345 //y=4.79 //x2=35.42 //y2=4.865
r315 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=35.345 //y=4.79 //x2=35.055 //y2=4.79
r316 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.01 //y=1.22 //x2=34.97 //y2=1.375
r317 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.01 //y=0.875 //x2=34.97 //y2=0.72
r318 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=35.01 //y=0.875 //x2=35.01 //y2=1.22
r319 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=34.98 //y=4.865 //x2=35.055 //y2=4.79
r320 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=34.98 //y=4.865 //x2=34.78 //y2=4.7
r321 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.635 //y=1.375 //x2=34.52 //y2=1.375
r322 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.855 //y=1.375 //x2=34.97 //y2=1.375
r323 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.635 //y=0.72 //x2=34.52 //y2=0.72
r324 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.855 //y=0.72 //x2=34.97 //y2=0.72
r325 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=34.855 //y=0.72 //x2=34.635 //y2=0.72
r326 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.915 //x2=34.78 //y2=2.08
r327 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.53 //x2=34.52 //y2=1.375
r328 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.53 //x2=34.48 //y2=1.915
r329 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.22 //x2=34.52 //y2=1.375
r330 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.48 //y=0.875 //x2=34.52 //y2=0.72
r331 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=34.48 //y=0.875 //x2=34.48 //y2=1.22
r332 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=40.23 //y=6.02 //x2=40.23 //y2=4.865
r333 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=39.79 //y=6.02 //x2=39.79 //y2=4.865
r334 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.42 //y=6.02 //x2=35.42 //y2=4.865
r335 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.98 //y=6.02 //x2=34.98 //y2=4.865
r336 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.555 //y=1.375 //x2=39.665 //y2=1.375
r337 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.555 //y=1.375 //x2=39.445 //y2=1.375
r338 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.745 //y=1.375 //x2=34.855 //y2=1.375
r339 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.745 //y=1.375 //x2=34.635 //y2=1.375
r340 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.59 //y=4.7 //x2=39.59 //y2=4.7
r341 (  57 59 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=39.59 //y=2.59 //x2=39.59 //y2=4.7
r342 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.59 //y=2.08 //x2=39.59 //y2=2.08
r343 (  54 57 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=39.59 //y=2.08 //x2=39.59 //y2=2.59
r344 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.78 //y=4.7 //x2=34.78 //y2=4.7
r345 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=34.78 //y=2.59 //x2=34.78 //y2=4.7
r346 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.78 //y=2.08 //x2=34.78 //y2=2.08
r347 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=34.78 //y=2.08 //x2=34.78 //y2=2.59
r348 (  42 44 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=32.93 //y=5.07 //x2=32.93 //y2=2.59
r349 (  41 44 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=32.93 //y=1.75 //x2=32.93 //y2=2.59
r350 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.845 //y=1.665 //x2=32.93 //y2=1.75
r351 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=32.845 //y=1.665 //x2=32.53 //y2=1.665
r352 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.445 //y=1.58 //x2=32.53 //y2=1.665
r353 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=32.445 //y=1.58 //x2=32.445 //y2=1.01
r354 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.235 //y=5.155 //x2=32.15 //y2=5.155
r355 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.845 //y=5.155 //x2=32.93 //y2=5.07
r356 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=32.845 //y=5.155 //x2=32.235 //y2=5.155
r357 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.15 //y=5.24 //x2=32.15 //y2=5.155
r358 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=32.15 //y=5.24 //x2=32.15 //y2=5.725
r359 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.355 //y=5.155 //x2=31.27 //y2=5.155
r360 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.065 //y=5.155 //x2=32.15 //y2=5.155
r361 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=32.065 //y=5.155 //x2=31.355 //y2=5.155
r362 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.27 //y=5.24 //x2=31.27 //y2=5.155
r363 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.27 //y=5.24 //x2=31.27 //y2=5.725
r364 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.185 //y=5.155 //x2=31.27 //y2=5.155
r365 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=31.185 //y=5.155 //x2=30.475 //y2=5.155
r366 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=30.39 //y=5.24 //x2=30.475 //y2=5.155
r367 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=30.39 //y=5.24 //x2=30.39 //y2=5.725
r368 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=39.59 //y=2.59 //x2=39.59 //y2=2.59
r369 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=34.78 //y=2.59 //x2=34.78 //y2=2.59
r370 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=32.93 //y=2.59 //x2=32.93 //y2=2.59
r371 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.895 //y=2.59 //x2=34.78 //y2=2.59
r372 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=39.475 //y=2.59 //x2=39.59 //y2=2.59
r373 (  3 4 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=39.475 //y=2.59 //x2=34.895 //y2=2.59
r374 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=33.045 //y=2.59 //x2=32.93 //y2=2.59
r375 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=2.59 //x2=34.78 //y2=2.59
r376 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=34.665 //y=2.59 //x2=33.045 //y2=2.59
ends PM_TMRDFFSNRNQNX1\%noxref_9

subckt PM_TMRDFFSNRNQNX1\%noxref_10 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 \
 53 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c169 ( 85 0 ) capacitor c=0.023087f //x=41.625 //y=5.02
c170 ( 84 0 ) capacitor c=0.023519f //x=40.745 //y=5.02
c171 ( 83 0 ) capacitor c=0.0224735f //x=39.865 //y=5.02
c172 ( 81 0 ) capacitor c=0.00853354f //x=41.875 //y=0.915
c173 ( 69 0 ) capacitor c=0.0549166f //x=44.675 //y=4.79
c174 ( 68 0 ) capacitor c=0.0294456f //x=44.965 //y=4.79
c175 ( 67 0 ) capacitor c=0.0347816f //x=44.63 //y=1.22
c176 ( 66 0 ) capacitor c=0.0187487f //x=44.63 //y=0.875
c177 ( 60 0 ) capacitor c=0.0137055f //x=44.475 //y=1.375
c178 ( 58 0 ) capacitor c=0.0149861f //x=44.475 //y=0.72
c179 ( 57 0 ) capacitor c=0.096037f //x=44.1 //y=1.915
c180 ( 56 0 ) capacitor c=0.0228993f //x=44.1 //y=1.53
c181 ( 55 0 ) capacitor c=0.0234352f //x=44.1 //y=1.22
c182 ( 54 0 ) capacitor c=0.0198724f //x=44.1 //y=0.875
c183 ( 53 0 ) capacitor c=0.109949f //x=45.04 //y=6.02
c184 ( 52 0 ) capacitor c=0.158483f //x=44.6 //y=6.02
c185 ( 50 0 ) capacitor c=9.74268e-19 //x=41.77 //y=5.155
c186 ( 49 0 ) capacitor c=0.00191414f //x=40.89 //y=5.155
c187 ( 42 0 ) capacitor c=0.0911502f //x=44.4 //y=2.08
c188 ( 40 0 ) capacitor c=0.103494f //x=42.55 //y=2.59
c189 ( 36 0 ) capacitor c=0.00398962f //x=42.15 //y=1.665
c190 ( 35 0 ) capacitor c=0.0137288f //x=42.465 //y=1.665
c191 ( 29 0 ) capacitor c=0.0276208f //x=42.465 //y=5.155
c192 ( 21 0 ) capacitor c=0.0169868f //x=41.685 //y=5.155
c193 ( 14 0 ) capacitor c=0.00316998f //x=40.095 //y=5.155
c194 ( 13 0 ) capacitor c=0.014258f //x=40.805 //y=5.155
c195 ( 2 0 ) capacitor c=0.00808366f //x=42.665 //y=2.59
c196 ( 1 0 ) capacitor c=0.0351856f //x=44.285 //y=2.59
r197 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=44.965 //y=4.79 //x2=45.04 //y2=4.865
r198 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=44.965 //y=4.79 //x2=44.675 //y2=4.79
r199 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.63 //y=1.22 //x2=44.59 //y2=1.375
r200 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.63 //y=0.875 //x2=44.59 //y2=0.72
r201 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=44.63 //y=0.875 //x2=44.63 //y2=1.22
r202 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=44.6 //y=4.865 //x2=44.675 //y2=4.79
r203 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=44.6 //y=4.865 //x2=44.4 //y2=4.7
r204 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.255 //y=1.375 //x2=44.14 //y2=1.375
r205 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.475 //y=1.375 //x2=44.59 //y2=1.375
r206 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.255 //y=0.72 //x2=44.14 //y2=0.72
r207 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.475 //y=0.72 //x2=44.59 //y2=0.72
r208 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=44.475 //y=0.72 //x2=44.255 //y2=0.72
r209 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=44.1 //y=1.915 //x2=44.4 //y2=2.08
r210 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.1 //y=1.53 //x2=44.14 //y2=1.375
r211 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=44.1 //y=1.53 //x2=44.1 //y2=1.915
r212 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.1 //y=1.22 //x2=44.14 //y2=1.375
r213 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.1 //y=0.875 //x2=44.14 //y2=0.72
r214 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=44.1 //y=0.875 //x2=44.1 //y2=1.22
r215 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.04 //y=6.02 //x2=45.04 //y2=4.865
r216 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=44.6 //y=6.02 //x2=44.6 //y2=4.865
r217 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=44.365 //y=1.375 //x2=44.475 //y2=1.375
r218 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=44.365 //y=1.375 //x2=44.255 //y2=1.375
r219 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=44.4 //y=4.7 //x2=44.4 //y2=4.7
r220 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=44.4 //y=2.59 //x2=44.4 //y2=4.7
r221 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=44.4 //y=2.08 //x2=44.4 //y2=2.08
r222 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=44.4 //y=2.08 //x2=44.4 //y2=2.59
r223 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=42.55 //y=5.07 //x2=42.55 //y2=2.59
r224 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=42.55 //y=1.75 //x2=42.55 //y2=2.59
r225 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.465 //y=1.665 //x2=42.55 //y2=1.75
r226 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=42.465 //y=1.665 //x2=42.15 //y2=1.665
r227 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.065 //y=1.58 //x2=42.15 //y2=1.665
r228 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=42.065 //y=1.58 //x2=42.065 //y2=1.01
r229 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.855 //y=5.155 //x2=41.77 //y2=5.155
r230 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.465 //y=5.155 //x2=42.55 //y2=5.07
r231 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=42.465 //y=5.155 //x2=41.855 //y2=5.155
r232 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.77 //y=5.24 //x2=41.77 //y2=5.155
r233 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=41.77 //y=5.24 //x2=41.77 //y2=5.725
r234 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.975 //y=5.155 //x2=40.89 //y2=5.155
r235 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.685 //y=5.155 //x2=41.77 //y2=5.155
r236 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=41.685 //y=5.155 //x2=40.975 //y2=5.155
r237 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.89 //y=5.24 //x2=40.89 //y2=5.155
r238 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=40.89 //y=5.24 //x2=40.89 //y2=5.725
r239 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.805 //y=5.155 //x2=40.89 //y2=5.155
r240 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=40.805 //y=5.155 //x2=40.095 //y2=5.155
r241 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=40.01 //y=5.24 //x2=40.095 //y2=5.155
r242 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=40.01 //y=5.24 //x2=40.01 //y2=5.725
r243 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=44.4 //y=2.59 //x2=44.4 //y2=2.59
r244 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=42.55 //y=2.59 //x2=42.55 //y2=2.59
r245 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=42.665 //y=2.59 //x2=42.55 //y2=2.59
r246 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=44.285 //y=2.59 //x2=44.4 //y2=2.59
r247 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=44.285 //y=2.59 //x2=42.665 //y2=2.59
ends PM_TMRDFFSNRNQNX1\%noxref_10

subckt PM_TMRDFFSNRNQNX1\%noxref_11 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 \
 63 64 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 90 92 98 99 100 101 106 \
 107 112 123 125 126 127 )
c281 ( 127 0 ) capacitor c=0.023087f //x=36.815 //y=5.02
c282 ( 126 0 ) capacitor c=0.023519f //x=35.935 //y=5.02
c283 ( 125 0 ) capacitor c=0.0224735f //x=35.055 //y=5.02
c284 ( 123 0 ) capacitor c=0.00853354f //x=37.065 //y=0.915
c285 ( 112 0 ) capacitor c=0.0588394f //x=32.19 //y=4.7
c286 ( 107 0 ) capacitor c=0.0273931f //x=32.19 //y=1.915
c287 ( 106 0 ) capacitor c=0.0456313f //x=32.19 //y=2.08
c288 ( 101 0 ) capacitor c=0.0547611f //x=49.485 //y=4.79
c289 ( 100 0 ) capacitor c=0.0294456f //x=49.775 //y=4.79
c290 ( 99 0 ) capacitor c=0.0347816f //x=49.44 //y=1.22
c291 ( 98 0 ) capacitor c=0.0187487f //x=49.44 //y=0.875
c292 ( 92 0 ) capacitor c=0.0137055f //x=49.285 //y=1.375
c293 ( 90 0 ) capacitor c=0.0149861f //x=49.285 //y=0.72
c294 ( 89 0 ) capacitor c=0.096037f //x=48.91 //y=1.915
c295 ( 88 0 ) capacitor c=0.0228993f //x=48.91 //y=1.53
c296 ( 87 0 ) capacitor c=0.0234352f //x=48.91 //y=1.22
c297 ( 86 0 ) capacitor c=0.0198724f //x=48.91 //y=0.875
c298 ( 85 0 ) capacitor c=0.0432517f //x=32.71 //y=1.26
c299 ( 84 0 ) capacitor c=0.0200379f //x=32.71 //y=0.915
c300 ( 81 0 ) capacitor c=0.0148873f //x=32.555 //y=1.415
c301 ( 79 0 ) capacitor c=0.0157803f //x=32.555 //y=0.76
c302 ( 74 0 ) capacitor c=0.0218028f //x=32.18 //y=1.57
c303 ( 73 0 ) capacitor c=0.0207459f //x=32.18 //y=1.26
c304 ( 72 0 ) capacitor c=0.0194308f //x=32.18 //y=0.915
c305 ( 68 0 ) capacitor c=0.109949f //x=49.85 //y=6.02
c306 ( 67 0 ) capacitor c=0.158483f //x=49.41 //y=6.02
c307 ( 66 0 ) capacitor c=0.158754f //x=32.37 //y=6.02
c308 ( 65 0 ) capacitor c=0.109949f //x=31.93 //y=6.02
c309 ( 62 0 ) capacitor c=9.74268e-19 //x=36.96 //y=5.155
c310 ( 61 0 ) capacitor c=0.00191414f //x=36.08 //y=5.155
c311 ( 54 0 ) capacitor c=0.0937531f //x=49.21 //y=2.08
c312 ( 52 0 ) capacitor c=0.103032f //x=37.74 //y=3.33
c313 ( 48 0 ) capacitor c=0.00398962f //x=37.34 //y=1.665
c314 ( 47 0 ) capacitor c=0.0137288f //x=37.655 //y=1.665
c315 ( 41 0 ) capacitor c=0.0276208f //x=37.655 //y=5.155
c316 ( 33 0 ) capacitor c=0.0169868f //x=36.875 //y=5.155
c317 ( 26 0 ) capacitor c=0.00316998f //x=35.285 //y=5.155
c318 ( 25 0 ) capacitor c=0.014258f //x=35.995 //y=5.155
c319 ( 12 0 ) capacitor c=0.0816952f //x=32.19 //y=2.08
c320 ( 4 0 ) capacitor c=0.00551333f //x=37.855 //y=3.33
c321 ( 3 0 ) capacitor c=0.173933f //x=49.095 //y=3.33
c322 ( 2 0 ) capacitor c=0.0108616f //x=32.305 //y=3.33
c323 ( 1 0 ) capacitor c=0.0905825f //x=37.625 //y=3.33
r324 (  106 107 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=32.19 //y=2.08 //x2=32.19 //y2=1.915
r325 (  100 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=49.775 //y=4.79 //x2=49.85 //y2=4.865
r326 (  100 101 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=49.775 //y=4.79 //x2=49.485 //y2=4.79
r327 (  99 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.44 //y=1.22 //x2=49.4 //y2=1.375
r328 (  98 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.44 //y=0.875 //x2=49.4 //y2=0.72
r329 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=49.44 //y=0.875 //x2=49.44 //y2=1.22
r330 (  95 101 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=49.41 //y=4.865 //x2=49.485 //y2=4.79
r331 (  95 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=49.41 //y=4.865 //x2=49.21 //y2=4.7
r332 (  93 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.065 //y=1.375 //x2=48.95 //y2=1.375
r333 (  92 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.285 //y=1.375 //x2=49.4 //y2=1.375
r334 (  91 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.065 //y=0.72 //x2=48.95 //y2=0.72
r335 (  90 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.285 //y=0.72 //x2=49.4 //y2=0.72
r336 (  90 91 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=49.285 //y=0.72 //x2=49.065 //y2=0.72
r337 (  89 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.915 //x2=49.21 //y2=2.08
r338 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.53 //x2=48.95 //y2=1.375
r339 (  88 89 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.53 //x2=48.91 //y2=1.915
r340 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.22 //x2=48.95 //y2=1.375
r341 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=48.91 //y=0.875 //x2=48.95 //y2=0.72
r342 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=48.91 //y=0.875 //x2=48.91 //y2=1.22
r343 (  85 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.71 //y=1.26 //x2=32.67 //y2=1.415
r344 (  84 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.71 //y=0.915 //x2=32.67 //y2=0.76
r345 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=32.71 //y=0.915 //x2=32.71 //y2=1.26
r346 (  82 110 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.335 //y=1.415 //x2=32.22 //y2=1.415
r347 (  81 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.555 //y=1.415 //x2=32.67 //y2=1.415
r348 (  80 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.335 //y=0.76 //x2=32.22 //y2=0.76
r349 (  79 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.555 //y=0.76 //x2=32.67 //y2=0.76
r350 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=32.555 //y=0.76 //x2=32.335 //y2=0.76
r351 (  76 112 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=32.37 //y=4.865 //x2=32.19 //y2=4.7
r352 (  74 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.18 //y=1.57 //x2=32.22 //y2=1.415
r353 (  74 107 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=32.18 //y=1.57 //x2=32.18 //y2=1.915
r354 (  73 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.18 //y=1.26 //x2=32.22 //y2=1.415
r355 (  72 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.18 //y=0.915 //x2=32.22 //y2=0.76
r356 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=32.18 //y=0.915 //x2=32.18 //y2=1.26
r357 (  69 112 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=31.93 //y=4.865 //x2=32.19 //y2=4.7
r358 (  68 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.85 //y=6.02 //x2=49.85 //y2=4.865
r359 (  67 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.41 //y=6.02 //x2=49.41 //y2=4.865
r360 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=32.37 //y=6.02 //x2=32.37 //y2=4.865
r361 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.93 //y=6.02 //x2=31.93 //y2=4.865
r362 (  64 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=49.175 //y=1.375 //x2=49.285 //y2=1.375
r363 (  64 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=49.175 //y=1.375 //x2=49.065 //y2=1.375
r364 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=32.445 //y=1.415 //x2=32.555 //y2=1.415
r365 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=32.445 //y=1.415 //x2=32.335 //y2=1.415
r366 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.21 //y=4.7 //x2=49.21 //y2=4.7
r367 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=49.21 //y=3.33 //x2=49.21 //y2=4.7
r368 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.21 //y=2.08 //x2=49.21 //y2=2.08
r369 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=49.21 //y=2.08 //x2=49.21 //y2=3.33
r370 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=37.74 //y=5.07 //x2=37.74 //y2=3.33
r371 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=37.74 //y=1.75 //x2=37.74 //y2=3.33
r372 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.655 //y=1.665 //x2=37.74 //y2=1.75
r373 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=37.655 //y=1.665 //x2=37.34 //y2=1.665
r374 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.255 //y=1.58 //x2=37.34 //y2=1.665
r375 (  43 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=37.255 //y=1.58 //x2=37.255 //y2=1.01
r376 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.045 //y=5.155 //x2=36.96 //y2=5.155
r377 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.655 //y=5.155 //x2=37.74 //y2=5.07
r378 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=37.655 //y=5.155 //x2=37.045 //y2=5.155
r379 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.96 //y=5.24 //x2=36.96 //y2=5.155
r380 (  35 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=36.96 //y=5.24 //x2=36.96 //y2=5.725
r381 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.165 //y=5.155 //x2=36.08 //y2=5.155
r382 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.875 //y=5.155 //x2=36.96 //y2=5.155
r383 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=36.875 //y=5.155 //x2=36.165 //y2=5.155
r384 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.08 //y=5.24 //x2=36.08 //y2=5.155
r385 (  27 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=36.08 //y=5.24 //x2=36.08 //y2=5.725
r386 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.995 //y=5.155 //x2=36.08 //y2=5.155
r387 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=35.995 //y=5.155 //x2=35.285 //y2=5.155
r388 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=35.2 //y=5.24 //x2=35.285 //y2=5.155
r389 (  19 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.2 //y=5.24 //x2=35.2 //y2=5.725
r390 (  17 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=32.19 //y=4.7 //x2=32.19 //y2=4.7
r391 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=32.19 //y=3.33 //x2=32.19 //y2=4.7
r392 (  12 106 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=32.19 //y=2.08 //x2=32.19 //y2=2.08
r393 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=32.19 //y=2.08 //x2=32.19 //y2=3.33
r394 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=49.21 //y=3.33 //x2=49.21 //y2=3.33
r395 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=37.74 //y=3.33 //x2=37.74 //y2=3.33
r396 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=32.19 //y=3.33 //x2=32.19 //y2=3.33
r397 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.855 //y=3.33 //x2=37.74 //y2=3.33
r398 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=49.095 //y=3.33 //x2=49.21 //y2=3.33
r399 (  3 4 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=49.095 //y=3.33 //x2=37.855 //y2=3.33
r400 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=32.305 //y=3.33 //x2=32.19 //y2=3.33
r401 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.625 //y=3.33 //x2=37.74 //y2=3.33
r402 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=37.625 //y=3.33 //x2=32.305 //y2=3.33
ends PM_TMRDFFSNRNQNX1\%noxref_11

subckt PM_TMRDFFSNRNQNX1\%noxref_12 ( 1 2 3 4 5 6 16 24 37 38 45 53 59 60 64 \
 66 73 74 75 76 77 78 79 80 81 82 83 87 88 89 94 96 99 100 104 105 106 111 113 \
 116 117 121 122 123 128 130 133 134 136 137 142 146 147 152 156 157 162 165 \
 167 168 169 )
c354 ( 169 0 ) capacitor c=0.023087f //x=46.435 //y=5.02
c355 ( 168 0 ) capacitor c=0.023519f //x=45.555 //y=5.02
c356 ( 167 0 ) capacitor c=0.0224735f //x=44.675 //y=5.02
c357 ( 165 0 ) capacitor c=0.00853354f //x=46.685 //y=0.915
c358 ( 162 0 ) capacitor c=0.0588394f //x=56.24 //y=4.7
c359 ( 157 0 ) capacitor c=0.0273931f //x=56.24 //y=1.915
c360 ( 156 0 ) capacitor c=0.0456313f //x=56.24 //y=2.08
c361 ( 152 0 ) capacitor c=0.0588394f //x=41.81 //y=4.7
c362 ( 147 0 ) capacitor c=0.0273931f //x=41.81 //y=1.915
c363 ( 146 0 ) capacitor c=0.0456313f //x=41.81 //y=2.08
c364 ( 142 0 ) capacitor c=0.0589949f //x=37 //y=4.7
c365 ( 137 0 ) capacitor c=0.0273931f //x=37 //y=1.915
c366 ( 136 0 ) capacitor c=0.0456313f //x=37 //y=2.08
c367 ( 134 0 ) capacitor c=0.0432517f //x=56.76 //y=1.26
c368 ( 133 0 ) capacitor c=0.0200379f //x=56.76 //y=0.915
c369 ( 130 0 ) capacitor c=0.0148873f //x=56.605 //y=1.415
c370 ( 128 0 ) capacitor c=0.0157803f //x=56.605 //y=0.76
c371 ( 123 0 ) capacitor c=0.0218028f //x=56.23 //y=1.57
c372 ( 122 0 ) capacitor c=0.0207459f //x=56.23 //y=1.26
c373 ( 121 0 ) capacitor c=0.0194308f //x=56.23 //y=0.915
c374 ( 117 0 ) capacitor c=0.0432517f //x=42.33 //y=1.26
c375 ( 116 0 ) capacitor c=0.0200379f //x=42.33 //y=0.915
c376 ( 113 0 ) capacitor c=0.0148873f //x=42.175 //y=1.415
c377 ( 111 0 ) capacitor c=0.0157803f //x=42.175 //y=0.76
c378 ( 106 0 ) capacitor c=0.0218028f //x=41.8 //y=1.57
c379 ( 105 0 ) capacitor c=0.0207459f //x=41.8 //y=1.26
c380 ( 104 0 ) capacitor c=0.0194308f //x=41.8 //y=0.915
c381 ( 100 0 ) capacitor c=0.0432517f //x=37.52 //y=1.26
c382 ( 99 0 ) capacitor c=0.0200379f //x=37.52 //y=0.915
c383 ( 96 0 ) capacitor c=0.0148873f //x=37.365 //y=1.415
c384 ( 94 0 ) capacitor c=0.0157803f //x=37.365 //y=0.76
c385 ( 89 0 ) capacitor c=0.0218028f //x=36.99 //y=1.57
c386 ( 88 0 ) capacitor c=0.0207459f //x=36.99 //y=1.26
c387 ( 87 0 ) capacitor c=0.0194308f //x=36.99 //y=0.915
c388 ( 83 0 ) capacitor c=0.158754f //x=56.42 //y=6.02
c389 ( 82 0 ) capacitor c=0.109949f //x=55.98 //y=6.02
c390 ( 81 0 ) capacitor c=0.158754f //x=41.99 //y=6.02
c391 ( 80 0 ) capacitor c=0.109949f //x=41.55 //y=6.02
c392 ( 79 0 ) capacitor c=0.158754f //x=37.18 //y=6.02
c393 ( 78 0 ) capacitor c=0.109949f //x=36.74 //y=6.02
c394 ( 74 0 ) capacitor c=9.74268e-19 //x=46.58 //y=5.155
c395 ( 73 0 ) capacitor c=0.00191414f //x=45.7 //y=5.155
c396 ( 66 0 ) capacitor c=0.0770908f //x=56.24 //y=2.08
c397 ( 64 0 ) capacitor c=0.104892f //x=47.36 //y=3.7
c398 ( 60 0 ) capacitor c=0.00398962f //x=46.96 //y=1.665
c399 ( 59 0 ) capacitor c=0.0137288f //x=47.275 //y=1.665
c400 ( 53 0 ) capacitor c=0.0276208f //x=47.275 //y=5.155
c401 ( 45 0 ) capacitor c=0.0169868f //x=46.495 //y=5.155
c402 ( 38 0 ) capacitor c=0.00316998f //x=44.905 //y=5.155
c403 ( 37 0 ) capacitor c=0.014258f //x=45.615 //y=5.155
c404 ( 24 0 ) capacitor c=0.0790362f //x=41.81 //y=2.08
c405 ( 16 0 ) capacitor c=0.0776243f //x=37 //y=2.08
c406 ( 6 0 ) capacitor c=0.0055354f //x=47.475 //y=3.7
c407 ( 5 0 ) capacitor c=0.140148f //x=56.125 //y=3.7
c408 ( 4 0 ) capacitor c=0.00533183f //x=41.925 //y=3.7
c409 ( 3 0 ) capacitor c=0.0751185f //x=47.245 //y=3.7
c410 ( 2 0 ) capacitor c=0.01364f //x=37.115 //y=3.7
c411 ( 1 0 ) capacitor c=0.0665749f //x=41.695 //y=3.7
r412 (  156 157 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=56.24 //y=2.08 //x2=56.24 //y2=1.915
r413 (  146 147 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=41.81 //y=2.08 //x2=41.81 //y2=1.915
r414 (  136 137 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=37 //y=2.08 //x2=37 //y2=1.915
r415 (  134 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.76 //y=1.26 //x2=56.72 //y2=1.415
r416 (  133 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.76 //y=0.915 //x2=56.72 //y2=0.76
r417 (  133 134 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.76 //y=0.915 //x2=56.76 //y2=1.26
r418 (  131 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.385 //y=1.415 //x2=56.27 //y2=1.415
r419 (  130 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.605 //y=1.415 //x2=56.72 //y2=1.415
r420 (  129 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.385 //y=0.76 //x2=56.27 //y2=0.76
r421 (  128 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.605 //y=0.76 //x2=56.72 //y2=0.76
r422 (  128 129 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=56.605 //y=0.76 //x2=56.385 //y2=0.76
r423 (  125 162 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=56.42 //y=4.865 //x2=56.24 //y2=4.7
r424 (  123 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.23 //y=1.57 //x2=56.27 //y2=1.415
r425 (  123 157 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.23 //y=1.57 //x2=56.23 //y2=1.915
r426 (  122 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.23 //y=1.26 //x2=56.27 //y2=1.415
r427 (  121 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.23 //y=0.915 //x2=56.27 //y2=0.76
r428 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.23 //y=0.915 //x2=56.23 //y2=1.26
r429 (  118 162 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=55.98 //y=4.865 //x2=56.24 //y2=4.7
r430 (  117 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.33 //y=1.26 //x2=42.29 //y2=1.415
r431 (  116 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.33 //y=0.915 //x2=42.29 //y2=0.76
r432 (  116 117 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.33 //y=0.915 //x2=42.33 //y2=1.26
r433 (  114 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.955 //y=1.415 //x2=41.84 //y2=1.415
r434 (  113 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.175 //y=1.415 //x2=42.29 //y2=1.415
r435 (  112 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.955 //y=0.76 //x2=41.84 //y2=0.76
r436 (  111 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.175 //y=0.76 //x2=42.29 //y2=0.76
r437 (  111 112 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=42.175 //y=0.76 //x2=41.955 //y2=0.76
r438 (  108 152 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=41.99 //y=4.865 //x2=41.81 //y2=4.7
r439 (  106 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.8 //y=1.57 //x2=41.84 //y2=1.415
r440 (  106 147 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=41.8 //y=1.57 //x2=41.8 //y2=1.915
r441 (  105 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.8 //y=1.26 //x2=41.84 //y2=1.415
r442 (  104 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.8 //y=0.915 //x2=41.84 //y2=0.76
r443 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=41.8 //y=0.915 //x2=41.8 //y2=1.26
r444 (  101 152 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=41.55 //y=4.865 //x2=41.81 //y2=4.7
r445 (  100 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.52 //y=1.26 //x2=37.48 //y2=1.415
r446 (  99 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.52 //y=0.915 //x2=37.48 //y2=0.76
r447 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=37.52 //y=0.915 //x2=37.52 //y2=1.26
r448 (  97 140 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.145 //y=1.415 //x2=37.03 //y2=1.415
r449 (  96 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.365 //y=1.415 //x2=37.48 //y2=1.415
r450 (  95 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.145 //y=0.76 //x2=37.03 //y2=0.76
r451 (  94 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.365 //y=0.76 //x2=37.48 //y2=0.76
r452 (  94 95 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=37.365 //y=0.76 //x2=37.145 //y2=0.76
r453 (  91 142 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=37.18 //y=4.865 //x2=37 //y2=4.7
r454 (  89 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.99 //y=1.57 //x2=37.03 //y2=1.415
r455 (  89 137 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=36.99 //y=1.57 //x2=36.99 //y2=1.915
r456 (  88 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.99 //y=1.26 //x2=37.03 //y2=1.415
r457 (  87 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.99 //y=0.915 //x2=37.03 //y2=0.76
r458 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=36.99 //y=0.915 //x2=36.99 //y2=1.26
r459 (  84 142 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=36.74 //y=4.865 //x2=37 //y2=4.7
r460 (  83 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=56.42 //y=6.02 //x2=56.42 //y2=4.865
r461 (  82 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.98 //y=6.02 //x2=55.98 //y2=4.865
r462 (  81 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.99 //y=6.02 //x2=41.99 //y2=4.865
r463 (  80 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.55 //y=6.02 //x2=41.55 //y2=4.865
r464 (  79 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=37.18 //y=6.02 //x2=37.18 //y2=4.865
r465 (  78 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=36.74 //y=6.02 //x2=36.74 //y2=4.865
r466 (  77 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=56.495 //y=1.415 //x2=56.605 //y2=1.415
r467 (  77 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=56.495 //y=1.415 //x2=56.385 //y2=1.415
r468 (  76 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.065 //y=1.415 //x2=42.175 //y2=1.415
r469 (  76 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.065 //y=1.415 //x2=41.955 //y2=1.415
r470 (  75 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.255 //y=1.415 //x2=37.365 //y2=1.415
r471 (  75 97 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.255 //y=1.415 //x2=37.145 //y2=1.415
r472 (  71 162 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=56.24 //y=4.7 //x2=56.24 //y2=4.7
r473 (  69 71 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=56.24 //y=3.7 //x2=56.24 //y2=4.7
r474 (  66 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=56.24 //y=2.08 //x2=56.24 //y2=2.08
r475 (  66 69 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=56.24 //y=2.08 //x2=56.24 //y2=3.7
r476 (  62 64 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=47.36 //y=5.07 //x2=47.36 //y2=3.7
r477 (  61 64 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=47.36 //y=1.75 //x2=47.36 //y2=3.7
r478 (  59 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=47.275 //y=1.665 //x2=47.36 //y2=1.75
r479 (  59 60 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=47.275 //y=1.665 //x2=46.96 //y2=1.665
r480 (  55 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=46.875 //y=1.58 //x2=46.96 //y2=1.665
r481 (  55 165 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=46.875 //y=1.58 //x2=46.875 //y2=1.01
r482 (  54 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.665 //y=5.155 //x2=46.58 //y2=5.155
r483 (  53 62 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=47.275 //y=5.155 //x2=47.36 //y2=5.07
r484 (  53 54 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=47.275 //y=5.155 //x2=46.665 //y2=5.155
r485 (  47 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.58 //y=5.24 //x2=46.58 //y2=5.155
r486 (  47 169 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.58 //y=5.24 //x2=46.58 //y2=5.725
r487 (  46 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.785 //y=5.155 //x2=45.7 //y2=5.155
r488 (  45 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.495 //y=5.155 //x2=46.58 //y2=5.155
r489 (  45 46 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.495 //y=5.155 //x2=45.785 //y2=5.155
r490 (  39 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.7 //y=5.24 //x2=45.7 //y2=5.155
r491 (  39 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.7 //y=5.24 //x2=45.7 //y2=5.725
r492 (  37 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.615 //y=5.155 //x2=45.7 //y2=5.155
r493 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=45.615 //y=5.155 //x2=44.905 //y2=5.155
r494 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=44.82 //y=5.24 //x2=44.905 //y2=5.155
r495 (  31 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=44.82 //y=5.24 //x2=44.82 //y2=5.725
r496 (  29 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.81 //y=4.7 //x2=41.81 //y2=4.7
r497 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=41.81 //y=3.7 //x2=41.81 //y2=4.7
r498 (  24 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.81 //y=2.08 //x2=41.81 //y2=2.08
r499 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=41.81 //y=2.08 //x2=41.81 //y2=3.7
r500 (  21 142 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37 //y=4.7 //x2=37 //y2=4.7
r501 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=37 //y=3.7 //x2=37 //y2=4.7
r502 (  16 136 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37 //y=2.08 //x2=37 //y2=2.08
r503 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=37 //y=2.08 //x2=37 //y2=3.7
r504 (  14 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=56.24 //y=3.7 //x2=56.24 //y2=3.7
r505 (  12 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=47.36 //y=3.7 //x2=47.36 //y2=3.7
r506 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=41.81 //y=3.7 //x2=41.81 //y2=3.7
r507 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=37 \
 //y=3.7 //x2=37 //y2=3.7
r508 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.475 //y=3.7 //x2=47.36 //y2=3.7
r509 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.125 //y=3.7 //x2=56.24 //y2=3.7
r510 (  5 6 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=56.125 //y=3.7 //x2=47.475 //y2=3.7
r511 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=41.925 //y=3.7 //x2=41.81 //y2=3.7
r512 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.245 //y=3.7 //x2=47.36 //y2=3.7
r513 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=47.245 //y=3.7 //x2=41.925 //y2=3.7
r514 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.115 //y=3.7 //x2=37 //y2=3.7
r515 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=41.695 //y=3.7 //x2=41.81 //y2=3.7
r516 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=41.695 //y=3.7 //x2=37.115 //y2=3.7
ends PM_TMRDFFSNRNQNX1\%noxref_12

subckt PM_TMRDFFSNRNQNX1\%noxref_13 ( 1 2 8 21 22 29 37 43 44 48 49 50 51 52 \
 53 57 58 59 64 66 69 70 72 73 78 81 83 84 85 )
c178 ( 85 0 ) capacitor c=0.023087f //x=56.055 //y=5.02
c179 ( 84 0 ) capacitor c=0.023519f //x=55.175 //y=5.02
c180 ( 83 0 ) capacitor c=0.0224735f //x=54.295 //y=5.02
c181 ( 81 0 ) capacitor c=0.00853354f //x=56.305 //y=0.915
c182 ( 78 0 ) capacitor c=0.0588394f //x=51.43 //y=4.7
c183 ( 73 0 ) capacitor c=0.0273931f //x=51.43 //y=1.915
c184 ( 72 0 ) capacitor c=0.0456313f //x=51.43 //y=2.08
c185 ( 70 0 ) capacitor c=0.0432517f //x=51.95 //y=1.26
c186 ( 69 0 ) capacitor c=0.0200379f //x=51.95 //y=0.915
c187 ( 66 0 ) capacitor c=0.0148873f //x=51.795 //y=1.415
c188 ( 64 0 ) capacitor c=0.0157803f //x=51.795 //y=0.76
c189 ( 59 0 ) capacitor c=0.0218028f //x=51.42 //y=1.57
c190 ( 58 0 ) capacitor c=0.0207459f //x=51.42 //y=1.26
c191 ( 57 0 ) capacitor c=0.0194308f //x=51.42 //y=0.915
c192 ( 53 0 ) capacitor c=0.158754f //x=51.61 //y=6.02
c193 ( 52 0 ) capacitor c=0.109949f //x=51.17 //y=6.02
c194 ( 50 0 ) capacitor c=9.74268e-19 //x=56.2 //y=5.155
c195 ( 49 0 ) capacitor c=0.00191414f //x=55.32 //y=5.155
c196 ( 48 0 ) capacitor c=0.0997105f //x=56.98 //y=2.59
c197 ( 44 0 ) capacitor c=0.00398962f //x=56.58 //y=1.665
c198 ( 43 0 ) capacitor c=0.0137288f //x=56.895 //y=1.665
c199 ( 37 0 ) capacitor c=0.0276208f //x=56.895 //y=5.155
c200 ( 29 0 ) capacitor c=0.0169868f //x=56.115 //y=5.155
c201 ( 22 0 ) capacitor c=0.00316998f //x=54.525 //y=5.155
c202 ( 21 0 ) capacitor c=0.014258f //x=55.235 //y=5.155
c203 ( 8 0 ) capacitor c=0.0791424f //x=51.43 //y=2.08
c204 ( 2 0 ) capacitor c=0.0137813f //x=51.545 //y=2.59
c205 ( 1 0 ) capacitor c=0.0833895f //x=56.865 //y=2.59
r206 (  72 73 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=51.43 //y=2.08 //x2=51.43 //y2=1.915
r207 (  70 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.95 //y=1.26 //x2=51.91 //y2=1.415
r208 (  69 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.95 //y=0.915 //x2=51.91 //y2=0.76
r209 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=51.95 //y=0.915 //x2=51.95 //y2=1.26
r210 (  67 76 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.575 //y=1.415 //x2=51.46 //y2=1.415
r211 (  66 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.795 //y=1.415 //x2=51.91 //y2=1.415
r212 (  65 75 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.575 //y=0.76 //x2=51.46 //y2=0.76
r213 (  64 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.795 //y=0.76 //x2=51.91 //y2=0.76
r214 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=51.795 //y=0.76 //x2=51.575 //y2=0.76
r215 (  61 78 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=51.61 //y=4.865 //x2=51.43 //y2=4.7
r216 (  59 76 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.42 //y=1.57 //x2=51.46 //y2=1.415
r217 (  59 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=51.42 //y=1.57 //x2=51.42 //y2=1.915
r218 (  58 76 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.42 //y=1.26 //x2=51.46 //y2=1.415
r219 (  57 75 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.42 //y=0.915 //x2=51.46 //y2=0.76
r220 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=51.42 //y=0.915 //x2=51.42 //y2=1.26
r221 (  54 78 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=51.17 //y=4.865 //x2=51.43 //y2=4.7
r222 (  53 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=51.61 //y=6.02 //x2=51.61 //y2=4.865
r223 (  52 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=51.17 //y=6.02 //x2=51.17 //y2=4.865
r224 (  51 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=51.685 //y=1.415 //x2=51.795 //y2=1.415
r225 (  51 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=51.685 //y=1.415 //x2=51.575 //y2=1.415
r226 (  46 48 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=56.98 //y=5.07 //x2=56.98 //y2=2.59
r227 (  45 48 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=56.98 //y=1.75 //x2=56.98 //y2=2.59
r228 (  43 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.895 //y=1.665 //x2=56.98 //y2=1.75
r229 (  43 44 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=56.895 //y=1.665 //x2=56.58 //y2=1.665
r230 (  39 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.495 //y=1.58 //x2=56.58 //y2=1.665
r231 (  39 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=56.495 //y=1.58 //x2=56.495 //y2=1.01
r232 (  38 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.285 //y=5.155 //x2=56.2 //y2=5.155
r233 (  37 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.895 //y=5.155 //x2=56.98 //y2=5.07
r234 (  37 38 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=56.895 //y=5.155 //x2=56.285 //y2=5.155
r235 (  31 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.2 //y=5.24 //x2=56.2 //y2=5.155
r236 (  31 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=56.2 //y=5.24 //x2=56.2 //y2=5.725
r237 (  30 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.405 //y=5.155 //x2=55.32 //y2=5.155
r238 (  29 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.115 //y=5.155 //x2=56.2 //y2=5.155
r239 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=56.115 //y=5.155 //x2=55.405 //y2=5.155
r240 (  23 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.32 //y=5.24 //x2=55.32 //y2=5.155
r241 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.32 //y=5.24 //x2=55.32 //y2=5.725
r242 (  21 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.235 //y=5.155 //x2=55.32 //y2=5.155
r243 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=55.235 //y=5.155 //x2=54.525 //y2=5.155
r244 (  15 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=54.44 //y=5.24 //x2=54.525 //y2=5.155
r245 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.44 //y=5.24 //x2=54.44 //y2=5.725
r246 (  13 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=51.43 //y=4.7 //x2=51.43 //y2=4.7
r247 (  11 13 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=51.43 //y=2.59 //x2=51.43 //y2=4.7
r248 (  8 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=51.43 //y=2.08 //x2=51.43 //y2=2.08
r249 (  8 11 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=51.43 //y=2.08 //x2=51.43 //y2=2.59
r250 (  6 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=56.98 //y=2.59 //x2=56.98 //y2=2.59
r251 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=51.43 //y=2.59 //x2=51.43 //y2=2.59
r252 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=51.545 //y=2.59 //x2=51.43 //y2=2.59
r253 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.865 //y=2.59 //x2=56.98 //y2=2.59
r254 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=56.865 //y=2.59 //x2=51.545 //y2=2.59
ends PM_TMRDFFSNRNQNX1\%noxref_13

subckt PM_TMRDFFSNRNQNX1\%D ( 1 2 3 4 11 12 13 14 15 16 17 18 19 20 21 22 23 \
 24 26 40 51 60 61 62 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 \
 91 92 94 100 101 102 103 107 108 109 110 111 113 119 120 121 122 )
c342 ( 122 0 ) capacitor c=0.0547611f //x=59.105 //y=4.79
c343 ( 121 0 ) capacitor c=0.0294456f //x=59.395 //y=4.79
c344 ( 120 0 ) capacitor c=0.0347816f //x=59.06 //y=1.22
c345 ( 119 0 ) capacitor c=0.0187487f //x=59.06 //y=0.875
c346 ( 113 0 ) capacitor c=0.0137055f //x=58.905 //y=1.375
c347 ( 111 0 ) capacitor c=0.0149861f //x=58.905 //y=0.72
c348 ( 110 0 ) capacitor c=0.096037f //x=58.53 //y=1.915
c349 ( 109 0 ) capacitor c=0.0228993f //x=58.53 //y=1.53
c350 ( 108 0 ) capacitor c=0.0234352f //x=58.53 //y=1.22
c351 ( 107 0 ) capacitor c=0.0198724f //x=58.53 //y=0.875
c352 ( 103 0 ) capacitor c=0.0547611f //x=30.245 //y=4.79
c353 ( 102 0 ) capacitor c=0.0294456f //x=30.535 //y=4.79
c354 ( 101 0 ) capacitor c=0.0347816f //x=30.2 //y=1.22
c355 ( 100 0 ) capacitor c=0.0187487f //x=30.2 //y=0.875
c356 ( 94 0 ) capacitor c=0.0137055f //x=30.045 //y=1.375
c357 ( 92 0 ) capacitor c=0.0149861f //x=30.045 //y=0.72
c358 ( 91 0 ) capacitor c=0.096037f //x=29.67 //y=1.915
c359 ( 90 0 ) capacitor c=0.0228993f //x=29.67 //y=1.53
c360 ( 89 0 ) capacitor c=0.0234352f //x=29.67 //y=1.22
c361 ( 88 0 ) capacitor c=0.0198724f //x=29.67 //y=0.875
c362 ( 84 0 ) capacitor c=0.0558341f //x=1.385 //y=4.79
c363 ( 83 0 ) capacitor c=0.0298189f //x=1.675 //y=4.79
c364 ( 82 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c365 ( 81 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c366 ( 75 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c367 ( 73 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c368 ( 72 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c369 ( 71 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c370 ( 70 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c371 ( 69 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c372 ( 68 0 ) capacitor c=0.109949f //x=59.47 //y=6.02
c373 ( 67 0 ) capacitor c=0.158483f //x=59.03 //y=6.02
c374 ( 66 0 ) capacitor c=0.109949f //x=30.61 //y=6.02
c375 ( 65 0 ) capacitor c=0.158483f //x=30.17 //y=6.02
c376 ( 64 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c377 ( 63 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c378 ( 51 0 ) capacitor c=0.0952756f //x=58.83 //y=2.08
c379 ( 40 0 ) capacitor c=0.0991769f //x=29.97 //y=2.08
c380 ( 26 0 ) capacitor c=0.124371f //x=1.11 //y=2.08
c381 ( 4 0 ) capacitor c=0.00590384f //x=30.085 //y=4.07
c382 ( 3 0 ) capacitor c=0.426491f //x=58.715 //y=4.07
c383 ( 2 0 ) capacitor c=0.0231516f //x=1.225 //y=4.07
c384 ( 1 0 ) capacitor c=0.511583f //x=29.855 //y=4.07
r385 (  121 123 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=59.395 //y=4.79 //x2=59.47 //y2=4.865
r386 (  121 122 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=59.395 //y=4.79 //x2=59.105 //y2=4.79
r387 (  120 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.06 //y=1.22 //x2=59.02 //y2=1.375
r388 (  119 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.06 //y=0.875 //x2=59.02 //y2=0.72
r389 (  119 120 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=59.06 //y=0.875 //x2=59.06 //y2=1.22
r390 (  116 122 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=59.03 //y=4.865 //x2=59.105 //y2=4.79
r391 (  116 147 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=59.03 //y=4.865 //x2=58.83 //y2=4.7
r392 (  114 143 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.685 //y=1.375 //x2=58.57 //y2=1.375
r393 (  113 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.905 //y=1.375 //x2=59.02 //y2=1.375
r394 (  112 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.685 //y=0.72 //x2=58.57 //y2=0.72
r395 (  111 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.905 //y=0.72 //x2=59.02 //y2=0.72
r396 (  111 112 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=58.905 //y=0.72 //x2=58.685 //y2=0.72
r397 (  110 145 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=58.53 //y=1.915 //x2=58.83 //y2=2.08
r398 (  109 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.53 //y=1.53 //x2=58.57 //y2=1.375
r399 (  109 110 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=58.53 //y=1.53 //x2=58.53 //y2=1.915
r400 (  108 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.53 //y=1.22 //x2=58.57 //y2=1.375
r401 (  107 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.53 //y=0.875 //x2=58.57 //y2=0.72
r402 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=58.53 //y=0.875 //x2=58.53 //y2=1.22
r403 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=30.535 //y=4.79 //x2=30.61 //y2=4.865
r404 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=30.535 //y=4.79 //x2=30.245 //y2=4.79
r405 (  101 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.2 //y=1.22 //x2=30.16 //y2=1.375
r406 (  100 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.2 //y=0.875 //x2=30.16 //y2=0.72
r407 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=30.2 //y=0.875 //x2=30.2 //y2=1.22
r408 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=30.17 //y=4.865 //x2=30.245 //y2=4.79
r409 (  97 139 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=30.17 //y=4.865 //x2=29.97 //y2=4.7
r410 (  95 135 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.825 //y=1.375 //x2=29.71 //y2=1.375
r411 (  94 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.045 //y=1.375 //x2=30.16 //y2=1.375
r412 (  93 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.825 //y=0.72 //x2=29.71 //y2=0.72
r413 (  92 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.045 //y=0.72 //x2=30.16 //y2=0.72
r414 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=30.045 //y=0.72 //x2=29.825 //y2=0.72
r415 (  91 137 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=29.67 //y=1.915 //x2=29.97 //y2=2.08
r416 (  90 135 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.67 //y=1.53 //x2=29.71 //y2=1.375
r417 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=29.67 //y=1.53 //x2=29.67 //y2=1.915
r418 (  89 135 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.67 //y=1.22 //x2=29.71 //y2=1.375
r419 (  88 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.67 //y=0.875 //x2=29.71 //y2=0.72
r420 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=29.67 //y=0.875 //x2=29.67 //y2=1.22
r421 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r422 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r423 (  82 133 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r424 (  81 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r425 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r426 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r427 (  78 131 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r428 (  76 127 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r429 (  75 133 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r430 (  74 126 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r431 (  73 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r432 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r433 (  72 129 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r434 (  71 127 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r435 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r436 (  70 127 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r437 (  69 126 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r438 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r439 (  68 123 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.47 //y=6.02 //x2=59.47 //y2=4.865
r440 (  67 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.03 //y=6.02 //x2=59.03 //y2=4.865
r441 (  66 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.61 //y=6.02 //x2=30.61 //y2=4.865
r442 (  65 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.17 //y=6.02 //x2=30.17 //y2=4.865
r443 (  64 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r444 (  63 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r445 (  62 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.795 //y=1.375 //x2=58.905 //y2=1.375
r446 (  62 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.795 //y=1.375 //x2=58.685 //y2=1.375
r447 (  61 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=29.935 //y=1.375 //x2=30.045 //y2=1.375
r448 (  61 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=29.935 //y=1.375 //x2=29.825 //y2=1.375
r449 (  60 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r450 (  60 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r451 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.83 //y=4.7 //x2=58.83 //y2=4.7
r452 (  51 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.83 //y=2.08 //x2=58.83 //y2=2.08
r453 (  48 139 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.97 //y=4.7 //x2=29.97 //y2=4.7
r454 (  40 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.97 //y=2.08 //x2=29.97 //y2=2.08
r455 (  37 131 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r456 (  26 129 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r457 (  24 58 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=58.83 //y=4.07 //x2=58.83 //y2=4.7
r458 (  23 24 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=58.83 //y=3.33 //x2=58.83 //y2=4.07
r459 (  22 23 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=58.83 //y=2.59 //x2=58.83 //y2=3.33
r460 (  22 51 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=58.83 //y=2.59 //x2=58.83 //y2=2.08
r461 (  21 48 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=29.97 //y=4.07 //x2=29.97 //y2=4.7
r462 (  20 21 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=29.97 //y=3.7 //x2=29.97 //y2=4.07
r463 (  19 20 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=29.97 //y=3.33 //x2=29.97 //y2=3.7
r464 (  18 19 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=29.97 //y=2.59 //x2=29.97 //y2=3.33
r465 (  18 40 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=29.97 //y=2.59 //x2=29.97 //y2=2.08
r466 (  17 37 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.44 //x2=1.11 //y2=4.7
r467 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r468 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r469 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r470 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r471 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r472 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.22 //x2=1.11 //y2=2.59
r473 (  11 26 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.22 //x2=1.11 //y2=2.08
r474 (  10 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=58.83 //y=4.07 //x2=58.83 //y2=4.07
r475 (  8 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=29.97 //y=4.07 //x2=29.97 //y2=4.07
r476 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.07
r477 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=30.085 //y=4.07 //x2=29.97 //y2=4.07
r478 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=58.715 //y=4.07 //x2=58.83 //y2=4.07
r479 (  3 4 ) resistor r=27.3187 //w=0.131 //l=28.63 //layer=m1 \
 //thickness=0.36 //x=58.715 //y=4.07 //x2=30.085 //y2=4.07
r480 (  2 6 ) resistor r=0.0738079 //w=0.207 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=4.07 //x2=1.11 //y2=4.07
r481 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=29.855 //y=4.07 //x2=29.97 //y2=4.07
r482 (  1 2 ) resistor r=27.3187 //w=0.131 //l=28.63 //layer=m1 \
 //thickness=0.36 //x=29.855 //y=4.07 //x2=1.225 //y2=4.07
ends PM_TMRDFFSNRNQNX1\%D

subckt PM_TMRDFFSNRNQNX1\%noxref_15 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 \
 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c253 ( 127 0 ) capacitor c=0.023087f //x=60.865 //y=5.02
c254 ( 126 0 ) capacitor c=0.023519f //x=59.985 //y=5.02
c255 ( 125 0 ) capacitor c=0.0224735f //x=59.105 //y=5.02
c256 ( 123 0 ) capacitor c=0.00853354f //x=61.115 //y=0.915
c257 ( 103 0 ) capacitor c=0.0547611f //x=68.725 //y=4.79
c258 ( 102 0 ) capacitor c=0.0294456f //x=69.015 //y=4.79
c259 ( 101 0 ) capacitor c=0.0347816f //x=68.68 //y=1.22
c260 ( 100 0 ) capacitor c=0.0187487f //x=68.68 //y=0.875
c261 ( 94 0 ) capacitor c=0.0137055f //x=68.525 //y=1.375
c262 ( 92 0 ) capacitor c=0.0149861f //x=68.525 //y=0.72
c263 ( 91 0 ) capacitor c=0.096037f //x=68.15 //y=1.915
c264 ( 90 0 ) capacitor c=0.0228993f //x=68.15 //y=1.53
c265 ( 89 0 ) capacitor c=0.0234352f //x=68.15 //y=1.22
c266 ( 88 0 ) capacitor c=0.0198724f //x=68.15 //y=0.875
c267 ( 84 0 ) capacitor c=0.0549166f //x=63.915 //y=4.79
c268 ( 83 0 ) capacitor c=0.0294456f //x=64.205 //y=4.79
c269 ( 82 0 ) capacitor c=0.0347816f //x=63.87 //y=1.22
c270 ( 81 0 ) capacitor c=0.0187487f //x=63.87 //y=0.875
c271 ( 75 0 ) capacitor c=0.0137055f //x=63.715 //y=1.375
c272 ( 73 0 ) capacitor c=0.0149861f //x=63.715 //y=0.72
c273 ( 72 0 ) capacitor c=0.096037f //x=63.34 //y=1.915
c274 ( 71 0 ) capacitor c=0.0228993f //x=63.34 //y=1.53
c275 ( 70 0 ) capacitor c=0.0234352f //x=63.34 //y=1.22
c276 ( 69 0 ) capacitor c=0.0198724f //x=63.34 //y=0.875
c277 ( 68 0 ) capacitor c=0.109949f //x=69.09 //y=6.02
c278 ( 67 0 ) capacitor c=0.158483f //x=68.65 //y=6.02
c279 ( 66 0 ) capacitor c=0.109949f //x=64.28 //y=6.02
c280 ( 65 0 ) capacitor c=0.158483f //x=63.84 //y=6.02
c281 ( 62 0 ) capacitor c=9.74268e-19 //x=61.01 //y=5.155
c282 ( 61 0 ) capacitor c=0.00191414f //x=60.13 //y=5.155
c283 ( 54 0 ) capacitor c=0.0913827f //x=68.45 //y=2.08
c284 ( 46 0 ) capacitor c=0.093372f //x=63.64 //y=2.08
c285 ( 44 0 ) capacitor c=0.105725f //x=61.79 //y=2.59
c286 ( 40 0 ) capacitor c=0.00398962f //x=61.39 //y=1.665
c287 ( 39 0 ) capacitor c=0.0137288f //x=61.705 //y=1.665
c288 ( 33 0 ) capacitor c=0.0276208f //x=61.705 //y=5.155
c289 ( 25 0 ) capacitor c=0.0169868f //x=60.925 //y=5.155
c290 ( 18 0 ) capacitor c=0.00316998f //x=59.335 //y=5.155
c291 ( 17 0 ) capacitor c=0.014258f //x=60.045 //y=5.155
c292 ( 4 0 ) capacitor c=0.00401138f //x=63.755 //y=2.59
c293 ( 3 0 ) capacitor c=0.0706637f //x=68.335 //y=2.59
c294 ( 2 0 ) capacitor c=0.0120752f //x=61.905 //y=2.59
c295 ( 1 0 ) capacitor c=0.0233554f //x=63.525 //y=2.59
r296 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=69.015 //y=4.79 //x2=69.09 //y2=4.865
r297 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=69.015 //y=4.79 //x2=68.725 //y2=4.79
r298 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.68 //y=1.22 //x2=68.64 //y2=1.375
r299 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.68 //y=0.875 //x2=68.64 //y2=0.72
r300 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=68.68 //y=0.875 //x2=68.68 //y2=1.22
r301 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=68.65 //y=4.865 //x2=68.725 //y2=4.79
r302 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=68.65 //y=4.865 //x2=68.45 //y2=4.7
r303 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.305 //y=1.375 //x2=68.19 //y2=1.375
r304 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.525 //y=1.375 //x2=68.64 //y2=1.375
r305 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.305 //y=0.72 //x2=68.19 //y2=0.72
r306 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.525 //y=0.72 //x2=68.64 //y2=0.72
r307 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=68.525 //y=0.72 //x2=68.305 //y2=0.72
r308 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=68.15 //y=1.915 //x2=68.45 //y2=2.08
r309 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.15 //y=1.53 //x2=68.19 //y2=1.375
r310 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=68.15 //y=1.53 //x2=68.15 //y2=1.915
r311 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.15 //y=1.22 //x2=68.19 //y2=1.375
r312 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.15 //y=0.875 //x2=68.19 //y2=0.72
r313 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=68.15 //y=0.875 //x2=68.15 //y2=1.22
r314 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=64.205 //y=4.79 //x2=64.28 //y2=4.865
r315 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=64.205 //y=4.79 //x2=63.915 //y2=4.79
r316 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.87 //y=1.22 //x2=63.83 //y2=1.375
r317 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.87 //y=0.875 //x2=63.83 //y2=0.72
r318 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.87 //y=0.875 //x2=63.87 //y2=1.22
r319 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=63.84 //y=4.865 //x2=63.915 //y2=4.79
r320 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=63.84 //y=4.865 //x2=63.64 //y2=4.7
r321 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.495 //y=1.375 //x2=63.38 //y2=1.375
r322 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.715 //y=1.375 //x2=63.83 //y2=1.375
r323 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.495 //y=0.72 //x2=63.38 //y2=0.72
r324 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.715 //y=0.72 //x2=63.83 //y2=0.72
r325 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=63.715 //y=0.72 //x2=63.495 //y2=0.72
r326 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=63.34 //y=1.915 //x2=63.64 //y2=2.08
r327 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.34 //y=1.53 //x2=63.38 //y2=1.375
r328 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=63.34 //y=1.53 //x2=63.34 //y2=1.915
r329 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.34 //y=1.22 //x2=63.38 //y2=1.375
r330 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.34 //y=0.875 //x2=63.38 //y2=0.72
r331 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.34 //y=0.875 //x2=63.34 //y2=1.22
r332 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.09 //y=6.02 //x2=69.09 //y2=4.865
r333 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=68.65 //y=6.02 //x2=68.65 //y2=4.865
r334 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=64.28 //y=6.02 //x2=64.28 //y2=4.865
r335 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=63.84 //y=6.02 //x2=63.84 //y2=4.865
r336 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=68.415 //y=1.375 //x2=68.525 //y2=1.375
r337 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=68.415 //y=1.375 //x2=68.305 //y2=1.375
r338 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.605 //y=1.375 //x2=63.715 //y2=1.375
r339 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.605 //y=1.375 //x2=63.495 //y2=1.375
r340 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=68.45 //y=4.7 //x2=68.45 //y2=4.7
r341 (  57 59 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=68.45 //y=2.59 //x2=68.45 //y2=4.7
r342 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=68.45 //y=2.08 //x2=68.45 //y2=2.08
r343 (  54 57 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=68.45 //y=2.08 //x2=68.45 //y2=2.59
r344 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.64 //y=4.7 //x2=63.64 //y2=4.7
r345 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=63.64 //y=2.59 //x2=63.64 //y2=4.7
r346 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.64 //y=2.08 //x2=63.64 //y2=2.08
r347 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=63.64 //y=2.08 //x2=63.64 //y2=2.59
r348 (  42 44 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=61.79 //y=5.07 //x2=61.79 //y2=2.59
r349 (  41 44 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=61.79 //y=1.75 //x2=61.79 //y2=2.59
r350 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=61.705 //y=1.665 //x2=61.79 //y2=1.75
r351 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=61.705 //y=1.665 //x2=61.39 //y2=1.665
r352 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=61.305 //y=1.58 //x2=61.39 //y2=1.665
r353 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=61.305 //y=1.58 //x2=61.305 //y2=1.01
r354 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.095 //y=5.155 //x2=61.01 //y2=5.155
r355 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=61.705 //y=5.155 //x2=61.79 //y2=5.07
r356 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=61.705 //y=5.155 //x2=61.095 //y2=5.155
r357 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.01 //y=5.24 //x2=61.01 //y2=5.155
r358 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=61.01 //y=5.24 //x2=61.01 //y2=5.725
r359 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.215 //y=5.155 //x2=60.13 //y2=5.155
r360 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.925 //y=5.155 //x2=61.01 //y2=5.155
r361 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=60.925 //y=5.155 //x2=60.215 //y2=5.155
r362 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.13 //y=5.24 //x2=60.13 //y2=5.155
r363 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.13 //y=5.24 //x2=60.13 //y2=5.725
r364 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.045 //y=5.155 //x2=60.13 //y2=5.155
r365 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=60.045 //y=5.155 //x2=59.335 //y2=5.155
r366 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=59.25 //y=5.24 //x2=59.335 //y2=5.155
r367 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.25 //y=5.24 //x2=59.25 //y2=5.725
r368 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=68.45 //y=2.59 //x2=68.45 //y2=2.59
r369 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=63.64 //y=2.59 //x2=63.64 //y2=2.59
r370 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=61.79 //y=2.59 //x2=61.79 //y2=2.59
r371 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.755 //y=2.59 //x2=63.64 //y2=2.59
r372 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=68.335 //y=2.59 //x2=68.45 //y2=2.59
r373 (  3 4 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=68.335 //y=2.59 //x2=63.755 //y2=2.59
r374 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=61.905 //y=2.59 //x2=61.79 //y2=2.59
r375 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.525 //y=2.59 //x2=63.64 //y2=2.59
r376 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=63.525 //y=2.59 //x2=61.905 //y2=2.59
ends PM_TMRDFFSNRNQNX1\%noxref_15

subckt PM_TMRDFFSNRNQNX1\%noxref_16 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 \
 53 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c168 ( 85 0 ) capacitor c=0.023087f //x=70.485 //y=5.02
c169 ( 84 0 ) capacitor c=0.023519f //x=69.605 //y=5.02
c170 ( 83 0 ) capacitor c=0.0224735f //x=68.725 //y=5.02
c171 ( 81 0 ) capacitor c=0.00853354f //x=70.735 //y=0.915
c172 ( 69 0 ) capacitor c=0.0547611f //x=73.535 //y=4.79
c173 ( 68 0 ) capacitor c=0.0294456f //x=73.825 //y=4.79
c174 ( 67 0 ) capacitor c=0.0347816f //x=73.49 //y=1.22
c175 ( 66 0 ) capacitor c=0.0187487f //x=73.49 //y=0.875
c176 ( 60 0 ) capacitor c=0.0137055f //x=73.335 //y=1.375
c177 ( 58 0 ) capacitor c=0.0149861f //x=73.335 //y=0.72
c178 ( 57 0 ) capacitor c=0.096037f //x=72.96 //y=1.915
c179 ( 56 0 ) capacitor c=0.0228993f //x=72.96 //y=1.53
c180 ( 55 0 ) capacitor c=0.0234352f //x=72.96 //y=1.22
c181 ( 54 0 ) capacitor c=0.0198724f //x=72.96 //y=0.875
c182 ( 53 0 ) capacitor c=0.109949f //x=73.9 //y=6.02
c183 ( 52 0 ) capacitor c=0.158483f //x=73.46 //y=6.02
c184 ( 50 0 ) capacitor c=9.74268e-19 //x=70.63 //y=5.155
c185 ( 49 0 ) capacitor c=0.00191414f //x=69.75 //y=5.155
c186 ( 42 0 ) capacitor c=0.0911502f //x=73.26 //y=2.08
c187 ( 40 0 ) capacitor c=0.103494f //x=71.41 //y=2.59
c188 ( 36 0 ) capacitor c=0.00398962f //x=71.01 //y=1.665
c189 ( 35 0 ) capacitor c=0.0137288f //x=71.325 //y=1.665
c190 ( 29 0 ) capacitor c=0.0276208f //x=71.325 //y=5.155
c191 ( 21 0 ) capacitor c=0.0169868f //x=70.545 //y=5.155
c192 ( 14 0 ) capacitor c=0.00316998f //x=68.955 //y=5.155
c193 ( 13 0 ) capacitor c=0.014258f //x=69.665 //y=5.155
c194 ( 2 0 ) capacitor c=0.00808366f //x=71.525 //y=2.59
c195 ( 1 0 ) capacitor c=0.0351856f //x=73.145 //y=2.59
r196 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=73.825 //y=4.79 //x2=73.9 //y2=4.865
r197 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=73.825 //y=4.79 //x2=73.535 //y2=4.79
r198 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.49 //y=1.22 //x2=73.45 //y2=1.375
r199 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.49 //y=0.875 //x2=73.45 //y2=0.72
r200 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=73.49 //y=0.875 //x2=73.49 //y2=1.22
r201 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=73.46 //y=4.865 //x2=73.535 //y2=4.79
r202 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=73.46 //y=4.865 //x2=73.26 //y2=4.7
r203 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.115 //y=1.375 //x2=73 //y2=1.375
r204 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.335 //y=1.375 //x2=73.45 //y2=1.375
r205 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.115 //y=0.72 //x2=73 //y2=0.72
r206 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.335 //y=0.72 //x2=73.45 //y2=0.72
r207 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=73.335 //y=0.72 //x2=73.115 //y2=0.72
r208 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=72.96 //y=1.915 //x2=73.26 //y2=2.08
r209 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.96 //y=1.53 //x2=73 //y2=1.375
r210 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=72.96 //y=1.53 //x2=72.96 //y2=1.915
r211 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.96 //y=1.22 //x2=73 //y2=1.375
r212 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.96 //y=0.875 //x2=73 //y2=0.72
r213 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=72.96 //y=0.875 //x2=72.96 //y2=1.22
r214 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=73.9 //y=6.02 //x2=73.9 //y2=4.865
r215 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=73.46 //y=6.02 //x2=73.46 //y2=4.865
r216 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=73.225 //y=1.375 //x2=73.335 //y2=1.375
r217 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=73.225 //y=1.375 //x2=73.115 //y2=1.375
r218 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=73.26 //y=4.7 //x2=73.26 //y2=4.7
r219 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=73.26 //y=2.59 //x2=73.26 //y2=4.7
r220 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=73.26 //y=2.08 //x2=73.26 //y2=2.08
r221 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=73.26 //y=2.08 //x2=73.26 //y2=2.59
r222 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=71.41 //y=5.07 //x2=71.41 //y2=2.59
r223 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=71.41 //y=1.75 //x2=71.41 //y2=2.59
r224 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=71.325 //y=1.665 //x2=71.41 //y2=1.75
r225 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=71.325 //y=1.665 //x2=71.01 //y2=1.665
r226 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=70.925 //y=1.58 //x2=71.01 //y2=1.665
r227 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=70.925 //y=1.58 //x2=70.925 //y2=1.01
r228 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.715 //y=5.155 //x2=70.63 //y2=5.155
r229 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=71.325 //y=5.155 //x2=71.41 //y2=5.07
r230 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=71.325 //y=5.155 //x2=70.715 //y2=5.155
r231 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.63 //y=5.24 //x2=70.63 //y2=5.155
r232 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=70.63 //y=5.24 //x2=70.63 //y2=5.725
r233 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.835 //y=5.155 //x2=69.75 //y2=5.155
r234 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.545 //y=5.155 //x2=70.63 //y2=5.155
r235 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=70.545 //y=5.155 //x2=69.835 //y2=5.155
r236 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.75 //y=5.24 //x2=69.75 //y2=5.155
r237 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=69.75 //y=5.24 //x2=69.75 //y2=5.725
r238 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.665 //y=5.155 //x2=69.75 //y2=5.155
r239 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=69.665 //y=5.155 //x2=68.955 //y2=5.155
r240 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=68.87 //y=5.24 //x2=68.955 //y2=5.155
r241 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=68.87 //y=5.24 //x2=68.87 //y2=5.725
r242 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=73.26 //y=2.59 //x2=73.26 //y2=2.59
r243 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=71.41 //y=2.59 //x2=71.41 //y2=2.59
r244 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=71.525 //y=2.59 //x2=71.41 //y2=2.59
r245 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=73.145 //y=2.59 //x2=73.26 //y2=2.59
r246 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=73.145 //y=2.59 //x2=71.525 //y2=2.59
ends PM_TMRDFFSNRNQNX1\%noxref_16

subckt PM_TMRDFFSNRNQNX1\%CLK ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 \
 31 32 33 34 36 46 55 64 73 81 89 90 91 92 93 94 95 96 97 98 99 100 101 102 \
 103 104 105 106 107 108 109 111 117 118 119 120 121 126 127 128 130 136 137 \
 138 139 140 145 146 147 149 155 156 157 158 159 164 165 166 168 174 175 176 \
 177 178 183 184 185 187 193 194 195 196 197 202 203 204 206 212 213 214 215 \
 216 224 235 246 257 268 279 )
c707 ( 279 0 ) capacitor c=0.0333177f //x=74.37 //y=4.7
c708 ( 268 0 ) capacitor c=0.0333177f //x=64.75 //y=4.7
c709 ( 257 0 ) capacitor c=0.0333177f //x=45.51 //y=4.7
c710 ( 246 0 ) capacitor c=0.0333177f //x=35.89 //y=4.7
c711 ( 235 0 ) capacitor c=0.0334842f //x=16.65 //y=4.7
c712 ( 224 0 ) capacitor c=0.0334842f //x=7.03 //y=4.7
c713 ( 216 0 ) capacitor c=0.0252241f //x=74.705 //y=4.79
c714 ( 215 0 ) capacitor c=0.0825763f //x=74.46 //y=1.915
c715 ( 214 0 ) capacitor c=0.0170266f //x=74.46 //y=1.45
c716 ( 213 0 ) capacitor c=0.018609f //x=74.46 //y=1.22
c717 ( 212 0 ) capacitor c=0.0187309f //x=74.46 //y=0.91
c718 ( 206 0 ) capacitor c=0.014725f //x=74.305 //y=1.375
c719 ( 204 0 ) capacitor c=0.0146567f //x=74.305 //y=0.755
c720 ( 203 0 ) capacitor c=0.0335408f //x=73.935 //y=1.22
c721 ( 202 0 ) capacitor c=0.0173761f //x=73.935 //y=0.91
c722 ( 197 0 ) capacitor c=0.0246783f //x=65.085 //y=4.79
c723 ( 196 0 ) capacitor c=0.0825763f //x=64.84 //y=1.915
c724 ( 195 0 ) capacitor c=0.0170266f //x=64.84 //y=1.45
c725 ( 194 0 ) capacitor c=0.018609f //x=64.84 //y=1.22
c726 ( 193 0 ) capacitor c=0.0187309f //x=64.84 //y=0.91
c727 ( 187 0 ) capacitor c=0.014725f //x=64.685 //y=1.375
c728 ( 185 0 ) capacitor c=0.0146567f //x=64.685 //y=0.755
c729 ( 184 0 ) capacitor c=0.0335408f //x=64.315 //y=1.22
c730 ( 183 0 ) capacitor c=0.0173761f //x=64.315 //y=0.91
c731 ( 178 0 ) capacitor c=0.0246783f //x=45.845 //y=4.79
c732 ( 177 0 ) capacitor c=0.0825763f //x=45.6 //y=1.915
c733 ( 176 0 ) capacitor c=0.0170266f //x=45.6 //y=1.45
c734 ( 175 0 ) capacitor c=0.018609f //x=45.6 //y=1.22
c735 ( 174 0 ) capacitor c=0.0187309f //x=45.6 //y=0.91
c736 ( 168 0 ) capacitor c=0.014725f //x=45.445 //y=1.375
c737 ( 166 0 ) capacitor c=0.0146567f //x=45.445 //y=0.755
c738 ( 165 0 ) capacitor c=0.0335408f //x=45.075 //y=1.22
c739 ( 164 0 ) capacitor c=0.0173761f //x=45.075 //y=0.91
c740 ( 159 0 ) capacitor c=0.0246783f //x=36.225 //y=4.79
c741 ( 158 0 ) capacitor c=0.0825763f //x=35.98 //y=1.915
c742 ( 157 0 ) capacitor c=0.0170266f //x=35.98 //y=1.45
c743 ( 156 0 ) capacitor c=0.018609f //x=35.98 //y=1.22
c744 ( 155 0 ) capacitor c=0.0187309f //x=35.98 //y=0.91
c745 ( 149 0 ) capacitor c=0.014725f //x=35.825 //y=1.375
c746 ( 147 0 ) capacitor c=0.0146567f //x=35.825 //y=0.755
c747 ( 146 0 ) capacitor c=0.0335408f //x=35.455 //y=1.22
c748 ( 145 0 ) capacitor c=0.0173761f //x=35.455 //y=0.91
c749 ( 140 0 ) capacitor c=0.0245352f //x=16.985 //y=4.79
c750 ( 139 0 ) capacitor c=0.0825763f //x=16.74 //y=1.915
c751 ( 138 0 ) capacitor c=0.0170266f //x=16.74 //y=1.45
c752 ( 137 0 ) capacitor c=0.018609f //x=16.74 //y=1.22
c753 ( 136 0 ) capacitor c=0.0187309f //x=16.74 //y=0.91
c754 ( 130 0 ) capacitor c=0.014725f //x=16.585 //y=1.375
c755 ( 128 0 ) capacitor c=0.0146567f //x=16.585 //y=0.755
c756 ( 127 0 ) capacitor c=0.0335408f //x=16.215 //y=1.22
c757 ( 126 0 ) capacitor c=0.0173761f //x=16.215 //y=0.91
c758 ( 121 0 ) capacitor c=0.0245352f //x=7.365 //y=4.79
c759 ( 120 0 ) capacitor c=0.0825763f //x=7.12 //y=1.915
c760 ( 119 0 ) capacitor c=0.0170266f //x=7.12 //y=1.45
c761 ( 118 0 ) capacitor c=0.018609f //x=7.12 //y=1.22
c762 ( 117 0 ) capacitor c=0.0187309f //x=7.12 //y=0.91
c763 ( 111 0 ) capacitor c=0.014725f //x=6.965 //y=1.375
c764 ( 109 0 ) capacitor c=0.0146567f //x=6.965 //y=0.755
c765 ( 108 0 ) capacitor c=0.0335408f //x=6.595 //y=1.22
c766 ( 107 0 ) capacitor c=0.0173761f //x=6.595 //y=0.91
c767 ( 106 0 ) capacitor c=0.109949f //x=74.78 //y=6.02
c768 ( 105 0 ) capacitor c=0.109956f //x=74.34 //y=6.02
c769 ( 104 0 ) capacitor c=0.109949f //x=65.16 //y=6.02
c770 ( 103 0 ) capacitor c=0.109956f //x=64.72 //y=6.02
c771 ( 102 0 ) capacitor c=0.109949f //x=45.92 //y=6.02
c772 ( 101 0 ) capacitor c=0.109956f //x=45.48 //y=6.02
c773 ( 100 0 ) capacitor c=0.109949f //x=36.3 //y=6.02
c774 ( 99 0 ) capacitor c=0.109956f //x=35.86 //y=6.02
c775 ( 98 0 ) capacitor c=0.110114f //x=17.06 //y=6.02
c776 ( 97 0 ) capacitor c=0.11012f //x=16.62 //y=6.02
c777 ( 96 0 ) capacitor c=0.110114f //x=7.44 //y=6.02
c778 ( 95 0 ) capacitor c=0.11012f //x=7 //y=6.02
c779 ( 81 0 ) capacitor c=0.0880092f //x=74.37 //y=2.08
c780 ( 73 0 ) capacitor c=0.0867127f //x=64.75 //y=2.08
c781 ( 64 0 ) capacitor c=0.0882702f //x=45.51 //y=2.08
c782 ( 55 0 ) capacitor c=0.088164f //x=35.89 //y=2.08
c783 ( 46 0 ) capacitor c=0.0899873f //x=16.65 //y=2.08
c784 ( 36 0 ) capacitor c=0.0925246f //x=7.03 //y=2.08
c785 ( 10 0 ) capacitor c=0.0052048f //x=64.865 //y=4.44
c786 ( 9 0 ) capacitor c=0.124137f //x=74.255 //y=4.44
c787 ( 8 0 ) capacitor c=0.00494979f //x=45.625 //y=4.44
c788 ( 7 0 ) capacitor c=0.255004f //x=64.635 //y=4.44
c789 ( 6 0 ) capacitor c=0.00494979f //x=36.005 //y=4.44
c790 ( 5 0 ) capacitor c=0.117333f //x=45.395 //y=4.44
c791 ( 4 0 ) capacitor c=0.00697397f //x=16.765 //y=4.44
c792 ( 3 0 ) capacitor c=0.297275f //x=35.775 //y=4.44
c793 ( 2 0 ) capacitor c=0.0154455f //x=7.145 //y=4.44
c794 ( 1 0 ) capacitor c=0.212324f //x=16.535 //y=4.44
r795 (  281 282 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=74.37 //y=4.79 //x2=74.37 //y2=4.865
r796 (  279 281 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=74.37 //y=4.7 //x2=74.37 //y2=4.79
r797 (  270 271 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=64.75 //y=4.79 //x2=64.75 //y2=4.865
r798 (  268 270 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=64.75 //y=4.7 //x2=64.75 //y2=4.79
r799 (  259 260 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=45.51 //y=4.79 //x2=45.51 //y2=4.865
r800 (  257 259 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=45.51 //y=4.7 //x2=45.51 //y2=4.79
r801 (  248 249 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=35.89 //y=4.79 //x2=35.89 //y2=4.865
r802 (  246 248 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=35.89 //y=4.7 //x2=35.89 //y2=4.79
r803 (  237 238 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=16.65 //y=4.79 //x2=16.65 //y2=4.865
r804 (  235 237 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=16.65 //y=4.7 //x2=16.65 //y2=4.79
r805 (  226 227 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.79 //x2=7.03 //y2=4.865
r806 (  224 226 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.7 //x2=7.03 //y2=4.79
r807 (  217 281 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=74.505 //y=4.79 //x2=74.37 //y2=4.79
r808 (  216 218 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=74.705 //y=4.79 //x2=74.78 //y2=4.865
r809 (  216 217 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=74.705 //y=4.79 //x2=74.505 //y2=4.79
r810 (  215 286 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=74.46 //y=1.915 //x2=74.385 //y2=2.08
r811 (  214 284 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=74.46 //y=1.45 //x2=74.42 //y2=1.375
r812 (  214 215 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=74.46 //y=1.45 //x2=74.46 //y2=1.915
r813 (  213 284 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.46 //y=1.22 //x2=74.42 //y2=1.375
r814 (  212 283 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.46 //y=0.91 //x2=74.42 //y2=0.755
r815 (  212 213 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=74.46 //y=0.91 //x2=74.46 //y2=1.22
r816 (  207 277 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.09 //y=1.375 //x2=73.975 //y2=1.375
r817 (  206 284 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.305 //y=1.375 //x2=74.42 //y2=1.375
r818 (  205 276 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.09 //y=0.755 //x2=73.975 //y2=0.755
r819 (  204 283 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.305 //y=0.755 //x2=74.42 //y2=0.755
r820 (  204 205 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=74.305 //y=0.755 //x2=74.09 //y2=0.755
r821 (  203 277 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.935 //y=1.22 //x2=73.975 //y2=1.375
r822 (  202 276 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.935 //y=0.91 //x2=73.975 //y2=0.755
r823 (  202 203 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=73.935 //y=0.91 //x2=73.935 //y2=1.22
r824 (  198 270 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=64.885 //y=4.79 //x2=64.75 //y2=4.79
r825 (  197 199 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=65.085 //y=4.79 //x2=65.16 //y2=4.865
r826 (  197 198 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=65.085 //y=4.79 //x2=64.885 //y2=4.79
r827 (  196 275 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=64.84 //y=1.915 //x2=64.765 //y2=2.08
r828 (  195 273 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=64.84 //y=1.45 //x2=64.8 //y2=1.375
r829 (  195 196 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=64.84 //y=1.45 //x2=64.84 //y2=1.915
r830 (  194 273 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.84 //y=1.22 //x2=64.8 //y2=1.375
r831 (  193 272 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.84 //y=0.91 //x2=64.8 //y2=0.755
r832 (  193 194 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=64.84 //y=0.91 //x2=64.84 //y2=1.22
r833 (  188 266 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.47 //y=1.375 //x2=64.355 //y2=1.375
r834 (  187 273 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.685 //y=1.375 //x2=64.8 //y2=1.375
r835 (  186 265 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.47 //y=0.755 //x2=64.355 //y2=0.755
r836 (  185 272 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.685 //y=0.755 //x2=64.8 //y2=0.755
r837 (  185 186 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=64.685 //y=0.755 //x2=64.47 //y2=0.755
r838 (  184 266 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.315 //y=1.22 //x2=64.355 //y2=1.375
r839 (  183 265 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.315 //y=0.91 //x2=64.355 //y2=0.755
r840 (  183 184 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=64.315 //y=0.91 //x2=64.315 //y2=1.22
r841 (  179 259 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=45.645 //y=4.79 //x2=45.51 //y2=4.79
r842 (  178 180 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=45.845 //y=4.79 //x2=45.92 //y2=4.865
r843 (  178 179 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=45.845 //y=4.79 //x2=45.645 //y2=4.79
r844 (  177 264 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=45.6 //y=1.915 //x2=45.525 //y2=2.08
r845 (  176 262 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=45.6 //y=1.45 //x2=45.56 //y2=1.375
r846 (  176 177 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=45.6 //y=1.45 //x2=45.6 //y2=1.915
r847 (  175 262 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.6 //y=1.22 //x2=45.56 //y2=1.375
r848 (  174 261 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.6 //y=0.91 //x2=45.56 //y2=0.755
r849 (  174 175 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=45.6 //y=0.91 //x2=45.6 //y2=1.22
r850 (  169 255 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.23 //y=1.375 //x2=45.115 //y2=1.375
r851 (  168 262 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.445 //y=1.375 //x2=45.56 //y2=1.375
r852 (  167 254 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.23 //y=0.755 //x2=45.115 //y2=0.755
r853 (  166 261 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.445 //y=0.755 //x2=45.56 //y2=0.755
r854 (  166 167 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=45.445 //y=0.755 //x2=45.23 //y2=0.755
r855 (  165 255 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.075 //y=1.22 //x2=45.115 //y2=1.375
r856 (  164 254 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.075 //y=0.91 //x2=45.115 //y2=0.755
r857 (  164 165 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=45.075 //y=0.91 //x2=45.075 //y2=1.22
r858 (  160 248 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=36.025 //y=4.79 //x2=35.89 //y2=4.79
r859 (  159 161 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=36.225 //y=4.79 //x2=36.3 //y2=4.865
r860 (  159 160 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=36.225 //y=4.79 //x2=36.025 //y2=4.79
r861 (  158 253 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=35.98 //y=1.915 //x2=35.905 //y2=2.08
r862 (  157 251 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=35.98 //y=1.45 //x2=35.94 //y2=1.375
r863 (  157 158 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=35.98 //y=1.45 //x2=35.98 //y2=1.915
r864 (  156 251 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.98 //y=1.22 //x2=35.94 //y2=1.375
r865 (  155 250 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.98 //y=0.91 //x2=35.94 //y2=0.755
r866 (  155 156 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=35.98 //y=0.91 //x2=35.98 //y2=1.22
r867 (  150 244 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.61 //y=1.375 //x2=35.495 //y2=1.375
r868 (  149 251 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.825 //y=1.375 //x2=35.94 //y2=1.375
r869 (  148 243 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.61 //y=0.755 //x2=35.495 //y2=0.755
r870 (  147 250 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.825 //y=0.755 //x2=35.94 //y2=0.755
r871 (  147 148 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=35.825 //y=0.755 //x2=35.61 //y2=0.755
r872 (  146 244 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.455 //y=1.22 //x2=35.495 //y2=1.375
r873 (  145 243 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.455 //y=0.91 //x2=35.495 //y2=0.755
r874 (  145 146 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=35.455 //y=0.91 //x2=35.455 //y2=1.22
r875 (  141 237 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=16.785 //y=4.79 //x2=16.65 //y2=4.79
r876 (  140 142 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=16.985 //y=4.79 //x2=17.06 //y2=4.865
r877 (  140 141 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=16.985 //y=4.79 //x2=16.785 //y2=4.79
r878 (  139 242 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.915 //x2=16.665 //y2=2.08
r879 (  138 240 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.45 //x2=16.7 //y2=1.375
r880 (  138 139 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.45 //x2=16.74 //y2=1.915
r881 (  137 240 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.22 //x2=16.7 //y2=1.375
r882 (  136 239 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.74 //y=0.91 //x2=16.7 //y2=0.755
r883 (  136 137 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=16.74 //y=0.91 //x2=16.74 //y2=1.22
r884 (  131 233 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.37 //y=1.375 //x2=16.255 //y2=1.375
r885 (  130 240 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.585 //y=1.375 //x2=16.7 //y2=1.375
r886 (  129 232 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.37 //y=0.755 //x2=16.255 //y2=0.755
r887 (  128 239 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.585 //y=0.755 //x2=16.7 //y2=0.755
r888 (  128 129 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=16.585 //y=0.755 //x2=16.37 //y2=0.755
r889 (  127 233 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.215 //y=1.22 //x2=16.255 //y2=1.375
r890 (  126 232 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.215 //y=0.91 //x2=16.255 //y2=0.755
r891 (  126 127 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=16.215 //y=0.91 //x2=16.215 //y2=1.22
r892 (  122 226 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=7.165 //y=4.79 //x2=7.03 //y2=4.79
r893 (  121 123 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.44 //y2=4.865
r894 (  121 122 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.165 //y2=4.79
r895 (  120 231 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.915 //x2=7.045 //y2=2.08
r896 (  119 229 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.08 //y2=1.375
r897 (  119 120 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.12 //y2=1.915
r898 (  118 229 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.22 //x2=7.08 //y2=1.375
r899 (  117 228 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.08 //y2=0.755
r900 (  117 118 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.12 //y2=1.22
r901 (  112 222 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=1.375 //x2=6.635 //y2=1.375
r902 (  111 229 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=1.375 //x2=7.08 //y2=1.375
r903 (  110 221 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=0.755 //x2=6.635 //y2=0.755
r904 (  109 228 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=7.08 //y2=0.755
r905 (  109 110 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=6.75 //y2=0.755
r906 (  108 222 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=1.22 //x2=6.635 //y2=1.375
r907 (  107 221 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.635 //y2=0.755
r908 (  107 108 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.595 //y2=1.22
r909 (  106 218 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=74.78 //y=6.02 //x2=74.78 //y2=4.865
r910 (  105 282 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=74.34 //y=6.02 //x2=74.34 //y2=4.865
r911 (  104 199 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=65.16 //y=6.02 //x2=65.16 //y2=4.865
r912 (  103 271 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=64.72 //y=6.02 //x2=64.72 //y2=4.865
r913 (  102 180 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.92 //y=6.02 //x2=45.92 //y2=4.865
r914 (  101 260 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.48 //y=6.02 //x2=45.48 //y2=4.865
r915 (  100 161 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=36.3 //y=6.02 //x2=36.3 //y2=4.865
r916 (  99 249 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.86 //y=6.02 //x2=35.86 //y2=4.865
r917 (  98 142 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.06 //y=6.02 //x2=17.06 //y2=4.865
r918 (  97 238 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.62 //y=6.02 //x2=16.62 //y2=4.865
r919 (  96 123 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.44 //y=6.02 //x2=7.44 //y2=4.865
r920 (  95 227 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7 //y=6.02 //x2=7 //y2=4.865
r921 (  94 206 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=74.197 //y=1.375 //x2=74.305 //y2=1.375
r922 (  94 207 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=74.197 //y=1.375 //x2=74.09 //y2=1.375
r923 (  93 187 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=64.577 //y=1.375 //x2=64.685 //y2=1.375
r924 (  93 188 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=64.577 //y=1.375 //x2=64.47 //y2=1.375
r925 (  92 168 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=45.337 //y=1.375 //x2=45.445 //y2=1.375
r926 (  92 169 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=45.337 //y=1.375 //x2=45.23 //y2=1.375
r927 (  91 149 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=35.717 //y=1.375 //x2=35.825 //y2=1.375
r928 (  91 150 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=35.717 //y=1.375 //x2=35.61 //y2=1.375
r929 (  90 130 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=16.477 //y=1.375 //x2=16.585 //y2=1.375
r930 (  90 131 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=16.477 //y=1.375 //x2=16.37 //y2=1.375
r931 (  89 111 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.965 //y2=1.375
r932 (  89 112 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.75 //y2=1.375
r933 (  87 279 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=74.37 //y=4.7 //x2=74.37 //y2=4.7
r934 (  81 286 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=74.37 //y=2.08 //x2=74.37 //y2=2.08
r935 (  78 268 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=64.75 //y=4.7 //x2=64.75 //y2=4.7
r936 (  73 275 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=64.75 //y=2.08 //x2=64.75 //y2=2.08
r937 (  70 257 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.51 //y=4.7 //x2=45.51 //y2=4.7
r938 (  64 264 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.51 //y=2.08 //x2=45.51 //y2=2.08
r939 (  61 246 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.89 //y=4.7 //x2=35.89 //y2=4.7
r940 (  55 253 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.89 //y=2.08 //x2=35.89 //y2=2.08
r941 (  52 235 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=4.7 //x2=16.65 //y2=4.7
r942 (  46 242 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=2.08 //x2=16.65 //y2=2.08
r943 (  43 224 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=4.7 //x2=7.03 //y2=4.7
r944 (  36 231 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=2.08 //x2=7.03 //y2=2.08
r945 (  34 87 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=74.37 //y=4.44 //x2=74.37 //y2=4.7
r946 (  33 34 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=74.37 //y=2.59 //x2=74.37 //y2=4.44
r947 (  33 81 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=74.37 //y=2.59 //x2=74.37 //y2=2.08
r948 (  32 78 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=64.75 //y=4.44 //x2=64.75 //y2=4.7
r949 (  32 73 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=64.75 //y=4.44 //x2=64.75 //y2=2.08
r950 (  31 70 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=45.51 //y=4.44 //x2=45.51 //y2=4.7
r951 (  30 31 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=45.51 //y=2.59 //x2=45.51 //y2=4.44
r952 (  30 64 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=45.51 //y=2.59 //x2=45.51 //y2=2.08
r953 (  29 61 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=35.89 //y=4.44 //x2=35.89 //y2=4.7
r954 (  28 29 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=35.89 //y=3.7 //x2=35.89 //y2=4.44
r955 (  28 55 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=35.89 //y=3.7 //x2=35.89 //y2=2.08
r956 (  27 52 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.44 //x2=16.65 //y2=4.7
r957 (  26 27 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.59 //x2=16.65 //y2=4.44
r958 (  26 46 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.59 //x2=16.65 //y2=2.08
r959 (  25 43 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=7.03 //y=4.44 //x2=7.03 //y2=4.7
r960 (  24 25 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=7.03 //y=3.7 //x2=7.03 //y2=4.44
r961 (  23 24 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.96 //x2=7.03 //y2=3.7
r962 (  23 36 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.96 //x2=7.03 //y2=2.08
r963 (  22 34 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=74.37 //y=4.44 //x2=74.37 //y2=4.44
r964 (  20 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=64.75 //y=4.44 //x2=64.75 //y2=4.44
r965 (  18 31 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=45.51 //y=4.44 //x2=45.51 //y2=4.44
r966 (  16 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=35.89 //y=4.44 //x2=35.89 //y2=4.44
r967 (  14 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=16.65 //y=4.44 //x2=16.65 //y2=4.44
r968 (  12 25 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.03 //y=4.44 //x2=7.03 //y2=4.44
r969 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=64.865 //y=4.44 //x2=64.75 //y2=4.44
r970 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=74.255 //y=4.44 //x2=74.37 //y2=4.44
r971 (  9 10 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=74.255 //y=4.44 //x2=64.865 //y2=4.44
r972 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.625 //y=4.44 //x2=45.51 //y2=4.44
r973 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=64.635 //y=4.44 //x2=64.75 //y2=4.44
r974 (  7 8 ) resistor r=18.1393 //w=0.131 //l=19.01 //layer=m1 \
 //thickness=0.36 //x=64.635 //y=4.44 //x2=45.625 //y2=4.44
r975 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=36.005 //y=4.44 //x2=35.89 //y2=4.44
r976 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.395 //y=4.44 //x2=45.51 //y2=4.44
r977 (  5 6 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=45.395 //y=4.44 //x2=36.005 //y2=4.44
r978 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.765 //y=4.44 //x2=16.65 //y2=4.44
r979 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=35.775 //y=4.44 //x2=35.89 //y2=4.44
r980 (  3 4 ) resistor r=18.1393 //w=0.131 //l=19.01 //layer=m1 \
 //thickness=0.36 //x=35.775 //y=4.44 //x2=16.765 //y2=4.44
r981 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.145 //y=4.44 //x2=7.03 //y2=4.44
r982 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.535 //y=4.44 //x2=16.65 //y2=4.44
r983 (  1 2 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=16.535 //y=4.44 //x2=7.145 //y2=4.44
ends PM_TMRDFFSNRNQNX1\%CLK

subckt PM_TMRDFFSNRNQNX1\%noxref_18 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 \
 63 64 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 90 92 98 99 100 101 106 \
 107 112 123 125 126 127 )
c274 ( 127 0 ) capacitor c=0.023087f //x=65.675 //y=5.02
c275 ( 126 0 ) capacitor c=0.023519f //x=64.795 //y=5.02
c276 ( 125 0 ) capacitor c=0.0224735f //x=63.915 //y=5.02
c277 ( 123 0 ) capacitor c=0.00853354f //x=65.925 //y=0.915
c278 ( 112 0 ) capacitor c=0.0588394f //x=61.05 //y=4.7
c279 ( 107 0 ) capacitor c=0.0273931f //x=61.05 //y=1.915
c280 ( 106 0 ) capacitor c=0.0456313f //x=61.05 //y=2.08
c281 ( 101 0 ) capacitor c=0.0556143f //x=78.345 //y=4.79
c282 ( 100 0 ) capacitor c=0.0293157f //x=78.635 //y=4.79
c283 ( 99 0 ) capacitor c=0.0347816f //x=78.3 //y=1.22
c284 ( 98 0 ) capacitor c=0.0187487f //x=78.3 //y=0.875
c285 ( 92 0 ) capacitor c=0.0137055f //x=78.145 //y=1.375
c286 ( 90 0 ) capacitor c=0.0149861f //x=78.145 //y=0.72
c287 ( 89 0 ) capacitor c=0.096037f //x=77.77 //y=1.915
c288 ( 88 0 ) capacitor c=0.0228993f //x=77.77 //y=1.53
c289 ( 87 0 ) capacitor c=0.0234352f //x=77.77 //y=1.22
c290 ( 86 0 ) capacitor c=0.0198724f //x=77.77 //y=0.875
c291 ( 85 0 ) capacitor c=0.0432517f //x=61.57 //y=1.26
c292 ( 84 0 ) capacitor c=0.0200379f //x=61.57 //y=0.915
c293 ( 81 0 ) capacitor c=0.0148873f //x=61.415 //y=1.415
c294 ( 79 0 ) capacitor c=0.0157803f //x=61.415 //y=0.76
c295 ( 74 0 ) capacitor c=0.0218028f //x=61.04 //y=1.57
c296 ( 73 0 ) capacitor c=0.0207459f //x=61.04 //y=1.26
c297 ( 72 0 ) capacitor c=0.0194308f //x=61.04 //y=0.915
c298 ( 68 0 ) capacitor c=0.110114f //x=78.71 //y=6.02
c299 ( 67 0 ) capacitor c=0.158956f //x=78.27 //y=6.02
c300 ( 66 0 ) capacitor c=0.158754f //x=61.23 //y=6.02
c301 ( 65 0 ) capacitor c=0.109949f //x=60.79 //y=6.02
c302 ( 62 0 ) capacitor c=9.74268e-19 //x=65.82 //y=5.155
c303 ( 61 0 ) capacitor c=0.00191414f //x=64.94 //y=5.155
c304 ( 54 0 ) capacitor c=0.0958029f //x=78.07 //y=2.08
c305 ( 52 0 ) capacitor c=0.1027f //x=66.6 //y=3.33
c306 ( 48 0 ) capacitor c=0.00398962f //x=66.2 //y=1.665
c307 ( 47 0 ) capacitor c=0.0137288f //x=66.515 //y=1.665
c308 ( 41 0 ) capacitor c=0.0276208f //x=66.515 //y=5.155
c309 ( 33 0 ) capacitor c=0.0169868f //x=65.735 //y=5.155
c310 ( 26 0 ) capacitor c=0.00316998f //x=64.145 //y=5.155
c311 ( 25 0 ) capacitor c=0.014258f //x=64.855 //y=5.155
c312 ( 12 0 ) capacitor c=0.0814556f //x=61.05 //y=2.08
c313 ( 4 0 ) capacitor c=0.00551333f //x=66.715 //y=3.33
c314 ( 3 0 ) capacitor c=0.17826f //x=77.955 //y=3.33
c315 ( 2 0 ) capacitor c=0.0109971f //x=61.165 //y=3.33
c316 ( 1 0 ) capacitor c=0.077341f //x=66.485 //y=3.33
r317 (  106 107 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=61.05 //y=2.08 //x2=61.05 //y2=1.915
r318 (  100 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=78.635 //y=4.79 //x2=78.71 //y2=4.865
r319 (  100 101 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=78.635 //y=4.79 //x2=78.345 //y2=4.79
r320 (  99 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.3 //y=1.22 //x2=78.26 //y2=1.375
r321 (  98 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.3 //y=0.875 //x2=78.26 //y2=0.72
r322 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=78.3 //y=0.875 //x2=78.3 //y2=1.22
r323 (  95 101 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=78.27 //y=4.865 //x2=78.345 //y2=4.79
r324 (  95 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=78.27 //y=4.865 //x2=78.07 //y2=4.7
r325 (  93 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.925 //y=1.375 //x2=77.81 //y2=1.375
r326 (  92 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.145 //y=1.375 //x2=78.26 //y2=1.375
r327 (  91 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.925 //y=0.72 //x2=77.81 //y2=0.72
r328 (  90 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.145 //y=0.72 //x2=78.26 //y2=0.72
r329 (  90 91 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=78.145 //y=0.72 //x2=77.925 //y2=0.72
r330 (  89 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.915 //x2=78.07 //y2=2.08
r331 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.53 //x2=77.81 //y2=1.375
r332 (  88 89 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.53 //x2=77.77 //y2=1.915
r333 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.22 //x2=77.81 //y2=1.375
r334 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.77 //y=0.875 //x2=77.81 //y2=0.72
r335 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=77.77 //y=0.875 //x2=77.77 //y2=1.22
r336 (  85 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.57 //y=1.26 //x2=61.53 //y2=1.415
r337 (  84 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.57 //y=0.915 //x2=61.53 //y2=0.76
r338 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=61.57 //y=0.915 //x2=61.57 //y2=1.26
r339 (  82 110 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=61.195 //y=1.415 //x2=61.08 //y2=1.415
r340 (  81 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=61.415 //y=1.415 //x2=61.53 //y2=1.415
r341 (  80 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=61.195 //y=0.76 //x2=61.08 //y2=0.76
r342 (  79 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=61.415 //y=0.76 //x2=61.53 //y2=0.76
r343 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=61.415 //y=0.76 //x2=61.195 //y2=0.76
r344 (  76 112 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=61.23 //y=4.865 //x2=61.05 //y2=4.7
r345 (  74 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.04 //y=1.57 //x2=61.08 //y2=1.415
r346 (  74 107 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=61.04 //y=1.57 //x2=61.04 //y2=1.915
r347 (  73 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.04 //y=1.26 //x2=61.08 //y2=1.415
r348 (  72 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.04 //y=0.915 //x2=61.08 //y2=0.76
r349 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=61.04 //y=0.915 //x2=61.04 //y2=1.26
r350 (  69 112 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=60.79 //y=4.865 //x2=61.05 //y2=4.7
r351 (  68 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.71 //y=6.02 //x2=78.71 //y2=4.865
r352 (  67 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.27 //y=6.02 //x2=78.27 //y2=4.865
r353 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=61.23 //y=6.02 //x2=61.23 //y2=4.865
r354 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.79 //y=6.02 //x2=60.79 //y2=4.865
r355 (  64 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.035 //y=1.375 //x2=78.145 //y2=1.375
r356 (  64 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.035 //y=1.375 //x2=77.925 //y2=1.375
r357 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=61.305 //y=1.415 //x2=61.415 //y2=1.415
r358 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=61.305 //y=1.415 //x2=61.195 //y2=1.415
r359 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=78.07 //y=4.7 //x2=78.07 //y2=4.7
r360 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=78.07 //y=3.33 //x2=78.07 //y2=4.7
r361 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=78.07 //y=2.08 //x2=78.07 //y2=2.08
r362 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=78.07 //y=2.08 //x2=78.07 //y2=3.33
r363 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=66.6 //y=5.07 //x2=66.6 //y2=3.33
r364 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=66.6 //y=1.75 //x2=66.6 //y2=3.33
r365 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=66.515 //y=1.665 //x2=66.6 //y2=1.75
r366 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=66.515 //y=1.665 //x2=66.2 //y2=1.665
r367 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=66.115 //y=1.58 //x2=66.2 //y2=1.665
r368 (  43 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=66.115 //y=1.58 //x2=66.115 //y2=1.01
r369 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.905 //y=5.155 //x2=65.82 //y2=5.155
r370 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=66.515 //y=5.155 //x2=66.6 //y2=5.07
r371 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=66.515 //y=5.155 //x2=65.905 //y2=5.155
r372 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.82 //y=5.24 //x2=65.82 //y2=5.155
r373 (  35 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=65.82 //y=5.24 //x2=65.82 //y2=5.725
r374 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.025 //y=5.155 //x2=64.94 //y2=5.155
r375 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.735 //y=5.155 //x2=65.82 //y2=5.155
r376 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=65.735 //y=5.155 //x2=65.025 //y2=5.155
r377 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.94 //y=5.24 //x2=64.94 //y2=5.155
r378 (  27 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=64.94 //y=5.24 //x2=64.94 //y2=5.725
r379 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.855 //y=5.155 //x2=64.94 //y2=5.155
r380 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=64.855 //y=5.155 //x2=64.145 //y2=5.155
r381 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=64.06 //y=5.24 //x2=64.145 //y2=5.155
r382 (  19 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=64.06 //y=5.24 //x2=64.06 //y2=5.725
r383 (  17 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=61.05 //y=4.7 //x2=61.05 //y2=4.7
r384 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=61.05 //y=3.33 //x2=61.05 //y2=4.7
r385 (  12 106 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=61.05 //y=2.08 //x2=61.05 //y2=2.08
r386 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=61.05 //y=2.08 //x2=61.05 //y2=3.33
r387 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=78.07 //y=3.33 //x2=78.07 //y2=3.33
r388 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.6 //y=3.33 //x2=66.6 //y2=3.33
r389 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=61.05 //y=3.33 //x2=61.05 //y2=3.33
r390 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.715 //y=3.33 //x2=66.6 //y2=3.33
r391 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=77.955 //y=3.33 //x2=78.07 //y2=3.33
r392 (  3 4 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=77.955 //y=3.33 //x2=66.715 //y2=3.33
r393 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=61.165 //y=3.33 //x2=61.05 //y2=3.33
r394 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.485 //y=3.33 //x2=66.6 //y2=3.33
r395 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=66.485 //y=3.33 //x2=61.165 //y2=3.33
ends PM_TMRDFFSNRNQNX1\%noxref_18

subckt PM_TMRDFFSNRNQNX1\%RN ( 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 35 36 37 \
 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 \
 65 78 87 97 108 117 127 138 147 156 157 158 159 160 161 162 163 164 165 166 \
 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 \
 187 193 194 195 196 197 205 206 207 212 214 217 218 219 220 221 223 229 230 \
 231 232 233 238 239 240 242 248 249 250 251 252 260 261 262 267 269 272 273 \
 274 275 276 278 284 285 286 287 288 293 294 295 297 303 304 305 306 307 315 \
 316 317 322 324 327 328 329 330 331 333 339 340 341 342 343 351 360 361 366 \
 372 383 392 393 398 404 415 424 425 430 436 )
c1108 ( 436 0 ) capacitor c=0.0335551f //x=79.18 //y=4.7
c1109 ( 430 0 ) capacitor c=0.0584472f //x=75.48 //y=4.7
c1110 ( 425 0 ) capacitor c=0.0273931f //x=75.48 //y=1.915
c1111 ( 424 0 ) capacitor c=0.0455604f //x=75.48 //y=2.08
c1112 ( 415 0 ) capacitor c=0.0333886f //x=59.94 //y=4.7
c1113 ( 404 0 ) capacitor c=0.0333886f //x=50.32 //y=4.7
c1114 ( 398 0 ) capacitor c=0.0589949f //x=46.62 //y=4.7
c1115 ( 393 0 ) capacitor c=0.0273931f //x=46.62 //y=1.915
c1116 ( 392 0 ) capacitor c=0.0455604f //x=46.62 //y=2.08
c1117 ( 383 0 ) capacitor c=0.0333886f //x=31.08 //y=4.7
c1118 ( 372 0 ) capacitor c=0.0335551f //x=21.46 //y=4.7
c1119 ( 366 0 ) capacitor c=0.058931f //x=17.76 //y=4.7
c1120 ( 361 0 ) capacitor c=0.0273931f //x=17.76 //y=1.915
c1121 ( 360 0 ) capacitor c=0.0455604f //x=17.76 //y=2.08
c1122 ( 351 0 ) capacitor c=0.0336203f //x=2.22 //y=4.7
c1123 ( 343 0 ) capacitor c=0.0245352f //x=79.515 //y=4.79
c1124 ( 342 0 ) capacitor c=0.0827272f //x=79.27 //y=1.915
c1125 ( 341 0 ) capacitor c=0.0170266f //x=79.27 //y=1.45
c1126 ( 340 0 ) capacitor c=0.018609f //x=79.27 //y=1.22
c1127 ( 339 0 ) capacitor c=0.0187309f //x=79.27 //y=0.91
c1128 ( 333 0 ) capacitor c=0.014725f //x=79.115 //y=1.375
c1129 ( 331 0 ) capacitor c=0.0146567f //x=79.115 //y=0.755
c1130 ( 330 0 ) capacitor c=0.0335408f //x=78.745 //y=1.22
c1131 ( 329 0 ) capacitor c=0.0173761f //x=78.745 //y=0.91
c1132 ( 328 0 ) capacitor c=0.0432517f //x=76 //y=1.26
c1133 ( 327 0 ) capacitor c=0.0200379f //x=76 //y=0.915
c1134 ( 324 0 ) capacitor c=0.0148873f //x=75.845 //y=1.415
c1135 ( 322 0 ) capacitor c=0.0157803f //x=75.845 //y=0.76
c1136 ( 317 0 ) capacitor c=0.0218028f //x=75.47 //y=1.57
c1137 ( 316 0 ) capacitor c=0.0207459f //x=75.47 //y=1.26
c1138 ( 315 0 ) capacitor c=0.0194308f //x=75.47 //y=0.915
c1139 ( 307 0 ) capacitor c=0.0246783f //x=60.275 //y=4.79
c1140 ( 306 0 ) capacitor c=0.0825033f //x=60.03 //y=1.915
c1141 ( 305 0 ) capacitor c=0.0170266f //x=60.03 //y=1.45
c1142 ( 304 0 ) capacitor c=0.018609f //x=60.03 //y=1.22
c1143 ( 303 0 ) capacitor c=0.0187309f //x=60.03 //y=0.91
c1144 ( 297 0 ) capacitor c=0.014725f //x=59.875 //y=1.375
c1145 ( 295 0 ) capacitor c=0.0146567f //x=59.875 //y=0.755
c1146 ( 294 0 ) capacitor c=0.0335408f //x=59.505 //y=1.22
c1147 ( 293 0 ) capacitor c=0.0173761f //x=59.505 //y=0.91
c1148 ( 288 0 ) capacitor c=0.0246783f //x=50.655 //y=4.79
c1149 ( 287 0 ) capacitor c=0.0825033f //x=50.41 //y=1.915
c1150 ( 286 0 ) capacitor c=0.0170266f //x=50.41 //y=1.45
c1151 ( 285 0 ) capacitor c=0.018609f //x=50.41 //y=1.22
c1152 ( 284 0 ) capacitor c=0.0187309f //x=50.41 //y=0.91
c1153 ( 278 0 ) capacitor c=0.014725f //x=50.255 //y=1.375
c1154 ( 276 0 ) capacitor c=0.0146567f //x=50.255 //y=0.755
c1155 ( 275 0 ) capacitor c=0.0335408f //x=49.885 //y=1.22
c1156 ( 274 0 ) capacitor c=0.0173761f //x=49.885 //y=0.91
c1157 ( 273 0 ) capacitor c=0.0432517f //x=47.14 //y=1.26
c1158 ( 272 0 ) capacitor c=0.0200379f //x=47.14 //y=0.915
c1159 ( 269 0 ) capacitor c=0.0148873f //x=46.985 //y=1.415
c1160 ( 267 0 ) capacitor c=0.0157803f //x=46.985 //y=0.76
c1161 ( 262 0 ) capacitor c=0.0218028f //x=46.61 //y=1.57
c1162 ( 261 0 ) capacitor c=0.0207459f //x=46.61 //y=1.26
c1163 ( 260 0 ) capacitor c=0.0194308f //x=46.61 //y=0.915
c1164 ( 252 0 ) capacitor c=0.0246783f //x=31.415 //y=4.79
c1165 ( 251 0 ) capacitor c=0.0825033f //x=31.17 //y=1.915
c1166 ( 250 0 ) capacitor c=0.0170266f //x=31.17 //y=1.45
c1167 ( 249 0 ) capacitor c=0.018609f //x=31.17 //y=1.22
c1168 ( 248 0 ) capacitor c=0.0187309f //x=31.17 //y=0.91
c1169 ( 242 0 ) capacitor c=0.014725f //x=31.015 //y=1.375
c1170 ( 240 0 ) capacitor c=0.0146567f //x=31.015 //y=0.755
c1171 ( 239 0 ) capacitor c=0.0335408f //x=30.645 //y=1.22
c1172 ( 238 0 ) capacitor c=0.0173761f //x=30.645 //y=0.91
c1173 ( 233 0 ) capacitor c=0.0245352f //x=21.795 //y=4.79
c1174 ( 232 0 ) capacitor c=0.0825033f //x=21.55 //y=1.915
c1175 ( 231 0 ) capacitor c=0.0170266f //x=21.55 //y=1.45
c1176 ( 230 0 ) capacitor c=0.018609f //x=21.55 //y=1.22
c1177 ( 229 0 ) capacitor c=0.0187309f //x=21.55 //y=0.91
c1178 ( 223 0 ) capacitor c=0.014725f //x=21.395 //y=1.375
c1179 ( 221 0 ) capacitor c=0.0146567f //x=21.395 //y=0.755
c1180 ( 220 0 ) capacitor c=0.0335408f //x=21.025 //y=1.22
c1181 ( 219 0 ) capacitor c=0.0173761f //x=21.025 //y=0.91
c1182 ( 218 0 ) capacitor c=0.0432517f //x=18.28 //y=1.26
c1183 ( 217 0 ) capacitor c=0.0200379f //x=18.28 //y=0.915
c1184 ( 214 0 ) capacitor c=0.0148873f //x=18.125 //y=1.415
c1185 ( 212 0 ) capacitor c=0.0157803f //x=18.125 //y=0.76
c1186 ( 207 0 ) capacitor c=0.0218028f //x=17.75 //y=1.57
c1187 ( 206 0 ) capacitor c=0.0207459f //x=17.75 //y=1.26
c1188 ( 205 0 ) capacitor c=0.0194308f //x=17.75 //y=0.915
c1189 ( 197 0 ) capacitor c=0.024933f //x=2.555 //y=4.79
c1190 ( 196 0 ) capacitor c=0.0826756f //x=2.31 //y=1.915
c1191 ( 195 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c1192 ( 194 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c1193 ( 193 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c1194 ( 187 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c1195 ( 185 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c1196 ( 184 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c1197 ( 183 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c1198 ( 182 0 ) capacitor c=0.110114f //x=79.59 //y=6.02
c1199 ( 181 0 ) capacitor c=0.11012f //x=79.15 //y=6.02
c1200 ( 180 0 ) capacitor c=0.158794f //x=75.66 //y=6.02
c1201 ( 179 0 ) capacitor c=0.11002f //x=75.22 //y=6.02
c1202 ( 178 0 ) capacitor c=0.109949f //x=60.35 //y=6.02
c1203 ( 177 0 ) capacitor c=0.109956f //x=59.91 //y=6.02
c1204 ( 176 0 ) capacitor c=0.109949f //x=50.73 //y=6.02
c1205 ( 175 0 ) capacitor c=0.109956f //x=50.29 //y=6.02
c1206 ( 174 0 ) capacitor c=0.158754f //x=46.8 //y=6.02
c1207 ( 173 0 ) capacitor c=0.109949f //x=46.36 //y=6.02
c1208 ( 172 0 ) capacitor c=0.109949f //x=31.49 //y=6.02
c1209 ( 171 0 ) capacitor c=0.109956f //x=31.05 //y=6.02
c1210 ( 170 0 ) capacitor c=0.110114f //x=21.87 //y=6.02
c1211 ( 169 0 ) capacitor c=0.11012f //x=21.43 //y=6.02
c1212 ( 168 0 ) capacitor c=0.158794f //x=17.94 //y=6.02
c1213 ( 167 0 ) capacitor c=0.110114f //x=17.5 //y=6.02
c1214 ( 166 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c1215 ( 165 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c1216 ( 147 0 ) capacitor c=0.0921679f //x=79.18 //y=2.08
c1217 ( 138 0 ) capacitor c=0.0818106f //x=75.48 //y=2.08
c1218 ( 127 0 ) capacitor c=0.0920722f //x=59.94 //y=2.08
c1219 ( 117 0 ) capacitor c=0.0898148f //x=50.32 //y=2.08
c1220 ( 108 0 ) capacitor c=0.0797966f //x=46.62 //y=2.08
c1221 ( 97 0 ) capacitor c=0.092949f //x=31.08 //y=2.08
c1222 ( 87 0 ) capacitor c=0.0915318f //x=21.46 //y=2.08
c1223 ( 78 0 ) capacitor c=0.081834f //x=17.76 //y=2.08
c1224 ( 65 0 ) capacitor c=0.100124f //x=2.22 //y=2.08
c1225 ( 16 0 ) capacitor c=0.00626813f //x=75.595 //y=2.22
c1226 ( 15 0 ) capacitor c=0.0896247f //x=79.065 //y=2.22
c1227 ( 14 0 ) capacitor c=0.00683472f //x=60.055 //y=2.22
c1228 ( 13 0 ) capacitor c=0.318477f //x=75.365 //y=2.22
c1229 ( 12 0 ) capacitor c=0.0059254f //x=50.435 //y=2.22
c1230 ( 11 0 ) capacitor c=0.196303f //x=59.825 //y=2.22
c1231 ( 10 0 ) capacitor c=0.00618148f //x=46.735 //y=2.22
c1232 ( 9 0 ) capacitor c=0.0804516f //x=50.205 //y=2.22
c1233 ( 8 0 ) capacitor c=0.00683472f //x=31.195 //y=2.22
c1234 ( 7 0 ) capacitor c=0.318477f //x=46.505 //y=2.22
c1235 ( 6 0 ) capacitor c=0.00601205f //x=21.575 //y=2.22
c1236 ( 5 0 ) capacitor c=0.20788f //x=30.965 //y=2.22
c1237 ( 4 0 ) capacitor c=0.00626813f //x=17.875 //y=2.22
c1238 ( 3 0 ) capacitor c=0.0805381f //x=21.345 //y=2.22
c1239 ( 2 0 ) capacitor c=0.0163048f //x=2.335 //y=2.22
c1240 ( 1 0 ) capacitor c=0.330466f //x=17.645 //y=2.22
r1241 (  438 439 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=79.18 //y=4.79 //x2=79.18 //y2=4.865
r1242 (  436 438 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=79.18 //y=4.7 //x2=79.18 //y2=4.79
r1243 (  424 425 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=75.48 //y=2.08 //x2=75.48 //y2=1.915
r1244 (  417 418 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=59.94 //y=4.79 //x2=59.94 //y2=4.865
r1245 (  415 417 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=59.94 //y=4.7 //x2=59.94 //y2=4.79
r1246 (  406 407 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=50.32 //y=4.79 //x2=50.32 //y2=4.865
r1247 (  404 406 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=50.32 //y=4.7 //x2=50.32 //y2=4.79
r1248 (  392 393 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=46.62 //y=2.08 //x2=46.62 //y2=1.915
r1249 (  385 386 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=31.08 //y=4.79 //x2=31.08 //y2=4.865
r1250 (  383 385 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=31.08 //y=4.7 //x2=31.08 //y2=4.79
r1251 (  374 375 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=21.46 //y=4.79 //x2=21.46 //y2=4.865
r1252 (  372 374 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=21.46 //y=4.7 //x2=21.46 //y2=4.79
r1253 (  360 361 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.76 //y=2.08 //x2=17.76 //y2=1.915
r1254 (  353 354 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r1255 (  351 353 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r1256 (  344 438 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=79.315 //y=4.79 //x2=79.18 //y2=4.79
r1257 (  343 345 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=79.515 //y=4.79 //x2=79.59 //y2=4.865
r1258 (  343 344 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=79.515 //y=4.79 //x2=79.315 //y2=4.79
r1259 (  342 443 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=79.27 //y=1.915 //x2=79.195 //y2=2.08
r1260 (  341 441 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=79.27 //y=1.45 //x2=79.23 //y2=1.375
r1261 (  341 342 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=79.27 //y=1.45 //x2=79.27 //y2=1.915
r1262 (  340 441 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.27 //y=1.22 //x2=79.23 //y2=1.375
r1263 (  339 440 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.27 //y=0.91 //x2=79.23 //y2=0.755
r1264 (  339 340 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=79.27 //y=0.91 //x2=79.27 //y2=1.22
r1265 (  334 434 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.9 //y=1.375 //x2=78.785 //y2=1.375
r1266 (  333 441 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=79.115 //y=1.375 //x2=79.23 //y2=1.375
r1267 (  332 433 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.9 //y=0.755 //x2=78.785 //y2=0.755
r1268 (  331 440 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=79.115 //y=0.755 //x2=79.23 //y2=0.755
r1269 (  331 332 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=79.115 //y=0.755 //x2=78.9 //y2=0.755
r1270 (  330 434 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.745 //y=1.22 //x2=78.785 //y2=1.375
r1271 (  329 433 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.745 //y=0.91 //x2=78.785 //y2=0.755
r1272 (  329 330 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=78.745 //y=0.91 //x2=78.745 //y2=1.22
r1273 (  328 432 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=76 //y=1.26 //x2=75.96 //y2=1.415
r1274 (  327 431 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=76 //y=0.915 //x2=75.96 //y2=0.76
r1275 (  327 328 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=76 //y=0.915 //x2=76 //y2=1.26
r1276 (  325 428 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.625 //y=1.415 //x2=75.51 //y2=1.415
r1277 (  324 432 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.845 //y=1.415 //x2=75.96 //y2=1.415
r1278 (  323 427 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.625 //y=0.76 //x2=75.51 //y2=0.76
r1279 (  322 431 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.845 //y=0.76 //x2=75.96 //y2=0.76
r1280 (  322 323 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=75.845 //y=0.76 //x2=75.625 //y2=0.76
r1281 (  319 430 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=75.66 //y=4.865 //x2=75.48 //y2=4.7
r1282 (  317 428 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.47 //y=1.57 //x2=75.51 //y2=1.415
r1283 (  317 425 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.47 //y=1.57 //x2=75.47 //y2=1.915
r1284 (  316 428 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.47 //y=1.26 //x2=75.51 //y2=1.415
r1285 (  315 427 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.47 //y=0.915 //x2=75.51 //y2=0.76
r1286 (  315 316 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.47 //y=0.915 //x2=75.47 //y2=1.26
r1287 (  312 430 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=75.22 //y=4.865 //x2=75.48 //y2=4.7
r1288 (  308 417 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=60.075 //y=4.79 //x2=59.94 //y2=4.79
r1289 (  307 309 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=60.275 //y=4.79 //x2=60.35 //y2=4.865
r1290 (  307 308 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=60.275 //y=4.79 //x2=60.075 //y2=4.79
r1291 (  306 422 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=60.03 //y=1.915 //x2=59.955 //y2=2.08
r1292 (  305 420 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=60.03 //y=1.45 //x2=59.99 //y2=1.375
r1293 (  305 306 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=60.03 //y=1.45 //x2=60.03 //y2=1.915
r1294 (  304 420 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.03 //y=1.22 //x2=59.99 //y2=1.375
r1295 (  303 419 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.03 //y=0.91 //x2=59.99 //y2=0.755
r1296 (  303 304 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=60.03 //y=0.91 //x2=60.03 //y2=1.22
r1297 (  298 413 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.66 //y=1.375 //x2=59.545 //y2=1.375
r1298 (  297 420 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.875 //y=1.375 //x2=59.99 //y2=1.375
r1299 (  296 412 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.66 //y=0.755 //x2=59.545 //y2=0.755
r1300 (  295 419 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.875 //y=0.755 //x2=59.99 //y2=0.755
r1301 (  295 296 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=59.875 //y=0.755 //x2=59.66 //y2=0.755
r1302 (  294 413 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.505 //y=1.22 //x2=59.545 //y2=1.375
r1303 (  293 412 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.505 //y=0.91 //x2=59.545 //y2=0.755
r1304 (  293 294 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=59.505 //y=0.91 //x2=59.505 //y2=1.22
r1305 (  289 406 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=50.455 //y=4.79 //x2=50.32 //y2=4.79
r1306 (  288 290 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=50.655 //y=4.79 //x2=50.73 //y2=4.865
r1307 (  288 289 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=50.655 //y=4.79 //x2=50.455 //y2=4.79
r1308 (  287 411 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=50.41 //y=1.915 //x2=50.335 //y2=2.08
r1309 (  286 409 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=50.41 //y=1.45 //x2=50.37 //y2=1.375
r1310 (  286 287 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=50.41 //y=1.45 //x2=50.41 //y2=1.915
r1311 (  285 409 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.41 //y=1.22 //x2=50.37 //y2=1.375
r1312 (  284 408 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.41 //y=0.91 //x2=50.37 //y2=0.755
r1313 (  284 285 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=50.41 //y=0.91 //x2=50.41 //y2=1.22
r1314 (  279 402 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.04 //y=1.375 //x2=49.925 //y2=1.375
r1315 (  278 409 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.255 //y=1.375 //x2=50.37 //y2=1.375
r1316 (  277 401 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.04 //y=0.755 //x2=49.925 //y2=0.755
r1317 (  276 408 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.255 //y=0.755 //x2=50.37 //y2=0.755
r1318 (  276 277 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=50.255 //y=0.755 //x2=50.04 //y2=0.755
r1319 (  275 402 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.885 //y=1.22 //x2=49.925 //y2=1.375
r1320 (  274 401 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.885 //y=0.91 //x2=49.925 //y2=0.755
r1321 (  274 275 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=49.885 //y=0.91 //x2=49.885 //y2=1.22
r1322 (  273 400 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.14 //y=1.26 //x2=47.1 //y2=1.415
r1323 (  272 399 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.14 //y=0.915 //x2=47.1 //y2=0.76
r1324 (  272 273 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=47.14 //y=0.915 //x2=47.14 //y2=1.26
r1325 (  270 396 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.765 //y=1.415 //x2=46.65 //y2=1.415
r1326 (  269 400 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.985 //y=1.415 //x2=47.1 //y2=1.415
r1327 (  268 395 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.765 //y=0.76 //x2=46.65 //y2=0.76
r1328 (  267 399 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.985 //y=0.76 //x2=47.1 //y2=0.76
r1329 (  267 268 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=46.985 //y=0.76 //x2=46.765 //y2=0.76
r1330 (  264 398 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=46.8 //y=4.865 //x2=46.62 //y2=4.7
r1331 (  262 396 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.61 //y=1.57 //x2=46.65 //y2=1.415
r1332 (  262 393 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=46.61 //y=1.57 //x2=46.61 //y2=1.915
r1333 (  261 396 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.61 //y=1.26 //x2=46.65 //y2=1.415
r1334 (  260 395 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.61 //y=0.915 //x2=46.65 //y2=0.76
r1335 (  260 261 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=46.61 //y=0.915 //x2=46.61 //y2=1.26
r1336 (  257 398 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=46.36 //y=4.865 //x2=46.62 //y2=4.7
r1337 (  253 385 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=31.215 //y=4.79 //x2=31.08 //y2=4.79
r1338 (  252 254 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=31.415 //y=4.79 //x2=31.49 //y2=4.865
r1339 (  252 253 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=31.415 //y=4.79 //x2=31.215 //y2=4.79
r1340 (  251 390 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=31.17 //y=1.915 //x2=31.095 //y2=2.08
r1341 (  250 388 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=31.17 //y=1.45 //x2=31.13 //y2=1.375
r1342 (  250 251 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=31.17 //y=1.45 //x2=31.17 //y2=1.915
r1343 (  249 388 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.17 //y=1.22 //x2=31.13 //y2=1.375
r1344 (  248 387 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.17 //y=0.91 //x2=31.13 //y2=0.755
r1345 (  248 249 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=31.17 //y=0.91 //x2=31.17 //y2=1.22
r1346 (  243 381 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.8 //y=1.375 //x2=30.685 //y2=1.375
r1347 (  242 388 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.015 //y=1.375 //x2=31.13 //y2=1.375
r1348 (  241 380 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.8 //y=0.755 //x2=30.685 //y2=0.755
r1349 (  240 387 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.015 //y=0.755 //x2=31.13 //y2=0.755
r1350 (  240 241 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=31.015 //y=0.755 //x2=30.8 //y2=0.755
r1351 (  239 381 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.645 //y=1.22 //x2=30.685 //y2=1.375
r1352 (  238 380 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.645 //y=0.91 //x2=30.685 //y2=0.755
r1353 (  238 239 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=30.645 //y=0.91 //x2=30.645 //y2=1.22
r1354 (  234 374 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=21.595 //y=4.79 //x2=21.46 //y2=4.79
r1355 (  233 235 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.795 //y=4.79 //x2=21.87 //y2=4.865
r1356 (  233 234 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=21.795 //y=4.79 //x2=21.595 //y2=4.79
r1357 (  232 379 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.915 //x2=21.475 //y2=2.08
r1358 (  231 377 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.45 //x2=21.51 //y2=1.375
r1359 (  231 232 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.45 //x2=21.55 //y2=1.915
r1360 (  230 377 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.22 //x2=21.51 //y2=1.375
r1361 (  229 376 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.91 //x2=21.51 //y2=0.755
r1362 (  229 230 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.91 //x2=21.55 //y2=1.22
r1363 (  224 370 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.18 //y=1.375 //x2=21.065 //y2=1.375
r1364 (  223 377 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.395 //y=1.375 //x2=21.51 //y2=1.375
r1365 (  222 369 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.18 //y=0.755 //x2=21.065 //y2=0.755
r1366 (  221 376 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.755 //x2=21.51 //y2=0.755
r1367 (  221 222 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.755 //x2=21.18 //y2=0.755
r1368 (  220 370 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.025 //y=1.22 //x2=21.065 //y2=1.375
r1369 (  219 369 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.025 //y=0.91 //x2=21.065 //y2=0.755
r1370 (  219 220 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.025 //y=0.91 //x2=21.025 //y2=1.22
r1371 (  218 368 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.28 //y=1.26 //x2=18.24 //y2=1.415
r1372 (  217 367 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.28 //y=0.915 //x2=18.24 //y2=0.76
r1373 (  217 218 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.28 //y=0.915 //x2=18.28 //y2=1.26
r1374 (  215 364 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.905 //y=1.415 //x2=17.79 //y2=1.415
r1375 (  214 368 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.125 //y=1.415 //x2=18.24 //y2=1.415
r1376 (  213 363 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.905 //y=0.76 //x2=17.79 //y2=0.76
r1377 (  212 367 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.125 //y=0.76 //x2=18.24 //y2=0.76
r1378 (  212 213 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.125 //y=0.76 //x2=17.905 //y2=0.76
r1379 (  209 366 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=17.94 //y=4.865 //x2=17.76 //y2=4.7
r1380 (  207 364 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.57 //x2=17.79 //y2=1.415
r1381 (  207 361 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.57 //x2=17.75 //y2=1.915
r1382 (  206 364 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.26 //x2=17.79 //y2=1.415
r1383 (  205 363 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=0.915 //x2=17.79 //y2=0.76
r1384 (  205 206 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.75 //y=0.915 //x2=17.75 //y2=1.26
r1385 (  202 366 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=17.5 //y=4.865 //x2=17.76 //y2=4.7
r1386 (  198 353 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r1387 (  197 199 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r1388 (  197 198 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r1389 (  196 358 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r1390 (  195 356 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r1391 (  195 196 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r1392 (  194 356 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r1393 (  193 355 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r1394 (  193 194 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r1395 (  188 349 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r1396 (  187 356 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r1397 (  186 348 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r1398 (  185 355 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r1399 (  185 186 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r1400 (  184 349 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r1401 (  183 348 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r1402 (  183 184 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r1403 (  182 345 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=79.59 //y=6.02 //x2=79.59 //y2=4.865
r1404 (  181 439 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=79.15 //y=6.02 //x2=79.15 //y2=4.865
r1405 (  180 319 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.66 //y=6.02 //x2=75.66 //y2=4.865
r1406 (  179 312 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.22 //y=6.02 //x2=75.22 //y2=4.865
r1407 (  178 309 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.35 //y=6.02 //x2=60.35 //y2=4.865
r1408 (  177 418 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.91 //y=6.02 //x2=59.91 //y2=4.865
r1409 (  176 290 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.73 //y=6.02 //x2=50.73 //y2=4.865
r1410 (  175 407 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.29 //y=6.02 //x2=50.29 //y2=4.865
r1411 (  174 264 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.8 //y=6.02 //x2=46.8 //y2=4.865
r1412 (  173 257 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.36 //y=6.02 //x2=46.36 //y2=4.865
r1413 (  172 254 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.49 //y=6.02 //x2=31.49 //y2=4.865
r1414 (  171 386 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.05 //y=6.02 //x2=31.05 //y2=4.865
r1415 (  170 235 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.87 //y=6.02 //x2=21.87 //y2=4.865
r1416 (  169 375 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.43 //y=6.02 //x2=21.43 //y2=4.865
r1417 (  168 209 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.94 //y=6.02 //x2=17.94 //y2=4.865
r1418 (  167 202 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.5 //y=6.02 //x2=17.5 //y2=4.865
r1419 (  166 199 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r1420 (  165 354 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r1421 (  164 333 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=79.007 //y=1.375 //x2=79.115 //y2=1.375
r1422 (  164 334 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=79.007 //y=1.375 //x2=78.9 //y2=1.375
r1423 (  163 324 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.735 //y=1.415 //x2=75.845 //y2=1.415
r1424 (  163 325 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.735 //y=1.415 //x2=75.625 //y2=1.415
r1425 (  162 297 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=59.767 //y=1.375 //x2=59.875 //y2=1.375
r1426 (  162 298 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=59.767 //y=1.375 //x2=59.66 //y2=1.375
r1427 (  161 278 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=50.147 //y=1.375 //x2=50.255 //y2=1.375
r1428 (  161 279 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=50.147 //y=1.375 //x2=50.04 //y2=1.375
r1429 (  160 269 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=46.875 //y=1.415 //x2=46.985 //y2=1.415
r1430 (  160 270 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=46.875 //y=1.415 //x2=46.765 //y2=1.415
r1431 (  159 242 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=30.907 //y=1.375 //x2=31.015 //y2=1.375
r1432 (  159 243 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=30.907 //y=1.375 //x2=30.8 //y2=1.375
r1433 (  158 223 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=21.287 //y=1.375 //x2=21.395 //y2=1.375
r1434 (  158 224 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=21.287 //y=1.375 //x2=21.18 //y2=1.375
r1435 (  157 214 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.015 //y=1.415 //x2=18.125 //y2=1.415
r1436 (  157 215 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.015 //y=1.415 //x2=17.905 //y2=1.415
r1437 (  156 187 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r1438 (  156 188 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r1439 (  154 436 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.18 //y=4.7 //x2=79.18 //y2=4.7
r1440 (  147 443 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.18 //y=2.08 //x2=79.18 //y2=2.08
r1441 (  144 430 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.48 //y=4.7 //x2=75.48 //y2=4.7
r1442 (  138 424 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.48 //y=2.08 //x2=75.48 //y2=2.08
r1443 (  135 415 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.94 //y=4.7 //x2=59.94 //y2=4.7
r1444 (  127 422 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.94 //y=2.08 //x2=59.94 //y2=2.08
r1445 (  124 404 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.32 //y=4.7 //x2=50.32 //y2=4.7
r1446 (  117 411 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.32 //y=2.08 //x2=50.32 //y2=2.08
r1447 (  114 398 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.62 //y=4.7 //x2=46.62 //y2=4.7
r1448 (  108 392 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.62 //y=2.08 //x2=46.62 //y2=2.08
r1449 (  105 383 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.08 //y=4.7 //x2=31.08 //y2=4.7
r1450 (  97 390 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.08 //y=2.08 //x2=31.08 //y2=2.08
r1451 (  94 372 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=4.7 //x2=21.46 //y2=4.7
r1452 (  87 379 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=2.08 //x2=21.46 //y2=2.08
r1453 (  84 366 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=4.7 //x2=17.76 //y2=4.7
r1454 (  78 360 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=2.08 //x2=17.76 //y2=2.08
r1455 (  75 351 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r1456 (  65 358 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r1457 (  63 154 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=79.18 //y=3.33 //x2=79.18 //y2=4.7
r1458 (  62 63 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=79.18 //y=2.59 //x2=79.18 //y2=3.33
r1459 (  61 62 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=79.18 //y=2.22 //x2=79.18 //y2=2.59
r1460 (  61 147 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=79.18 //y=2.22 //x2=79.18 //y2=2.08
r1461 (  60 144 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=75.48 //y=2.59 //x2=75.48 //y2=4.7
r1462 (  59 60 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=75.48 //y=2.22 //x2=75.48 //y2=2.59
r1463 (  59 138 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=75.48 //y=2.22 //x2=75.48 //y2=2.08
r1464 (  58 135 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=59.94 //y=4.07 //x2=59.94 //y2=4.7
r1465 (  57 58 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=59.94 //y=3.33 //x2=59.94 //y2=4.07
r1466 (  56 57 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=59.94 //y=2.59 //x2=59.94 //y2=3.33
r1467 (  55 56 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=59.94 //y=2.22 //x2=59.94 //y2=2.59
r1468 (  55 127 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=59.94 //y=2.22 //x2=59.94 //y2=2.08
r1469 (  54 124 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=50.32 //y=3.33 //x2=50.32 //y2=4.7
r1470 (  53 54 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=50.32 //y=2.59 //x2=50.32 //y2=3.33
r1471 (  52 53 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=50.32 //y=2.22 //x2=50.32 //y2=2.59
r1472 (  52 117 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=50.32 //y=2.22 //x2=50.32 //y2=2.08
r1473 (  51 114 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=46.62 //y=2.59 //x2=46.62 //y2=4.7
r1474 (  50 51 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=46.62 //y=2.22 //x2=46.62 //y2=2.59
r1475 (  50 108 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=46.62 //y=2.22 //x2=46.62 //y2=2.08
r1476 (  49 105 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li \
 //thickness=0.1 //x=31.08 //y=3.7 //x2=31.08 //y2=4.7
r1477 (  48 49 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=31.08 //y=3.33 //x2=31.08 //y2=3.7
r1478 (  47 48 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=31.08 //y=2.59 //x2=31.08 //y2=3.33
r1479 (  46 47 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=31.08 //y=2.22 //x2=31.08 //y2=2.59
r1480 (  46 97 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=31.08 //y=2.22 //x2=31.08 //y2=2.08
r1481 (  45 94 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=3.33 //x2=21.46 //y2=4.7
r1482 (  44 45 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.59 //x2=21.46 //y2=3.33
r1483 (  43 44 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.22 //x2=21.46 //y2=2.59
r1484 (  43 87 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.22 //x2=21.46 //y2=2.08
r1485 (  42 84 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.59 //x2=17.76 //y2=4.7
r1486 (  41 42 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.22 //x2=17.76 //y2=2.59
r1487 (  41 78 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.22 //x2=17.76 //y2=2.08
r1488 (  40 75 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=2.22 //y=4.44 //x2=2.22 //y2=4.7
r1489 (  39 40 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.7 //x2=2.22 //y2=4.44
r1490 (  38 39 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.33 //x2=2.22 //y2=3.7
r1491 (  37 38 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.96 //x2=2.22 //y2=3.33
r1492 (  36 37 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.59 //x2=2.22 //y2=2.96
r1493 (  35 36 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.22 //x2=2.22 //y2=2.59
r1494 (  35 65 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.22 //x2=2.22 //y2=2.08
r1495 (  34 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.18 //y=2.22 //x2=79.18 //y2=2.22
r1496 (  32 59 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.48 //y=2.22 //x2=75.48 //y2=2.22
r1497 (  30 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=59.94 //y=2.22 //x2=59.94 //y2=2.22
r1498 (  28 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=50.32 //y=2.22 //x2=50.32 //y2=2.22
r1499 (  26 50 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=46.62 //y=2.22 //x2=46.62 //y2=2.22
r1500 (  24 46 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=31.08 //y=2.22 //x2=31.08 //y2=2.22
r1501 (  22 43 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.46 //y=2.22 //x2=21.46 //y2=2.22
r1502 (  20 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.76 //y=2.22 //x2=17.76 //y2=2.22
r1503 (  18 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.22 //y=2.22 //x2=2.22 //y2=2.22
r1504 (  16 32 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.595 //y=2.22 //x2=75.48 //y2=2.22
r1505 (  15 34 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.065 //y=2.22 //x2=79.18 //y2=2.22
r1506 (  15 16 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=79.065 //y=2.22 //x2=75.595 //y2=2.22
r1507 (  14 30 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.055 //y=2.22 //x2=59.94 //y2=2.22
r1508 (  13 32 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.365 //y=2.22 //x2=75.48 //y2=2.22
r1509 (  13 14 ) resistor r=14.6088 //w=0.131 //l=15.31 //layer=m1 \
 //thickness=0.36 //x=75.365 //y=2.22 //x2=60.055 //y2=2.22
r1510 (  12 28 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.435 //y=2.22 //x2=50.32 //y2=2.22
r1511 (  11 30 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=59.825 //y=2.22 //x2=59.94 //y2=2.22
r1512 (  11 12 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=59.825 //y=2.22 //x2=50.435 //y2=2.22
r1513 (  10 26 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=46.735 //y=2.22 //x2=46.62 //y2=2.22
r1514 (  9 28 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.205 //y=2.22 //x2=50.32 //y2=2.22
r1515 (  9 10 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=50.205 //y=2.22 //x2=46.735 //y2=2.22
r1516 (  8 24 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.195 //y=2.22 //x2=31.08 //y2=2.22
r1517 (  7 26 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=46.505 //y=2.22 //x2=46.62 //y2=2.22
r1518 (  7 8 ) resistor r=14.6088 //w=0.131 //l=15.31 //layer=m1 \
 //thickness=0.36 //x=46.505 //y=2.22 //x2=31.195 //y2=2.22
r1519 (  6 22 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.575 //y=2.22 //x2=21.46 //y2=2.22
r1520 (  5 24 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=30.965 //y=2.22 //x2=31.08 //y2=2.22
r1521 (  5 6 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=30.965 //y=2.22 //x2=21.575 //y2=2.22
r1522 (  4 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.875 //y=2.22 //x2=17.76 //y2=2.22
r1523 (  3 22 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=2.22 //x2=21.46 //y2=2.22
r1524 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=2.22 //x2=17.875 //y2=2.22
r1525 (  2 18 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.335 //y=2.22 //x2=2.22 //y2=2.22
r1526 (  1 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.645 //y=2.22 //x2=17.76 //y2=2.22
r1527 (  1 2 ) resistor r=14.6088 //w=0.131 //l=15.31 //layer=m1 \
 //thickness=0.36 //x=17.645 //y=2.22 //x2=2.335 //y2=2.22
ends PM_TMRDFFSNRNQNX1\%RN

subckt PM_TMRDFFSNRNQNX1\%SN ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 31 \
 33 42 51 60 68 77 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 \
 103 104 106 112 113 114 115 116 121 122 123 125 131 132 133 134 135 140 141 \
 142 144 150 151 152 153 154 159 160 161 163 169 170 171 172 173 178 179 180 \
 182 188 189 190 191 192 197 198 199 201 207 208 209 210 211 219 230 241 252 \
 263 274 )
c699 ( 274 0 ) capacitor c=0.0335551f //x=83.99 //y=4.7
c700 ( 263 0 ) capacitor c=0.0333886f //x=69.56 //y=4.7
c701 ( 252 0 ) capacitor c=0.0333886f //x=55.13 //y=4.7
c702 ( 241 0 ) capacitor c=0.0333886f //x=40.7 //y=4.7
c703 ( 230 0 ) capacitor c=0.0333886f //x=26.27 //y=4.7
c704 ( 219 0 ) capacitor c=0.0335551f //x=11.84 //y=4.7
c705 ( 211 0 ) capacitor c=0.0245352f //x=84.325 //y=4.79
c706 ( 210 0 ) capacitor c=0.0825763f //x=84.08 //y=1.915
c707 ( 209 0 ) capacitor c=0.0170266f //x=84.08 //y=1.45
c708 ( 208 0 ) capacitor c=0.018609f //x=84.08 //y=1.22
c709 ( 207 0 ) capacitor c=0.0187309f //x=84.08 //y=0.91
c710 ( 201 0 ) capacitor c=0.014725f //x=83.925 //y=1.375
c711 ( 199 0 ) capacitor c=0.0146567f //x=83.925 //y=0.755
c712 ( 198 0 ) capacitor c=0.0335408f //x=83.555 //y=1.22
c713 ( 197 0 ) capacitor c=0.0173761f //x=83.555 //y=0.91
c714 ( 192 0 ) capacitor c=0.0246783f //x=69.895 //y=4.79
c715 ( 191 0 ) capacitor c=0.0825763f //x=69.65 //y=1.915
c716 ( 190 0 ) capacitor c=0.0170266f //x=69.65 //y=1.45
c717 ( 189 0 ) capacitor c=0.018609f //x=69.65 //y=1.22
c718 ( 188 0 ) capacitor c=0.0187309f //x=69.65 //y=0.91
c719 ( 182 0 ) capacitor c=0.014725f //x=69.495 //y=1.375
c720 ( 180 0 ) capacitor c=0.0146567f //x=69.495 //y=0.755
c721 ( 179 0 ) capacitor c=0.0335408f //x=69.125 //y=1.22
c722 ( 178 0 ) capacitor c=0.0173761f //x=69.125 //y=0.91
c723 ( 173 0 ) capacitor c=0.0246783f //x=55.465 //y=4.79
c724 ( 172 0 ) capacitor c=0.0825763f //x=55.22 //y=1.915
c725 ( 171 0 ) capacitor c=0.0170266f //x=55.22 //y=1.45
c726 ( 170 0 ) capacitor c=0.018609f //x=55.22 //y=1.22
c727 ( 169 0 ) capacitor c=0.0187309f //x=55.22 //y=0.91
c728 ( 163 0 ) capacitor c=0.014725f //x=55.065 //y=1.375
c729 ( 161 0 ) capacitor c=0.0146567f //x=55.065 //y=0.755
c730 ( 160 0 ) capacitor c=0.0335408f //x=54.695 //y=1.22
c731 ( 159 0 ) capacitor c=0.0173761f //x=54.695 //y=0.91
c732 ( 154 0 ) capacitor c=0.0246783f //x=41.035 //y=4.79
c733 ( 153 0 ) capacitor c=0.0825763f //x=40.79 //y=1.915
c734 ( 152 0 ) capacitor c=0.0170266f //x=40.79 //y=1.45
c735 ( 151 0 ) capacitor c=0.018609f //x=40.79 //y=1.22
c736 ( 150 0 ) capacitor c=0.0187309f //x=40.79 //y=0.91
c737 ( 144 0 ) capacitor c=0.014725f //x=40.635 //y=1.375
c738 ( 142 0 ) capacitor c=0.0146567f //x=40.635 //y=0.755
c739 ( 141 0 ) capacitor c=0.0335408f //x=40.265 //y=1.22
c740 ( 140 0 ) capacitor c=0.0173761f //x=40.265 //y=0.91
c741 ( 135 0 ) capacitor c=0.0246783f //x=26.605 //y=4.79
c742 ( 134 0 ) capacitor c=0.0825763f //x=26.36 //y=1.915
c743 ( 133 0 ) capacitor c=0.0170266f //x=26.36 //y=1.45
c744 ( 132 0 ) capacitor c=0.018609f //x=26.36 //y=1.22
c745 ( 131 0 ) capacitor c=0.0187309f //x=26.36 //y=0.91
c746 ( 125 0 ) capacitor c=0.014725f //x=26.205 //y=1.375
c747 ( 123 0 ) capacitor c=0.0146567f //x=26.205 //y=0.755
c748 ( 122 0 ) capacitor c=0.0335408f //x=25.835 //y=1.22
c749 ( 121 0 ) capacitor c=0.0173761f //x=25.835 //y=0.91
c750 ( 116 0 ) capacitor c=0.0245352f //x=12.175 //y=4.79
c751 ( 115 0 ) capacitor c=0.0825763f //x=11.93 //y=1.915
c752 ( 114 0 ) capacitor c=0.0170266f //x=11.93 //y=1.45
c753 ( 113 0 ) capacitor c=0.018609f //x=11.93 //y=1.22
c754 ( 112 0 ) capacitor c=0.0187309f //x=11.93 //y=0.91
c755 ( 106 0 ) capacitor c=0.014725f //x=11.775 //y=1.375
c756 ( 104 0 ) capacitor c=0.0146567f //x=11.775 //y=0.755
c757 ( 103 0 ) capacitor c=0.0335408f //x=11.405 //y=1.22
c758 ( 102 0 ) capacitor c=0.0173761f //x=11.405 //y=0.91
c759 ( 101 0 ) capacitor c=0.110114f //x=84.4 //y=6.02
c760 ( 100 0 ) capacitor c=0.11012f //x=83.96 //y=6.02
c761 ( 99 0 ) capacitor c=0.109949f //x=69.97 //y=6.02
c762 ( 98 0 ) capacitor c=0.109956f //x=69.53 //y=6.02
c763 ( 97 0 ) capacitor c=0.109949f //x=55.54 //y=6.02
c764 ( 96 0 ) capacitor c=0.109956f //x=55.1 //y=6.02
c765 ( 95 0 ) capacitor c=0.109949f //x=41.11 //y=6.02
c766 ( 94 0 ) capacitor c=0.109956f //x=40.67 //y=6.02
c767 ( 93 0 ) capacitor c=0.109949f //x=26.68 //y=6.02
c768 ( 92 0 ) capacitor c=0.109956f //x=26.24 //y=6.02
c769 ( 91 0 ) capacitor c=0.110114f //x=12.25 //y=6.02
c770 ( 90 0 ) capacitor c=0.11012f //x=11.81 //y=6.02
c771 ( 77 0 ) capacitor c=0.0905889f //x=83.99 //y=2.08
c772 ( 68 0 ) capacitor c=0.0877968f //x=69.56 //y=2.08
c773 ( 60 0 ) capacitor c=0.0858298f //x=55.13 //y=2.08
c774 ( 51 0 ) capacitor c=0.0877968f //x=40.7 //y=2.08
c775 ( 42 0 ) capacitor c=0.0881699f //x=26.27 //y=2.08
c776 ( 33 0 ) capacitor c=0.0895139f //x=11.84 //y=2.08
c777 ( 10 0 ) capacitor c=0.00568147f //x=69.675 //y=2.96
c778 ( 9 0 ) capacitor c=0.263037f //x=83.875 //y=2.96
c779 ( 8 0 ) capacitor c=0.00539919f //x=55.245 //y=2.96
c780 ( 7 0 ) capacitor c=0.22725f //x=69.445 //y=2.96
c781 ( 6 0 ) capacitor c=0.00568147f //x=40.815 //y=2.96
c782 ( 5 0 ) capacitor c=0.228822f //x=55.015 //y=2.96
c783 ( 4 0 ) capacitor c=0.00568147f //x=26.385 //y=2.96
c784 ( 3 0 ) capacitor c=0.242055f //x=40.585 //y=2.96
c785 ( 2 0 ) capacitor c=0.0141295f //x=11.955 //y=2.96
c786 ( 1 0 ) capacitor c=0.231676f //x=26.155 //y=2.96
r787 (  276 277 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=83.99 //y=4.79 //x2=83.99 //y2=4.865
r788 (  274 276 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=83.99 //y=4.7 //x2=83.99 //y2=4.79
r789 (  265 266 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=69.56 //y=4.79 //x2=69.56 //y2=4.865
r790 (  263 265 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=69.56 //y=4.7 //x2=69.56 //y2=4.79
r791 (  254 255 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=55.13 //y=4.79 //x2=55.13 //y2=4.865
r792 (  252 254 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=55.13 //y=4.7 //x2=55.13 //y2=4.79
r793 (  243 244 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=40.7 //y=4.79 //x2=40.7 //y2=4.865
r794 (  241 243 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=40.7 //y=4.7 //x2=40.7 //y2=4.79
r795 (  232 233 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=26.27 //y=4.79 //x2=26.27 //y2=4.865
r796 (  230 232 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=26.27 //y=4.7 //x2=26.27 //y2=4.79
r797 (  221 222 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=11.84 //y=4.79 //x2=11.84 //y2=4.865
r798 (  219 221 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=11.84 //y=4.7 //x2=11.84 //y2=4.79
r799 (  212 276 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=84.125 //y=4.79 //x2=83.99 //y2=4.79
r800 (  211 213 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=84.325 //y=4.79 //x2=84.4 //y2=4.865
r801 (  211 212 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=84.325 //y=4.79 //x2=84.125 //y2=4.79
r802 (  210 281 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=84.08 //y=1.915 //x2=84.005 //y2=2.08
r803 (  209 279 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=84.08 //y=1.45 //x2=84.04 //y2=1.375
r804 (  209 210 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=84.08 //y=1.45 //x2=84.08 //y2=1.915
r805 (  208 279 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=84.08 //y=1.22 //x2=84.04 //y2=1.375
r806 (  207 278 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=84.08 //y=0.91 //x2=84.04 //y2=0.755
r807 (  207 208 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=84.08 //y=0.91 //x2=84.08 //y2=1.22
r808 (  202 272 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.71 //y=1.375 //x2=83.595 //y2=1.375
r809 (  201 279 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.925 //y=1.375 //x2=84.04 //y2=1.375
r810 (  200 271 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.71 //y=0.755 //x2=83.595 //y2=0.755
r811 (  199 278 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.925 //y=0.755 //x2=84.04 //y2=0.755
r812 (  199 200 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=83.925 //y=0.755 //x2=83.71 //y2=0.755
r813 (  198 272 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.555 //y=1.22 //x2=83.595 //y2=1.375
r814 (  197 271 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.555 //y=0.91 //x2=83.595 //y2=0.755
r815 (  197 198 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=83.555 //y=0.91 //x2=83.555 //y2=1.22
r816 (  193 265 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=69.695 //y=4.79 //x2=69.56 //y2=4.79
r817 (  192 194 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=69.895 //y=4.79 //x2=69.97 //y2=4.865
r818 (  192 193 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=69.895 //y=4.79 //x2=69.695 //y2=4.79
r819 (  191 270 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=69.65 //y=1.915 //x2=69.575 //y2=2.08
r820 (  190 268 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=69.65 //y=1.45 //x2=69.61 //y2=1.375
r821 (  190 191 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=69.65 //y=1.45 //x2=69.65 //y2=1.915
r822 (  189 268 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.65 //y=1.22 //x2=69.61 //y2=1.375
r823 (  188 267 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.65 //y=0.91 //x2=69.61 //y2=0.755
r824 (  188 189 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=69.65 //y=0.91 //x2=69.65 //y2=1.22
r825 (  183 261 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.28 //y=1.375 //x2=69.165 //y2=1.375
r826 (  182 268 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.495 //y=1.375 //x2=69.61 //y2=1.375
r827 (  181 260 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.28 //y=0.755 //x2=69.165 //y2=0.755
r828 (  180 267 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.495 //y=0.755 //x2=69.61 //y2=0.755
r829 (  180 181 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=69.495 //y=0.755 //x2=69.28 //y2=0.755
r830 (  179 261 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.125 //y=1.22 //x2=69.165 //y2=1.375
r831 (  178 260 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.125 //y=0.91 //x2=69.165 //y2=0.755
r832 (  178 179 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=69.125 //y=0.91 //x2=69.125 //y2=1.22
r833 (  174 254 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=55.265 //y=4.79 //x2=55.13 //y2=4.79
r834 (  173 175 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=55.465 //y=4.79 //x2=55.54 //y2=4.865
r835 (  173 174 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=55.465 //y=4.79 //x2=55.265 //y2=4.79
r836 (  172 259 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=55.22 //y=1.915 //x2=55.145 //y2=2.08
r837 (  171 257 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=55.22 //y=1.45 //x2=55.18 //y2=1.375
r838 (  171 172 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=55.22 //y=1.45 //x2=55.22 //y2=1.915
r839 (  170 257 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.22 //y=1.22 //x2=55.18 //y2=1.375
r840 (  169 256 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.22 //y=0.91 //x2=55.18 //y2=0.755
r841 (  169 170 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=55.22 //y=0.91 //x2=55.22 //y2=1.22
r842 (  164 250 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.85 //y=1.375 //x2=54.735 //y2=1.375
r843 (  163 257 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.065 //y=1.375 //x2=55.18 //y2=1.375
r844 (  162 249 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.85 //y=0.755 //x2=54.735 //y2=0.755
r845 (  161 256 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.065 //y=0.755 //x2=55.18 //y2=0.755
r846 (  161 162 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=55.065 //y=0.755 //x2=54.85 //y2=0.755
r847 (  160 250 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.695 //y=1.22 //x2=54.735 //y2=1.375
r848 (  159 249 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.695 //y=0.91 //x2=54.735 //y2=0.755
r849 (  159 160 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=54.695 //y=0.91 //x2=54.695 //y2=1.22
r850 (  155 243 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=40.835 //y=4.79 //x2=40.7 //y2=4.79
r851 (  154 156 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=41.035 //y=4.79 //x2=41.11 //y2=4.865
r852 (  154 155 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=41.035 //y=4.79 //x2=40.835 //y2=4.79
r853 (  153 248 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=40.79 //y=1.915 //x2=40.715 //y2=2.08
r854 (  152 246 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=40.79 //y=1.45 //x2=40.75 //y2=1.375
r855 (  152 153 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=40.79 //y=1.45 //x2=40.79 //y2=1.915
r856 (  151 246 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.79 //y=1.22 //x2=40.75 //y2=1.375
r857 (  150 245 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.79 //y=0.91 //x2=40.75 //y2=0.755
r858 (  150 151 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=40.79 //y=0.91 //x2=40.79 //y2=1.22
r859 (  145 239 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.42 //y=1.375 //x2=40.305 //y2=1.375
r860 (  144 246 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.635 //y=1.375 //x2=40.75 //y2=1.375
r861 (  143 238 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.42 //y=0.755 //x2=40.305 //y2=0.755
r862 (  142 245 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.635 //y=0.755 //x2=40.75 //y2=0.755
r863 (  142 143 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=40.635 //y=0.755 //x2=40.42 //y2=0.755
r864 (  141 239 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.265 //y=1.22 //x2=40.305 //y2=1.375
r865 (  140 238 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.265 //y=0.91 //x2=40.305 //y2=0.755
r866 (  140 141 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=40.265 //y=0.91 //x2=40.265 //y2=1.22
r867 (  136 232 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=26.405 //y=4.79 //x2=26.27 //y2=4.79
r868 (  135 137 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=26.605 //y=4.79 //x2=26.68 //y2=4.865
r869 (  135 136 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=26.605 //y=4.79 //x2=26.405 //y2=4.79
r870 (  134 237 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.915 //x2=26.285 //y2=2.08
r871 (  133 235 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.45 //x2=26.32 //y2=1.375
r872 (  133 134 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.45 //x2=26.36 //y2=1.915
r873 (  132 235 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.22 //x2=26.32 //y2=1.375
r874 (  131 234 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.36 //y=0.91 //x2=26.32 //y2=0.755
r875 (  131 132 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=26.36 //y=0.91 //x2=26.36 //y2=1.22
r876 (  126 228 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.99 //y=1.375 //x2=25.875 //y2=1.375
r877 (  125 235 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.205 //y=1.375 //x2=26.32 //y2=1.375
r878 (  124 227 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.99 //y=0.755 //x2=25.875 //y2=0.755
r879 (  123 234 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.205 //y=0.755 //x2=26.32 //y2=0.755
r880 (  123 124 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=26.205 //y=0.755 //x2=25.99 //y2=0.755
r881 (  122 228 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.835 //y=1.22 //x2=25.875 //y2=1.375
r882 (  121 227 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.835 //y=0.91 //x2=25.875 //y2=0.755
r883 (  121 122 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=25.835 //y=0.91 //x2=25.835 //y2=1.22
r884 (  117 221 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=11.975 //y=4.79 //x2=11.84 //y2=4.79
r885 (  116 118 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=12.175 //y=4.79 //x2=12.25 //y2=4.865
r886 (  116 117 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=12.175 //y=4.79 //x2=11.975 //y2=4.79
r887 (  115 226 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.915 //x2=11.855 //y2=2.08
r888 (  114 224 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.45 //x2=11.89 //y2=1.375
r889 (  114 115 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.45 //x2=11.93 //y2=1.915
r890 (  113 224 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.22 //x2=11.89 //y2=1.375
r891 (  112 223 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.93 //y=0.91 //x2=11.89 //y2=0.755
r892 (  112 113 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=11.93 //y=0.91 //x2=11.93 //y2=1.22
r893 (  107 217 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.56 //y=1.375 //x2=11.445 //y2=1.375
r894 (  106 224 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.775 //y=1.375 //x2=11.89 //y2=1.375
r895 (  105 216 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.56 //y=0.755 //x2=11.445 //y2=0.755
r896 (  104 223 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.775 //y=0.755 //x2=11.89 //y2=0.755
r897 (  104 105 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=11.775 //y=0.755 //x2=11.56 //y2=0.755
r898 (  103 217 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.405 //y=1.22 //x2=11.445 //y2=1.375
r899 (  102 216 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.405 //y=0.91 //x2=11.445 //y2=0.755
r900 (  102 103 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=11.405 //y=0.91 //x2=11.405 //y2=1.22
r901 (  101 213 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=84.4 //y=6.02 //x2=84.4 //y2=4.865
r902 (  100 277 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=83.96 //y=6.02 //x2=83.96 //y2=4.865
r903 (  99 194 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.97 //y=6.02 //x2=69.97 //y2=4.865
r904 (  98 266 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.53 //y=6.02 //x2=69.53 //y2=4.865
r905 (  97 175 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.54 //y=6.02 //x2=55.54 //y2=4.865
r906 (  96 255 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.1 //y=6.02 //x2=55.1 //y2=4.865
r907 (  95 156 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.11 //y=6.02 //x2=41.11 //y2=4.865
r908 (  94 244 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=40.67 //y=6.02 //x2=40.67 //y2=4.865
r909 (  93 137 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.68 //y=6.02 //x2=26.68 //y2=4.865
r910 (  92 233 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.24 //y=6.02 //x2=26.24 //y2=4.865
r911 (  91 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.25 //y=6.02 //x2=12.25 //y2=4.865
r912 (  90 222 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.81 //y=6.02 //x2=11.81 //y2=4.865
r913 (  89 201 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=83.817 //y=1.375 //x2=83.925 //y2=1.375
r914 (  89 202 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=83.817 //y=1.375 //x2=83.71 //y2=1.375
r915 (  88 182 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=69.387 //y=1.375 //x2=69.495 //y2=1.375
r916 (  88 183 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=69.387 //y=1.375 //x2=69.28 //y2=1.375
r917 (  87 163 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=54.957 //y=1.375 //x2=55.065 //y2=1.375
r918 (  87 164 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=54.957 //y=1.375 //x2=54.85 //y2=1.375
r919 (  86 144 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=40.527 //y=1.375 //x2=40.635 //y2=1.375
r920 (  86 145 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=40.527 //y=1.375 //x2=40.42 //y2=1.375
r921 (  85 125 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=26.097 //y=1.375 //x2=26.205 //y2=1.375
r922 (  85 126 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=26.097 //y=1.375 //x2=25.99 //y2=1.375
r923 (  84 106 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=11.667 //y=1.375 //x2=11.775 //y2=1.375
r924 (  84 107 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=11.667 //y=1.375 //x2=11.56 //y2=1.375
r925 (  82 274 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=83.99 //y=4.7 //x2=83.99 //y2=4.7
r926 (  80 82 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=83.99 //y=2.96 //x2=83.99 //y2=4.7
r927 (  77 281 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=83.99 //y=2.08 //x2=83.99 //y2=2.08
r928 (  77 80 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=83.99 //y=2.08 //x2=83.99 //y2=2.96
r929 (  74 263 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=69.56 //y=4.7 //x2=69.56 //y2=4.7
r930 (  68 270 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=69.56 //y=2.08 //x2=69.56 //y2=2.08
r931 (  65 252 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.13 //y=4.7 //x2=55.13 //y2=4.7
r932 (  60 259 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.13 //y=2.08 //x2=55.13 //y2=2.08
r933 (  57 241 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=40.7 //y=4.7 //x2=40.7 //y2=4.7
r934 (  51 248 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=40.7 //y=2.08 //x2=40.7 //y2=2.08
r935 (  48 230 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=4.7 //x2=26.27 //y2=4.7
r936 (  42 237 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=2.08 //x2=26.27 //y2=2.08
r937 (  39 219 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=4.7 //x2=11.84 //y2=4.7
r938 (  33 226 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=2.08 //x2=11.84 //y2=2.08
r939 (  31 74 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=69.56 //y=2.96 //x2=69.56 //y2=4.7
r940 (  30 31 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=69.56 //y=2.59 //x2=69.56 //y2=2.96
r941 (  30 68 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=69.56 //y=2.59 //x2=69.56 //y2=2.08
r942 (  29 65 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=55.13 //y=2.96 //x2=55.13 //y2=4.7
r943 (  29 60 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=55.13 //y=2.96 //x2=55.13 //y2=2.08
r944 (  28 57 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=40.7 //y=2.96 //x2=40.7 //y2=4.7
r945 (  27 28 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=40.7 //y=2.59 //x2=40.7 //y2=2.96
r946 (  27 51 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=40.7 //y=2.59 //x2=40.7 //y2=2.08
r947 (  26 48 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.96 //x2=26.27 //y2=4.7
r948 (  25 26 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.59 //x2=26.27 //y2=2.96
r949 (  25 42 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.59 //x2=26.27 //y2=2.08
r950 (  24 39 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.96 //x2=11.84 //y2=4.7
r951 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.59 //x2=11.84 //y2=2.96
r952 (  23 33 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.59 //x2=11.84 //y2=2.08
r953 (  22 80 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=83.99 //y=2.96 //x2=83.99 //y2=2.96
r954 (  20 31 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=69.56 //y=2.96 //x2=69.56 //y2=2.96
r955 (  18 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=55.13 //y=2.96 //x2=55.13 //y2=2.96
r956 (  16 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=40.7 //y=2.96 //x2=40.7 //y2=2.96
r957 (  14 26 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=26.27 //y=2.96 //x2=26.27 //y2=2.96
r958 (  12 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.84 //y=2.96 //x2=11.84 //y2=2.96
r959 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.675 //y=2.96 //x2=69.56 //y2=2.96
r960 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=83.875 //y=2.96 //x2=83.99 //y2=2.96
r961 (  9 10 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=83.875 //y=2.96 //x2=69.675 //y2=2.96
r962 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.245 //y=2.96 //x2=55.13 //y2=2.96
r963 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.445 //y=2.96 //x2=69.56 //y2=2.96
r964 (  7 8 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=69.445 //y=2.96 //x2=55.245 //y2=2.96
r965 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=40.815 //y=2.96 //x2=40.7 //y2=2.96
r966 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.015 //y=2.96 //x2=55.13 //y2=2.96
r967 (  5 6 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=55.015 //y=2.96 //x2=40.815 //y2=2.96
r968 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=26.385 //y=2.96 //x2=26.27 //y2=2.96
r969 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=40.585 //y=2.96 //x2=40.7 //y2=2.96
r970 (  3 4 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=40.585 //y=2.96 //x2=26.385 //y2=2.96
r971 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.955 //y=2.96 //x2=11.84 //y2=2.96
r972 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=2.96 //x2=26.27 //y2=2.96
r973 (  1 2 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=2.96 //x2=11.955 //y2=2.96
ends PM_TMRDFFSNRNQNX1\%SN

subckt PM_TMRDFFSNRNQNX1\%noxref_21 ( 1 2 3 4 5 6 16 24 37 38 45 53 59 60 64 \
 66 73 74 75 76 77 78 79 80 81 82 83 87 88 89 94 96 99 100 104 105 106 111 113 \
 116 117 121 122 123 128 130 133 134 136 137 142 146 147 152 156 157 162 165 \
 167 168 169 )
c343 ( 169 0 ) capacitor c=0.023087f //x=75.295 //y=5.02
c344 ( 168 0 ) capacitor c=0.023519f //x=74.415 //y=5.02
c345 ( 167 0 ) capacitor c=0.0224735f //x=73.535 //y=5.02
c346 ( 165 0 ) capacitor c=0.00853354f //x=75.545 //y=0.915
c347 ( 162 0 ) capacitor c=0.0587755f //x=85.1 //y=4.7
c348 ( 157 0 ) capacitor c=0.0273931f //x=85.1 //y=1.915
c349 ( 156 0 ) capacitor c=0.0456313f //x=85.1 //y=2.08
c350 ( 152 0 ) capacitor c=0.0588394f //x=70.67 //y=4.7
c351 ( 147 0 ) capacitor c=0.0273931f //x=70.67 //y=1.915
c352 ( 146 0 ) capacitor c=0.0456313f //x=70.67 //y=2.08
c353 ( 142 0 ) capacitor c=0.0589949f //x=65.86 //y=4.7
c354 ( 137 0 ) capacitor c=0.0273931f //x=65.86 //y=1.915
c355 ( 136 0 ) capacitor c=0.0456313f //x=65.86 //y=2.08
c356 ( 134 0 ) capacitor c=0.0432517f //x=85.62 //y=1.26
c357 ( 133 0 ) capacitor c=0.0200379f //x=85.62 //y=0.915
c358 ( 130 0 ) capacitor c=0.0148873f //x=85.465 //y=1.415
c359 ( 128 0 ) capacitor c=0.0157803f //x=85.465 //y=0.76
c360 ( 123 0 ) capacitor c=0.0218028f //x=85.09 //y=1.57
c361 ( 122 0 ) capacitor c=0.0207459f //x=85.09 //y=1.26
c362 ( 121 0 ) capacitor c=0.0194308f //x=85.09 //y=0.915
c363 ( 117 0 ) capacitor c=0.0432517f //x=71.19 //y=1.26
c364 ( 116 0 ) capacitor c=0.0200379f //x=71.19 //y=0.915
c365 ( 113 0 ) capacitor c=0.0148873f //x=71.035 //y=1.415
c366 ( 111 0 ) capacitor c=0.0157803f //x=71.035 //y=0.76
c367 ( 106 0 ) capacitor c=0.0218028f //x=70.66 //y=1.57
c368 ( 105 0 ) capacitor c=0.0207459f //x=70.66 //y=1.26
c369 ( 104 0 ) capacitor c=0.0194308f //x=70.66 //y=0.915
c370 ( 100 0 ) capacitor c=0.0432517f //x=66.38 //y=1.26
c371 ( 99 0 ) capacitor c=0.0200379f //x=66.38 //y=0.915
c372 ( 96 0 ) capacitor c=0.0148873f //x=66.225 //y=1.415
c373 ( 94 0 ) capacitor c=0.0157803f //x=66.225 //y=0.76
c374 ( 89 0 ) capacitor c=0.0218028f //x=65.85 //y=1.57
c375 ( 88 0 ) capacitor c=0.0207459f //x=65.85 //y=1.26
c376 ( 87 0 ) capacitor c=0.0194308f //x=65.85 //y=0.915
c377 ( 83 0 ) capacitor c=0.158794f //x=85.28 //y=6.02
c378 ( 82 0 ) capacitor c=0.110114f //x=84.84 //y=6.02
c379 ( 81 0 ) capacitor c=0.158754f //x=70.85 //y=6.02
c380 ( 80 0 ) capacitor c=0.109949f //x=70.41 //y=6.02
c381 ( 79 0 ) capacitor c=0.158754f //x=66.04 //y=6.02
c382 ( 78 0 ) capacitor c=0.109949f //x=65.6 //y=6.02
c383 ( 74 0 ) capacitor c=0.00106608f //x=75.44 //y=5.155
c384 ( 73 0 ) capacitor c=0.00191414f //x=74.56 //y=5.155
c385 ( 66 0 ) capacitor c=0.0836242f //x=85.1 //y=2.08
c386 ( 64 0 ) capacitor c=0.10494f //x=76.22 //y=3.7
c387 ( 60 0 ) capacitor c=0.00398962f //x=75.82 //y=1.665
c388 ( 59 0 ) capacitor c=0.0137288f //x=76.135 //y=1.665
c389 ( 53 0 ) capacitor c=0.0283082f //x=76.135 //y=5.155
c390 ( 45 0 ) capacitor c=0.0170864f //x=75.355 //y=5.155
c391 ( 38 0 ) capacitor c=0.00316998f //x=73.765 //y=5.155
c392 ( 37 0 ) capacitor c=0.014258f //x=74.475 //y=5.155
c393 ( 24 0 ) capacitor c=0.0790362f //x=70.67 //y=2.08
c394 ( 16 0 ) capacitor c=0.076565f //x=65.86 //y=2.08
c395 ( 6 0 ) capacitor c=0.0055354f //x=76.335 //y=3.7
c396 ( 5 0 ) capacitor c=0.164574f //x=84.985 //y=3.7
c397 ( 4 0 ) capacitor c=0.00533183f //x=70.785 //y=3.7
c398 ( 3 0 ) capacitor c=0.0753575f //x=76.105 //y=3.7
c399 ( 2 0 ) capacitor c=0.00692093f //x=65.975 //y=3.7
c400 ( 1 0 ) capacitor c=0.0665749f //x=70.555 //y=3.7
r401 (  156 157 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=85.1 //y=2.08 //x2=85.1 //y2=1.915
r402 (  146 147 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=70.67 //y=2.08 //x2=70.67 //y2=1.915
r403 (  136 137 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=65.86 //y=2.08 //x2=65.86 //y2=1.915
r404 (  134 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.62 //y=1.26 //x2=85.58 //y2=1.415
r405 (  133 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.62 //y=0.915 //x2=85.58 //y2=0.76
r406 (  133 134 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=85.62 //y=0.915 //x2=85.62 //y2=1.26
r407 (  131 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.245 //y=1.415 //x2=85.13 //y2=1.415
r408 (  130 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.465 //y=1.415 //x2=85.58 //y2=1.415
r409 (  129 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.245 //y=0.76 //x2=85.13 //y2=0.76
r410 (  128 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.465 //y=0.76 //x2=85.58 //y2=0.76
r411 (  128 129 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=85.465 //y=0.76 //x2=85.245 //y2=0.76
r412 (  125 162 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=85.28 //y=4.865 //x2=85.1 //y2=4.7
r413 (  123 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.09 //y=1.57 //x2=85.13 //y2=1.415
r414 (  123 157 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=85.09 //y=1.57 //x2=85.09 //y2=1.915
r415 (  122 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.09 //y=1.26 //x2=85.13 //y2=1.415
r416 (  121 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.09 //y=0.915 //x2=85.13 //y2=0.76
r417 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=85.09 //y=0.915 //x2=85.09 //y2=1.26
r418 (  118 162 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=84.84 //y=4.865 //x2=85.1 //y2=4.7
r419 (  117 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.19 //y=1.26 //x2=71.15 //y2=1.415
r420 (  116 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.19 //y=0.915 //x2=71.15 //y2=0.76
r421 (  116 117 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=71.19 //y=0.915 //x2=71.19 //y2=1.26
r422 (  114 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.815 //y=1.415 //x2=70.7 //y2=1.415
r423 (  113 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.035 //y=1.415 //x2=71.15 //y2=1.415
r424 (  112 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.815 //y=0.76 //x2=70.7 //y2=0.76
r425 (  111 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.035 //y=0.76 //x2=71.15 //y2=0.76
r426 (  111 112 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=71.035 //y=0.76 //x2=70.815 //y2=0.76
r427 (  108 152 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=70.85 //y=4.865 //x2=70.67 //y2=4.7
r428 (  106 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.66 //y=1.57 //x2=70.7 //y2=1.415
r429 (  106 147 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=70.66 //y=1.57 //x2=70.66 //y2=1.915
r430 (  105 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.66 //y=1.26 //x2=70.7 //y2=1.415
r431 (  104 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.66 //y=0.915 //x2=70.7 //y2=0.76
r432 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=70.66 //y=0.915 //x2=70.66 //y2=1.26
r433 (  101 152 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=70.41 //y=4.865 //x2=70.67 //y2=4.7
r434 (  100 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.38 //y=1.26 //x2=66.34 //y2=1.415
r435 (  99 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.38 //y=0.915 //x2=66.34 //y2=0.76
r436 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=66.38 //y=0.915 //x2=66.38 //y2=1.26
r437 (  97 140 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.005 //y=1.415 //x2=65.89 //y2=1.415
r438 (  96 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.225 //y=1.415 //x2=66.34 //y2=1.415
r439 (  95 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.005 //y=0.76 //x2=65.89 //y2=0.76
r440 (  94 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.225 //y=0.76 //x2=66.34 //y2=0.76
r441 (  94 95 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=66.225 //y=0.76 //x2=66.005 //y2=0.76
r442 (  91 142 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=66.04 //y=4.865 //x2=65.86 //y2=4.7
r443 (  89 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.85 //y=1.57 //x2=65.89 //y2=1.415
r444 (  89 137 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=65.85 //y=1.57 //x2=65.85 //y2=1.915
r445 (  88 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.85 //y=1.26 //x2=65.89 //y2=1.415
r446 (  87 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.85 //y=0.915 //x2=65.89 //y2=0.76
r447 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=65.85 //y=0.915 //x2=65.85 //y2=1.26
r448 (  84 142 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=65.6 //y=4.865 //x2=65.86 //y2=4.7
r449 (  83 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=85.28 //y=6.02 //x2=85.28 //y2=4.865
r450 (  82 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=84.84 //y=6.02 //x2=84.84 //y2=4.865
r451 (  81 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.85 //y=6.02 //x2=70.85 //y2=4.865
r452 (  80 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.41 //y=6.02 //x2=70.41 //y2=4.865
r453 (  79 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.04 //y=6.02 //x2=66.04 //y2=4.865
r454 (  78 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=65.6 //y=6.02 //x2=65.6 //y2=4.865
r455 (  77 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=85.355 //y=1.415 //x2=85.465 //y2=1.415
r456 (  77 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=85.355 //y=1.415 //x2=85.245 //y2=1.415
r457 (  76 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=70.925 //y=1.415 //x2=71.035 //y2=1.415
r458 (  76 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=70.925 //y=1.415 //x2=70.815 //y2=1.415
r459 (  75 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.115 //y=1.415 //x2=66.225 //y2=1.415
r460 (  75 97 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.115 //y=1.415 //x2=66.005 //y2=1.415
r461 (  71 162 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=85.1 //y=4.7 //x2=85.1 //y2=4.7
r462 (  69 71 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=85.1 //y=3.7 //x2=85.1 //y2=4.7
r463 (  66 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=85.1 //y=2.08 //x2=85.1 //y2=2.08
r464 (  66 69 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=85.1 //y=2.08 //x2=85.1 //y2=3.7
r465 (  62 64 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=76.22 //y=5.07 //x2=76.22 //y2=3.7
r466 (  61 64 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=76.22 //y=1.75 //x2=76.22 //y2=3.7
r467 (  59 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=76.135 //y=1.665 //x2=76.22 //y2=1.75
r468 (  59 60 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=76.135 //y=1.665 //x2=75.82 //y2=1.665
r469 (  55 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=75.735 //y=1.58 //x2=75.82 //y2=1.665
r470 (  55 165 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=75.735 //y=1.58 //x2=75.735 //y2=1.01
r471 (  54 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.525 //y=5.155 //x2=75.44 //y2=5.155
r472 (  53 62 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=76.135 //y=5.155 //x2=76.22 //y2=5.07
r473 (  53 54 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=76.135 //y=5.155 //x2=75.525 //y2=5.155
r474 (  47 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.44 //y=5.24 //x2=75.44 //y2=5.155
r475 (  47 169 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=75.44 //y=5.24 //x2=75.44 //y2=5.725
r476 (  46 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.645 //y=5.155 //x2=74.56 //y2=5.155
r477 (  45 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.355 //y=5.155 //x2=75.44 //y2=5.155
r478 (  45 46 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=75.355 //y=5.155 //x2=74.645 //y2=5.155
r479 (  39 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.56 //y=5.24 //x2=74.56 //y2=5.155
r480 (  39 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=74.56 //y=5.24 //x2=74.56 //y2=5.725
r481 (  37 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.475 //y=5.155 //x2=74.56 //y2=5.155
r482 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=74.475 //y=5.155 //x2=73.765 //y2=5.155
r483 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=73.68 //y=5.24 //x2=73.765 //y2=5.155
r484 (  31 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=73.68 //y=5.24 //x2=73.68 //y2=5.725
r485 (  29 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=4.7 //x2=70.67 //y2=4.7
r486 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=70.67 //y=3.7 //x2=70.67 //y2=4.7
r487 (  24 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=2.08 //x2=70.67 //y2=2.08
r488 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=70.67 //y=2.08 //x2=70.67 //y2=3.7
r489 (  21 142 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=65.86 //y=4.7 //x2=65.86 //y2=4.7
r490 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=65.86 //y=3.7 //x2=65.86 //y2=4.7
r491 (  16 136 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=65.86 //y=2.08 //x2=65.86 //y2=2.08
r492 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=65.86 //y=2.08 //x2=65.86 //y2=3.7
r493 (  14 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=85.1 //y=3.7 //x2=85.1 //y2=3.7
r494 (  12 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=76.22 //y=3.7 //x2=76.22 //y2=3.7
r495 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=70.67 //y=3.7 //x2=70.67 //y2=3.7
r496 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=65.86 //y=3.7 //x2=65.86 //y2=3.7
r497 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=76.335 //y=3.7 //x2=76.22 //y2=3.7
r498 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=84.985 //y=3.7 //x2=85.1 //y2=3.7
r499 (  5 6 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=84.985 //y=3.7 //x2=76.335 //y2=3.7
r500 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=70.785 //y=3.7 //x2=70.67 //y2=3.7
r501 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=76.105 //y=3.7 //x2=76.22 //y2=3.7
r502 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=76.105 //y=3.7 //x2=70.785 //y2=3.7
r503 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=65.975 //y=3.7 //x2=65.86 //y2=3.7
r504 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=3.7 //x2=70.67 //y2=3.7
r505 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=3.7 //x2=65.975 //y2=3.7
ends PM_TMRDFFSNRNQNX1\%noxref_21

subckt PM_TMRDFFSNRNQNX1\%noxref_22 ( 1 2 8 21 22 29 37 43 44 48 49 50 51 52 \
 53 57 58 59 64 66 69 70 72 73 78 81 83 84 85 )
c171 ( 85 0 ) capacitor c=0.023087f //x=84.915 //y=5.02
c172 ( 84 0 ) capacitor c=0.023519f //x=84.035 //y=5.02
c173 ( 83 0 ) capacitor c=0.0224735f //x=83.155 //y=5.02
c174 ( 81 0 ) capacitor c=0.0087111f //x=85.165 //y=0.915
c175 ( 78 0 ) capacitor c=0.0587755f //x=80.29 //y=4.7
c176 ( 73 0 ) capacitor c=0.0273931f //x=80.29 //y=1.915
c177 ( 72 0 ) capacitor c=0.0457015f //x=80.29 //y=2.08
c178 ( 70 0 ) capacitor c=0.0432517f //x=80.81 //y=1.26
c179 ( 69 0 ) capacitor c=0.0200379f //x=80.81 //y=0.915
c180 ( 66 0 ) capacitor c=0.0158629f //x=80.655 //y=1.415
c181 ( 64 0 ) capacitor c=0.0157803f //x=80.655 //y=0.76
c182 ( 59 0 ) capacitor c=0.0218028f //x=80.28 //y=1.57
c183 ( 58 0 ) capacitor c=0.0207459f //x=80.28 //y=1.26
c184 ( 57 0 ) capacitor c=0.0194308f //x=80.28 //y=0.915
c185 ( 53 0 ) capacitor c=0.158794f //x=80.47 //y=6.02
c186 ( 52 0 ) capacitor c=0.110114f //x=80.03 //y=6.02
c187 ( 50 0 ) capacitor c=0.00106608f //x=85.06 //y=5.155
c188 ( 49 0 ) capacitor c=0.00207319f //x=84.18 //y=5.155
c189 ( 48 0 ) capacitor c=0.108549f //x=85.84 //y=2.59
c190 ( 44 0 ) capacitor c=0.00398962f //x=85.44 //y=1.665
c191 ( 43 0 ) capacitor c=0.0137288f //x=85.755 //y=1.665
c192 ( 37 0 ) capacitor c=0.0281866f //x=85.755 //y=5.155
c193 ( 29 0 ) capacitor c=0.0176454f //x=84.975 //y=5.155
c194 ( 22 0 ) capacitor c=0.00332903f //x=83.385 //y=5.155
c195 ( 21 0 ) capacitor c=0.0148427f //x=84.095 //y=5.155
c196 ( 8 0 ) capacitor c=0.0838166f //x=80.29 //y=2.08
c197 ( 2 0 ) capacitor c=0.0158526f //x=80.405 //y=2.59
c198 ( 1 0 ) capacitor c=0.0993317f //x=85.725 //y=2.59
r199 (  72 73 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=80.29 //y=2.08 //x2=80.29 //y2=1.915
r200 (  70 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.81 //y=1.26 //x2=80.77 //y2=1.415
r201 (  69 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.81 //y=0.915 //x2=80.77 //y2=0.76
r202 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=80.81 //y=0.915 //x2=80.81 //y2=1.26
r203 (  67 76 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.435 //y=1.415 //x2=80.32 //y2=1.415
r204 (  66 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.655 //y=1.415 //x2=80.77 //y2=1.415
r205 (  65 75 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.435 //y=0.76 //x2=80.32 //y2=0.76
r206 (  64 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.655 //y=0.76 //x2=80.77 //y2=0.76
r207 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=80.655 //y=0.76 //x2=80.435 //y2=0.76
r208 (  61 78 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=80.47 //y=4.865 //x2=80.29 //y2=4.7
r209 (  59 76 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.28 //y=1.57 //x2=80.32 //y2=1.415
r210 (  59 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=80.28 //y=1.57 //x2=80.28 //y2=1.915
r211 (  58 76 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.28 //y=1.26 //x2=80.32 //y2=1.415
r212 (  57 75 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.28 //y=0.915 //x2=80.32 //y2=0.76
r213 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=80.28 //y=0.915 //x2=80.28 //y2=1.26
r214 (  54 78 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=80.03 //y=4.865 //x2=80.29 //y2=4.7
r215 (  53 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=80.47 //y=6.02 //x2=80.47 //y2=4.865
r216 (  52 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=80.03 //y=6.02 //x2=80.03 //y2=4.865
r217 (  51 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=80.545 //y=1.415 //x2=80.655 //y2=1.415
r218 (  51 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=80.545 //y=1.415 //x2=80.435 //y2=1.415
r219 (  46 48 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=85.84 //y=5.07 //x2=85.84 //y2=2.59
r220 (  45 48 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=85.84 //y=1.75 //x2=85.84 //y2=2.59
r221 (  43 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=85.755 //y=1.665 //x2=85.84 //y2=1.75
r222 (  43 44 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=85.755 //y=1.665 //x2=85.44 //y2=1.665
r223 (  39 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=85.355 //y=1.58 //x2=85.44 //y2=1.665
r224 (  39 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=85.355 //y=1.58 //x2=85.355 //y2=1.01
r225 (  38 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.145 //y=5.155 //x2=85.06 //y2=5.155
r226 (  37 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=85.755 //y=5.155 //x2=85.84 //y2=5.07
r227 (  37 38 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=85.755 //y=5.155 //x2=85.145 //y2=5.155
r228 (  31 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.06 //y=5.24 //x2=85.06 //y2=5.155
r229 (  31 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=85.06 //y=5.24 //x2=85.06 //y2=5.725
r230 (  30 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.265 //y=5.155 //x2=84.18 //y2=5.155
r231 (  29 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.975 //y=5.155 //x2=85.06 //y2=5.155
r232 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=84.975 //y=5.155 //x2=84.265 //y2=5.155
r233 (  23 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.18 //y=5.24 //x2=84.18 //y2=5.155
r234 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=84.18 //y=5.24 //x2=84.18 //y2=5.725
r235 (  21 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.095 //y=5.155 //x2=84.18 //y2=5.155
r236 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=84.095 //y=5.155 //x2=83.385 //y2=5.155
r237 (  15 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=83.3 //y=5.24 //x2=83.385 //y2=5.155
r238 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=83.3 //y=5.24 //x2=83.3 //y2=5.725
r239 (  13 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=80.29 //y=4.7 //x2=80.29 //y2=4.7
r240 (  11 13 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=80.29 //y=2.59 //x2=80.29 //y2=4.7
r241 (  8 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=80.29 //y=2.08 //x2=80.29 //y2=2.08
r242 (  8 11 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=80.29 //y=2.08 //x2=80.29 //y2=2.59
r243 (  6 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=85.84 //y=2.59 //x2=85.84 //y2=2.59
r244 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=80.29 //y=2.59 //x2=80.29 //y2=2.59
r245 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=80.405 //y=2.59 //x2=80.29 //y2=2.59
r246 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=85.725 //y=2.59 //x2=85.84 //y2=2.59
r247 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=85.725 //y=2.59 //x2=80.405 //y2=2.59
ends PM_TMRDFFSNRNQNX1\%noxref_22

subckt PM_TMRDFFSNRNQNX1\%noxref_23 ( 1 2 13 14 15 23 29 30 37 50 51 52 53 54 )
c91 ( 54 0 ) capacitor c=0.034295f //x=92.305 //y=5.025
c92 ( 53 0 ) capacitor c=0.0174957f //x=91.425 //y=5.025
c93 ( 51 0 ) capacitor c=0.0214849f //x=88.545 //y=5.025
c94 ( 50 0 ) capacitor c=0.0217161f //x=87.665 //y=5.025
c95 ( 49 0 ) capacitor c=0.00115294f //x=91.57 //y=6.91
c96 ( 37 0 ) capacitor c=0.0131238f //x=92.365 //y=6.91
c97 ( 30 0 ) capacitor c=0.00386507f //x=90.775 //y=6.91
c98 ( 29 0 ) capacitor c=0.00951687f //x=91.485 //y=6.91
c99 ( 23 0 ) capacitor c=0.0455351f //x=90.69 //y=5.21
c100 ( 15 0 ) capacitor c=0.00871244f //x=88.69 //y=5.295
c101 ( 14 0 ) capacitor c=0.00290434f //x=87.895 //y=5.21
c102 ( 13 0 ) capacitor c=0.0139202f //x=88.605 //y=5.21
c103 ( 2 0 ) capacitor c=0.0091252f //x=88.805 //y=5.21
c104 ( 1 0 ) capacitor c=0.0484159f //x=90.575 //y=5.21
r105 (  39 54 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=92.45 //y=6.825 //x2=92.45 //y2=6.74
r106 (  38 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.655 //y=6.91 //x2=91.57 //y2=6.91
r107 (  37 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=92.365 //y=6.91 //x2=92.45 //y2=6.825
r108 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=92.365 //y=6.91 //x2=91.655 //y2=6.91
r109 (  31 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.57 //y=6.825 //x2=91.57 //y2=6.91
r110 (  31 53 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.57 //y=6.825 //x2=91.57 //y2=6.74
r111 (  29 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.485 //y=6.91 //x2=91.57 //y2=6.91
r112 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=91.485 //y=6.91 //x2=90.775 //y2=6.91
r113 (  23 52 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=90.69 //y=5.21 //x2=90.69 //y2=6.06
r114 (  21 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=90.69 //y=6.825 //x2=90.775 //y2=6.91
r115 (  21 52 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=90.69 //y=6.825 //x2=90.69 //y2=6.74
r116 (  15 48 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=88.69 //y=5.295 //x2=88.69 //y2=5.17
r117 (  15 51 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=88.69 //y=5.295 //x2=88.69 //y2=6.06
r118 (  13 48 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=88.605 //y=5.21 //x2=88.69 //y2=5.17
r119 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=88.605 //y=5.21 //x2=87.895 //y2=5.21
r120 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=87.81 //y=5.295 //x2=87.895 //y2=5.21
r121 (  7 50 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=87.81 //y=5.295 //x2=87.81 //y2=5.72
r122 (  6 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=90.69 //y=5.21 //x2=90.69 //y2=5.21
r123 (  4 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=88.69 //y=5.21 //x2=88.69 //y2=5.21
r124 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=88.805 //y=5.21 //x2=88.69 //y2=5.21
r125 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=90.575 //y=5.21 //x2=90.69 //y2=5.21
r126 (  1 2 ) resistor r=1.68893 //w=0.131 //l=1.77 //layer=m1 \
 //thickness=0.36 //x=90.575 //y=5.21 //x2=88.805 //y2=5.21
ends PM_TMRDFFSNRNQNX1\%noxref_23

subckt PM_TMRDFFSNRNQNX1\%noxref_24 ( 1 2 3 4 5 12 22 23 30 38 44 45 49 51 59 \
 66 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 89 95 96 97 98 105 106 107 \
 108 109 111 114 117 118 119 120 121 122 123 124 128 130 133 134 135 136 157 \
 164 166 167 168 )
c390 ( 168 0 ) capacitor c=0.023087f //x=80.105 //y=5.02
c391 ( 167 0 ) capacitor c=0.023519f //x=79.225 //y=5.02
c392 ( 166 0 ) capacitor c=0.0224735f //x=78.345 //y=5.02
c393 ( 164 0 ) capacitor c=0.00853354f //x=80.355 //y=0.915
c394 ( 157 0 ) capacitor c=0.0583848f //x=93.98 //y=2.08
c395 ( 136 0 ) capacitor c=0.0316774f //x=94.685 //y=1.21
c396 ( 135 0 ) capacitor c=0.0187384f //x=94.685 //y=0.865
c397 ( 134 0 ) capacitor c=0.0590362f //x=94.325 //y=4.795
c398 ( 133 0 ) capacitor c=0.0296075f //x=94.615 //y=4.795
c399 ( 130 0 ) capacitor c=0.0157912f //x=94.53 //y=1.365
c400 ( 128 0 ) capacitor c=0.0149844f //x=94.53 //y=0.71
c401 ( 124 0 ) capacitor c=0.0302441f //x=94.155 //y=1.915
c402 ( 123 0 ) capacitor c=0.0234157f //x=94.155 //y=1.52
c403 ( 122 0 ) capacitor c=0.0234376f //x=94.155 //y=1.21
c404 ( 121 0 ) capacitor c=0.0199931f //x=94.155 //y=0.865
c405 ( 120 0 ) capacitor c=0.092271f //x=92.325 //y=1.915
c406 ( 119 0 ) capacitor c=0.0249466f //x=92.325 //y=1.56
c407 ( 118 0 ) capacitor c=0.0234397f //x=92.325 //y=1.25
c408 ( 117 0 ) capacitor c=0.0193195f //x=92.325 //y=0.905
c409 ( 114 0 ) capacitor c=0.0631944f //x=92.23 //y=4.87
c410 ( 111 0 ) capacitor c=0.0164325f //x=92.17 //y=1.405
c411 ( 109 0 ) capacitor c=0.0157803f //x=92.17 //y=0.75
c412 ( 108 0 ) capacitor c=0.010629f //x=91.865 //y=4.795
c413 ( 107 0 ) capacitor c=0.0194269f //x=92.155 //y=4.795
c414 ( 106 0 ) capacitor c=0.0353695f //x=91.795 //y=1.25
c415 ( 105 0 ) capacitor c=0.0175988f //x=91.795 //y=0.905
c416 ( 98 0 ) capacitor c=0.0556143f //x=83.155 //y=4.79
c417 ( 97 0 ) capacitor c=0.0293157f //x=83.445 //y=4.79
c418 ( 96 0 ) capacitor c=0.0347816f //x=83.11 //y=1.22
c419 ( 95 0 ) capacitor c=0.0187487f //x=83.11 //y=0.875
c420 ( 89 0 ) capacitor c=0.0137055f //x=82.955 //y=1.375
c421 ( 87 0 ) capacitor c=0.0149861f //x=82.955 //y=0.72
c422 ( 86 0 ) capacitor c=0.095966f //x=82.58 //y=1.915
c423 ( 85 0 ) capacitor c=0.0228993f //x=82.58 //y=1.53
c424 ( 84 0 ) capacitor c=0.0234352f //x=82.58 //y=1.22
c425 ( 83 0 ) capacitor c=0.0198724f //x=82.58 //y=0.875
c426 ( 82 0 ) capacitor c=0.110622f //x=94.69 //y=6.025
c427 ( 81 0 ) capacitor c=0.154068f //x=94.25 //y=6.025
c428 ( 80 0 ) capacitor c=0.154291f //x=92.23 //y=6.025
c429 ( 79 0 ) capacitor c=0.110404f //x=91.79 //y=6.025
c430 ( 78 0 ) capacitor c=0.110114f //x=83.52 //y=6.02
c431 ( 77 0 ) capacitor c=0.158956f //x=83.08 //y=6.02
c432 ( 73 0 ) capacitor c=0.00106608f //x=80.25 //y=5.155
c433 ( 72 0 ) capacitor c=0.00207319f //x=79.37 //y=5.155
c434 ( 66 0 ) capacitor c=0.100793f //x=93.98 //y=2.08
c435 ( 59 0 ) capacitor c=0.107544f //x=92.5 //y=2.08
c436 ( 51 0 ) capacitor c=0.0970431f //x=82.88 //y=2.08
c437 ( 49 0 ) capacitor c=0.107181f //x=81.03 //y=2.22
c438 ( 45 0 ) capacitor c=0.00431225f //x=80.63 //y=1.665
c439 ( 44 0 ) capacitor c=0.0141892f //x=80.945 //y=1.665
c440 ( 38 0 ) capacitor c=0.0283082f //x=80.945 //y=5.155
c441 ( 30 0 ) capacitor c=0.0176454f //x=80.165 //y=5.155
c442 ( 23 0 ) capacitor c=0.00332903f //x=78.575 //y=5.155
c443 ( 22 0 ) capacitor c=0.0148427f //x=79.285 //y=5.155
c444 ( 12 0 ) capacitor c=0.0148272f //x=92.5 //y=2.08
c445 ( 5 0 ) capacitor c=0.0465668f //x=93.865 //y=2.08
c446 ( 4 0 ) capacitor c=0.00560639f //x=82.995 //y=2.22
c447 ( 3 0 ) capacitor c=0.244868f //x=92.355 //y=2.22
c448 ( 2 0 ) capacitor c=0.00833032f //x=81.145 //y=2.22
c449 ( 1 0 ) capacitor c=0.0348685f //x=82.765 //y=2.22
r450 (  136 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.685 //y=1.21 //x2=94.645 //y2=1.365
r451 (  135 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.685 //y=0.865 //x2=94.645 //y2=0.71
r452 (  135 136 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=94.685 //y=0.865 //x2=94.685 //y2=1.21
r453 (  133 137 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=94.615 //y=4.795 //x2=94.69 //y2=4.87
r454 (  133 134 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=94.615 //y=4.795 //x2=94.325 //y2=4.795
r455 (  131 161 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=94.31 //y=1.365 //x2=94.195 //y2=1.365
r456 (  130 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=94.53 //y=1.365 //x2=94.645 //y2=1.365
r457 (  129 160 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=94.31 //y=0.71 //x2=94.195 //y2=0.71
r458 (  128 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=94.53 //y=0.71 //x2=94.645 //y2=0.71
r459 (  128 129 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=94.53 //y=0.71 //x2=94.31 //y2=0.71
r460 (  125 134 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=94.25 //y=4.87 //x2=94.325 //y2=4.795
r461 (  125 159 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=94.25 //y=4.87 //x2=93.98 //y2=4.705
r462 (  124 157 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=94.155 //y=1.915 //x2=93.98 //y2=2.08
r463 (  123 161 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.155 //y=1.52 //x2=94.195 //y2=1.365
r464 (  123 124 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=94.155 //y=1.52 //x2=94.155 //y2=1.915
r465 (  122 161 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.155 //y=1.21 //x2=94.195 //y2=1.365
r466 (  121 160 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.155 //y=0.865 //x2=94.195 //y2=0.71
r467 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=94.155 //y=0.865 //x2=94.155 //y2=1.21
r468 (  120 153 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=92.325 //y=1.915 //x2=92.5 //y2=2.08
r469 (  119 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=92.325 //y=1.56 //x2=92.285 //y2=1.405
r470 (  119 120 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=92.325 //y=1.56 //x2=92.325 //y2=1.915
r471 (  118 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=92.325 //y=1.25 //x2=92.285 //y2=1.405
r472 (  117 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=92.325 //y=0.905 //x2=92.285 //y2=0.75
r473 (  117 118 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=92.325 //y=0.905 //x2=92.325 //y2=1.25
r474 (  114 155 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=92.23 //y=4.87 //x2=92.5 //y2=4.705
r475 (  112 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=91.95 //y=1.405 //x2=91.835 //y2=1.405
r476 (  111 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=92.17 //y=1.405 //x2=92.285 //y2=1.405
r477 (  110 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=91.95 //y=0.75 //x2=91.835 //y2=0.75
r478 (  109 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=92.17 //y=0.75 //x2=92.285 //y2=0.75
r479 (  109 110 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=92.17 //y=0.75 //x2=91.95 //y2=0.75
r480 (  107 114 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=92.155 //y=4.795 //x2=92.23 //y2=4.87
r481 (  107 108 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=92.155 //y=4.795 //x2=91.865 //y2=4.795
r482 (  106 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=91.795 //y=1.25 //x2=91.835 //y2=1.405
r483 (  105 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=91.795 //y=0.905 //x2=91.835 //y2=0.75
r484 (  105 106 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=91.795 //y=0.905 //x2=91.795 //y2=1.25
r485 (  102 108 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=91.79 //y=4.87 //x2=91.865 //y2=4.795
r486 (  97 99 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=83.445 //y=4.79 //x2=83.52 //y2=4.865
r487 (  97 98 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=83.445 //y=4.79 //x2=83.155 //y2=4.79
r488 (  96 147 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.11 //y=1.22 //x2=83.07 //y2=1.375
r489 (  95 146 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.11 //y=0.875 //x2=83.07 //y2=0.72
r490 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=83.11 //y=0.875 //x2=83.11 //y2=1.22
r491 (  92 98 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=83.08 //y=4.865 //x2=83.155 //y2=4.79
r492 (  92 145 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=83.08 //y=4.865 //x2=82.88 //y2=4.7
r493 (  90 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.735 //y=1.375 //x2=82.62 //y2=1.375
r494 (  89 147 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.955 //y=1.375 //x2=83.07 //y2=1.375
r495 (  88 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.735 //y=0.72 //x2=82.62 //y2=0.72
r496 (  87 146 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.955 //y=0.72 //x2=83.07 //y2=0.72
r497 (  87 88 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=82.955 //y=0.72 //x2=82.735 //y2=0.72
r498 (  86 143 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=82.58 //y=1.915 //x2=82.88 //y2=2.08
r499 (  85 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.58 //y=1.53 //x2=82.62 //y2=1.375
r500 (  85 86 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=82.58 //y=1.53 //x2=82.58 //y2=1.915
r501 (  84 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.58 //y=1.22 //x2=82.62 //y2=1.375
r502 (  83 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.58 //y=0.875 //x2=82.62 //y2=0.72
r503 (  83 84 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=82.58 //y=0.875 //x2=82.58 //y2=1.22
r504 (  82 137 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=94.69 //y=6.025 //x2=94.69 //y2=4.87
r505 (  81 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=94.25 //y=6.025 //x2=94.25 //y2=4.87
r506 (  80 114 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=92.23 //y=6.025 //x2=92.23 //y2=4.87
r507 (  79 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=91.79 //y=6.025 //x2=91.79 //y2=4.87
r508 (  78 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=83.52 //y=6.02 //x2=83.52 //y2=4.865
r509 (  77 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=83.08 //y=6.02 //x2=83.08 //y2=4.865
r510 (  76 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=94.42 //y=1.365 //x2=94.53 //y2=1.365
r511 (  76 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=94.42 //y=1.365 //x2=94.31 //y2=1.365
r512 (  75 111 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=92.06 //y=1.405 //x2=92.17 //y2=1.405
r513 (  75 112 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=92.06 //y=1.405 //x2=91.95 //y2=1.405
r514 (  74 89 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.845 //y=1.375 //x2=82.955 //y2=1.375
r515 (  74 90 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.845 //y=1.375 //x2=82.735 //y2=1.375
r516 (  70 159 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=93.98 //y=4.705 //x2=93.98 //y2=4.705
r517 (  66 157 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=93.98 //y=2.08 //x2=93.98 //y2=2.08
r518 (  66 70 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=93.98 //y=2.08 //x2=93.98 //y2=4.705
r519 (  63 155 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=92.5 //y=4.705 //x2=92.5 //y2=4.705
r520 (  59 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=92.5 //y=2.08 //x2=92.5 //y2=2.08
r521 (  59 63 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=92.5 //y=2.08 //x2=92.5 //y2=4.705
r522 (  56 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=82.88 //y=4.7 //x2=82.88 //y2=4.7
r523 (  54 56 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=82.88 //y=2.22 //x2=82.88 //y2=4.7
r524 (  51 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=82.88 //y=2.08 //x2=82.88 //y2=2.08
r525 (  51 54 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=82.88 //y=2.08 //x2=82.88 //y2=2.22
r526 (  47 49 ) resistor r=195.08 //w=0.187 //l=2.85 //layer=li \
 //thickness=0.1 //x=81.03 //y=5.07 //x2=81.03 //y2=2.22
r527 (  46 49 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=81.03 //y=1.75 //x2=81.03 //y2=2.22
r528 (  44 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=80.945 //y=1.665 //x2=81.03 //y2=1.75
r529 (  44 45 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=80.945 //y=1.665 //x2=80.63 //y2=1.665
r530 (  40 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=80.545 //y=1.58 //x2=80.63 //y2=1.665
r531 (  40 164 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=80.545 //y=1.58 //x2=80.545 //y2=1.01
r532 (  39 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.335 //y=5.155 //x2=80.25 //y2=5.155
r533 (  38 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=80.945 //y=5.155 //x2=81.03 //y2=5.07
r534 (  38 39 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=80.945 //y=5.155 //x2=80.335 //y2=5.155
r535 (  32 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.25 //y=5.24 //x2=80.25 //y2=5.155
r536 (  32 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=80.25 //y=5.24 //x2=80.25 //y2=5.725
r537 (  31 72 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.455 //y=5.155 //x2=79.37 //y2=5.155
r538 (  30 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.165 //y=5.155 //x2=80.25 //y2=5.155
r539 (  30 31 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=80.165 //y=5.155 //x2=79.455 //y2=5.155
r540 (  24 72 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.37 //y=5.24 //x2=79.37 //y2=5.155
r541 (  24 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=79.37 //y=5.24 //x2=79.37 //y2=5.725
r542 (  22 72 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.285 //y=5.155 //x2=79.37 //y2=5.155
r543 (  22 23 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=79.285 //y=5.155 //x2=78.575 //y2=5.155
r544 (  16 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=78.49 //y=5.24 //x2=78.575 //y2=5.155
r545 (  16 166 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=78.49 //y=5.24 //x2=78.49 //y2=5.725
r546 (  15 66 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=93.98 //y=2.08 //x2=93.98 //y2=2.08
r547 (  12 59 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=92.5 //y=2.08 //x2=92.5 //y2=2.08
r548 (  12 13 ) resistor r=0.0678295 //w=0.258 //l=0.14 //layer=m1 \
 //thickness=0.36 //x=92.485 //y=2.08 //x2=92.485 //y2=2.22
r549 (  10 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=82.88 //y=2.22 //x2=82.88 //y2=2.22
r550 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=81.03 //y=2.22 //x2=81.03 //y2=2.22
r551 (  6 12 ) resistor r=0.032569 //w=0.258 //l=0.13 //layer=m1 \
 //thickness=0.36 //x=92.615 //y=2.08 //x2=92.485 //y2=2.08
r552 (  5 15 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=93.865 //y=2.08 //x2=93.98 //y2=2.08
r553 (  5 6 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=93.865 //y=2.08 //x2=92.615 //y2=2.08
r554 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=82.995 //y=2.22 //x2=82.88 //y2=2.22
r555 (  3 13 ) resistor r=0.032569 //w=0.258 //l=0.13 //layer=m1 \
 //thickness=0.36 //x=92.355 //y=2.22 //x2=92.485 //y2=2.22
r556 (  3 4 ) resistor r=8.9313 //w=0.131 //l=9.36 //layer=m1 //thickness=0.36 \
 //x=92.355 //y=2.22 //x2=82.995 //y2=2.22
r557 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=81.145 //y=2.22 //x2=81.03 //y2=2.22
r558 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=82.765 //y=2.22 //x2=82.88 //y2=2.22
r559 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=82.765 //y=2.22 //x2=81.145 //y2=2.22
ends PM_TMRDFFSNRNQNX1\%noxref_24

subckt PM_TMRDFFSNRNQNX1\%noxref_25 ( 1 2 13 14 15 21 27 28 35 46 47 48 49 50 )
c89 ( 50 0 ) capacitor c=0.0306574f //x=95.645 //y=5.025
c90 ( 49 0 ) capacitor c=0.0173945f //x=94.765 //y=5.025
c91 ( 47 0 ) capacitor c=0.0169278f //x=91.865 //y=5.025
c92 ( 46 0 ) capacitor c=0.0166762f //x=90.985 //y=5.025
c93 ( 45 0 ) capacitor c=0.00115294f //x=94.91 //y=6.91
c94 ( 35 0 ) capacitor c=0.0132983f //x=95.705 //y=6.91
c95 ( 28 0 ) capacitor c=0.00388794f //x=94.115 //y=6.91
c96 ( 27 0 ) capacitor c=0.00985708f //x=94.825 //y=6.91
c97 ( 21 0 ) capacitor c=0.0442221f //x=94.03 //y=5.21
c98 ( 15 0 ) capacitor c=0.0105083f //x=92.01 //y=5.295
c99 ( 14 0 ) capacitor c=0.00227812f //x=91.215 //y=5.21
c100 ( 13 0 ) capacitor c=0.0174384f //x=91.925 //y=5.21
c101 ( 2 0 ) capacitor c=0.00682032f //x=92.125 //y=5.21
c102 ( 1 0 ) capacitor c=0.0574911f //x=93.915 //y=5.21
r103 (  37 50 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=95.79 //y=6.825 //x2=95.79 //y2=6.74
r104 (  36 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.995 //y=6.91 //x2=94.91 //y2=6.91
r105 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=95.705 //y=6.91 //x2=95.79 //y2=6.825
r106 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=95.705 //y=6.91 //x2=94.995 //y2=6.91
r107 (  29 45 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.91 //y=6.825 //x2=94.91 //y2=6.91
r108 (  29 49 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.91 //y=6.825 //x2=94.91 //y2=6.74
r109 (  27 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.825 //y=6.91 //x2=94.91 //y2=6.91
r110 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=94.825 //y=6.91 //x2=94.115 //y2=6.91
r111 (  21 48 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=94.03 //y=5.21 //x2=94.03 //y2=6.06
r112 (  19 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=94.03 //y=6.825 //x2=94.115 //y2=6.91
r113 (  19 48 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.03 //y=6.825 //x2=94.03 //y2=6.74
r114 (  15 44 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=92.01 //y=5.295 //x2=92.01 //y2=5.17
r115 (  15 47 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=92.01 //y=5.295 //x2=92.01 //y2=6.06
r116 (  13 44 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=91.925 //y=5.21 //x2=92.01 //y2=5.17
r117 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=91.925 //y=5.21 //x2=91.215 //y2=5.21
r118 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=91.13 //y=5.295 //x2=91.215 //y2=5.21
r119 (  7 46 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=91.13 //y=5.295 //x2=91.13 //y2=5.72
r120 (  6 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=94.03 //y=5.21 //x2=94.03 //y2=5.21
r121 (  4 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=92.01 //y=5.21 //x2=92.01 //y2=5.21
r122 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=92.125 //y=5.21 //x2=92.01 //y2=5.21
r123 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=93.915 //y=5.21 //x2=94.03 //y2=5.21
r124 (  1 2 ) resistor r=1.70802 //w=0.131 //l=1.79 //layer=m1 \
 //thickness=0.36 //x=93.915 //y=5.21 //x2=92.125 //y2=5.21
ends PM_TMRDFFSNRNQNX1\%noxref_25

subckt PM_TMRDFFSNRNQNX1\%noxref_26 ( 1 2 3 4 6 7 8 10 11 12 13 14 29 30 37 45 \
 51 52 56 58 65 67 73 77 78 82 85 86 87 88 89 90 91 92 93 94 95 96 97 98 100 \
 106 107 108 109 113 114 115 120 122 124 130 131 132 133 134 139 141 143 149 \
 150 160 161 164 172 173 176 184 186 187 188 )
c455 ( 188 0 ) capacitor c=0.023087f //x=51.245 //y=5.02
c456 ( 187 0 ) capacitor c=0.023519f //x=50.365 //y=5.02
c457 ( 186 0 ) capacitor c=0.0224735f //x=49.485 //y=5.02
c458 ( 184 0 ) capacitor c=0.00853354f //x=51.495 //y=0.915
c459 ( 176 0 ) capacitor c=0.0352016f //x=95.11 //y=4.705
c460 ( 173 0 ) capacitor c=0.0279733f //x=95.09 //y=1.915
c461 ( 172 0 ) capacitor c=0.0467621f //x=95.09 //y=2.08
c462 ( 164 0 ) capacitor c=0.03845f //x=88.47 //y=4.705
c463 ( 161 0 ) capacitor c=0.0300885f //x=88.43 //y=1.915
c464 ( 160 0 ) capacitor c=0.0504818f //x=88.43 //y=2.08
c465 ( 150 0 ) capacitor c=0.0237734f //x=95.655 //y=1.255
c466 ( 149 0 ) capacitor c=0.0191782f //x=95.655 //y=0.905
c467 ( 143 0 ) capacitor c=0.0351663f //x=95.5 //y=1.405
c468 ( 141 0 ) capacitor c=0.0157803f //x=95.5 //y=0.75
c469 ( 139 0 ) capacitor c=0.0373879f //x=95.495 //y=4.795
c470 ( 134 0 ) capacitor c=0.0200628f //x=95.125 //y=1.56
c471 ( 133 0 ) capacitor c=0.0168575f //x=95.125 //y=1.255
c472 ( 132 0 ) capacitor c=0.0174993f //x=95.125 //y=0.905
c473 ( 131 0 ) capacitor c=0.0435065f //x=88.995 //y=1.25
c474 ( 130 0 ) capacitor c=0.019286f //x=88.995 //y=0.905
c475 ( 124 0 ) capacitor c=0.0164316f //x=88.84 //y=1.405
c476 ( 122 0 ) capacitor c=0.0157795f //x=88.84 //y=0.75
c477 ( 120 0 ) capacitor c=0.029531f //x=88.835 //y=4.795
c478 ( 115 0 ) capacitor c=0.0206178f //x=88.465 //y=1.56
c479 ( 114 0 ) capacitor c=0.016848f //x=88.465 //y=1.25
c480 ( 113 0 ) capacitor c=0.0174777f //x=88.465 //y=0.905
c481 ( 109 0 ) capacitor c=0.0547611f //x=54.295 //y=4.79
c482 ( 108 0 ) capacitor c=0.0294456f //x=54.585 //y=4.79
c483 ( 107 0 ) capacitor c=0.0347816f //x=54.25 //y=1.22
c484 ( 106 0 ) capacitor c=0.0187487f //x=54.25 //y=0.875
c485 ( 100 0 ) capacitor c=0.0137055f //x=54.095 //y=1.375
c486 ( 98 0 ) capacitor c=0.0149861f //x=54.095 //y=0.72
c487 ( 97 0 ) capacitor c=0.096037f //x=53.72 //y=1.915
c488 ( 96 0 ) capacitor c=0.0228993f //x=53.72 //y=1.53
c489 ( 95 0 ) capacitor c=0.0234352f //x=53.72 //y=1.22
c490 ( 94 0 ) capacitor c=0.0198724f //x=53.72 //y=0.875
c491 ( 93 0 ) capacitor c=0.15325f //x=95.57 //y=6.025
c492 ( 92 0 ) capacitor c=0.110411f //x=95.13 //y=6.025
c493 ( 91 0 ) capacitor c=0.154236f //x=88.91 //y=6.025
c494 ( 90 0 ) capacitor c=0.110294f //x=88.47 //y=6.025
c495 ( 89 0 ) capacitor c=0.109949f //x=54.66 //y=6.02
c496 ( 88 0 ) capacitor c=0.158483f //x=54.22 //y=6.02
c497 ( 82 0 ) capacitor c=0.00501304f //x=95.11 //y=4.705
c498 ( 78 0 ) capacitor c=9.74268e-19 //x=51.39 //y=5.155
c499 ( 77 0 ) capacitor c=0.00191414f //x=50.51 //y=5.155
c500 ( 73 0 ) capacitor c=0.0903046f //x=95.09 //y=2.08
c501 ( 67 0 ) capacitor c=0.11005f //x=88.43 //y=2.08
c502 ( 65 0 ) capacitor c=0.00669947f //x=88.43 //y=4.54
c503 ( 58 0 ) capacitor c=0.0907522f //x=54.02 //y=2.08
c504 ( 56 0 ) capacitor c=0.103749f //x=52.17 //y=3.33
c505 ( 52 0 ) capacitor c=0.00398962f //x=51.77 //y=1.665
c506 ( 51 0 ) capacitor c=0.0137288f //x=52.085 //y=1.665
c507 ( 45 0 ) capacitor c=0.0276208f //x=52.085 //y=5.155
c508 ( 37 0 ) capacitor c=0.0169868f //x=51.305 //y=5.155
c509 ( 30 0 ) capacitor c=0.00316998f //x=49.715 //y=5.155
c510 ( 29 0 ) capacitor c=0.014258f //x=50.425 //y=5.155
c511 ( 14 0 ) capacitor c=0.00672327f //x=88.545 //y=4.07
c512 ( 13 0 ) capacitor c=0.212984f //x=94.975 //y=4.07
c513 ( 12 0 ) capacitor c=0.004561f //x=65.205 //y=4.07
c514 ( 11 0 ) capacitor c=0.345736f //x=88.315 //y=4.07
c515 ( 10 0 ) capacitor c=0.00784097f //x=65.12 //y=3.985
c516 ( 8 0 ) capacitor c=1.67157e-19 //x=57.065 //y=3.7
c517 ( 7 0 ) capacitor c=0.146519f //x=65.035 //y=3.7
c518 ( 6 0 ) capacitor c=0.0049602f //x=56.98 //y=3.615
c519 ( 4 0 ) capacitor c=0.00349717f //x=54.135 //y=3.33
c520 ( 3 0 ) capacitor c=0.0428789f //x=56.895 //y=3.33
c521 ( 2 0 ) capacitor c=0.00852385f //x=52.285 //y=3.33
c522 ( 1 0 ) capacitor c=0.0280751f //x=53.905 //y=3.33
r523 (  178 179 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=95.11 //y=4.795 //x2=95.11 //y2=4.87
r524 (  176 178 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=95.11 //y=4.705 //x2=95.11 //y2=4.795
r525 (  172 173 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=95.09 //y=2.08 //x2=95.09 //y2=1.915
r526 (  164 166 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=88.47 //y=4.705 //x2=88.47 //y2=4.795
r527 (  160 161 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=88.43 //y=2.08 //x2=88.43 //y2=1.915
r528 (  150 183 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=95.655 //y=1.255 //x2=95.655 //y2=1.367
r529 (  149 182 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=95.655 //y=0.905 //x2=95.615 //y2=0.75
r530 (  149 150 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=95.655 //y=0.905 //x2=95.655 //y2=1.255
r531 (  144 181 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=95.28 //y=1.405 //x2=95.165 //y2=1.405
r532 (  143 183 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=95.5 //y=1.405 //x2=95.655 //y2=1.367
r533 (  142 180 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=95.28 //y=0.75 //x2=95.165 //y2=0.75
r534 (  141 182 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=95.5 //y=0.75 //x2=95.615 //y2=0.75
r535 (  141 142 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=95.5 //y=0.75 //x2=95.28 //y2=0.75
r536 (  140 178 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=95.245 //y=4.795 //x2=95.11 //y2=4.795
r537 (  139 146 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=95.495 //y=4.795 //x2=95.57 //y2=4.87
r538 (  139 140 ) resistor r=128.191 //w=0.094 //l=0.25 //layer=ply \
 //thickness=0.18 //x=95.495 //y=4.795 //x2=95.245 //y2=4.795
r539 (  134 181 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=95.125 //y=1.56 //x2=95.165 //y2=1.405
r540 (  134 173 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=95.125 //y=1.56 //x2=95.125 //y2=1.915
r541 (  133 181 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=95.125 //y=1.255 //x2=95.165 //y2=1.405
r542 (  132 180 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=95.125 //y=0.905 //x2=95.165 //y2=0.75
r543 (  132 133 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=95.125 //y=0.905 //x2=95.125 //y2=1.255
r544 (  131 170 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.995 //y=1.25 //x2=88.955 //y2=1.405
r545 (  130 169 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.995 //y=0.905 //x2=88.955 //y2=0.75
r546 (  130 131 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=88.995 //y=0.905 //x2=88.995 //y2=1.25
r547 (  125 168 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=88.62 //y=1.405 //x2=88.505 //y2=1.405
r548 (  124 170 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=88.84 //y=1.405 //x2=88.955 //y2=1.405
r549 (  123 167 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=88.62 //y=0.75 //x2=88.505 //y2=0.75
r550 (  122 169 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=88.84 //y=0.75 //x2=88.955 //y2=0.75
r551 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=88.84 //y=0.75 //x2=88.62 //y2=0.75
r552 (  121 166 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=88.605 //y=4.795 //x2=88.47 //y2=4.795
r553 (  120 127 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=88.835 //y=4.795 //x2=88.91 //y2=4.87
r554 (  120 121 ) resistor r=117.936 //w=0.094 //l=0.23 //layer=ply \
 //thickness=0.18 //x=88.835 //y=4.795 //x2=88.605 //y2=4.795
r555 (  117 166 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=88.47 //y=4.87 //x2=88.47 //y2=4.795
r556 (  115 168 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.465 //y=1.56 //x2=88.505 //y2=1.405
r557 (  115 161 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=88.465 //y=1.56 //x2=88.465 //y2=1.915
r558 (  114 168 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.465 //y=1.25 //x2=88.505 //y2=1.405
r559 (  113 167 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.465 //y=0.905 //x2=88.505 //y2=0.75
r560 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=88.465 //y=0.905 //x2=88.465 //y2=1.25
r561 (  108 110 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=54.585 //y=4.79 //x2=54.66 //y2=4.865
r562 (  108 109 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=54.585 //y=4.79 //x2=54.295 //y2=4.79
r563 (  107 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.25 //y=1.22 //x2=54.21 //y2=1.375
r564 (  106 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.25 //y=0.875 //x2=54.21 //y2=0.72
r565 (  106 107 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=54.25 //y=0.875 //x2=54.25 //y2=1.22
r566 (  103 109 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=54.22 //y=4.865 //x2=54.295 //y2=4.79
r567 (  103 156 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=54.22 //y=4.865 //x2=54.02 //y2=4.7
r568 (  101 152 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.875 //y=1.375 //x2=53.76 //y2=1.375
r569 (  100 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.095 //y=1.375 //x2=54.21 //y2=1.375
r570 (  99 151 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.875 //y=0.72 //x2=53.76 //y2=0.72
r571 (  98 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.095 //y=0.72 //x2=54.21 //y2=0.72
r572 (  98 99 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=54.095 //y=0.72 //x2=53.875 //y2=0.72
r573 (  97 154 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=53.72 //y=1.915 //x2=54.02 //y2=2.08
r574 (  96 152 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.72 //y=1.53 //x2=53.76 //y2=1.375
r575 (  96 97 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=53.72 //y=1.53 //x2=53.72 //y2=1.915
r576 (  95 152 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.72 //y=1.22 //x2=53.76 //y2=1.375
r577 (  94 151 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.72 //y=0.875 //x2=53.76 //y2=0.72
r578 (  94 95 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=53.72 //y=0.875 //x2=53.72 //y2=1.22
r579 (  93 146 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=95.57 //y=6.025 //x2=95.57 //y2=4.87
r580 (  92 179 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=95.13 //y=6.025 //x2=95.13 //y2=4.87
r581 (  91 127 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=88.91 //y=6.025 //x2=88.91 //y2=4.87
r582 (  90 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=88.47 //y=6.025 //x2=88.47 //y2=4.87
r583 (  89 110 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.66 //y=6.02 //x2=54.66 //y2=4.865
r584 (  88 103 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.22 //y=6.02 //x2=54.22 //y2=4.865
r585 (  87 143 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=95.39 //y=1.405 //x2=95.5 //y2=1.405
r586 (  87 144 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=95.39 //y=1.405 //x2=95.28 //y2=1.405
r587 (  86 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=88.73 //y=1.405 //x2=88.84 //y2=1.405
r588 (  86 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=88.73 //y=1.405 //x2=88.62 //y2=1.405
r589 (  85 100 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.985 //y=1.375 //x2=54.095 //y2=1.375
r590 (  85 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.985 //y=1.375 //x2=53.875 //y2=1.375
r591 (  82 176 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=95.11 //y=4.705 //x2=95.11 //y2=4.705
r592 (  82 83 ) resistor r=10.3507 //w=0.207 //l=0.165 //layer=li \
 //thickness=0.1 //x=95.1 //y=4.705 //x2=95.1 //y2=4.54
r593 (  80 164 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=88.47 //y=4.705 //x2=88.47 //y2=4.705
r594 (  76 83 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=95.09 //y=4.07 //x2=95.09 //y2=4.54
r595 (  73 172 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=95.09 //y=2.08 //x2=95.09 //y2=2.08
r596 (  73 76 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=95.09 //y=2.08 //x2=95.09 //y2=4.07
r597 (  67 160 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=88.43 //y=2.08 //x2=88.43 //y2=2.08
r598 (  67 70 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=88.43 //y=2.08 //x2=88.43 //y2=4.07
r599 (  65 80 ) resistor r=11.2426 //w=0.191 //l=0.174714 //layer=li \
 //thickness=0.1 //x=88.43 //y=4.54 //x2=88.45 //y2=4.705
r600 (  65 70 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=88.43 //y=4.54 //x2=88.43 //y2=4.07
r601 (  63 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.02 //y=4.7 //x2=54.02 //y2=4.7
r602 (  61 63 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=54.02 //y=3.33 //x2=54.02 //y2=4.7
r603 (  58 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.02 //y=2.08 //x2=54.02 //y2=2.08
r604 (  58 61 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=54.02 //y=2.08 //x2=54.02 //y2=3.33
r605 (  54 56 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=52.17 //y=5.07 //x2=52.17 //y2=3.33
r606 (  53 56 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=52.17 //y=1.75 //x2=52.17 //y2=3.33
r607 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=52.085 //y=1.665 //x2=52.17 //y2=1.75
r608 (  51 52 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=52.085 //y=1.665 //x2=51.77 //y2=1.665
r609 (  47 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=51.685 //y=1.58 //x2=51.77 //y2=1.665
r610 (  47 184 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=51.685 //y=1.58 //x2=51.685 //y2=1.01
r611 (  46 78 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.475 //y=5.155 //x2=51.39 //y2=5.155
r612 (  45 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=52.085 //y=5.155 //x2=52.17 //y2=5.07
r613 (  45 46 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=52.085 //y=5.155 //x2=51.475 //y2=5.155
r614 (  39 78 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.39 //y=5.24 //x2=51.39 //y2=5.155
r615 (  39 188 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=51.39 //y=5.24 //x2=51.39 //y2=5.725
r616 (  38 77 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.595 //y=5.155 //x2=50.51 //y2=5.155
r617 (  37 78 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.305 //y=5.155 //x2=51.39 //y2=5.155
r618 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=51.305 //y=5.155 //x2=50.595 //y2=5.155
r619 (  31 77 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.51 //y=5.24 //x2=50.51 //y2=5.155
r620 (  31 187 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.51 //y=5.24 //x2=50.51 //y2=5.725
r621 (  29 77 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.425 //y=5.155 //x2=50.51 //y2=5.155
r622 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.425 //y=5.155 //x2=49.715 //y2=5.155
r623 (  23 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=49.63 //y=5.24 //x2=49.715 //y2=5.155
r624 (  23 186 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=49.63 //y=5.24 //x2=49.63 //y2=5.725
r625 (  22 76 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=95.09 //y=4.07 //x2=95.09 //y2=4.07
r626 (  20 70 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=88.43 //y=4.07 //x2=88.43 //y2=4.07
r627 (  18 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=54.02 //y=3.33 //x2=54.02 //y2=3.33
r628 (  16 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=52.17 //y=3.33 //x2=52.17 //y2=3.33
r629 (  14 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=88.545 //y=4.07 //x2=88.43 //y2=4.07
r630 (  13 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=94.975 //y=4.07 //x2=95.09 //y2=4.07
r631 (  13 14 ) resistor r=6.1355 //w=0.131 //l=6.43 //layer=m1 \
 //thickness=0.36 //x=94.975 //y=4.07 //x2=88.545 //y2=4.07
r632 (  11 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=88.315 //y=4.07 //x2=88.43 //y2=4.07
r633 (  11 12 ) resistor r=22.0515 //w=0.131 //l=23.11 //layer=m1 \
 //thickness=0.36 //x=88.315 //y=4.07 //x2=65.205 //y2=4.07
r634 (  10 12 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=65.12 //y=3.985 //x2=65.205 //y2=4.07
r635 (  9 10 ) resistor r=0.19084 //w=0.131 //l=0.2 //layer=m1 \
 //thickness=0.36 //x=65.12 //y=3.785 //x2=65.12 //y2=3.985
r636 (  7 9 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=65.035 //y=3.7 //x2=65.12 //y2=3.785
r637 (  7 8 ) resistor r=7.60496 //w=0.131 //l=7.97 //layer=m1 \
 //thickness=0.36 //x=65.035 //y=3.7 //x2=57.065 //y2=3.7
r638 (  6 8 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=56.98 //y=3.615 //x2=57.065 //y2=3.7
r639 (  5 6 ) resistor r=0.19084 //w=0.131 //l=0.2 //layer=m1 //thickness=0.36 \
 //x=56.98 //y=3.415 //x2=56.98 //y2=3.615
r640 (  4 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=54.135 //y=3.33 //x2=54.02 //y2=3.33
r641 (  3 5 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=56.895 //y=3.33 //x2=56.98 //y2=3.415
r642 (  3 4 ) resistor r=2.63359 //w=0.131 //l=2.76 //layer=m1 \
 //thickness=0.36 //x=56.895 //y=3.33 //x2=54.135 //y2=3.33
r643 (  2 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=52.285 //y=3.33 //x2=52.17 //y2=3.33
r644 (  1 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=53.905 //y=3.33 //x2=54.02 //y2=3.33
r645 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=53.905 //y=3.33 //x2=52.285 //y2=3.33
ends PM_TMRDFFSNRNQNX1\%noxref_26

subckt PM_TMRDFFSNRNQNX1\%Q ( 1 2 3 4 5 26 27 40 42 43 47 52 53 54 55 59 60 )
c175 ( 60 0 ) capacitor c=0.0167617f //x=95.205 //y=5.025
c176 ( 59 0 ) capacitor c=0.0164812f //x=94.325 //y=5.025
c177 ( 55 0 ) capacitor c=0.0108176f //x=95.2 //y=0.905
c178 ( 54 0 ) capacitor c=0.0131637f //x=91.87 //y=0.905
c179 ( 53 0 ) capacitor c=0.0131367f //x=88.54 //y=0.905
c180 ( 52 0 ) capacitor c=0.00421476f //x=95.35 //y=5.21
c181 ( 47 0 ) capacitor c=0.13039f //x=95.83 //y=4.07
c182 ( 43 0 ) capacitor c=0.00775877f //x=95.475 //y=1.645
c183 ( 42 0 ) capacitor c=0.0161066f //x=95.745 //y=1.645
c184 ( 40 0 ) capacitor c=0.0151634f //x=95.745 //y=5.21
c185 ( 27 0 ) capacitor c=0.0029383f //x=94.555 //y=5.21
c186 ( 26 0 ) capacitor c=0.0155464f //x=95.265 //y=5.21
c187 ( 5 0 ) capacitor c=0.00436966f //x=92.175 //y=1.18
c188 ( 4 0 ) capacitor c=0.069473f //x=95.275 //y=1.18
c189 ( 3 0 ) capacitor c=0.0141674f //x=88.845 //y=1.18
c190 ( 2 0 ) capacitor c=0.0494873f //x=91.945 //y=1.18
c191 ( 1 0 ) capacitor c=0.0241378f //x=95.83 //y=4.07
r192 (  51 53 ) resistor r=13.3953 //w=0.172 //l=0.18 //layer=li \
 //thickness=0.1 //x=88.727 //y=1.18 //x2=88.727 //y2=1
r193 (  45 47 ) resistor r=72.2139 //w=0.187 //l=1.055 //layer=li \
 //thickness=0.1 //x=95.83 //y=5.125 //x2=95.83 //y2=4.07
r194 (  44 47 ) resistor r=160.171 //w=0.187 //l=2.34 //layer=li \
 //thickness=0.1 //x=95.83 //y=1.73 //x2=95.83 //y2=4.07
r195 (  42 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=95.745 //y=1.645 //x2=95.83 //y2=1.73
r196 (  42 43 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=95.745 //y=1.645 //x2=95.475 //y2=1.645
r197 (  41 52 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=95.435 //y=5.21 //x2=95.35 //y2=5.21
r198 (  40 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=95.745 //y=5.21 //x2=95.83 //y2=5.125
r199 (  40 41 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=95.745 //y=5.21 //x2=95.435 //y2=5.21
r200 (  39 55 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=95.39 //y=1.18 //x2=95.39 //y2=1
r201 (  34 43 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=95.39 //y=1.56 //x2=95.475 //y2=1.645
r202 (  34 39 ) resistor r=26.0107 //w=0.187 //l=0.38 //layer=li \
 //thickness=0.1 //x=95.39 //y=1.56 //x2=95.39 //y2=1.18
r203 (  28 52 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=95.35 //y=5.295 //x2=95.35 //y2=5.21
r204 (  28 60 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=95.35 //y=5.295 //x2=95.35 //y2=5.72
r205 (  26 52 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=95.265 //y=5.21 //x2=95.35 //y2=5.21
r206 (  26 27 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=95.265 //y=5.21 //x2=94.555 //y2=5.21
r207 (  20 27 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=94.47 //y=5.295 //x2=94.555 //y2=5.21
r208 (  20 59 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=94.47 //y=5.295 //x2=94.47 //y2=5.72
r209 (  18 54 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=92.06 //y=1.18 //x2=92.06 //y2=1
r210 (  11 39 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=95.39 //y=1.18 //x2=95.39 //y2=1.18
r211 (  9 18 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=92.06 //y=1.18 //x2=92.06 //y2=1.18
r212 (  7 51 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=88.73 //y=1.18 //x2=88.73 //y2=1.18
r213 (  5 9 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=92.175 //y=1.18 //x2=92.06 //y2=1.18
r214 (  4 11 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=95.275 //y=1.18 //x2=95.39 //y2=1.18
r215 (  4 5 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=95.275 //y=1.18 //x2=92.175 //y2=1.18
r216 (  3 7 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=88.845 //y=1.18 //x2=88.73 //y2=1.18
r217 (  2 9 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=91.945 //y=1.18 //x2=92.06 //y2=1.18
r218 (  2 3 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=91.945 //y=1.18 //x2=88.845 //y2=1.18
r219 (  1 47 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=95.83 //y=4.07 //x2=95.83 //y2=4.07
ends PM_TMRDFFSNRNQNX1\%Q

subckt PM_TMRDFFSNRNQNX1\%noxref_28 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0687824f //x=0.455 //y=0.375
c50 ( 17 0 ) capacitor c=0.0213512f //x=2.445 //y=1.59
c51 ( 13 0 ) capacitor c=0.015523f //x=2.445 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c53 ( 5 0 ) capacitor c=0.0204181f //x=1.475 //y=1.59
c54 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_28

subckt PM_TMRDFFSNRNQNX1\%noxref_29 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=2.965 //y=0.375
c53 ( 28 0 ) capacitor c=0.00462395f //x=1.86 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=3.985 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=3.015 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_29

subckt PM_TMRDFFSNRNQNX1\%noxref_30 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=5.265 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=7.255 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=7.255 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=6.37 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=6.285 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=5.4 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=1.59 //x2=6.37 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=1.59 //x2=6.855 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=1.59 //x2=7.34 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=1.59 //x2=6.855 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=0.54 //x2=6.37 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=0.54 //x2=6.855 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=0.54 //x2=7.34 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=0.54 //x2=6.855 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.485 //y=1.59 //x2=5.4 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.485 //y=1.59 //x2=5.885 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.285 //y=1.59 //x2=6.37 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.285 //y=1.59 //x2=5.885 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.4 //y=1.505 //x2=5.4 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.4 //y=1.505 //x2=5.4 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_30

subckt PM_TMRDFFSNRNQNX1\%noxref_31 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=7.775 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=6.67 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=7.91 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=8.88 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=8.795 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=7.91 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=7.825 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.995 //y=0.54 //x2=7.91 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.995 //y=0.54 //x2=8.395 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.795 //y=0.54 //x2=8.88 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.795 //y=0.54 //x2=8.395 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.945 //y=0.995 //x2=6.86 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=7.91 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=6.945 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_31

subckt PM_TMRDFFSNRNQNX1\%noxref_32 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=10.075 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=12.065 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=12.065 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=11.18 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=11.095 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=10.21 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.265 //y=1.59 //x2=11.18 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.265 //y=1.59 //x2=11.665 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.065 //y=1.59 //x2=12.15 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.065 //y=1.59 //x2=11.665 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.265 //y=0.54 //x2=11.18 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.265 //y=0.54 //x2=11.665 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.065 //y=0.54 //x2=12.15 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.065 //y=0.54 //x2=11.665 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=11.18 //y=1.505 //x2=11.18 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=11.18 //y=1.505 //x2=11.18 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.18 //y=0.625 //x2=11.18 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.18 //y=0.625 //x2=11.18 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.295 //y=1.59 //x2=10.21 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.295 //y=1.59 //x2=10.695 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.095 //y=1.59 //x2=11.18 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.095 //y=1.59 //x2=10.695 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=10.21 //y=1.505 //x2=10.21 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.21 //y=1.505 //x2=10.21 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_32

subckt PM_TMRDFFSNRNQNX1\%noxref_33 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=12.585 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=11.48 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=12.72 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=13.69 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=13.605 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=12.72 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=12.635 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=13.69 //y=0.625 //x2=13.69 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=13.69 //y=0.625 //x2=13.69 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.805 //y=0.54 //x2=12.72 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.805 //y=0.54 //x2=13.205 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.605 //y=0.54 //x2=13.69 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.605 //y=0.54 //x2=13.205 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.72 //y=1.08 //x2=12.72 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=12.72 //y=1.08 //x2=12.72 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.91 //x2=12.72 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.91 //x2=12.72 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.625 //x2=12.72 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.625 //x2=12.72 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.755 //y=0.995 //x2=11.67 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.635 //y=0.995 //x2=12.72 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=12.635 //y=0.995 //x2=11.755 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_33

subckt PM_TMRDFFSNRNQNX1\%noxref_34 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=14.885 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=16.875 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=16.875 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=15.99 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=15.905 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=15.02 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.075 //y=1.59 //x2=15.99 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.075 //y=1.59 //x2=16.475 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.875 //y=1.59 //x2=16.96 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.875 //y=1.59 //x2=16.475 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.075 //y=0.54 //x2=15.99 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.075 //y=0.54 //x2=16.475 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.875 //y=0.54 //x2=16.96 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.875 //y=0.54 //x2=16.475 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=15.99 //y=1.505 //x2=15.99 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.99 //y=1.505 //x2=15.99 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.99 //y=0.625 //x2=15.99 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=15.99 //y=0.625 //x2=15.99 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.105 //y=1.59 //x2=15.02 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.105 //y=1.59 //x2=15.505 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.905 //y=1.59 //x2=15.99 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.905 //y=1.59 //x2=15.505 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.02 //y=1.505 //x2=15.02 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.02 //y=1.505 //x2=15.02 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_34

subckt PM_TMRDFFSNRNQNX1\%noxref_35 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=17.395 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=16.29 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=17.53 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=18.5 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=18.415 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=17.53 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=17.445 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=18.5 //y=0.625 //x2=18.5 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.5 //y=0.625 //x2=18.5 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.615 //y=0.54 //x2=17.53 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.615 //y=0.54 //x2=18.015 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.415 //y=0.54 //x2=18.5 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.415 //y=0.54 //x2=18.015 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.53 //y=1.08 //x2=17.53 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=17.53 //y=1.08 //x2=17.53 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.91 //x2=17.53 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.91 //x2=17.53 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.625 //x2=17.53 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.625 //x2=17.53 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.565 //y=0.995 //x2=16.48 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.445 //y=0.995 //x2=17.53 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=17.445 //y=0.995 //x2=16.565 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_35

subckt PM_TMRDFFSNRNQNX1\%noxref_36 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=19.695 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=21.685 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=21.685 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=20.8 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=20.715 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=19.83 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.885 //y=1.59 //x2=20.8 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.885 //y=1.59 //x2=21.285 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.685 //y=1.59 //x2=21.77 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.685 //y=1.59 //x2=21.285 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.885 //y=0.54 //x2=20.8 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.885 //y=0.54 //x2=21.285 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.685 //y=0.54 //x2=21.77 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.685 //y=0.54 //x2=21.285 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=20.8 //y=1.505 //x2=20.8 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=20.8 //y=1.505 //x2=20.8 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.8 //y=0.625 //x2=20.8 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=20.8 //y=0.625 //x2=20.8 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.915 //y=1.59 //x2=19.83 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.915 //y=1.59 //x2=20.315 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.715 //y=1.59 //x2=20.8 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.715 //y=1.59 //x2=20.315 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=19.83 //y=1.505 //x2=19.83 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=19.83 //y=1.505 //x2=19.83 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_36

subckt PM_TMRDFFSNRNQNX1\%noxref_37 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=22.205 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=21.1 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=22.34 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=23.31 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=23.225 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=22.34 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=22.255 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.31 //y=0.625 //x2=23.31 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=23.31 //y=0.625 //x2=23.31 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.425 //y=0.54 //x2=22.34 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.425 //y=0.54 //x2=22.825 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.225 //y=0.54 //x2=23.31 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.225 //y=0.54 //x2=22.825 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.34 //y=1.08 //x2=22.34 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=22.34 //y=1.08 //x2=22.34 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.91 //x2=22.34 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.91 //x2=22.34 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.625 //x2=22.34 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.625 //x2=22.34 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.375 //y=0.995 //x2=21.29 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.255 //y=0.995 //x2=22.34 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=22.255 //y=0.995 //x2=21.375 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_37

subckt PM_TMRDFFSNRNQNX1\%noxref_38 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=24.505 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=26.495 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=26.495 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=25.61 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=25.525 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=24.64 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.695 //y=1.59 //x2=25.61 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.695 //y=1.59 //x2=26.095 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.495 //y=1.59 //x2=26.58 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.495 //y=1.59 //x2=26.095 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.695 //y=0.54 //x2=25.61 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.695 //y=0.54 //x2=26.095 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.495 //y=0.54 //x2=26.58 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.495 //y=0.54 //x2=26.095 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=25.61 //y=1.505 //x2=25.61 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=25.61 //y=1.505 //x2=25.61 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=25.61 //y=0.625 //x2=25.61 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=25.61 //y=0.625 //x2=25.61 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.725 //y=1.59 //x2=24.64 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.725 //y=1.59 //x2=25.125 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.525 //y=1.59 //x2=25.61 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.525 //y=1.59 //x2=25.125 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=24.64 //y=1.505 //x2=24.64 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=24.64 //y=1.505 //x2=24.64 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_38

subckt PM_TMRDFFSNRNQNX1\%noxref_39 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=27.015 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=25.91 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=27.15 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=28.12 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=28.035 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=27.15 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=27.065 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=28.12 //y=0.625 //x2=28.12 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=28.12 //y=0.625 //x2=28.12 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=27.235 //y=0.54 //x2=27.15 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=27.235 //y=0.54 //x2=27.635 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=28.035 //y=0.54 //x2=28.12 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.035 //y=0.54 //x2=27.635 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.15 //y=1.08 //x2=27.15 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=27.15 //y=1.08 //x2=27.15 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.91 //x2=27.15 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.91 //x2=27.15 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.625 //x2=27.15 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.625 //x2=27.15 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.185 //y=0.995 //x2=26.1 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.065 //y=0.995 //x2=27.15 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=27.065 //y=0.995 //x2=26.185 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_39

subckt PM_TMRDFFSNRNQNX1\%noxref_40 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=29.315 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=31.305 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=31.305 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=30.42 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=30.335 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=29.45 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.505 //y=1.59 //x2=30.42 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.505 //y=1.59 //x2=30.905 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.305 //y=1.59 //x2=31.39 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=31.305 //y=1.59 //x2=30.905 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.505 //y=0.54 //x2=30.42 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.505 //y=0.54 //x2=30.905 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.305 //y=0.54 //x2=31.39 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=31.305 //y=0.54 //x2=30.905 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=30.42 //y=1.505 //x2=30.42 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=30.42 //y=1.505 //x2=30.42 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=30.42 //y=0.625 //x2=30.42 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=30.42 //y=0.625 //x2=30.42 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.535 //y=1.59 //x2=29.45 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.535 //y=1.59 //x2=29.935 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.335 //y=1.59 //x2=30.42 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.335 //y=1.59 //x2=29.935 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=29.45 //y=1.505 //x2=29.45 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=29.45 //y=1.505 //x2=29.45 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_40

subckt PM_TMRDFFSNRNQNX1\%noxref_41 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=31.825 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=30.72 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=31.96 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=32.93 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=32.845 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=31.96 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=31.875 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=32.93 //y=0.625 //x2=32.93 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=32.93 //y=0.625 //x2=32.93 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=32.045 //y=0.54 //x2=31.96 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=32.045 //y=0.54 //x2=32.445 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=32.845 //y=0.54 //x2=32.93 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=32.845 //y=0.54 //x2=32.445 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=31.96 //y=1.08 //x2=31.96 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=31.96 //y=1.08 //x2=31.96 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=31.96 //y=0.91 //x2=31.96 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=31.96 //y=0.91 //x2=31.96 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=31.96 //y=0.625 //x2=31.96 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=31.96 //y=0.625 //x2=31.96 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.995 //y=0.995 //x2=30.91 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=31.875 //y=0.995 //x2=31.96 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=31.875 //y=0.995 //x2=30.995 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_41

subckt PM_TMRDFFSNRNQNX1\%noxref_42 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=34.125 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=36.115 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=36.115 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=35.23 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=35.145 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=34.26 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=35.315 //y=1.59 //x2=35.23 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.315 //y=1.59 //x2=35.715 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.115 //y=1.59 //x2=36.2 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=36.115 //y=1.59 //x2=35.715 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=35.315 //y=0.54 //x2=35.23 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.315 //y=0.54 //x2=35.715 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.115 //y=0.54 //x2=36.2 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=36.115 //y=0.54 //x2=35.715 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=35.23 //y=1.505 //x2=35.23 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=35.23 //y=1.505 //x2=35.23 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=35.23 //y=0.625 //x2=35.23 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=35.23 //y=0.625 //x2=35.23 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.345 //y=1.59 //x2=34.26 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.345 //y=1.59 //x2=34.745 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=35.145 //y=1.59 //x2=35.23 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.145 //y=1.59 //x2=34.745 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=34.26 //y=1.505 //x2=34.26 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=34.26 //y=1.505 //x2=34.26 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_42

subckt PM_TMRDFFSNRNQNX1\%noxref_43 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=36.635 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=35.53 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=36.77 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=37.74 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=37.655 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=36.77 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=36.685 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=37.74 //y=0.625 //x2=37.74 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=37.74 //y=0.625 //x2=37.74 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=36.855 //y=0.54 //x2=36.77 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=36.855 //y=0.54 //x2=37.255 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=37.655 //y=0.54 //x2=37.74 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=37.655 //y=0.54 //x2=37.255 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=36.77 //y=1.08 //x2=36.77 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=36.77 //y=1.08 //x2=36.77 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=36.77 //y=0.91 //x2=36.77 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=36.77 //y=0.91 //x2=36.77 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=36.77 //y=0.625 //x2=36.77 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=36.77 //y=0.625 //x2=36.77 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.805 //y=0.995 //x2=35.72 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=36.685 //y=0.995 //x2=36.77 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=36.685 //y=0.995 //x2=35.805 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_43

subckt PM_TMRDFFSNRNQNX1\%noxref_44 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=38.935 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=40.925 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=40.925 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=40.04 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=39.955 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=39.07 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=40.125 //y=1.59 //x2=40.04 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.125 //y=1.59 //x2=40.525 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.925 //y=1.59 //x2=41.01 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.925 //y=1.59 //x2=40.525 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=40.125 //y=0.54 //x2=40.04 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.125 //y=0.54 //x2=40.525 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.925 //y=0.54 //x2=41.01 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.925 //y=0.54 //x2=40.525 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=40.04 //y=1.505 //x2=40.04 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=40.04 //y=1.505 //x2=40.04 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=40.04 //y=0.625 //x2=40.04 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=40.04 //y=0.625 //x2=40.04 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=39.155 //y=1.59 //x2=39.07 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=39.155 //y=1.59 //x2=39.555 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=39.955 //y=1.59 //x2=40.04 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=39.955 //y=1.59 //x2=39.555 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=39.07 //y=1.505 //x2=39.07 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=39.07 //y=1.505 //x2=39.07 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_44

subckt PM_TMRDFFSNRNQNX1\%noxref_45 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=41.445 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=40.34 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=41.58 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=42.55 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=42.465 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=41.58 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=41.495 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=42.55 //y=0.625 //x2=42.55 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=42.55 //y=0.625 //x2=42.55 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=41.665 //y=0.54 //x2=41.58 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=41.665 //y=0.54 //x2=42.065 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=42.465 //y=0.54 //x2=42.55 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=42.465 //y=0.54 //x2=42.065 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=41.58 //y=1.08 //x2=41.58 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=41.58 //y=1.08 //x2=41.58 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=41.58 //y=0.91 //x2=41.58 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=41.58 //y=0.91 //x2=41.58 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=41.58 //y=0.625 //x2=41.58 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=41.58 //y=0.625 //x2=41.58 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.615 //y=0.995 //x2=40.53 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=41.495 //y=0.995 //x2=41.58 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=41.495 //y=0.995 //x2=40.615 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_45

subckt PM_TMRDFFSNRNQNX1\%noxref_46 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=43.745 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=45.735 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=45.735 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=44.85 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=44.765 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=43.88 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.935 //y=1.59 //x2=44.85 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.935 //y=1.59 //x2=45.335 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.735 //y=1.59 //x2=45.82 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.735 //y=1.59 //x2=45.335 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.935 //y=0.54 //x2=44.85 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.935 //y=0.54 //x2=45.335 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.735 //y=0.54 //x2=45.82 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.735 //y=0.54 //x2=45.335 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=44.85 //y=1.505 //x2=44.85 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=44.85 //y=1.505 //x2=44.85 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=44.85 //y=0.625 //x2=44.85 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=44.85 //y=0.625 //x2=44.85 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=43.965 //y=1.59 //x2=43.88 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=43.965 //y=1.59 //x2=44.365 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.765 //y=1.59 //x2=44.85 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.765 //y=1.59 //x2=44.365 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=43.88 //y=1.505 //x2=43.88 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=43.88 //y=1.505 //x2=43.88 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_46

subckt PM_TMRDFFSNRNQNX1\%noxref_47 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=46.255 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=45.15 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=46.39 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=47.36 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=47.275 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=46.39 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=46.305 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=47.36 //y=0.625 //x2=47.36 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=47.36 //y=0.625 //x2=47.36 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=46.475 //y=0.54 //x2=46.39 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.475 //y=0.54 //x2=46.875 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=47.275 //y=0.54 //x2=47.36 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=47.275 //y=0.54 //x2=46.875 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.39 //y=1.08 //x2=46.39 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=46.39 //y=1.08 //x2=46.39 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.39 //y=0.91 //x2=46.39 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=46.39 //y=0.91 //x2=46.39 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=46.39 //y=0.625 //x2=46.39 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=46.39 //y=0.625 //x2=46.39 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.425 //y=0.995 //x2=45.34 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.305 //y=0.995 //x2=46.39 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=46.305 //y=0.995 //x2=45.425 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_47

subckt PM_TMRDFFSNRNQNX1\%noxref_48 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=48.555 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=50.545 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=50.545 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=49.66 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=49.575 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=48.69 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.745 //y=1.59 //x2=49.66 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.745 //y=1.59 //x2=50.145 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.545 //y=1.59 //x2=50.63 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.545 //y=1.59 //x2=50.145 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.745 //y=0.54 //x2=49.66 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.745 //y=0.54 //x2=50.145 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.545 //y=0.54 //x2=50.63 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.545 //y=0.54 //x2=50.145 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=49.66 //y=1.505 //x2=49.66 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=49.66 //y=1.505 //x2=49.66 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=49.66 //y=0.625 //x2=49.66 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=49.66 //y=0.625 //x2=49.66 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=48.775 //y=1.59 //x2=48.69 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=48.775 //y=1.59 //x2=49.175 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.575 //y=1.59 //x2=49.66 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.575 //y=1.59 //x2=49.175 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=48.69 //y=1.505 //x2=48.69 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=48.69 //y=1.505 //x2=48.69 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_48

subckt PM_TMRDFFSNRNQNX1\%noxref_49 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=51.065 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=49.96 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=51.2 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=52.17 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=52.085 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=51.2 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=51.115 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=52.17 //y=0.625 //x2=52.17 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=52.17 //y=0.625 //x2=52.17 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=51.285 //y=0.54 //x2=51.2 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=51.285 //y=0.54 //x2=51.685 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=52.085 //y=0.54 //x2=52.17 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=52.085 //y=0.54 //x2=51.685 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=51.2 //y=1.08 //x2=51.2 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=51.2 //y=1.08 //x2=51.2 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=51.2 //y=0.91 //x2=51.2 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=51.2 //y=0.91 //x2=51.2 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=51.2 //y=0.625 //x2=51.2 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=51.2 //y=0.625 //x2=51.2 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.235 //y=0.995 //x2=50.15 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=51.115 //y=0.995 //x2=51.2 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=51.115 //y=0.995 //x2=50.235 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_49

subckt PM_TMRDFFSNRNQNX1\%noxref_50 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=53.365 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=55.355 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=55.355 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=54.47 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=54.385 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=53.5 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=54.555 //y=1.59 //x2=54.47 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.555 //y=1.59 //x2=54.955 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.355 //y=1.59 //x2=55.44 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=55.355 //y=1.59 //x2=54.955 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=54.555 //y=0.54 //x2=54.47 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.555 //y=0.54 //x2=54.955 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.355 //y=0.54 //x2=55.44 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=55.355 //y=0.54 //x2=54.955 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=54.47 //y=1.505 //x2=54.47 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=54.47 //y=1.505 //x2=54.47 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=54.47 //y=0.625 //x2=54.47 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=54.47 //y=0.625 //x2=54.47 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.585 //y=1.59 //x2=53.5 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.585 //y=1.59 //x2=53.985 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=54.385 //y=1.59 //x2=54.47 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.385 //y=1.59 //x2=53.985 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=53.5 //y=1.505 //x2=53.5 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=53.5 //y=1.505 //x2=53.5 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_50

subckt PM_TMRDFFSNRNQNX1\%noxref_51 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=55.875 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=54.77 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=56.01 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=56.98 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=56.895 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=56.01 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=55.925 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=56.98 //y=0.625 //x2=56.98 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=56.98 //y=0.625 //x2=56.98 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=56.095 //y=0.54 //x2=56.01 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=56.095 //y=0.54 //x2=56.495 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=56.895 //y=0.54 //x2=56.98 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=56.895 //y=0.54 //x2=56.495 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=56.01 //y=1.08 //x2=56.01 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=56.01 //y=1.08 //x2=56.01 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=56.01 //y=0.91 //x2=56.01 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=56.01 //y=0.91 //x2=56.01 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=56.01 //y=0.625 //x2=56.01 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=56.01 //y=0.625 //x2=56.01 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.045 //y=0.995 //x2=54.96 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=55.925 //y=0.995 //x2=56.01 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=55.925 //y=0.995 //x2=55.045 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_51

subckt PM_TMRDFFSNRNQNX1\%noxref_52 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=58.175 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=60.165 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=60.165 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=59.28 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=59.195 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=58.31 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=59.365 //y=1.59 //x2=59.28 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.365 //y=1.59 //x2=59.765 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.165 //y=1.59 //x2=60.25 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.165 //y=1.59 //x2=59.765 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=59.365 //y=0.54 //x2=59.28 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.365 //y=0.54 //x2=59.765 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.165 //y=0.54 //x2=60.25 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.165 //y=0.54 //x2=59.765 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=59.28 //y=1.505 //x2=59.28 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=59.28 //y=1.505 //x2=59.28 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=59.28 //y=0.625 //x2=59.28 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=59.28 //y=0.625 //x2=59.28 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.395 //y=1.59 //x2=58.31 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.395 //y=1.59 //x2=58.795 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=59.195 //y=1.59 //x2=59.28 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.195 //y=1.59 //x2=58.795 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=58.31 //y=1.505 //x2=58.31 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=58.31 //y=1.505 //x2=58.31 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_52

subckt PM_TMRDFFSNRNQNX1\%noxref_53 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=60.685 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=59.58 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=60.82 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=61.79 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=61.705 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=60.82 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=60.735 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=61.79 //y=0.625 //x2=61.79 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=61.79 //y=0.625 //x2=61.79 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=60.905 //y=0.54 //x2=60.82 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.905 //y=0.54 //x2=61.305 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=61.705 //y=0.54 //x2=61.79 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=61.705 //y=0.54 //x2=61.305 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.82 //y=1.08 //x2=60.82 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=60.82 //y=1.08 //x2=60.82 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.82 //y=0.91 //x2=60.82 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=60.82 //y=0.91 //x2=60.82 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=60.82 //y=0.625 //x2=60.82 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=60.82 //y=0.625 //x2=60.82 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.855 //y=0.995 //x2=59.77 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.735 //y=0.995 //x2=60.82 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=60.735 //y=0.995 //x2=59.855 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_53

subckt PM_TMRDFFSNRNQNX1\%noxref_54 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=62.985 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=64.975 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=64.975 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=64.09 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=64.005 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=63.12 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=64.175 //y=1.59 //x2=64.09 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.175 //y=1.59 //x2=64.575 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.975 //y=1.59 //x2=65.06 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.975 //y=1.59 //x2=64.575 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=64.175 //y=0.54 //x2=64.09 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.175 //y=0.54 //x2=64.575 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.975 //y=0.54 //x2=65.06 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.975 //y=0.54 //x2=64.575 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=64.09 //y=1.505 //x2=64.09 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=64.09 //y=1.505 //x2=64.09 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=64.09 //y=0.625 //x2=64.09 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=64.09 //y=0.625 //x2=64.09 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63.205 //y=1.59 //x2=63.12 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63.205 //y=1.59 //x2=63.605 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=64.005 //y=1.59 //x2=64.09 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.005 //y=1.59 //x2=63.605 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=63.12 //y=1.505 //x2=63.12 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=63.12 //y=1.505 //x2=63.12 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_54

subckt PM_TMRDFFSNRNQNX1\%noxref_55 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=65.495 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=64.39 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=65.63 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=66.6 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=66.515 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=65.63 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=65.545 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=66.6 //y=0.625 //x2=66.6 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=66.6 //y=0.625 //x2=66.6 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=65.715 //y=0.54 //x2=65.63 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=65.715 //y=0.54 //x2=66.115 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.515 //y=0.54 //x2=66.6 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=66.515 //y=0.54 //x2=66.115 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=65.63 //y=1.08 //x2=65.63 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=65.63 //y=1.08 //x2=65.63 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=65.63 //y=0.91 //x2=65.63 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=65.63 //y=0.91 //x2=65.63 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=65.63 //y=0.625 //x2=65.63 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=65.63 //y=0.625 //x2=65.63 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.665 //y=0.995 //x2=64.58 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=65.545 //y=0.995 //x2=65.63 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=65.545 //y=0.995 //x2=64.665 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_55

subckt PM_TMRDFFSNRNQNX1\%noxref_56 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=67.795 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=69.785 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=69.785 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=68.9 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=68.815 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=67.93 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.985 //y=1.59 //x2=68.9 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.985 //y=1.59 //x2=69.385 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.785 //y=1.59 //x2=69.87 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.785 //y=1.59 //x2=69.385 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.985 //y=0.54 //x2=68.9 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.985 //y=0.54 //x2=69.385 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.785 //y=0.54 //x2=69.87 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.785 //y=0.54 //x2=69.385 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=68.9 //y=1.505 //x2=68.9 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=68.9 //y=1.505 //x2=68.9 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=68.9 //y=0.625 //x2=68.9 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=68.9 //y=0.625 //x2=68.9 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.015 //y=1.59 //x2=67.93 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.015 //y=1.59 //x2=68.415 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.815 //y=1.59 //x2=68.9 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.815 //y=1.59 //x2=68.415 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=67.93 //y=1.505 //x2=67.93 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=67.93 //y=1.505 //x2=67.93 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_56

subckt PM_TMRDFFSNRNQNX1\%noxref_57 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=70.305 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=69.2 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=70.44 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=71.41 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=71.325 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=70.44 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=70.355 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=71.41 //y=0.625 //x2=71.41 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=71.41 //y=0.625 //x2=71.41 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=70.525 //y=0.54 //x2=70.44 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.525 //y=0.54 //x2=70.925 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=71.325 //y=0.54 //x2=71.41 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=71.325 //y=0.54 //x2=70.925 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=70.44 //y=1.08 //x2=70.44 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=70.44 //y=1.08 //x2=70.44 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=70.44 //y=0.91 //x2=70.44 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=70.44 //y=0.91 //x2=70.44 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=70.44 //y=0.625 //x2=70.44 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=70.44 //y=0.625 //x2=70.44 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.475 //y=0.995 //x2=69.39 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=70.355 //y=0.995 //x2=70.44 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=70.355 //y=0.995 //x2=69.475 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_57

subckt PM_TMRDFFSNRNQNX1\%noxref_58 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=72.605 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=74.595 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=74.595 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=73.71 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=73.625 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=72.74 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=73.795 //y=1.59 //x2=73.71 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=73.795 //y=1.59 //x2=74.195 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.595 //y=1.59 //x2=74.68 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=74.595 //y=1.59 //x2=74.195 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=73.795 //y=0.54 //x2=73.71 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=73.795 //y=0.54 //x2=74.195 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.595 //y=0.54 //x2=74.68 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=74.595 //y=0.54 //x2=74.195 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=73.71 //y=1.505 //x2=73.71 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=73.71 //y=1.505 //x2=73.71 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=73.71 //y=0.625 //x2=73.71 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=73.71 //y=0.625 //x2=73.71 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=72.825 //y=1.59 //x2=72.74 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=72.825 //y=1.59 //x2=73.225 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=73.625 //y=1.59 //x2=73.71 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=73.625 //y=1.59 //x2=73.225 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=72.74 //y=1.505 //x2=72.74 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=72.74 //y=1.505 //x2=72.74 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_58

subckt PM_TMRDFFSNRNQNX1\%noxref_59 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=75.115 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=74.01 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=75.25 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=76.22 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=76.135 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=75.25 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=75.165 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=76.22 //y=0.625 //x2=76.22 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=76.22 //y=0.625 //x2=76.22 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.335 //y=0.54 //x2=75.25 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=75.335 //y=0.54 //x2=75.735 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=76.135 //y=0.54 //x2=76.22 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=76.135 //y=0.54 //x2=75.735 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=75.25 //y=1.08 //x2=75.25 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=75.25 //y=1.08 //x2=75.25 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=75.25 //y=0.91 //x2=75.25 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=75.25 //y=0.91 //x2=75.25 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=75.25 //y=0.625 //x2=75.25 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=75.25 //y=0.625 //x2=75.25 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.285 //y=0.995 //x2=74.2 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=75.165 //y=0.995 //x2=75.25 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=75.165 //y=0.995 //x2=74.285 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_59

subckt PM_TMRDFFSNRNQNX1\%noxref_60 ( 1 5 9 13 17 35 )
c51 ( 35 0 ) capacitor c=0.0680259f //x=77.415 //y=0.375
c52 ( 17 0 ) capacitor c=0.0180446f //x=79.405 //y=1.59
c53 ( 13 0 ) capacitor c=0.0155283f //x=79.405 //y=0.54
c54 ( 9 0 ) capacitor c=0.00678203f //x=78.52 //y=0.625
c55 ( 5 0 ) capacitor c=0.0164013f //x=78.435 //y=1.59
c56 ( 1 0 ) capacitor c=0.00696517f //x=77.55 //y=1.505
r57 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.605 //y=1.59 //x2=78.52 //y2=1.63
r58 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.605 //y=1.59 //x2=79.005 //y2=1.59
r59 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.405 //y=1.59 //x2=79.49 //y2=1.59
r60 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=79.405 //y=1.59 //x2=79.005 //y2=1.59
r61 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.605 //y=0.54 //x2=78.52 //y2=0.5
r62 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.605 //y=0.54 //x2=79.005 //y2=0.54
r63 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.405 //y=0.54 //x2=79.49 //y2=0.54
r64 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=79.405 //y=0.54 //x2=79.005 //y2=0.54
r65 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=78.52 //y=1.505 //x2=78.52 //y2=1.63
r66 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=78.52 //y=1.505 //x2=78.52 //y2=0.89
r67 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=78.52 //y=0.625 //x2=78.52 //y2=0.5
r68 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=78.52 //y=0.625 //x2=78.52 //y2=0.89
r69 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=77.635 //y=1.59 //x2=77.55 //y2=1.63
r70 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=77.635 //y=1.59 //x2=78.035 //y2=1.59
r71 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.435 //y=1.59 //x2=78.52 //y2=1.63
r72 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.435 //y=1.59 //x2=78.035 //y2=1.59
r73 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=77.55 //y=1.505 //x2=77.55 //y2=1.63
r74 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=77.55 //y=1.505 //x2=77.55 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_60

subckt PM_TMRDFFSNRNQNX1\%noxref_61 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0420321f //x=79.925 //y=0.375
c55 ( 28 0 ) capacitor c=0.00457437f //x=78.82 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=80.06 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=81.03 //y=0.625
c58 ( 11 0 ) capacitor c=0.0145658f //x=80.945 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=80.06 //y=0.625
c60 ( 1 0 ) capacitor c=0.0234159f //x=79.975 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=81.03 //y=0.625 //x2=81.03 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=81.03 //y=0.625 //x2=81.03 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=80.145 //y=0.54 //x2=80.06 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=80.145 //y=0.54 //x2=80.545 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=80.945 //y=0.54 //x2=81.03 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=80.945 //y=0.54 //x2=80.545 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=80.06 //y=1.08 //x2=80.06 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=80.06 //y=1.08 //x2=80.06 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=80.06 //y=0.91 //x2=80.06 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=80.06 //y=0.91 //x2=80.06 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=80.06 //y=0.625 //x2=80.06 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=80.06 //y=0.625 //x2=80.06 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.095 //y=0.995 //x2=79.01 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=79.975 //y=0.995 //x2=80.06 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=79.975 //y=0.995 //x2=79.095 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_61

subckt PM_TMRDFFSNRNQNX1\%noxref_62 ( 1 5 9 13 17 35 )
c51 ( 35 0 ) capacitor c=0.0673029f //x=82.225 //y=0.375
c52 ( 17 0 ) capacitor c=0.0178317f //x=84.215 //y=1.59
c53 ( 13 0 ) capacitor c=0.0154936f //x=84.215 //y=0.54
c54 ( 9 0 ) capacitor c=0.00678203f //x=83.33 //y=0.625
c55 ( 5 0 ) capacitor c=0.0163955f //x=83.245 //y=1.59
c56 ( 1 0 ) capacitor c=0.00696517f //x=82.36 //y=1.505
r57 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=83.415 //y=1.59 //x2=83.33 //y2=1.63
r58 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=83.415 //y=1.59 //x2=83.815 //y2=1.59
r59 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.215 //y=1.59 //x2=84.3 //y2=1.59
r60 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=84.215 //y=1.59 //x2=83.815 //y2=1.59
r61 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=83.415 //y=0.54 //x2=83.33 //y2=0.5
r62 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=83.415 //y=0.54 //x2=83.815 //y2=0.54
r63 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.215 //y=0.54 //x2=84.3 //y2=0.54
r64 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=84.215 //y=0.54 //x2=83.815 //y2=0.54
r65 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=83.33 //y=1.505 //x2=83.33 //y2=1.63
r66 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=83.33 //y=1.505 //x2=83.33 //y2=0.89
r67 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=83.33 //y=0.625 //x2=83.33 //y2=0.5
r68 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=83.33 //y=0.625 //x2=83.33 //y2=0.89
r69 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=82.445 //y=1.59 //x2=82.36 //y2=1.63
r70 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=82.445 //y=1.59 //x2=82.845 //y2=1.59
r71 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=83.245 //y=1.59 //x2=83.33 //y2=1.63
r72 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=83.245 //y=1.59 //x2=82.845 //y2=1.59
r73 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=82.36 //y=1.505 //x2=82.36 //y2=1.63
r74 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=82.36 //y=1.505 //x2=82.36 //y2=0.89
ends PM_TMRDFFSNRNQNX1\%noxref_62

subckt PM_TMRDFFSNRNQNX1\%noxref_63 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.041346f //x=84.735 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=83.63 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=84.87 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=85.84 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=85.755 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=84.87 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=84.785 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=85.84 //y=0.625 //x2=85.84 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=85.84 //y=0.625 //x2=85.84 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=84.955 //y=0.54 //x2=84.87 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=84.955 //y=0.54 //x2=85.355 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=85.755 //y=0.54 //x2=85.84 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=85.755 //y=0.54 //x2=85.355 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=84.87 //y=1.08 //x2=84.87 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=84.87 //y=1.08 //x2=84.87 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=84.87 //y=0.91 //x2=84.87 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=84.87 //y=0.91 //x2=84.87 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=84.87 //y=0.625 //x2=84.87 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=84.87 //y=0.625 //x2=84.87 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.905 //y=0.995 //x2=83.82 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=84.785 //y=0.995 //x2=84.87 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=84.785 //y=0.995 //x2=83.905 //y2=0.995
ends PM_TMRDFFSNRNQNX1\%noxref_63

subckt PM_TMRDFFSNRNQNX1\%noxref_64 ( 1 5 9 10 13 17 29 )
c57 ( 29 0 ) capacitor c=0.0751624f //x=87.14 //y=0.365
c58 ( 17 0 ) capacitor c=0.0072249f //x=89.215 //y=0.615
c59 ( 13 0 ) capacitor c=0.0152499f //x=89.13 //y=0.53
c60 ( 10 0 ) capacitor c=0.00698291f //x=88.245 //y=1.495
c61 ( 9 0 ) capacitor c=0.006761f //x=88.245 //y=0.615
c62 ( 5 0 ) capacitor c=0.0191191f //x=88.16 //y=1.58
c63 ( 1 0 ) capacitor c=0.00483164f //x=87.275 //y=1.495
r64 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=89.215 //y=0.615 //x2=89.215 //y2=0.49
r65 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=89.215 //y=0.615 //x2=89.215 //y2=1.22
r66 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=88.33 //y=0.53 //x2=88.245 //y2=0.49
r67 (  14 29 ) resistor r=27.0374 //w=0.187 //l=0.395 //layer=li \
 //thickness=0.1 //x=88.33 //y=0.53 //x2=88.725 //y2=0.53
r68 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=89.13 //y=0.53 //x2=89.215 //y2=0.49
r69 (  13 29 ) resistor r=27.7219 //w=0.187 //l=0.405 //layer=li \
 //thickness=0.1 //x=89.13 //y=0.53 //x2=88.725 //y2=0.53
r70 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=88.245 //y=1.495 //x2=88.245 //y2=1.62
r71 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=88.245 //y=1.495 //x2=88.245 //y2=0.88
r72 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=88.245 //y=0.615 //x2=88.245 //y2=0.49
r73 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=88.245 //y=0.615 //x2=88.245 //y2=0.88
r74 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=87.36 //y=1.58 //x2=87.275 //y2=1.62
r75 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=87.36 //y=1.58 //x2=87.76 //y2=1.58
r76 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=88.16 //y=1.58 //x2=88.245 //y2=1.62
r77 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=88.16 //y=1.58 //x2=87.76 //y2=1.58
r78 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=87.275 //y=1.495 //x2=87.275 //y2=1.62
r79 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=87.275 //y=1.495 //x2=87.275 //y2=0.88
ends PM_TMRDFFSNRNQNX1\%noxref_64

subckt PM_TMRDFFSNRNQNX1\%noxref_65 ( 1 5 9 10 13 17 29 )
c55 ( 29 0 ) capacitor c=0.0723103f //x=90.47 //y=0.365
c56 ( 17 0 ) capacitor c=0.0072249f //x=92.545 //y=0.615
c57 ( 13 0 ) capacitor c=0.0155051f //x=92.46 //y=0.53
c58 ( 10 0 ) capacitor c=0.00811719f //x=91.575 //y=1.495
c59 ( 9 0 ) capacitor c=0.006761f //x=91.575 //y=0.615
c60 ( 5 0 ) capacitor c=0.0166789f //x=91.49 //y=1.58
c61 ( 1 0 ) capacitor c=0.00788388f //x=90.605 //y=1.495
r62 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=92.545 //y=0.615 //x2=92.545 //y2=0.49
r63 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=92.545 //y=0.615 //x2=92.545 //y2=1.22
r64 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=91.66 //y=0.53 //x2=91.575 //y2=0.49
r65 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=91.66 //y=0.53 //x2=92.06 //y2=0.53
r66 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=92.46 //y=0.53 //x2=92.545 //y2=0.49
r67 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=92.46 //y=0.53 //x2=92.06 //y2=0.53
r68 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=91.575 //y=1.495 //x2=91.575 //y2=1.62
r69 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=91.575 //y=1.495 //x2=91.575 //y2=0.88
r70 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=91.575 //y=0.615 //x2=91.575 //y2=0.49
r71 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=91.575 //y=0.615 //x2=91.575 //y2=0.88
r72 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=90.69 //y=1.58 //x2=90.605 //y2=1.62
r73 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=90.69 //y=1.58 //x2=91.09 //y2=1.58
r74 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=91.49 //y=1.58 //x2=91.575 //y2=1.62
r75 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=91.49 //y=1.58 //x2=91.09 //y2=1.58
r76 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=90.605 //y=1.495 //x2=90.605 //y2=1.62
r77 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=90.605 //y=1.495 //x2=90.605 //y2=0.88
ends PM_TMRDFFSNRNQNX1\%noxref_65

subckt PM_TMRDFFSNRNQNX1\%noxref_66 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0637439f //x=93.8 //y=0.365
c55 ( 17 0 ) capacitor c=0.00722228f //x=95.875 //y=0.615
c56 ( 13 0 ) capacitor c=0.0141607f //x=95.79 //y=0.53
c57 ( 10 0 ) capacitor c=0.00712138f //x=94.905 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=94.905 //y=0.615
c59 ( 5 0 ) capacitor c=0.0233454f //x=94.82 //y=1.58
c60 ( 1 0 ) capacitor c=0.00481264f //x=93.935 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=95.875 //y=0.615 //x2=95.875 //y2=0.49
r62 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=95.875 //y=0.615 //x2=95.875 //y2=0.88
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=94.99 //y=0.53 //x2=94.905 //y2=0.49
r64 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=94.99 //y=0.53 //x2=95.39 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=95.79 //y=0.53 //x2=95.875 //y2=0.49
r66 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=95.79 //y=0.53 //x2=95.39 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=94.905 //y=1.495 //x2=94.905 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=94.905 //y=1.495 //x2=94.905 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=94.905 //y=0.615 //x2=94.905 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=94.905 //y=0.615 //x2=94.905 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=94.02 //y=1.58 //x2=93.935 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=94.02 //y=1.58 //x2=94.42 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=94.82 //y=1.58 //x2=94.905 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=94.82 //y=1.58 //x2=94.42 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=93.935 //y=1.495 //x2=93.935 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=93.935 //y=1.495 //x2=93.935 //y2=0.88
ends PM_TMRDFFSNRNQNX1\%noxref_66

