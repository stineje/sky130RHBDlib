magic
tech sky130A
magscale 1 2
timestamp 1669564325
<< nwell >>
rect -87 786 19401 1550
<< pwell >>
rect -34 -34 19348 544
<< nmos >>
rect 147 290 177 351
tri 177 290 193 306 sw
rect 447 290 477 351
rect 147 260 253 290
tri 253 260 283 290 sw
rect 147 159 177 260
tri 177 244 193 260 nw
tri 237 244 253 260 ne
tri 177 159 193 175 sw
tri 237 159 253 175 se
rect 253 159 283 260
tri 342 260 372 290 se
rect 372 260 477 290
rect 342 166 372 260
tri 372 244 388 260 nw
tri 431 244 447 260 ne
tri 372 166 388 182 sw
tri 431 166 447 182 se
rect 447 166 477 260
tri 147 129 177 159 ne
rect 177 129 253 159
tri 253 129 283 159 nw
tri 342 136 372 166 ne
rect 372 136 447 166
tri 447 136 477 166 nw
rect 649 298 679 351
tri 679 298 695 314 sw
rect 649 268 755 298
tri 755 268 785 298 sw
rect 649 167 679 268
tri 679 252 695 268 nw
tri 739 252 755 268 ne
tri 679 167 695 183 sw
tri 739 167 755 183 se
rect 755 167 785 268
tri 649 137 679 167 ne
rect 679 137 755 167
tri 755 137 785 167 nw
rect 1109 290 1139 351
tri 1139 290 1155 306 sw
rect 1409 290 1439 351
rect 1109 260 1215 290
tri 1215 260 1245 290 sw
rect 1109 159 1139 260
tri 1139 244 1155 260 nw
tri 1199 244 1215 260 ne
tri 1139 159 1155 175 sw
tri 1199 159 1215 175 se
rect 1215 159 1245 260
tri 1304 260 1334 290 se
rect 1334 260 1439 290
rect 1304 166 1334 260
tri 1334 244 1350 260 nw
tri 1393 244 1409 260 ne
tri 1334 166 1350 182 sw
tri 1393 166 1409 182 se
rect 1409 166 1439 260
tri 1109 129 1139 159 ne
rect 1139 129 1215 159
tri 1215 129 1245 159 nw
tri 1304 136 1334 166 ne
rect 1334 136 1409 166
tri 1409 136 1439 166 nw
rect 1611 298 1641 351
tri 1641 298 1657 314 sw
rect 1611 268 1717 298
tri 1717 268 1747 298 sw
rect 1611 167 1641 268
tri 1641 252 1657 268 nw
tri 1701 252 1717 268 ne
tri 1641 167 1657 183 sw
tri 1701 167 1717 183 se
rect 1717 167 1747 268
tri 1611 137 1641 167 ne
rect 1641 137 1717 167
tri 1717 137 1747 167 nw
rect 2071 290 2101 351
tri 2101 290 2117 306 sw
rect 2371 290 2401 351
rect 2071 260 2177 290
tri 2177 260 2207 290 sw
rect 2071 159 2101 260
tri 2101 244 2117 260 nw
tri 2161 244 2177 260 ne
tri 2101 159 2117 175 sw
tri 2161 159 2177 175 se
rect 2177 159 2207 260
tri 2266 260 2296 290 se
rect 2296 260 2401 290
rect 2266 166 2296 260
tri 2296 244 2312 260 nw
tri 2355 244 2371 260 ne
tri 2296 166 2312 182 sw
tri 2355 166 2371 182 se
rect 2371 166 2401 260
tri 2071 129 2101 159 ne
rect 2101 129 2177 159
tri 2177 129 2207 159 nw
tri 2266 136 2296 166 ne
rect 2296 136 2371 166
tri 2371 136 2401 166 nw
rect 2573 298 2603 351
tri 2603 298 2619 314 sw
rect 2573 268 2679 298
tri 2679 268 2709 298 sw
rect 2573 167 2603 268
tri 2603 252 2619 268 nw
tri 2663 252 2679 268 ne
tri 2603 167 2619 183 sw
tri 2663 167 2679 183 se
rect 2679 167 2709 268
tri 2573 137 2603 167 ne
rect 2603 137 2679 167
tri 2679 137 2709 167 nw
rect 3033 290 3063 351
tri 3063 290 3079 306 sw
rect 3333 290 3363 351
rect 3033 260 3139 290
tri 3139 260 3169 290 sw
rect 3033 159 3063 260
tri 3063 244 3079 260 nw
tri 3123 244 3139 260 ne
tri 3063 159 3079 175 sw
tri 3123 159 3139 175 se
rect 3139 159 3169 260
tri 3228 260 3258 290 se
rect 3258 260 3363 290
rect 3228 166 3258 260
tri 3258 244 3274 260 nw
tri 3317 244 3333 260 ne
tri 3258 166 3274 182 sw
tri 3317 166 3333 182 se
rect 3333 166 3363 260
tri 3033 129 3063 159 ne
rect 3063 129 3139 159
tri 3139 129 3169 159 nw
tri 3228 136 3258 166 ne
rect 3258 136 3333 166
tri 3333 136 3363 166 nw
rect 3535 298 3565 351
tri 3565 298 3581 314 sw
rect 3535 268 3641 298
tri 3641 268 3671 298 sw
rect 3535 167 3565 268
tri 3565 252 3581 268 nw
tri 3625 252 3641 268 ne
tri 3565 167 3581 183 sw
tri 3625 167 3641 183 se
rect 3641 167 3671 268
tri 3535 137 3565 167 ne
rect 3565 137 3641 167
tri 3641 137 3671 167 nw
rect 3995 290 4025 351
tri 4025 290 4041 306 sw
rect 4295 290 4325 351
rect 3995 260 4101 290
tri 4101 260 4131 290 sw
rect 3995 159 4025 260
tri 4025 244 4041 260 nw
tri 4085 244 4101 260 ne
tri 4025 159 4041 175 sw
tri 4085 159 4101 175 se
rect 4101 159 4131 260
tri 4190 260 4220 290 se
rect 4220 260 4325 290
rect 4190 166 4220 260
tri 4220 244 4236 260 nw
tri 4279 244 4295 260 ne
tri 4220 166 4236 182 sw
tri 4279 166 4295 182 se
rect 4295 166 4325 260
tri 3995 129 4025 159 ne
rect 4025 129 4101 159
tri 4101 129 4131 159 nw
tri 4190 136 4220 166 ne
rect 4220 136 4295 166
tri 4295 136 4325 166 nw
rect 4497 298 4527 351
tri 4527 298 4543 314 sw
rect 4497 268 4603 298
tri 4603 268 4633 298 sw
rect 4497 167 4527 268
tri 4527 252 4543 268 nw
tri 4587 252 4603 268 ne
tri 4527 167 4543 183 sw
tri 4587 167 4603 183 se
rect 4603 167 4633 268
tri 4497 137 4527 167 ne
rect 4527 137 4603 167
tri 4603 137 4633 167 nw
rect 4957 290 4987 351
tri 4987 290 5003 306 sw
rect 5257 290 5287 351
rect 4957 260 5063 290
tri 5063 260 5093 290 sw
rect 4957 159 4987 260
tri 4987 244 5003 260 nw
tri 5047 244 5063 260 ne
tri 4987 159 5003 175 sw
tri 5047 159 5063 175 se
rect 5063 159 5093 260
tri 5152 260 5182 290 se
rect 5182 260 5287 290
rect 5152 166 5182 260
tri 5182 244 5198 260 nw
tri 5241 244 5257 260 ne
tri 5182 166 5198 182 sw
tri 5241 166 5257 182 se
rect 5257 166 5287 260
tri 4957 129 4987 159 ne
rect 4987 129 5063 159
tri 5063 129 5093 159 nw
tri 5152 136 5182 166 ne
rect 5182 136 5257 166
tri 5257 136 5287 166 nw
rect 5459 298 5489 351
tri 5489 298 5505 314 sw
rect 5459 268 5565 298
tri 5565 268 5595 298 sw
rect 5459 167 5489 268
tri 5489 252 5505 268 nw
tri 5549 252 5565 268 ne
tri 5489 167 5505 183 sw
tri 5549 167 5565 183 se
rect 5565 167 5595 268
tri 5459 137 5489 167 ne
rect 5489 137 5565 167
tri 5565 137 5595 167 nw
rect 5919 290 5949 351
tri 5949 290 5965 306 sw
rect 6219 290 6249 351
rect 5919 260 6025 290
tri 6025 260 6055 290 sw
rect 5919 159 5949 260
tri 5949 244 5965 260 nw
tri 6009 244 6025 260 ne
tri 5949 159 5965 175 sw
tri 6009 159 6025 175 se
rect 6025 159 6055 260
tri 6114 260 6144 290 se
rect 6144 260 6249 290
rect 6114 166 6144 260
tri 6144 244 6160 260 nw
tri 6203 244 6219 260 ne
tri 6144 166 6160 182 sw
tri 6203 166 6219 182 se
rect 6219 166 6249 260
tri 5919 129 5949 159 ne
rect 5949 129 6025 159
tri 6025 129 6055 159 nw
tri 6114 136 6144 166 ne
rect 6144 136 6219 166
tri 6219 136 6249 166 nw
rect 6421 298 6451 351
tri 6451 298 6467 314 sw
rect 6421 268 6527 298
tri 6527 268 6557 298 sw
rect 6421 167 6451 268
tri 6451 252 6467 268 nw
tri 6511 252 6527 268 ne
tri 6451 167 6467 183 sw
tri 6511 167 6527 183 se
rect 6527 167 6557 268
tri 6421 137 6451 167 ne
rect 6451 137 6527 167
tri 6527 137 6557 167 nw
rect 6881 290 6911 351
tri 6911 290 6927 306 sw
rect 7181 290 7211 351
rect 6881 260 6987 290
tri 6987 260 7017 290 sw
rect 6881 159 6911 260
tri 6911 244 6927 260 nw
tri 6971 244 6987 260 ne
tri 6911 159 6927 175 sw
tri 6971 159 6987 175 se
rect 6987 159 7017 260
tri 7076 260 7106 290 se
rect 7106 260 7211 290
rect 7076 166 7106 260
tri 7106 244 7122 260 nw
tri 7165 244 7181 260 ne
tri 7106 166 7122 182 sw
tri 7165 166 7181 182 se
rect 7181 166 7211 260
tri 6881 129 6911 159 ne
rect 6911 129 6987 159
tri 6987 129 7017 159 nw
tri 7076 136 7106 166 ne
rect 7106 136 7181 166
tri 7181 136 7211 166 nw
rect 7383 298 7413 351
tri 7413 298 7429 314 sw
rect 7383 268 7489 298
tri 7489 268 7519 298 sw
rect 7383 167 7413 268
tri 7413 252 7429 268 nw
tri 7473 252 7489 268 ne
tri 7413 167 7429 183 sw
tri 7473 167 7489 183 se
rect 7489 167 7519 268
tri 7383 137 7413 167 ne
rect 7413 137 7489 167
tri 7489 137 7519 167 nw
rect 7843 290 7873 351
tri 7873 290 7889 306 sw
rect 8143 290 8173 351
rect 7843 260 7949 290
tri 7949 260 7979 290 sw
rect 7843 159 7873 260
tri 7873 244 7889 260 nw
tri 7933 244 7949 260 ne
tri 7873 159 7889 175 sw
tri 7933 159 7949 175 se
rect 7949 159 7979 260
tri 8038 260 8068 290 se
rect 8068 260 8173 290
rect 8038 166 8068 260
tri 8068 244 8084 260 nw
tri 8127 244 8143 260 ne
tri 8068 166 8084 182 sw
tri 8127 166 8143 182 se
rect 8143 166 8173 260
tri 7843 129 7873 159 ne
rect 7873 129 7949 159
tri 7949 129 7979 159 nw
tri 8038 136 8068 166 ne
rect 8068 136 8143 166
tri 8143 136 8173 166 nw
rect 8345 298 8375 351
tri 8375 298 8391 314 sw
rect 8345 268 8451 298
tri 8451 268 8481 298 sw
rect 8345 167 8375 268
tri 8375 252 8391 268 nw
tri 8435 252 8451 268 ne
tri 8375 167 8391 183 sw
tri 8435 167 8451 183 se
rect 8451 167 8481 268
tri 8345 137 8375 167 ne
rect 8375 137 8451 167
tri 8451 137 8481 167 nw
rect 8805 290 8835 351
tri 8835 290 8851 306 sw
rect 9105 290 9135 351
rect 8805 260 8911 290
tri 8911 260 8941 290 sw
rect 8805 159 8835 260
tri 8835 244 8851 260 nw
tri 8895 244 8911 260 ne
tri 8835 159 8851 175 sw
tri 8895 159 8911 175 se
rect 8911 159 8941 260
tri 9000 260 9030 290 se
rect 9030 260 9135 290
rect 9000 166 9030 260
tri 9030 244 9046 260 nw
tri 9089 244 9105 260 ne
tri 9030 166 9046 182 sw
tri 9089 166 9105 182 se
rect 9105 166 9135 260
tri 8805 129 8835 159 ne
rect 8835 129 8911 159
tri 8911 129 8941 159 nw
tri 9000 136 9030 166 ne
rect 9030 136 9105 166
tri 9105 136 9135 166 nw
rect 9307 298 9337 351
tri 9337 298 9353 314 sw
rect 9307 268 9413 298
tri 9413 268 9443 298 sw
rect 9307 167 9337 268
tri 9337 252 9353 268 nw
tri 9397 252 9413 268 ne
tri 9337 167 9353 183 sw
tri 9397 167 9413 183 se
rect 9413 167 9443 268
tri 9307 137 9337 167 ne
rect 9337 137 9413 167
tri 9413 137 9443 167 nw
rect 9767 290 9797 351
tri 9797 290 9813 306 sw
rect 10067 290 10097 351
rect 9767 260 9873 290
tri 9873 260 9903 290 sw
rect 9767 159 9797 260
tri 9797 244 9813 260 nw
tri 9857 244 9873 260 ne
tri 9797 159 9813 175 sw
tri 9857 159 9873 175 se
rect 9873 159 9903 260
tri 9962 260 9992 290 se
rect 9992 260 10097 290
rect 9962 166 9992 260
tri 9992 244 10008 260 nw
tri 10051 244 10067 260 ne
tri 9992 166 10008 182 sw
tri 10051 166 10067 182 se
rect 10067 166 10097 260
tri 9767 129 9797 159 ne
rect 9797 129 9873 159
tri 9873 129 9903 159 nw
tri 9962 136 9992 166 ne
rect 9992 136 10067 166
tri 10067 136 10097 166 nw
rect 10269 298 10299 351
tri 10299 298 10315 314 sw
rect 10269 268 10375 298
tri 10375 268 10405 298 sw
rect 10269 167 10299 268
tri 10299 252 10315 268 nw
tri 10359 252 10375 268 ne
tri 10299 167 10315 183 sw
tri 10359 167 10375 183 se
rect 10375 167 10405 268
tri 10269 137 10299 167 ne
rect 10299 137 10375 167
tri 10375 137 10405 167 nw
rect 10729 290 10759 351
tri 10759 290 10775 306 sw
rect 11029 290 11059 351
rect 10729 260 10835 290
tri 10835 260 10865 290 sw
rect 10729 159 10759 260
tri 10759 244 10775 260 nw
tri 10819 244 10835 260 ne
tri 10759 159 10775 175 sw
tri 10819 159 10835 175 se
rect 10835 159 10865 260
tri 10924 260 10954 290 se
rect 10954 260 11059 290
rect 10924 166 10954 260
tri 10954 244 10970 260 nw
tri 11013 244 11029 260 ne
tri 10954 166 10970 182 sw
tri 11013 166 11029 182 se
rect 11029 166 11059 260
tri 10729 129 10759 159 ne
rect 10759 129 10835 159
tri 10835 129 10865 159 nw
tri 10924 136 10954 166 ne
rect 10954 136 11029 166
tri 11029 136 11059 166 nw
rect 11231 298 11261 351
tri 11261 298 11277 314 sw
rect 11231 268 11337 298
tri 11337 268 11367 298 sw
rect 11231 167 11261 268
tri 11261 252 11277 268 nw
tri 11321 252 11337 268 ne
tri 11261 167 11277 183 sw
tri 11321 167 11337 183 se
rect 11337 167 11367 268
tri 11231 137 11261 167 ne
rect 11261 137 11337 167
tri 11337 137 11367 167 nw
rect 11691 290 11721 351
tri 11721 290 11737 306 sw
rect 11991 290 12021 351
rect 11691 260 11797 290
tri 11797 260 11827 290 sw
rect 11691 159 11721 260
tri 11721 244 11737 260 nw
tri 11781 244 11797 260 ne
tri 11721 159 11737 175 sw
tri 11781 159 11797 175 se
rect 11797 159 11827 260
tri 11886 260 11916 290 se
rect 11916 260 12021 290
rect 11886 166 11916 260
tri 11916 244 11932 260 nw
tri 11975 244 11991 260 ne
tri 11916 166 11932 182 sw
tri 11975 166 11991 182 se
rect 11991 166 12021 260
tri 11691 129 11721 159 ne
rect 11721 129 11797 159
tri 11797 129 11827 159 nw
tri 11886 136 11916 166 ne
rect 11916 136 11991 166
tri 11991 136 12021 166 nw
rect 12193 298 12223 351
tri 12223 298 12239 314 sw
rect 12193 268 12299 298
tri 12299 268 12329 298 sw
rect 12193 167 12223 268
tri 12223 252 12239 268 nw
tri 12283 252 12299 268 ne
tri 12223 167 12239 183 sw
tri 12283 167 12299 183 se
rect 12299 167 12329 268
tri 12193 137 12223 167 ne
rect 12223 137 12299 167
tri 12299 137 12329 167 nw
rect 12653 290 12683 351
tri 12683 290 12699 306 sw
rect 12953 290 12983 351
rect 12653 260 12759 290
tri 12759 260 12789 290 sw
rect 12653 159 12683 260
tri 12683 244 12699 260 nw
tri 12743 244 12759 260 ne
tri 12683 159 12699 175 sw
tri 12743 159 12759 175 se
rect 12759 159 12789 260
tri 12848 260 12878 290 se
rect 12878 260 12983 290
rect 12848 166 12878 260
tri 12878 244 12894 260 nw
tri 12937 244 12953 260 ne
tri 12878 166 12894 182 sw
tri 12937 166 12953 182 se
rect 12953 166 12983 260
tri 12653 129 12683 159 ne
rect 12683 129 12759 159
tri 12759 129 12789 159 nw
tri 12848 136 12878 166 ne
rect 12878 136 12953 166
tri 12953 136 12983 166 nw
rect 13155 298 13185 351
tri 13185 298 13201 314 sw
rect 13155 268 13261 298
tri 13261 268 13291 298 sw
rect 13155 167 13185 268
tri 13185 252 13201 268 nw
tri 13245 252 13261 268 ne
tri 13185 167 13201 183 sw
tri 13245 167 13261 183 se
rect 13261 167 13291 268
tri 13155 137 13185 167 ne
rect 13185 137 13261 167
tri 13261 137 13291 167 nw
rect 13615 290 13645 351
tri 13645 290 13661 306 sw
rect 13915 290 13945 351
rect 13615 260 13721 290
tri 13721 260 13751 290 sw
rect 13615 159 13645 260
tri 13645 244 13661 260 nw
tri 13705 244 13721 260 ne
tri 13645 159 13661 175 sw
tri 13705 159 13721 175 se
rect 13721 159 13751 260
tri 13810 260 13840 290 se
rect 13840 260 13945 290
rect 13810 166 13840 260
tri 13840 244 13856 260 nw
tri 13899 244 13915 260 ne
tri 13840 166 13856 182 sw
tri 13899 166 13915 182 se
rect 13915 166 13945 260
tri 13615 129 13645 159 ne
rect 13645 129 13721 159
tri 13721 129 13751 159 nw
tri 13810 136 13840 166 ne
rect 13840 136 13915 166
tri 13915 136 13945 166 nw
rect 14117 298 14147 351
tri 14147 298 14163 314 sw
rect 14117 268 14223 298
tri 14223 268 14253 298 sw
rect 14117 167 14147 268
tri 14147 252 14163 268 nw
tri 14207 252 14223 268 ne
tri 14147 167 14163 183 sw
tri 14207 167 14223 183 se
rect 14223 167 14253 268
tri 14117 137 14147 167 ne
rect 14147 137 14223 167
tri 14223 137 14253 167 nw
rect 14577 290 14607 351
tri 14607 290 14623 306 sw
rect 14877 290 14907 351
rect 14577 260 14683 290
tri 14683 260 14713 290 sw
rect 14577 159 14607 260
tri 14607 244 14623 260 nw
tri 14667 244 14683 260 ne
tri 14607 159 14623 175 sw
tri 14667 159 14683 175 se
rect 14683 159 14713 260
tri 14772 260 14802 290 se
rect 14802 260 14907 290
rect 14772 166 14802 260
tri 14802 244 14818 260 nw
tri 14861 244 14877 260 ne
tri 14802 166 14818 182 sw
tri 14861 166 14877 182 se
rect 14877 166 14907 260
tri 14577 129 14607 159 ne
rect 14607 129 14683 159
tri 14683 129 14713 159 nw
tri 14772 136 14802 166 ne
rect 14802 136 14877 166
tri 14877 136 14907 166 nw
rect 15079 298 15109 351
tri 15109 298 15125 314 sw
rect 15079 268 15185 298
tri 15185 268 15215 298 sw
rect 15079 167 15109 268
tri 15109 252 15125 268 nw
tri 15169 252 15185 268 ne
tri 15109 167 15125 183 sw
tri 15169 167 15185 183 se
rect 15185 167 15215 268
tri 15079 137 15109 167 ne
rect 15109 137 15185 167
tri 15185 137 15215 167 nw
rect 15539 290 15569 351
tri 15569 290 15585 306 sw
rect 15839 290 15869 351
rect 15539 260 15645 290
tri 15645 260 15675 290 sw
rect 15539 159 15569 260
tri 15569 244 15585 260 nw
tri 15629 244 15645 260 ne
tri 15569 159 15585 175 sw
tri 15629 159 15645 175 se
rect 15645 159 15675 260
tri 15734 260 15764 290 se
rect 15764 260 15869 290
rect 15734 166 15764 260
tri 15764 244 15780 260 nw
tri 15823 244 15839 260 ne
tri 15764 166 15780 182 sw
tri 15823 166 15839 182 se
rect 15839 166 15869 260
tri 15539 129 15569 159 ne
rect 15569 129 15645 159
tri 15645 129 15675 159 nw
tri 15734 136 15764 166 ne
rect 15764 136 15839 166
tri 15839 136 15869 166 nw
rect 16041 298 16071 351
tri 16071 298 16087 314 sw
rect 16041 268 16147 298
tri 16147 268 16177 298 sw
rect 16041 167 16071 268
tri 16071 252 16087 268 nw
tri 16131 252 16147 268 ne
tri 16071 167 16087 183 sw
tri 16131 167 16147 183 se
rect 16147 167 16177 268
tri 16041 137 16071 167 ne
rect 16071 137 16147 167
tri 16147 137 16177 167 nw
rect 16501 290 16531 351
tri 16531 290 16547 306 sw
rect 16801 290 16831 351
rect 16501 260 16607 290
tri 16607 260 16637 290 sw
rect 16501 159 16531 260
tri 16531 244 16547 260 nw
tri 16591 244 16607 260 ne
tri 16531 159 16547 175 sw
tri 16591 159 16607 175 se
rect 16607 159 16637 260
tri 16696 260 16726 290 se
rect 16726 260 16831 290
rect 16696 166 16726 260
tri 16726 244 16742 260 nw
tri 16785 244 16801 260 ne
tri 16726 166 16742 182 sw
tri 16785 166 16801 182 se
rect 16801 166 16831 260
tri 16501 129 16531 159 ne
rect 16531 129 16607 159
tri 16607 129 16637 159 nw
tri 16696 136 16726 166 ne
rect 16726 136 16801 166
tri 16801 136 16831 166 nw
rect 17003 298 17033 351
tri 17033 298 17049 314 sw
rect 17003 268 17109 298
tri 17109 268 17139 298 sw
rect 17003 167 17033 268
tri 17033 252 17049 268 nw
tri 17093 252 17109 268 ne
tri 17033 167 17049 183 sw
tri 17093 167 17109 183 se
rect 17109 167 17139 268
tri 17003 137 17033 167 ne
rect 17033 137 17109 167
tri 17109 137 17139 167 nw
rect 17484 288 17514 349
tri 17514 288 17530 304 sw
rect 17678 296 17708 349
tri 17708 296 17724 312 sw
rect 17484 258 17590 288
tri 17590 258 17620 288 sw
rect 17678 266 17784 296
tri 17784 266 17814 296 sw
rect 17484 157 17514 258
tri 17514 242 17530 258 nw
tri 17574 242 17590 258 ne
tri 17514 157 17530 173 sw
tri 17574 157 17590 173 se
rect 17590 157 17620 258
rect 17678 165 17708 266
tri 17708 250 17724 266 nw
tri 17768 250 17784 266 ne
tri 17708 165 17724 181 sw
tri 17768 165 17784 181 se
rect 17784 165 17814 266
tri 17484 127 17514 157 ne
rect 17514 127 17590 157
tri 17590 127 17620 157 nw
tri 17678 135 17708 165 ne
rect 17708 135 17784 165
tri 17784 135 17814 165 nw
rect 18150 288 18180 349
tri 18180 288 18196 304 sw
tri 18434 296 18450 312 se
rect 18450 296 18480 349
rect 18150 258 18256 288
tri 18256 258 18286 288 sw
tri 18344 266 18374 296 se
rect 18374 266 18480 296
rect 18150 157 18180 258
tri 18180 242 18196 258 nw
tri 18240 242 18256 258 ne
tri 18180 157 18196 173 sw
tri 18240 157 18256 173 se
rect 18256 157 18286 258
rect 18344 165 18374 266
tri 18374 250 18390 266 nw
tri 18434 250 18450 266 ne
tri 18374 165 18390 181 sw
tri 18434 165 18450 181 se
rect 18450 165 18480 266
tri 18150 127 18180 157 ne
rect 18180 127 18256 157
tri 18256 127 18286 157 nw
tri 18344 135 18374 165 ne
rect 18374 135 18450 165
tri 18450 135 18480 165 nw
rect 18816 288 18846 349
tri 18846 288 18862 304 sw
rect 19010 296 19040 349
tri 19040 296 19056 312 sw
rect 18816 258 18922 288
tri 18922 258 18952 288 sw
rect 19010 266 19116 296
tri 19116 266 19146 296 sw
rect 18816 157 18846 258
tri 18846 242 18862 258 nw
tri 18906 242 18922 258 ne
tri 18846 157 18862 173 sw
tri 18906 157 18922 173 se
rect 18922 157 18952 258
rect 19010 251 19041 266
tri 19041 251 19056 266 nw
tri 19100 251 19115 266 ne
rect 19115 251 19146 266
rect 19010 165 19040 251
tri 19040 165 19056 181 sw
tri 19100 165 19116 181 se
rect 19116 165 19146 251
tri 18816 127 18846 157 ne
rect 18846 127 18922 157
tri 18922 127 18952 157 nw
tri 19010 135 19040 165 ne
rect 19040 135 19116 165
tri 19116 135 19146 165 nw
<< pmos >>
rect 247 1004 277 1404
rect 335 1004 365 1404
rect 423 1004 453 1404
rect 511 1004 541 1404
rect 599 1004 629 1404
rect 687 1004 717 1404
rect 1209 1004 1239 1404
rect 1297 1004 1327 1404
rect 1385 1004 1415 1404
rect 1473 1004 1503 1404
rect 1561 1004 1591 1404
rect 1649 1004 1679 1404
rect 2171 1004 2201 1404
rect 2259 1004 2289 1404
rect 2347 1004 2377 1404
rect 2435 1004 2465 1404
rect 2523 1004 2553 1404
rect 2611 1004 2641 1404
rect 3133 1004 3163 1404
rect 3221 1004 3251 1404
rect 3309 1004 3339 1404
rect 3397 1004 3427 1404
rect 3485 1004 3515 1404
rect 3573 1004 3603 1404
rect 4095 1004 4125 1404
rect 4183 1004 4213 1404
rect 4271 1004 4301 1404
rect 4359 1004 4389 1404
rect 4447 1004 4477 1404
rect 4535 1004 4565 1404
rect 5057 1004 5087 1404
rect 5145 1004 5175 1404
rect 5233 1004 5263 1404
rect 5321 1004 5351 1404
rect 5409 1004 5439 1404
rect 5497 1004 5527 1404
rect 6019 1004 6049 1404
rect 6107 1004 6137 1404
rect 6195 1004 6225 1404
rect 6283 1004 6313 1404
rect 6371 1004 6401 1404
rect 6459 1004 6489 1404
rect 6981 1004 7011 1404
rect 7069 1004 7099 1404
rect 7157 1004 7187 1404
rect 7245 1004 7275 1404
rect 7333 1004 7363 1404
rect 7421 1004 7451 1404
rect 7943 1004 7973 1404
rect 8031 1004 8061 1404
rect 8119 1004 8149 1404
rect 8207 1004 8237 1404
rect 8295 1004 8325 1404
rect 8383 1004 8413 1404
rect 8905 1004 8935 1404
rect 8993 1004 9023 1404
rect 9081 1004 9111 1404
rect 9169 1004 9199 1404
rect 9257 1004 9287 1404
rect 9345 1004 9375 1404
rect 9867 1004 9897 1404
rect 9955 1004 9985 1404
rect 10043 1004 10073 1404
rect 10131 1004 10161 1404
rect 10219 1004 10249 1404
rect 10307 1004 10337 1404
rect 10829 1004 10859 1404
rect 10917 1004 10947 1404
rect 11005 1004 11035 1404
rect 11093 1004 11123 1404
rect 11181 1004 11211 1404
rect 11269 1004 11299 1404
rect 11791 1004 11821 1404
rect 11879 1004 11909 1404
rect 11967 1004 11997 1404
rect 12055 1004 12085 1404
rect 12143 1004 12173 1404
rect 12231 1004 12261 1404
rect 12753 1004 12783 1404
rect 12841 1004 12871 1404
rect 12929 1004 12959 1404
rect 13017 1004 13047 1404
rect 13105 1004 13135 1404
rect 13193 1004 13223 1404
rect 13715 1004 13745 1404
rect 13803 1004 13833 1404
rect 13891 1004 13921 1404
rect 13979 1004 14009 1404
rect 14067 1004 14097 1404
rect 14155 1004 14185 1404
rect 14677 1004 14707 1404
rect 14765 1004 14795 1404
rect 14853 1004 14883 1404
rect 14941 1004 14971 1404
rect 15029 1004 15059 1404
rect 15117 1004 15147 1404
rect 15639 1004 15669 1404
rect 15727 1004 15757 1404
rect 15815 1004 15845 1404
rect 15903 1004 15933 1404
rect 15991 1004 16021 1404
rect 16079 1004 16109 1404
rect 16601 1004 16631 1404
rect 16689 1004 16719 1404
rect 16777 1004 16807 1404
rect 16865 1004 16895 1404
rect 16953 1004 16983 1404
rect 17041 1004 17071 1404
rect 17503 1005 17533 1405
rect 17591 1005 17621 1405
rect 17679 1005 17709 1405
rect 17767 1005 17797 1405
rect 18167 1005 18197 1405
rect 18255 1005 18285 1405
rect 18343 1005 18373 1405
rect 18431 1005 18461 1405
rect 18835 1005 18865 1405
rect 18923 1005 18953 1405
rect 19011 1005 19041 1405
rect 19099 1005 19129 1405
<< ndiff >>
rect 91 335 147 351
rect 91 301 101 335
rect 135 301 147 335
rect 91 263 147 301
rect 177 335 447 351
rect 177 306 198 335
tri 177 290 193 306 ne
rect 193 301 198 306
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 447 335
rect 193 290 447 301
rect 477 335 533 351
rect 477 301 489 335
rect 523 301 533 335
rect 91 229 101 263
rect 135 229 147 263
tri 253 260 283 290 ne
rect 283 263 342 290
rect 91 195 147 229
rect 91 161 101 195
rect 135 161 147 195
rect 91 129 147 161
tri 177 244 193 260 se
rect 193 244 237 260
tri 237 244 253 260 sw
rect 177 210 253 244
rect 177 176 198 210
rect 232 176 253 210
rect 177 175 253 176
tri 177 159 193 175 ne
rect 193 159 237 175
tri 237 159 253 175 nw
rect 283 229 295 263
rect 329 229 342 263
tri 342 260 372 290 nw
rect 283 195 342 229
rect 283 161 295 195
rect 329 161 342 195
tri 372 244 388 260 se
rect 388 244 431 260
tri 431 244 447 260 sw
rect 372 216 447 244
rect 372 182 393 216
rect 427 182 447 216
tri 372 166 388 182 ne
rect 388 166 431 182
tri 431 166 447 182 nw
tri 147 129 177 159 sw
tri 253 129 283 159 se
rect 283 136 342 161
tri 342 136 372 166 sw
tri 447 136 477 166 se
rect 477 136 533 301
rect 283 129 533 136
rect 91 125 533 129
rect 91 91 101 125
rect 135 91 295 125
rect 329 91 392 125
rect 426 91 489 125
rect 523 91 533 125
rect 91 75 533 91
rect 593 335 649 351
rect 593 301 603 335
rect 637 301 649 335
rect 593 263 649 301
rect 679 314 841 351
tri 679 298 695 314 ne
rect 695 298 841 314
tri 755 268 785 298 ne
rect 593 229 603 263
rect 637 229 649 263
rect 593 195 649 229
rect 593 161 603 195
rect 637 161 649 195
tri 679 252 695 268 se
rect 695 252 739 268
tri 739 252 755 268 sw
rect 679 219 755 252
rect 679 185 700 219
rect 734 185 755 219
rect 679 183 755 185
tri 679 167 695 183 ne
rect 695 167 739 183
tri 739 167 755 183 nw
rect 785 263 841 298
rect 785 229 797 263
rect 831 229 841 263
rect 785 195 841 229
rect 593 137 649 161
tri 649 137 679 167 sw
tri 755 137 785 167 se
rect 785 161 797 195
rect 831 161 841 195
rect 785 137 841 161
rect 593 125 841 137
rect 593 91 603 125
rect 637 91 700 125
rect 734 91 797 125
rect 831 91 841 125
rect 593 75 841 91
rect 1053 335 1109 351
rect 1053 301 1063 335
rect 1097 301 1109 335
rect 1053 263 1109 301
rect 1139 335 1409 351
rect 1139 306 1160 335
tri 1139 290 1155 306 ne
rect 1155 301 1160 306
rect 1194 301 1257 335
rect 1291 301 1354 335
rect 1388 301 1409 335
rect 1155 290 1409 301
rect 1439 335 1495 351
rect 1439 301 1451 335
rect 1485 301 1495 335
rect 1053 229 1063 263
rect 1097 229 1109 263
tri 1215 260 1245 290 ne
rect 1245 263 1304 290
rect 1053 195 1109 229
rect 1053 161 1063 195
rect 1097 161 1109 195
rect 1053 129 1109 161
tri 1139 244 1155 260 se
rect 1155 244 1199 260
tri 1199 244 1215 260 sw
rect 1139 210 1215 244
rect 1139 176 1160 210
rect 1194 176 1215 210
rect 1139 175 1215 176
tri 1139 159 1155 175 ne
rect 1155 159 1199 175
tri 1199 159 1215 175 nw
rect 1245 229 1257 263
rect 1291 229 1304 263
tri 1304 260 1334 290 nw
rect 1245 195 1304 229
rect 1245 161 1257 195
rect 1291 161 1304 195
tri 1334 244 1350 260 se
rect 1350 244 1393 260
tri 1393 244 1409 260 sw
rect 1334 216 1409 244
rect 1334 182 1355 216
rect 1389 182 1409 216
tri 1334 166 1350 182 ne
rect 1350 166 1393 182
tri 1393 166 1409 182 nw
tri 1109 129 1139 159 sw
tri 1215 129 1245 159 se
rect 1245 136 1304 161
tri 1304 136 1334 166 sw
tri 1409 136 1439 166 se
rect 1439 136 1495 301
rect 1245 129 1495 136
rect 1053 125 1495 129
rect 1053 91 1063 125
rect 1097 91 1257 125
rect 1291 91 1354 125
rect 1388 91 1451 125
rect 1485 91 1495 125
rect 1053 75 1495 91
rect 1555 335 1611 351
rect 1555 301 1565 335
rect 1599 301 1611 335
rect 1555 263 1611 301
rect 1641 314 1803 351
tri 1641 298 1657 314 ne
rect 1657 298 1803 314
tri 1717 268 1747 298 ne
rect 1555 229 1565 263
rect 1599 229 1611 263
rect 1555 195 1611 229
rect 1555 161 1565 195
rect 1599 161 1611 195
tri 1641 252 1657 268 se
rect 1657 252 1701 268
tri 1701 252 1717 268 sw
rect 1641 219 1717 252
rect 1641 185 1662 219
rect 1696 185 1717 219
rect 1641 183 1717 185
tri 1641 167 1657 183 ne
rect 1657 167 1701 183
tri 1701 167 1717 183 nw
rect 1747 263 1803 298
rect 1747 229 1759 263
rect 1793 229 1803 263
rect 1747 195 1803 229
rect 1555 137 1611 161
tri 1611 137 1641 167 sw
tri 1717 137 1747 167 se
rect 1747 161 1759 195
rect 1793 161 1803 195
rect 1747 137 1803 161
rect 1555 125 1803 137
rect 1555 91 1565 125
rect 1599 91 1662 125
rect 1696 91 1759 125
rect 1793 91 1803 125
rect 1555 75 1803 91
rect 2015 335 2071 351
rect 2015 301 2025 335
rect 2059 301 2071 335
rect 2015 263 2071 301
rect 2101 335 2371 351
rect 2101 306 2122 335
tri 2101 290 2117 306 ne
rect 2117 301 2122 306
rect 2156 301 2219 335
rect 2253 301 2316 335
rect 2350 301 2371 335
rect 2117 290 2371 301
rect 2401 335 2457 351
rect 2401 301 2413 335
rect 2447 301 2457 335
rect 2015 229 2025 263
rect 2059 229 2071 263
tri 2177 260 2207 290 ne
rect 2207 263 2266 290
rect 2015 195 2071 229
rect 2015 161 2025 195
rect 2059 161 2071 195
rect 2015 129 2071 161
tri 2101 244 2117 260 se
rect 2117 244 2161 260
tri 2161 244 2177 260 sw
rect 2101 210 2177 244
rect 2101 176 2122 210
rect 2156 176 2177 210
rect 2101 175 2177 176
tri 2101 159 2117 175 ne
rect 2117 159 2161 175
tri 2161 159 2177 175 nw
rect 2207 229 2219 263
rect 2253 229 2266 263
tri 2266 260 2296 290 nw
rect 2207 195 2266 229
rect 2207 161 2219 195
rect 2253 161 2266 195
tri 2296 244 2312 260 se
rect 2312 244 2355 260
tri 2355 244 2371 260 sw
rect 2296 216 2371 244
rect 2296 182 2317 216
rect 2351 182 2371 216
tri 2296 166 2312 182 ne
rect 2312 166 2355 182
tri 2355 166 2371 182 nw
tri 2071 129 2101 159 sw
tri 2177 129 2207 159 se
rect 2207 136 2266 161
tri 2266 136 2296 166 sw
tri 2371 136 2401 166 se
rect 2401 136 2457 301
rect 2207 129 2457 136
rect 2015 125 2457 129
rect 2015 91 2025 125
rect 2059 91 2219 125
rect 2253 91 2316 125
rect 2350 91 2413 125
rect 2447 91 2457 125
rect 2015 75 2457 91
rect 2517 335 2573 351
rect 2517 301 2527 335
rect 2561 301 2573 335
rect 2517 263 2573 301
rect 2603 314 2765 351
tri 2603 298 2619 314 ne
rect 2619 298 2765 314
tri 2679 268 2709 298 ne
rect 2517 229 2527 263
rect 2561 229 2573 263
rect 2517 195 2573 229
rect 2517 161 2527 195
rect 2561 161 2573 195
tri 2603 252 2619 268 se
rect 2619 252 2663 268
tri 2663 252 2679 268 sw
rect 2603 219 2679 252
rect 2603 185 2624 219
rect 2658 185 2679 219
rect 2603 183 2679 185
tri 2603 167 2619 183 ne
rect 2619 167 2663 183
tri 2663 167 2679 183 nw
rect 2709 263 2765 298
rect 2709 229 2721 263
rect 2755 229 2765 263
rect 2709 195 2765 229
rect 2517 137 2573 161
tri 2573 137 2603 167 sw
tri 2679 137 2709 167 se
rect 2709 161 2721 195
rect 2755 161 2765 195
rect 2709 137 2765 161
rect 2517 125 2765 137
rect 2517 91 2527 125
rect 2561 91 2624 125
rect 2658 91 2721 125
rect 2755 91 2765 125
rect 2517 75 2765 91
rect 2977 335 3033 351
rect 2977 301 2987 335
rect 3021 301 3033 335
rect 2977 263 3033 301
rect 3063 335 3333 351
rect 3063 306 3084 335
tri 3063 290 3079 306 ne
rect 3079 301 3084 306
rect 3118 301 3181 335
rect 3215 301 3278 335
rect 3312 301 3333 335
rect 3079 290 3333 301
rect 3363 335 3419 351
rect 3363 301 3375 335
rect 3409 301 3419 335
rect 2977 229 2987 263
rect 3021 229 3033 263
tri 3139 260 3169 290 ne
rect 3169 263 3228 290
rect 2977 195 3033 229
rect 2977 161 2987 195
rect 3021 161 3033 195
rect 2977 129 3033 161
tri 3063 244 3079 260 se
rect 3079 244 3123 260
tri 3123 244 3139 260 sw
rect 3063 210 3139 244
rect 3063 176 3084 210
rect 3118 176 3139 210
rect 3063 175 3139 176
tri 3063 159 3079 175 ne
rect 3079 159 3123 175
tri 3123 159 3139 175 nw
rect 3169 229 3181 263
rect 3215 229 3228 263
tri 3228 260 3258 290 nw
rect 3169 195 3228 229
rect 3169 161 3181 195
rect 3215 161 3228 195
tri 3258 244 3274 260 se
rect 3274 244 3317 260
tri 3317 244 3333 260 sw
rect 3258 216 3333 244
rect 3258 182 3279 216
rect 3313 182 3333 216
tri 3258 166 3274 182 ne
rect 3274 166 3317 182
tri 3317 166 3333 182 nw
tri 3033 129 3063 159 sw
tri 3139 129 3169 159 se
rect 3169 136 3228 161
tri 3228 136 3258 166 sw
tri 3333 136 3363 166 se
rect 3363 136 3419 301
rect 3169 129 3419 136
rect 2977 125 3419 129
rect 2977 91 2987 125
rect 3021 91 3181 125
rect 3215 91 3278 125
rect 3312 91 3375 125
rect 3409 91 3419 125
rect 2977 75 3419 91
rect 3479 335 3535 351
rect 3479 301 3489 335
rect 3523 301 3535 335
rect 3479 263 3535 301
rect 3565 314 3727 351
tri 3565 298 3581 314 ne
rect 3581 298 3727 314
tri 3641 268 3671 298 ne
rect 3479 229 3489 263
rect 3523 229 3535 263
rect 3479 195 3535 229
rect 3479 161 3489 195
rect 3523 161 3535 195
tri 3565 252 3581 268 se
rect 3581 252 3625 268
tri 3625 252 3641 268 sw
rect 3565 219 3641 252
rect 3565 185 3586 219
rect 3620 185 3641 219
rect 3565 183 3641 185
tri 3565 167 3581 183 ne
rect 3581 167 3625 183
tri 3625 167 3641 183 nw
rect 3671 263 3727 298
rect 3671 229 3683 263
rect 3717 229 3727 263
rect 3671 195 3727 229
rect 3479 137 3535 161
tri 3535 137 3565 167 sw
tri 3641 137 3671 167 se
rect 3671 161 3683 195
rect 3717 161 3727 195
rect 3671 137 3727 161
rect 3479 125 3727 137
rect 3479 91 3489 125
rect 3523 91 3586 125
rect 3620 91 3683 125
rect 3717 91 3727 125
rect 3479 75 3727 91
rect 3939 335 3995 351
rect 3939 301 3949 335
rect 3983 301 3995 335
rect 3939 263 3995 301
rect 4025 335 4295 351
rect 4025 306 4046 335
tri 4025 290 4041 306 ne
rect 4041 301 4046 306
rect 4080 301 4143 335
rect 4177 301 4240 335
rect 4274 301 4295 335
rect 4041 290 4295 301
rect 4325 335 4381 351
rect 4325 301 4337 335
rect 4371 301 4381 335
rect 3939 229 3949 263
rect 3983 229 3995 263
tri 4101 260 4131 290 ne
rect 4131 263 4190 290
rect 3939 195 3995 229
rect 3939 161 3949 195
rect 3983 161 3995 195
rect 3939 129 3995 161
tri 4025 244 4041 260 se
rect 4041 244 4085 260
tri 4085 244 4101 260 sw
rect 4025 210 4101 244
rect 4025 176 4046 210
rect 4080 176 4101 210
rect 4025 175 4101 176
tri 4025 159 4041 175 ne
rect 4041 159 4085 175
tri 4085 159 4101 175 nw
rect 4131 229 4143 263
rect 4177 229 4190 263
tri 4190 260 4220 290 nw
rect 4131 195 4190 229
rect 4131 161 4143 195
rect 4177 161 4190 195
tri 4220 244 4236 260 se
rect 4236 244 4279 260
tri 4279 244 4295 260 sw
rect 4220 216 4295 244
rect 4220 182 4241 216
rect 4275 182 4295 216
tri 4220 166 4236 182 ne
rect 4236 166 4279 182
tri 4279 166 4295 182 nw
tri 3995 129 4025 159 sw
tri 4101 129 4131 159 se
rect 4131 136 4190 161
tri 4190 136 4220 166 sw
tri 4295 136 4325 166 se
rect 4325 136 4381 301
rect 4131 129 4381 136
rect 3939 125 4381 129
rect 3939 91 3949 125
rect 3983 91 4143 125
rect 4177 91 4240 125
rect 4274 91 4337 125
rect 4371 91 4381 125
rect 3939 75 4381 91
rect 4441 335 4497 351
rect 4441 301 4451 335
rect 4485 301 4497 335
rect 4441 263 4497 301
rect 4527 314 4689 351
tri 4527 298 4543 314 ne
rect 4543 298 4689 314
tri 4603 268 4633 298 ne
rect 4441 229 4451 263
rect 4485 229 4497 263
rect 4441 195 4497 229
rect 4441 161 4451 195
rect 4485 161 4497 195
tri 4527 252 4543 268 se
rect 4543 252 4587 268
tri 4587 252 4603 268 sw
rect 4527 219 4603 252
rect 4527 185 4548 219
rect 4582 185 4603 219
rect 4527 183 4603 185
tri 4527 167 4543 183 ne
rect 4543 167 4587 183
tri 4587 167 4603 183 nw
rect 4633 263 4689 298
rect 4633 229 4645 263
rect 4679 229 4689 263
rect 4633 195 4689 229
rect 4441 137 4497 161
tri 4497 137 4527 167 sw
tri 4603 137 4633 167 se
rect 4633 161 4645 195
rect 4679 161 4689 195
rect 4633 137 4689 161
rect 4441 125 4689 137
rect 4441 91 4451 125
rect 4485 91 4548 125
rect 4582 91 4645 125
rect 4679 91 4689 125
rect 4441 75 4689 91
rect 4901 335 4957 351
rect 4901 301 4911 335
rect 4945 301 4957 335
rect 4901 263 4957 301
rect 4987 335 5257 351
rect 4987 306 5008 335
tri 4987 290 5003 306 ne
rect 5003 301 5008 306
rect 5042 301 5105 335
rect 5139 301 5202 335
rect 5236 301 5257 335
rect 5003 290 5257 301
rect 5287 335 5343 351
rect 5287 301 5299 335
rect 5333 301 5343 335
rect 4901 229 4911 263
rect 4945 229 4957 263
tri 5063 260 5093 290 ne
rect 5093 263 5152 290
rect 4901 195 4957 229
rect 4901 161 4911 195
rect 4945 161 4957 195
rect 4901 129 4957 161
tri 4987 244 5003 260 se
rect 5003 244 5047 260
tri 5047 244 5063 260 sw
rect 4987 210 5063 244
rect 4987 176 5008 210
rect 5042 176 5063 210
rect 4987 175 5063 176
tri 4987 159 5003 175 ne
rect 5003 159 5047 175
tri 5047 159 5063 175 nw
rect 5093 229 5105 263
rect 5139 229 5152 263
tri 5152 260 5182 290 nw
rect 5093 195 5152 229
rect 5093 161 5105 195
rect 5139 161 5152 195
tri 5182 244 5198 260 se
rect 5198 244 5241 260
tri 5241 244 5257 260 sw
rect 5182 216 5257 244
rect 5182 182 5203 216
rect 5237 182 5257 216
tri 5182 166 5198 182 ne
rect 5198 166 5241 182
tri 5241 166 5257 182 nw
tri 4957 129 4987 159 sw
tri 5063 129 5093 159 se
rect 5093 136 5152 161
tri 5152 136 5182 166 sw
tri 5257 136 5287 166 se
rect 5287 136 5343 301
rect 5093 129 5343 136
rect 4901 125 5343 129
rect 4901 91 4911 125
rect 4945 91 5105 125
rect 5139 91 5202 125
rect 5236 91 5299 125
rect 5333 91 5343 125
rect 4901 75 5343 91
rect 5403 335 5459 351
rect 5403 301 5413 335
rect 5447 301 5459 335
rect 5403 263 5459 301
rect 5489 314 5651 351
tri 5489 298 5505 314 ne
rect 5505 298 5651 314
tri 5565 268 5595 298 ne
rect 5403 229 5413 263
rect 5447 229 5459 263
rect 5403 195 5459 229
rect 5403 161 5413 195
rect 5447 161 5459 195
tri 5489 252 5505 268 se
rect 5505 252 5549 268
tri 5549 252 5565 268 sw
rect 5489 219 5565 252
rect 5489 185 5510 219
rect 5544 185 5565 219
rect 5489 183 5565 185
tri 5489 167 5505 183 ne
rect 5505 167 5549 183
tri 5549 167 5565 183 nw
rect 5595 263 5651 298
rect 5595 229 5607 263
rect 5641 229 5651 263
rect 5595 195 5651 229
rect 5403 137 5459 161
tri 5459 137 5489 167 sw
tri 5565 137 5595 167 se
rect 5595 161 5607 195
rect 5641 161 5651 195
rect 5595 137 5651 161
rect 5403 125 5651 137
rect 5403 91 5413 125
rect 5447 91 5510 125
rect 5544 91 5607 125
rect 5641 91 5651 125
rect 5403 75 5651 91
rect 5863 335 5919 351
rect 5863 301 5873 335
rect 5907 301 5919 335
rect 5863 263 5919 301
rect 5949 335 6219 351
rect 5949 306 5970 335
tri 5949 290 5965 306 ne
rect 5965 301 5970 306
rect 6004 301 6067 335
rect 6101 301 6164 335
rect 6198 301 6219 335
rect 5965 290 6219 301
rect 6249 335 6305 351
rect 6249 301 6261 335
rect 6295 301 6305 335
rect 5863 229 5873 263
rect 5907 229 5919 263
tri 6025 260 6055 290 ne
rect 6055 263 6114 290
rect 5863 195 5919 229
rect 5863 161 5873 195
rect 5907 161 5919 195
rect 5863 129 5919 161
tri 5949 244 5965 260 se
rect 5965 244 6009 260
tri 6009 244 6025 260 sw
rect 5949 210 6025 244
rect 5949 176 5970 210
rect 6004 176 6025 210
rect 5949 175 6025 176
tri 5949 159 5965 175 ne
rect 5965 159 6009 175
tri 6009 159 6025 175 nw
rect 6055 229 6067 263
rect 6101 229 6114 263
tri 6114 260 6144 290 nw
rect 6055 195 6114 229
rect 6055 161 6067 195
rect 6101 161 6114 195
tri 6144 244 6160 260 se
rect 6160 244 6203 260
tri 6203 244 6219 260 sw
rect 6144 216 6219 244
rect 6144 182 6165 216
rect 6199 182 6219 216
tri 6144 166 6160 182 ne
rect 6160 166 6203 182
tri 6203 166 6219 182 nw
tri 5919 129 5949 159 sw
tri 6025 129 6055 159 se
rect 6055 136 6114 161
tri 6114 136 6144 166 sw
tri 6219 136 6249 166 se
rect 6249 136 6305 301
rect 6055 129 6305 136
rect 5863 125 6305 129
rect 5863 91 5873 125
rect 5907 91 6067 125
rect 6101 91 6164 125
rect 6198 91 6261 125
rect 6295 91 6305 125
rect 5863 75 6305 91
rect 6365 335 6421 351
rect 6365 301 6375 335
rect 6409 301 6421 335
rect 6365 263 6421 301
rect 6451 314 6613 351
tri 6451 298 6467 314 ne
rect 6467 298 6613 314
tri 6527 268 6557 298 ne
rect 6365 229 6375 263
rect 6409 229 6421 263
rect 6365 195 6421 229
rect 6365 161 6375 195
rect 6409 161 6421 195
tri 6451 252 6467 268 se
rect 6467 252 6511 268
tri 6511 252 6527 268 sw
rect 6451 219 6527 252
rect 6451 185 6472 219
rect 6506 185 6527 219
rect 6451 183 6527 185
tri 6451 167 6467 183 ne
rect 6467 167 6511 183
tri 6511 167 6527 183 nw
rect 6557 263 6613 298
rect 6557 229 6569 263
rect 6603 229 6613 263
rect 6557 195 6613 229
rect 6365 137 6421 161
tri 6421 137 6451 167 sw
tri 6527 137 6557 167 se
rect 6557 161 6569 195
rect 6603 161 6613 195
rect 6557 137 6613 161
rect 6365 125 6613 137
rect 6365 91 6375 125
rect 6409 91 6472 125
rect 6506 91 6569 125
rect 6603 91 6613 125
rect 6365 75 6613 91
rect 6825 335 6881 351
rect 6825 301 6835 335
rect 6869 301 6881 335
rect 6825 263 6881 301
rect 6911 335 7181 351
rect 6911 306 6932 335
tri 6911 290 6927 306 ne
rect 6927 301 6932 306
rect 6966 301 7029 335
rect 7063 301 7126 335
rect 7160 301 7181 335
rect 6927 290 7181 301
rect 7211 335 7267 351
rect 7211 301 7223 335
rect 7257 301 7267 335
rect 6825 229 6835 263
rect 6869 229 6881 263
tri 6987 260 7017 290 ne
rect 7017 263 7076 290
rect 6825 195 6881 229
rect 6825 161 6835 195
rect 6869 161 6881 195
rect 6825 129 6881 161
tri 6911 244 6927 260 se
rect 6927 244 6971 260
tri 6971 244 6987 260 sw
rect 6911 210 6987 244
rect 6911 176 6932 210
rect 6966 176 6987 210
rect 6911 175 6987 176
tri 6911 159 6927 175 ne
rect 6927 159 6971 175
tri 6971 159 6987 175 nw
rect 7017 229 7029 263
rect 7063 229 7076 263
tri 7076 260 7106 290 nw
rect 7017 195 7076 229
rect 7017 161 7029 195
rect 7063 161 7076 195
tri 7106 244 7122 260 se
rect 7122 244 7165 260
tri 7165 244 7181 260 sw
rect 7106 216 7181 244
rect 7106 182 7127 216
rect 7161 182 7181 216
tri 7106 166 7122 182 ne
rect 7122 166 7165 182
tri 7165 166 7181 182 nw
tri 6881 129 6911 159 sw
tri 6987 129 7017 159 se
rect 7017 136 7076 161
tri 7076 136 7106 166 sw
tri 7181 136 7211 166 se
rect 7211 136 7267 301
rect 7017 129 7267 136
rect 6825 125 7267 129
rect 6825 91 6835 125
rect 6869 91 7029 125
rect 7063 91 7126 125
rect 7160 91 7223 125
rect 7257 91 7267 125
rect 6825 75 7267 91
rect 7327 335 7383 351
rect 7327 301 7337 335
rect 7371 301 7383 335
rect 7327 263 7383 301
rect 7413 314 7575 351
tri 7413 298 7429 314 ne
rect 7429 298 7575 314
tri 7489 268 7519 298 ne
rect 7327 229 7337 263
rect 7371 229 7383 263
rect 7327 195 7383 229
rect 7327 161 7337 195
rect 7371 161 7383 195
tri 7413 252 7429 268 se
rect 7429 252 7473 268
tri 7473 252 7489 268 sw
rect 7413 219 7489 252
rect 7413 185 7434 219
rect 7468 185 7489 219
rect 7413 183 7489 185
tri 7413 167 7429 183 ne
rect 7429 167 7473 183
tri 7473 167 7489 183 nw
rect 7519 263 7575 298
rect 7519 229 7531 263
rect 7565 229 7575 263
rect 7519 195 7575 229
rect 7327 137 7383 161
tri 7383 137 7413 167 sw
tri 7489 137 7519 167 se
rect 7519 161 7531 195
rect 7565 161 7575 195
rect 7519 137 7575 161
rect 7327 125 7575 137
rect 7327 91 7337 125
rect 7371 91 7434 125
rect 7468 91 7531 125
rect 7565 91 7575 125
rect 7327 75 7575 91
rect 7787 335 7843 351
rect 7787 301 7797 335
rect 7831 301 7843 335
rect 7787 263 7843 301
rect 7873 335 8143 351
rect 7873 306 7894 335
tri 7873 290 7889 306 ne
rect 7889 301 7894 306
rect 7928 301 7991 335
rect 8025 301 8088 335
rect 8122 301 8143 335
rect 7889 290 8143 301
rect 8173 335 8229 351
rect 8173 301 8185 335
rect 8219 301 8229 335
rect 7787 229 7797 263
rect 7831 229 7843 263
tri 7949 260 7979 290 ne
rect 7979 263 8038 290
rect 7787 195 7843 229
rect 7787 161 7797 195
rect 7831 161 7843 195
rect 7787 129 7843 161
tri 7873 244 7889 260 se
rect 7889 244 7933 260
tri 7933 244 7949 260 sw
rect 7873 210 7949 244
rect 7873 176 7894 210
rect 7928 176 7949 210
rect 7873 175 7949 176
tri 7873 159 7889 175 ne
rect 7889 159 7933 175
tri 7933 159 7949 175 nw
rect 7979 229 7991 263
rect 8025 229 8038 263
tri 8038 260 8068 290 nw
rect 7979 195 8038 229
rect 7979 161 7991 195
rect 8025 161 8038 195
tri 8068 244 8084 260 se
rect 8084 244 8127 260
tri 8127 244 8143 260 sw
rect 8068 216 8143 244
rect 8068 182 8089 216
rect 8123 182 8143 216
tri 8068 166 8084 182 ne
rect 8084 166 8127 182
tri 8127 166 8143 182 nw
tri 7843 129 7873 159 sw
tri 7949 129 7979 159 se
rect 7979 136 8038 161
tri 8038 136 8068 166 sw
tri 8143 136 8173 166 se
rect 8173 136 8229 301
rect 7979 129 8229 136
rect 7787 125 8229 129
rect 7787 91 7797 125
rect 7831 91 7991 125
rect 8025 91 8088 125
rect 8122 91 8185 125
rect 8219 91 8229 125
rect 7787 75 8229 91
rect 8289 335 8345 351
rect 8289 301 8299 335
rect 8333 301 8345 335
rect 8289 263 8345 301
rect 8375 314 8537 351
tri 8375 298 8391 314 ne
rect 8391 298 8537 314
tri 8451 268 8481 298 ne
rect 8289 229 8299 263
rect 8333 229 8345 263
rect 8289 195 8345 229
rect 8289 161 8299 195
rect 8333 161 8345 195
tri 8375 252 8391 268 se
rect 8391 252 8435 268
tri 8435 252 8451 268 sw
rect 8375 219 8451 252
rect 8375 185 8396 219
rect 8430 185 8451 219
rect 8375 183 8451 185
tri 8375 167 8391 183 ne
rect 8391 167 8435 183
tri 8435 167 8451 183 nw
rect 8481 263 8537 298
rect 8481 229 8493 263
rect 8527 229 8537 263
rect 8481 195 8537 229
rect 8289 137 8345 161
tri 8345 137 8375 167 sw
tri 8451 137 8481 167 se
rect 8481 161 8493 195
rect 8527 161 8537 195
rect 8481 137 8537 161
rect 8289 125 8537 137
rect 8289 91 8299 125
rect 8333 91 8396 125
rect 8430 91 8493 125
rect 8527 91 8537 125
rect 8289 75 8537 91
rect 8749 335 8805 351
rect 8749 301 8759 335
rect 8793 301 8805 335
rect 8749 263 8805 301
rect 8835 335 9105 351
rect 8835 306 8856 335
tri 8835 290 8851 306 ne
rect 8851 301 8856 306
rect 8890 301 8953 335
rect 8987 301 9050 335
rect 9084 301 9105 335
rect 8851 290 9105 301
rect 9135 335 9191 351
rect 9135 301 9147 335
rect 9181 301 9191 335
rect 8749 229 8759 263
rect 8793 229 8805 263
tri 8911 260 8941 290 ne
rect 8941 263 9000 290
rect 8749 195 8805 229
rect 8749 161 8759 195
rect 8793 161 8805 195
rect 8749 129 8805 161
tri 8835 244 8851 260 se
rect 8851 244 8895 260
tri 8895 244 8911 260 sw
rect 8835 210 8911 244
rect 8835 176 8856 210
rect 8890 176 8911 210
rect 8835 175 8911 176
tri 8835 159 8851 175 ne
rect 8851 159 8895 175
tri 8895 159 8911 175 nw
rect 8941 229 8953 263
rect 8987 229 9000 263
tri 9000 260 9030 290 nw
rect 8941 195 9000 229
rect 8941 161 8953 195
rect 8987 161 9000 195
tri 9030 244 9046 260 se
rect 9046 244 9089 260
tri 9089 244 9105 260 sw
rect 9030 216 9105 244
rect 9030 182 9051 216
rect 9085 182 9105 216
tri 9030 166 9046 182 ne
rect 9046 166 9089 182
tri 9089 166 9105 182 nw
tri 8805 129 8835 159 sw
tri 8911 129 8941 159 se
rect 8941 136 9000 161
tri 9000 136 9030 166 sw
tri 9105 136 9135 166 se
rect 9135 136 9191 301
rect 8941 129 9191 136
rect 8749 125 9191 129
rect 8749 91 8759 125
rect 8793 91 8953 125
rect 8987 91 9050 125
rect 9084 91 9147 125
rect 9181 91 9191 125
rect 8749 75 9191 91
rect 9251 335 9307 351
rect 9251 301 9261 335
rect 9295 301 9307 335
rect 9251 263 9307 301
rect 9337 314 9499 351
tri 9337 298 9353 314 ne
rect 9353 298 9499 314
tri 9413 268 9443 298 ne
rect 9251 229 9261 263
rect 9295 229 9307 263
rect 9251 195 9307 229
rect 9251 161 9261 195
rect 9295 161 9307 195
tri 9337 252 9353 268 se
rect 9353 252 9397 268
tri 9397 252 9413 268 sw
rect 9337 219 9413 252
rect 9337 185 9358 219
rect 9392 185 9413 219
rect 9337 183 9413 185
tri 9337 167 9353 183 ne
rect 9353 167 9397 183
tri 9397 167 9413 183 nw
rect 9443 263 9499 298
rect 9443 229 9455 263
rect 9489 229 9499 263
rect 9443 195 9499 229
rect 9251 137 9307 161
tri 9307 137 9337 167 sw
tri 9413 137 9443 167 se
rect 9443 161 9455 195
rect 9489 161 9499 195
rect 9443 137 9499 161
rect 9251 125 9499 137
rect 9251 91 9261 125
rect 9295 91 9358 125
rect 9392 91 9455 125
rect 9489 91 9499 125
rect 9251 75 9499 91
rect 9711 335 9767 351
rect 9711 301 9721 335
rect 9755 301 9767 335
rect 9711 263 9767 301
rect 9797 335 10067 351
rect 9797 306 9818 335
tri 9797 290 9813 306 ne
rect 9813 301 9818 306
rect 9852 301 9915 335
rect 9949 301 10012 335
rect 10046 301 10067 335
rect 9813 290 10067 301
rect 10097 335 10153 351
rect 10097 301 10109 335
rect 10143 301 10153 335
rect 9711 229 9721 263
rect 9755 229 9767 263
tri 9873 260 9903 290 ne
rect 9903 263 9962 290
rect 9711 195 9767 229
rect 9711 161 9721 195
rect 9755 161 9767 195
rect 9711 129 9767 161
tri 9797 244 9813 260 se
rect 9813 244 9857 260
tri 9857 244 9873 260 sw
rect 9797 210 9873 244
rect 9797 176 9818 210
rect 9852 176 9873 210
rect 9797 175 9873 176
tri 9797 159 9813 175 ne
rect 9813 159 9857 175
tri 9857 159 9873 175 nw
rect 9903 229 9915 263
rect 9949 229 9962 263
tri 9962 260 9992 290 nw
rect 9903 195 9962 229
rect 9903 161 9915 195
rect 9949 161 9962 195
tri 9992 244 10008 260 se
rect 10008 244 10051 260
tri 10051 244 10067 260 sw
rect 9992 216 10067 244
rect 9992 182 10013 216
rect 10047 182 10067 216
tri 9992 166 10008 182 ne
rect 10008 166 10051 182
tri 10051 166 10067 182 nw
tri 9767 129 9797 159 sw
tri 9873 129 9903 159 se
rect 9903 136 9962 161
tri 9962 136 9992 166 sw
tri 10067 136 10097 166 se
rect 10097 136 10153 301
rect 9903 129 10153 136
rect 9711 125 10153 129
rect 9711 91 9721 125
rect 9755 91 9915 125
rect 9949 91 10012 125
rect 10046 91 10109 125
rect 10143 91 10153 125
rect 9711 75 10153 91
rect 10213 335 10269 351
rect 10213 301 10223 335
rect 10257 301 10269 335
rect 10213 263 10269 301
rect 10299 314 10461 351
tri 10299 298 10315 314 ne
rect 10315 298 10461 314
tri 10375 268 10405 298 ne
rect 10213 229 10223 263
rect 10257 229 10269 263
rect 10213 195 10269 229
rect 10213 161 10223 195
rect 10257 161 10269 195
tri 10299 252 10315 268 se
rect 10315 252 10359 268
tri 10359 252 10375 268 sw
rect 10299 219 10375 252
rect 10299 185 10320 219
rect 10354 185 10375 219
rect 10299 183 10375 185
tri 10299 167 10315 183 ne
rect 10315 167 10359 183
tri 10359 167 10375 183 nw
rect 10405 263 10461 298
rect 10405 229 10417 263
rect 10451 229 10461 263
rect 10405 195 10461 229
rect 10213 137 10269 161
tri 10269 137 10299 167 sw
tri 10375 137 10405 167 se
rect 10405 161 10417 195
rect 10451 161 10461 195
rect 10405 137 10461 161
rect 10213 125 10461 137
rect 10213 91 10223 125
rect 10257 91 10320 125
rect 10354 91 10417 125
rect 10451 91 10461 125
rect 10213 75 10461 91
rect 10673 335 10729 351
rect 10673 301 10683 335
rect 10717 301 10729 335
rect 10673 263 10729 301
rect 10759 335 11029 351
rect 10759 306 10780 335
tri 10759 290 10775 306 ne
rect 10775 301 10780 306
rect 10814 301 10877 335
rect 10911 301 10974 335
rect 11008 301 11029 335
rect 10775 290 11029 301
rect 11059 335 11115 351
rect 11059 301 11071 335
rect 11105 301 11115 335
rect 10673 229 10683 263
rect 10717 229 10729 263
tri 10835 260 10865 290 ne
rect 10865 263 10924 290
rect 10673 195 10729 229
rect 10673 161 10683 195
rect 10717 161 10729 195
rect 10673 129 10729 161
tri 10759 244 10775 260 se
rect 10775 244 10819 260
tri 10819 244 10835 260 sw
rect 10759 210 10835 244
rect 10759 176 10780 210
rect 10814 176 10835 210
rect 10759 175 10835 176
tri 10759 159 10775 175 ne
rect 10775 159 10819 175
tri 10819 159 10835 175 nw
rect 10865 229 10877 263
rect 10911 229 10924 263
tri 10924 260 10954 290 nw
rect 10865 195 10924 229
rect 10865 161 10877 195
rect 10911 161 10924 195
tri 10954 244 10970 260 se
rect 10970 244 11013 260
tri 11013 244 11029 260 sw
rect 10954 216 11029 244
rect 10954 182 10975 216
rect 11009 182 11029 216
tri 10954 166 10970 182 ne
rect 10970 166 11013 182
tri 11013 166 11029 182 nw
tri 10729 129 10759 159 sw
tri 10835 129 10865 159 se
rect 10865 136 10924 161
tri 10924 136 10954 166 sw
tri 11029 136 11059 166 se
rect 11059 136 11115 301
rect 10865 129 11115 136
rect 10673 125 11115 129
rect 10673 91 10683 125
rect 10717 91 10877 125
rect 10911 91 10974 125
rect 11008 91 11071 125
rect 11105 91 11115 125
rect 10673 75 11115 91
rect 11175 335 11231 351
rect 11175 301 11185 335
rect 11219 301 11231 335
rect 11175 263 11231 301
rect 11261 314 11423 351
tri 11261 298 11277 314 ne
rect 11277 298 11423 314
tri 11337 268 11367 298 ne
rect 11175 229 11185 263
rect 11219 229 11231 263
rect 11175 195 11231 229
rect 11175 161 11185 195
rect 11219 161 11231 195
tri 11261 252 11277 268 se
rect 11277 252 11321 268
tri 11321 252 11337 268 sw
rect 11261 219 11337 252
rect 11261 185 11282 219
rect 11316 185 11337 219
rect 11261 183 11337 185
tri 11261 167 11277 183 ne
rect 11277 167 11321 183
tri 11321 167 11337 183 nw
rect 11367 263 11423 298
rect 11367 229 11379 263
rect 11413 229 11423 263
rect 11367 195 11423 229
rect 11175 137 11231 161
tri 11231 137 11261 167 sw
tri 11337 137 11367 167 se
rect 11367 161 11379 195
rect 11413 161 11423 195
rect 11367 137 11423 161
rect 11175 125 11423 137
rect 11175 91 11185 125
rect 11219 91 11282 125
rect 11316 91 11379 125
rect 11413 91 11423 125
rect 11175 75 11423 91
rect 11635 335 11691 351
rect 11635 301 11645 335
rect 11679 301 11691 335
rect 11635 263 11691 301
rect 11721 335 11991 351
rect 11721 306 11742 335
tri 11721 290 11737 306 ne
rect 11737 301 11742 306
rect 11776 301 11839 335
rect 11873 301 11936 335
rect 11970 301 11991 335
rect 11737 290 11991 301
rect 12021 335 12077 351
rect 12021 301 12033 335
rect 12067 301 12077 335
rect 11635 229 11645 263
rect 11679 229 11691 263
tri 11797 260 11827 290 ne
rect 11827 263 11886 290
rect 11635 195 11691 229
rect 11635 161 11645 195
rect 11679 161 11691 195
rect 11635 129 11691 161
tri 11721 244 11737 260 se
rect 11737 244 11781 260
tri 11781 244 11797 260 sw
rect 11721 210 11797 244
rect 11721 176 11742 210
rect 11776 176 11797 210
rect 11721 175 11797 176
tri 11721 159 11737 175 ne
rect 11737 159 11781 175
tri 11781 159 11797 175 nw
rect 11827 229 11839 263
rect 11873 229 11886 263
tri 11886 260 11916 290 nw
rect 11827 195 11886 229
rect 11827 161 11839 195
rect 11873 161 11886 195
tri 11916 244 11932 260 se
rect 11932 244 11975 260
tri 11975 244 11991 260 sw
rect 11916 216 11991 244
rect 11916 182 11937 216
rect 11971 182 11991 216
tri 11916 166 11932 182 ne
rect 11932 166 11975 182
tri 11975 166 11991 182 nw
tri 11691 129 11721 159 sw
tri 11797 129 11827 159 se
rect 11827 136 11886 161
tri 11886 136 11916 166 sw
tri 11991 136 12021 166 se
rect 12021 136 12077 301
rect 11827 129 12077 136
rect 11635 125 12077 129
rect 11635 91 11645 125
rect 11679 91 11839 125
rect 11873 91 11936 125
rect 11970 91 12033 125
rect 12067 91 12077 125
rect 11635 75 12077 91
rect 12137 335 12193 351
rect 12137 301 12147 335
rect 12181 301 12193 335
rect 12137 263 12193 301
rect 12223 314 12385 351
tri 12223 298 12239 314 ne
rect 12239 298 12385 314
tri 12299 268 12329 298 ne
rect 12137 229 12147 263
rect 12181 229 12193 263
rect 12137 195 12193 229
rect 12137 161 12147 195
rect 12181 161 12193 195
tri 12223 252 12239 268 se
rect 12239 252 12283 268
tri 12283 252 12299 268 sw
rect 12223 219 12299 252
rect 12223 185 12244 219
rect 12278 185 12299 219
rect 12223 183 12299 185
tri 12223 167 12239 183 ne
rect 12239 167 12283 183
tri 12283 167 12299 183 nw
rect 12329 263 12385 298
rect 12329 229 12341 263
rect 12375 229 12385 263
rect 12329 195 12385 229
rect 12137 137 12193 161
tri 12193 137 12223 167 sw
tri 12299 137 12329 167 se
rect 12329 161 12341 195
rect 12375 161 12385 195
rect 12329 137 12385 161
rect 12137 125 12385 137
rect 12137 91 12147 125
rect 12181 91 12244 125
rect 12278 91 12341 125
rect 12375 91 12385 125
rect 12137 75 12385 91
rect 12597 335 12653 351
rect 12597 301 12607 335
rect 12641 301 12653 335
rect 12597 263 12653 301
rect 12683 335 12953 351
rect 12683 306 12704 335
tri 12683 290 12699 306 ne
rect 12699 301 12704 306
rect 12738 301 12801 335
rect 12835 301 12898 335
rect 12932 301 12953 335
rect 12699 290 12953 301
rect 12983 335 13039 351
rect 12983 301 12995 335
rect 13029 301 13039 335
rect 12597 229 12607 263
rect 12641 229 12653 263
tri 12759 260 12789 290 ne
rect 12789 263 12848 290
rect 12597 195 12653 229
rect 12597 161 12607 195
rect 12641 161 12653 195
rect 12597 129 12653 161
tri 12683 244 12699 260 se
rect 12699 244 12743 260
tri 12743 244 12759 260 sw
rect 12683 210 12759 244
rect 12683 176 12704 210
rect 12738 176 12759 210
rect 12683 175 12759 176
tri 12683 159 12699 175 ne
rect 12699 159 12743 175
tri 12743 159 12759 175 nw
rect 12789 229 12801 263
rect 12835 229 12848 263
tri 12848 260 12878 290 nw
rect 12789 195 12848 229
rect 12789 161 12801 195
rect 12835 161 12848 195
tri 12878 244 12894 260 se
rect 12894 244 12937 260
tri 12937 244 12953 260 sw
rect 12878 216 12953 244
rect 12878 182 12899 216
rect 12933 182 12953 216
tri 12878 166 12894 182 ne
rect 12894 166 12937 182
tri 12937 166 12953 182 nw
tri 12653 129 12683 159 sw
tri 12759 129 12789 159 se
rect 12789 136 12848 161
tri 12848 136 12878 166 sw
tri 12953 136 12983 166 se
rect 12983 136 13039 301
rect 12789 129 13039 136
rect 12597 125 13039 129
rect 12597 91 12607 125
rect 12641 91 12801 125
rect 12835 91 12898 125
rect 12932 91 12995 125
rect 13029 91 13039 125
rect 12597 75 13039 91
rect 13099 335 13155 351
rect 13099 301 13109 335
rect 13143 301 13155 335
rect 13099 263 13155 301
rect 13185 314 13347 351
tri 13185 298 13201 314 ne
rect 13201 298 13347 314
tri 13261 268 13291 298 ne
rect 13099 229 13109 263
rect 13143 229 13155 263
rect 13099 195 13155 229
rect 13099 161 13109 195
rect 13143 161 13155 195
tri 13185 252 13201 268 se
rect 13201 252 13245 268
tri 13245 252 13261 268 sw
rect 13185 219 13261 252
rect 13185 185 13206 219
rect 13240 185 13261 219
rect 13185 183 13261 185
tri 13185 167 13201 183 ne
rect 13201 167 13245 183
tri 13245 167 13261 183 nw
rect 13291 263 13347 298
rect 13291 229 13303 263
rect 13337 229 13347 263
rect 13291 195 13347 229
rect 13099 137 13155 161
tri 13155 137 13185 167 sw
tri 13261 137 13291 167 se
rect 13291 161 13303 195
rect 13337 161 13347 195
rect 13291 137 13347 161
rect 13099 125 13347 137
rect 13099 91 13109 125
rect 13143 91 13206 125
rect 13240 91 13303 125
rect 13337 91 13347 125
rect 13099 75 13347 91
rect 13559 335 13615 351
rect 13559 301 13569 335
rect 13603 301 13615 335
rect 13559 263 13615 301
rect 13645 335 13915 351
rect 13645 306 13666 335
tri 13645 290 13661 306 ne
rect 13661 301 13666 306
rect 13700 301 13763 335
rect 13797 301 13860 335
rect 13894 301 13915 335
rect 13661 290 13915 301
rect 13945 335 14001 351
rect 13945 301 13957 335
rect 13991 301 14001 335
rect 13559 229 13569 263
rect 13603 229 13615 263
tri 13721 260 13751 290 ne
rect 13751 263 13810 290
rect 13559 195 13615 229
rect 13559 161 13569 195
rect 13603 161 13615 195
rect 13559 129 13615 161
tri 13645 244 13661 260 se
rect 13661 244 13705 260
tri 13705 244 13721 260 sw
rect 13645 210 13721 244
rect 13645 176 13666 210
rect 13700 176 13721 210
rect 13645 175 13721 176
tri 13645 159 13661 175 ne
rect 13661 159 13705 175
tri 13705 159 13721 175 nw
rect 13751 229 13763 263
rect 13797 229 13810 263
tri 13810 260 13840 290 nw
rect 13751 195 13810 229
rect 13751 161 13763 195
rect 13797 161 13810 195
tri 13840 244 13856 260 se
rect 13856 244 13899 260
tri 13899 244 13915 260 sw
rect 13840 216 13915 244
rect 13840 182 13861 216
rect 13895 182 13915 216
tri 13840 166 13856 182 ne
rect 13856 166 13899 182
tri 13899 166 13915 182 nw
tri 13615 129 13645 159 sw
tri 13721 129 13751 159 se
rect 13751 136 13810 161
tri 13810 136 13840 166 sw
tri 13915 136 13945 166 se
rect 13945 136 14001 301
rect 13751 129 14001 136
rect 13559 125 14001 129
rect 13559 91 13569 125
rect 13603 91 13763 125
rect 13797 91 13860 125
rect 13894 91 13957 125
rect 13991 91 14001 125
rect 13559 75 14001 91
rect 14061 335 14117 351
rect 14061 301 14071 335
rect 14105 301 14117 335
rect 14061 263 14117 301
rect 14147 314 14309 351
tri 14147 298 14163 314 ne
rect 14163 298 14309 314
tri 14223 268 14253 298 ne
rect 14061 229 14071 263
rect 14105 229 14117 263
rect 14061 195 14117 229
rect 14061 161 14071 195
rect 14105 161 14117 195
tri 14147 252 14163 268 se
rect 14163 252 14207 268
tri 14207 252 14223 268 sw
rect 14147 219 14223 252
rect 14147 185 14168 219
rect 14202 185 14223 219
rect 14147 183 14223 185
tri 14147 167 14163 183 ne
rect 14163 167 14207 183
tri 14207 167 14223 183 nw
rect 14253 263 14309 298
rect 14253 229 14265 263
rect 14299 229 14309 263
rect 14253 195 14309 229
rect 14061 137 14117 161
tri 14117 137 14147 167 sw
tri 14223 137 14253 167 se
rect 14253 161 14265 195
rect 14299 161 14309 195
rect 14253 137 14309 161
rect 14061 125 14309 137
rect 14061 91 14071 125
rect 14105 91 14168 125
rect 14202 91 14265 125
rect 14299 91 14309 125
rect 14061 75 14309 91
rect 14521 335 14577 351
rect 14521 301 14531 335
rect 14565 301 14577 335
rect 14521 263 14577 301
rect 14607 335 14877 351
rect 14607 306 14628 335
tri 14607 290 14623 306 ne
rect 14623 301 14628 306
rect 14662 301 14725 335
rect 14759 301 14822 335
rect 14856 301 14877 335
rect 14623 290 14877 301
rect 14907 335 14963 351
rect 14907 301 14919 335
rect 14953 301 14963 335
rect 14521 229 14531 263
rect 14565 229 14577 263
tri 14683 260 14713 290 ne
rect 14713 263 14772 290
rect 14521 195 14577 229
rect 14521 161 14531 195
rect 14565 161 14577 195
rect 14521 129 14577 161
tri 14607 244 14623 260 se
rect 14623 244 14667 260
tri 14667 244 14683 260 sw
rect 14607 210 14683 244
rect 14607 176 14628 210
rect 14662 176 14683 210
rect 14607 175 14683 176
tri 14607 159 14623 175 ne
rect 14623 159 14667 175
tri 14667 159 14683 175 nw
rect 14713 229 14725 263
rect 14759 229 14772 263
tri 14772 260 14802 290 nw
rect 14713 195 14772 229
rect 14713 161 14725 195
rect 14759 161 14772 195
tri 14802 244 14818 260 se
rect 14818 244 14861 260
tri 14861 244 14877 260 sw
rect 14802 216 14877 244
rect 14802 182 14823 216
rect 14857 182 14877 216
tri 14802 166 14818 182 ne
rect 14818 166 14861 182
tri 14861 166 14877 182 nw
tri 14577 129 14607 159 sw
tri 14683 129 14713 159 se
rect 14713 136 14772 161
tri 14772 136 14802 166 sw
tri 14877 136 14907 166 se
rect 14907 136 14963 301
rect 14713 129 14963 136
rect 14521 125 14963 129
rect 14521 91 14531 125
rect 14565 91 14725 125
rect 14759 91 14822 125
rect 14856 91 14919 125
rect 14953 91 14963 125
rect 14521 75 14963 91
rect 15023 335 15079 351
rect 15023 301 15033 335
rect 15067 301 15079 335
rect 15023 263 15079 301
rect 15109 314 15271 351
tri 15109 298 15125 314 ne
rect 15125 298 15271 314
tri 15185 268 15215 298 ne
rect 15023 229 15033 263
rect 15067 229 15079 263
rect 15023 195 15079 229
rect 15023 161 15033 195
rect 15067 161 15079 195
tri 15109 252 15125 268 se
rect 15125 252 15169 268
tri 15169 252 15185 268 sw
rect 15109 219 15185 252
rect 15109 185 15130 219
rect 15164 185 15185 219
rect 15109 183 15185 185
tri 15109 167 15125 183 ne
rect 15125 167 15169 183
tri 15169 167 15185 183 nw
rect 15215 263 15271 298
rect 15215 229 15227 263
rect 15261 229 15271 263
rect 15215 195 15271 229
rect 15023 137 15079 161
tri 15079 137 15109 167 sw
tri 15185 137 15215 167 se
rect 15215 161 15227 195
rect 15261 161 15271 195
rect 15215 137 15271 161
rect 15023 125 15271 137
rect 15023 91 15033 125
rect 15067 91 15130 125
rect 15164 91 15227 125
rect 15261 91 15271 125
rect 15023 75 15271 91
rect 15483 335 15539 351
rect 15483 301 15493 335
rect 15527 301 15539 335
rect 15483 263 15539 301
rect 15569 335 15839 351
rect 15569 306 15590 335
tri 15569 290 15585 306 ne
rect 15585 301 15590 306
rect 15624 301 15687 335
rect 15721 301 15784 335
rect 15818 301 15839 335
rect 15585 290 15839 301
rect 15869 335 15925 351
rect 15869 301 15881 335
rect 15915 301 15925 335
rect 15483 229 15493 263
rect 15527 229 15539 263
tri 15645 260 15675 290 ne
rect 15675 263 15734 290
rect 15483 195 15539 229
rect 15483 161 15493 195
rect 15527 161 15539 195
rect 15483 129 15539 161
tri 15569 244 15585 260 se
rect 15585 244 15629 260
tri 15629 244 15645 260 sw
rect 15569 210 15645 244
rect 15569 176 15590 210
rect 15624 176 15645 210
rect 15569 175 15645 176
tri 15569 159 15585 175 ne
rect 15585 159 15629 175
tri 15629 159 15645 175 nw
rect 15675 229 15687 263
rect 15721 229 15734 263
tri 15734 260 15764 290 nw
rect 15675 195 15734 229
rect 15675 161 15687 195
rect 15721 161 15734 195
tri 15764 244 15780 260 se
rect 15780 244 15823 260
tri 15823 244 15839 260 sw
rect 15764 216 15839 244
rect 15764 182 15785 216
rect 15819 182 15839 216
tri 15764 166 15780 182 ne
rect 15780 166 15823 182
tri 15823 166 15839 182 nw
tri 15539 129 15569 159 sw
tri 15645 129 15675 159 se
rect 15675 136 15734 161
tri 15734 136 15764 166 sw
tri 15839 136 15869 166 se
rect 15869 136 15925 301
rect 15675 129 15925 136
rect 15483 125 15925 129
rect 15483 91 15493 125
rect 15527 91 15687 125
rect 15721 91 15784 125
rect 15818 91 15881 125
rect 15915 91 15925 125
rect 15483 75 15925 91
rect 15985 335 16041 351
rect 15985 301 15995 335
rect 16029 301 16041 335
rect 15985 263 16041 301
rect 16071 314 16233 351
tri 16071 298 16087 314 ne
rect 16087 298 16233 314
tri 16147 268 16177 298 ne
rect 15985 229 15995 263
rect 16029 229 16041 263
rect 15985 195 16041 229
rect 15985 161 15995 195
rect 16029 161 16041 195
tri 16071 252 16087 268 se
rect 16087 252 16131 268
tri 16131 252 16147 268 sw
rect 16071 219 16147 252
rect 16071 185 16092 219
rect 16126 185 16147 219
rect 16071 183 16147 185
tri 16071 167 16087 183 ne
rect 16087 167 16131 183
tri 16131 167 16147 183 nw
rect 16177 263 16233 298
rect 16177 229 16189 263
rect 16223 229 16233 263
rect 16177 195 16233 229
rect 15985 137 16041 161
tri 16041 137 16071 167 sw
tri 16147 137 16177 167 se
rect 16177 161 16189 195
rect 16223 161 16233 195
rect 16177 137 16233 161
rect 15985 125 16233 137
rect 15985 91 15995 125
rect 16029 91 16092 125
rect 16126 91 16189 125
rect 16223 91 16233 125
rect 15985 75 16233 91
rect 16445 335 16501 351
rect 16445 301 16455 335
rect 16489 301 16501 335
rect 16445 263 16501 301
rect 16531 335 16801 351
rect 16531 306 16552 335
tri 16531 290 16547 306 ne
rect 16547 301 16552 306
rect 16586 301 16649 335
rect 16683 301 16746 335
rect 16780 301 16801 335
rect 16547 290 16801 301
rect 16831 335 16887 351
rect 16831 301 16843 335
rect 16877 301 16887 335
rect 16445 229 16455 263
rect 16489 229 16501 263
tri 16607 260 16637 290 ne
rect 16637 263 16696 290
rect 16445 195 16501 229
rect 16445 161 16455 195
rect 16489 161 16501 195
rect 16445 129 16501 161
tri 16531 244 16547 260 se
rect 16547 244 16591 260
tri 16591 244 16607 260 sw
rect 16531 210 16607 244
rect 16531 176 16552 210
rect 16586 176 16607 210
rect 16531 175 16607 176
tri 16531 159 16547 175 ne
rect 16547 159 16591 175
tri 16591 159 16607 175 nw
rect 16637 229 16649 263
rect 16683 229 16696 263
tri 16696 260 16726 290 nw
rect 16637 195 16696 229
rect 16637 161 16649 195
rect 16683 161 16696 195
tri 16726 244 16742 260 se
rect 16742 244 16785 260
tri 16785 244 16801 260 sw
rect 16726 216 16801 244
rect 16726 182 16747 216
rect 16781 182 16801 216
tri 16726 166 16742 182 ne
rect 16742 166 16785 182
tri 16785 166 16801 182 nw
tri 16501 129 16531 159 sw
tri 16607 129 16637 159 se
rect 16637 136 16696 161
tri 16696 136 16726 166 sw
tri 16801 136 16831 166 se
rect 16831 136 16887 301
rect 16637 129 16887 136
rect 16445 125 16887 129
rect 16445 91 16455 125
rect 16489 91 16649 125
rect 16683 91 16746 125
rect 16780 91 16843 125
rect 16877 91 16887 125
rect 16445 75 16887 91
rect 16947 335 17003 351
rect 16947 301 16957 335
rect 16991 301 17003 335
rect 16947 263 17003 301
rect 17033 314 17195 351
tri 17033 298 17049 314 ne
rect 17049 298 17195 314
tri 17109 268 17139 298 ne
rect 16947 229 16957 263
rect 16991 229 17003 263
rect 16947 195 17003 229
rect 16947 161 16957 195
rect 16991 161 17003 195
tri 17033 252 17049 268 se
rect 17049 252 17093 268
tri 17093 252 17109 268 sw
rect 17033 219 17109 252
rect 17033 185 17054 219
rect 17088 185 17109 219
rect 17033 183 17109 185
tri 17033 167 17049 183 ne
rect 17049 167 17093 183
tri 17093 167 17109 183 nw
rect 17139 263 17195 298
rect 17139 229 17151 263
rect 17185 229 17195 263
rect 17139 195 17195 229
rect 16947 137 17003 161
tri 17003 137 17033 167 sw
tri 17109 137 17139 167 se
rect 17139 161 17151 195
rect 17185 161 17195 195
rect 17139 137 17195 161
rect 16947 125 17195 137
rect 16947 91 16957 125
rect 16991 91 17054 125
rect 17088 91 17151 125
rect 17185 91 17195 125
rect 16947 75 17195 91
rect 17428 333 17484 349
rect 17428 299 17438 333
rect 17472 299 17484 333
rect 17428 261 17484 299
rect 17514 333 17678 349
rect 17514 304 17535 333
tri 17514 288 17530 304 ne
rect 17530 299 17535 304
rect 17569 299 17632 333
rect 17666 299 17678 333
rect 17530 288 17678 299
rect 17708 333 17868 349
rect 17708 312 17826 333
tri 17708 296 17724 312 ne
rect 17724 299 17826 312
rect 17860 299 17868 333
rect 17724 296 17868 299
rect 17428 227 17438 261
rect 17472 227 17484 261
tri 17590 258 17620 288 ne
rect 17620 261 17678 288
tri 17784 266 17814 296 ne
rect 17428 193 17484 227
rect 17428 159 17438 193
rect 17472 159 17484 193
rect 17428 127 17484 159
tri 17514 242 17530 258 se
rect 17530 242 17574 258
tri 17574 242 17590 258 sw
rect 17514 208 17590 242
rect 17514 174 17535 208
rect 17569 174 17590 208
rect 17514 173 17590 174
tri 17514 157 17530 173 ne
rect 17530 157 17574 173
tri 17574 157 17590 173 nw
rect 17620 227 17632 261
rect 17666 227 17678 261
rect 17620 193 17678 227
rect 17620 159 17632 193
rect 17666 159 17678 193
tri 17708 250 17724 266 se
rect 17724 250 17768 266
tri 17768 250 17784 266 sw
rect 17708 217 17784 250
rect 17708 183 17728 217
rect 17762 183 17784 217
rect 17708 181 17784 183
tri 17708 165 17724 181 ne
rect 17724 165 17768 181
tri 17768 165 17784 181 nw
rect 17814 261 17868 296
rect 17814 227 17826 261
rect 17860 227 17868 261
rect 17814 193 17868 227
tri 17484 127 17514 157 sw
tri 17590 127 17620 157 se
rect 17620 135 17678 159
tri 17678 135 17708 165 sw
tri 17784 135 17814 165 se
rect 17814 159 17826 193
rect 17860 159 17868 193
rect 17814 135 17868 159
rect 17620 127 17868 135
rect 17428 123 17868 127
rect 17428 89 17438 123
rect 17472 89 17632 123
rect 17666 89 17728 123
rect 17762 89 17826 123
rect 17860 89 17868 123
rect 17428 73 17868 89
rect 18094 333 18150 349
rect 18094 299 18104 333
rect 18138 299 18150 333
rect 18094 261 18150 299
rect 18180 333 18450 349
rect 18180 304 18201 333
tri 18180 288 18196 304 ne
rect 18196 299 18201 304
rect 18235 299 18298 333
rect 18332 312 18450 333
rect 18332 299 18434 312
rect 18196 296 18434 299
tri 18434 296 18450 312 nw
rect 18480 333 18536 349
rect 18480 299 18492 333
rect 18526 299 18536 333
rect 18196 288 18344 296
rect 18094 227 18104 261
rect 18138 227 18150 261
tri 18256 258 18286 288 ne
rect 18286 261 18344 288
tri 18344 266 18374 296 nw
rect 18094 193 18150 227
rect 18094 159 18104 193
rect 18138 159 18150 193
rect 18094 127 18150 159
tri 18180 242 18196 258 se
rect 18196 242 18240 258
tri 18240 242 18256 258 sw
rect 18180 208 18256 242
rect 18180 174 18201 208
rect 18235 174 18256 208
rect 18180 173 18256 174
tri 18180 157 18196 173 ne
rect 18196 157 18240 173
tri 18240 157 18256 173 nw
rect 18286 227 18298 261
rect 18332 227 18344 261
rect 18286 193 18344 227
rect 18286 159 18298 193
rect 18332 159 18344 193
tri 18374 250 18390 266 se
rect 18390 250 18434 266
tri 18434 250 18450 266 sw
rect 18374 217 18450 250
rect 18374 183 18395 217
rect 18429 183 18450 217
rect 18374 181 18450 183
tri 18374 165 18390 181 ne
rect 18390 165 18434 181
tri 18434 165 18450 181 nw
rect 18480 261 18536 299
rect 18480 227 18492 261
rect 18526 227 18536 261
rect 18480 193 18536 227
tri 18150 127 18180 157 sw
tri 18256 127 18286 157 se
rect 18286 135 18344 159
tri 18344 135 18374 165 sw
tri 18450 135 18480 165 se
rect 18480 159 18492 193
rect 18526 159 18536 193
rect 18480 135 18536 159
rect 18286 127 18536 135
rect 18094 123 18536 127
rect 18094 89 18104 123
rect 18138 89 18298 123
rect 18332 89 18395 123
rect 18429 89 18492 123
rect 18526 89 18536 123
rect 18094 73 18536 89
rect 18760 333 18816 349
rect 18760 299 18770 333
rect 18804 299 18816 333
rect 18760 261 18816 299
rect 18846 333 19010 349
rect 18846 304 18867 333
tri 18846 288 18862 304 ne
rect 18862 299 18867 304
rect 18901 299 18964 333
rect 18998 299 19010 333
rect 18862 288 19010 299
rect 19040 312 19202 349
tri 19040 296 19056 312 ne
rect 19056 296 19202 312
rect 18760 227 18770 261
rect 18804 227 18816 261
tri 18922 258 18952 288 ne
rect 18952 261 19010 288
tri 19116 266 19146 296 ne
rect 18760 193 18816 227
rect 18760 159 18770 193
rect 18804 159 18816 193
rect 18760 127 18816 159
tri 18846 242 18862 258 se
rect 18862 242 18906 258
tri 18906 242 18922 258 sw
rect 18846 208 18922 242
rect 18846 174 18867 208
rect 18901 174 18922 208
rect 18846 173 18922 174
tri 18846 157 18862 173 ne
rect 18862 157 18906 173
tri 18906 157 18922 173 nw
rect 18952 227 18964 261
rect 18998 227 19010 261
tri 19041 251 19056 266 se
rect 19056 251 19100 266
tri 19100 251 19115 266 sw
rect 19146 261 19202 296
rect 18952 193 19010 227
rect 18952 159 18964 193
rect 18998 159 19010 193
rect 19040 217 19116 251
rect 19040 183 19061 217
rect 19095 183 19116 217
rect 19040 181 19116 183
tri 19040 165 19056 181 ne
rect 19056 165 19100 181
tri 19100 165 19116 181 nw
rect 19146 227 19158 261
rect 19192 227 19202 261
rect 19146 193 19202 227
tri 18816 127 18846 157 sw
tri 18922 127 18952 157 se
rect 18952 135 19010 159
tri 19010 135 19040 165 sw
tri 19116 135 19146 165 se
rect 19146 159 19158 193
rect 19192 159 19202 193
rect 19146 135 19202 159
rect 18952 127 19202 135
rect 18760 123 19202 127
rect 18760 89 18770 123
rect 18804 89 18964 123
rect 18998 89 19061 123
rect 19095 89 19158 123
rect 19192 89 19202 123
rect 18760 73 19202 89
<< pdiff >>
rect 191 1366 247 1404
rect 191 1332 201 1366
rect 235 1332 247 1366
rect 191 1298 247 1332
rect 191 1264 201 1298
rect 235 1264 247 1298
rect 191 1230 247 1264
rect 191 1196 201 1230
rect 235 1196 247 1230
rect 191 1162 247 1196
rect 191 1128 201 1162
rect 235 1128 247 1162
rect 191 1093 247 1128
rect 191 1059 201 1093
rect 235 1059 247 1093
rect 191 1004 247 1059
rect 277 1366 335 1404
rect 277 1332 289 1366
rect 323 1332 335 1366
rect 277 1298 335 1332
rect 277 1264 289 1298
rect 323 1264 335 1298
rect 277 1230 335 1264
rect 277 1196 289 1230
rect 323 1196 335 1230
rect 277 1162 335 1196
rect 277 1128 289 1162
rect 323 1128 335 1162
rect 277 1093 335 1128
rect 277 1059 289 1093
rect 323 1059 335 1093
rect 277 1004 335 1059
rect 365 1366 423 1404
rect 365 1332 377 1366
rect 411 1332 423 1366
rect 365 1298 423 1332
rect 365 1264 377 1298
rect 411 1264 423 1298
rect 365 1230 423 1264
rect 365 1196 377 1230
rect 411 1196 423 1230
rect 365 1162 423 1196
rect 365 1128 377 1162
rect 411 1128 423 1162
rect 365 1004 423 1128
rect 453 1366 511 1404
rect 453 1332 465 1366
rect 499 1332 511 1366
rect 453 1298 511 1332
rect 453 1264 465 1298
rect 499 1264 511 1298
rect 453 1230 511 1264
rect 453 1196 465 1230
rect 499 1196 511 1230
rect 453 1162 511 1196
rect 453 1128 465 1162
rect 499 1128 511 1162
rect 453 1093 511 1128
rect 453 1059 465 1093
rect 499 1059 511 1093
rect 453 1004 511 1059
rect 541 1366 599 1404
rect 541 1332 553 1366
rect 587 1332 599 1366
rect 541 1298 599 1332
rect 541 1264 553 1298
rect 587 1264 599 1298
rect 541 1230 599 1264
rect 541 1196 553 1230
rect 587 1196 599 1230
rect 541 1162 599 1196
rect 541 1128 553 1162
rect 587 1128 599 1162
rect 541 1004 599 1128
rect 629 1366 687 1404
rect 629 1332 641 1366
rect 675 1332 687 1366
rect 629 1298 687 1332
rect 629 1264 641 1298
rect 675 1264 687 1298
rect 629 1230 687 1264
rect 629 1196 641 1230
rect 675 1196 687 1230
rect 629 1162 687 1196
rect 629 1128 641 1162
rect 675 1128 687 1162
rect 629 1093 687 1128
rect 629 1059 641 1093
rect 675 1059 687 1093
rect 629 1004 687 1059
rect 717 1366 771 1404
rect 717 1332 729 1366
rect 763 1332 771 1366
rect 717 1298 771 1332
rect 717 1264 729 1298
rect 763 1264 771 1298
rect 717 1230 771 1264
rect 717 1196 729 1230
rect 763 1196 771 1230
rect 717 1162 771 1196
rect 717 1128 729 1162
rect 763 1128 771 1162
rect 717 1004 771 1128
rect 1153 1366 1209 1404
rect 1153 1332 1163 1366
rect 1197 1332 1209 1366
rect 1153 1298 1209 1332
rect 1153 1264 1163 1298
rect 1197 1264 1209 1298
rect 1153 1230 1209 1264
rect 1153 1196 1163 1230
rect 1197 1196 1209 1230
rect 1153 1162 1209 1196
rect 1153 1128 1163 1162
rect 1197 1128 1209 1162
rect 1153 1093 1209 1128
rect 1153 1059 1163 1093
rect 1197 1059 1209 1093
rect 1153 1004 1209 1059
rect 1239 1366 1297 1404
rect 1239 1332 1251 1366
rect 1285 1332 1297 1366
rect 1239 1298 1297 1332
rect 1239 1264 1251 1298
rect 1285 1264 1297 1298
rect 1239 1230 1297 1264
rect 1239 1196 1251 1230
rect 1285 1196 1297 1230
rect 1239 1162 1297 1196
rect 1239 1128 1251 1162
rect 1285 1128 1297 1162
rect 1239 1093 1297 1128
rect 1239 1059 1251 1093
rect 1285 1059 1297 1093
rect 1239 1004 1297 1059
rect 1327 1366 1385 1404
rect 1327 1332 1339 1366
rect 1373 1332 1385 1366
rect 1327 1298 1385 1332
rect 1327 1264 1339 1298
rect 1373 1264 1385 1298
rect 1327 1230 1385 1264
rect 1327 1196 1339 1230
rect 1373 1196 1385 1230
rect 1327 1162 1385 1196
rect 1327 1128 1339 1162
rect 1373 1128 1385 1162
rect 1327 1004 1385 1128
rect 1415 1366 1473 1404
rect 1415 1332 1427 1366
rect 1461 1332 1473 1366
rect 1415 1298 1473 1332
rect 1415 1264 1427 1298
rect 1461 1264 1473 1298
rect 1415 1230 1473 1264
rect 1415 1196 1427 1230
rect 1461 1196 1473 1230
rect 1415 1162 1473 1196
rect 1415 1128 1427 1162
rect 1461 1128 1473 1162
rect 1415 1093 1473 1128
rect 1415 1059 1427 1093
rect 1461 1059 1473 1093
rect 1415 1004 1473 1059
rect 1503 1366 1561 1404
rect 1503 1332 1515 1366
rect 1549 1332 1561 1366
rect 1503 1298 1561 1332
rect 1503 1264 1515 1298
rect 1549 1264 1561 1298
rect 1503 1230 1561 1264
rect 1503 1196 1515 1230
rect 1549 1196 1561 1230
rect 1503 1162 1561 1196
rect 1503 1128 1515 1162
rect 1549 1128 1561 1162
rect 1503 1004 1561 1128
rect 1591 1366 1649 1404
rect 1591 1332 1603 1366
rect 1637 1332 1649 1366
rect 1591 1298 1649 1332
rect 1591 1264 1603 1298
rect 1637 1264 1649 1298
rect 1591 1230 1649 1264
rect 1591 1196 1603 1230
rect 1637 1196 1649 1230
rect 1591 1162 1649 1196
rect 1591 1128 1603 1162
rect 1637 1128 1649 1162
rect 1591 1093 1649 1128
rect 1591 1059 1603 1093
rect 1637 1059 1649 1093
rect 1591 1004 1649 1059
rect 1679 1366 1733 1404
rect 1679 1332 1691 1366
rect 1725 1332 1733 1366
rect 1679 1298 1733 1332
rect 1679 1264 1691 1298
rect 1725 1264 1733 1298
rect 1679 1230 1733 1264
rect 1679 1196 1691 1230
rect 1725 1196 1733 1230
rect 1679 1162 1733 1196
rect 1679 1128 1691 1162
rect 1725 1128 1733 1162
rect 1679 1004 1733 1128
rect 2115 1366 2171 1404
rect 2115 1332 2125 1366
rect 2159 1332 2171 1366
rect 2115 1298 2171 1332
rect 2115 1264 2125 1298
rect 2159 1264 2171 1298
rect 2115 1230 2171 1264
rect 2115 1196 2125 1230
rect 2159 1196 2171 1230
rect 2115 1162 2171 1196
rect 2115 1128 2125 1162
rect 2159 1128 2171 1162
rect 2115 1093 2171 1128
rect 2115 1059 2125 1093
rect 2159 1059 2171 1093
rect 2115 1004 2171 1059
rect 2201 1366 2259 1404
rect 2201 1332 2213 1366
rect 2247 1332 2259 1366
rect 2201 1298 2259 1332
rect 2201 1264 2213 1298
rect 2247 1264 2259 1298
rect 2201 1230 2259 1264
rect 2201 1196 2213 1230
rect 2247 1196 2259 1230
rect 2201 1162 2259 1196
rect 2201 1128 2213 1162
rect 2247 1128 2259 1162
rect 2201 1093 2259 1128
rect 2201 1059 2213 1093
rect 2247 1059 2259 1093
rect 2201 1004 2259 1059
rect 2289 1366 2347 1404
rect 2289 1332 2301 1366
rect 2335 1332 2347 1366
rect 2289 1298 2347 1332
rect 2289 1264 2301 1298
rect 2335 1264 2347 1298
rect 2289 1230 2347 1264
rect 2289 1196 2301 1230
rect 2335 1196 2347 1230
rect 2289 1162 2347 1196
rect 2289 1128 2301 1162
rect 2335 1128 2347 1162
rect 2289 1004 2347 1128
rect 2377 1366 2435 1404
rect 2377 1332 2389 1366
rect 2423 1332 2435 1366
rect 2377 1298 2435 1332
rect 2377 1264 2389 1298
rect 2423 1264 2435 1298
rect 2377 1230 2435 1264
rect 2377 1196 2389 1230
rect 2423 1196 2435 1230
rect 2377 1162 2435 1196
rect 2377 1128 2389 1162
rect 2423 1128 2435 1162
rect 2377 1093 2435 1128
rect 2377 1059 2389 1093
rect 2423 1059 2435 1093
rect 2377 1004 2435 1059
rect 2465 1366 2523 1404
rect 2465 1332 2477 1366
rect 2511 1332 2523 1366
rect 2465 1298 2523 1332
rect 2465 1264 2477 1298
rect 2511 1264 2523 1298
rect 2465 1230 2523 1264
rect 2465 1196 2477 1230
rect 2511 1196 2523 1230
rect 2465 1162 2523 1196
rect 2465 1128 2477 1162
rect 2511 1128 2523 1162
rect 2465 1004 2523 1128
rect 2553 1366 2611 1404
rect 2553 1332 2565 1366
rect 2599 1332 2611 1366
rect 2553 1298 2611 1332
rect 2553 1264 2565 1298
rect 2599 1264 2611 1298
rect 2553 1230 2611 1264
rect 2553 1196 2565 1230
rect 2599 1196 2611 1230
rect 2553 1162 2611 1196
rect 2553 1128 2565 1162
rect 2599 1128 2611 1162
rect 2553 1093 2611 1128
rect 2553 1059 2565 1093
rect 2599 1059 2611 1093
rect 2553 1004 2611 1059
rect 2641 1366 2695 1404
rect 2641 1332 2653 1366
rect 2687 1332 2695 1366
rect 2641 1298 2695 1332
rect 2641 1264 2653 1298
rect 2687 1264 2695 1298
rect 2641 1230 2695 1264
rect 2641 1196 2653 1230
rect 2687 1196 2695 1230
rect 2641 1162 2695 1196
rect 2641 1128 2653 1162
rect 2687 1128 2695 1162
rect 2641 1004 2695 1128
rect 3077 1366 3133 1404
rect 3077 1332 3087 1366
rect 3121 1332 3133 1366
rect 3077 1298 3133 1332
rect 3077 1264 3087 1298
rect 3121 1264 3133 1298
rect 3077 1230 3133 1264
rect 3077 1196 3087 1230
rect 3121 1196 3133 1230
rect 3077 1162 3133 1196
rect 3077 1128 3087 1162
rect 3121 1128 3133 1162
rect 3077 1093 3133 1128
rect 3077 1059 3087 1093
rect 3121 1059 3133 1093
rect 3077 1004 3133 1059
rect 3163 1366 3221 1404
rect 3163 1332 3175 1366
rect 3209 1332 3221 1366
rect 3163 1298 3221 1332
rect 3163 1264 3175 1298
rect 3209 1264 3221 1298
rect 3163 1230 3221 1264
rect 3163 1196 3175 1230
rect 3209 1196 3221 1230
rect 3163 1162 3221 1196
rect 3163 1128 3175 1162
rect 3209 1128 3221 1162
rect 3163 1093 3221 1128
rect 3163 1059 3175 1093
rect 3209 1059 3221 1093
rect 3163 1004 3221 1059
rect 3251 1366 3309 1404
rect 3251 1332 3263 1366
rect 3297 1332 3309 1366
rect 3251 1298 3309 1332
rect 3251 1264 3263 1298
rect 3297 1264 3309 1298
rect 3251 1230 3309 1264
rect 3251 1196 3263 1230
rect 3297 1196 3309 1230
rect 3251 1162 3309 1196
rect 3251 1128 3263 1162
rect 3297 1128 3309 1162
rect 3251 1004 3309 1128
rect 3339 1366 3397 1404
rect 3339 1332 3351 1366
rect 3385 1332 3397 1366
rect 3339 1298 3397 1332
rect 3339 1264 3351 1298
rect 3385 1264 3397 1298
rect 3339 1230 3397 1264
rect 3339 1196 3351 1230
rect 3385 1196 3397 1230
rect 3339 1162 3397 1196
rect 3339 1128 3351 1162
rect 3385 1128 3397 1162
rect 3339 1093 3397 1128
rect 3339 1059 3351 1093
rect 3385 1059 3397 1093
rect 3339 1004 3397 1059
rect 3427 1366 3485 1404
rect 3427 1332 3439 1366
rect 3473 1332 3485 1366
rect 3427 1298 3485 1332
rect 3427 1264 3439 1298
rect 3473 1264 3485 1298
rect 3427 1230 3485 1264
rect 3427 1196 3439 1230
rect 3473 1196 3485 1230
rect 3427 1162 3485 1196
rect 3427 1128 3439 1162
rect 3473 1128 3485 1162
rect 3427 1004 3485 1128
rect 3515 1366 3573 1404
rect 3515 1332 3527 1366
rect 3561 1332 3573 1366
rect 3515 1298 3573 1332
rect 3515 1264 3527 1298
rect 3561 1264 3573 1298
rect 3515 1230 3573 1264
rect 3515 1196 3527 1230
rect 3561 1196 3573 1230
rect 3515 1162 3573 1196
rect 3515 1128 3527 1162
rect 3561 1128 3573 1162
rect 3515 1093 3573 1128
rect 3515 1059 3527 1093
rect 3561 1059 3573 1093
rect 3515 1004 3573 1059
rect 3603 1366 3657 1404
rect 3603 1332 3615 1366
rect 3649 1332 3657 1366
rect 3603 1298 3657 1332
rect 3603 1264 3615 1298
rect 3649 1264 3657 1298
rect 3603 1230 3657 1264
rect 3603 1196 3615 1230
rect 3649 1196 3657 1230
rect 3603 1162 3657 1196
rect 3603 1128 3615 1162
rect 3649 1128 3657 1162
rect 3603 1004 3657 1128
rect 4039 1366 4095 1404
rect 4039 1332 4049 1366
rect 4083 1332 4095 1366
rect 4039 1298 4095 1332
rect 4039 1264 4049 1298
rect 4083 1264 4095 1298
rect 4039 1230 4095 1264
rect 4039 1196 4049 1230
rect 4083 1196 4095 1230
rect 4039 1162 4095 1196
rect 4039 1128 4049 1162
rect 4083 1128 4095 1162
rect 4039 1093 4095 1128
rect 4039 1059 4049 1093
rect 4083 1059 4095 1093
rect 4039 1004 4095 1059
rect 4125 1366 4183 1404
rect 4125 1332 4137 1366
rect 4171 1332 4183 1366
rect 4125 1298 4183 1332
rect 4125 1264 4137 1298
rect 4171 1264 4183 1298
rect 4125 1230 4183 1264
rect 4125 1196 4137 1230
rect 4171 1196 4183 1230
rect 4125 1162 4183 1196
rect 4125 1128 4137 1162
rect 4171 1128 4183 1162
rect 4125 1093 4183 1128
rect 4125 1059 4137 1093
rect 4171 1059 4183 1093
rect 4125 1004 4183 1059
rect 4213 1366 4271 1404
rect 4213 1332 4225 1366
rect 4259 1332 4271 1366
rect 4213 1298 4271 1332
rect 4213 1264 4225 1298
rect 4259 1264 4271 1298
rect 4213 1230 4271 1264
rect 4213 1196 4225 1230
rect 4259 1196 4271 1230
rect 4213 1162 4271 1196
rect 4213 1128 4225 1162
rect 4259 1128 4271 1162
rect 4213 1004 4271 1128
rect 4301 1366 4359 1404
rect 4301 1332 4313 1366
rect 4347 1332 4359 1366
rect 4301 1298 4359 1332
rect 4301 1264 4313 1298
rect 4347 1264 4359 1298
rect 4301 1230 4359 1264
rect 4301 1196 4313 1230
rect 4347 1196 4359 1230
rect 4301 1162 4359 1196
rect 4301 1128 4313 1162
rect 4347 1128 4359 1162
rect 4301 1093 4359 1128
rect 4301 1059 4313 1093
rect 4347 1059 4359 1093
rect 4301 1004 4359 1059
rect 4389 1366 4447 1404
rect 4389 1332 4401 1366
rect 4435 1332 4447 1366
rect 4389 1298 4447 1332
rect 4389 1264 4401 1298
rect 4435 1264 4447 1298
rect 4389 1230 4447 1264
rect 4389 1196 4401 1230
rect 4435 1196 4447 1230
rect 4389 1162 4447 1196
rect 4389 1128 4401 1162
rect 4435 1128 4447 1162
rect 4389 1004 4447 1128
rect 4477 1366 4535 1404
rect 4477 1332 4489 1366
rect 4523 1332 4535 1366
rect 4477 1298 4535 1332
rect 4477 1264 4489 1298
rect 4523 1264 4535 1298
rect 4477 1230 4535 1264
rect 4477 1196 4489 1230
rect 4523 1196 4535 1230
rect 4477 1162 4535 1196
rect 4477 1128 4489 1162
rect 4523 1128 4535 1162
rect 4477 1093 4535 1128
rect 4477 1059 4489 1093
rect 4523 1059 4535 1093
rect 4477 1004 4535 1059
rect 4565 1366 4619 1404
rect 4565 1332 4577 1366
rect 4611 1332 4619 1366
rect 4565 1298 4619 1332
rect 4565 1264 4577 1298
rect 4611 1264 4619 1298
rect 4565 1230 4619 1264
rect 4565 1196 4577 1230
rect 4611 1196 4619 1230
rect 4565 1162 4619 1196
rect 4565 1128 4577 1162
rect 4611 1128 4619 1162
rect 4565 1004 4619 1128
rect 5001 1366 5057 1404
rect 5001 1332 5011 1366
rect 5045 1332 5057 1366
rect 5001 1298 5057 1332
rect 5001 1264 5011 1298
rect 5045 1264 5057 1298
rect 5001 1230 5057 1264
rect 5001 1196 5011 1230
rect 5045 1196 5057 1230
rect 5001 1162 5057 1196
rect 5001 1128 5011 1162
rect 5045 1128 5057 1162
rect 5001 1093 5057 1128
rect 5001 1059 5011 1093
rect 5045 1059 5057 1093
rect 5001 1004 5057 1059
rect 5087 1366 5145 1404
rect 5087 1332 5099 1366
rect 5133 1332 5145 1366
rect 5087 1298 5145 1332
rect 5087 1264 5099 1298
rect 5133 1264 5145 1298
rect 5087 1230 5145 1264
rect 5087 1196 5099 1230
rect 5133 1196 5145 1230
rect 5087 1162 5145 1196
rect 5087 1128 5099 1162
rect 5133 1128 5145 1162
rect 5087 1093 5145 1128
rect 5087 1059 5099 1093
rect 5133 1059 5145 1093
rect 5087 1004 5145 1059
rect 5175 1366 5233 1404
rect 5175 1332 5187 1366
rect 5221 1332 5233 1366
rect 5175 1298 5233 1332
rect 5175 1264 5187 1298
rect 5221 1264 5233 1298
rect 5175 1230 5233 1264
rect 5175 1196 5187 1230
rect 5221 1196 5233 1230
rect 5175 1162 5233 1196
rect 5175 1128 5187 1162
rect 5221 1128 5233 1162
rect 5175 1004 5233 1128
rect 5263 1366 5321 1404
rect 5263 1332 5275 1366
rect 5309 1332 5321 1366
rect 5263 1298 5321 1332
rect 5263 1264 5275 1298
rect 5309 1264 5321 1298
rect 5263 1230 5321 1264
rect 5263 1196 5275 1230
rect 5309 1196 5321 1230
rect 5263 1162 5321 1196
rect 5263 1128 5275 1162
rect 5309 1128 5321 1162
rect 5263 1093 5321 1128
rect 5263 1059 5275 1093
rect 5309 1059 5321 1093
rect 5263 1004 5321 1059
rect 5351 1366 5409 1404
rect 5351 1332 5363 1366
rect 5397 1332 5409 1366
rect 5351 1298 5409 1332
rect 5351 1264 5363 1298
rect 5397 1264 5409 1298
rect 5351 1230 5409 1264
rect 5351 1196 5363 1230
rect 5397 1196 5409 1230
rect 5351 1162 5409 1196
rect 5351 1128 5363 1162
rect 5397 1128 5409 1162
rect 5351 1004 5409 1128
rect 5439 1366 5497 1404
rect 5439 1332 5451 1366
rect 5485 1332 5497 1366
rect 5439 1298 5497 1332
rect 5439 1264 5451 1298
rect 5485 1264 5497 1298
rect 5439 1230 5497 1264
rect 5439 1196 5451 1230
rect 5485 1196 5497 1230
rect 5439 1162 5497 1196
rect 5439 1128 5451 1162
rect 5485 1128 5497 1162
rect 5439 1093 5497 1128
rect 5439 1059 5451 1093
rect 5485 1059 5497 1093
rect 5439 1004 5497 1059
rect 5527 1366 5581 1404
rect 5527 1332 5539 1366
rect 5573 1332 5581 1366
rect 5527 1298 5581 1332
rect 5527 1264 5539 1298
rect 5573 1264 5581 1298
rect 5527 1230 5581 1264
rect 5527 1196 5539 1230
rect 5573 1196 5581 1230
rect 5527 1162 5581 1196
rect 5527 1128 5539 1162
rect 5573 1128 5581 1162
rect 5527 1004 5581 1128
rect 5963 1366 6019 1404
rect 5963 1332 5973 1366
rect 6007 1332 6019 1366
rect 5963 1298 6019 1332
rect 5963 1264 5973 1298
rect 6007 1264 6019 1298
rect 5963 1230 6019 1264
rect 5963 1196 5973 1230
rect 6007 1196 6019 1230
rect 5963 1162 6019 1196
rect 5963 1128 5973 1162
rect 6007 1128 6019 1162
rect 5963 1093 6019 1128
rect 5963 1059 5973 1093
rect 6007 1059 6019 1093
rect 5963 1004 6019 1059
rect 6049 1366 6107 1404
rect 6049 1332 6061 1366
rect 6095 1332 6107 1366
rect 6049 1298 6107 1332
rect 6049 1264 6061 1298
rect 6095 1264 6107 1298
rect 6049 1230 6107 1264
rect 6049 1196 6061 1230
rect 6095 1196 6107 1230
rect 6049 1162 6107 1196
rect 6049 1128 6061 1162
rect 6095 1128 6107 1162
rect 6049 1093 6107 1128
rect 6049 1059 6061 1093
rect 6095 1059 6107 1093
rect 6049 1004 6107 1059
rect 6137 1366 6195 1404
rect 6137 1332 6149 1366
rect 6183 1332 6195 1366
rect 6137 1298 6195 1332
rect 6137 1264 6149 1298
rect 6183 1264 6195 1298
rect 6137 1230 6195 1264
rect 6137 1196 6149 1230
rect 6183 1196 6195 1230
rect 6137 1162 6195 1196
rect 6137 1128 6149 1162
rect 6183 1128 6195 1162
rect 6137 1004 6195 1128
rect 6225 1366 6283 1404
rect 6225 1332 6237 1366
rect 6271 1332 6283 1366
rect 6225 1298 6283 1332
rect 6225 1264 6237 1298
rect 6271 1264 6283 1298
rect 6225 1230 6283 1264
rect 6225 1196 6237 1230
rect 6271 1196 6283 1230
rect 6225 1162 6283 1196
rect 6225 1128 6237 1162
rect 6271 1128 6283 1162
rect 6225 1093 6283 1128
rect 6225 1059 6237 1093
rect 6271 1059 6283 1093
rect 6225 1004 6283 1059
rect 6313 1366 6371 1404
rect 6313 1332 6325 1366
rect 6359 1332 6371 1366
rect 6313 1298 6371 1332
rect 6313 1264 6325 1298
rect 6359 1264 6371 1298
rect 6313 1230 6371 1264
rect 6313 1196 6325 1230
rect 6359 1196 6371 1230
rect 6313 1162 6371 1196
rect 6313 1128 6325 1162
rect 6359 1128 6371 1162
rect 6313 1004 6371 1128
rect 6401 1366 6459 1404
rect 6401 1332 6413 1366
rect 6447 1332 6459 1366
rect 6401 1298 6459 1332
rect 6401 1264 6413 1298
rect 6447 1264 6459 1298
rect 6401 1230 6459 1264
rect 6401 1196 6413 1230
rect 6447 1196 6459 1230
rect 6401 1162 6459 1196
rect 6401 1128 6413 1162
rect 6447 1128 6459 1162
rect 6401 1093 6459 1128
rect 6401 1059 6413 1093
rect 6447 1059 6459 1093
rect 6401 1004 6459 1059
rect 6489 1366 6543 1404
rect 6489 1332 6501 1366
rect 6535 1332 6543 1366
rect 6489 1298 6543 1332
rect 6489 1264 6501 1298
rect 6535 1264 6543 1298
rect 6489 1230 6543 1264
rect 6489 1196 6501 1230
rect 6535 1196 6543 1230
rect 6489 1162 6543 1196
rect 6489 1128 6501 1162
rect 6535 1128 6543 1162
rect 6489 1004 6543 1128
rect 6925 1366 6981 1404
rect 6925 1332 6935 1366
rect 6969 1332 6981 1366
rect 6925 1298 6981 1332
rect 6925 1264 6935 1298
rect 6969 1264 6981 1298
rect 6925 1230 6981 1264
rect 6925 1196 6935 1230
rect 6969 1196 6981 1230
rect 6925 1162 6981 1196
rect 6925 1128 6935 1162
rect 6969 1128 6981 1162
rect 6925 1093 6981 1128
rect 6925 1059 6935 1093
rect 6969 1059 6981 1093
rect 6925 1004 6981 1059
rect 7011 1366 7069 1404
rect 7011 1332 7023 1366
rect 7057 1332 7069 1366
rect 7011 1298 7069 1332
rect 7011 1264 7023 1298
rect 7057 1264 7069 1298
rect 7011 1230 7069 1264
rect 7011 1196 7023 1230
rect 7057 1196 7069 1230
rect 7011 1162 7069 1196
rect 7011 1128 7023 1162
rect 7057 1128 7069 1162
rect 7011 1093 7069 1128
rect 7011 1059 7023 1093
rect 7057 1059 7069 1093
rect 7011 1004 7069 1059
rect 7099 1366 7157 1404
rect 7099 1332 7111 1366
rect 7145 1332 7157 1366
rect 7099 1298 7157 1332
rect 7099 1264 7111 1298
rect 7145 1264 7157 1298
rect 7099 1230 7157 1264
rect 7099 1196 7111 1230
rect 7145 1196 7157 1230
rect 7099 1162 7157 1196
rect 7099 1128 7111 1162
rect 7145 1128 7157 1162
rect 7099 1004 7157 1128
rect 7187 1366 7245 1404
rect 7187 1332 7199 1366
rect 7233 1332 7245 1366
rect 7187 1298 7245 1332
rect 7187 1264 7199 1298
rect 7233 1264 7245 1298
rect 7187 1230 7245 1264
rect 7187 1196 7199 1230
rect 7233 1196 7245 1230
rect 7187 1162 7245 1196
rect 7187 1128 7199 1162
rect 7233 1128 7245 1162
rect 7187 1093 7245 1128
rect 7187 1059 7199 1093
rect 7233 1059 7245 1093
rect 7187 1004 7245 1059
rect 7275 1366 7333 1404
rect 7275 1332 7287 1366
rect 7321 1332 7333 1366
rect 7275 1298 7333 1332
rect 7275 1264 7287 1298
rect 7321 1264 7333 1298
rect 7275 1230 7333 1264
rect 7275 1196 7287 1230
rect 7321 1196 7333 1230
rect 7275 1162 7333 1196
rect 7275 1128 7287 1162
rect 7321 1128 7333 1162
rect 7275 1004 7333 1128
rect 7363 1366 7421 1404
rect 7363 1332 7375 1366
rect 7409 1332 7421 1366
rect 7363 1298 7421 1332
rect 7363 1264 7375 1298
rect 7409 1264 7421 1298
rect 7363 1230 7421 1264
rect 7363 1196 7375 1230
rect 7409 1196 7421 1230
rect 7363 1162 7421 1196
rect 7363 1128 7375 1162
rect 7409 1128 7421 1162
rect 7363 1093 7421 1128
rect 7363 1059 7375 1093
rect 7409 1059 7421 1093
rect 7363 1004 7421 1059
rect 7451 1366 7505 1404
rect 7451 1332 7463 1366
rect 7497 1332 7505 1366
rect 7451 1298 7505 1332
rect 7451 1264 7463 1298
rect 7497 1264 7505 1298
rect 7451 1230 7505 1264
rect 7451 1196 7463 1230
rect 7497 1196 7505 1230
rect 7451 1162 7505 1196
rect 7451 1128 7463 1162
rect 7497 1128 7505 1162
rect 7451 1004 7505 1128
rect 7887 1366 7943 1404
rect 7887 1332 7897 1366
rect 7931 1332 7943 1366
rect 7887 1298 7943 1332
rect 7887 1264 7897 1298
rect 7931 1264 7943 1298
rect 7887 1230 7943 1264
rect 7887 1196 7897 1230
rect 7931 1196 7943 1230
rect 7887 1162 7943 1196
rect 7887 1128 7897 1162
rect 7931 1128 7943 1162
rect 7887 1093 7943 1128
rect 7887 1059 7897 1093
rect 7931 1059 7943 1093
rect 7887 1004 7943 1059
rect 7973 1366 8031 1404
rect 7973 1332 7985 1366
rect 8019 1332 8031 1366
rect 7973 1298 8031 1332
rect 7973 1264 7985 1298
rect 8019 1264 8031 1298
rect 7973 1230 8031 1264
rect 7973 1196 7985 1230
rect 8019 1196 8031 1230
rect 7973 1162 8031 1196
rect 7973 1128 7985 1162
rect 8019 1128 8031 1162
rect 7973 1093 8031 1128
rect 7973 1059 7985 1093
rect 8019 1059 8031 1093
rect 7973 1004 8031 1059
rect 8061 1366 8119 1404
rect 8061 1332 8073 1366
rect 8107 1332 8119 1366
rect 8061 1298 8119 1332
rect 8061 1264 8073 1298
rect 8107 1264 8119 1298
rect 8061 1230 8119 1264
rect 8061 1196 8073 1230
rect 8107 1196 8119 1230
rect 8061 1162 8119 1196
rect 8061 1128 8073 1162
rect 8107 1128 8119 1162
rect 8061 1004 8119 1128
rect 8149 1366 8207 1404
rect 8149 1332 8161 1366
rect 8195 1332 8207 1366
rect 8149 1298 8207 1332
rect 8149 1264 8161 1298
rect 8195 1264 8207 1298
rect 8149 1230 8207 1264
rect 8149 1196 8161 1230
rect 8195 1196 8207 1230
rect 8149 1162 8207 1196
rect 8149 1128 8161 1162
rect 8195 1128 8207 1162
rect 8149 1093 8207 1128
rect 8149 1059 8161 1093
rect 8195 1059 8207 1093
rect 8149 1004 8207 1059
rect 8237 1366 8295 1404
rect 8237 1332 8249 1366
rect 8283 1332 8295 1366
rect 8237 1298 8295 1332
rect 8237 1264 8249 1298
rect 8283 1264 8295 1298
rect 8237 1230 8295 1264
rect 8237 1196 8249 1230
rect 8283 1196 8295 1230
rect 8237 1162 8295 1196
rect 8237 1128 8249 1162
rect 8283 1128 8295 1162
rect 8237 1004 8295 1128
rect 8325 1366 8383 1404
rect 8325 1332 8337 1366
rect 8371 1332 8383 1366
rect 8325 1298 8383 1332
rect 8325 1264 8337 1298
rect 8371 1264 8383 1298
rect 8325 1230 8383 1264
rect 8325 1196 8337 1230
rect 8371 1196 8383 1230
rect 8325 1162 8383 1196
rect 8325 1128 8337 1162
rect 8371 1128 8383 1162
rect 8325 1093 8383 1128
rect 8325 1059 8337 1093
rect 8371 1059 8383 1093
rect 8325 1004 8383 1059
rect 8413 1366 8467 1404
rect 8413 1332 8425 1366
rect 8459 1332 8467 1366
rect 8413 1298 8467 1332
rect 8413 1264 8425 1298
rect 8459 1264 8467 1298
rect 8413 1230 8467 1264
rect 8413 1196 8425 1230
rect 8459 1196 8467 1230
rect 8413 1162 8467 1196
rect 8413 1128 8425 1162
rect 8459 1128 8467 1162
rect 8413 1004 8467 1128
rect 8849 1366 8905 1404
rect 8849 1332 8859 1366
rect 8893 1332 8905 1366
rect 8849 1298 8905 1332
rect 8849 1264 8859 1298
rect 8893 1264 8905 1298
rect 8849 1230 8905 1264
rect 8849 1196 8859 1230
rect 8893 1196 8905 1230
rect 8849 1162 8905 1196
rect 8849 1128 8859 1162
rect 8893 1128 8905 1162
rect 8849 1093 8905 1128
rect 8849 1059 8859 1093
rect 8893 1059 8905 1093
rect 8849 1004 8905 1059
rect 8935 1366 8993 1404
rect 8935 1332 8947 1366
rect 8981 1332 8993 1366
rect 8935 1298 8993 1332
rect 8935 1264 8947 1298
rect 8981 1264 8993 1298
rect 8935 1230 8993 1264
rect 8935 1196 8947 1230
rect 8981 1196 8993 1230
rect 8935 1162 8993 1196
rect 8935 1128 8947 1162
rect 8981 1128 8993 1162
rect 8935 1093 8993 1128
rect 8935 1059 8947 1093
rect 8981 1059 8993 1093
rect 8935 1004 8993 1059
rect 9023 1366 9081 1404
rect 9023 1332 9035 1366
rect 9069 1332 9081 1366
rect 9023 1298 9081 1332
rect 9023 1264 9035 1298
rect 9069 1264 9081 1298
rect 9023 1230 9081 1264
rect 9023 1196 9035 1230
rect 9069 1196 9081 1230
rect 9023 1162 9081 1196
rect 9023 1128 9035 1162
rect 9069 1128 9081 1162
rect 9023 1004 9081 1128
rect 9111 1366 9169 1404
rect 9111 1332 9123 1366
rect 9157 1332 9169 1366
rect 9111 1298 9169 1332
rect 9111 1264 9123 1298
rect 9157 1264 9169 1298
rect 9111 1230 9169 1264
rect 9111 1196 9123 1230
rect 9157 1196 9169 1230
rect 9111 1162 9169 1196
rect 9111 1128 9123 1162
rect 9157 1128 9169 1162
rect 9111 1093 9169 1128
rect 9111 1059 9123 1093
rect 9157 1059 9169 1093
rect 9111 1004 9169 1059
rect 9199 1366 9257 1404
rect 9199 1332 9211 1366
rect 9245 1332 9257 1366
rect 9199 1298 9257 1332
rect 9199 1264 9211 1298
rect 9245 1264 9257 1298
rect 9199 1230 9257 1264
rect 9199 1196 9211 1230
rect 9245 1196 9257 1230
rect 9199 1162 9257 1196
rect 9199 1128 9211 1162
rect 9245 1128 9257 1162
rect 9199 1004 9257 1128
rect 9287 1366 9345 1404
rect 9287 1332 9299 1366
rect 9333 1332 9345 1366
rect 9287 1298 9345 1332
rect 9287 1264 9299 1298
rect 9333 1264 9345 1298
rect 9287 1230 9345 1264
rect 9287 1196 9299 1230
rect 9333 1196 9345 1230
rect 9287 1162 9345 1196
rect 9287 1128 9299 1162
rect 9333 1128 9345 1162
rect 9287 1093 9345 1128
rect 9287 1059 9299 1093
rect 9333 1059 9345 1093
rect 9287 1004 9345 1059
rect 9375 1366 9429 1404
rect 9375 1332 9387 1366
rect 9421 1332 9429 1366
rect 9375 1298 9429 1332
rect 9375 1264 9387 1298
rect 9421 1264 9429 1298
rect 9375 1230 9429 1264
rect 9375 1196 9387 1230
rect 9421 1196 9429 1230
rect 9375 1162 9429 1196
rect 9375 1128 9387 1162
rect 9421 1128 9429 1162
rect 9375 1004 9429 1128
rect 9811 1366 9867 1404
rect 9811 1332 9821 1366
rect 9855 1332 9867 1366
rect 9811 1298 9867 1332
rect 9811 1264 9821 1298
rect 9855 1264 9867 1298
rect 9811 1230 9867 1264
rect 9811 1196 9821 1230
rect 9855 1196 9867 1230
rect 9811 1162 9867 1196
rect 9811 1128 9821 1162
rect 9855 1128 9867 1162
rect 9811 1093 9867 1128
rect 9811 1059 9821 1093
rect 9855 1059 9867 1093
rect 9811 1004 9867 1059
rect 9897 1366 9955 1404
rect 9897 1332 9909 1366
rect 9943 1332 9955 1366
rect 9897 1298 9955 1332
rect 9897 1264 9909 1298
rect 9943 1264 9955 1298
rect 9897 1230 9955 1264
rect 9897 1196 9909 1230
rect 9943 1196 9955 1230
rect 9897 1162 9955 1196
rect 9897 1128 9909 1162
rect 9943 1128 9955 1162
rect 9897 1093 9955 1128
rect 9897 1059 9909 1093
rect 9943 1059 9955 1093
rect 9897 1004 9955 1059
rect 9985 1366 10043 1404
rect 9985 1332 9997 1366
rect 10031 1332 10043 1366
rect 9985 1298 10043 1332
rect 9985 1264 9997 1298
rect 10031 1264 10043 1298
rect 9985 1230 10043 1264
rect 9985 1196 9997 1230
rect 10031 1196 10043 1230
rect 9985 1162 10043 1196
rect 9985 1128 9997 1162
rect 10031 1128 10043 1162
rect 9985 1004 10043 1128
rect 10073 1366 10131 1404
rect 10073 1332 10085 1366
rect 10119 1332 10131 1366
rect 10073 1298 10131 1332
rect 10073 1264 10085 1298
rect 10119 1264 10131 1298
rect 10073 1230 10131 1264
rect 10073 1196 10085 1230
rect 10119 1196 10131 1230
rect 10073 1162 10131 1196
rect 10073 1128 10085 1162
rect 10119 1128 10131 1162
rect 10073 1093 10131 1128
rect 10073 1059 10085 1093
rect 10119 1059 10131 1093
rect 10073 1004 10131 1059
rect 10161 1366 10219 1404
rect 10161 1332 10173 1366
rect 10207 1332 10219 1366
rect 10161 1298 10219 1332
rect 10161 1264 10173 1298
rect 10207 1264 10219 1298
rect 10161 1230 10219 1264
rect 10161 1196 10173 1230
rect 10207 1196 10219 1230
rect 10161 1162 10219 1196
rect 10161 1128 10173 1162
rect 10207 1128 10219 1162
rect 10161 1004 10219 1128
rect 10249 1366 10307 1404
rect 10249 1332 10261 1366
rect 10295 1332 10307 1366
rect 10249 1298 10307 1332
rect 10249 1264 10261 1298
rect 10295 1264 10307 1298
rect 10249 1230 10307 1264
rect 10249 1196 10261 1230
rect 10295 1196 10307 1230
rect 10249 1162 10307 1196
rect 10249 1128 10261 1162
rect 10295 1128 10307 1162
rect 10249 1093 10307 1128
rect 10249 1059 10261 1093
rect 10295 1059 10307 1093
rect 10249 1004 10307 1059
rect 10337 1366 10391 1404
rect 10337 1332 10349 1366
rect 10383 1332 10391 1366
rect 10337 1298 10391 1332
rect 10337 1264 10349 1298
rect 10383 1264 10391 1298
rect 10337 1230 10391 1264
rect 10337 1196 10349 1230
rect 10383 1196 10391 1230
rect 10337 1162 10391 1196
rect 10337 1128 10349 1162
rect 10383 1128 10391 1162
rect 10337 1004 10391 1128
rect 10773 1366 10829 1404
rect 10773 1332 10783 1366
rect 10817 1332 10829 1366
rect 10773 1298 10829 1332
rect 10773 1264 10783 1298
rect 10817 1264 10829 1298
rect 10773 1230 10829 1264
rect 10773 1196 10783 1230
rect 10817 1196 10829 1230
rect 10773 1162 10829 1196
rect 10773 1128 10783 1162
rect 10817 1128 10829 1162
rect 10773 1093 10829 1128
rect 10773 1059 10783 1093
rect 10817 1059 10829 1093
rect 10773 1004 10829 1059
rect 10859 1366 10917 1404
rect 10859 1332 10871 1366
rect 10905 1332 10917 1366
rect 10859 1298 10917 1332
rect 10859 1264 10871 1298
rect 10905 1264 10917 1298
rect 10859 1230 10917 1264
rect 10859 1196 10871 1230
rect 10905 1196 10917 1230
rect 10859 1162 10917 1196
rect 10859 1128 10871 1162
rect 10905 1128 10917 1162
rect 10859 1093 10917 1128
rect 10859 1059 10871 1093
rect 10905 1059 10917 1093
rect 10859 1004 10917 1059
rect 10947 1366 11005 1404
rect 10947 1332 10959 1366
rect 10993 1332 11005 1366
rect 10947 1298 11005 1332
rect 10947 1264 10959 1298
rect 10993 1264 11005 1298
rect 10947 1230 11005 1264
rect 10947 1196 10959 1230
rect 10993 1196 11005 1230
rect 10947 1162 11005 1196
rect 10947 1128 10959 1162
rect 10993 1128 11005 1162
rect 10947 1004 11005 1128
rect 11035 1366 11093 1404
rect 11035 1332 11047 1366
rect 11081 1332 11093 1366
rect 11035 1298 11093 1332
rect 11035 1264 11047 1298
rect 11081 1264 11093 1298
rect 11035 1230 11093 1264
rect 11035 1196 11047 1230
rect 11081 1196 11093 1230
rect 11035 1162 11093 1196
rect 11035 1128 11047 1162
rect 11081 1128 11093 1162
rect 11035 1093 11093 1128
rect 11035 1059 11047 1093
rect 11081 1059 11093 1093
rect 11035 1004 11093 1059
rect 11123 1366 11181 1404
rect 11123 1332 11135 1366
rect 11169 1332 11181 1366
rect 11123 1298 11181 1332
rect 11123 1264 11135 1298
rect 11169 1264 11181 1298
rect 11123 1230 11181 1264
rect 11123 1196 11135 1230
rect 11169 1196 11181 1230
rect 11123 1162 11181 1196
rect 11123 1128 11135 1162
rect 11169 1128 11181 1162
rect 11123 1004 11181 1128
rect 11211 1366 11269 1404
rect 11211 1332 11223 1366
rect 11257 1332 11269 1366
rect 11211 1298 11269 1332
rect 11211 1264 11223 1298
rect 11257 1264 11269 1298
rect 11211 1230 11269 1264
rect 11211 1196 11223 1230
rect 11257 1196 11269 1230
rect 11211 1162 11269 1196
rect 11211 1128 11223 1162
rect 11257 1128 11269 1162
rect 11211 1093 11269 1128
rect 11211 1059 11223 1093
rect 11257 1059 11269 1093
rect 11211 1004 11269 1059
rect 11299 1366 11353 1404
rect 11299 1332 11311 1366
rect 11345 1332 11353 1366
rect 11299 1298 11353 1332
rect 11299 1264 11311 1298
rect 11345 1264 11353 1298
rect 11299 1230 11353 1264
rect 11299 1196 11311 1230
rect 11345 1196 11353 1230
rect 11299 1162 11353 1196
rect 11299 1128 11311 1162
rect 11345 1128 11353 1162
rect 11299 1004 11353 1128
rect 11735 1366 11791 1404
rect 11735 1332 11745 1366
rect 11779 1332 11791 1366
rect 11735 1298 11791 1332
rect 11735 1264 11745 1298
rect 11779 1264 11791 1298
rect 11735 1230 11791 1264
rect 11735 1196 11745 1230
rect 11779 1196 11791 1230
rect 11735 1162 11791 1196
rect 11735 1128 11745 1162
rect 11779 1128 11791 1162
rect 11735 1093 11791 1128
rect 11735 1059 11745 1093
rect 11779 1059 11791 1093
rect 11735 1004 11791 1059
rect 11821 1366 11879 1404
rect 11821 1332 11833 1366
rect 11867 1332 11879 1366
rect 11821 1298 11879 1332
rect 11821 1264 11833 1298
rect 11867 1264 11879 1298
rect 11821 1230 11879 1264
rect 11821 1196 11833 1230
rect 11867 1196 11879 1230
rect 11821 1162 11879 1196
rect 11821 1128 11833 1162
rect 11867 1128 11879 1162
rect 11821 1093 11879 1128
rect 11821 1059 11833 1093
rect 11867 1059 11879 1093
rect 11821 1004 11879 1059
rect 11909 1366 11967 1404
rect 11909 1332 11921 1366
rect 11955 1332 11967 1366
rect 11909 1298 11967 1332
rect 11909 1264 11921 1298
rect 11955 1264 11967 1298
rect 11909 1230 11967 1264
rect 11909 1196 11921 1230
rect 11955 1196 11967 1230
rect 11909 1162 11967 1196
rect 11909 1128 11921 1162
rect 11955 1128 11967 1162
rect 11909 1004 11967 1128
rect 11997 1366 12055 1404
rect 11997 1332 12009 1366
rect 12043 1332 12055 1366
rect 11997 1298 12055 1332
rect 11997 1264 12009 1298
rect 12043 1264 12055 1298
rect 11997 1230 12055 1264
rect 11997 1196 12009 1230
rect 12043 1196 12055 1230
rect 11997 1162 12055 1196
rect 11997 1128 12009 1162
rect 12043 1128 12055 1162
rect 11997 1093 12055 1128
rect 11997 1059 12009 1093
rect 12043 1059 12055 1093
rect 11997 1004 12055 1059
rect 12085 1366 12143 1404
rect 12085 1332 12097 1366
rect 12131 1332 12143 1366
rect 12085 1298 12143 1332
rect 12085 1264 12097 1298
rect 12131 1264 12143 1298
rect 12085 1230 12143 1264
rect 12085 1196 12097 1230
rect 12131 1196 12143 1230
rect 12085 1162 12143 1196
rect 12085 1128 12097 1162
rect 12131 1128 12143 1162
rect 12085 1004 12143 1128
rect 12173 1366 12231 1404
rect 12173 1332 12185 1366
rect 12219 1332 12231 1366
rect 12173 1298 12231 1332
rect 12173 1264 12185 1298
rect 12219 1264 12231 1298
rect 12173 1230 12231 1264
rect 12173 1196 12185 1230
rect 12219 1196 12231 1230
rect 12173 1162 12231 1196
rect 12173 1128 12185 1162
rect 12219 1128 12231 1162
rect 12173 1093 12231 1128
rect 12173 1059 12185 1093
rect 12219 1059 12231 1093
rect 12173 1004 12231 1059
rect 12261 1366 12315 1404
rect 12261 1332 12273 1366
rect 12307 1332 12315 1366
rect 12261 1298 12315 1332
rect 12261 1264 12273 1298
rect 12307 1264 12315 1298
rect 12261 1230 12315 1264
rect 12261 1196 12273 1230
rect 12307 1196 12315 1230
rect 12261 1162 12315 1196
rect 12261 1128 12273 1162
rect 12307 1128 12315 1162
rect 12261 1004 12315 1128
rect 12697 1366 12753 1404
rect 12697 1332 12707 1366
rect 12741 1332 12753 1366
rect 12697 1298 12753 1332
rect 12697 1264 12707 1298
rect 12741 1264 12753 1298
rect 12697 1230 12753 1264
rect 12697 1196 12707 1230
rect 12741 1196 12753 1230
rect 12697 1162 12753 1196
rect 12697 1128 12707 1162
rect 12741 1128 12753 1162
rect 12697 1093 12753 1128
rect 12697 1059 12707 1093
rect 12741 1059 12753 1093
rect 12697 1004 12753 1059
rect 12783 1366 12841 1404
rect 12783 1332 12795 1366
rect 12829 1332 12841 1366
rect 12783 1298 12841 1332
rect 12783 1264 12795 1298
rect 12829 1264 12841 1298
rect 12783 1230 12841 1264
rect 12783 1196 12795 1230
rect 12829 1196 12841 1230
rect 12783 1162 12841 1196
rect 12783 1128 12795 1162
rect 12829 1128 12841 1162
rect 12783 1093 12841 1128
rect 12783 1059 12795 1093
rect 12829 1059 12841 1093
rect 12783 1004 12841 1059
rect 12871 1366 12929 1404
rect 12871 1332 12883 1366
rect 12917 1332 12929 1366
rect 12871 1298 12929 1332
rect 12871 1264 12883 1298
rect 12917 1264 12929 1298
rect 12871 1230 12929 1264
rect 12871 1196 12883 1230
rect 12917 1196 12929 1230
rect 12871 1162 12929 1196
rect 12871 1128 12883 1162
rect 12917 1128 12929 1162
rect 12871 1004 12929 1128
rect 12959 1366 13017 1404
rect 12959 1332 12971 1366
rect 13005 1332 13017 1366
rect 12959 1298 13017 1332
rect 12959 1264 12971 1298
rect 13005 1264 13017 1298
rect 12959 1230 13017 1264
rect 12959 1196 12971 1230
rect 13005 1196 13017 1230
rect 12959 1162 13017 1196
rect 12959 1128 12971 1162
rect 13005 1128 13017 1162
rect 12959 1093 13017 1128
rect 12959 1059 12971 1093
rect 13005 1059 13017 1093
rect 12959 1004 13017 1059
rect 13047 1366 13105 1404
rect 13047 1332 13059 1366
rect 13093 1332 13105 1366
rect 13047 1298 13105 1332
rect 13047 1264 13059 1298
rect 13093 1264 13105 1298
rect 13047 1230 13105 1264
rect 13047 1196 13059 1230
rect 13093 1196 13105 1230
rect 13047 1162 13105 1196
rect 13047 1128 13059 1162
rect 13093 1128 13105 1162
rect 13047 1004 13105 1128
rect 13135 1366 13193 1404
rect 13135 1332 13147 1366
rect 13181 1332 13193 1366
rect 13135 1298 13193 1332
rect 13135 1264 13147 1298
rect 13181 1264 13193 1298
rect 13135 1230 13193 1264
rect 13135 1196 13147 1230
rect 13181 1196 13193 1230
rect 13135 1162 13193 1196
rect 13135 1128 13147 1162
rect 13181 1128 13193 1162
rect 13135 1093 13193 1128
rect 13135 1059 13147 1093
rect 13181 1059 13193 1093
rect 13135 1004 13193 1059
rect 13223 1366 13277 1404
rect 13223 1332 13235 1366
rect 13269 1332 13277 1366
rect 13223 1298 13277 1332
rect 13223 1264 13235 1298
rect 13269 1264 13277 1298
rect 13223 1230 13277 1264
rect 13223 1196 13235 1230
rect 13269 1196 13277 1230
rect 13223 1162 13277 1196
rect 13223 1128 13235 1162
rect 13269 1128 13277 1162
rect 13223 1004 13277 1128
rect 13659 1366 13715 1404
rect 13659 1332 13669 1366
rect 13703 1332 13715 1366
rect 13659 1298 13715 1332
rect 13659 1264 13669 1298
rect 13703 1264 13715 1298
rect 13659 1230 13715 1264
rect 13659 1196 13669 1230
rect 13703 1196 13715 1230
rect 13659 1162 13715 1196
rect 13659 1128 13669 1162
rect 13703 1128 13715 1162
rect 13659 1093 13715 1128
rect 13659 1059 13669 1093
rect 13703 1059 13715 1093
rect 13659 1004 13715 1059
rect 13745 1366 13803 1404
rect 13745 1332 13757 1366
rect 13791 1332 13803 1366
rect 13745 1298 13803 1332
rect 13745 1264 13757 1298
rect 13791 1264 13803 1298
rect 13745 1230 13803 1264
rect 13745 1196 13757 1230
rect 13791 1196 13803 1230
rect 13745 1162 13803 1196
rect 13745 1128 13757 1162
rect 13791 1128 13803 1162
rect 13745 1093 13803 1128
rect 13745 1059 13757 1093
rect 13791 1059 13803 1093
rect 13745 1004 13803 1059
rect 13833 1366 13891 1404
rect 13833 1332 13845 1366
rect 13879 1332 13891 1366
rect 13833 1298 13891 1332
rect 13833 1264 13845 1298
rect 13879 1264 13891 1298
rect 13833 1230 13891 1264
rect 13833 1196 13845 1230
rect 13879 1196 13891 1230
rect 13833 1162 13891 1196
rect 13833 1128 13845 1162
rect 13879 1128 13891 1162
rect 13833 1004 13891 1128
rect 13921 1366 13979 1404
rect 13921 1332 13933 1366
rect 13967 1332 13979 1366
rect 13921 1298 13979 1332
rect 13921 1264 13933 1298
rect 13967 1264 13979 1298
rect 13921 1230 13979 1264
rect 13921 1196 13933 1230
rect 13967 1196 13979 1230
rect 13921 1162 13979 1196
rect 13921 1128 13933 1162
rect 13967 1128 13979 1162
rect 13921 1093 13979 1128
rect 13921 1059 13933 1093
rect 13967 1059 13979 1093
rect 13921 1004 13979 1059
rect 14009 1366 14067 1404
rect 14009 1332 14021 1366
rect 14055 1332 14067 1366
rect 14009 1298 14067 1332
rect 14009 1264 14021 1298
rect 14055 1264 14067 1298
rect 14009 1230 14067 1264
rect 14009 1196 14021 1230
rect 14055 1196 14067 1230
rect 14009 1162 14067 1196
rect 14009 1128 14021 1162
rect 14055 1128 14067 1162
rect 14009 1004 14067 1128
rect 14097 1366 14155 1404
rect 14097 1332 14109 1366
rect 14143 1332 14155 1366
rect 14097 1298 14155 1332
rect 14097 1264 14109 1298
rect 14143 1264 14155 1298
rect 14097 1230 14155 1264
rect 14097 1196 14109 1230
rect 14143 1196 14155 1230
rect 14097 1162 14155 1196
rect 14097 1128 14109 1162
rect 14143 1128 14155 1162
rect 14097 1093 14155 1128
rect 14097 1059 14109 1093
rect 14143 1059 14155 1093
rect 14097 1004 14155 1059
rect 14185 1366 14239 1404
rect 14185 1332 14197 1366
rect 14231 1332 14239 1366
rect 14185 1298 14239 1332
rect 14185 1264 14197 1298
rect 14231 1264 14239 1298
rect 14185 1230 14239 1264
rect 14185 1196 14197 1230
rect 14231 1196 14239 1230
rect 14185 1162 14239 1196
rect 14185 1128 14197 1162
rect 14231 1128 14239 1162
rect 14185 1004 14239 1128
rect 14621 1366 14677 1404
rect 14621 1332 14631 1366
rect 14665 1332 14677 1366
rect 14621 1298 14677 1332
rect 14621 1264 14631 1298
rect 14665 1264 14677 1298
rect 14621 1230 14677 1264
rect 14621 1196 14631 1230
rect 14665 1196 14677 1230
rect 14621 1162 14677 1196
rect 14621 1128 14631 1162
rect 14665 1128 14677 1162
rect 14621 1093 14677 1128
rect 14621 1059 14631 1093
rect 14665 1059 14677 1093
rect 14621 1004 14677 1059
rect 14707 1366 14765 1404
rect 14707 1332 14719 1366
rect 14753 1332 14765 1366
rect 14707 1298 14765 1332
rect 14707 1264 14719 1298
rect 14753 1264 14765 1298
rect 14707 1230 14765 1264
rect 14707 1196 14719 1230
rect 14753 1196 14765 1230
rect 14707 1162 14765 1196
rect 14707 1128 14719 1162
rect 14753 1128 14765 1162
rect 14707 1093 14765 1128
rect 14707 1059 14719 1093
rect 14753 1059 14765 1093
rect 14707 1004 14765 1059
rect 14795 1366 14853 1404
rect 14795 1332 14807 1366
rect 14841 1332 14853 1366
rect 14795 1298 14853 1332
rect 14795 1264 14807 1298
rect 14841 1264 14853 1298
rect 14795 1230 14853 1264
rect 14795 1196 14807 1230
rect 14841 1196 14853 1230
rect 14795 1162 14853 1196
rect 14795 1128 14807 1162
rect 14841 1128 14853 1162
rect 14795 1004 14853 1128
rect 14883 1366 14941 1404
rect 14883 1332 14895 1366
rect 14929 1332 14941 1366
rect 14883 1298 14941 1332
rect 14883 1264 14895 1298
rect 14929 1264 14941 1298
rect 14883 1230 14941 1264
rect 14883 1196 14895 1230
rect 14929 1196 14941 1230
rect 14883 1162 14941 1196
rect 14883 1128 14895 1162
rect 14929 1128 14941 1162
rect 14883 1093 14941 1128
rect 14883 1059 14895 1093
rect 14929 1059 14941 1093
rect 14883 1004 14941 1059
rect 14971 1366 15029 1404
rect 14971 1332 14983 1366
rect 15017 1332 15029 1366
rect 14971 1298 15029 1332
rect 14971 1264 14983 1298
rect 15017 1264 15029 1298
rect 14971 1230 15029 1264
rect 14971 1196 14983 1230
rect 15017 1196 15029 1230
rect 14971 1162 15029 1196
rect 14971 1128 14983 1162
rect 15017 1128 15029 1162
rect 14971 1004 15029 1128
rect 15059 1366 15117 1404
rect 15059 1332 15071 1366
rect 15105 1332 15117 1366
rect 15059 1298 15117 1332
rect 15059 1264 15071 1298
rect 15105 1264 15117 1298
rect 15059 1230 15117 1264
rect 15059 1196 15071 1230
rect 15105 1196 15117 1230
rect 15059 1162 15117 1196
rect 15059 1128 15071 1162
rect 15105 1128 15117 1162
rect 15059 1093 15117 1128
rect 15059 1059 15071 1093
rect 15105 1059 15117 1093
rect 15059 1004 15117 1059
rect 15147 1366 15201 1404
rect 15147 1332 15159 1366
rect 15193 1332 15201 1366
rect 15147 1298 15201 1332
rect 15147 1264 15159 1298
rect 15193 1264 15201 1298
rect 15147 1230 15201 1264
rect 15147 1196 15159 1230
rect 15193 1196 15201 1230
rect 15147 1162 15201 1196
rect 15147 1128 15159 1162
rect 15193 1128 15201 1162
rect 15147 1004 15201 1128
rect 15583 1366 15639 1404
rect 15583 1332 15593 1366
rect 15627 1332 15639 1366
rect 15583 1298 15639 1332
rect 15583 1264 15593 1298
rect 15627 1264 15639 1298
rect 15583 1230 15639 1264
rect 15583 1196 15593 1230
rect 15627 1196 15639 1230
rect 15583 1162 15639 1196
rect 15583 1128 15593 1162
rect 15627 1128 15639 1162
rect 15583 1093 15639 1128
rect 15583 1059 15593 1093
rect 15627 1059 15639 1093
rect 15583 1004 15639 1059
rect 15669 1366 15727 1404
rect 15669 1332 15681 1366
rect 15715 1332 15727 1366
rect 15669 1298 15727 1332
rect 15669 1264 15681 1298
rect 15715 1264 15727 1298
rect 15669 1230 15727 1264
rect 15669 1196 15681 1230
rect 15715 1196 15727 1230
rect 15669 1162 15727 1196
rect 15669 1128 15681 1162
rect 15715 1128 15727 1162
rect 15669 1093 15727 1128
rect 15669 1059 15681 1093
rect 15715 1059 15727 1093
rect 15669 1004 15727 1059
rect 15757 1366 15815 1404
rect 15757 1332 15769 1366
rect 15803 1332 15815 1366
rect 15757 1298 15815 1332
rect 15757 1264 15769 1298
rect 15803 1264 15815 1298
rect 15757 1230 15815 1264
rect 15757 1196 15769 1230
rect 15803 1196 15815 1230
rect 15757 1162 15815 1196
rect 15757 1128 15769 1162
rect 15803 1128 15815 1162
rect 15757 1004 15815 1128
rect 15845 1366 15903 1404
rect 15845 1332 15857 1366
rect 15891 1332 15903 1366
rect 15845 1298 15903 1332
rect 15845 1264 15857 1298
rect 15891 1264 15903 1298
rect 15845 1230 15903 1264
rect 15845 1196 15857 1230
rect 15891 1196 15903 1230
rect 15845 1162 15903 1196
rect 15845 1128 15857 1162
rect 15891 1128 15903 1162
rect 15845 1093 15903 1128
rect 15845 1059 15857 1093
rect 15891 1059 15903 1093
rect 15845 1004 15903 1059
rect 15933 1366 15991 1404
rect 15933 1332 15945 1366
rect 15979 1332 15991 1366
rect 15933 1298 15991 1332
rect 15933 1264 15945 1298
rect 15979 1264 15991 1298
rect 15933 1230 15991 1264
rect 15933 1196 15945 1230
rect 15979 1196 15991 1230
rect 15933 1162 15991 1196
rect 15933 1128 15945 1162
rect 15979 1128 15991 1162
rect 15933 1004 15991 1128
rect 16021 1366 16079 1404
rect 16021 1332 16033 1366
rect 16067 1332 16079 1366
rect 16021 1298 16079 1332
rect 16021 1264 16033 1298
rect 16067 1264 16079 1298
rect 16021 1230 16079 1264
rect 16021 1196 16033 1230
rect 16067 1196 16079 1230
rect 16021 1162 16079 1196
rect 16021 1128 16033 1162
rect 16067 1128 16079 1162
rect 16021 1093 16079 1128
rect 16021 1059 16033 1093
rect 16067 1059 16079 1093
rect 16021 1004 16079 1059
rect 16109 1366 16163 1404
rect 16109 1332 16121 1366
rect 16155 1332 16163 1366
rect 16109 1298 16163 1332
rect 16109 1264 16121 1298
rect 16155 1264 16163 1298
rect 16109 1230 16163 1264
rect 16109 1196 16121 1230
rect 16155 1196 16163 1230
rect 16109 1162 16163 1196
rect 16109 1128 16121 1162
rect 16155 1128 16163 1162
rect 16109 1004 16163 1128
rect 16545 1366 16601 1404
rect 16545 1332 16555 1366
rect 16589 1332 16601 1366
rect 16545 1298 16601 1332
rect 16545 1264 16555 1298
rect 16589 1264 16601 1298
rect 16545 1230 16601 1264
rect 16545 1196 16555 1230
rect 16589 1196 16601 1230
rect 16545 1162 16601 1196
rect 16545 1128 16555 1162
rect 16589 1128 16601 1162
rect 16545 1093 16601 1128
rect 16545 1059 16555 1093
rect 16589 1059 16601 1093
rect 16545 1004 16601 1059
rect 16631 1366 16689 1404
rect 16631 1332 16643 1366
rect 16677 1332 16689 1366
rect 16631 1298 16689 1332
rect 16631 1264 16643 1298
rect 16677 1264 16689 1298
rect 16631 1230 16689 1264
rect 16631 1196 16643 1230
rect 16677 1196 16689 1230
rect 16631 1162 16689 1196
rect 16631 1128 16643 1162
rect 16677 1128 16689 1162
rect 16631 1093 16689 1128
rect 16631 1059 16643 1093
rect 16677 1059 16689 1093
rect 16631 1004 16689 1059
rect 16719 1366 16777 1404
rect 16719 1332 16731 1366
rect 16765 1332 16777 1366
rect 16719 1298 16777 1332
rect 16719 1264 16731 1298
rect 16765 1264 16777 1298
rect 16719 1230 16777 1264
rect 16719 1196 16731 1230
rect 16765 1196 16777 1230
rect 16719 1162 16777 1196
rect 16719 1128 16731 1162
rect 16765 1128 16777 1162
rect 16719 1004 16777 1128
rect 16807 1366 16865 1404
rect 16807 1332 16819 1366
rect 16853 1332 16865 1366
rect 16807 1298 16865 1332
rect 16807 1264 16819 1298
rect 16853 1264 16865 1298
rect 16807 1230 16865 1264
rect 16807 1196 16819 1230
rect 16853 1196 16865 1230
rect 16807 1162 16865 1196
rect 16807 1128 16819 1162
rect 16853 1128 16865 1162
rect 16807 1093 16865 1128
rect 16807 1059 16819 1093
rect 16853 1059 16865 1093
rect 16807 1004 16865 1059
rect 16895 1366 16953 1404
rect 16895 1332 16907 1366
rect 16941 1332 16953 1366
rect 16895 1298 16953 1332
rect 16895 1264 16907 1298
rect 16941 1264 16953 1298
rect 16895 1230 16953 1264
rect 16895 1196 16907 1230
rect 16941 1196 16953 1230
rect 16895 1162 16953 1196
rect 16895 1128 16907 1162
rect 16941 1128 16953 1162
rect 16895 1004 16953 1128
rect 16983 1366 17041 1404
rect 16983 1332 16995 1366
rect 17029 1332 17041 1366
rect 16983 1298 17041 1332
rect 16983 1264 16995 1298
rect 17029 1264 17041 1298
rect 16983 1230 17041 1264
rect 16983 1196 16995 1230
rect 17029 1196 17041 1230
rect 16983 1162 17041 1196
rect 16983 1128 16995 1162
rect 17029 1128 17041 1162
rect 16983 1093 17041 1128
rect 16983 1059 16995 1093
rect 17029 1059 17041 1093
rect 16983 1004 17041 1059
rect 17071 1366 17125 1404
rect 17071 1332 17083 1366
rect 17117 1332 17125 1366
rect 17071 1298 17125 1332
rect 17071 1264 17083 1298
rect 17117 1264 17125 1298
rect 17071 1230 17125 1264
rect 17071 1196 17083 1230
rect 17117 1196 17125 1230
rect 17071 1162 17125 1196
rect 17071 1128 17083 1162
rect 17117 1128 17125 1162
rect 17071 1004 17125 1128
rect 17447 1365 17503 1405
rect 17447 1331 17457 1365
rect 17491 1331 17503 1365
rect 17447 1297 17503 1331
rect 17447 1263 17457 1297
rect 17491 1263 17503 1297
rect 17447 1229 17503 1263
rect 17447 1195 17457 1229
rect 17491 1195 17503 1229
rect 17447 1161 17503 1195
rect 17447 1127 17457 1161
rect 17491 1127 17503 1161
rect 17447 1093 17503 1127
rect 17447 1059 17457 1093
rect 17491 1059 17503 1093
rect 17447 1005 17503 1059
rect 17533 1365 17591 1405
rect 17533 1331 17545 1365
rect 17579 1331 17591 1365
rect 17533 1297 17591 1331
rect 17533 1263 17545 1297
rect 17579 1263 17591 1297
rect 17533 1229 17591 1263
rect 17533 1195 17545 1229
rect 17579 1195 17591 1229
rect 17533 1161 17591 1195
rect 17533 1127 17545 1161
rect 17579 1127 17591 1161
rect 17533 1093 17591 1127
rect 17533 1059 17545 1093
rect 17579 1059 17591 1093
rect 17533 1005 17591 1059
rect 17621 1365 17679 1405
rect 17621 1331 17633 1365
rect 17667 1331 17679 1365
rect 17621 1297 17679 1331
rect 17621 1263 17633 1297
rect 17667 1263 17679 1297
rect 17621 1229 17679 1263
rect 17621 1195 17633 1229
rect 17667 1195 17679 1229
rect 17621 1161 17679 1195
rect 17621 1127 17633 1161
rect 17667 1127 17679 1161
rect 17621 1005 17679 1127
rect 17709 1365 17767 1405
rect 17709 1331 17721 1365
rect 17755 1331 17767 1365
rect 17709 1297 17767 1331
rect 17709 1263 17721 1297
rect 17755 1263 17767 1297
rect 17709 1229 17767 1263
rect 17709 1195 17721 1229
rect 17755 1195 17767 1229
rect 17709 1161 17767 1195
rect 17709 1127 17721 1161
rect 17755 1127 17767 1161
rect 17709 1005 17767 1127
rect 17797 1365 17851 1405
rect 17797 1331 17809 1365
rect 17843 1331 17851 1365
rect 17797 1297 17851 1331
rect 17797 1263 17809 1297
rect 17843 1263 17851 1297
rect 17797 1229 17851 1263
rect 17797 1195 17809 1229
rect 17843 1195 17851 1229
rect 17797 1161 17851 1195
rect 17797 1127 17809 1161
rect 17843 1127 17851 1161
rect 17797 1093 17851 1127
rect 17797 1059 17809 1093
rect 17843 1059 17851 1093
rect 17797 1005 17851 1059
rect 18113 1365 18167 1405
rect 18113 1331 18121 1365
rect 18155 1331 18167 1365
rect 18113 1297 18167 1331
rect 18113 1263 18121 1297
rect 18155 1263 18167 1297
rect 18113 1229 18167 1263
rect 18113 1195 18121 1229
rect 18155 1195 18167 1229
rect 18113 1161 18167 1195
rect 18113 1127 18121 1161
rect 18155 1127 18167 1161
rect 18113 1005 18167 1127
rect 18197 1297 18255 1405
rect 18197 1263 18209 1297
rect 18243 1263 18255 1297
rect 18197 1229 18255 1263
rect 18197 1195 18209 1229
rect 18243 1195 18255 1229
rect 18197 1161 18255 1195
rect 18197 1127 18209 1161
rect 18243 1127 18255 1161
rect 18197 1093 18255 1127
rect 18197 1059 18209 1093
rect 18243 1059 18255 1093
rect 18197 1005 18255 1059
rect 18285 1365 18343 1405
rect 18285 1331 18297 1365
rect 18331 1331 18343 1365
rect 18285 1297 18343 1331
rect 18285 1263 18297 1297
rect 18331 1263 18343 1297
rect 18285 1229 18343 1263
rect 18285 1195 18297 1229
rect 18331 1195 18343 1229
rect 18285 1161 18343 1195
rect 18285 1127 18297 1161
rect 18331 1127 18343 1161
rect 18285 1005 18343 1127
rect 18373 1297 18431 1405
rect 18373 1263 18385 1297
rect 18419 1263 18431 1297
rect 18373 1229 18431 1263
rect 18373 1195 18385 1229
rect 18419 1195 18431 1229
rect 18373 1161 18431 1195
rect 18373 1127 18385 1161
rect 18419 1127 18431 1161
rect 18373 1005 18431 1127
rect 18461 1365 18517 1405
rect 18461 1331 18473 1365
rect 18507 1331 18517 1365
rect 18461 1297 18517 1331
rect 18461 1263 18473 1297
rect 18507 1263 18517 1297
rect 18461 1229 18517 1263
rect 18461 1195 18473 1229
rect 18507 1195 18517 1229
rect 18461 1161 18517 1195
rect 18461 1127 18473 1161
rect 18507 1127 18517 1161
rect 18461 1005 18517 1127
rect 18779 1365 18835 1405
rect 18779 1331 18789 1365
rect 18823 1331 18835 1365
rect 18779 1297 18835 1331
rect 18779 1263 18789 1297
rect 18823 1263 18835 1297
rect 18779 1229 18835 1263
rect 18779 1195 18789 1229
rect 18823 1195 18835 1229
rect 18779 1161 18835 1195
rect 18779 1127 18789 1161
rect 18823 1127 18835 1161
rect 18779 1005 18835 1127
rect 18865 1297 18923 1405
rect 18865 1263 18877 1297
rect 18911 1263 18923 1297
rect 18865 1229 18923 1263
rect 18865 1195 18877 1229
rect 18911 1195 18923 1229
rect 18865 1161 18923 1195
rect 18865 1127 18877 1161
rect 18911 1127 18923 1161
rect 18865 1093 18923 1127
rect 18865 1059 18877 1093
rect 18911 1059 18923 1093
rect 18865 1005 18923 1059
rect 18953 1365 19011 1405
rect 18953 1331 18965 1365
rect 18999 1331 19011 1365
rect 18953 1297 19011 1331
rect 18953 1263 18965 1297
rect 18999 1263 19011 1297
rect 18953 1229 19011 1263
rect 18953 1195 18965 1229
rect 18999 1195 19011 1229
rect 18953 1161 19011 1195
rect 18953 1127 18965 1161
rect 18999 1127 19011 1161
rect 18953 1005 19011 1127
rect 19041 1297 19099 1405
rect 19041 1263 19053 1297
rect 19087 1263 19099 1297
rect 19041 1229 19099 1263
rect 19041 1195 19053 1229
rect 19087 1195 19099 1229
rect 19041 1161 19099 1195
rect 19041 1127 19053 1161
rect 19087 1127 19099 1161
rect 19041 1093 19099 1127
rect 19041 1059 19053 1093
rect 19087 1059 19099 1093
rect 19041 1005 19099 1059
rect 19129 1365 19183 1405
rect 19129 1331 19141 1365
rect 19175 1331 19183 1365
rect 19129 1297 19183 1331
rect 19129 1263 19141 1297
rect 19175 1263 19183 1297
rect 19129 1229 19183 1263
rect 19129 1195 19141 1229
rect 19175 1195 19183 1229
rect 19129 1161 19183 1195
rect 19129 1127 19141 1161
rect 19175 1127 19183 1161
rect 19129 1005 19183 1127
<< ndiffc >>
rect 101 301 135 335
rect 198 301 232 335
rect 295 301 329 335
rect 392 301 426 335
rect 489 301 523 335
rect 101 229 135 263
rect 101 161 135 195
rect 198 176 232 210
rect 295 229 329 263
rect 295 161 329 195
rect 393 182 427 216
rect 101 91 135 125
rect 295 91 329 125
rect 392 91 426 125
rect 489 91 523 125
rect 603 301 637 335
rect 603 229 637 263
rect 603 161 637 195
rect 700 185 734 219
rect 797 229 831 263
rect 797 161 831 195
rect 603 91 637 125
rect 700 91 734 125
rect 797 91 831 125
rect 1063 301 1097 335
rect 1160 301 1194 335
rect 1257 301 1291 335
rect 1354 301 1388 335
rect 1451 301 1485 335
rect 1063 229 1097 263
rect 1063 161 1097 195
rect 1160 176 1194 210
rect 1257 229 1291 263
rect 1257 161 1291 195
rect 1355 182 1389 216
rect 1063 91 1097 125
rect 1257 91 1291 125
rect 1354 91 1388 125
rect 1451 91 1485 125
rect 1565 301 1599 335
rect 1565 229 1599 263
rect 1565 161 1599 195
rect 1662 185 1696 219
rect 1759 229 1793 263
rect 1759 161 1793 195
rect 1565 91 1599 125
rect 1662 91 1696 125
rect 1759 91 1793 125
rect 2025 301 2059 335
rect 2122 301 2156 335
rect 2219 301 2253 335
rect 2316 301 2350 335
rect 2413 301 2447 335
rect 2025 229 2059 263
rect 2025 161 2059 195
rect 2122 176 2156 210
rect 2219 229 2253 263
rect 2219 161 2253 195
rect 2317 182 2351 216
rect 2025 91 2059 125
rect 2219 91 2253 125
rect 2316 91 2350 125
rect 2413 91 2447 125
rect 2527 301 2561 335
rect 2527 229 2561 263
rect 2527 161 2561 195
rect 2624 185 2658 219
rect 2721 229 2755 263
rect 2721 161 2755 195
rect 2527 91 2561 125
rect 2624 91 2658 125
rect 2721 91 2755 125
rect 2987 301 3021 335
rect 3084 301 3118 335
rect 3181 301 3215 335
rect 3278 301 3312 335
rect 3375 301 3409 335
rect 2987 229 3021 263
rect 2987 161 3021 195
rect 3084 176 3118 210
rect 3181 229 3215 263
rect 3181 161 3215 195
rect 3279 182 3313 216
rect 2987 91 3021 125
rect 3181 91 3215 125
rect 3278 91 3312 125
rect 3375 91 3409 125
rect 3489 301 3523 335
rect 3489 229 3523 263
rect 3489 161 3523 195
rect 3586 185 3620 219
rect 3683 229 3717 263
rect 3683 161 3717 195
rect 3489 91 3523 125
rect 3586 91 3620 125
rect 3683 91 3717 125
rect 3949 301 3983 335
rect 4046 301 4080 335
rect 4143 301 4177 335
rect 4240 301 4274 335
rect 4337 301 4371 335
rect 3949 229 3983 263
rect 3949 161 3983 195
rect 4046 176 4080 210
rect 4143 229 4177 263
rect 4143 161 4177 195
rect 4241 182 4275 216
rect 3949 91 3983 125
rect 4143 91 4177 125
rect 4240 91 4274 125
rect 4337 91 4371 125
rect 4451 301 4485 335
rect 4451 229 4485 263
rect 4451 161 4485 195
rect 4548 185 4582 219
rect 4645 229 4679 263
rect 4645 161 4679 195
rect 4451 91 4485 125
rect 4548 91 4582 125
rect 4645 91 4679 125
rect 4911 301 4945 335
rect 5008 301 5042 335
rect 5105 301 5139 335
rect 5202 301 5236 335
rect 5299 301 5333 335
rect 4911 229 4945 263
rect 4911 161 4945 195
rect 5008 176 5042 210
rect 5105 229 5139 263
rect 5105 161 5139 195
rect 5203 182 5237 216
rect 4911 91 4945 125
rect 5105 91 5139 125
rect 5202 91 5236 125
rect 5299 91 5333 125
rect 5413 301 5447 335
rect 5413 229 5447 263
rect 5413 161 5447 195
rect 5510 185 5544 219
rect 5607 229 5641 263
rect 5607 161 5641 195
rect 5413 91 5447 125
rect 5510 91 5544 125
rect 5607 91 5641 125
rect 5873 301 5907 335
rect 5970 301 6004 335
rect 6067 301 6101 335
rect 6164 301 6198 335
rect 6261 301 6295 335
rect 5873 229 5907 263
rect 5873 161 5907 195
rect 5970 176 6004 210
rect 6067 229 6101 263
rect 6067 161 6101 195
rect 6165 182 6199 216
rect 5873 91 5907 125
rect 6067 91 6101 125
rect 6164 91 6198 125
rect 6261 91 6295 125
rect 6375 301 6409 335
rect 6375 229 6409 263
rect 6375 161 6409 195
rect 6472 185 6506 219
rect 6569 229 6603 263
rect 6569 161 6603 195
rect 6375 91 6409 125
rect 6472 91 6506 125
rect 6569 91 6603 125
rect 6835 301 6869 335
rect 6932 301 6966 335
rect 7029 301 7063 335
rect 7126 301 7160 335
rect 7223 301 7257 335
rect 6835 229 6869 263
rect 6835 161 6869 195
rect 6932 176 6966 210
rect 7029 229 7063 263
rect 7029 161 7063 195
rect 7127 182 7161 216
rect 6835 91 6869 125
rect 7029 91 7063 125
rect 7126 91 7160 125
rect 7223 91 7257 125
rect 7337 301 7371 335
rect 7337 229 7371 263
rect 7337 161 7371 195
rect 7434 185 7468 219
rect 7531 229 7565 263
rect 7531 161 7565 195
rect 7337 91 7371 125
rect 7434 91 7468 125
rect 7531 91 7565 125
rect 7797 301 7831 335
rect 7894 301 7928 335
rect 7991 301 8025 335
rect 8088 301 8122 335
rect 8185 301 8219 335
rect 7797 229 7831 263
rect 7797 161 7831 195
rect 7894 176 7928 210
rect 7991 229 8025 263
rect 7991 161 8025 195
rect 8089 182 8123 216
rect 7797 91 7831 125
rect 7991 91 8025 125
rect 8088 91 8122 125
rect 8185 91 8219 125
rect 8299 301 8333 335
rect 8299 229 8333 263
rect 8299 161 8333 195
rect 8396 185 8430 219
rect 8493 229 8527 263
rect 8493 161 8527 195
rect 8299 91 8333 125
rect 8396 91 8430 125
rect 8493 91 8527 125
rect 8759 301 8793 335
rect 8856 301 8890 335
rect 8953 301 8987 335
rect 9050 301 9084 335
rect 9147 301 9181 335
rect 8759 229 8793 263
rect 8759 161 8793 195
rect 8856 176 8890 210
rect 8953 229 8987 263
rect 8953 161 8987 195
rect 9051 182 9085 216
rect 8759 91 8793 125
rect 8953 91 8987 125
rect 9050 91 9084 125
rect 9147 91 9181 125
rect 9261 301 9295 335
rect 9261 229 9295 263
rect 9261 161 9295 195
rect 9358 185 9392 219
rect 9455 229 9489 263
rect 9455 161 9489 195
rect 9261 91 9295 125
rect 9358 91 9392 125
rect 9455 91 9489 125
rect 9721 301 9755 335
rect 9818 301 9852 335
rect 9915 301 9949 335
rect 10012 301 10046 335
rect 10109 301 10143 335
rect 9721 229 9755 263
rect 9721 161 9755 195
rect 9818 176 9852 210
rect 9915 229 9949 263
rect 9915 161 9949 195
rect 10013 182 10047 216
rect 9721 91 9755 125
rect 9915 91 9949 125
rect 10012 91 10046 125
rect 10109 91 10143 125
rect 10223 301 10257 335
rect 10223 229 10257 263
rect 10223 161 10257 195
rect 10320 185 10354 219
rect 10417 229 10451 263
rect 10417 161 10451 195
rect 10223 91 10257 125
rect 10320 91 10354 125
rect 10417 91 10451 125
rect 10683 301 10717 335
rect 10780 301 10814 335
rect 10877 301 10911 335
rect 10974 301 11008 335
rect 11071 301 11105 335
rect 10683 229 10717 263
rect 10683 161 10717 195
rect 10780 176 10814 210
rect 10877 229 10911 263
rect 10877 161 10911 195
rect 10975 182 11009 216
rect 10683 91 10717 125
rect 10877 91 10911 125
rect 10974 91 11008 125
rect 11071 91 11105 125
rect 11185 301 11219 335
rect 11185 229 11219 263
rect 11185 161 11219 195
rect 11282 185 11316 219
rect 11379 229 11413 263
rect 11379 161 11413 195
rect 11185 91 11219 125
rect 11282 91 11316 125
rect 11379 91 11413 125
rect 11645 301 11679 335
rect 11742 301 11776 335
rect 11839 301 11873 335
rect 11936 301 11970 335
rect 12033 301 12067 335
rect 11645 229 11679 263
rect 11645 161 11679 195
rect 11742 176 11776 210
rect 11839 229 11873 263
rect 11839 161 11873 195
rect 11937 182 11971 216
rect 11645 91 11679 125
rect 11839 91 11873 125
rect 11936 91 11970 125
rect 12033 91 12067 125
rect 12147 301 12181 335
rect 12147 229 12181 263
rect 12147 161 12181 195
rect 12244 185 12278 219
rect 12341 229 12375 263
rect 12341 161 12375 195
rect 12147 91 12181 125
rect 12244 91 12278 125
rect 12341 91 12375 125
rect 12607 301 12641 335
rect 12704 301 12738 335
rect 12801 301 12835 335
rect 12898 301 12932 335
rect 12995 301 13029 335
rect 12607 229 12641 263
rect 12607 161 12641 195
rect 12704 176 12738 210
rect 12801 229 12835 263
rect 12801 161 12835 195
rect 12899 182 12933 216
rect 12607 91 12641 125
rect 12801 91 12835 125
rect 12898 91 12932 125
rect 12995 91 13029 125
rect 13109 301 13143 335
rect 13109 229 13143 263
rect 13109 161 13143 195
rect 13206 185 13240 219
rect 13303 229 13337 263
rect 13303 161 13337 195
rect 13109 91 13143 125
rect 13206 91 13240 125
rect 13303 91 13337 125
rect 13569 301 13603 335
rect 13666 301 13700 335
rect 13763 301 13797 335
rect 13860 301 13894 335
rect 13957 301 13991 335
rect 13569 229 13603 263
rect 13569 161 13603 195
rect 13666 176 13700 210
rect 13763 229 13797 263
rect 13763 161 13797 195
rect 13861 182 13895 216
rect 13569 91 13603 125
rect 13763 91 13797 125
rect 13860 91 13894 125
rect 13957 91 13991 125
rect 14071 301 14105 335
rect 14071 229 14105 263
rect 14071 161 14105 195
rect 14168 185 14202 219
rect 14265 229 14299 263
rect 14265 161 14299 195
rect 14071 91 14105 125
rect 14168 91 14202 125
rect 14265 91 14299 125
rect 14531 301 14565 335
rect 14628 301 14662 335
rect 14725 301 14759 335
rect 14822 301 14856 335
rect 14919 301 14953 335
rect 14531 229 14565 263
rect 14531 161 14565 195
rect 14628 176 14662 210
rect 14725 229 14759 263
rect 14725 161 14759 195
rect 14823 182 14857 216
rect 14531 91 14565 125
rect 14725 91 14759 125
rect 14822 91 14856 125
rect 14919 91 14953 125
rect 15033 301 15067 335
rect 15033 229 15067 263
rect 15033 161 15067 195
rect 15130 185 15164 219
rect 15227 229 15261 263
rect 15227 161 15261 195
rect 15033 91 15067 125
rect 15130 91 15164 125
rect 15227 91 15261 125
rect 15493 301 15527 335
rect 15590 301 15624 335
rect 15687 301 15721 335
rect 15784 301 15818 335
rect 15881 301 15915 335
rect 15493 229 15527 263
rect 15493 161 15527 195
rect 15590 176 15624 210
rect 15687 229 15721 263
rect 15687 161 15721 195
rect 15785 182 15819 216
rect 15493 91 15527 125
rect 15687 91 15721 125
rect 15784 91 15818 125
rect 15881 91 15915 125
rect 15995 301 16029 335
rect 15995 229 16029 263
rect 15995 161 16029 195
rect 16092 185 16126 219
rect 16189 229 16223 263
rect 16189 161 16223 195
rect 15995 91 16029 125
rect 16092 91 16126 125
rect 16189 91 16223 125
rect 16455 301 16489 335
rect 16552 301 16586 335
rect 16649 301 16683 335
rect 16746 301 16780 335
rect 16843 301 16877 335
rect 16455 229 16489 263
rect 16455 161 16489 195
rect 16552 176 16586 210
rect 16649 229 16683 263
rect 16649 161 16683 195
rect 16747 182 16781 216
rect 16455 91 16489 125
rect 16649 91 16683 125
rect 16746 91 16780 125
rect 16843 91 16877 125
rect 16957 301 16991 335
rect 16957 229 16991 263
rect 16957 161 16991 195
rect 17054 185 17088 219
rect 17151 229 17185 263
rect 17151 161 17185 195
rect 16957 91 16991 125
rect 17054 91 17088 125
rect 17151 91 17185 125
rect 17438 299 17472 333
rect 17535 299 17569 333
rect 17632 299 17666 333
rect 17826 299 17860 333
rect 17438 227 17472 261
rect 17438 159 17472 193
rect 17535 174 17569 208
rect 17632 227 17666 261
rect 17632 159 17666 193
rect 17728 183 17762 217
rect 17826 227 17860 261
rect 17826 159 17860 193
rect 17438 89 17472 123
rect 17632 89 17666 123
rect 17728 89 17762 123
rect 17826 89 17860 123
rect 18104 299 18138 333
rect 18201 299 18235 333
rect 18298 299 18332 333
rect 18492 299 18526 333
rect 18104 227 18138 261
rect 18104 159 18138 193
rect 18201 174 18235 208
rect 18298 227 18332 261
rect 18298 159 18332 193
rect 18395 183 18429 217
rect 18492 227 18526 261
rect 18492 159 18526 193
rect 18104 89 18138 123
rect 18298 89 18332 123
rect 18395 89 18429 123
rect 18492 89 18526 123
rect 18770 299 18804 333
rect 18867 299 18901 333
rect 18964 299 18998 333
rect 18770 227 18804 261
rect 18770 159 18804 193
rect 18867 174 18901 208
rect 18964 227 18998 261
rect 18964 159 18998 193
rect 19061 183 19095 217
rect 19158 227 19192 261
rect 19158 159 19192 193
rect 18770 89 18804 123
rect 18964 89 18998 123
rect 19061 89 19095 123
rect 19158 89 19192 123
<< pdiffc >>
rect 201 1332 235 1366
rect 201 1264 235 1298
rect 201 1196 235 1230
rect 201 1128 235 1162
rect 201 1059 235 1093
rect 289 1332 323 1366
rect 289 1264 323 1298
rect 289 1196 323 1230
rect 289 1128 323 1162
rect 289 1059 323 1093
rect 377 1332 411 1366
rect 377 1264 411 1298
rect 377 1196 411 1230
rect 377 1128 411 1162
rect 465 1332 499 1366
rect 465 1264 499 1298
rect 465 1196 499 1230
rect 465 1128 499 1162
rect 465 1059 499 1093
rect 553 1332 587 1366
rect 553 1264 587 1298
rect 553 1196 587 1230
rect 553 1128 587 1162
rect 641 1332 675 1366
rect 641 1264 675 1298
rect 641 1196 675 1230
rect 641 1128 675 1162
rect 641 1059 675 1093
rect 729 1332 763 1366
rect 729 1264 763 1298
rect 729 1196 763 1230
rect 729 1128 763 1162
rect 1163 1332 1197 1366
rect 1163 1264 1197 1298
rect 1163 1196 1197 1230
rect 1163 1128 1197 1162
rect 1163 1059 1197 1093
rect 1251 1332 1285 1366
rect 1251 1264 1285 1298
rect 1251 1196 1285 1230
rect 1251 1128 1285 1162
rect 1251 1059 1285 1093
rect 1339 1332 1373 1366
rect 1339 1264 1373 1298
rect 1339 1196 1373 1230
rect 1339 1128 1373 1162
rect 1427 1332 1461 1366
rect 1427 1264 1461 1298
rect 1427 1196 1461 1230
rect 1427 1128 1461 1162
rect 1427 1059 1461 1093
rect 1515 1332 1549 1366
rect 1515 1264 1549 1298
rect 1515 1196 1549 1230
rect 1515 1128 1549 1162
rect 1603 1332 1637 1366
rect 1603 1264 1637 1298
rect 1603 1196 1637 1230
rect 1603 1128 1637 1162
rect 1603 1059 1637 1093
rect 1691 1332 1725 1366
rect 1691 1264 1725 1298
rect 1691 1196 1725 1230
rect 1691 1128 1725 1162
rect 2125 1332 2159 1366
rect 2125 1264 2159 1298
rect 2125 1196 2159 1230
rect 2125 1128 2159 1162
rect 2125 1059 2159 1093
rect 2213 1332 2247 1366
rect 2213 1264 2247 1298
rect 2213 1196 2247 1230
rect 2213 1128 2247 1162
rect 2213 1059 2247 1093
rect 2301 1332 2335 1366
rect 2301 1264 2335 1298
rect 2301 1196 2335 1230
rect 2301 1128 2335 1162
rect 2389 1332 2423 1366
rect 2389 1264 2423 1298
rect 2389 1196 2423 1230
rect 2389 1128 2423 1162
rect 2389 1059 2423 1093
rect 2477 1332 2511 1366
rect 2477 1264 2511 1298
rect 2477 1196 2511 1230
rect 2477 1128 2511 1162
rect 2565 1332 2599 1366
rect 2565 1264 2599 1298
rect 2565 1196 2599 1230
rect 2565 1128 2599 1162
rect 2565 1059 2599 1093
rect 2653 1332 2687 1366
rect 2653 1264 2687 1298
rect 2653 1196 2687 1230
rect 2653 1128 2687 1162
rect 3087 1332 3121 1366
rect 3087 1264 3121 1298
rect 3087 1196 3121 1230
rect 3087 1128 3121 1162
rect 3087 1059 3121 1093
rect 3175 1332 3209 1366
rect 3175 1264 3209 1298
rect 3175 1196 3209 1230
rect 3175 1128 3209 1162
rect 3175 1059 3209 1093
rect 3263 1332 3297 1366
rect 3263 1264 3297 1298
rect 3263 1196 3297 1230
rect 3263 1128 3297 1162
rect 3351 1332 3385 1366
rect 3351 1264 3385 1298
rect 3351 1196 3385 1230
rect 3351 1128 3385 1162
rect 3351 1059 3385 1093
rect 3439 1332 3473 1366
rect 3439 1264 3473 1298
rect 3439 1196 3473 1230
rect 3439 1128 3473 1162
rect 3527 1332 3561 1366
rect 3527 1264 3561 1298
rect 3527 1196 3561 1230
rect 3527 1128 3561 1162
rect 3527 1059 3561 1093
rect 3615 1332 3649 1366
rect 3615 1264 3649 1298
rect 3615 1196 3649 1230
rect 3615 1128 3649 1162
rect 4049 1332 4083 1366
rect 4049 1264 4083 1298
rect 4049 1196 4083 1230
rect 4049 1128 4083 1162
rect 4049 1059 4083 1093
rect 4137 1332 4171 1366
rect 4137 1264 4171 1298
rect 4137 1196 4171 1230
rect 4137 1128 4171 1162
rect 4137 1059 4171 1093
rect 4225 1332 4259 1366
rect 4225 1264 4259 1298
rect 4225 1196 4259 1230
rect 4225 1128 4259 1162
rect 4313 1332 4347 1366
rect 4313 1264 4347 1298
rect 4313 1196 4347 1230
rect 4313 1128 4347 1162
rect 4313 1059 4347 1093
rect 4401 1332 4435 1366
rect 4401 1264 4435 1298
rect 4401 1196 4435 1230
rect 4401 1128 4435 1162
rect 4489 1332 4523 1366
rect 4489 1264 4523 1298
rect 4489 1196 4523 1230
rect 4489 1128 4523 1162
rect 4489 1059 4523 1093
rect 4577 1332 4611 1366
rect 4577 1264 4611 1298
rect 4577 1196 4611 1230
rect 4577 1128 4611 1162
rect 5011 1332 5045 1366
rect 5011 1264 5045 1298
rect 5011 1196 5045 1230
rect 5011 1128 5045 1162
rect 5011 1059 5045 1093
rect 5099 1332 5133 1366
rect 5099 1264 5133 1298
rect 5099 1196 5133 1230
rect 5099 1128 5133 1162
rect 5099 1059 5133 1093
rect 5187 1332 5221 1366
rect 5187 1264 5221 1298
rect 5187 1196 5221 1230
rect 5187 1128 5221 1162
rect 5275 1332 5309 1366
rect 5275 1264 5309 1298
rect 5275 1196 5309 1230
rect 5275 1128 5309 1162
rect 5275 1059 5309 1093
rect 5363 1332 5397 1366
rect 5363 1264 5397 1298
rect 5363 1196 5397 1230
rect 5363 1128 5397 1162
rect 5451 1332 5485 1366
rect 5451 1264 5485 1298
rect 5451 1196 5485 1230
rect 5451 1128 5485 1162
rect 5451 1059 5485 1093
rect 5539 1332 5573 1366
rect 5539 1264 5573 1298
rect 5539 1196 5573 1230
rect 5539 1128 5573 1162
rect 5973 1332 6007 1366
rect 5973 1264 6007 1298
rect 5973 1196 6007 1230
rect 5973 1128 6007 1162
rect 5973 1059 6007 1093
rect 6061 1332 6095 1366
rect 6061 1264 6095 1298
rect 6061 1196 6095 1230
rect 6061 1128 6095 1162
rect 6061 1059 6095 1093
rect 6149 1332 6183 1366
rect 6149 1264 6183 1298
rect 6149 1196 6183 1230
rect 6149 1128 6183 1162
rect 6237 1332 6271 1366
rect 6237 1264 6271 1298
rect 6237 1196 6271 1230
rect 6237 1128 6271 1162
rect 6237 1059 6271 1093
rect 6325 1332 6359 1366
rect 6325 1264 6359 1298
rect 6325 1196 6359 1230
rect 6325 1128 6359 1162
rect 6413 1332 6447 1366
rect 6413 1264 6447 1298
rect 6413 1196 6447 1230
rect 6413 1128 6447 1162
rect 6413 1059 6447 1093
rect 6501 1332 6535 1366
rect 6501 1264 6535 1298
rect 6501 1196 6535 1230
rect 6501 1128 6535 1162
rect 6935 1332 6969 1366
rect 6935 1264 6969 1298
rect 6935 1196 6969 1230
rect 6935 1128 6969 1162
rect 6935 1059 6969 1093
rect 7023 1332 7057 1366
rect 7023 1264 7057 1298
rect 7023 1196 7057 1230
rect 7023 1128 7057 1162
rect 7023 1059 7057 1093
rect 7111 1332 7145 1366
rect 7111 1264 7145 1298
rect 7111 1196 7145 1230
rect 7111 1128 7145 1162
rect 7199 1332 7233 1366
rect 7199 1264 7233 1298
rect 7199 1196 7233 1230
rect 7199 1128 7233 1162
rect 7199 1059 7233 1093
rect 7287 1332 7321 1366
rect 7287 1264 7321 1298
rect 7287 1196 7321 1230
rect 7287 1128 7321 1162
rect 7375 1332 7409 1366
rect 7375 1264 7409 1298
rect 7375 1196 7409 1230
rect 7375 1128 7409 1162
rect 7375 1059 7409 1093
rect 7463 1332 7497 1366
rect 7463 1264 7497 1298
rect 7463 1196 7497 1230
rect 7463 1128 7497 1162
rect 7897 1332 7931 1366
rect 7897 1264 7931 1298
rect 7897 1196 7931 1230
rect 7897 1128 7931 1162
rect 7897 1059 7931 1093
rect 7985 1332 8019 1366
rect 7985 1264 8019 1298
rect 7985 1196 8019 1230
rect 7985 1128 8019 1162
rect 7985 1059 8019 1093
rect 8073 1332 8107 1366
rect 8073 1264 8107 1298
rect 8073 1196 8107 1230
rect 8073 1128 8107 1162
rect 8161 1332 8195 1366
rect 8161 1264 8195 1298
rect 8161 1196 8195 1230
rect 8161 1128 8195 1162
rect 8161 1059 8195 1093
rect 8249 1332 8283 1366
rect 8249 1264 8283 1298
rect 8249 1196 8283 1230
rect 8249 1128 8283 1162
rect 8337 1332 8371 1366
rect 8337 1264 8371 1298
rect 8337 1196 8371 1230
rect 8337 1128 8371 1162
rect 8337 1059 8371 1093
rect 8425 1332 8459 1366
rect 8425 1264 8459 1298
rect 8425 1196 8459 1230
rect 8425 1128 8459 1162
rect 8859 1332 8893 1366
rect 8859 1264 8893 1298
rect 8859 1196 8893 1230
rect 8859 1128 8893 1162
rect 8859 1059 8893 1093
rect 8947 1332 8981 1366
rect 8947 1264 8981 1298
rect 8947 1196 8981 1230
rect 8947 1128 8981 1162
rect 8947 1059 8981 1093
rect 9035 1332 9069 1366
rect 9035 1264 9069 1298
rect 9035 1196 9069 1230
rect 9035 1128 9069 1162
rect 9123 1332 9157 1366
rect 9123 1264 9157 1298
rect 9123 1196 9157 1230
rect 9123 1128 9157 1162
rect 9123 1059 9157 1093
rect 9211 1332 9245 1366
rect 9211 1264 9245 1298
rect 9211 1196 9245 1230
rect 9211 1128 9245 1162
rect 9299 1332 9333 1366
rect 9299 1264 9333 1298
rect 9299 1196 9333 1230
rect 9299 1128 9333 1162
rect 9299 1059 9333 1093
rect 9387 1332 9421 1366
rect 9387 1264 9421 1298
rect 9387 1196 9421 1230
rect 9387 1128 9421 1162
rect 9821 1332 9855 1366
rect 9821 1264 9855 1298
rect 9821 1196 9855 1230
rect 9821 1128 9855 1162
rect 9821 1059 9855 1093
rect 9909 1332 9943 1366
rect 9909 1264 9943 1298
rect 9909 1196 9943 1230
rect 9909 1128 9943 1162
rect 9909 1059 9943 1093
rect 9997 1332 10031 1366
rect 9997 1264 10031 1298
rect 9997 1196 10031 1230
rect 9997 1128 10031 1162
rect 10085 1332 10119 1366
rect 10085 1264 10119 1298
rect 10085 1196 10119 1230
rect 10085 1128 10119 1162
rect 10085 1059 10119 1093
rect 10173 1332 10207 1366
rect 10173 1264 10207 1298
rect 10173 1196 10207 1230
rect 10173 1128 10207 1162
rect 10261 1332 10295 1366
rect 10261 1264 10295 1298
rect 10261 1196 10295 1230
rect 10261 1128 10295 1162
rect 10261 1059 10295 1093
rect 10349 1332 10383 1366
rect 10349 1264 10383 1298
rect 10349 1196 10383 1230
rect 10349 1128 10383 1162
rect 10783 1332 10817 1366
rect 10783 1264 10817 1298
rect 10783 1196 10817 1230
rect 10783 1128 10817 1162
rect 10783 1059 10817 1093
rect 10871 1332 10905 1366
rect 10871 1264 10905 1298
rect 10871 1196 10905 1230
rect 10871 1128 10905 1162
rect 10871 1059 10905 1093
rect 10959 1332 10993 1366
rect 10959 1264 10993 1298
rect 10959 1196 10993 1230
rect 10959 1128 10993 1162
rect 11047 1332 11081 1366
rect 11047 1264 11081 1298
rect 11047 1196 11081 1230
rect 11047 1128 11081 1162
rect 11047 1059 11081 1093
rect 11135 1332 11169 1366
rect 11135 1264 11169 1298
rect 11135 1196 11169 1230
rect 11135 1128 11169 1162
rect 11223 1332 11257 1366
rect 11223 1264 11257 1298
rect 11223 1196 11257 1230
rect 11223 1128 11257 1162
rect 11223 1059 11257 1093
rect 11311 1332 11345 1366
rect 11311 1264 11345 1298
rect 11311 1196 11345 1230
rect 11311 1128 11345 1162
rect 11745 1332 11779 1366
rect 11745 1264 11779 1298
rect 11745 1196 11779 1230
rect 11745 1128 11779 1162
rect 11745 1059 11779 1093
rect 11833 1332 11867 1366
rect 11833 1264 11867 1298
rect 11833 1196 11867 1230
rect 11833 1128 11867 1162
rect 11833 1059 11867 1093
rect 11921 1332 11955 1366
rect 11921 1264 11955 1298
rect 11921 1196 11955 1230
rect 11921 1128 11955 1162
rect 12009 1332 12043 1366
rect 12009 1264 12043 1298
rect 12009 1196 12043 1230
rect 12009 1128 12043 1162
rect 12009 1059 12043 1093
rect 12097 1332 12131 1366
rect 12097 1264 12131 1298
rect 12097 1196 12131 1230
rect 12097 1128 12131 1162
rect 12185 1332 12219 1366
rect 12185 1264 12219 1298
rect 12185 1196 12219 1230
rect 12185 1128 12219 1162
rect 12185 1059 12219 1093
rect 12273 1332 12307 1366
rect 12273 1264 12307 1298
rect 12273 1196 12307 1230
rect 12273 1128 12307 1162
rect 12707 1332 12741 1366
rect 12707 1264 12741 1298
rect 12707 1196 12741 1230
rect 12707 1128 12741 1162
rect 12707 1059 12741 1093
rect 12795 1332 12829 1366
rect 12795 1264 12829 1298
rect 12795 1196 12829 1230
rect 12795 1128 12829 1162
rect 12795 1059 12829 1093
rect 12883 1332 12917 1366
rect 12883 1264 12917 1298
rect 12883 1196 12917 1230
rect 12883 1128 12917 1162
rect 12971 1332 13005 1366
rect 12971 1264 13005 1298
rect 12971 1196 13005 1230
rect 12971 1128 13005 1162
rect 12971 1059 13005 1093
rect 13059 1332 13093 1366
rect 13059 1264 13093 1298
rect 13059 1196 13093 1230
rect 13059 1128 13093 1162
rect 13147 1332 13181 1366
rect 13147 1264 13181 1298
rect 13147 1196 13181 1230
rect 13147 1128 13181 1162
rect 13147 1059 13181 1093
rect 13235 1332 13269 1366
rect 13235 1264 13269 1298
rect 13235 1196 13269 1230
rect 13235 1128 13269 1162
rect 13669 1332 13703 1366
rect 13669 1264 13703 1298
rect 13669 1196 13703 1230
rect 13669 1128 13703 1162
rect 13669 1059 13703 1093
rect 13757 1332 13791 1366
rect 13757 1264 13791 1298
rect 13757 1196 13791 1230
rect 13757 1128 13791 1162
rect 13757 1059 13791 1093
rect 13845 1332 13879 1366
rect 13845 1264 13879 1298
rect 13845 1196 13879 1230
rect 13845 1128 13879 1162
rect 13933 1332 13967 1366
rect 13933 1264 13967 1298
rect 13933 1196 13967 1230
rect 13933 1128 13967 1162
rect 13933 1059 13967 1093
rect 14021 1332 14055 1366
rect 14021 1264 14055 1298
rect 14021 1196 14055 1230
rect 14021 1128 14055 1162
rect 14109 1332 14143 1366
rect 14109 1264 14143 1298
rect 14109 1196 14143 1230
rect 14109 1128 14143 1162
rect 14109 1059 14143 1093
rect 14197 1332 14231 1366
rect 14197 1264 14231 1298
rect 14197 1196 14231 1230
rect 14197 1128 14231 1162
rect 14631 1332 14665 1366
rect 14631 1264 14665 1298
rect 14631 1196 14665 1230
rect 14631 1128 14665 1162
rect 14631 1059 14665 1093
rect 14719 1332 14753 1366
rect 14719 1264 14753 1298
rect 14719 1196 14753 1230
rect 14719 1128 14753 1162
rect 14719 1059 14753 1093
rect 14807 1332 14841 1366
rect 14807 1264 14841 1298
rect 14807 1196 14841 1230
rect 14807 1128 14841 1162
rect 14895 1332 14929 1366
rect 14895 1264 14929 1298
rect 14895 1196 14929 1230
rect 14895 1128 14929 1162
rect 14895 1059 14929 1093
rect 14983 1332 15017 1366
rect 14983 1264 15017 1298
rect 14983 1196 15017 1230
rect 14983 1128 15017 1162
rect 15071 1332 15105 1366
rect 15071 1264 15105 1298
rect 15071 1196 15105 1230
rect 15071 1128 15105 1162
rect 15071 1059 15105 1093
rect 15159 1332 15193 1366
rect 15159 1264 15193 1298
rect 15159 1196 15193 1230
rect 15159 1128 15193 1162
rect 15593 1332 15627 1366
rect 15593 1264 15627 1298
rect 15593 1196 15627 1230
rect 15593 1128 15627 1162
rect 15593 1059 15627 1093
rect 15681 1332 15715 1366
rect 15681 1264 15715 1298
rect 15681 1196 15715 1230
rect 15681 1128 15715 1162
rect 15681 1059 15715 1093
rect 15769 1332 15803 1366
rect 15769 1264 15803 1298
rect 15769 1196 15803 1230
rect 15769 1128 15803 1162
rect 15857 1332 15891 1366
rect 15857 1264 15891 1298
rect 15857 1196 15891 1230
rect 15857 1128 15891 1162
rect 15857 1059 15891 1093
rect 15945 1332 15979 1366
rect 15945 1264 15979 1298
rect 15945 1196 15979 1230
rect 15945 1128 15979 1162
rect 16033 1332 16067 1366
rect 16033 1264 16067 1298
rect 16033 1196 16067 1230
rect 16033 1128 16067 1162
rect 16033 1059 16067 1093
rect 16121 1332 16155 1366
rect 16121 1264 16155 1298
rect 16121 1196 16155 1230
rect 16121 1128 16155 1162
rect 16555 1332 16589 1366
rect 16555 1264 16589 1298
rect 16555 1196 16589 1230
rect 16555 1128 16589 1162
rect 16555 1059 16589 1093
rect 16643 1332 16677 1366
rect 16643 1264 16677 1298
rect 16643 1196 16677 1230
rect 16643 1128 16677 1162
rect 16643 1059 16677 1093
rect 16731 1332 16765 1366
rect 16731 1264 16765 1298
rect 16731 1196 16765 1230
rect 16731 1128 16765 1162
rect 16819 1332 16853 1366
rect 16819 1264 16853 1298
rect 16819 1196 16853 1230
rect 16819 1128 16853 1162
rect 16819 1059 16853 1093
rect 16907 1332 16941 1366
rect 16907 1264 16941 1298
rect 16907 1196 16941 1230
rect 16907 1128 16941 1162
rect 16995 1332 17029 1366
rect 16995 1264 17029 1298
rect 16995 1196 17029 1230
rect 16995 1128 17029 1162
rect 16995 1059 17029 1093
rect 17083 1332 17117 1366
rect 17083 1264 17117 1298
rect 17083 1196 17117 1230
rect 17083 1128 17117 1162
rect 17457 1331 17491 1365
rect 17457 1263 17491 1297
rect 17457 1195 17491 1229
rect 17457 1127 17491 1161
rect 17457 1059 17491 1093
rect 17545 1331 17579 1365
rect 17545 1263 17579 1297
rect 17545 1195 17579 1229
rect 17545 1127 17579 1161
rect 17545 1059 17579 1093
rect 17633 1331 17667 1365
rect 17633 1263 17667 1297
rect 17633 1195 17667 1229
rect 17633 1127 17667 1161
rect 17721 1331 17755 1365
rect 17721 1263 17755 1297
rect 17721 1195 17755 1229
rect 17721 1127 17755 1161
rect 17809 1331 17843 1365
rect 17809 1263 17843 1297
rect 17809 1195 17843 1229
rect 17809 1127 17843 1161
rect 17809 1059 17843 1093
rect 18121 1331 18155 1365
rect 18121 1263 18155 1297
rect 18121 1195 18155 1229
rect 18121 1127 18155 1161
rect 18209 1263 18243 1297
rect 18209 1195 18243 1229
rect 18209 1127 18243 1161
rect 18209 1059 18243 1093
rect 18297 1331 18331 1365
rect 18297 1263 18331 1297
rect 18297 1195 18331 1229
rect 18297 1127 18331 1161
rect 18385 1263 18419 1297
rect 18385 1195 18419 1229
rect 18385 1127 18419 1161
rect 18473 1331 18507 1365
rect 18473 1263 18507 1297
rect 18473 1195 18507 1229
rect 18473 1127 18507 1161
rect 18789 1331 18823 1365
rect 18789 1263 18823 1297
rect 18789 1195 18823 1229
rect 18789 1127 18823 1161
rect 18877 1263 18911 1297
rect 18877 1195 18911 1229
rect 18877 1127 18911 1161
rect 18877 1059 18911 1093
rect 18965 1331 18999 1365
rect 18965 1263 18999 1297
rect 18965 1195 18999 1229
rect 18965 1127 18999 1161
rect 19053 1263 19087 1297
rect 19053 1195 19087 1229
rect 19053 1127 19087 1161
rect 19053 1059 19087 1093
rect 19141 1331 19175 1365
rect 19141 1263 19175 1297
rect 19141 1195 19175 1229
rect 19141 1127 19175 1161
<< psubdiff >>
rect -34 482 19348 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 928 461 996 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 928 427 945 461
rect 979 427 996 461
rect 1890 461 1958 482
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 928 313 996 353
rect 1890 427 1907 461
rect 1941 427 1958 461
rect 2852 461 2920 482
rect 1890 387 1958 427
rect 1890 353 1907 387
rect 1941 353 1958 387
rect 928 279 945 313
rect 979 279 996 313
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect -34 17 34 57
rect 928 57 945 91
rect 979 57 996 91
rect 1890 313 1958 353
rect 2852 427 2869 461
rect 2903 427 2920 461
rect 3814 461 3882 482
rect 2852 387 2920 427
rect 2852 353 2869 387
rect 2903 353 2920 387
rect 1890 279 1907 313
rect 1941 279 1958 313
rect 1890 239 1958 279
rect 1890 205 1907 239
rect 1941 205 1958 239
rect 1890 165 1958 205
rect 1890 131 1907 165
rect 1941 131 1958 165
rect 1890 91 1958 131
rect 928 17 996 57
rect 1890 57 1907 91
rect 1941 57 1958 91
rect 2852 313 2920 353
rect 3814 427 3831 461
rect 3865 427 3882 461
rect 4776 461 4844 482
rect 3814 387 3882 427
rect 3814 353 3831 387
rect 3865 353 3882 387
rect 2852 279 2869 313
rect 2903 279 2920 313
rect 2852 239 2920 279
rect 2852 205 2869 239
rect 2903 205 2920 239
rect 2852 165 2920 205
rect 2852 131 2869 165
rect 2903 131 2920 165
rect 2852 91 2920 131
rect 1890 17 1958 57
rect 2852 57 2869 91
rect 2903 57 2920 91
rect 3814 313 3882 353
rect 4776 427 4793 461
rect 4827 427 4844 461
rect 5738 461 5806 482
rect 4776 387 4844 427
rect 4776 353 4793 387
rect 4827 353 4844 387
rect 3814 279 3831 313
rect 3865 279 3882 313
rect 3814 239 3882 279
rect 3814 205 3831 239
rect 3865 205 3882 239
rect 3814 165 3882 205
rect 3814 131 3831 165
rect 3865 131 3882 165
rect 3814 91 3882 131
rect 2852 17 2920 57
rect 3814 57 3831 91
rect 3865 57 3882 91
rect 4776 313 4844 353
rect 5738 427 5755 461
rect 5789 427 5806 461
rect 6700 461 6768 482
rect 5738 387 5806 427
rect 5738 353 5755 387
rect 5789 353 5806 387
rect 4776 279 4793 313
rect 4827 279 4844 313
rect 4776 239 4844 279
rect 4776 205 4793 239
rect 4827 205 4844 239
rect 4776 165 4844 205
rect 4776 131 4793 165
rect 4827 131 4844 165
rect 4776 91 4844 131
rect 3814 17 3882 57
rect 4776 57 4793 91
rect 4827 57 4844 91
rect 5738 313 5806 353
rect 6700 427 6717 461
rect 6751 427 6768 461
rect 7662 461 7730 482
rect 6700 387 6768 427
rect 6700 353 6717 387
rect 6751 353 6768 387
rect 5738 279 5755 313
rect 5789 279 5806 313
rect 5738 239 5806 279
rect 5738 205 5755 239
rect 5789 205 5806 239
rect 5738 165 5806 205
rect 5738 131 5755 165
rect 5789 131 5806 165
rect 5738 91 5806 131
rect 4776 17 4844 57
rect 5738 57 5755 91
rect 5789 57 5806 91
rect 6700 313 6768 353
rect 7662 427 7679 461
rect 7713 427 7730 461
rect 8624 461 8692 482
rect 7662 387 7730 427
rect 7662 353 7679 387
rect 7713 353 7730 387
rect 6700 279 6717 313
rect 6751 279 6768 313
rect 6700 239 6768 279
rect 6700 205 6717 239
rect 6751 205 6768 239
rect 6700 165 6768 205
rect 6700 131 6717 165
rect 6751 131 6768 165
rect 6700 91 6768 131
rect 5738 17 5806 57
rect 6700 57 6717 91
rect 6751 57 6768 91
rect 7662 313 7730 353
rect 8624 427 8641 461
rect 8675 427 8692 461
rect 9586 461 9654 482
rect 8624 387 8692 427
rect 8624 353 8641 387
rect 8675 353 8692 387
rect 7662 279 7679 313
rect 7713 279 7730 313
rect 7662 239 7730 279
rect 7662 205 7679 239
rect 7713 205 7730 239
rect 7662 165 7730 205
rect 7662 131 7679 165
rect 7713 131 7730 165
rect 7662 91 7730 131
rect 6700 17 6768 57
rect 7662 57 7679 91
rect 7713 57 7730 91
rect 8624 313 8692 353
rect 9586 427 9603 461
rect 9637 427 9654 461
rect 10548 461 10616 482
rect 9586 387 9654 427
rect 9586 353 9603 387
rect 9637 353 9654 387
rect 8624 279 8641 313
rect 8675 279 8692 313
rect 8624 239 8692 279
rect 8624 205 8641 239
rect 8675 205 8692 239
rect 8624 165 8692 205
rect 8624 131 8641 165
rect 8675 131 8692 165
rect 8624 91 8692 131
rect 7662 17 7730 57
rect 8624 57 8641 91
rect 8675 57 8692 91
rect 9586 313 9654 353
rect 10548 427 10565 461
rect 10599 427 10616 461
rect 11510 461 11578 482
rect 10548 387 10616 427
rect 10548 353 10565 387
rect 10599 353 10616 387
rect 9586 279 9603 313
rect 9637 279 9654 313
rect 9586 239 9654 279
rect 9586 205 9603 239
rect 9637 205 9654 239
rect 9586 165 9654 205
rect 9586 131 9603 165
rect 9637 131 9654 165
rect 9586 91 9654 131
rect 8624 17 8692 57
rect 9586 57 9603 91
rect 9637 57 9654 91
rect 10548 313 10616 353
rect 11510 427 11527 461
rect 11561 427 11578 461
rect 12472 461 12540 482
rect 11510 387 11578 427
rect 11510 353 11527 387
rect 11561 353 11578 387
rect 10548 279 10565 313
rect 10599 279 10616 313
rect 10548 239 10616 279
rect 10548 205 10565 239
rect 10599 205 10616 239
rect 10548 165 10616 205
rect 10548 131 10565 165
rect 10599 131 10616 165
rect 10548 91 10616 131
rect 9586 17 9654 57
rect 10548 57 10565 91
rect 10599 57 10616 91
rect 11510 313 11578 353
rect 12472 427 12489 461
rect 12523 427 12540 461
rect 13434 461 13502 482
rect 12472 387 12540 427
rect 12472 353 12489 387
rect 12523 353 12540 387
rect 11510 279 11527 313
rect 11561 279 11578 313
rect 11510 239 11578 279
rect 11510 205 11527 239
rect 11561 205 11578 239
rect 11510 165 11578 205
rect 11510 131 11527 165
rect 11561 131 11578 165
rect 11510 91 11578 131
rect 10548 17 10616 57
rect 11510 57 11527 91
rect 11561 57 11578 91
rect 12472 313 12540 353
rect 13434 427 13451 461
rect 13485 427 13502 461
rect 14396 461 14464 482
rect 13434 387 13502 427
rect 13434 353 13451 387
rect 13485 353 13502 387
rect 12472 279 12489 313
rect 12523 279 12540 313
rect 12472 239 12540 279
rect 12472 205 12489 239
rect 12523 205 12540 239
rect 12472 165 12540 205
rect 12472 131 12489 165
rect 12523 131 12540 165
rect 12472 91 12540 131
rect 11510 17 11578 57
rect 12472 57 12489 91
rect 12523 57 12540 91
rect 13434 313 13502 353
rect 14396 427 14413 461
rect 14447 427 14464 461
rect 15358 461 15426 482
rect 14396 387 14464 427
rect 14396 353 14413 387
rect 14447 353 14464 387
rect 13434 279 13451 313
rect 13485 279 13502 313
rect 13434 239 13502 279
rect 13434 205 13451 239
rect 13485 205 13502 239
rect 13434 165 13502 205
rect 13434 131 13451 165
rect 13485 131 13502 165
rect 13434 91 13502 131
rect 12472 17 12540 57
rect 13434 57 13451 91
rect 13485 57 13502 91
rect 14396 313 14464 353
rect 15358 427 15375 461
rect 15409 427 15426 461
rect 16320 461 16388 482
rect 15358 387 15426 427
rect 15358 353 15375 387
rect 15409 353 15426 387
rect 14396 279 14413 313
rect 14447 279 14464 313
rect 14396 239 14464 279
rect 14396 205 14413 239
rect 14447 205 14464 239
rect 14396 165 14464 205
rect 14396 131 14413 165
rect 14447 131 14464 165
rect 14396 91 14464 131
rect 13434 17 13502 57
rect 14396 57 14413 91
rect 14447 57 14464 91
rect 15358 313 15426 353
rect 16320 427 16337 461
rect 16371 427 16388 461
rect 17282 461 17350 482
rect 16320 387 16388 427
rect 16320 353 16337 387
rect 16371 353 16388 387
rect 15358 279 15375 313
rect 15409 279 15426 313
rect 15358 239 15426 279
rect 15358 205 15375 239
rect 15409 205 15426 239
rect 15358 165 15426 205
rect 15358 131 15375 165
rect 15409 131 15426 165
rect 15358 91 15426 131
rect 14396 17 14464 57
rect 15358 57 15375 91
rect 15409 57 15426 91
rect 16320 313 16388 353
rect 17282 427 17299 461
rect 17333 427 17350 461
rect 17948 461 18016 482
rect 17282 387 17350 427
rect 17282 353 17299 387
rect 17333 353 17350 387
rect 17948 427 17965 461
rect 17999 427 18016 461
rect 18614 461 18682 482
rect 17948 387 18016 427
rect 16320 279 16337 313
rect 16371 279 16388 313
rect 16320 239 16388 279
rect 16320 205 16337 239
rect 16371 205 16388 239
rect 16320 165 16388 205
rect 16320 131 16337 165
rect 16371 131 16388 165
rect 16320 91 16388 131
rect 15358 17 15426 57
rect 16320 57 16337 91
rect 16371 57 16388 91
rect 17282 313 17350 353
rect 17948 353 17965 387
rect 17999 353 18016 387
rect 17282 279 17299 313
rect 17333 279 17350 313
rect 17282 239 17350 279
rect 17282 205 17299 239
rect 17333 205 17350 239
rect 17282 165 17350 205
rect 17282 131 17299 165
rect 17333 131 17350 165
rect 17282 91 17350 131
rect 16320 17 16388 57
rect 17282 57 17299 91
rect 17333 57 17350 91
rect 17948 313 18016 353
rect 18614 427 18631 461
rect 18665 427 18682 461
rect 19280 461 19348 482
rect 18614 387 18682 427
rect 18614 353 18631 387
rect 18665 353 18682 387
rect 19280 427 19297 461
rect 19331 427 19348 461
rect 19280 387 19348 427
rect 17948 279 17965 313
rect 17999 279 18016 313
rect 17948 239 18016 279
rect 17948 205 17965 239
rect 17999 205 18016 239
rect 17948 165 18016 205
rect 17948 131 17965 165
rect 17999 131 18016 165
rect 17948 91 18016 131
rect 17282 17 17350 57
rect 17948 57 17965 91
rect 17999 57 18016 91
rect 18614 313 18682 353
rect 19280 353 19297 387
rect 19331 353 19348 387
rect 18614 279 18631 313
rect 18665 279 18682 313
rect 18614 239 18682 279
rect 18614 205 18631 239
rect 18665 205 18682 239
rect 18614 165 18682 205
rect 18614 131 18631 165
rect 18665 131 18682 165
rect 18614 91 18682 131
rect 17948 17 18016 57
rect 18614 57 18631 91
rect 18665 57 18682 91
rect 19280 313 19348 353
rect 19280 279 19297 313
rect 19331 279 19348 313
rect 19280 239 19348 279
rect 19280 205 19297 239
rect 19331 205 19348 239
rect 19280 165 19348 205
rect 19280 131 19297 165
rect 19331 131 19348 165
rect 19280 91 19348 131
rect 18614 17 18682 57
rect 19280 57 19297 91
rect 19331 57 19348 91
rect 19280 17 19348 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6569 17
rect 6603 -17 6643 17
rect 6677 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7753 17
rect 7787 -17 7827 17
rect 7861 -17 7901 17
rect 7935 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8123 17
rect 8157 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8567 17
rect 8601 -17 8715 17
rect 8749 -17 8789 17
rect 8823 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9529 17
rect 9563 -17 9677 17
rect 9711 -17 9751 17
rect 9785 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10195 17
rect 10229 -17 10269 17
rect 10303 -17 10343 17
rect 10377 -17 10417 17
rect 10451 -17 10491 17
rect 10525 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10861 17
rect 10895 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11305 17
rect 11339 -17 11379 17
rect 11413 -17 11453 17
rect 11487 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12193 17
rect 12227 -17 12267 17
rect 12301 -17 12341 17
rect 12375 -17 12415 17
rect 12449 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12859 17
rect 12893 -17 12933 17
rect 12967 -17 13007 17
rect 13041 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13525 17
rect 13559 -17 13599 17
rect 13633 -17 13673 17
rect 13707 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13895 17
rect 13929 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14191 17
rect 14225 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14635 17
rect 14669 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14857 17
rect 14891 -17 14931 17
rect 14965 -17 15005 17
rect 15039 -17 15079 17
rect 15113 -17 15153 17
rect 15187 -17 15227 17
rect 15261 -17 15301 17
rect 15335 -17 15449 17
rect 15483 -17 15523 17
rect 15557 -17 15597 17
rect 15631 -17 15671 17
rect 15705 -17 15745 17
rect 15779 -17 15819 17
rect 15853 -17 15893 17
rect 15927 -17 15967 17
rect 16001 -17 16041 17
rect 16075 -17 16115 17
rect 16149 -17 16189 17
rect 16223 -17 16263 17
rect 16297 -17 16411 17
rect 16445 -17 16485 17
rect 16519 -17 16559 17
rect 16593 -17 16633 17
rect 16667 -17 16707 17
rect 16741 -17 16781 17
rect 16815 -17 16855 17
rect 16889 -17 16929 17
rect 16963 -17 17003 17
rect 17037 -17 17077 17
rect 17111 -17 17151 17
rect 17185 -17 17225 17
rect 17259 -17 17373 17
rect 17407 -17 17447 17
rect 17481 -17 17521 17
rect 17555 -17 17595 17
rect 17629 -17 17669 17
rect 17703 -17 17743 17
rect 17777 -17 17817 17
rect 17851 -17 17891 17
rect 17925 -17 18039 17
rect 18073 -17 18113 17
rect 18147 -17 18187 17
rect 18221 -17 18261 17
rect 18295 -17 18335 17
rect 18369 -17 18409 17
rect 18443 -17 18483 17
rect 18517 -17 18557 17
rect 18591 -17 18705 17
rect 18739 -17 18779 17
rect 18813 -17 18853 17
rect 18887 -17 18927 17
rect 18961 -17 19001 17
rect 19035 -17 19075 17
rect 19109 -17 19149 17
rect 19183 -17 19223 17
rect 19257 -17 19348 17
rect -34 -34 19348 -17
<< nsubdiff >>
rect -34 1497 19348 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6569 1497
rect 6603 1463 6643 1497
rect 6677 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7753 1497
rect 7787 1463 7827 1497
rect 7861 1463 7901 1497
rect 7935 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8123 1497
rect 8157 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8567 1497
rect 8601 1463 8715 1497
rect 8749 1463 8789 1497
rect 8823 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9529 1497
rect 9563 1463 9677 1497
rect 9711 1463 9751 1497
rect 9785 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10195 1497
rect 10229 1463 10269 1497
rect 10303 1463 10343 1497
rect 10377 1463 10417 1497
rect 10451 1463 10491 1497
rect 10525 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10861 1497
rect 10895 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11305 1497
rect 11339 1463 11379 1497
rect 11413 1463 11453 1497
rect 11487 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12193 1497
rect 12227 1463 12267 1497
rect 12301 1463 12341 1497
rect 12375 1463 12415 1497
rect 12449 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12859 1497
rect 12893 1463 12933 1497
rect 12967 1463 13007 1497
rect 13041 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13525 1497
rect 13559 1463 13599 1497
rect 13633 1463 13673 1497
rect 13707 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13895 1497
rect 13929 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14191 1497
rect 14225 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14635 1497
rect 14669 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14857 1497
rect 14891 1463 14931 1497
rect 14965 1463 15005 1497
rect 15039 1463 15079 1497
rect 15113 1463 15153 1497
rect 15187 1463 15227 1497
rect 15261 1463 15301 1497
rect 15335 1463 15449 1497
rect 15483 1463 15523 1497
rect 15557 1463 15597 1497
rect 15631 1463 15671 1497
rect 15705 1463 15745 1497
rect 15779 1463 15819 1497
rect 15853 1463 15893 1497
rect 15927 1463 15967 1497
rect 16001 1463 16041 1497
rect 16075 1463 16115 1497
rect 16149 1463 16189 1497
rect 16223 1463 16263 1497
rect 16297 1463 16411 1497
rect 16445 1463 16485 1497
rect 16519 1463 16559 1497
rect 16593 1463 16633 1497
rect 16667 1463 16707 1497
rect 16741 1463 16781 1497
rect 16815 1463 16855 1497
rect 16889 1463 16929 1497
rect 16963 1463 17003 1497
rect 17037 1463 17077 1497
rect 17111 1463 17151 1497
rect 17185 1463 17225 1497
rect 17259 1463 17373 1497
rect 17407 1463 17447 1497
rect 17481 1463 17521 1497
rect 17555 1463 17595 1497
rect 17629 1463 17669 1497
rect 17703 1463 17743 1497
rect 17777 1463 17817 1497
rect 17851 1463 17891 1497
rect 17925 1463 18039 1497
rect 18073 1463 18113 1497
rect 18147 1463 18187 1497
rect 18221 1463 18261 1497
rect 18295 1463 18335 1497
rect 18369 1463 18409 1497
rect 18443 1463 18483 1497
rect 18517 1463 18557 1497
rect 18591 1463 18705 1497
rect 18739 1463 18779 1497
rect 18813 1463 18853 1497
rect 18887 1463 18927 1497
rect 18961 1463 19001 1497
rect 19035 1463 19075 1497
rect 19109 1463 19149 1497
rect 19183 1463 19223 1497
rect 19257 1463 19348 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 928 1423 996 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 1890 1423 1958 1463
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect 928 1019 945 1053
rect 979 1019 996 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 928 979 996 1019
rect 1890 1389 1907 1423
rect 1941 1389 1958 1423
rect 2852 1423 2920 1463
rect 1890 1349 1958 1389
rect 1890 1315 1907 1349
rect 1941 1315 1958 1349
rect 1890 1275 1958 1315
rect 1890 1241 1907 1275
rect 1941 1241 1958 1275
rect 1890 1201 1958 1241
rect 1890 1167 1907 1201
rect 1941 1167 1958 1201
rect 1890 1127 1958 1167
rect 1890 1093 1907 1127
rect 1941 1093 1958 1127
rect 1890 1053 1958 1093
rect 1890 1019 1907 1053
rect 1941 1019 1958 1053
rect 928 945 945 979
rect 979 945 996 979
rect -34 871 -17 905
rect 17 884 34 905
rect 928 905 996 945
rect 1890 979 1958 1019
rect 2852 1389 2869 1423
rect 2903 1389 2920 1423
rect 3814 1423 3882 1463
rect 2852 1349 2920 1389
rect 2852 1315 2869 1349
rect 2903 1315 2920 1349
rect 2852 1275 2920 1315
rect 2852 1241 2869 1275
rect 2903 1241 2920 1275
rect 2852 1201 2920 1241
rect 2852 1167 2869 1201
rect 2903 1167 2920 1201
rect 2852 1127 2920 1167
rect 2852 1093 2869 1127
rect 2903 1093 2920 1127
rect 2852 1053 2920 1093
rect 2852 1019 2869 1053
rect 2903 1019 2920 1053
rect 1890 945 1907 979
rect 1941 945 1958 979
rect 928 884 945 905
rect 17 871 945 884
rect 979 884 996 905
rect 1890 905 1958 945
rect 2852 979 2920 1019
rect 3814 1389 3831 1423
rect 3865 1389 3882 1423
rect 4776 1423 4844 1463
rect 3814 1349 3882 1389
rect 3814 1315 3831 1349
rect 3865 1315 3882 1349
rect 3814 1275 3882 1315
rect 3814 1241 3831 1275
rect 3865 1241 3882 1275
rect 3814 1201 3882 1241
rect 3814 1167 3831 1201
rect 3865 1167 3882 1201
rect 3814 1127 3882 1167
rect 3814 1093 3831 1127
rect 3865 1093 3882 1127
rect 3814 1053 3882 1093
rect 3814 1019 3831 1053
rect 3865 1019 3882 1053
rect 2852 945 2869 979
rect 2903 945 2920 979
rect 1890 884 1907 905
rect 979 871 1907 884
rect 1941 884 1958 905
rect 2852 905 2920 945
rect 3814 979 3882 1019
rect 4776 1389 4793 1423
rect 4827 1389 4844 1423
rect 5738 1423 5806 1463
rect 4776 1349 4844 1389
rect 4776 1315 4793 1349
rect 4827 1315 4844 1349
rect 4776 1275 4844 1315
rect 4776 1241 4793 1275
rect 4827 1241 4844 1275
rect 4776 1201 4844 1241
rect 4776 1167 4793 1201
rect 4827 1167 4844 1201
rect 4776 1127 4844 1167
rect 4776 1093 4793 1127
rect 4827 1093 4844 1127
rect 4776 1053 4844 1093
rect 4776 1019 4793 1053
rect 4827 1019 4844 1053
rect 3814 945 3831 979
rect 3865 945 3882 979
rect 2852 884 2869 905
rect 1941 871 2869 884
rect 2903 884 2920 905
rect 3814 905 3882 945
rect 4776 979 4844 1019
rect 5738 1389 5755 1423
rect 5789 1389 5806 1423
rect 6700 1423 6768 1463
rect 5738 1349 5806 1389
rect 5738 1315 5755 1349
rect 5789 1315 5806 1349
rect 5738 1275 5806 1315
rect 5738 1241 5755 1275
rect 5789 1241 5806 1275
rect 5738 1201 5806 1241
rect 5738 1167 5755 1201
rect 5789 1167 5806 1201
rect 5738 1127 5806 1167
rect 5738 1093 5755 1127
rect 5789 1093 5806 1127
rect 5738 1053 5806 1093
rect 5738 1019 5755 1053
rect 5789 1019 5806 1053
rect 4776 945 4793 979
rect 4827 945 4844 979
rect 3814 884 3831 905
rect 2903 871 3831 884
rect 3865 884 3882 905
rect 4776 905 4844 945
rect 5738 979 5806 1019
rect 6700 1389 6717 1423
rect 6751 1389 6768 1423
rect 7662 1423 7730 1463
rect 6700 1349 6768 1389
rect 6700 1315 6717 1349
rect 6751 1315 6768 1349
rect 6700 1275 6768 1315
rect 6700 1241 6717 1275
rect 6751 1241 6768 1275
rect 6700 1201 6768 1241
rect 6700 1167 6717 1201
rect 6751 1167 6768 1201
rect 6700 1127 6768 1167
rect 6700 1093 6717 1127
rect 6751 1093 6768 1127
rect 6700 1053 6768 1093
rect 6700 1019 6717 1053
rect 6751 1019 6768 1053
rect 5738 945 5755 979
rect 5789 945 5806 979
rect 4776 884 4793 905
rect 3865 871 4793 884
rect 4827 884 4844 905
rect 5738 905 5806 945
rect 6700 979 6768 1019
rect 7662 1389 7679 1423
rect 7713 1389 7730 1423
rect 8624 1423 8692 1463
rect 7662 1349 7730 1389
rect 7662 1315 7679 1349
rect 7713 1315 7730 1349
rect 7662 1275 7730 1315
rect 7662 1241 7679 1275
rect 7713 1241 7730 1275
rect 7662 1201 7730 1241
rect 7662 1167 7679 1201
rect 7713 1167 7730 1201
rect 7662 1127 7730 1167
rect 7662 1093 7679 1127
rect 7713 1093 7730 1127
rect 7662 1053 7730 1093
rect 7662 1019 7679 1053
rect 7713 1019 7730 1053
rect 6700 945 6717 979
rect 6751 945 6768 979
rect 5738 884 5755 905
rect 4827 871 5755 884
rect 5789 884 5806 905
rect 6700 905 6768 945
rect 7662 979 7730 1019
rect 8624 1389 8641 1423
rect 8675 1389 8692 1423
rect 9586 1423 9654 1463
rect 8624 1349 8692 1389
rect 8624 1315 8641 1349
rect 8675 1315 8692 1349
rect 8624 1275 8692 1315
rect 8624 1241 8641 1275
rect 8675 1241 8692 1275
rect 8624 1201 8692 1241
rect 8624 1167 8641 1201
rect 8675 1167 8692 1201
rect 8624 1127 8692 1167
rect 8624 1093 8641 1127
rect 8675 1093 8692 1127
rect 8624 1053 8692 1093
rect 8624 1019 8641 1053
rect 8675 1019 8692 1053
rect 7662 945 7679 979
rect 7713 945 7730 979
rect 6700 884 6717 905
rect 5789 871 6717 884
rect 6751 884 6768 905
rect 7662 905 7730 945
rect 8624 979 8692 1019
rect 9586 1389 9603 1423
rect 9637 1389 9654 1423
rect 10548 1423 10616 1463
rect 9586 1349 9654 1389
rect 9586 1315 9603 1349
rect 9637 1315 9654 1349
rect 9586 1275 9654 1315
rect 9586 1241 9603 1275
rect 9637 1241 9654 1275
rect 9586 1201 9654 1241
rect 9586 1167 9603 1201
rect 9637 1167 9654 1201
rect 9586 1127 9654 1167
rect 9586 1093 9603 1127
rect 9637 1093 9654 1127
rect 9586 1053 9654 1093
rect 9586 1019 9603 1053
rect 9637 1019 9654 1053
rect 8624 945 8641 979
rect 8675 945 8692 979
rect 7662 884 7679 905
rect 6751 871 7679 884
rect 7713 884 7730 905
rect 8624 905 8692 945
rect 9586 979 9654 1019
rect 10548 1389 10565 1423
rect 10599 1389 10616 1423
rect 11510 1423 11578 1463
rect 10548 1349 10616 1389
rect 10548 1315 10565 1349
rect 10599 1315 10616 1349
rect 10548 1275 10616 1315
rect 10548 1241 10565 1275
rect 10599 1241 10616 1275
rect 10548 1201 10616 1241
rect 10548 1167 10565 1201
rect 10599 1167 10616 1201
rect 10548 1127 10616 1167
rect 10548 1093 10565 1127
rect 10599 1093 10616 1127
rect 10548 1053 10616 1093
rect 10548 1019 10565 1053
rect 10599 1019 10616 1053
rect 9586 945 9603 979
rect 9637 945 9654 979
rect 8624 884 8641 905
rect 7713 871 8641 884
rect 8675 884 8692 905
rect 9586 905 9654 945
rect 10548 979 10616 1019
rect 11510 1389 11527 1423
rect 11561 1389 11578 1423
rect 12472 1423 12540 1463
rect 11510 1349 11578 1389
rect 11510 1315 11527 1349
rect 11561 1315 11578 1349
rect 11510 1275 11578 1315
rect 11510 1241 11527 1275
rect 11561 1241 11578 1275
rect 11510 1201 11578 1241
rect 11510 1167 11527 1201
rect 11561 1167 11578 1201
rect 11510 1127 11578 1167
rect 11510 1093 11527 1127
rect 11561 1093 11578 1127
rect 11510 1053 11578 1093
rect 11510 1019 11527 1053
rect 11561 1019 11578 1053
rect 10548 945 10565 979
rect 10599 945 10616 979
rect 9586 884 9603 905
rect 8675 871 9603 884
rect 9637 884 9654 905
rect 10548 905 10616 945
rect 11510 979 11578 1019
rect 12472 1389 12489 1423
rect 12523 1389 12540 1423
rect 13434 1423 13502 1463
rect 12472 1349 12540 1389
rect 12472 1315 12489 1349
rect 12523 1315 12540 1349
rect 12472 1275 12540 1315
rect 12472 1241 12489 1275
rect 12523 1241 12540 1275
rect 12472 1201 12540 1241
rect 12472 1167 12489 1201
rect 12523 1167 12540 1201
rect 12472 1127 12540 1167
rect 12472 1093 12489 1127
rect 12523 1093 12540 1127
rect 12472 1053 12540 1093
rect 12472 1019 12489 1053
rect 12523 1019 12540 1053
rect 11510 945 11527 979
rect 11561 945 11578 979
rect 10548 884 10565 905
rect 9637 871 10565 884
rect 10599 884 10616 905
rect 11510 905 11578 945
rect 12472 979 12540 1019
rect 13434 1389 13451 1423
rect 13485 1389 13502 1423
rect 14396 1423 14464 1463
rect 13434 1349 13502 1389
rect 13434 1315 13451 1349
rect 13485 1315 13502 1349
rect 13434 1275 13502 1315
rect 13434 1241 13451 1275
rect 13485 1241 13502 1275
rect 13434 1201 13502 1241
rect 13434 1167 13451 1201
rect 13485 1167 13502 1201
rect 13434 1127 13502 1167
rect 13434 1093 13451 1127
rect 13485 1093 13502 1127
rect 13434 1053 13502 1093
rect 13434 1019 13451 1053
rect 13485 1019 13502 1053
rect 12472 945 12489 979
rect 12523 945 12540 979
rect 11510 884 11527 905
rect 10599 871 11527 884
rect 11561 884 11578 905
rect 12472 905 12540 945
rect 13434 979 13502 1019
rect 14396 1389 14413 1423
rect 14447 1389 14464 1423
rect 15358 1423 15426 1463
rect 14396 1349 14464 1389
rect 14396 1315 14413 1349
rect 14447 1315 14464 1349
rect 14396 1275 14464 1315
rect 14396 1241 14413 1275
rect 14447 1241 14464 1275
rect 14396 1201 14464 1241
rect 14396 1167 14413 1201
rect 14447 1167 14464 1201
rect 14396 1127 14464 1167
rect 14396 1093 14413 1127
rect 14447 1093 14464 1127
rect 14396 1053 14464 1093
rect 14396 1019 14413 1053
rect 14447 1019 14464 1053
rect 13434 945 13451 979
rect 13485 945 13502 979
rect 12472 884 12489 905
rect 11561 871 12489 884
rect 12523 884 12540 905
rect 13434 905 13502 945
rect 14396 979 14464 1019
rect 15358 1389 15375 1423
rect 15409 1389 15426 1423
rect 16320 1423 16388 1463
rect 15358 1349 15426 1389
rect 15358 1315 15375 1349
rect 15409 1315 15426 1349
rect 15358 1275 15426 1315
rect 15358 1241 15375 1275
rect 15409 1241 15426 1275
rect 15358 1201 15426 1241
rect 15358 1167 15375 1201
rect 15409 1167 15426 1201
rect 15358 1127 15426 1167
rect 15358 1093 15375 1127
rect 15409 1093 15426 1127
rect 15358 1053 15426 1093
rect 15358 1019 15375 1053
rect 15409 1019 15426 1053
rect 14396 945 14413 979
rect 14447 945 14464 979
rect 13434 884 13451 905
rect 12523 871 13451 884
rect 13485 884 13502 905
rect 14396 905 14464 945
rect 15358 979 15426 1019
rect 16320 1389 16337 1423
rect 16371 1389 16388 1423
rect 17282 1423 17350 1463
rect 16320 1349 16388 1389
rect 16320 1315 16337 1349
rect 16371 1315 16388 1349
rect 16320 1275 16388 1315
rect 16320 1241 16337 1275
rect 16371 1241 16388 1275
rect 16320 1201 16388 1241
rect 16320 1167 16337 1201
rect 16371 1167 16388 1201
rect 16320 1127 16388 1167
rect 16320 1093 16337 1127
rect 16371 1093 16388 1127
rect 16320 1053 16388 1093
rect 16320 1019 16337 1053
rect 16371 1019 16388 1053
rect 15358 945 15375 979
rect 15409 945 15426 979
rect 14396 884 14413 905
rect 13485 871 14413 884
rect 14447 884 14464 905
rect 15358 905 15426 945
rect 16320 979 16388 1019
rect 17282 1389 17299 1423
rect 17333 1389 17350 1423
rect 17948 1423 18016 1463
rect 17282 1349 17350 1389
rect 17282 1315 17299 1349
rect 17333 1315 17350 1349
rect 17282 1275 17350 1315
rect 17282 1241 17299 1275
rect 17333 1241 17350 1275
rect 17282 1201 17350 1241
rect 17282 1167 17299 1201
rect 17333 1167 17350 1201
rect 17282 1127 17350 1167
rect 17282 1093 17299 1127
rect 17333 1093 17350 1127
rect 17282 1053 17350 1093
rect 17282 1019 17299 1053
rect 17333 1019 17350 1053
rect 16320 945 16337 979
rect 16371 945 16388 979
rect 15358 884 15375 905
rect 14447 871 15375 884
rect 15409 884 15426 905
rect 16320 905 16388 945
rect 17282 979 17350 1019
rect 17948 1389 17965 1423
rect 17999 1389 18016 1423
rect 18614 1423 18682 1463
rect 19262 1459 19348 1463
rect 17948 1349 18016 1389
rect 17948 1315 17965 1349
rect 17999 1315 18016 1349
rect 17948 1275 18016 1315
rect 17948 1241 17965 1275
rect 17999 1241 18016 1275
rect 17948 1201 18016 1241
rect 17948 1167 17965 1201
rect 17999 1167 18016 1201
rect 17948 1127 18016 1167
rect 17948 1093 17965 1127
rect 17999 1093 18016 1127
rect 17948 1053 18016 1093
rect 17948 1019 17965 1053
rect 17999 1019 18016 1053
rect 17282 945 17299 979
rect 17333 945 17350 979
rect 16320 884 16337 905
rect 15409 871 16337 884
rect 16371 884 16388 905
rect 17282 905 17350 945
rect 17948 979 18016 1019
rect 18614 1389 18631 1423
rect 18665 1389 18682 1423
rect 19280 1423 19348 1459
rect 18614 1349 18682 1389
rect 18614 1315 18631 1349
rect 18665 1315 18682 1349
rect 18614 1275 18682 1315
rect 18614 1241 18631 1275
rect 18665 1241 18682 1275
rect 18614 1201 18682 1241
rect 18614 1167 18631 1201
rect 18665 1167 18682 1201
rect 18614 1127 18682 1167
rect 18614 1093 18631 1127
rect 18665 1093 18682 1127
rect 18614 1053 18682 1093
rect 18614 1019 18631 1053
rect 18665 1019 18682 1053
rect 17948 945 17965 979
rect 17999 945 18016 979
rect 17282 884 17299 905
rect 16371 871 17299 884
rect 17333 884 17350 905
rect 17948 905 18016 945
rect 18614 979 18682 1019
rect 19280 1389 19297 1423
rect 19331 1389 19348 1423
rect 19280 1349 19348 1389
rect 19280 1315 19297 1349
rect 19331 1315 19348 1349
rect 19280 1275 19348 1315
rect 19280 1241 19297 1275
rect 19331 1241 19348 1275
rect 19280 1201 19348 1241
rect 19280 1167 19297 1201
rect 19331 1167 19348 1201
rect 19280 1127 19348 1167
rect 19280 1093 19297 1127
rect 19331 1093 19348 1127
rect 19280 1053 19348 1093
rect 19280 1019 19297 1053
rect 19331 1019 19348 1053
rect 18614 945 18631 979
rect 18665 945 18682 979
rect 17948 884 17965 905
rect 17333 871 17965 884
rect 17999 884 18016 905
rect 18614 905 18682 945
rect 19280 979 19348 1019
rect 19280 945 19297 979
rect 19331 945 19348 979
rect 18614 884 18631 905
rect 17999 871 18631 884
rect 18665 884 18682 905
rect 19280 905 19348 945
rect 19280 884 19297 905
rect 18665 871 19297 884
rect 19331 871 19348 905
rect -34 822 19348 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 945 427 979 461
rect 945 353 979 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1907 427 1941 461
rect 1907 353 1941 387
rect 945 279 979 313
rect 945 205 979 239
rect 945 131 979 165
rect 945 57 979 91
rect 2869 427 2903 461
rect 2869 353 2903 387
rect 1907 279 1941 313
rect 1907 205 1941 239
rect 1907 131 1941 165
rect 1907 57 1941 91
rect 3831 427 3865 461
rect 3831 353 3865 387
rect 2869 279 2903 313
rect 2869 205 2903 239
rect 2869 131 2903 165
rect 2869 57 2903 91
rect 4793 427 4827 461
rect 4793 353 4827 387
rect 3831 279 3865 313
rect 3831 205 3865 239
rect 3831 131 3865 165
rect 3831 57 3865 91
rect 5755 427 5789 461
rect 5755 353 5789 387
rect 4793 279 4827 313
rect 4793 205 4827 239
rect 4793 131 4827 165
rect 4793 57 4827 91
rect 6717 427 6751 461
rect 6717 353 6751 387
rect 5755 279 5789 313
rect 5755 205 5789 239
rect 5755 131 5789 165
rect 5755 57 5789 91
rect 7679 427 7713 461
rect 7679 353 7713 387
rect 6717 279 6751 313
rect 6717 205 6751 239
rect 6717 131 6751 165
rect 6717 57 6751 91
rect 8641 427 8675 461
rect 8641 353 8675 387
rect 7679 279 7713 313
rect 7679 205 7713 239
rect 7679 131 7713 165
rect 7679 57 7713 91
rect 9603 427 9637 461
rect 9603 353 9637 387
rect 8641 279 8675 313
rect 8641 205 8675 239
rect 8641 131 8675 165
rect 8641 57 8675 91
rect 10565 427 10599 461
rect 10565 353 10599 387
rect 9603 279 9637 313
rect 9603 205 9637 239
rect 9603 131 9637 165
rect 9603 57 9637 91
rect 11527 427 11561 461
rect 11527 353 11561 387
rect 10565 279 10599 313
rect 10565 205 10599 239
rect 10565 131 10599 165
rect 10565 57 10599 91
rect 12489 427 12523 461
rect 12489 353 12523 387
rect 11527 279 11561 313
rect 11527 205 11561 239
rect 11527 131 11561 165
rect 11527 57 11561 91
rect 13451 427 13485 461
rect 13451 353 13485 387
rect 12489 279 12523 313
rect 12489 205 12523 239
rect 12489 131 12523 165
rect 12489 57 12523 91
rect 14413 427 14447 461
rect 14413 353 14447 387
rect 13451 279 13485 313
rect 13451 205 13485 239
rect 13451 131 13485 165
rect 13451 57 13485 91
rect 15375 427 15409 461
rect 15375 353 15409 387
rect 14413 279 14447 313
rect 14413 205 14447 239
rect 14413 131 14447 165
rect 14413 57 14447 91
rect 16337 427 16371 461
rect 16337 353 16371 387
rect 15375 279 15409 313
rect 15375 205 15409 239
rect 15375 131 15409 165
rect 15375 57 15409 91
rect 17299 427 17333 461
rect 17299 353 17333 387
rect 17965 427 17999 461
rect 16337 279 16371 313
rect 16337 205 16371 239
rect 16337 131 16371 165
rect 16337 57 16371 91
rect 17965 353 17999 387
rect 17299 279 17333 313
rect 17299 205 17333 239
rect 17299 131 17333 165
rect 17299 57 17333 91
rect 18631 427 18665 461
rect 18631 353 18665 387
rect 19297 427 19331 461
rect 17965 279 17999 313
rect 17965 205 17999 239
rect 17965 131 17999 165
rect 17965 57 17999 91
rect 19297 353 19331 387
rect 18631 279 18665 313
rect 18631 205 18665 239
rect 18631 131 18665 165
rect 18631 57 18665 91
rect 19297 279 19331 313
rect 19297 205 19331 239
rect 19297 131 19331 165
rect 19297 57 19331 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5163 -17 5197 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5533 -17 5567 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5829 -17 5863 17
rect 5903 -17 5937 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6125 -17 6159 17
rect 6199 -17 6233 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6495 -17 6529 17
rect 6569 -17 6603 17
rect 6643 -17 6677 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7087 -17 7121 17
rect 7161 -17 7195 17
rect 7235 -17 7269 17
rect 7309 -17 7343 17
rect 7383 -17 7417 17
rect 7457 -17 7491 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7753 -17 7787 17
rect 7827 -17 7861 17
rect 7901 -17 7935 17
rect 7975 -17 8009 17
rect 8049 -17 8083 17
rect 8123 -17 8157 17
rect 8197 -17 8231 17
rect 8271 -17 8305 17
rect 8345 -17 8379 17
rect 8419 -17 8453 17
rect 8493 -17 8527 17
rect 8567 -17 8601 17
rect 8715 -17 8749 17
rect 8789 -17 8823 17
rect 8863 -17 8897 17
rect 8937 -17 8971 17
rect 9011 -17 9045 17
rect 9085 -17 9119 17
rect 9159 -17 9193 17
rect 9233 -17 9267 17
rect 9307 -17 9341 17
rect 9381 -17 9415 17
rect 9455 -17 9489 17
rect 9529 -17 9563 17
rect 9677 -17 9711 17
rect 9751 -17 9785 17
rect 9825 -17 9859 17
rect 9899 -17 9933 17
rect 9973 -17 10007 17
rect 10047 -17 10081 17
rect 10121 -17 10155 17
rect 10195 -17 10229 17
rect 10269 -17 10303 17
rect 10343 -17 10377 17
rect 10417 -17 10451 17
rect 10491 -17 10525 17
rect 10639 -17 10673 17
rect 10713 -17 10747 17
rect 10787 -17 10821 17
rect 10861 -17 10895 17
rect 10935 -17 10969 17
rect 11009 -17 11043 17
rect 11083 -17 11117 17
rect 11157 -17 11191 17
rect 11231 -17 11265 17
rect 11305 -17 11339 17
rect 11379 -17 11413 17
rect 11453 -17 11487 17
rect 11601 -17 11635 17
rect 11675 -17 11709 17
rect 11749 -17 11783 17
rect 11823 -17 11857 17
rect 11897 -17 11931 17
rect 11971 -17 12005 17
rect 12045 -17 12079 17
rect 12119 -17 12153 17
rect 12193 -17 12227 17
rect 12267 -17 12301 17
rect 12341 -17 12375 17
rect 12415 -17 12449 17
rect 12563 -17 12597 17
rect 12637 -17 12671 17
rect 12711 -17 12745 17
rect 12785 -17 12819 17
rect 12859 -17 12893 17
rect 12933 -17 12967 17
rect 13007 -17 13041 17
rect 13081 -17 13115 17
rect 13155 -17 13189 17
rect 13229 -17 13263 17
rect 13303 -17 13337 17
rect 13377 -17 13411 17
rect 13525 -17 13559 17
rect 13599 -17 13633 17
rect 13673 -17 13707 17
rect 13747 -17 13781 17
rect 13821 -17 13855 17
rect 13895 -17 13929 17
rect 13969 -17 14003 17
rect 14043 -17 14077 17
rect 14117 -17 14151 17
rect 14191 -17 14225 17
rect 14265 -17 14299 17
rect 14339 -17 14373 17
rect 14487 -17 14521 17
rect 14561 -17 14595 17
rect 14635 -17 14669 17
rect 14709 -17 14743 17
rect 14783 -17 14817 17
rect 14857 -17 14891 17
rect 14931 -17 14965 17
rect 15005 -17 15039 17
rect 15079 -17 15113 17
rect 15153 -17 15187 17
rect 15227 -17 15261 17
rect 15301 -17 15335 17
rect 15449 -17 15483 17
rect 15523 -17 15557 17
rect 15597 -17 15631 17
rect 15671 -17 15705 17
rect 15745 -17 15779 17
rect 15819 -17 15853 17
rect 15893 -17 15927 17
rect 15967 -17 16001 17
rect 16041 -17 16075 17
rect 16115 -17 16149 17
rect 16189 -17 16223 17
rect 16263 -17 16297 17
rect 16411 -17 16445 17
rect 16485 -17 16519 17
rect 16559 -17 16593 17
rect 16633 -17 16667 17
rect 16707 -17 16741 17
rect 16781 -17 16815 17
rect 16855 -17 16889 17
rect 16929 -17 16963 17
rect 17003 -17 17037 17
rect 17077 -17 17111 17
rect 17151 -17 17185 17
rect 17225 -17 17259 17
rect 17373 -17 17407 17
rect 17447 -17 17481 17
rect 17521 -17 17555 17
rect 17595 -17 17629 17
rect 17669 -17 17703 17
rect 17743 -17 17777 17
rect 17817 -17 17851 17
rect 17891 -17 17925 17
rect 18039 -17 18073 17
rect 18113 -17 18147 17
rect 18187 -17 18221 17
rect 18261 -17 18295 17
rect 18335 -17 18369 17
rect 18409 -17 18443 17
rect 18483 -17 18517 17
rect 18557 -17 18591 17
rect 18705 -17 18739 17
rect 18779 -17 18813 17
rect 18853 -17 18887 17
rect 18927 -17 18961 17
rect 19001 -17 19035 17
rect 19075 -17 19109 17
rect 19149 -17 19183 17
rect 19223 -17 19257 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5163 1463 5197 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5533 1463 5567 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5829 1463 5863 1497
rect 5903 1463 5937 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6125 1463 6159 1497
rect 6199 1463 6233 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6495 1463 6529 1497
rect 6569 1463 6603 1497
rect 6643 1463 6677 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7087 1463 7121 1497
rect 7161 1463 7195 1497
rect 7235 1463 7269 1497
rect 7309 1463 7343 1497
rect 7383 1463 7417 1497
rect 7457 1463 7491 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7753 1463 7787 1497
rect 7827 1463 7861 1497
rect 7901 1463 7935 1497
rect 7975 1463 8009 1497
rect 8049 1463 8083 1497
rect 8123 1463 8157 1497
rect 8197 1463 8231 1497
rect 8271 1463 8305 1497
rect 8345 1463 8379 1497
rect 8419 1463 8453 1497
rect 8493 1463 8527 1497
rect 8567 1463 8601 1497
rect 8715 1463 8749 1497
rect 8789 1463 8823 1497
rect 8863 1463 8897 1497
rect 8937 1463 8971 1497
rect 9011 1463 9045 1497
rect 9085 1463 9119 1497
rect 9159 1463 9193 1497
rect 9233 1463 9267 1497
rect 9307 1463 9341 1497
rect 9381 1463 9415 1497
rect 9455 1463 9489 1497
rect 9529 1463 9563 1497
rect 9677 1463 9711 1497
rect 9751 1463 9785 1497
rect 9825 1463 9859 1497
rect 9899 1463 9933 1497
rect 9973 1463 10007 1497
rect 10047 1463 10081 1497
rect 10121 1463 10155 1497
rect 10195 1463 10229 1497
rect 10269 1463 10303 1497
rect 10343 1463 10377 1497
rect 10417 1463 10451 1497
rect 10491 1463 10525 1497
rect 10639 1463 10673 1497
rect 10713 1463 10747 1497
rect 10787 1463 10821 1497
rect 10861 1463 10895 1497
rect 10935 1463 10969 1497
rect 11009 1463 11043 1497
rect 11083 1463 11117 1497
rect 11157 1463 11191 1497
rect 11231 1463 11265 1497
rect 11305 1463 11339 1497
rect 11379 1463 11413 1497
rect 11453 1463 11487 1497
rect 11601 1463 11635 1497
rect 11675 1463 11709 1497
rect 11749 1463 11783 1497
rect 11823 1463 11857 1497
rect 11897 1463 11931 1497
rect 11971 1463 12005 1497
rect 12045 1463 12079 1497
rect 12119 1463 12153 1497
rect 12193 1463 12227 1497
rect 12267 1463 12301 1497
rect 12341 1463 12375 1497
rect 12415 1463 12449 1497
rect 12563 1463 12597 1497
rect 12637 1463 12671 1497
rect 12711 1463 12745 1497
rect 12785 1463 12819 1497
rect 12859 1463 12893 1497
rect 12933 1463 12967 1497
rect 13007 1463 13041 1497
rect 13081 1463 13115 1497
rect 13155 1463 13189 1497
rect 13229 1463 13263 1497
rect 13303 1463 13337 1497
rect 13377 1463 13411 1497
rect 13525 1463 13559 1497
rect 13599 1463 13633 1497
rect 13673 1463 13707 1497
rect 13747 1463 13781 1497
rect 13821 1463 13855 1497
rect 13895 1463 13929 1497
rect 13969 1463 14003 1497
rect 14043 1463 14077 1497
rect 14117 1463 14151 1497
rect 14191 1463 14225 1497
rect 14265 1463 14299 1497
rect 14339 1463 14373 1497
rect 14487 1463 14521 1497
rect 14561 1463 14595 1497
rect 14635 1463 14669 1497
rect 14709 1463 14743 1497
rect 14783 1463 14817 1497
rect 14857 1463 14891 1497
rect 14931 1463 14965 1497
rect 15005 1463 15039 1497
rect 15079 1463 15113 1497
rect 15153 1463 15187 1497
rect 15227 1463 15261 1497
rect 15301 1463 15335 1497
rect 15449 1463 15483 1497
rect 15523 1463 15557 1497
rect 15597 1463 15631 1497
rect 15671 1463 15705 1497
rect 15745 1463 15779 1497
rect 15819 1463 15853 1497
rect 15893 1463 15927 1497
rect 15967 1463 16001 1497
rect 16041 1463 16075 1497
rect 16115 1463 16149 1497
rect 16189 1463 16223 1497
rect 16263 1463 16297 1497
rect 16411 1463 16445 1497
rect 16485 1463 16519 1497
rect 16559 1463 16593 1497
rect 16633 1463 16667 1497
rect 16707 1463 16741 1497
rect 16781 1463 16815 1497
rect 16855 1463 16889 1497
rect 16929 1463 16963 1497
rect 17003 1463 17037 1497
rect 17077 1463 17111 1497
rect 17151 1463 17185 1497
rect 17225 1463 17259 1497
rect 17373 1463 17407 1497
rect 17447 1463 17481 1497
rect 17521 1463 17555 1497
rect 17595 1463 17629 1497
rect 17669 1463 17703 1497
rect 17743 1463 17777 1497
rect 17817 1463 17851 1497
rect 17891 1463 17925 1497
rect 18039 1463 18073 1497
rect 18113 1463 18147 1497
rect 18187 1463 18221 1497
rect 18261 1463 18295 1497
rect 18335 1463 18369 1497
rect 18409 1463 18443 1497
rect 18483 1463 18517 1497
rect 18557 1463 18591 1497
rect 18705 1463 18739 1497
rect 18779 1463 18813 1497
rect 18853 1463 18887 1497
rect 18927 1463 18961 1497
rect 19001 1463 19035 1497
rect 19075 1463 19109 1497
rect 19149 1463 19183 1497
rect 19223 1463 19257 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 945 1389 979 1423
rect 945 1315 979 1349
rect 945 1241 979 1275
rect 945 1167 979 1201
rect 945 1093 979 1127
rect 945 1019 979 1053
rect -17 945 17 979
rect 1907 1389 1941 1423
rect 1907 1315 1941 1349
rect 1907 1241 1941 1275
rect 1907 1167 1941 1201
rect 1907 1093 1941 1127
rect 1907 1019 1941 1053
rect 945 945 979 979
rect -17 871 17 905
rect 2869 1389 2903 1423
rect 2869 1315 2903 1349
rect 2869 1241 2903 1275
rect 2869 1167 2903 1201
rect 2869 1093 2903 1127
rect 2869 1019 2903 1053
rect 1907 945 1941 979
rect 945 871 979 905
rect 3831 1389 3865 1423
rect 3831 1315 3865 1349
rect 3831 1241 3865 1275
rect 3831 1167 3865 1201
rect 3831 1093 3865 1127
rect 3831 1019 3865 1053
rect 2869 945 2903 979
rect 1907 871 1941 905
rect 4793 1389 4827 1423
rect 4793 1315 4827 1349
rect 4793 1241 4827 1275
rect 4793 1167 4827 1201
rect 4793 1093 4827 1127
rect 4793 1019 4827 1053
rect 3831 945 3865 979
rect 2869 871 2903 905
rect 5755 1389 5789 1423
rect 5755 1315 5789 1349
rect 5755 1241 5789 1275
rect 5755 1167 5789 1201
rect 5755 1093 5789 1127
rect 5755 1019 5789 1053
rect 4793 945 4827 979
rect 3831 871 3865 905
rect 6717 1389 6751 1423
rect 6717 1315 6751 1349
rect 6717 1241 6751 1275
rect 6717 1167 6751 1201
rect 6717 1093 6751 1127
rect 6717 1019 6751 1053
rect 5755 945 5789 979
rect 4793 871 4827 905
rect 7679 1389 7713 1423
rect 7679 1315 7713 1349
rect 7679 1241 7713 1275
rect 7679 1167 7713 1201
rect 7679 1093 7713 1127
rect 7679 1019 7713 1053
rect 6717 945 6751 979
rect 5755 871 5789 905
rect 8641 1389 8675 1423
rect 8641 1315 8675 1349
rect 8641 1241 8675 1275
rect 8641 1167 8675 1201
rect 8641 1093 8675 1127
rect 8641 1019 8675 1053
rect 7679 945 7713 979
rect 6717 871 6751 905
rect 9603 1389 9637 1423
rect 9603 1315 9637 1349
rect 9603 1241 9637 1275
rect 9603 1167 9637 1201
rect 9603 1093 9637 1127
rect 9603 1019 9637 1053
rect 8641 945 8675 979
rect 7679 871 7713 905
rect 10565 1389 10599 1423
rect 10565 1315 10599 1349
rect 10565 1241 10599 1275
rect 10565 1167 10599 1201
rect 10565 1093 10599 1127
rect 10565 1019 10599 1053
rect 9603 945 9637 979
rect 8641 871 8675 905
rect 11527 1389 11561 1423
rect 11527 1315 11561 1349
rect 11527 1241 11561 1275
rect 11527 1167 11561 1201
rect 11527 1093 11561 1127
rect 11527 1019 11561 1053
rect 10565 945 10599 979
rect 9603 871 9637 905
rect 12489 1389 12523 1423
rect 12489 1315 12523 1349
rect 12489 1241 12523 1275
rect 12489 1167 12523 1201
rect 12489 1093 12523 1127
rect 12489 1019 12523 1053
rect 11527 945 11561 979
rect 10565 871 10599 905
rect 13451 1389 13485 1423
rect 13451 1315 13485 1349
rect 13451 1241 13485 1275
rect 13451 1167 13485 1201
rect 13451 1093 13485 1127
rect 13451 1019 13485 1053
rect 12489 945 12523 979
rect 11527 871 11561 905
rect 14413 1389 14447 1423
rect 14413 1315 14447 1349
rect 14413 1241 14447 1275
rect 14413 1167 14447 1201
rect 14413 1093 14447 1127
rect 14413 1019 14447 1053
rect 13451 945 13485 979
rect 12489 871 12523 905
rect 15375 1389 15409 1423
rect 15375 1315 15409 1349
rect 15375 1241 15409 1275
rect 15375 1167 15409 1201
rect 15375 1093 15409 1127
rect 15375 1019 15409 1053
rect 14413 945 14447 979
rect 13451 871 13485 905
rect 16337 1389 16371 1423
rect 16337 1315 16371 1349
rect 16337 1241 16371 1275
rect 16337 1167 16371 1201
rect 16337 1093 16371 1127
rect 16337 1019 16371 1053
rect 15375 945 15409 979
rect 14413 871 14447 905
rect 17299 1389 17333 1423
rect 17299 1315 17333 1349
rect 17299 1241 17333 1275
rect 17299 1167 17333 1201
rect 17299 1093 17333 1127
rect 17299 1019 17333 1053
rect 16337 945 16371 979
rect 15375 871 15409 905
rect 17965 1389 17999 1423
rect 17965 1315 17999 1349
rect 17965 1241 17999 1275
rect 17965 1167 17999 1201
rect 17965 1093 17999 1127
rect 17965 1019 17999 1053
rect 17299 945 17333 979
rect 16337 871 16371 905
rect 18631 1389 18665 1423
rect 18631 1315 18665 1349
rect 18631 1241 18665 1275
rect 18631 1167 18665 1201
rect 18631 1093 18665 1127
rect 18631 1019 18665 1053
rect 17965 945 17999 979
rect 17299 871 17333 905
rect 19297 1389 19331 1423
rect 19297 1315 19331 1349
rect 19297 1241 19331 1275
rect 19297 1167 19331 1201
rect 19297 1093 19331 1127
rect 19297 1019 19331 1053
rect 18631 945 18665 979
rect 17965 871 17999 905
rect 19297 945 19331 979
rect 18631 871 18665 905
rect 19297 871 19331 905
<< poly >>
rect 247 1404 277 1430
rect 335 1404 365 1430
rect 423 1404 453 1430
rect 511 1404 541 1430
rect 599 1404 629 1430
rect 687 1404 717 1430
rect 1209 1404 1239 1430
rect 1297 1404 1327 1430
rect 1385 1404 1415 1430
rect 1473 1404 1503 1430
rect 1561 1404 1591 1430
rect 1649 1404 1679 1430
rect 247 973 277 1004
rect 335 973 365 1004
rect 423 973 453 1004
rect 511 973 541 1004
rect 195 957 365 973
rect 195 923 205 957
rect 239 943 365 957
rect 417 957 541 973
rect 239 923 249 943
rect 195 907 249 923
rect 417 923 427 957
rect 461 943 541 957
rect 599 973 629 1004
rect 687 973 717 1004
rect 599 957 717 973
rect 599 943 649 957
rect 461 923 471 943
rect 417 907 471 923
rect 639 923 649 943
rect 683 943 717 957
rect 2171 1404 2201 1430
rect 2259 1404 2289 1430
rect 2347 1404 2377 1430
rect 2435 1404 2465 1430
rect 2523 1404 2553 1430
rect 2611 1404 2641 1430
rect 1209 973 1239 1004
rect 1297 973 1327 1004
rect 1385 973 1415 1004
rect 1473 973 1503 1004
rect 683 923 693 943
rect 639 907 693 923
rect 1157 957 1327 973
rect 1157 923 1167 957
rect 1201 943 1327 957
rect 1379 957 1503 973
rect 1201 923 1211 943
rect 1157 907 1211 923
rect 1379 923 1389 957
rect 1423 943 1503 957
rect 1561 973 1591 1004
rect 1649 973 1679 1004
rect 1561 957 1679 973
rect 1561 943 1611 957
rect 1423 923 1433 943
rect 1379 907 1433 923
rect 1601 923 1611 943
rect 1645 943 1679 957
rect 3133 1404 3163 1430
rect 3221 1404 3251 1430
rect 3309 1404 3339 1430
rect 3397 1404 3427 1430
rect 3485 1404 3515 1430
rect 3573 1404 3603 1430
rect 2171 973 2201 1004
rect 2259 973 2289 1004
rect 2347 973 2377 1004
rect 2435 973 2465 1004
rect 1645 923 1655 943
rect 1601 907 1655 923
rect 2119 957 2289 973
rect 2119 923 2129 957
rect 2163 943 2289 957
rect 2341 957 2465 973
rect 2163 923 2173 943
rect 2119 907 2173 923
rect 2341 923 2351 957
rect 2385 943 2465 957
rect 2523 973 2553 1004
rect 2611 973 2641 1004
rect 2523 957 2641 973
rect 2523 943 2573 957
rect 2385 923 2395 943
rect 2341 907 2395 923
rect 2563 923 2573 943
rect 2607 943 2641 957
rect 4095 1404 4125 1430
rect 4183 1404 4213 1430
rect 4271 1404 4301 1430
rect 4359 1404 4389 1430
rect 4447 1404 4477 1430
rect 4535 1404 4565 1430
rect 3133 973 3163 1004
rect 3221 973 3251 1004
rect 3309 973 3339 1004
rect 3397 973 3427 1004
rect 2607 923 2617 943
rect 2563 907 2617 923
rect 3081 957 3251 973
rect 3081 923 3091 957
rect 3125 943 3251 957
rect 3303 957 3427 973
rect 3125 923 3135 943
rect 3081 907 3135 923
rect 3303 923 3313 957
rect 3347 943 3427 957
rect 3485 973 3515 1004
rect 3573 973 3603 1004
rect 3485 957 3603 973
rect 3485 943 3535 957
rect 3347 923 3357 943
rect 3303 907 3357 923
rect 3525 923 3535 943
rect 3569 943 3603 957
rect 5057 1404 5087 1430
rect 5145 1404 5175 1430
rect 5233 1404 5263 1430
rect 5321 1404 5351 1430
rect 5409 1404 5439 1430
rect 5497 1404 5527 1430
rect 4095 973 4125 1004
rect 4183 973 4213 1004
rect 4271 973 4301 1004
rect 4359 973 4389 1004
rect 3569 923 3579 943
rect 3525 907 3579 923
rect 4043 957 4213 973
rect 4043 923 4053 957
rect 4087 943 4213 957
rect 4265 957 4389 973
rect 4087 923 4097 943
rect 4043 907 4097 923
rect 4265 923 4275 957
rect 4309 943 4389 957
rect 4447 973 4477 1004
rect 4535 973 4565 1004
rect 4447 957 4565 973
rect 4447 943 4497 957
rect 4309 923 4319 943
rect 4265 907 4319 923
rect 4487 923 4497 943
rect 4531 943 4565 957
rect 6019 1404 6049 1430
rect 6107 1404 6137 1430
rect 6195 1404 6225 1430
rect 6283 1404 6313 1430
rect 6371 1404 6401 1430
rect 6459 1404 6489 1430
rect 5057 973 5087 1004
rect 5145 973 5175 1004
rect 5233 973 5263 1004
rect 5321 973 5351 1004
rect 4531 923 4541 943
rect 4487 907 4541 923
rect 5005 957 5175 973
rect 5005 923 5015 957
rect 5049 943 5175 957
rect 5227 957 5351 973
rect 5049 923 5059 943
rect 5005 907 5059 923
rect 5227 923 5237 957
rect 5271 943 5351 957
rect 5409 973 5439 1004
rect 5497 973 5527 1004
rect 5409 957 5527 973
rect 5409 943 5459 957
rect 5271 923 5281 943
rect 5227 907 5281 923
rect 5449 923 5459 943
rect 5493 943 5527 957
rect 6981 1404 7011 1430
rect 7069 1404 7099 1430
rect 7157 1404 7187 1430
rect 7245 1404 7275 1430
rect 7333 1404 7363 1430
rect 7421 1404 7451 1430
rect 6019 973 6049 1004
rect 6107 973 6137 1004
rect 6195 973 6225 1004
rect 6283 973 6313 1004
rect 5493 923 5503 943
rect 5449 907 5503 923
rect 5967 957 6137 973
rect 5967 923 5977 957
rect 6011 943 6137 957
rect 6189 957 6313 973
rect 6011 923 6021 943
rect 5967 907 6021 923
rect 6189 923 6199 957
rect 6233 943 6313 957
rect 6371 973 6401 1004
rect 6459 973 6489 1004
rect 6371 957 6489 973
rect 6371 943 6421 957
rect 6233 923 6243 943
rect 6189 907 6243 923
rect 6411 923 6421 943
rect 6455 943 6489 957
rect 7943 1404 7973 1430
rect 8031 1404 8061 1430
rect 8119 1404 8149 1430
rect 8207 1404 8237 1430
rect 8295 1404 8325 1430
rect 8383 1404 8413 1430
rect 6981 973 7011 1004
rect 7069 973 7099 1004
rect 7157 973 7187 1004
rect 7245 973 7275 1004
rect 6455 923 6465 943
rect 6411 907 6465 923
rect 6929 957 7099 973
rect 6929 923 6939 957
rect 6973 943 7099 957
rect 7151 957 7275 973
rect 6973 923 6983 943
rect 6929 907 6983 923
rect 7151 923 7161 957
rect 7195 943 7275 957
rect 7333 973 7363 1004
rect 7421 973 7451 1004
rect 7333 957 7451 973
rect 7333 943 7383 957
rect 7195 923 7205 943
rect 7151 907 7205 923
rect 7373 923 7383 943
rect 7417 943 7451 957
rect 8905 1404 8935 1430
rect 8993 1404 9023 1430
rect 9081 1404 9111 1430
rect 9169 1404 9199 1430
rect 9257 1404 9287 1430
rect 9345 1404 9375 1430
rect 7943 973 7973 1004
rect 8031 973 8061 1004
rect 8119 973 8149 1004
rect 8207 973 8237 1004
rect 7417 923 7427 943
rect 7373 907 7427 923
rect 7891 957 8061 973
rect 7891 923 7901 957
rect 7935 943 8061 957
rect 8113 957 8237 973
rect 7935 923 7945 943
rect 7891 907 7945 923
rect 8113 923 8123 957
rect 8157 943 8237 957
rect 8295 973 8325 1004
rect 8383 973 8413 1004
rect 8295 957 8413 973
rect 8295 943 8345 957
rect 8157 923 8167 943
rect 8113 907 8167 923
rect 8335 923 8345 943
rect 8379 943 8413 957
rect 9867 1404 9897 1430
rect 9955 1404 9985 1430
rect 10043 1404 10073 1430
rect 10131 1404 10161 1430
rect 10219 1404 10249 1430
rect 10307 1404 10337 1430
rect 8905 973 8935 1004
rect 8993 973 9023 1004
rect 9081 973 9111 1004
rect 9169 973 9199 1004
rect 8379 923 8389 943
rect 8335 907 8389 923
rect 8853 957 9023 973
rect 8853 923 8863 957
rect 8897 943 9023 957
rect 9075 957 9199 973
rect 8897 923 8907 943
rect 8853 907 8907 923
rect 9075 923 9085 957
rect 9119 943 9199 957
rect 9257 973 9287 1004
rect 9345 973 9375 1004
rect 9257 957 9375 973
rect 9257 943 9307 957
rect 9119 923 9129 943
rect 9075 907 9129 923
rect 9297 923 9307 943
rect 9341 943 9375 957
rect 10829 1404 10859 1430
rect 10917 1404 10947 1430
rect 11005 1404 11035 1430
rect 11093 1404 11123 1430
rect 11181 1404 11211 1430
rect 11269 1404 11299 1430
rect 9867 973 9897 1004
rect 9955 973 9985 1004
rect 10043 973 10073 1004
rect 10131 973 10161 1004
rect 9341 923 9351 943
rect 9297 907 9351 923
rect 9815 957 9985 973
rect 9815 923 9825 957
rect 9859 943 9985 957
rect 10037 957 10161 973
rect 9859 923 9869 943
rect 9815 907 9869 923
rect 10037 923 10047 957
rect 10081 943 10161 957
rect 10219 973 10249 1004
rect 10307 973 10337 1004
rect 10219 957 10337 973
rect 10219 943 10269 957
rect 10081 923 10091 943
rect 10037 907 10091 923
rect 10259 923 10269 943
rect 10303 943 10337 957
rect 11791 1404 11821 1430
rect 11879 1404 11909 1430
rect 11967 1404 11997 1430
rect 12055 1404 12085 1430
rect 12143 1404 12173 1430
rect 12231 1404 12261 1430
rect 10829 973 10859 1004
rect 10917 973 10947 1004
rect 11005 973 11035 1004
rect 11093 973 11123 1004
rect 10303 923 10313 943
rect 10259 907 10313 923
rect 10777 957 10947 973
rect 10777 923 10787 957
rect 10821 943 10947 957
rect 10999 957 11123 973
rect 10821 923 10831 943
rect 10777 907 10831 923
rect 10999 923 11009 957
rect 11043 943 11123 957
rect 11181 973 11211 1004
rect 11269 973 11299 1004
rect 11181 957 11299 973
rect 11181 943 11231 957
rect 11043 923 11053 943
rect 10999 907 11053 923
rect 11221 923 11231 943
rect 11265 943 11299 957
rect 12753 1404 12783 1430
rect 12841 1404 12871 1430
rect 12929 1404 12959 1430
rect 13017 1404 13047 1430
rect 13105 1404 13135 1430
rect 13193 1404 13223 1430
rect 11791 973 11821 1004
rect 11879 973 11909 1004
rect 11967 973 11997 1004
rect 12055 973 12085 1004
rect 11265 923 11275 943
rect 11221 907 11275 923
rect 11739 957 11909 973
rect 11739 923 11749 957
rect 11783 943 11909 957
rect 11961 957 12085 973
rect 11783 923 11793 943
rect 11739 907 11793 923
rect 11961 923 11971 957
rect 12005 943 12085 957
rect 12143 973 12173 1004
rect 12231 973 12261 1004
rect 12143 957 12261 973
rect 12143 943 12193 957
rect 12005 923 12015 943
rect 11961 907 12015 923
rect 12183 923 12193 943
rect 12227 943 12261 957
rect 13715 1404 13745 1430
rect 13803 1404 13833 1430
rect 13891 1404 13921 1430
rect 13979 1404 14009 1430
rect 14067 1404 14097 1430
rect 14155 1404 14185 1430
rect 12753 973 12783 1004
rect 12841 973 12871 1004
rect 12929 973 12959 1004
rect 13017 973 13047 1004
rect 12227 923 12237 943
rect 12183 907 12237 923
rect 12701 957 12871 973
rect 12701 923 12711 957
rect 12745 943 12871 957
rect 12923 957 13047 973
rect 12745 923 12755 943
rect 12701 907 12755 923
rect 12923 923 12933 957
rect 12967 943 13047 957
rect 13105 973 13135 1004
rect 13193 973 13223 1004
rect 13105 957 13223 973
rect 13105 943 13155 957
rect 12967 923 12977 943
rect 12923 907 12977 923
rect 13145 923 13155 943
rect 13189 943 13223 957
rect 14677 1404 14707 1430
rect 14765 1404 14795 1430
rect 14853 1404 14883 1430
rect 14941 1404 14971 1430
rect 15029 1404 15059 1430
rect 15117 1404 15147 1430
rect 13715 973 13745 1004
rect 13803 973 13833 1004
rect 13891 973 13921 1004
rect 13979 973 14009 1004
rect 13189 923 13199 943
rect 13145 907 13199 923
rect 13663 957 13833 973
rect 13663 923 13673 957
rect 13707 943 13833 957
rect 13885 957 14009 973
rect 13707 923 13717 943
rect 13663 907 13717 923
rect 13885 923 13895 957
rect 13929 943 14009 957
rect 14067 973 14097 1004
rect 14155 973 14185 1004
rect 14067 957 14185 973
rect 14067 943 14117 957
rect 13929 923 13939 943
rect 13885 907 13939 923
rect 14107 923 14117 943
rect 14151 943 14185 957
rect 15639 1404 15669 1430
rect 15727 1404 15757 1430
rect 15815 1404 15845 1430
rect 15903 1404 15933 1430
rect 15991 1404 16021 1430
rect 16079 1404 16109 1430
rect 14677 973 14707 1004
rect 14765 973 14795 1004
rect 14853 973 14883 1004
rect 14941 973 14971 1004
rect 14151 923 14161 943
rect 14107 907 14161 923
rect 14625 957 14795 973
rect 14625 923 14635 957
rect 14669 943 14795 957
rect 14847 957 14971 973
rect 14669 923 14679 943
rect 14625 907 14679 923
rect 14847 923 14857 957
rect 14891 943 14971 957
rect 15029 973 15059 1004
rect 15117 973 15147 1004
rect 15029 957 15147 973
rect 15029 943 15079 957
rect 14891 923 14901 943
rect 14847 907 14901 923
rect 15069 923 15079 943
rect 15113 943 15147 957
rect 16601 1404 16631 1430
rect 16689 1404 16719 1430
rect 16777 1404 16807 1430
rect 16865 1404 16895 1430
rect 16953 1404 16983 1430
rect 17041 1404 17071 1430
rect 15639 973 15669 1004
rect 15727 973 15757 1004
rect 15815 973 15845 1004
rect 15903 973 15933 1004
rect 15113 923 15123 943
rect 15069 907 15123 923
rect 15587 957 15757 973
rect 15587 923 15597 957
rect 15631 943 15757 957
rect 15809 957 15933 973
rect 15631 923 15641 943
rect 15587 907 15641 923
rect 15809 923 15819 957
rect 15853 943 15933 957
rect 15991 973 16021 1004
rect 16079 973 16109 1004
rect 15991 957 16109 973
rect 15991 943 16041 957
rect 15853 923 15863 943
rect 15809 907 15863 923
rect 16031 923 16041 943
rect 16075 943 16109 957
rect 17503 1405 17533 1431
rect 17591 1405 17621 1431
rect 17679 1405 17709 1431
rect 17767 1405 17797 1431
rect 16601 973 16631 1004
rect 16689 973 16719 1004
rect 16777 973 16807 1004
rect 16865 973 16895 1004
rect 16075 923 16085 943
rect 16031 907 16085 923
rect 16549 957 16719 973
rect 16549 923 16559 957
rect 16593 943 16719 957
rect 16771 957 16895 973
rect 16593 923 16603 943
rect 16549 907 16603 923
rect 16771 923 16781 957
rect 16815 943 16895 957
rect 16953 973 16983 1004
rect 17041 973 17071 1004
rect 16953 957 17071 973
rect 16953 943 17003 957
rect 16815 923 16825 943
rect 16771 907 16825 923
rect 16993 923 17003 943
rect 17037 943 17071 957
rect 18167 1405 18197 1431
rect 18255 1405 18285 1431
rect 18343 1405 18373 1431
rect 18431 1405 18461 1431
rect 17503 974 17533 1005
rect 17591 974 17621 1005
rect 17679 974 17709 1005
rect 17767 974 17797 1005
rect 17037 923 17047 943
rect 16993 907 17047 923
rect 17437 958 17621 974
rect 17437 924 17447 958
rect 17481 944 17621 958
rect 17667 958 17797 974
rect 17481 924 17491 944
rect 17437 908 17491 924
rect 17667 924 17677 958
rect 17711 944 17797 958
rect 18835 1405 18865 1431
rect 18923 1405 18953 1431
rect 19011 1405 19041 1431
rect 19099 1405 19129 1431
rect 17711 924 17721 944
rect 17667 908 17721 924
rect 18167 974 18197 1005
rect 18255 974 18285 1005
rect 18167 958 18285 974
rect 18167 944 18187 958
rect 18177 924 18187 944
rect 18221 944 18285 958
rect 18343 974 18373 1005
rect 18431 974 18461 1005
rect 18343 958 18527 974
rect 18343 944 18483 958
rect 18221 924 18231 944
rect 18177 908 18231 924
rect 18473 924 18483 944
rect 18517 924 18527 958
rect 18473 908 18527 924
rect 18835 974 18865 1005
rect 18923 974 18953 1005
rect 19011 974 19041 1005
rect 19099 974 19129 1005
rect 18769 958 18953 974
rect 18769 924 18779 958
rect 18813 944 18953 958
rect 18995 958 19129 974
rect 18813 924 18823 944
rect 18769 908 18823 924
rect 18995 924 19005 958
rect 19039 944 19129 958
rect 19039 924 19049 944
rect 18995 908 19049 924
rect 195 433 249 449
rect 195 413 205 433
rect 147 399 205 413
rect 239 399 249 433
rect 147 383 249 399
rect 417 433 471 449
rect 417 399 427 433
rect 461 413 471 433
rect 639 433 693 449
rect 461 399 477 413
rect 417 383 477 399
rect 639 399 649 433
rect 683 399 693 433
rect 639 383 693 399
rect 1157 433 1211 449
rect 1157 413 1167 433
rect 147 351 177 383
rect 447 351 477 383
rect 649 351 679 383
rect 1109 399 1167 413
rect 1201 399 1211 433
rect 1109 383 1211 399
rect 1379 433 1433 449
rect 1379 399 1389 433
rect 1423 413 1433 433
rect 1601 433 1655 449
rect 1423 399 1439 413
rect 1379 383 1439 399
rect 1601 399 1611 433
rect 1645 399 1655 433
rect 1601 383 1655 399
rect 2119 433 2173 449
rect 2119 413 2129 433
rect 1109 351 1139 383
rect 1409 351 1439 383
rect 1611 351 1641 383
rect 2071 399 2129 413
rect 2163 399 2173 433
rect 2071 383 2173 399
rect 2341 433 2395 449
rect 2341 399 2351 433
rect 2385 413 2395 433
rect 2563 433 2617 449
rect 2385 399 2401 413
rect 2341 383 2401 399
rect 2563 399 2573 433
rect 2607 399 2617 433
rect 2563 383 2617 399
rect 3081 433 3135 449
rect 3081 413 3091 433
rect 2071 351 2101 383
rect 2371 351 2401 383
rect 2573 351 2603 383
rect 3033 399 3091 413
rect 3125 399 3135 433
rect 3033 383 3135 399
rect 3303 433 3357 449
rect 3303 399 3313 433
rect 3347 413 3357 433
rect 3525 433 3579 449
rect 3347 399 3363 413
rect 3303 383 3363 399
rect 3525 399 3535 433
rect 3569 399 3579 433
rect 3525 383 3579 399
rect 4043 433 4097 449
rect 4043 413 4053 433
rect 3033 351 3063 383
rect 3333 351 3363 383
rect 3535 351 3565 383
rect 3995 399 4053 413
rect 4087 399 4097 433
rect 3995 383 4097 399
rect 4265 433 4319 449
rect 4265 399 4275 433
rect 4309 413 4319 433
rect 4487 433 4541 449
rect 4309 399 4325 413
rect 4265 383 4325 399
rect 4487 399 4497 433
rect 4531 399 4541 433
rect 4487 383 4541 399
rect 5005 433 5059 449
rect 5005 413 5015 433
rect 3995 351 4025 383
rect 4295 351 4325 383
rect 4497 351 4527 383
rect 4957 399 5015 413
rect 5049 399 5059 433
rect 4957 383 5059 399
rect 5227 433 5281 449
rect 5227 399 5237 433
rect 5271 413 5281 433
rect 5449 433 5503 449
rect 5271 399 5287 413
rect 5227 383 5287 399
rect 5449 399 5459 433
rect 5493 399 5503 433
rect 5449 383 5503 399
rect 5967 433 6021 449
rect 5967 413 5977 433
rect 4957 351 4987 383
rect 5257 351 5287 383
rect 5459 351 5489 383
rect 5919 399 5977 413
rect 6011 399 6021 433
rect 5919 383 6021 399
rect 6189 433 6243 449
rect 6189 399 6199 433
rect 6233 413 6243 433
rect 6411 433 6465 449
rect 6233 399 6249 413
rect 6189 383 6249 399
rect 6411 399 6421 433
rect 6455 399 6465 433
rect 6411 383 6465 399
rect 6929 433 6983 449
rect 6929 413 6939 433
rect 5919 351 5949 383
rect 6219 351 6249 383
rect 6421 351 6451 383
rect 6881 399 6939 413
rect 6973 399 6983 433
rect 6881 383 6983 399
rect 7151 433 7205 449
rect 7151 399 7161 433
rect 7195 413 7205 433
rect 7373 433 7427 449
rect 7195 399 7211 413
rect 7151 383 7211 399
rect 7373 399 7383 433
rect 7417 399 7427 433
rect 7373 383 7427 399
rect 7891 433 7945 449
rect 7891 413 7901 433
rect 6881 351 6911 383
rect 7181 351 7211 383
rect 7383 351 7413 383
rect 7843 399 7901 413
rect 7935 399 7945 433
rect 7843 383 7945 399
rect 8113 433 8167 449
rect 8113 399 8123 433
rect 8157 413 8167 433
rect 8335 433 8389 449
rect 8157 399 8173 413
rect 8113 383 8173 399
rect 8335 399 8345 433
rect 8379 399 8389 433
rect 8335 383 8389 399
rect 8853 433 8907 449
rect 8853 413 8863 433
rect 7843 351 7873 383
rect 8143 351 8173 383
rect 8345 351 8375 383
rect 8805 399 8863 413
rect 8897 399 8907 433
rect 8805 383 8907 399
rect 9075 433 9129 449
rect 9075 399 9085 433
rect 9119 413 9129 433
rect 9297 433 9351 449
rect 9119 399 9135 413
rect 9075 383 9135 399
rect 9297 399 9307 433
rect 9341 399 9351 433
rect 9297 383 9351 399
rect 9815 433 9869 449
rect 9815 413 9825 433
rect 8805 351 8835 383
rect 9105 351 9135 383
rect 9307 351 9337 383
rect 9767 399 9825 413
rect 9859 399 9869 433
rect 9767 383 9869 399
rect 10037 433 10091 449
rect 10037 399 10047 433
rect 10081 413 10091 433
rect 10259 433 10313 449
rect 10081 399 10097 413
rect 10037 383 10097 399
rect 10259 399 10269 433
rect 10303 399 10313 433
rect 10259 383 10313 399
rect 10777 433 10831 449
rect 10777 413 10787 433
rect 9767 351 9797 383
rect 10067 351 10097 383
rect 10269 351 10299 383
rect 10729 399 10787 413
rect 10821 399 10831 433
rect 10729 383 10831 399
rect 10999 433 11053 449
rect 10999 399 11009 433
rect 11043 413 11053 433
rect 11221 433 11275 449
rect 11043 399 11059 413
rect 10999 383 11059 399
rect 11221 399 11231 433
rect 11265 399 11275 433
rect 11221 383 11275 399
rect 11739 433 11793 449
rect 11739 413 11749 433
rect 10729 351 10759 383
rect 11029 351 11059 383
rect 11231 351 11261 383
rect 11691 399 11749 413
rect 11783 399 11793 433
rect 11691 383 11793 399
rect 11961 433 12015 449
rect 11961 399 11971 433
rect 12005 413 12015 433
rect 12183 433 12237 449
rect 12005 399 12021 413
rect 11961 383 12021 399
rect 12183 399 12193 433
rect 12227 399 12237 433
rect 12183 383 12237 399
rect 12701 433 12755 449
rect 12701 413 12711 433
rect 11691 351 11721 383
rect 11991 351 12021 383
rect 12193 351 12223 383
rect 12653 399 12711 413
rect 12745 399 12755 433
rect 12653 383 12755 399
rect 12923 433 12977 449
rect 12923 399 12933 433
rect 12967 413 12977 433
rect 13145 433 13199 449
rect 12967 399 12983 413
rect 12923 383 12983 399
rect 13145 399 13155 433
rect 13189 399 13199 433
rect 13145 383 13199 399
rect 13663 433 13717 449
rect 13663 413 13673 433
rect 12653 351 12683 383
rect 12953 351 12983 383
rect 13155 351 13185 383
rect 13615 399 13673 413
rect 13707 399 13717 433
rect 13615 383 13717 399
rect 13885 433 13939 449
rect 13885 399 13895 433
rect 13929 413 13939 433
rect 14107 433 14161 449
rect 13929 399 13945 413
rect 13885 383 13945 399
rect 14107 399 14117 433
rect 14151 399 14161 433
rect 14107 383 14161 399
rect 14625 433 14679 449
rect 14625 413 14635 433
rect 13615 351 13645 383
rect 13915 351 13945 383
rect 14117 351 14147 383
rect 14577 399 14635 413
rect 14669 399 14679 433
rect 14577 383 14679 399
rect 14847 433 14901 449
rect 14847 399 14857 433
rect 14891 413 14901 433
rect 15069 433 15123 449
rect 14891 399 14907 413
rect 14847 383 14907 399
rect 15069 399 15079 433
rect 15113 399 15123 433
rect 15069 383 15123 399
rect 15587 433 15641 449
rect 15587 413 15597 433
rect 14577 351 14607 383
rect 14877 351 14907 383
rect 15079 351 15109 383
rect 15539 399 15597 413
rect 15631 399 15641 433
rect 15539 383 15641 399
rect 15809 433 15863 449
rect 15809 399 15819 433
rect 15853 413 15863 433
rect 16031 433 16085 449
rect 15853 399 15869 413
rect 15809 383 15869 399
rect 16031 399 16041 433
rect 16075 399 16085 433
rect 16031 383 16085 399
rect 16549 433 16603 449
rect 16549 413 16559 433
rect 15539 351 15569 383
rect 15839 351 15869 383
rect 16041 351 16071 383
rect 16501 399 16559 413
rect 16593 399 16603 433
rect 16501 383 16603 399
rect 16771 433 16825 449
rect 16771 399 16781 433
rect 16815 413 16825 433
rect 16993 433 17047 449
rect 16815 399 16831 413
rect 16771 383 16831 399
rect 16993 399 17003 433
rect 17037 399 17047 433
rect 16993 383 17047 399
rect 16501 351 16531 383
rect 16801 351 16831 383
rect 17003 351 17033 383
rect 17437 433 17491 449
rect 17437 399 17447 433
rect 17481 413 17491 433
rect 17659 433 17713 449
rect 17481 399 17514 413
rect 17437 383 17514 399
rect 17659 399 17669 433
rect 17703 399 17713 433
rect 17659 383 17713 399
rect 18177 433 18231 449
rect 18177 413 18187 433
rect 17484 349 17514 383
rect 17678 349 17708 383
rect 18150 399 18187 413
rect 18221 399 18231 433
rect 18473 433 18527 449
rect 18473 413 18483 433
rect 18150 383 18231 399
rect 18450 399 18483 413
rect 18517 399 18527 433
rect 18450 383 18527 399
rect 18150 349 18180 383
rect 18450 349 18480 383
rect 18769 433 18823 449
rect 18769 399 18779 433
rect 18813 413 18823 433
rect 18991 433 19045 449
rect 18813 399 18846 413
rect 18769 383 18846 399
rect 18991 399 19001 433
rect 19035 399 19045 433
rect 18991 383 19045 399
rect 18816 349 18846 383
rect 19010 349 19040 383
<< polycont >>
rect 205 923 239 957
rect 427 923 461 957
rect 649 923 683 957
rect 1167 923 1201 957
rect 1389 923 1423 957
rect 1611 923 1645 957
rect 2129 923 2163 957
rect 2351 923 2385 957
rect 2573 923 2607 957
rect 3091 923 3125 957
rect 3313 923 3347 957
rect 3535 923 3569 957
rect 4053 923 4087 957
rect 4275 923 4309 957
rect 4497 923 4531 957
rect 5015 923 5049 957
rect 5237 923 5271 957
rect 5459 923 5493 957
rect 5977 923 6011 957
rect 6199 923 6233 957
rect 6421 923 6455 957
rect 6939 923 6973 957
rect 7161 923 7195 957
rect 7383 923 7417 957
rect 7901 923 7935 957
rect 8123 923 8157 957
rect 8345 923 8379 957
rect 8863 923 8897 957
rect 9085 923 9119 957
rect 9307 923 9341 957
rect 9825 923 9859 957
rect 10047 923 10081 957
rect 10269 923 10303 957
rect 10787 923 10821 957
rect 11009 923 11043 957
rect 11231 923 11265 957
rect 11749 923 11783 957
rect 11971 923 12005 957
rect 12193 923 12227 957
rect 12711 923 12745 957
rect 12933 923 12967 957
rect 13155 923 13189 957
rect 13673 923 13707 957
rect 13895 923 13929 957
rect 14117 923 14151 957
rect 14635 923 14669 957
rect 14857 923 14891 957
rect 15079 923 15113 957
rect 15597 923 15631 957
rect 15819 923 15853 957
rect 16041 923 16075 957
rect 16559 923 16593 957
rect 16781 923 16815 957
rect 17003 923 17037 957
rect 17447 924 17481 958
rect 17677 924 17711 958
rect 18187 924 18221 958
rect 18483 924 18517 958
rect 18779 924 18813 958
rect 19005 924 19039 958
rect 205 399 239 433
rect 427 399 461 433
rect 649 399 683 433
rect 1167 399 1201 433
rect 1389 399 1423 433
rect 1611 399 1645 433
rect 2129 399 2163 433
rect 2351 399 2385 433
rect 2573 399 2607 433
rect 3091 399 3125 433
rect 3313 399 3347 433
rect 3535 399 3569 433
rect 4053 399 4087 433
rect 4275 399 4309 433
rect 4497 399 4531 433
rect 5015 399 5049 433
rect 5237 399 5271 433
rect 5459 399 5493 433
rect 5977 399 6011 433
rect 6199 399 6233 433
rect 6421 399 6455 433
rect 6939 399 6973 433
rect 7161 399 7195 433
rect 7383 399 7417 433
rect 7901 399 7935 433
rect 8123 399 8157 433
rect 8345 399 8379 433
rect 8863 399 8897 433
rect 9085 399 9119 433
rect 9307 399 9341 433
rect 9825 399 9859 433
rect 10047 399 10081 433
rect 10269 399 10303 433
rect 10787 399 10821 433
rect 11009 399 11043 433
rect 11231 399 11265 433
rect 11749 399 11783 433
rect 11971 399 12005 433
rect 12193 399 12227 433
rect 12711 399 12745 433
rect 12933 399 12967 433
rect 13155 399 13189 433
rect 13673 399 13707 433
rect 13895 399 13929 433
rect 14117 399 14151 433
rect 14635 399 14669 433
rect 14857 399 14891 433
rect 15079 399 15113 433
rect 15597 399 15631 433
rect 15819 399 15853 433
rect 16041 399 16075 433
rect 16559 399 16593 433
rect 16781 399 16815 433
rect 17003 399 17037 433
rect 17447 399 17481 433
rect 17669 399 17703 433
rect 18187 399 18221 433
rect 18483 399 18517 433
rect 18779 399 18813 433
rect 19001 399 19035 433
<< locali >>
rect -34 1497 19348 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6569 1497
rect 6603 1463 6643 1497
rect 6677 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7753 1497
rect 7787 1463 7827 1497
rect 7861 1463 7901 1497
rect 7935 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8123 1497
rect 8157 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8567 1497
rect 8601 1463 8715 1497
rect 8749 1463 8789 1497
rect 8823 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9529 1497
rect 9563 1463 9677 1497
rect 9711 1463 9751 1497
rect 9785 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10195 1497
rect 10229 1463 10269 1497
rect 10303 1463 10343 1497
rect 10377 1463 10417 1497
rect 10451 1463 10491 1497
rect 10525 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10861 1497
rect 10895 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11305 1497
rect 11339 1463 11379 1497
rect 11413 1463 11453 1497
rect 11487 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12193 1497
rect 12227 1463 12267 1497
rect 12301 1463 12341 1497
rect 12375 1463 12415 1497
rect 12449 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12859 1497
rect 12893 1463 12933 1497
rect 12967 1463 13007 1497
rect 13041 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13525 1497
rect 13559 1463 13599 1497
rect 13633 1463 13673 1497
rect 13707 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13895 1497
rect 13929 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14191 1497
rect 14225 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14635 1497
rect 14669 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14857 1497
rect 14891 1463 14931 1497
rect 14965 1463 15005 1497
rect 15039 1463 15079 1497
rect 15113 1463 15153 1497
rect 15187 1463 15227 1497
rect 15261 1463 15301 1497
rect 15335 1463 15449 1497
rect 15483 1463 15523 1497
rect 15557 1463 15597 1497
rect 15631 1463 15671 1497
rect 15705 1463 15745 1497
rect 15779 1463 15819 1497
rect 15853 1463 15893 1497
rect 15927 1463 15967 1497
rect 16001 1463 16041 1497
rect 16075 1463 16115 1497
rect 16149 1463 16189 1497
rect 16223 1463 16263 1497
rect 16297 1463 16411 1497
rect 16445 1463 16485 1497
rect 16519 1463 16559 1497
rect 16593 1463 16633 1497
rect 16667 1463 16707 1497
rect 16741 1463 16781 1497
rect 16815 1463 16855 1497
rect 16889 1463 16929 1497
rect 16963 1463 17003 1497
rect 17037 1463 17077 1497
rect 17111 1463 17151 1497
rect 17185 1463 17225 1497
rect 17259 1463 17373 1497
rect 17407 1463 17447 1497
rect 17481 1463 17521 1497
rect 17555 1463 17595 1497
rect 17629 1463 17669 1497
rect 17703 1463 17743 1497
rect 17777 1463 17817 1497
rect 17851 1463 17891 1497
rect 17925 1463 18039 1497
rect 18073 1463 18113 1497
rect 18147 1463 18187 1497
rect 18221 1463 18261 1497
rect 18295 1463 18335 1497
rect 18369 1463 18409 1497
rect 18443 1463 18483 1497
rect 18517 1463 18557 1497
rect 18591 1463 18705 1497
rect 18739 1463 18779 1497
rect 18813 1463 18853 1497
rect 18887 1463 18927 1497
rect 18961 1463 19001 1497
rect 19035 1463 19075 1497
rect 19109 1463 19149 1497
rect 19183 1463 19223 1497
rect 19257 1463 19348 1497
rect -34 1446 19348 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 201 1366 235 1446
rect 201 1298 235 1332
rect 201 1230 235 1264
rect 201 1162 235 1196
rect 201 1093 235 1128
rect 201 1043 235 1059
rect 289 1366 323 1404
rect 289 1298 323 1332
rect 289 1230 323 1264
rect 289 1162 323 1196
rect 289 1093 323 1128
rect 377 1366 411 1446
rect 377 1298 411 1332
rect 377 1230 411 1264
rect 377 1162 411 1196
rect 377 1111 411 1128
rect 465 1366 499 1404
rect 465 1298 499 1332
rect 465 1230 499 1264
rect 465 1162 499 1196
rect 289 1048 323 1059
rect 465 1093 499 1128
rect 553 1366 587 1446
rect 553 1298 587 1332
rect 553 1230 587 1264
rect 553 1162 587 1196
rect 553 1111 587 1128
rect 641 1366 675 1404
rect 641 1298 675 1332
rect 641 1230 675 1264
rect 641 1162 675 1196
rect 465 1048 499 1059
rect 641 1093 675 1128
rect 729 1366 763 1446
rect 729 1298 763 1332
rect 729 1230 763 1264
rect 729 1162 763 1196
rect 729 1111 763 1128
rect 928 1423 996 1446
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 641 1048 675 1059
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect -34 979 34 1019
rect 289 1014 831 1048
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 205 831 239 923
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 797
rect 205 383 239 399
rect 427 957 461 973
rect 427 461 461 923
rect 427 383 461 399
rect 649 957 683 973
rect 649 683 683 923
rect 649 433 683 649
rect 649 383 683 399
rect 797 535 831 1014
rect 928 1019 945 1053
rect 979 1019 996 1053
rect 1163 1366 1197 1446
rect 1163 1298 1197 1332
rect 1163 1230 1197 1264
rect 1163 1162 1197 1196
rect 1163 1093 1197 1128
rect 1163 1043 1197 1059
rect 1251 1366 1285 1404
rect 1251 1298 1285 1332
rect 1251 1230 1285 1264
rect 1251 1162 1285 1196
rect 1251 1093 1285 1128
rect 1339 1366 1373 1446
rect 1339 1298 1373 1332
rect 1339 1230 1373 1264
rect 1339 1162 1373 1196
rect 1339 1111 1373 1128
rect 1427 1366 1461 1404
rect 1427 1298 1461 1332
rect 1427 1230 1461 1264
rect 1427 1162 1461 1196
rect 1251 1048 1285 1059
rect 1427 1093 1461 1128
rect 1515 1366 1549 1446
rect 1515 1298 1549 1332
rect 1515 1230 1549 1264
rect 1515 1162 1549 1196
rect 1515 1111 1549 1128
rect 1603 1366 1637 1404
rect 1603 1298 1637 1332
rect 1603 1230 1637 1264
rect 1603 1162 1637 1196
rect 1427 1048 1461 1059
rect 1603 1093 1637 1128
rect 1691 1366 1725 1446
rect 1691 1298 1725 1332
rect 1691 1230 1725 1264
rect 1691 1162 1725 1196
rect 1691 1111 1725 1128
rect 1890 1423 1958 1446
rect 1890 1389 1907 1423
rect 1941 1389 1958 1423
rect 1890 1349 1958 1389
rect 1890 1315 1907 1349
rect 1941 1315 1958 1349
rect 1890 1275 1958 1315
rect 1890 1241 1907 1275
rect 1941 1241 1958 1275
rect 1890 1201 1958 1241
rect 1890 1167 1907 1201
rect 1941 1167 1958 1201
rect 1890 1127 1958 1167
rect 1603 1048 1637 1059
rect 1890 1093 1907 1127
rect 1941 1093 1958 1127
rect 1890 1053 1958 1093
rect 928 979 996 1019
rect 1251 1014 1793 1048
rect 928 945 945 979
rect 979 945 996 979
rect 928 905 996 945
rect 928 871 945 905
rect 979 871 996 905
rect 928 822 996 871
rect 1167 957 1201 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 101 335 135 351
rect 295 335 329 351
rect 489 335 523 351
rect 135 301 198 335
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 489 335
rect 101 263 135 301
rect 101 195 135 229
rect 295 263 329 301
rect 489 285 523 301
rect 603 335 637 351
rect 797 350 831 501
rect 603 263 637 301
rect 101 125 135 161
rect 101 75 135 91
rect 198 210 232 226
rect -34 34 34 57
rect 198 34 232 176
rect 295 195 329 229
rect 393 216 427 232
rect 603 216 637 229
rect 427 195 637 216
rect 427 182 603 195
rect 393 166 427 182
rect 295 125 329 161
rect 700 316 831 350
rect 928 461 996 544
rect 928 427 945 461
rect 979 427 996 461
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect 1167 535 1201 923
rect 1167 433 1201 501
rect 1167 383 1201 399
rect 1389 957 1423 973
rect 1389 905 1423 923
rect 1389 433 1423 871
rect 1389 383 1423 399
rect 1611 957 1645 973
rect 1611 757 1645 923
rect 1611 433 1645 723
rect 1611 383 1645 399
rect 1759 683 1793 1014
rect 1890 1019 1907 1053
rect 1941 1019 1958 1053
rect 2125 1366 2159 1446
rect 2125 1298 2159 1332
rect 2125 1230 2159 1264
rect 2125 1162 2159 1196
rect 2125 1093 2159 1128
rect 2125 1043 2159 1059
rect 2213 1366 2247 1404
rect 2213 1298 2247 1332
rect 2213 1230 2247 1264
rect 2213 1162 2247 1196
rect 2213 1093 2247 1128
rect 2301 1366 2335 1446
rect 2301 1298 2335 1332
rect 2301 1230 2335 1264
rect 2301 1162 2335 1196
rect 2301 1111 2335 1128
rect 2389 1366 2423 1404
rect 2389 1298 2423 1332
rect 2389 1230 2423 1264
rect 2389 1162 2423 1196
rect 2213 1048 2247 1059
rect 2389 1093 2423 1128
rect 2477 1366 2511 1446
rect 2477 1298 2511 1332
rect 2477 1230 2511 1264
rect 2477 1162 2511 1196
rect 2477 1111 2511 1128
rect 2565 1366 2599 1404
rect 2565 1298 2599 1332
rect 2565 1230 2599 1264
rect 2565 1162 2599 1196
rect 2389 1048 2423 1059
rect 2565 1093 2599 1128
rect 2653 1366 2687 1446
rect 2653 1298 2687 1332
rect 2653 1230 2687 1264
rect 2653 1162 2687 1196
rect 2653 1111 2687 1128
rect 2852 1423 2920 1446
rect 2852 1389 2869 1423
rect 2903 1389 2920 1423
rect 2852 1349 2920 1389
rect 2852 1315 2869 1349
rect 2903 1315 2920 1349
rect 2852 1275 2920 1315
rect 2852 1241 2869 1275
rect 2903 1241 2920 1275
rect 2852 1201 2920 1241
rect 2852 1167 2869 1201
rect 2903 1167 2920 1201
rect 2852 1127 2920 1167
rect 2565 1048 2599 1059
rect 2852 1093 2869 1127
rect 2903 1093 2920 1127
rect 2852 1053 2920 1093
rect 1890 979 1958 1019
rect 2213 1014 2755 1048
rect 1890 945 1907 979
rect 1941 945 1958 979
rect 1890 905 1958 945
rect 1890 871 1907 905
rect 1941 871 1958 905
rect 1890 822 1958 871
rect 2129 957 2163 973
rect 700 219 734 316
rect 928 313 996 353
rect 928 279 945 313
rect 979 279 996 313
rect 700 169 734 185
rect 797 263 831 279
rect 797 195 831 229
rect 489 125 523 141
rect 329 91 392 125
rect 426 91 489 125
rect 295 75 329 91
rect 489 75 523 91
rect 603 125 637 161
rect 797 125 831 161
rect 637 91 700 125
rect 734 91 797 125
rect 603 75 637 91
rect 797 75 831 91
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect 928 57 945 91
rect 979 57 996 91
rect 1063 335 1097 351
rect 1257 335 1291 351
rect 1451 335 1485 351
rect 1097 301 1160 335
rect 1194 301 1257 335
rect 1291 301 1354 335
rect 1388 301 1451 335
rect 1063 263 1097 301
rect 1063 195 1097 229
rect 1257 263 1291 301
rect 1451 285 1485 301
rect 1565 335 1599 351
rect 1759 350 1793 649
rect 1565 263 1599 301
rect 1063 125 1097 161
rect 1063 75 1097 91
rect 1160 210 1194 226
rect 928 34 996 57
rect 1160 34 1194 176
rect 1257 195 1291 229
rect 1355 216 1389 232
rect 1565 216 1599 229
rect 1389 195 1599 216
rect 1389 182 1565 195
rect 1355 166 1389 182
rect 1257 125 1291 161
rect 1662 316 1793 350
rect 1890 461 1958 544
rect 1890 427 1907 461
rect 1941 427 1958 461
rect 1890 387 1958 427
rect 1890 353 1907 387
rect 1941 353 1958 387
rect 2129 535 2163 923
rect 2129 433 2163 501
rect 2129 383 2163 399
rect 2351 957 2385 973
rect 2351 609 2385 923
rect 2351 433 2385 575
rect 2351 383 2385 399
rect 2573 957 2607 973
rect 2573 757 2607 923
rect 2573 433 2607 723
rect 2573 383 2607 399
rect 2721 535 2755 1014
rect 2852 1019 2869 1053
rect 2903 1019 2920 1053
rect 3087 1366 3121 1446
rect 3087 1298 3121 1332
rect 3087 1230 3121 1264
rect 3087 1162 3121 1196
rect 3087 1093 3121 1128
rect 3087 1043 3121 1059
rect 3175 1366 3209 1404
rect 3175 1298 3209 1332
rect 3175 1230 3209 1264
rect 3175 1162 3209 1196
rect 3175 1093 3209 1128
rect 3263 1366 3297 1446
rect 3263 1298 3297 1332
rect 3263 1230 3297 1264
rect 3263 1162 3297 1196
rect 3263 1111 3297 1128
rect 3351 1366 3385 1404
rect 3351 1298 3385 1332
rect 3351 1230 3385 1264
rect 3351 1162 3385 1196
rect 3175 1048 3209 1059
rect 3351 1093 3385 1128
rect 3439 1366 3473 1446
rect 3439 1298 3473 1332
rect 3439 1230 3473 1264
rect 3439 1162 3473 1196
rect 3439 1111 3473 1128
rect 3527 1366 3561 1404
rect 3527 1298 3561 1332
rect 3527 1230 3561 1264
rect 3527 1162 3561 1196
rect 3351 1048 3385 1059
rect 3527 1093 3561 1128
rect 3615 1366 3649 1446
rect 3615 1298 3649 1332
rect 3615 1230 3649 1264
rect 3615 1162 3649 1196
rect 3615 1111 3649 1128
rect 3814 1423 3882 1446
rect 3814 1389 3831 1423
rect 3865 1389 3882 1423
rect 3814 1349 3882 1389
rect 3814 1315 3831 1349
rect 3865 1315 3882 1349
rect 3814 1275 3882 1315
rect 3814 1241 3831 1275
rect 3865 1241 3882 1275
rect 3814 1201 3882 1241
rect 3814 1167 3831 1201
rect 3865 1167 3882 1201
rect 3814 1127 3882 1167
rect 3527 1048 3561 1059
rect 3814 1093 3831 1127
rect 3865 1093 3882 1127
rect 3814 1053 3882 1093
rect 2852 979 2920 1019
rect 3175 1014 3717 1048
rect 2852 945 2869 979
rect 2903 945 2920 979
rect 2852 905 2920 945
rect 2852 871 2869 905
rect 2903 871 2920 905
rect 2852 822 2920 871
rect 3091 957 3125 973
rect 1662 219 1696 316
rect 1890 313 1958 353
rect 1890 279 1907 313
rect 1941 279 1958 313
rect 1662 169 1696 185
rect 1759 263 1793 279
rect 1759 195 1793 229
rect 1451 125 1485 141
rect 1291 91 1354 125
rect 1388 91 1451 125
rect 1257 75 1291 91
rect 1451 75 1485 91
rect 1565 125 1599 161
rect 1759 125 1793 161
rect 1599 91 1662 125
rect 1696 91 1759 125
rect 1565 75 1599 91
rect 1759 75 1793 91
rect 1890 239 1958 279
rect 1890 205 1907 239
rect 1941 205 1958 239
rect 1890 165 1958 205
rect 1890 131 1907 165
rect 1941 131 1958 165
rect 1890 91 1958 131
rect 1890 57 1907 91
rect 1941 57 1958 91
rect 2025 335 2059 351
rect 2219 335 2253 351
rect 2413 335 2447 351
rect 2059 301 2122 335
rect 2156 301 2219 335
rect 2253 301 2316 335
rect 2350 301 2413 335
rect 2025 263 2059 301
rect 2025 195 2059 229
rect 2219 263 2253 301
rect 2413 285 2447 301
rect 2527 335 2561 351
rect 2721 350 2755 501
rect 2527 263 2561 301
rect 2025 125 2059 161
rect 2025 75 2059 91
rect 2122 210 2156 226
rect 1890 34 1958 57
rect 2122 34 2156 176
rect 2219 195 2253 229
rect 2317 216 2351 232
rect 2527 216 2561 229
rect 2351 195 2561 216
rect 2351 182 2527 195
rect 2317 166 2351 182
rect 2219 125 2253 161
rect 2624 316 2755 350
rect 2852 461 2920 544
rect 2852 427 2869 461
rect 2903 427 2920 461
rect 2852 387 2920 427
rect 2852 353 2869 387
rect 2903 353 2920 387
rect 3091 535 3125 923
rect 3091 433 3125 501
rect 3091 383 3125 399
rect 3313 957 3347 973
rect 3313 905 3347 923
rect 3313 433 3347 871
rect 3313 383 3347 399
rect 3535 957 3569 973
rect 3535 461 3569 923
rect 3535 383 3569 399
rect 3683 757 3717 1014
rect 3814 1019 3831 1053
rect 3865 1019 3882 1053
rect 4049 1366 4083 1446
rect 4049 1298 4083 1332
rect 4049 1230 4083 1264
rect 4049 1162 4083 1196
rect 4049 1093 4083 1128
rect 4049 1043 4083 1059
rect 4137 1366 4171 1404
rect 4137 1298 4171 1332
rect 4137 1230 4171 1264
rect 4137 1162 4171 1196
rect 4137 1093 4171 1128
rect 4225 1366 4259 1446
rect 4225 1298 4259 1332
rect 4225 1230 4259 1264
rect 4225 1162 4259 1196
rect 4225 1111 4259 1128
rect 4313 1366 4347 1404
rect 4313 1298 4347 1332
rect 4313 1230 4347 1264
rect 4313 1162 4347 1196
rect 4137 1048 4171 1059
rect 4313 1093 4347 1128
rect 4401 1366 4435 1446
rect 4401 1298 4435 1332
rect 4401 1230 4435 1264
rect 4401 1162 4435 1196
rect 4401 1111 4435 1128
rect 4489 1366 4523 1404
rect 4489 1298 4523 1332
rect 4489 1230 4523 1264
rect 4489 1162 4523 1196
rect 4313 1048 4347 1059
rect 4489 1093 4523 1128
rect 4577 1366 4611 1446
rect 4577 1298 4611 1332
rect 4577 1230 4611 1264
rect 4577 1162 4611 1196
rect 4577 1111 4611 1128
rect 4776 1423 4844 1446
rect 4776 1389 4793 1423
rect 4827 1389 4844 1423
rect 4776 1349 4844 1389
rect 4776 1315 4793 1349
rect 4827 1315 4844 1349
rect 4776 1275 4844 1315
rect 4776 1241 4793 1275
rect 4827 1241 4844 1275
rect 4776 1201 4844 1241
rect 4776 1167 4793 1201
rect 4827 1167 4844 1201
rect 4776 1127 4844 1167
rect 4489 1048 4523 1059
rect 4776 1093 4793 1127
rect 4827 1093 4844 1127
rect 4776 1053 4844 1093
rect 3814 979 3882 1019
rect 4137 1014 4679 1048
rect 3814 945 3831 979
rect 3865 945 3882 979
rect 4645 979 4679 1014
rect 3814 905 3882 945
rect 3814 871 3831 905
rect 3865 871 3882 905
rect 3814 822 3882 871
rect 4053 957 4087 973
rect 2624 219 2658 316
rect 2852 313 2920 353
rect 2852 279 2869 313
rect 2903 279 2920 313
rect 2624 169 2658 185
rect 2721 263 2755 279
rect 2721 195 2755 229
rect 2413 125 2447 141
rect 2253 91 2316 125
rect 2350 91 2413 125
rect 2219 75 2253 91
rect 2413 75 2447 91
rect 2527 125 2561 161
rect 2721 125 2755 161
rect 2561 91 2624 125
rect 2658 91 2721 125
rect 2527 75 2561 91
rect 2721 75 2755 91
rect 2852 239 2920 279
rect 2852 205 2869 239
rect 2903 205 2920 239
rect 2852 165 2920 205
rect 2852 131 2869 165
rect 2903 131 2920 165
rect 2852 91 2920 131
rect 2852 57 2869 91
rect 2903 57 2920 91
rect 2987 335 3021 351
rect 3181 335 3215 351
rect 3375 335 3409 351
rect 3021 301 3084 335
rect 3118 301 3181 335
rect 3215 301 3278 335
rect 3312 301 3375 335
rect 2987 263 3021 301
rect 2987 195 3021 229
rect 3181 263 3215 301
rect 3375 285 3409 301
rect 3489 335 3523 351
rect 3683 350 3717 723
rect 4053 683 4087 923
rect 3489 263 3523 301
rect 2987 125 3021 161
rect 2987 75 3021 91
rect 3084 210 3118 226
rect 2852 34 2920 57
rect 3084 34 3118 176
rect 3181 195 3215 229
rect 3279 216 3313 232
rect 3489 216 3523 229
rect 3313 195 3523 216
rect 3313 182 3489 195
rect 3279 166 3313 182
rect 3181 125 3215 161
rect 3586 316 3717 350
rect 3814 461 3882 544
rect 3814 427 3831 461
rect 3865 427 3882 461
rect 3814 387 3882 427
rect 3814 353 3831 387
rect 3865 353 3882 387
rect 4053 433 4087 649
rect 4053 383 4087 399
rect 4275 957 4309 973
rect 4275 461 4309 923
rect 4275 383 4309 399
rect 4497 957 4531 973
rect 4497 683 4531 923
rect 4497 433 4531 649
rect 4497 383 4531 399
rect 4645 535 4679 945
rect 4776 1019 4793 1053
rect 4827 1019 4844 1053
rect 5011 1366 5045 1446
rect 5011 1298 5045 1332
rect 5011 1230 5045 1264
rect 5011 1162 5045 1196
rect 5011 1093 5045 1128
rect 5011 1043 5045 1059
rect 5099 1366 5133 1404
rect 5099 1298 5133 1332
rect 5099 1230 5133 1264
rect 5099 1162 5133 1196
rect 5099 1093 5133 1128
rect 5187 1366 5221 1446
rect 5187 1298 5221 1332
rect 5187 1230 5221 1264
rect 5187 1162 5221 1196
rect 5187 1111 5221 1128
rect 5275 1366 5309 1404
rect 5275 1298 5309 1332
rect 5275 1230 5309 1264
rect 5275 1162 5309 1196
rect 5099 1048 5133 1059
rect 5275 1093 5309 1128
rect 5363 1366 5397 1446
rect 5363 1298 5397 1332
rect 5363 1230 5397 1264
rect 5363 1162 5397 1196
rect 5363 1111 5397 1128
rect 5451 1366 5485 1404
rect 5451 1298 5485 1332
rect 5451 1230 5485 1264
rect 5451 1162 5485 1196
rect 5275 1048 5309 1059
rect 5451 1093 5485 1128
rect 5539 1366 5573 1446
rect 5539 1298 5573 1332
rect 5539 1230 5573 1264
rect 5539 1162 5573 1196
rect 5539 1111 5573 1128
rect 5738 1423 5806 1446
rect 5738 1389 5755 1423
rect 5789 1389 5806 1423
rect 5738 1349 5806 1389
rect 5738 1315 5755 1349
rect 5789 1315 5806 1349
rect 5738 1275 5806 1315
rect 5738 1241 5755 1275
rect 5789 1241 5806 1275
rect 5738 1201 5806 1241
rect 5738 1167 5755 1201
rect 5789 1167 5806 1201
rect 5738 1127 5806 1167
rect 5451 1048 5485 1059
rect 5738 1093 5755 1127
rect 5789 1093 5806 1127
rect 5738 1053 5806 1093
rect 4776 979 4844 1019
rect 5099 1014 5641 1048
rect 4776 945 4793 979
rect 4827 945 4844 979
rect 4776 905 4844 945
rect 4776 871 4793 905
rect 4827 871 4844 905
rect 4776 822 4844 871
rect 5015 957 5049 973
rect 3586 219 3620 316
rect 3814 313 3882 353
rect 3814 279 3831 313
rect 3865 279 3882 313
rect 3586 169 3620 185
rect 3683 263 3717 279
rect 3683 195 3717 229
rect 3375 125 3409 141
rect 3215 91 3278 125
rect 3312 91 3375 125
rect 3181 75 3215 91
rect 3375 75 3409 91
rect 3489 125 3523 161
rect 3683 125 3717 161
rect 3523 91 3586 125
rect 3620 91 3683 125
rect 3489 75 3523 91
rect 3683 75 3717 91
rect 3814 239 3882 279
rect 3814 205 3831 239
rect 3865 205 3882 239
rect 3814 165 3882 205
rect 3814 131 3831 165
rect 3865 131 3882 165
rect 3814 91 3882 131
rect 3814 57 3831 91
rect 3865 57 3882 91
rect 3949 335 3983 351
rect 4143 335 4177 351
rect 4337 335 4371 351
rect 3983 301 4046 335
rect 4080 301 4143 335
rect 4177 301 4240 335
rect 4274 301 4337 335
rect 3949 263 3983 301
rect 3949 195 3983 229
rect 4143 263 4177 301
rect 4337 285 4371 301
rect 4451 335 4485 351
rect 4645 350 4679 501
rect 4451 263 4485 301
rect 3949 125 3983 161
rect 3949 75 3983 91
rect 4046 210 4080 226
rect 3814 34 3882 57
rect 4046 34 4080 176
rect 4143 195 4177 229
rect 4241 216 4275 232
rect 4451 216 4485 229
rect 4275 195 4485 216
rect 4275 182 4451 195
rect 4241 166 4275 182
rect 4143 125 4177 161
rect 4548 316 4679 350
rect 4776 461 4844 544
rect 4776 427 4793 461
rect 4827 427 4844 461
rect 4776 387 4844 427
rect 4776 353 4793 387
rect 4827 353 4844 387
rect 5015 535 5049 923
rect 5015 433 5049 501
rect 5015 383 5049 399
rect 5237 957 5271 973
rect 5237 609 5271 923
rect 5237 433 5271 575
rect 5237 383 5271 399
rect 5459 957 5493 973
rect 5459 757 5493 923
rect 5459 433 5493 723
rect 5459 383 5493 399
rect 5607 683 5641 1014
rect 5738 1019 5755 1053
rect 5789 1019 5806 1053
rect 5973 1366 6007 1446
rect 5973 1298 6007 1332
rect 5973 1230 6007 1264
rect 5973 1162 6007 1196
rect 5973 1093 6007 1128
rect 5973 1043 6007 1059
rect 6061 1366 6095 1404
rect 6061 1298 6095 1332
rect 6061 1230 6095 1264
rect 6061 1162 6095 1196
rect 6061 1093 6095 1128
rect 6149 1366 6183 1446
rect 6149 1298 6183 1332
rect 6149 1230 6183 1264
rect 6149 1162 6183 1196
rect 6149 1111 6183 1128
rect 6237 1366 6271 1404
rect 6237 1298 6271 1332
rect 6237 1230 6271 1264
rect 6237 1162 6271 1196
rect 6061 1048 6095 1059
rect 6237 1093 6271 1128
rect 6325 1366 6359 1446
rect 6325 1298 6359 1332
rect 6325 1230 6359 1264
rect 6325 1162 6359 1196
rect 6325 1111 6359 1128
rect 6413 1366 6447 1404
rect 6413 1298 6447 1332
rect 6413 1230 6447 1264
rect 6413 1162 6447 1196
rect 6237 1048 6271 1059
rect 6413 1093 6447 1128
rect 6501 1366 6535 1446
rect 6501 1298 6535 1332
rect 6501 1230 6535 1264
rect 6501 1162 6535 1196
rect 6501 1111 6535 1128
rect 6700 1423 6768 1446
rect 6700 1389 6717 1423
rect 6751 1389 6768 1423
rect 6700 1349 6768 1389
rect 6700 1315 6717 1349
rect 6751 1315 6768 1349
rect 6700 1275 6768 1315
rect 6700 1241 6717 1275
rect 6751 1241 6768 1275
rect 6700 1201 6768 1241
rect 6700 1167 6717 1201
rect 6751 1167 6768 1201
rect 6700 1127 6768 1167
rect 6413 1048 6447 1059
rect 6700 1093 6717 1127
rect 6751 1093 6768 1127
rect 6700 1053 6768 1093
rect 5738 979 5806 1019
rect 6061 1014 6603 1048
rect 5738 945 5755 979
rect 5789 945 5806 979
rect 5738 905 5806 945
rect 5738 871 5755 905
rect 5789 871 5806 905
rect 5738 822 5806 871
rect 5977 957 6011 973
rect 5977 831 6011 923
rect 4548 219 4582 316
rect 4776 313 4844 353
rect 4776 279 4793 313
rect 4827 279 4844 313
rect 4548 169 4582 185
rect 4645 263 4679 279
rect 4645 195 4679 229
rect 4337 125 4371 141
rect 4177 91 4240 125
rect 4274 91 4337 125
rect 4143 75 4177 91
rect 4337 75 4371 91
rect 4451 125 4485 161
rect 4645 125 4679 161
rect 4485 91 4548 125
rect 4582 91 4645 125
rect 4451 75 4485 91
rect 4645 75 4679 91
rect 4776 239 4844 279
rect 4776 205 4793 239
rect 4827 205 4844 239
rect 4776 165 4844 205
rect 4776 131 4793 165
rect 4827 131 4844 165
rect 4776 91 4844 131
rect 4776 57 4793 91
rect 4827 57 4844 91
rect 4911 335 4945 351
rect 5105 335 5139 351
rect 5299 335 5333 351
rect 4945 301 5008 335
rect 5042 301 5105 335
rect 5139 301 5202 335
rect 5236 301 5299 335
rect 4911 263 4945 301
rect 4911 195 4945 229
rect 5105 263 5139 301
rect 5299 285 5333 301
rect 5413 335 5447 351
rect 5607 350 5641 649
rect 5413 263 5447 301
rect 4911 125 4945 161
rect 4911 75 4945 91
rect 5008 210 5042 226
rect 4776 34 4844 57
rect 5008 34 5042 176
rect 5105 195 5139 229
rect 5203 216 5237 232
rect 5413 216 5447 229
rect 5237 195 5447 216
rect 5237 182 5413 195
rect 5203 166 5237 182
rect 5105 125 5139 161
rect 5510 316 5641 350
rect 5738 461 5806 544
rect 5738 427 5755 461
rect 5789 427 5806 461
rect 5738 387 5806 427
rect 5738 353 5755 387
rect 5789 353 5806 387
rect 5977 433 6011 797
rect 5977 383 6011 399
rect 6199 957 6233 973
rect 6199 461 6233 923
rect 6199 383 6233 399
rect 6421 957 6455 973
rect 6421 683 6455 923
rect 6421 433 6455 649
rect 6421 383 6455 399
rect 6569 535 6603 1014
rect 6700 1019 6717 1053
rect 6751 1019 6768 1053
rect 6935 1366 6969 1446
rect 6935 1298 6969 1332
rect 6935 1230 6969 1264
rect 6935 1162 6969 1196
rect 6935 1093 6969 1128
rect 6935 1043 6969 1059
rect 7023 1366 7057 1404
rect 7023 1298 7057 1332
rect 7023 1230 7057 1264
rect 7023 1162 7057 1196
rect 7023 1093 7057 1128
rect 7111 1366 7145 1446
rect 7111 1298 7145 1332
rect 7111 1230 7145 1264
rect 7111 1162 7145 1196
rect 7111 1111 7145 1128
rect 7199 1366 7233 1404
rect 7199 1298 7233 1332
rect 7199 1230 7233 1264
rect 7199 1162 7233 1196
rect 7023 1048 7057 1059
rect 7199 1093 7233 1128
rect 7287 1366 7321 1446
rect 7287 1298 7321 1332
rect 7287 1230 7321 1264
rect 7287 1162 7321 1196
rect 7287 1111 7321 1128
rect 7375 1366 7409 1404
rect 7375 1298 7409 1332
rect 7375 1230 7409 1264
rect 7375 1162 7409 1196
rect 7199 1048 7233 1059
rect 7375 1093 7409 1128
rect 7463 1366 7497 1446
rect 7463 1298 7497 1332
rect 7463 1230 7497 1264
rect 7463 1162 7497 1196
rect 7463 1111 7497 1128
rect 7662 1423 7730 1446
rect 7662 1389 7679 1423
rect 7713 1389 7730 1423
rect 7662 1349 7730 1389
rect 7662 1315 7679 1349
rect 7713 1315 7730 1349
rect 7662 1275 7730 1315
rect 7662 1241 7679 1275
rect 7713 1241 7730 1275
rect 7662 1201 7730 1241
rect 7662 1167 7679 1201
rect 7713 1167 7730 1201
rect 7662 1127 7730 1167
rect 7375 1048 7409 1059
rect 7662 1093 7679 1127
rect 7713 1093 7730 1127
rect 7662 1053 7730 1093
rect 6700 979 6768 1019
rect 7023 1014 7565 1048
rect 6700 945 6717 979
rect 6751 945 6768 979
rect 6700 905 6768 945
rect 6700 871 6717 905
rect 6751 871 6768 905
rect 6700 822 6768 871
rect 6939 957 6973 973
rect 5510 219 5544 316
rect 5738 313 5806 353
rect 5738 279 5755 313
rect 5789 279 5806 313
rect 5510 169 5544 185
rect 5607 263 5641 279
rect 5607 195 5641 229
rect 5299 125 5333 141
rect 5139 91 5202 125
rect 5236 91 5299 125
rect 5105 75 5139 91
rect 5299 75 5333 91
rect 5413 125 5447 161
rect 5607 125 5641 161
rect 5447 91 5510 125
rect 5544 91 5607 125
rect 5413 75 5447 91
rect 5607 75 5641 91
rect 5738 239 5806 279
rect 5738 205 5755 239
rect 5789 205 5806 239
rect 5738 165 5806 205
rect 5738 131 5755 165
rect 5789 131 5806 165
rect 5738 91 5806 131
rect 5738 57 5755 91
rect 5789 57 5806 91
rect 5873 335 5907 351
rect 6067 335 6101 351
rect 6261 335 6295 351
rect 5907 301 5970 335
rect 6004 301 6067 335
rect 6101 301 6164 335
rect 6198 301 6261 335
rect 5873 263 5907 301
rect 5873 195 5907 229
rect 6067 263 6101 301
rect 6261 285 6295 301
rect 6375 335 6409 351
rect 6569 350 6603 501
rect 6375 263 6409 301
rect 5873 125 5907 161
rect 5873 75 5907 91
rect 5970 210 6004 226
rect 5738 34 5806 57
rect 5970 34 6004 176
rect 6067 195 6101 229
rect 6165 216 6199 232
rect 6375 216 6409 229
rect 6199 195 6409 216
rect 6199 182 6375 195
rect 6165 166 6199 182
rect 6067 125 6101 161
rect 6472 316 6603 350
rect 6700 461 6768 544
rect 6700 427 6717 461
rect 6751 427 6768 461
rect 6700 387 6768 427
rect 6700 353 6717 387
rect 6751 353 6768 387
rect 6939 535 6973 923
rect 6939 433 6973 501
rect 6939 383 6973 399
rect 7161 957 7195 973
rect 7161 905 7195 923
rect 7161 433 7195 871
rect 7161 383 7195 399
rect 7383 957 7417 973
rect 7383 757 7417 923
rect 7383 433 7417 723
rect 7383 383 7417 399
rect 7531 683 7565 1014
rect 7662 1019 7679 1053
rect 7713 1019 7730 1053
rect 7897 1366 7931 1446
rect 7897 1298 7931 1332
rect 7897 1230 7931 1264
rect 7897 1162 7931 1196
rect 7897 1093 7931 1128
rect 7897 1043 7931 1059
rect 7985 1366 8019 1404
rect 7985 1298 8019 1332
rect 7985 1230 8019 1264
rect 7985 1162 8019 1196
rect 7985 1093 8019 1128
rect 8073 1366 8107 1446
rect 8073 1298 8107 1332
rect 8073 1230 8107 1264
rect 8073 1162 8107 1196
rect 8073 1111 8107 1128
rect 8161 1366 8195 1404
rect 8161 1298 8195 1332
rect 8161 1230 8195 1264
rect 8161 1162 8195 1196
rect 7985 1048 8019 1059
rect 8161 1093 8195 1128
rect 8249 1366 8283 1446
rect 8249 1298 8283 1332
rect 8249 1230 8283 1264
rect 8249 1162 8283 1196
rect 8249 1111 8283 1128
rect 8337 1366 8371 1404
rect 8337 1298 8371 1332
rect 8337 1230 8371 1264
rect 8337 1162 8371 1196
rect 8161 1048 8195 1059
rect 8337 1093 8371 1128
rect 8425 1366 8459 1446
rect 8425 1298 8459 1332
rect 8425 1230 8459 1264
rect 8425 1162 8459 1196
rect 8425 1111 8459 1128
rect 8624 1423 8692 1446
rect 8624 1389 8641 1423
rect 8675 1389 8692 1423
rect 8624 1349 8692 1389
rect 8624 1315 8641 1349
rect 8675 1315 8692 1349
rect 8624 1275 8692 1315
rect 8624 1241 8641 1275
rect 8675 1241 8692 1275
rect 8624 1201 8692 1241
rect 8624 1167 8641 1201
rect 8675 1167 8692 1201
rect 8624 1127 8692 1167
rect 8337 1048 8371 1059
rect 8624 1093 8641 1127
rect 8675 1093 8692 1127
rect 8624 1053 8692 1093
rect 7662 979 7730 1019
rect 7985 1014 8527 1048
rect 7662 945 7679 979
rect 7713 945 7730 979
rect 7662 905 7730 945
rect 7662 871 7679 905
rect 7713 871 7730 905
rect 7662 822 7730 871
rect 7901 957 7935 973
rect 6472 219 6506 316
rect 6700 313 6768 353
rect 6700 279 6717 313
rect 6751 279 6768 313
rect 6472 169 6506 185
rect 6569 263 6603 279
rect 6569 195 6603 229
rect 6261 125 6295 141
rect 6101 91 6164 125
rect 6198 91 6261 125
rect 6067 75 6101 91
rect 6261 75 6295 91
rect 6375 125 6409 161
rect 6569 125 6603 161
rect 6409 91 6472 125
rect 6506 91 6569 125
rect 6375 75 6409 91
rect 6569 75 6603 91
rect 6700 239 6768 279
rect 6700 205 6717 239
rect 6751 205 6768 239
rect 6700 165 6768 205
rect 6700 131 6717 165
rect 6751 131 6768 165
rect 6700 91 6768 131
rect 6700 57 6717 91
rect 6751 57 6768 91
rect 6835 335 6869 351
rect 7029 335 7063 351
rect 7223 335 7257 351
rect 6869 301 6932 335
rect 6966 301 7029 335
rect 7063 301 7126 335
rect 7160 301 7223 335
rect 6835 263 6869 301
rect 6835 195 6869 229
rect 7029 263 7063 301
rect 7223 285 7257 301
rect 7337 335 7371 351
rect 7531 350 7565 649
rect 7337 263 7371 301
rect 6835 125 6869 161
rect 6835 75 6869 91
rect 6932 210 6966 226
rect 6700 34 6768 57
rect 6932 34 6966 176
rect 7029 195 7063 229
rect 7127 216 7161 232
rect 7337 216 7371 229
rect 7161 195 7371 216
rect 7161 182 7337 195
rect 7127 166 7161 182
rect 7029 125 7063 161
rect 7434 316 7565 350
rect 7662 461 7730 544
rect 7662 427 7679 461
rect 7713 427 7730 461
rect 7662 387 7730 427
rect 7662 353 7679 387
rect 7713 353 7730 387
rect 7901 535 7935 923
rect 7901 433 7935 501
rect 7901 383 7935 399
rect 8123 957 8157 973
rect 8123 609 8157 923
rect 8123 433 8157 575
rect 8123 383 8157 399
rect 8345 957 8379 973
rect 8345 757 8379 923
rect 8345 433 8379 723
rect 8345 383 8379 399
rect 8493 535 8527 1014
rect 8624 1019 8641 1053
rect 8675 1019 8692 1053
rect 8859 1366 8893 1446
rect 8859 1298 8893 1332
rect 8859 1230 8893 1264
rect 8859 1162 8893 1196
rect 8859 1093 8893 1128
rect 8859 1043 8893 1059
rect 8947 1366 8981 1404
rect 8947 1298 8981 1332
rect 8947 1230 8981 1264
rect 8947 1162 8981 1196
rect 8947 1093 8981 1128
rect 9035 1366 9069 1446
rect 9035 1298 9069 1332
rect 9035 1230 9069 1264
rect 9035 1162 9069 1196
rect 9035 1111 9069 1128
rect 9123 1366 9157 1404
rect 9123 1298 9157 1332
rect 9123 1230 9157 1264
rect 9123 1162 9157 1196
rect 8947 1048 8981 1059
rect 9123 1093 9157 1128
rect 9211 1366 9245 1446
rect 9211 1298 9245 1332
rect 9211 1230 9245 1264
rect 9211 1162 9245 1196
rect 9211 1111 9245 1128
rect 9299 1366 9333 1404
rect 9299 1298 9333 1332
rect 9299 1230 9333 1264
rect 9299 1162 9333 1196
rect 9123 1048 9157 1059
rect 9299 1093 9333 1128
rect 9387 1366 9421 1446
rect 9387 1298 9421 1332
rect 9387 1230 9421 1264
rect 9387 1162 9421 1196
rect 9387 1111 9421 1128
rect 9586 1423 9654 1446
rect 9586 1389 9603 1423
rect 9637 1389 9654 1423
rect 9586 1349 9654 1389
rect 9586 1315 9603 1349
rect 9637 1315 9654 1349
rect 9586 1275 9654 1315
rect 9586 1241 9603 1275
rect 9637 1241 9654 1275
rect 9586 1201 9654 1241
rect 9586 1167 9603 1201
rect 9637 1167 9654 1201
rect 9586 1127 9654 1167
rect 9299 1048 9333 1059
rect 9586 1093 9603 1127
rect 9637 1093 9654 1127
rect 9586 1053 9654 1093
rect 8624 979 8692 1019
rect 8947 1014 9489 1048
rect 8624 945 8641 979
rect 8675 945 8692 979
rect 8624 905 8692 945
rect 8624 871 8641 905
rect 8675 871 8692 905
rect 8624 822 8692 871
rect 8863 957 8897 973
rect 7434 219 7468 316
rect 7662 313 7730 353
rect 7662 279 7679 313
rect 7713 279 7730 313
rect 7434 169 7468 185
rect 7531 263 7565 279
rect 7531 195 7565 229
rect 7223 125 7257 141
rect 7063 91 7126 125
rect 7160 91 7223 125
rect 7029 75 7063 91
rect 7223 75 7257 91
rect 7337 125 7371 161
rect 7531 125 7565 161
rect 7371 91 7434 125
rect 7468 91 7531 125
rect 7337 75 7371 91
rect 7531 75 7565 91
rect 7662 239 7730 279
rect 7662 205 7679 239
rect 7713 205 7730 239
rect 7662 165 7730 205
rect 7662 131 7679 165
rect 7713 131 7730 165
rect 7662 91 7730 131
rect 7662 57 7679 91
rect 7713 57 7730 91
rect 7797 335 7831 351
rect 7991 335 8025 351
rect 8185 335 8219 351
rect 7831 301 7894 335
rect 7928 301 7991 335
rect 8025 301 8088 335
rect 8122 301 8185 335
rect 7797 263 7831 301
rect 7797 195 7831 229
rect 7991 263 8025 301
rect 8185 285 8219 301
rect 8299 335 8333 351
rect 8493 350 8527 501
rect 8299 263 8333 301
rect 7797 125 7831 161
rect 7797 75 7831 91
rect 7894 210 7928 226
rect 7662 34 7730 57
rect 7894 34 7928 176
rect 7991 195 8025 229
rect 8089 216 8123 232
rect 8299 216 8333 229
rect 8123 195 8333 216
rect 8123 182 8299 195
rect 8089 166 8123 182
rect 7991 125 8025 161
rect 8396 316 8527 350
rect 8624 461 8692 544
rect 8624 427 8641 461
rect 8675 427 8692 461
rect 8624 387 8692 427
rect 8624 353 8641 387
rect 8675 353 8692 387
rect 8863 535 8897 923
rect 8863 433 8897 501
rect 8863 383 8897 399
rect 9085 957 9119 973
rect 9085 905 9119 923
rect 9085 433 9119 871
rect 9085 383 9119 399
rect 9307 957 9341 973
rect 9307 461 9341 923
rect 9307 383 9341 399
rect 9455 757 9489 1014
rect 9586 1019 9603 1053
rect 9637 1019 9654 1053
rect 9821 1366 9855 1446
rect 9821 1298 9855 1332
rect 9821 1230 9855 1264
rect 9821 1162 9855 1196
rect 9821 1093 9855 1128
rect 9821 1043 9855 1059
rect 9909 1366 9943 1404
rect 9909 1298 9943 1332
rect 9909 1230 9943 1264
rect 9909 1162 9943 1196
rect 9909 1093 9943 1128
rect 9997 1366 10031 1446
rect 9997 1298 10031 1332
rect 9997 1230 10031 1264
rect 9997 1162 10031 1196
rect 9997 1111 10031 1128
rect 10085 1366 10119 1404
rect 10085 1298 10119 1332
rect 10085 1230 10119 1264
rect 10085 1162 10119 1196
rect 9909 1048 9943 1059
rect 10085 1093 10119 1128
rect 10173 1366 10207 1446
rect 10173 1298 10207 1332
rect 10173 1230 10207 1264
rect 10173 1162 10207 1196
rect 10173 1111 10207 1128
rect 10261 1366 10295 1404
rect 10261 1298 10295 1332
rect 10261 1230 10295 1264
rect 10261 1162 10295 1196
rect 10085 1048 10119 1059
rect 10261 1093 10295 1128
rect 10349 1366 10383 1446
rect 10349 1298 10383 1332
rect 10349 1230 10383 1264
rect 10349 1162 10383 1196
rect 10349 1111 10383 1128
rect 10548 1423 10616 1446
rect 10548 1389 10565 1423
rect 10599 1389 10616 1423
rect 10548 1349 10616 1389
rect 10548 1315 10565 1349
rect 10599 1315 10616 1349
rect 10548 1275 10616 1315
rect 10548 1241 10565 1275
rect 10599 1241 10616 1275
rect 10548 1201 10616 1241
rect 10548 1167 10565 1201
rect 10599 1167 10616 1201
rect 10548 1127 10616 1167
rect 10261 1048 10295 1059
rect 10548 1093 10565 1127
rect 10599 1093 10616 1127
rect 10548 1053 10616 1093
rect 9586 979 9654 1019
rect 9909 1014 10451 1048
rect 9586 945 9603 979
rect 9637 945 9654 979
rect 9586 905 9654 945
rect 9586 871 9603 905
rect 9637 871 9654 905
rect 9586 822 9654 871
rect 9825 957 9859 973
rect 8396 219 8430 316
rect 8624 313 8692 353
rect 8624 279 8641 313
rect 8675 279 8692 313
rect 8396 169 8430 185
rect 8493 263 8527 279
rect 8493 195 8527 229
rect 8185 125 8219 141
rect 8025 91 8088 125
rect 8122 91 8185 125
rect 7991 75 8025 91
rect 8185 75 8219 91
rect 8299 125 8333 161
rect 8493 125 8527 161
rect 8333 91 8396 125
rect 8430 91 8493 125
rect 8299 75 8333 91
rect 8493 75 8527 91
rect 8624 239 8692 279
rect 8624 205 8641 239
rect 8675 205 8692 239
rect 8624 165 8692 205
rect 8624 131 8641 165
rect 8675 131 8692 165
rect 8624 91 8692 131
rect 8624 57 8641 91
rect 8675 57 8692 91
rect 8759 335 8793 351
rect 8953 335 8987 351
rect 9147 335 9181 351
rect 8793 301 8856 335
rect 8890 301 8953 335
rect 8987 301 9050 335
rect 9084 301 9147 335
rect 8759 263 8793 301
rect 8759 195 8793 229
rect 8953 263 8987 301
rect 9147 285 9181 301
rect 9261 335 9295 351
rect 9455 350 9489 723
rect 9825 683 9859 923
rect 9261 263 9295 301
rect 8759 125 8793 161
rect 8759 75 8793 91
rect 8856 210 8890 226
rect 8624 34 8692 57
rect 8856 34 8890 176
rect 8953 195 8987 229
rect 9051 216 9085 232
rect 9261 216 9295 229
rect 9085 195 9295 216
rect 9085 182 9261 195
rect 9051 166 9085 182
rect 8953 125 8987 161
rect 9358 316 9489 350
rect 9586 461 9654 544
rect 9586 427 9603 461
rect 9637 427 9654 461
rect 9586 387 9654 427
rect 9586 353 9603 387
rect 9637 353 9654 387
rect 9825 433 9859 649
rect 9825 383 9859 399
rect 10047 957 10081 973
rect 10047 461 10081 923
rect 10047 383 10081 399
rect 10269 957 10303 973
rect 10269 535 10303 923
rect 10269 433 10303 501
rect 10269 383 10303 399
rect 10417 683 10451 1014
rect 10548 1019 10565 1053
rect 10599 1019 10616 1053
rect 10783 1366 10817 1446
rect 10783 1298 10817 1332
rect 10783 1230 10817 1264
rect 10783 1162 10817 1196
rect 10783 1093 10817 1128
rect 10783 1043 10817 1059
rect 10871 1366 10905 1404
rect 10871 1298 10905 1332
rect 10871 1230 10905 1264
rect 10871 1162 10905 1196
rect 10871 1093 10905 1128
rect 10959 1366 10993 1446
rect 10959 1298 10993 1332
rect 10959 1230 10993 1264
rect 10959 1162 10993 1196
rect 10959 1111 10993 1128
rect 11047 1366 11081 1404
rect 11047 1298 11081 1332
rect 11047 1230 11081 1264
rect 11047 1162 11081 1196
rect 10871 1048 10905 1059
rect 11047 1093 11081 1128
rect 11135 1366 11169 1446
rect 11135 1298 11169 1332
rect 11135 1230 11169 1264
rect 11135 1162 11169 1196
rect 11135 1111 11169 1128
rect 11223 1366 11257 1404
rect 11223 1298 11257 1332
rect 11223 1230 11257 1264
rect 11223 1162 11257 1196
rect 11047 1048 11081 1059
rect 11223 1093 11257 1128
rect 11311 1366 11345 1446
rect 11311 1298 11345 1332
rect 11311 1230 11345 1264
rect 11311 1162 11345 1196
rect 11311 1111 11345 1128
rect 11510 1423 11578 1446
rect 11510 1389 11527 1423
rect 11561 1389 11578 1423
rect 11510 1349 11578 1389
rect 11510 1315 11527 1349
rect 11561 1315 11578 1349
rect 11510 1275 11578 1315
rect 11510 1241 11527 1275
rect 11561 1241 11578 1275
rect 11510 1201 11578 1241
rect 11510 1167 11527 1201
rect 11561 1167 11578 1201
rect 11510 1127 11578 1167
rect 11223 1048 11257 1059
rect 11510 1093 11527 1127
rect 11561 1093 11578 1127
rect 11510 1053 11578 1093
rect 10548 979 10616 1019
rect 10871 1014 11413 1048
rect 10548 945 10565 979
rect 10599 945 10616 979
rect 10548 905 10616 945
rect 10548 871 10565 905
rect 10599 871 10616 905
rect 10548 822 10616 871
rect 10787 957 10821 973
rect 9358 219 9392 316
rect 9586 313 9654 353
rect 9586 279 9603 313
rect 9637 279 9654 313
rect 9358 169 9392 185
rect 9455 263 9489 279
rect 9455 195 9489 229
rect 9147 125 9181 141
rect 8987 91 9050 125
rect 9084 91 9147 125
rect 8953 75 8987 91
rect 9147 75 9181 91
rect 9261 125 9295 161
rect 9455 125 9489 161
rect 9295 91 9358 125
rect 9392 91 9455 125
rect 9261 75 9295 91
rect 9455 75 9489 91
rect 9586 239 9654 279
rect 9586 205 9603 239
rect 9637 205 9654 239
rect 9586 165 9654 205
rect 9586 131 9603 165
rect 9637 131 9654 165
rect 9586 91 9654 131
rect 9586 57 9603 91
rect 9637 57 9654 91
rect 9721 335 9755 351
rect 9915 335 9949 351
rect 10109 335 10143 351
rect 9755 301 9818 335
rect 9852 301 9915 335
rect 9949 301 10012 335
rect 10046 301 10109 335
rect 9721 263 9755 301
rect 9721 195 9755 229
rect 9915 263 9949 301
rect 10109 285 10143 301
rect 10223 335 10257 351
rect 10417 350 10451 649
rect 10787 683 10821 923
rect 10223 263 10257 301
rect 9721 125 9755 161
rect 9721 75 9755 91
rect 9818 210 9852 226
rect 9586 34 9654 57
rect 9818 34 9852 176
rect 9915 195 9949 229
rect 10013 216 10047 232
rect 10223 216 10257 229
rect 10047 195 10257 216
rect 10047 182 10223 195
rect 10013 166 10047 182
rect 9915 125 9949 161
rect 10320 316 10451 350
rect 10548 461 10616 544
rect 10548 427 10565 461
rect 10599 427 10616 461
rect 10548 387 10616 427
rect 10548 353 10565 387
rect 10599 353 10616 387
rect 10787 433 10821 649
rect 10787 383 10821 399
rect 11009 957 11043 973
rect 11009 609 11043 923
rect 11009 433 11043 575
rect 11009 383 11043 399
rect 11231 957 11265 973
rect 11231 757 11265 923
rect 11231 433 11265 723
rect 11231 383 11265 399
rect 11379 535 11413 1014
rect 11510 1019 11527 1053
rect 11561 1019 11578 1053
rect 11745 1366 11779 1446
rect 11745 1298 11779 1332
rect 11745 1230 11779 1264
rect 11745 1162 11779 1196
rect 11745 1093 11779 1128
rect 11745 1043 11779 1059
rect 11833 1366 11867 1404
rect 11833 1298 11867 1332
rect 11833 1230 11867 1264
rect 11833 1162 11867 1196
rect 11833 1093 11867 1128
rect 11921 1366 11955 1446
rect 11921 1298 11955 1332
rect 11921 1230 11955 1264
rect 11921 1162 11955 1196
rect 11921 1111 11955 1128
rect 12009 1366 12043 1404
rect 12009 1298 12043 1332
rect 12009 1230 12043 1264
rect 12009 1162 12043 1196
rect 11833 1048 11867 1059
rect 12009 1093 12043 1128
rect 12097 1366 12131 1446
rect 12097 1298 12131 1332
rect 12097 1230 12131 1264
rect 12097 1162 12131 1196
rect 12097 1111 12131 1128
rect 12185 1366 12219 1404
rect 12185 1298 12219 1332
rect 12185 1230 12219 1264
rect 12185 1162 12219 1196
rect 12009 1048 12043 1059
rect 12185 1093 12219 1128
rect 12273 1366 12307 1446
rect 12273 1298 12307 1332
rect 12273 1230 12307 1264
rect 12273 1162 12307 1196
rect 12273 1111 12307 1128
rect 12472 1423 12540 1446
rect 12472 1389 12489 1423
rect 12523 1389 12540 1423
rect 12472 1349 12540 1389
rect 12472 1315 12489 1349
rect 12523 1315 12540 1349
rect 12472 1275 12540 1315
rect 12472 1241 12489 1275
rect 12523 1241 12540 1275
rect 12472 1201 12540 1241
rect 12472 1167 12489 1201
rect 12523 1167 12540 1201
rect 12472 1127 12540 1167
rect 12185 1048 12219 1059
rect 12472 1093 12489 1127
rect 12523 1093 12540 1127
rect 12472 1053 12540 1093
rect 11510 979 11578 1019
rect 11833 1014 12375 1048
rect 11510 945 11527 979
rect 11561 945 11578 979
rect 11510 905 11578 945
rect 11510 871 11527 905
rect 11561 871 11578 905
rect 11510 822 11578 871
rect 11749 957 11783 973
rect 11749 831 11783 923
rect 10320 219 10354 316
rect 10548 313 10616 353
rect 10548 279 10565 313
rect 10599 279 10616 313
rect 10320 169 10354 185
rect 10417 263 10451 279
rect 10417 195 10451 229
rect 10109 125 10143 141
rect 9949 91 10012 125
rect 10046 91 10109 125
rect 9915 75 9949 91
rect 10109 75 10143 91
rect 10223 125 10257 161
rect 10417 125 10451 161
rect 10257 91 10320 125
rect 10354 91 10417 125
rect 10223 75 10257 91
rect 10417 75 10451 91
rect 10548 239 10616 279
rect 10548 205 10565 239
rect 10599 205 10616 239
rect 10548 165 10616 205
rect 10548 131 10565 165
rect 10599 131 10616 165
rect 10548 91 10616 131
rect 10548 57 10565 91
rect 10599 57 10616 91
rect 10683 335 10717 351
rect 10877 335 10911 351
rect 11071 335 11105 351
rect 10717 301 10780 335
rect 10814 301 10877 335
rect 10911 301 10974 335
rect 11008 301 11071 335
rect 10683 263 10717 301
rect 10683 195 10717 229
rect 10877 263 10911 301
rect 11071 285 11105 301
rect 11185 335 11219 351
rect 11379 350 11413 501
rect 11185 263 11219 301
rect 10683 125 10717 161
rect 10683 75 10717 91
rect 10780 210 10814 226
rect 10548 34 10616 57
rect 10780 34 10814 176
rect 10877 195 10911 229
rect 10975 216 11009 232
rect 11185 216 11219 229
rect 11009 195 11219 216
rect 11009 182 11185 195
rect 10975 166 11009 182
rect 10877 125 10911 161
rect 11282 316 11413 350
rect 11510 461 11578 544
rect 11510 427 11527 461
rect 11561 427 11578 461
rect 11510 387 11578 427
rect 11510 353 11527 387
rect 11561 353 11578 387
rect 11749 433 11783 797
rect 11749 383 11783 399
rect 11971 957 12005 973
rect 11971 461 12005 923
rect 11971 383 12005 399
rect 12193 957 12227 973
rect 12193 683 12227 923
rect 12193 433 12227 649
rect 12193 383 12227 399
rect 12341 535 12375 1014
rect 12472 1019 12489 1053
rect 12523 1019 12540 1053
rect 12707 1366 12741 1446
rect 12707 1298 12741 1332
rect 12707 1230 12741 1264
rect 12707 1162 12741 1196
rect 12707 1093 12741 1128
rect 12707 1043 12741 1059
rect 12795 1366 12829 1404
rect 12795 1298 12829 1332
rect 12795 1230 12829 1264
rect 12795 1162 12829 1196
rect 12795 1093 12829 1128
rect 12883 1366 12917 1446
rect 12883 1298 12917 1332
rect 12883 1230 12917 1264
rect 12883 1162 12917 1196
rect 12883 1111 12917 1128
rect 12971 1366 13005 1404
rect 12971 1298 13005 1332
rect 12971 1230 13005 1264
rect 12971 1162 13005 1196
rect 12795 1048 12829 1059
rect 12971 1093 13005 1128
rect 13059 1366 13093 1446
rect 13059 1298 13093 1332
rect 13059 1230 13093 1264
rect 13059 1162 13093 1196
rect 13059 1111 13093 1128
rect 13147 1366 13181 1404
rect 13147 1298 13181 1332
rect 13147 1230 13181 1264
rect 13147 1162 13181 1196
rect 12971 1048 13005 1059
rect 13147 1093 13181 1128
rect 13235 1366 13269 1446
rect 13235 1298 13269 1332
rect 13235 1230 13269 1264
rect 13235 1162 13269 1196
rect 13235 1111 13269 1128
rect 13434 1423 13502 1446
rect 13434 1389 13451 1423
rect 13485 1389 13502 1423
rect 13434 1349 13502 1389
rect 13434 1315 13451 1349
rect 13485 1315 13502 1349
rect 13434 1275 13502 1315
rect 13434 1241 13451 1275
rect 13485 1241 13502 1275
rect 13434 1201 13502 1241
rect 13434 1167 13451 1201
rect 13485 1167 13502 1201
rect 13434 1127 13502 1167
rect 13147 1048 13181 1059
rect 13434 1093 13451 1127
rect 13485 1093 13502 1127
rect 13434 1053 13502 1093
rect 12472 979 12540 1019
rect 12795 1014 13337 1048
rect 12472 945 12489 979
rect 12523 945 12540 979
rect 12472 905 12540 945
rect 12472 871 12489 905
rect 12523 871 12540 905
rect 12472 822 12540 871
rect 12711 957 12745 973
rect 11282 219 11316 316
rect 11510 313 11578 353
rect 11510 279 11527 313
rect 11561 279 11578 313
rect 11282 169 11316 185
rect 11379 263 11413 279
rect 11379 195 11413 229
rect 11071 125 11105 141
rect 10911 91 10974 125
rect 11008 91 11071 125
rect 10877 75 10911 91
rect 11071 75 11105 91
rect 11185 125 11219 161
rect 11379 125 11413 161
rect 11219 91 11282 125
rect 11316 91 11379 125
rect 11185 75 11219 91
rect 11379 75 11413 91
rect 11510 239 11578 279
rect 11510 205 11527 239
rect 11561 205 11578 239
rect 11510 165 11578 205
rect 11510 131 11527 165
rect 11561 131 11578 165
rect 11510 91 11578 131
rect 11510 57 11527 91
rect 11561 57 11578 91
rect 11645 335 11679 351
rect 11839 335 11873 351
rect 12033 335 12067 351
rect 11679 301 11742 335
rect 11776 301 11839 335
rect 11873 301 11936 335
rect 11970 301 12033 335
rect 11645 263 11679 301
rect 11645 195 11679 229
rect 11839 263 11873 301
rect 12033 285 12067 301
rect 12147 335 12181 351
rect 12341 350 12375 501
rect 12147 263 12181 301
rect 11645 125 11679 161
rect 11645 75 11679 91
rect 11742 210 11776 226
rect 11510 34 11578 57
rect 11742 34 11776 176
rect 11839 195 11873 229
rect 11937 216 11971 232
rect 12147 216 12181 229
rect 11971 195 12181 216
rect 11971 182 12147 195
rect 11937 166 11971 182
rect 11839 125 11873 161
rect 12244 316 12375 350
rect 12472 461 12540 544
rect 12472 427 12489 461
rect 12523 427 12540 461
rect 12472 387 12540 427
rect 12472 353 12489 387
rect 12523 353 12540 387
rect 12711 535 12745 923
rect 12711 433 12745 501
rect 12711 383 12745 399
rect 12933 957 12967 973
rect 12933 905 12967 923
rect 12933 433 12967 871
rect 12933 383 12967 399
rect 13155 957 13189 973
rect 13155 757 13189 923
rect 13155 433 13189 723
rect 13155 383 13189 399
rect 13303 683 13337 1014
rect 13434 1019 13451 1053
rect 13485 1019 13502 1053
rect 13669 1366 13703 1446
rect 13669 1298 13703 1332
rect 13669 1230 13703 1264
rect 13669 1162 13703 1196
rect 13669 1093 13703 1128
rect 13669 1043 13703 1059
rect 13757 1366 13791 1404
rect 13757 1298 13791 1332
rect 13757 1230 13791 1264
rect 13757 1162 13791 1196
rect 13757 1093 13791 1128
rect 13845 1366 13879 1446
rect 13845 1298 13879 1332
rect 13845 1230 13879 1264
rect 13845 1162 13879 1196
rect 13845 1111 13879 1128
rect 13933 1366 13967 1404
rect 13933 1298 13967 1332
rect 13933 1230 13967 1264
rect 13933 1162 13967 1196
rect 13757 1048 13791 1059
rect 13933 1093 13967 1128
rect 14021 1366 14055 1446
rect 14021 1298 14055 1332
rect 14021 1230 14055 1264
rect 14021 1162 14055 1196
rect 14021 1111 14055 1128
rect 14109 1366 14143 1404
rect 14109 1298 14143 1332
rect 14109 1230 14143 1264
rect 14109 1162 14143 1196
rect 13933 1048 13967 1059
rect 14109 1093 14143 1128
rect 14197 1366 14231 1446
rect 14197 1298 14231 1332
rect 14197 1230 14231 1264
rect 14197 1162 14231 1196
rect 14197 1111 14231 1128
rect 14396 1423 14464 1446
rect 14396 1389 14413 1423
rect 14447 1389 14464 1423
rect 14396 1349 14464 1389
rect 14396 1315 14413 1349
rect 14447 1315 14464 1349
rect 14396 1275 14464 1315
rect 14396 1241 14413 1275
rect 14447 1241 14464 1275
rect 14396 1201 14464 1241
rect 14396 1167 14413 1201
rect 14447 1167 14464 1201
rect 14396 1127 14464 1167
rect 14109 1048 14143 1059
rect 14396 1093 14413 1127
rect 14447 1093 14464 1127
rect 14396 1053 14464 1093
rect 13434 979 13502 1019
rect 13757 1014 14299 1048
rect 13434 945 13451 979
rect 13485 945 13502 979
rect 13434 905 13502 945
rect 13434 871 13451 905
rect 13485 871 13502 905
rect 13434 822 13502 871
rect 13673 957 13707 973
rect 12244 219 12278 316
rect 12472 313 12540 353
rect 12472 279 12489 313
rect 12523 279 12540 313
rect 12244 169 12278 185
rect 12341 263 12375 279
rect 12341 195 12375 229
rect 12033 125 12067 141
rect 11873 91 11936 125
rect 11970 91 12033 125
rect 11839 75 11873 91
rect 12033 75 12067 91
rect 12147 125 12181 161
rect 12341 125 12375 161
rect 12181 91 12244 125
rect 12278 91 12341 125
rect 12147 75 12181 91
rect 12341 75 12375 91
rect 12472 239 12540 279
rect 12472 205 12489 239
rect 12523 205 12540 239
rect 12472 165 12540 205
rect 12472 131 12489 165
rect 12523 131 12540 165
rect 12472 91 12540 131
rect 12472 57 12489 91
rect 12523 57 12540 91
rect 12607 335 12641 351
rect 12801 335 12835 351
rect 12995 335 13029 351
rect 12641 301 12704 335
rect 12738 301 12801 335
rect 12835 301 12898 335
rect 12932 301 12995 335
rect 12607 263 12641 301
rect 12607 195 12641 229
rect 12801 263 12835 301
rect 12995 285 13029 301
rect 13109 335 13143 351
rect 13303 350 13337 649
rect 13109 263 13143 301
rect 12607 125 12641 161
rect 12607 75 12641 91
rect 12704 210 12738 226
rect 12472 34 12540 57
rect 12704 34 12738 176
rect 12801 195 12835 229
rect 12899 216 12933 232
rect 13109 216 13143 229
rect 12933 195 13143 216
rect 12933 182 13109 195
rect 12899 166 12933 182
rect 12801 125 12835 161
rect 13206 316 13337 350
rect 13434 461 13502 544
rect 13434 427 13451 461
rect 13485 427 13502 461
rect 13434 387 13502 427
rect 13434 353 13451 387
rect 13485 353 13502 387
rect 13673 535 13707 923
rect 13673 433 13707 501
rect 13673 383 13707 399
rect 13895 957 13929 973
rect 13895 609 13929 923
rect 13895 433 13929 575
rect 13895 383 13929 399
rect 14117 957 14151 973
rect 14117 757 14151 923
rect 14117 433 14151 723
rect 14117 383 14151 399
rect 14265 535 14299 1014
rect 14396 1019 14413 1053
rect 14447 1019 14464 1053
rect 14631 1366 14665 1446
rect 14631 1298 14665 1332
rect 14631 1230 14665 1264
rect 14631 1162 14665 1196
rect 14631 1093 14665 1128
rect 14631 1043 14665 1059
rect 14719 1366 14753 1404
rect 14719 1298 14753 1332
rect 14719 1230 14753 1264
rect 14719 1162 14753 1196
rect 14719 1093 14753 1128
rect 14807 1366 14841 1446
rect 14807 1298 14841 1332
rect 14807 1230 14841 1264
rect 14807 1162 14841 1196
rect 14807 1111 14841 1128
rect 14895 1366 14929 1404
rect 14895 1298 14929 1332
rect 14895 1230 14929 1264
rect 14895 1162 14929 1196
rect 14719 1048 14753 1059
rect 14895 1093 14929 1128
rect 14983 1366 15017 1446
rect 14983 1298 15017 1332
rect 14983 1230 15017 1264
rect 14983 1162 15017 1196
rect 14983 1111 15017 1128
rect 15071 1366 15105 1404
rect 15071 1298 15105 1332
rect 15071 1230 15105 1264
rect 15071 1162 15105 1196
rect 14895 1048 14929 1059
rect 15071 1093 15105 1128
rect 15159 1366 15193 1446
rect 15159 1298 15193 1332
rect 15159 1230 15193 1264
rect 15159 1162 15193 1196
rect 15159 1111 15193 1128
rect 15358 1423 15426 1446
rect 15358 1389 15375 1423
rect 15409 1389 15426 1423
rect 15358 1349 15426 1389
rect 15358 1315 15375 1349
rect 15409 1315 15426 1349
rect 15358 1275 15426 1315
rect 15358 1241 15375 1275
rect 15409 1241 15426 1275
rect 15358 1201 15426 1241
rect 15358 1167 15375 1201
rect 15409 1167 15426 1201
rect 15358 1127 15426 1167
rect 15071 1048 15105 1059
rect 15358 1093 15375 1127
rect 15409 1093 15426 1127
rect 15358 1053 15426 1093
rect 14396 979 14464 1019
rect 14719 1014 15261 1048
rect 14396 945 14413 979
rect 14447 945 14464 979
rect 14396 905 14464 945
rect 14396 871 14413 905
rect 14447 871 14464 905
rect 14396 822 14464 871
rect 14635 957 14669 973
rect 13206 219 13240 316
rect 13434 313 13502 353
rect 13434 279 13451 313
rect 13485 279 13502 313
rect 13206 169 13240 185
rect 13303 263 13337 279
rect 13303 195 13337 229
rect 12995 125 13029 141
rect 12835 91 12898 125
rect 12932 91 12995 125
rect 12801 75 12835 91
rect 12995 75 13029 91
rect 13109 125 13143 161
rect 13303 125 13337 161
rect 13143 91 13206 125
rect 13240 91 13303 125
rect 13109 75 13143 91
rect 13303 75 13337 91
rect 13434 239 13502 279
rect 13434 205 13451 239
rect 13485 205 13502 239
rect 13434 165 13502 205
rect 13434 131 13451 165
rect 13485 131 13502 165
rect 13434 91 13502 131
rect 13434 57 13451 91
rect 13485 57 13502 91
rect 13569 335 13603 351
rect 13763 335 13797 351
rect 13957 335 13991 351
rect 13603 301 13666 335
rect 13700 301 13763 335
rect 13797 301 13860 335
rect 13894 301 13957 335
rect 13569 263 13603 301
rect 13569 195 13603 229
rect 13763 263 13797 301
rect 13957 285 13991 301
rect 14071 335 14105 351
rect 14265 350 14299 501
rect 14071 263 14105 301
rect 13569 125 13603 161
rect 13569 75 13603 91
rect 13666 210 13700 226
rect 13434 34 13502 57
rect 13666 34 13700 176
rect 13763 195 13797 229
rect 13861 216 13895 232
rect 14071 216 14105 229
rect 13895 195 14105 216
rect 13895 182 14071 195
rect 13861 166 13895 182
rect 13763 125 13797 161
rect 14168 316 14299 350
rect 14396 461 14464 544
rect 14396 427 14413 461
rect 14447 427 14464 461
rect 14396 387 14464 427
rect 14396 353 14413 387
rect 14447 353 14464 387
rect 14635 535 14669 923
rect 14635 433 14669 501
rect 14635 383 14669 399
rect 14857 957 14891 973
rect 14857 905 14891 923
rect 14857 433 14891 871
rect 14857 383 14891 399
rect 15079 957 15113 973
rect 15079 461 15113 923
rect 15079 383 15113 399
rect 15227 757 15261 1014
rect 15358 1019 15375 1053
rect 15409 1019 15426 1053
rect 15593 1366 15627 1446
rect 15593 1298 15627 1332
rect 15593 1230 15627 1264
rect 15593 1162 15627 1196
rect 15593 1093 15627 1128
rect 15593 1043 15627 1059
rect 15681 1366 15715 1404
rect 15681 1298 15715 1332
rect 15681 1230 15715 1264
rect 15681 1162 15715 1196
rect 15681 1093 15715 1128
rect 15769 1366 15803 1446
rect 15769 1298 15803 1332
rect 15769 1230 15803 1264
rect 15769 1162 15803 1196
rect 15769 1111 15803 1128
rect 15857 1366 15891 1404
rect 15857 1298 15891 1332
rect 15857 1230 15891 1264
rect 15857 1162 15891 1196
rect 15681 1048 15715 1059
rect 15857 1093 15891 1128
rect 15945 1366 15979 1446
rect 15945 1298 15979 1332
rect 15945 1230 15979 1264
rect 15945 1162 15979 1196
rect 15945 1111 15979 1128
rect 16033 1366 16067 1404
rect 16033 1298 16067 1332
rect 16033 1230 16067 1264
rect 16033 1162 16067 1196
rect 15857 1048 15891 1059
rect 16033 1093 16067 1128
rect 16121 1366 16155 1446
rect 16121 1298 16155 1332
rect 16121 1230 16155 1264
rect 16121 1162 16155 1196
rect 16121 1111 16155 1128
rect 16320 1423 16388 1446
rect 16320 1389 16337 1423
rect 16371 1389 16388 1423
rect 16320 1349 16388 1389
rect 16320 1315 16337 1349
rect 16371 1315 16388 1349
rect 16320 1275 16388 1315
rect 16320 1241 16337 1275
rect 16371 1241 16388 1275
rect 16320 1201 16388 1241
rect 16320 1167 16337 1201
rect 16371 1167 16388 1201
rect 16320 1127 16388 1167
rect 16033 1048 16067 1059
rect 16320 1093 16337 1127
rect 16371 1093 16388 1127
rect 16320 1053 16388 1093
rect 15358 979 15426 1019
rect 15681 1014 16223 1048
rect 15358 945 15375 979
rect 15409 945 15426 979
rect 15358 905 15426 945
rect 15358 871 15375 905
rect 15409 871 15426 905
rect 15358 822 15426 871
rect 15597 957 15631 973
rect 14168 219 14202 316
rect 14396 313 14464 353
rect 14396 279 14413 313
rect 14447 279 14464 313
rect 14168 169 14202 185
rect 14265 263 14299 279
rect 14265 195 14299 229
rect 13957 125 13991 141
rect 13797 91 13860 125
rect 13894 91 13957 125
rect 13763 75 13797 91
rect 13957 75 13991 91
rect 14071 125 14105 161
rect 14265 125 14299 161
rect 14105 91 14168 125
rect 14202 91 14265 125
rect 14071 75 14105 91
rect 14265 75 14299 91
rect 14396 239 14464 279
rect 14396 205 14413 239
rect 14447 205 14464 239
rect 14396 165 14464 205
rect 14396 131 14413 165
rect 14447 131 14464 165
rect 14396 91 14464 131
rect 14396 57 14413 91
rect 14447 57 14464 91
rect 14531 335 14565 351
rect 14725 335 14759 351
rect 14919 335 14953 351
rect 14565 301 14628 335
rect 14662 301 14725 335
rect 14759 301 14822 335
rect 14856 301 14919 335
rect 14531 263 14565 301
rect 14531 195 14565 229
rect 14725 263 14759 301
rect 14919 285 14953 301
rect 15033 335 15067 351
rect 15227 350 15261 723
rect 15597 683 15631 923
rect 15033 263 15067 301
rect 14531 125 14565 161
rect 14531 75 14565 91
rect 14628 210 14662 226
rect 14396 34 14464 57
rect 14628 34 14662 176
rect 14725 195 14759 229
rect 14823 216 14857 232
rect 15033 216 15067 229
rect 14857 195 15067 216
rect 14857 182 15033 195
rect 14823 166 14857 182
rect 14725 125 14759 161
rect 15130 316 15261 350
rect 15358 461 15426 544
rect 15358 427 15375 461
rect 15409 427 15426 461
rect 15358 387 15426 427
rect 15358 353 15375 387
rect 15409 353 15426 387
rect 15597 433 15631 649
rect 15597 383 15631 399
rect 15819 957 15853 973
rect 15819 461 15853 923
rect 15819 383 15853 399
rect 16041 957 16075 973
rect 16041 535 16075 923
rect 16041 433 16075 501
rect 16041 383 16075 399
rect 16189 461 16223 1014
rect 16320 1019 16337 1053
rect 16371 1019 16388 1053
rect 16555 1366 16589 1446
rect 16555 1298 16589 1332
rect 16555 1230 16589 1264
rect 16555 1162 16589 1196
rect 16555 1093 16589 1128
rect 16555 1043 16589 1059
rect 16643 1366 16677 1404
rect 16643 1298 16677 1332
rect 16643 1230 16677 1264
rect 16643 1162 16677 1196
rect 16643 1093 16677 1128
rect 16731 1366 16765 1446
rect 16731 1298 16765 1332
rect 16731 1230 16765 1264
rect 16731 1162 16765 1196
rect 16731 1111 16765 1128
rect 16819 1366 16853 1404
rect 16819 1298 16853 1332
rect 16819 1230 16853 1264
rect 16819 1162 16853 1196
rect 16643 1048 16677 1059
rect 16819 1093 16853 1128
rect 16907 1366 16941 1446
rect 16907 1298 16941 1332
rect 16907 1230 16941 1264
rect 16907 1162 16941 1196
rect 16907 1111 16941 1128
rect 16995 1366 17029 1404
rect 16995 1298 17029 1332
rect 16995 1230 17029 1264
rect 16995 1162 17029 1196
rect 16819 1048 16853 1059
rect 16995 1093 17029 1128
rect 17083 1366 17117 1446
rect 17083 1298 17117 1332
rect 17083 1230 17117 1264
rect 17083 1162 17117 1196
rect 17083 1111 17117 1128
rect 17282 1423 17350 1446
rect 17282 1389 17299 1423
rect 17333 1389 17350 1423
rect 17282 1349 17350 1389
rect 17282 1315 17299 1349
rect 17333 1315 17350 1349
rect 17282 1275 17350 1315
rect 17282 1241 17299 1275
rect 17333 1241 17350 1275
rect 17282 1201 17350 1241
rect 17282 1167 17299 1201
rect 17333 1167 17350 1201
rect 17282 1127 17350 1167
rect 16995 1048 17029 1059
rect 17282 1093 17299 1127
rect 17333 1093 17350 1127
rect 17282 1053 17350 1093
rect 16320 979 16388 1019
rect 16643 1014 17185 1048
rect 16320 945 16337 979
rect 16371 945 16388 979
rect 16320 905 16388 945
rect 16320 871 16337 905
rect 16371 871 16388 905
rect 16320 822 16388 871
rect 16559 957 16593 973
rect 15130 219 15164 316
rect 15358 313 15426 353
rect 15358 279 15375 313
rect 15409 279 15426 313
rect 15130 169 15164 185
rect 15227 263 15261 279
rect 15227 195 15261 229
rect 14919 125 14953 141
rect 14759 91 14822 125
rect 14856 91 14919 125
rect 14725 75 14759 91
rect 14919 75 14953 91
rect 15033 125 15067 161
rect 15227 125 15261 161
rect 15067 91 15130 125
rect 15164 91 15227 125
rect 15033 75 15067 91
rect 15227 75 15261 91
rect 15358 239 15426 279
rect 15358 205 15375 239
rect 15409 205 15426 239
rect 15358 165 15426 205
rect 15358 131 15375 165
rect 15409 131 15426 165
rect 15358 91 15426 131
rect 15358 57 15375 91
rect 15409 57 15426 91
rect 15493 335 15527 351
rect 15687 335 15721 351
rect 15881 335 15915 351
rect 15527 301 15590 335
rect 15624 301 15687 335
rect 15721 301 15784 335
rect 15818 301 15881 335
rect 15493 263 15527 301
rect 15493 195 15527 229
rect 15687 263 15721 301
rect 15881 285 15915 301
rect 15995 335 16029 351
rect 16189 350 16223 427
rect 15995 263 16029 301
rect 15493 125 15527 161
rect 15493 75 15527 91
rect 15590 210 15624 226
rect 15358 34 15426 57
rect 15590 34 15624 176
rect 15687 195 15721 229
rect 15785 216 15819 232
rect 15995 216 16029 229
rect 15819 195 16029 216
rect 15819 182 15995 195
rect 15785 166 15819 182
rect 15687 125 15721 161
rect 16092 316 16223 350
rect 16320 461 16388 544
rect 16320 427 16337 461
rect 16371 427 16388 461
rect 16320 387 16388 427
rect 16320 353 16337 387
rect 16371 353 16388 387
rect 16559 461 16593 923
rect 16559 383 16593 399
rect 16781 957 16815 973
rect 16781 609 16815 923
rect 16781 433 16815 575
rect 16781 383 16815 399
rect 17003 957 17037 973
rect 17003 757 17037 923
rect 17003 433 17037 723
rect 17003 383 17037 399
rect 17151 535 17185 1014
rect 17282 1019 17299 1053
rect 17333 1019 17350 1053
rect 17457 1365 17491 1446
rect 17457 1297 17491 1331
rect 17457 1229 17491 1263
rect 17457 1161 17491 1195
rect 17457 1093 17491 1127
rect 17457 1025 17491 1059
rect 17545 1365 17581 1399
rect 17633 1365 17667 1446
rect 17545 1297 17579 1331
rect 17545 1229 17579 1263
rect 17545 1161 17579 1195
rect 17545 1093 17579 1127
rect 17633 1297 17667 1331
rect 17633 1229 17667 1263
rect 17633 1161 17667 1195
rect 17633 1111 17667 1127
rect 17721 1365 17755 1399
rect 17721 1297 17755 1331
rect 17721 1229 17755 1263
rect 17721 1161 17755 1195
rect 17721 1059 17755 1127
rect 17545 1025 17721 1059
rect 17809 1365 17843 1446
rect 17809 1297 17843 1331
rect 17809 1229 17843 1263
rect 17809 1161 17843 1195
rect 17809 1093 17843 1127
rect 17809 1025 17843 1059
rect 17948 1423 18016 1446
rect 17948 1389 17965 1423
rect 17999 1389 18016 1423
rect 18614 1423 18682 1446
rect 17948 1349 18016 1389
rect 17948 1315 17965 1349
rect 17999 1315 18016 1349
rect 17948 1275 18016 1315
rect 17948 1241 17965 1275
rect 17999 1241 18016 1275
rect 17948 1201 18016 1241
rect 17948 1167 17965 1201
rect 17999 1167 18016 1201
rect 17948 1127 18016 1167
rect 17948 1093 17965 1127
rect 17999 1093 18016 1127
rect 17948 1053 18016 1093
rect 17282 979 17350 1019
rect 17721 1009 17755 1025
rect 17948 1019 17965 1053
rect 17999 1019 18016 1053
rect 17282 945 17299 979
rect 17333 945 17350 979
rect 17948 979 18016 1019
rect 18121 1365 18507 1399
rect 18121 1297 18155 1331
rect 18121 1229 18155 1263
rect 18121 1161 18155 1195
rect 18121 1059 18155 1127
rect 18209 1297 18243 1313
rect 18209 1229 18243 1263
rect 18209 1161 18243 1195
rect 18209 1093 18243 1127
rect 18297 1297 18331 1331
rect 18297 1229 18331 1263
rect 18297 1161 18331 1195
rect 18297 1111 18331 1127
rect 18385 1297 18419 1313
rect 18385 1229 18419 1263
rect 18385 1161 18419 1195
rect 18385 1059 18419 1127
rect 18473 1297 18507 1331
rect 18473 1229 18507 1263
rect 18473 1161 18507 1195
rect 18473 1075 18507 1127
rect 18614 1389 18631 1423
rect 18665 1389 18682 1423
rect 19280 1423 19348 1446
rect 18614 1349 18682 1389
rect 18614 1315 18631 1349
rect 18665 1315 18682 1349
rect 18614 1275 18682 1315
rect 18614 1241 18631 1275
rect 18665 1241 18682 1275
rect 18614 1201 18682 1241
rect 18614 1167 18631 1201
rect 18665 1167 18682 1201
rect 18614 1127 18682 1167
rect 18614 1093 18631 1127
rect 18665 1093 18682 1127
rect 18209 1025 18385 1059
rect 18121 1009 18155 1025
rect 18385 1009 18419 1025
rect 18614 1053 18682 1093
rect 18614 1019 18631 1053
rect 18665 1019 18682 1053
rect 17282 905 17350 945
rect 17282 871 17299 905
rect 17333 871 17350 905
rect 17282 822 17350 871
rect 17447 958 17481 974
rect 17677 958 17711 974
rect 17447 905 17481 924
rect 16092 219 16126 316
rect 16320 313 16388 353
rect 16320 279 16337 313
rect 16371 279 16388 313
rect 16092 169 16126 185
rect 16189 263 16223 279
rect 16189 195 16223 229
rect 15881 125 15915 141
rect 15721 91 15784 125
rect 15818 91 15881 125
rect 15687 75 15721 91
rect 15881 75 15915 91
rect 15995 125 16029 161
rect 16189 125 16223 161
rect 16029 91 16092 125
rect 16126 91 16189 125
rect 15995 75 16029 91
rect 16189 75 16223 91
rect 16320 239 16388 279
rect 16320 205 16337 239
rect 16371 205 16388 239
rect 16320 165 16388 205
rect 16320 131 16337 165
rect 16371 131 16388 165
rect 16320 91 16388 131
rect 16320 57 16337 91
rect 16371 57 16388 91
rect 16455 335 16489 351
rect 16649 335 16683 351
rect 16843 335 16877 351
rect 16489 301 16552 335
rect 16586 301 16649 335
rect 16683 301 16746 335
rect 16780 301 16843 335
rect 16455 263 16489 301
rect 16455 195 16489 229
rect 16649 263 16683 301
rect 16843 285 16877 301
rect 16957 335 16991 351
rect 17151 350 17185 501
rect 16957 263 16991 301
rect 16455 125 16489 161
rect 16455 75 16489 91
rect 16552 210 16586 226
rect 16320 34 16388 57
rect 16552 34 16586 176
rect 16649 195 16683 229
rect 16747 216 16781 232
rect 16957 216 16991 229
rect 16781 195 16991 216
rect 16781 182 16957 195
rect 16747 166 16781 182
rect 16649 125 16683 161
rect 17054 316 17185 350
rect 17282 461 17350 544
rect 17282 427 17299 461
rect 17333 427 17350 461
rect 17282 387 17350 427
rect 17282 353 17299 387
rect 17333 353 17350 387
rect 17447 433 17481 871
rect 17447 383 17481 399
rect 17669 924 17677 942
rect 17669 908 17711 924
rect 17948 945 17965 979
rect 17999 945 18016 979
rect 18614 979 18682 1019
rect 18789 1365 19175 1399
rect 18789 1297 18823 1331
rect 18789 1229 18823 1263
rect 18789 1161 18823 1195
rect 18789 1059 18823 1127
rect 18877 1297 18911 1313
rect 18877 1229 18911 1263
rect 18877 1161 18911 1195
rect 18877 1093 18911 1127
rect 18965 1297 18999 1331
rect 18965 1229 18999 1263
rect 18965 1161 18999 1195
rect 18965 1111 18999 1127
rect 19053 1297 19087 1313
rect 19053 1229 19087 1263
rect 19053 1161 19087 1195
rect 19053 1093 19087 1127
rect 19141 1297 19175 1331
rect 19141 1229 19175 1263
rect 19141 1161 19175 1195
rect 19141 1111 19175 1127
rect 19280 1389 19297 1423
rect 19331 1389 19348 1423
rect 19280 1349 19348 1389
rect 19280 1315 19297 1349
rect 19331 1315 19348 1349
rect 19280 1275 19348 1315
rect 19280 1241 19297 1275
rect 19331 1241 19348 1275
rect 19280 1201 19348 1241
rect 19280 1167 19297 1201
rect 19331 1167 19348 1201
rect 19280 1127 19348 1167
rect 19280 1093 19297 1127
rect 19331 1093 19348 1127
rect 18877 1025 19183 1059
rect 18789 1009 18823 1025
rect 17669 831 17703 908
rect 17948 905 18016 945
rect 17948 871 17965 905
rect 17999 871 18016 905
rect 17948 822 18016 871
rect 18187 958 18221 974
rect 18187 905 18221 924
rect 17669 433 17703 797
rect 17669 383 17703 399
rect 17948 461 18016 544
rect 17948 427 17965 461
rect 17999 427 18016 461
rect 17948 387 18016 427
rect 17054 219 17088 316
rect 17282 313 17350 353
rect 17948 353 17965 387
rect 17999 353 18016 387
rect 18187 433 18221 871
rect 18187 383 18221 399
rect 18483 958 18517 974
rect 18483 433 18517 924
rect 18614 945 18631 979
rect 18665 945 18682 979
rect 18614 905 18682 945
rect 18614 871 18631 905
rect 18665 871 18682 905
rect 18614 822 18682 871
rect 18779 958 18813 974
rect 18483 383 18517 399
rect 18614 461 18682 544
rect 18614 427 18631 461
rect 18665 427 18682 461
rect 18614 387 18682 427
rect 17282 279 17299 313
rect 17333 279 17350 313
rect 17054 169 17088 185
rect 17151 263 17185 279
rect 17151 195 17185 229
rect 16843 125 16877 141
rect 16683 91 16746 125
rect 16780 91 16843 125
rect 16649 75 16683 91
rect 16843 75 16877 91
rect 16957 125 16991 161
rect 17151 125 17185 161
rect 16991 91 17054 125
rect 17088 91 17151 125
rect 16957 75 16991 91
rect 17151 75 17185 91
rect 17282 239 17350 279
rect 17282 205 17299 239
rect 17333 205 17350 239
rect 17282 165 17350 205
rect 17282 131 17299 165
rect 17333 131 17350 165
rect 17282 91 17350 131
rect 17282 57 17299 91
rect 17333 57 17350 91
rect 17438 333 17472 349
rect 17632 333 17666 349
rect 17472 299 17535 333
rect 17569 299 17632 333
rect 17438 261 17472 299
rect 17438 193 17472 227
rect 17632 261 17666 299
rect 17826 333 17860 349
rect 17729 253 17763 269
rect 17438 123 17472 159
rect 17438 73 17472 89
rect 17535 208 17569 224
rect 17282 34 17350 57
rect 17535 34 17569 174
rect 17632 193 17666 227
rect 17728 219 17729 234
rect 17728 217 17763 219
rect 17762 203 17763 217
rect 17826 261 17860 299
rect 17728 167 17762 183
rect 17826 193 17860 227
rect 17632 123 17666 159
rect 17826 123 17860 159
rect 17666 89 17728 123
rect 17762 89 17826 123
rect 17632 73 17666 89
rect 17826 73 17860 89
rect 17948 313 18016 353
rect 18614 353 18631 387
rect 18665 353 18682 387
rect 18779 433 18813 924
rect 18779 383 18813 399
rect 19001 958 19039 974
rect 19001 924 19005 958
rect 19001 908 19039 924
rect 19001 831 19035 908
rect 19001 433 19035 797
rect 19001 383 19035 399
rect 19149 831 19183 1025
rect 19280 1053 19348 1093
rect 19280 1019 19297 1053
rect 19331 1019 19348 1053
rect 19280 979 19348 1019
rect 19280 945 19297 979
rect 19331 945 19348 979
rect 19280 905 19348 945
rect 19280 871 19297 905
rect 19331 871 19348 905
rect 19280 822 19348 871
rect 17948 279 17965 313
rect 17999 279 18016 313
rect 17948 239 18016 279
rect 17948 205 17965 239
rect 17999 205 18016 239
rect 17948 165 18016 205
rect 17948 131 17965 165
rect 17999 131 18016 165
rect 17948 91 18016 131
rect 17948 57 17965 91
rect 17999 57 18016 91
rect 18104 333 18138 349
rect 18298 333 18332 349
rect 18138 299 18201 333
rect 18235 299 18298 333
rect 18104 261 18138 299
rect 18104 193 18138 227
rect 18298 261 18332 299
rect 18492 333 18526 349
rect 18104 123 18138 159
rect 18104 73 18138 89
rect 18201 208 18235 224
rect 17948 34 18016 57
rect 18201 34 18235 174
rect 18298 193 18332 227
rect 18395 253 18429 269
rect 18395 217 18429 219
rect 18395 167 18429 183
rect 18492 261 18526 299
rect 18492 193 18526 227
rect 18298 123 18332 159
rect 18492 123 18526 159
rect 18332 89 18395 123
rect 18429 89 18492 123
rect 18298 73 18332 89
rect 18492 73 18526 89
rect 18614 313 18682 353
rect 18614 279 18631 313
rect 18665 279 18682 313
rect 18614 239 18682 279
rect 18614 205 18631 239
rect 18665 205 18682 239
rect 18614 165 18682 205
rect 18614 131 18631 165
rect 18665 131 18682 165
rect 18614 91 18682 131
rect 18614 57 18631 91
rect 18665 57 18682 91
rect 18770 333 18804 349
rect 18964 333 18998 349
rect 19149 346 19183 797
rect 18804 299 18867 333
rect 18901 299 18964 333
rect 18770 261 18804 299
rect 18770 193 18804 227
rect 18964 261 18998 299
rect 18770 123 18804 159
rect 18770 73 18804 89
rect 18867 208 18901 224
rect 18614 34 18682 57
rect 18867 34 18901 174
rect 18964 193 18998 227
rect 19061 312 19183 346
rect 19280 461 19348 544
rect 19280 427 19297 461
rect 19331 427 19348 461
rect 19280 387 19348 427
rect 19280 353 19297 387
rect 19331 353 19348 387
rect 19280 313 19348 353
rect 19061 253 19095 312
rect 19280 279 19297 313
rect 19331 279 19348 313
rect 19061 217 19095 219
rect 19061 167 19095 183
rect 19158 261 19192 278
rect 19158 193 19192 227
rect 18964 123 18998 159
rect 19158 123 19192 159
rect 18998 89 19061 123
rect 19095 89 19158 123
rect 18964 73 18998 89
rect 19158 73 19192 89
rect 19280 239 19348 279
rect 19280 205 19297 239
rect 19331 205 19348 239
rect 19280 165 19348 205
rect 19280 131 19297 165
rect 19331 131 19348 165
rect 19280 91 19348 131
rect 19280 57 19297 91
rect 19331 57 19348 91
rect 19280 34 19348 57
rect -34 17 19348 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6569 17
rect 6603 -17 6643 17
rect 6677 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7753 17
rect 7787 -17 7827 17
rect 7861 -17 7901 17
rect 7935 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8123 17
rect 8157 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8567 17
rect 8601 -17 8715 17
rect 8749 -17 8789 17
rect 8823 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9529 17
rect 9563 -17 9677 17
rect 9711 -17 9751 17
rect 9785 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10195 17
rect 10229 -17 10269 17
rect 10303 -17 10343 17
rect 10377 -17 10417 17
rect 10451 -17 10491 17
rect 10525 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10861 17
rect 10895 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11305 17
rect 11339 -17 11379 17
rect 11413 -17 11453 17
rect 11487 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12193 17
rect 12227 -17 12267 17
rect 12301 -17 12341 17
rect 12375 -17 12415 17
rect 12449 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12859 17
rect 12893 -17 12933 17
rect 12967 -17 13007 17
rect 13041 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13525 17
rect 13559 -17 13599 17
rect 13633 -17 13673 17
rect 13707 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13895 17
rect 13929 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14191 17
rect 14225 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14635 17
rect 14669 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14857 17
rect 14891 -17 14931 17
rect 14965 -17 15005 17
rect 15039 -17 15079 17
rect 15113 -17 15153 17
rect 15187 -17 15227 17
rect 15261 -17 15301 17
rect 15335 -17 15449 17
rect 15483 -17 15523 17
rect 15557 -17 15597 17
rect 15631 -17 15671 17
rect 15705 -17 15745 17
rect 15779 -17 15819 17
rect 15853 -17 15893 17
rect 15927 -17 15967 17
rect 16001 -17 16041 17
rect 16075 -17 16115 17
rect 16149 -17 16189 17
rect 16223 -17 16263 17
rect 16297 -17 16411 17
rect 16445 -17 16485 17
rect 16519 -17 16559 17
rect 16593 -17 16633 17
rect 16667 -17 16707 17
rect 16741 -17 16781 17
rect 16815 -17 16855 17
rect 16889 -17 16929 17
rect 16963 -17 17003 17
rect 17037 -17 17077 17
rect 17111 -17 17151 17
rect 17185 -17 17225 17
rect 17259 -17 17373 17
rect 17407 -17 17447 17
rect 17481 -17 17521 17
rect 17555 -17 17595 17
rect 17629 -17 17669 17
rect 17703 -17 17743 17
rect 17777 -17 17817 17
rect 17851 -17 17891 17
rect 17925 -17 18039 17
rect 18073 -17 18113 17
rect 18147 -17 18187 17
rect 18221 -17 18261 17
rect 18295 -17 18335 17
rect 18369 -17 18409 17
rect 18443 -17 18483 17
rect 18517 -17 18557 17
rect 18591 -17 18705 17
rect 18739 -17 18779 17
rect 18813 -17 18853 17
rect 18887 -17 18927 17
rect 18961 -17 19001 17
rect 19035 -17 19075 17
rect 19109 -17 19149 17
rect 19183 -17 19223 17
rect 19257 -17 19348 17
rect -34 -34 19348 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5163 1463 5197 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5533 1463 5567 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5829 1463 5863 1497
rect 5903 1463 5937 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6125 1463 6159 1497
rect 6199 1463 6233 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6495 1463 6529 1497
rect 6569 1463 6603 1497
rect 6643 1463 6677 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7087 1463 7121 1497
rect 7161 1463 7195 1497
rect 7235 1463 7269 1497
rect 7309 1463 7343 1497
rect 7383 1463 7417 1497
rect 7457 1463 7491 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7753 1463 7787 1497
rect 7827 1463 7861 1497
rect 7901 1463 7935 1497
rect 7975 1463 8009 1497
rect 8049 1463 8083 1497
rect 8123 1463 8157 1497
rect 8197 1463 8231 1497
rect 8271 1463 8305 1497
rect 8345 1463 8379 1497
rect 8419 1463 8453 1497
rect 8493 1463 8527 1497
rect 8567 1463 8601 1497
rect 8715 1463 8749 1497
rect 8789 1463 8823 1497
rect 8863 1463 8897 1497
rect 8937 1463 8971 1497
rect 9011 1463 9045 1497
rect 9085 1463 9119 1497
rect 9159 1463 9193 1497
rect 9233 1463 9267 1497
rect 9307 1463 9341 1497
rect 9381 1463 9415 1497
rect 9455 1463 9489 1497
rect 9529 1463 9563 1497
rect 9677 1463 9711 1497
rect 9751 1463 9785 1497
rect 9825 1463 9859 1497
rect 9899 1463 9933 1497
rect 9973 1463 10007 1497
rect 10047 1463 10081 1497
rect 10121 1463 10155 1497
rect 10195 1463 10229 1497
rect 10269 1463 10303 1497
rect 10343 1463 10377 1497
rect 10417 1463 10451 1497
rect 10491 1463 10525 1497
rect 10639 1463 10673 1497
rect 10713 1463 10747 1497
rect 10787 1463 10821 1497
rect 10861 1463 10895 1497
rect 10935 1463 10969 1497
rect 11009 1463 11043 1497
rect 11083 1463 11117 1497
rect 11157 1463 11191 1497
rect 11231 1463 11265 1497
rect 11305 1463 11339 1497
rect 11379 1463 11413 1497
rect 11453 1463 11487 1497
rect 11601 1463 11635 1497
rect 11675 1463 11709 1497
rect 11749 1463 11783 1497
rect 11823 1463 11857 1497
rect 11897 1463 11931 1497
rect 11971 1463 12005 1497
rect 12045 1463 12079 1497
rect 12119 1463 12153 1497
rect 12193 1463 12227 1497
rect 12267 1463 12301 1497
rect 12341 1463 12375 1497
rect 12415 1463 12449 1497
rect 12563 1463 12597 1497
rect 12637 1463 12671 1497
rect 12711 1463 12745 1497
rect 12785 1463 12819 1497
rect 12859 1463 12893 1497
rect 12933 1463 12967 1497
rect 13007 1463 13041 1497
rect 13081 1463 13115 1497
rect 13155 1463 13189 1497
rect 13229 1463 13263 1497
rect 13303 1463 13337 1497
rect 13377 1463 13411 1497
rect 13525 1463 13559 1497
rect 13599 1463 13633 1497
rect 13673 1463 13707 1497
rect 13747 1463 13781 1497
rect 13821 1463 13855 1497
rect 13895 1463 13929 1497
rect 13969 1463 14003 1497
rect 14043 1463 14077 1497
rect 14117 1463 14151 1497
rect 14191 1463 14225 1497
rect 14265 1463 14299 1497
rect 14339 1463 14373 1497
rect 14487 1463 14521 1497
rect 14561 1463 14595 1497
rect 14635 1463 14669 1497
rect 14709 1463 14743 1497
rect 14783 1463 14817 1497
rect 14857 1463 14891 1497
rect 14931 1463 14965 1497
rect 15005 1463 15039 1497
rect 15079 1463 15113 1497
rect 15153 1463 15187 1497
rect 15227 1463 15261 1497
rect 15301 1463 15335 1497
rect 15449 1463 15483 1497
rect 15523 1463 15557 1497
rect 15597 1463 15631 1497
rect 15671 1463 15705 1497
rect 15745 1463 15779 1497
rect 15819 1463 15853 1497
rect 15893 1463 15927 1497
rect 15967 1463 16001 1497
rect 16041 1463 16075 1497
rect 16115 1463 16149 1497
rect 16189 1463 16223 1497
rect 16263 1463 16297 1497
rect 16411 1463 16445 1497
rect 16485 1463 16519 1497
rect 16559 1463 16593 1497
rect 16633 1463 16667 1497
rect 16707 1463 16741 1497
rect 16781 1463 16815 1497
rect 16855 1463 16889 1497
rect 16929 1463 16963 1497
rect 17003 1463 17037 1497
rect 17077 1463 17111 1497
rect 17151 1463 17185 1497
rect 17225 1463 17259 1497
rect 17373 1463 17407 1497
rect 17447 1463 17481 1497
rect 17521 1463 17555 1497
rect 17595 1463 17629 1497
rect 17669 1463 17703 1497
rect 17743 1463 17777 1497
rect 17817 1463 17851 1497
rect 17891 1463 17925 1497
rect 18039 1463 18073 1497
rect 18113 1463 18147 1497
rect 18187 1463 18221 1497
rect 18261 1463 18295 1497
rect 18335 1463 18369 1497
rect 18409 1463 18443 1497
rect 18483 1463 18517 1497
rect 18557 1463 18591 1497
rect 18705 1463 18739 1497
rect 18779 1463 18813 1497
rect 18853 1463 18887 1497
rect 18927 1463 18961 1497
rect 19001 1463 19035 1497
rect 19075 1463 19109 1497
rect 19149 1463 19183 1497
rect 19223 1463 19257 1497
rect 205 797 239 831
rect 427 433 461 461
rect 427 427 461 433
rect 649 649 683 683
rect 797 501 831 535
rect 1167 501 1201 535
rect 1389 871 1423 905
rect 1611 723 1645 757
rect 1759 649 1793 683
rect 2129 501 2163 535
rect 2351 575 2385 609
rect 2573 723 2607 757
rect 2721 501 2755 535
rect 3091 501 3125 535
rect 3313 871 3347 905
rect 3535 433 3569 461
rect 3535 427 3569 433
rect 3683 723 3717 757
rect 4053 649 4087 683
rect 4275 433 4309 461
rect 4275 427 4309 433
rect 4497 649 4531 683
rect 4645 945 4679 979
rect 4645 501 4679 535
rect 5015 501 5049 535
rect 5237 575 5271 609
rect 5459 723 5493 757
rect 5607 649 5641 683
rect 5977 797 6011 831
rect 6199 433 6233 461
rect 6199 427 6233 433
rect 6421 649 6455 683
rect 6569 501 6603 535
rect 6939 501 6973 535
rect 7161 871 7195 905
rect 7383 723 7417 757
rect 7531 649 7565 683
rect 7901 501 7935 535
rect 8123 575 8157 609
rect 8345 723 8379 757
rect 8493 501 8527 535
rect 8863 501 8897 535
rect 9085 871 9119 905
rect 9307 433 9341 461
rect 9307 427 9341 433
rect 9455 723 9489 757
rect 9825 649 9859 683
rect 10047 433 10081 461
rect 10047 427 10081 433
rect 10269 501 10303 535
rect 10417 649 10451 683
rect 10787 649 10821 683
rect 11009 575 11043 609
rect 11231 723 11265 757
rect 11749 797 11783 831
rect 11379 501 11413 535
rect 11971 433 12005 461
rect 11971 427 12005 433
rect 12193 649 12227 683
rect 12341 501 12375 535
rect 12711 501 12745 535
rect 12933 871 12967 905
rect 13155 723 13189 757
rect 13303 649 13337 683
rect 13673 501 13707 535
rect 13895 575 13929 609
rect 14117 723 14151 757
rect 14265 501 14299 535
rect 14635 501 14669 535
rect 14857 871 14891 905
rect 15079 433 15113 461
rect 15079 427 15113 433
rect 15227 723 15261 757
rect 15597 649 15631 683
rect 15819 433 15853 461
rect 15819 427 15853 433
rect 16041 501 16075 535
rect 16189 427 16223 461
rect 16559 433 16593 461
rect 16559 427 16593 433
rect 16781 575 16815 609
rect 17003 723 17037 757
rect 17721 1025 17755 1059
rect 18121 1025 18155 1059
rect 18385 1025 18419 1059
rect 17447 871 17481 905
rect 17151 501 17185 535
rect 18789 1025 18823 1059
rect 17669 797 17703 831
rect 18187 871 18221 905
rect 18483 399 18517 433
rect 17729 219 17763 253
rect 18779 399 18813 433
rect 19001 797 19035 831
rect 19149 797 19183 831
rect 18395 219 18429 253
rect 19061 219 19095 253
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5163 -17 5197 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5533 -17 5567 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5829 -17 5863 17
rect 5903 -17 5937 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6125 -17 6159 17
rect 6199 -17 6233 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6495 -17 6529 17
rect 6569 -17 6603 17
rect 6643 -17 6677 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7087 -17 7121 17
rect 7161 -17 7195 17
rect 7235 -17 7269 17
rect 7309 -17 7343 17
rect 7383 -17 7417 17
rect 7457 -17 7491 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7753 -17 7787 17
rect 7827 -17 7861 17
rect 7901 -17 7935 17
rect 7975 -17 8009 17
rect 8049 -17 8083 17
rect 8123 -17 8157 17
rect 8197 -17 8231 17
rect 8271 -17 8305 17
rect 8345 -17 8379 17
rect 8419 -17 8453 17
rect 8493 -17 8527 17
rect 8567 -17 8601 17
rect 8715 -17 8749 17
rect 8789 -17 8823 17
rect 8863 -17 8897 17
rect 8937 -17 8971 17
rect 9011 -17 9045 17
rect 9085 -17 9119 17
rect 9159 -17 9193 17
rect 9233 -17 9267 17
rect 9307 -17 9341 17
rect 9381 -17 9415 17
rect 9455 -17 9489 17
rect 9529 -17 9563 17
rect 9677 -17 9711 17
rect 9751 -17 9785 17
rect 9825 -17 9859 17
rect 9899 -17 9933 17
rect 9973 -17 10007 17
rect 10047 -17 10081 17
rect 10121 -17 10155 17
rect 10195 -17 10229 17
rect 10269 -17 10303 17
rect 10343 -17 10377 17
rect 10417 -17 10451 17
rect 10491 -17 10525 17
rect 10639 -17 10673 17
rect 10713 -17 10747 17
rect 10787 -17 10821 17
rect 10861 -17 10895 17
rect 10935 -17 10969 17
rect 11009 -17 11043 17
rect 11083 -17 11117 17
rect 11157 -17 11191 17
rect 11231 -17 11265 17
rect 11305 -17 11339 17
rect 11379 -17 11413 17
rect 11453 -17 11487 17
rect 11601 -17 11635 17
rect 11675 -17 11709 17
rect 11749 -17 11783 17
rect 11823 -17 11857 17
rect 11897 -17 11931 17
rect 11971 -17 12005 17
rect 12045 -17 12079 17
rect 12119 -17 12153 17
rect 12193 -17 12227 17
rect 12267 -17 12301 17
rect 12341 -17 12375 17
rect 12415 -17 12449 17
rect 12563 -17 12597 17
rect 12637 -17 12671 17
rect 12711 -17 12745 17
rect 12785 -17 12819 17
rect 12859 -17 12893 17
rect 12933 -17 12967 17
rect 13007 -17 13041 17
rect 13081 -17 13115 17
rect 13155 -17 13189 17
rect 13229 -17 13263 17
rect 13303 -17 13337 17
rect 13377 -17 13411 17
rect 13525 -17 13559 17
rect 13599 -17 13633 17
rect 13673 -17 13707 17
rect 13747 -17 13781 17
rect 13821 -17 13855 17
rect 13895 -17 13929 17
rect 13969 -17 14003 17
rect 14043 -17 14077 17
rect 14117 -17 14151 17
rect 14191 -17 14225 17
rect 14265 -17 14299 17
rect 14339 -17 14373 17
rect 14487 -17 14521 17
rect 14561 -17 14595 17
rect 14635 -17 14669 17
rect 14709 -17 14743 17
rect 14783 -17 14817 17
rect 14857 -17 14891 17
rect 14931 -17 14965 17
rect 15005 -17 15039 17
rect 15079 -17 15113 17
rect 15153 -17 15187 17
rect 15227 -17 15261 17
rect 15301 -17 15335 17
rect 15449 -17 15483 17
rect 15523 -17 15557 17
rect 15597 -17 15631 17
rect 15671 -17 15705 17
rect 15745 -17 15779 17
rect 15819 -17 15853 17
rect 15893 -17 15927 17
rect 15967 -17 16001 17
rect 16041 -17 16075 17
rect 16115 -17 16149 17
rect 16189 -17 16223 17
rect 16263 -17 16297 17
rect 16411 -17 16445 17
rect 16485 -17 16519 17
rect 16559 -17 16593 17
rect 16633 -17 16667 17
rect 16707 -17 16741 17
rect 16781 -17 16815 17
rect 16855 -17 16889 17
rect 16929 -17 16963 17
rect 17003 -17 17037 17
rect 17077 -17 17111 17
rect 17151 -17 17185 17
rect 17225 -17 17259 17
rect 17373 -17 17407 17
rect 17447 -17 17481 17
rect 17521 -17 17555 17
rect 17595 -17 17629 17
rect 17669 -17 17703 17
rect 17743 -17 17777 17
rect 17817 -17 17851 17
rect 17891 -17 17925 17
rect 18039 -17 18073 17
rect 18113 -17 18147 17
rect 18187 -17 18221 17
rect 18261 -17 18295 17
rect 18335 -17 18369 17
rect 18409 -17 18443 17
rect 18483 -17 18517 17
rect 18557 -17 18591 17
rect 18705 -17 18739 17
rect 18779 -17 18813 17
rect 18853 -17 18887 17
rect 18927 -17 18961 17
rect 19001 -17 19035 17
rect 19075 -17 19109 17
rect 19149 -17 19183 17
rect 19223 -17 19257 17
<< metal1 >>
rect -34 1497 19348 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6569 1497
rect 6603 1463 6643 1497
rect 6677 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7753 1497
rect 7787 1463 7827 1497
rect 7861 1463 7901 1497
rect 7935 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8123 1497
rect 8157 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8567 1497
rect 8601 1463 8715 1497
rect 8749 1463 8789 1497
rect 8823 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9529 1497
rect 9563 1463 9677 1497
rect 9711 1463 9751 1497
rect 9785 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10195 1497
rect 10229 1463 10269 1497
rect 10303 1463 10343 1497
rect 10377 1463 10417 1497
rect 10451 1463 10491 1497
rect 10525 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10861 1497
rect 10895 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11305 1497
rect 11339 1463 11379 1497
rect 11413 1463 11453 1497
rect 11487 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12193 1497
rect 12227 1463 12267 1497
rect 12301 1463 12341 1497
rect 12375 1463 12415 1497
rect 12449 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12859 1497
rect 12893 1463 12933 1497
rect 12967 1463 13007 1497
rect 13041 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13525 1497
rect 13559 1463 13599 1497
rect 13633 1463 13673 1497
rect 13707 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13895 1497
rect 13929 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14191 1497
rect 14225 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14635 1497
rect 14669 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14857 1497
rect 14891 1463 14931 1497
rect 14965 1463 15005 1497
rect 15039 1463 15079 1497
rect 15113 1463 15153 1497
rect 15187 1463 15227 1497
rect 15261 1463 15301 1497
rect 15335 1463 15449 1497
rect 15483 1463 15523 1497
rect 15557 1463 15597 1497
rect 15631 1463 15671 1497
rect 15705 1463 15745 1497
rect 15779 1463 15819 1497
rect 15853 1463 15893 1497
rect 15927 1463 15967 1497
rect 16001 1463 16041 1497
rect 16075 1463 16115 1497
rect 16149 1463 16189 1497
rect 16223 1463 16263 1497
rect 16297 1463 16411 1497
rect 16445 1463 16485 1497
rect 16519 1463 16559 1497
rect 16593 1463 16633 1497
rect 16667 1463 16707 1497
rect 16741 1463 16781 1497
rect 16815 1463 16855 1497
rect 16889 1463 16929 1497
rect 16963 1463 17003 1497
rect 17037 1463 17077 1497
rect 17111 1463 17151 1497
rect 17185 1463 17225 1497
rect 17259 1463 17373 1497
rect 17407 1463 17447 1497
rect 17481 1463 17521 1497
rect 17555 1463 17595 1497
rect 17629 1463 17669 1497
rect 17703 1463 17743 1497
rect 17777 1463 17817 1497
rect 17851 1463 17891 1497
rect 17925 1463 18039 1497
rect 18073 1463 18113 1497
rect 18147 1463 18187 1497
rect 18221 1463 18261 1497
rect 18295 1463 18335 1497
rect 18369 1463 18409 1497
rect 18443 1463 18483 1497
rect 18517 1463 18557 1497
rect 18591 1463 18705 1497
rect 18739 1463 18779 1497
rect 18813 1463 18853 1497
rect 18887 1463 18927 1497
rect 18961 1463 19001 1497
rect 19035 1463 19075 1497
rect 19109 1463 19149 1497
rect 19183 1463 19223 1497
rect 19257 1463 19348 1497
rect -34 1446 19348 1463
rect 17715 1059 17761 1065
rect 18115 1059 18161 1065
rect 18379 1059 18425 1065
rect 18783 1059 18829 1065
rect 17709 1025 17721 1059
rect 17755 1025 18121 1059
rect 18155 1025 18167 1059
rect 18373 1025 18385 1059
rect 18419 1025 18789 1059
rect 18823 1025 18835 1059
rect 17715 1019 17761 1025
rect 18115 1019 18161 1025
rect 18379 1019 18425 1025
rect 18783 1019 18829 1025
rect 4639 979 4685 985
rect 4633 945 4645 979
rect 4679 945 15039 979
rect 4639 939 4685 945
rect 1383 905 1429 911
rect 3307 905 3353 911
rect 7155 905 7201 911
rect 9079 905 9125 911
rect 12927 905 12973 911
rect 14851 905 14897 911
rect 15005 905 15039 945
rect 17441 905 17487 911
rect 18181 905 18227 911
rect 1377 871 1389 905
rect 1423 871 3313 905
rect 3347 871 7161 905
rect 7195 871 9085 905
rect 9119 871 12933 905
rect 12967 871 14857 905
rect 14891 871 14903 905
rect 15005 873 17447 905
rect 15021 871 17447 873
rect 17481 871 18187 905
rect 18221 871 18233 905
rect 1383 865 1429 871
rect 3307 865 3353 871
rect 7155 865 7201 871
rect 9079 865 9125 871
rect 12927 865 12973 871
rect 14851 865 14897 871
rect 17441 865 17487 871
rect 18181 865 18227 871
rect 199 831 245 837
rect 5971 831 6017 837
rect 11743 831 11789 837
rect 17663 831 17709 837
rect 18995 831 19041 837
rect 19143 831 19189 837
rect 169 797 205 831
rect 239 797 5977 831
rect 6011 797 11749 831
rect 11783 797 11795 831
rect 13007 797 17669 831
rect 17703 797 19001 831
rect 19035 797 19047 831
rect 19137 797 19149 831
rect 19183 797 19219 831
rect 199 791 245 797
rect 5971 791 6017 797
rect 11743 791 11789 797
rect 1605 757 1651 763
rect 2567 757 2613 763
rect 3677 757 3723 763
rect 5453 757 5499 763
rect 7377 757 7423 763
rect 8339 757 8385 763
rect 9449 757 9495 763
rect 11225 757 11271 763
rect 13007 757 13041 797
rect 17663 791 17709 797
rect 18995 791 19041 797
rect 19143 791 19189 797
rect 13149 757 13195 763
rect 14111 757 14157 763
rect 15221 757 15267 763
rect 16997 757 17043 763
rect 1599 723 1611 757
rect 1645 723 2573 757
rect 2607 723 3683 757
rect 3717 723 5459 757
rect 5493 723 5505 757
rect 7371 723 7383 757
rect 7417 723 8345 757
rect 8379 723 9455 757
rect 9489 723 11231 757
rect 11265 723 11277 757
rect 11379 723 13041 757
rect 13143 723 13155 757
rect 13189 723 14117 757
rect 14151 723 15227 757
rect 15261 723 17003 757
rect 17037 723 17049 757
rect 1605 717 1651 723
rect 2567 717 2613 723
rect 3677 717 3723 723
rect 5453 717 5499 723
rect 7377 717 7423 723
rect 8339 717 8385 723
rect 9449 717 9495 723
rect 11225 717 11271 723
rect 643 683 689 689
rect 1753 683 1799 689
rect 4047 683 4093 689
rect 4491 683 4537 689
rect 5601 683 5647 689
rect 6415 683 6461 689
rect 7525 683 7571 689
rect 9819 683 9865 689
rect 10411 683 10457 689
rect 10781 683 10827 689
rect 11379 683 11413 723
rect 13149 717 13195 723
rect 14111 717 14157 723
rect 15221 717 15267 723
rect 16997 717 17043 723
rect 12187 683 12233 689
rect 13297 683 13343 689
rect 15591 683 15637 689
rect 637 649 649 683
rect 683 649 1759 683
rect 1793 649 4053 683
rect 4087 649 4099 683
rect 4485 649 4497 683
rect 4531 649 5607 683
rect 5641 649 5653 683
rect 6409 649 6421 683
rect 6455 649 7531 683
rect 7565 649 9825 683
rect 9859 649 9871 683
rect 10405 649 10417 683
rect 10451 649 10787 683
rect 10821 649 11413 683
rect 12181 649 12193 683
rect 12227 649 13303 683
rect 13337 649 15597 683
rect 15631 649 15643 683
rect 643 643 689 649
rect 1753 643 1799 649
rect 4047 643 4093 649
rect 4491 643 4537 649
rect 5601 643 5647 649
rect 6415 643 6461 649
rect 7525 643 7571 649
rect 9819 643 9865 649
rect 10411 643 10457 649
rect 10781 643 10827 649
rect 12187 643 12233 649
rect 13297 643 13343 649
rect 15591 643 15637 649
rect 2345 609 2391 615
rect 5231 609 5277 615
rect 8117 609 8163 615
rect 11003 609 11049 615
rect 13889 609 13935 615
rect 16775 609 16821 615
rect 2339 575 2351 609
rect 2385 575 5237 609
rect 5271 575 8123 609
rect 8157 575 11009 609
rect 11043 575 13895 609
rect 13929 575 16781 609
rect 16815 575 16827 609
rect 2345 569 2391 575
rect 5231 569 5277 575
rect 8117 569 8163 575
rect 11003 569 11049 575
rect 13889 569 13935 575
rect 16775 569 16821 575
rect 791 535 837 541
rect 1161 535 1207 541
rect 2123 535 2169 541
rect 2715 535 2761 541
rect 3085 535 3131 541
rect 4639 535 4685 541
rect 5009 535 5055 541
rect 6563 535 6609 541
rect 6933 535 6979 541
rect 7895 535 7941 541
rect 8487 535 8533 541
rect 8857 535 8903 541
rect 10263 535 10309 541
rect 11373 535 11419 541
rect 12335 535 12381 541
rect 12705 535 12751 541
rect 13667 535 13713 541
rect 14259 535 14305 541
rect 14629 535 14675 541
rect 16035 535 16081 541
rect 17145 535 17191 541
rect 785 501 797 535
rect 831 501 1167 535
rect 1201 501 2129 535
rect 2163 501 2175 535
rect 2709 501 2721 535
rect 2755 501 3091 535
rect 3125 501 3137 535
rect 4633 501 4645 535
rect 4679 501 5015 535
rect 5049 501 5061 535
rect 6557 501 6569 535
rect 6603 501 6939 535
rect 6973 501 7901 535
rect 7935 501 7947 535
rect 8481 501 8493 535
rect 8527 501 8863 535
rect 8897 501 8909 535
rect 10257 501 10269 535
rect 10303 501 11379 535
rect 11413 501 11425 535
rect 12329 501 12341 535
rect 12375 501 12711 535
rect 12745 501 13673 535
rect 13707 501 13719 535
rect 14253 501 14265 535
rect 14299 501 14635 535
rect 14669 501 14681 535
rect 16029 501 16041 535
rect 16075 501 17151 535
rect 17185 501 17197 535
rect 791 495 837 501
rect 1161 495 1207 501
rect 2123 495 2169 501
rect 2715 495 2761 501
rect 3085 495 3131 501
rect 4639 495 4685 501
rect 5009 495 5055 501
rect 6563 495 6609 501
rect 6933 495 6979 501
rect 7895 495 7941 501
rect 8487 495 8533 501
rect 8857 495 8903 501
rect 10263 495 10309 501
rect 11373 495 11419 501
rect 12335 495 12381 501
rect 12705 495 12751 501
rect 13667 495 13713 501
rect 14259 495 14305 501
rect 14629 495 14675 501
rect 16035 495 16081 501
rect 17145 495 17191 501
rect 421 461 467 467
rect 3529 461 3575 467
rect 4269 461 4315 467
rect 6193 461 6239 467
rect 9301 461 9347 467
rect 10041 461 10087 467
rect 11965 461 12011 467
rect 15073 461 15119 467
rect 15813 461 15859 467
rect 16183 461 16229 467
rect 16553 461 16599 467
rect 415 427 427 461
rect 461 427 3535 461
rect 3569 427 4275 461
rect 4309 427 6199 461
rect 6233 427 9307 461
rect 9341 427 10047 461
rect 10081 427 11971 461
rect 12005 427 15079 461
rect 15113 427 15819 461
rect 15853 427 15865 461
rect 16177 427 16189 461
rect 16223 427 16559 461
rect 16593 433 18523 461
rect 18773 433 18819 439
rect 16593 427 18483 433
rect 421 421 467 427
rect 3529 421 3575 427
rect 4269 421 4315 427
rect 6193 421 6239 427
rect 9301 421 9347 427
rect 10041 421 10087 427
rect 11965 421 12011 427
rect 15073 421 15119 427
rect 15813 421 15859 427
rect 16183 421 16229 427
rect 16553 421 16599 427
rect 18471 399 18483 427
rect 18517 399 18779 433
rect 18813 399 18825 433
rect 18477 393 18523 399
rect 18773 393 18819 399
rect 17723 253 17769 259
rect 18389 253 18435 259
rect 19055 253 19101 259
rect 17717 219 17729 253
rect 17763 219 18395 253
rect 18429 219 19061 253
rect 19095 219 19107 253
rect 17723 213 17769 219
rect 18389 213 18435 219
rect 19055 213 19101 219
rect -34 17 19348 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6569 17
rect 6603 -17 6643 17
rect 6677 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7753 17
rect 7787 -17 7827 17
rect 7861 -17 7901 17
rect 7935 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8123 17
rect 8157 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8567 17
rect 8601 -17 8715 17
rect 8749 -17 8789 17
rect 8823 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9529 17
rect 9563 -17 9677 17
rect 9711 -17 9751 17
rect 9785 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10195 17
rect 10229 -17 10269 17
rect 10303 -17 10343 17
rect 10377 -17 10417 17
rect 10451 -17 10491 17
rect 10525 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10861 17
rect 10895 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11305 17
rect 11339 -17 11379 17
rect 11413 -17 11453 17
rect 11487 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12193 17
rect 12227 -17 12267 17
rect 12301 -17 12341 17
rect 12375 -17 12415 17
rect 12449 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12859 17
rect 12893 -17 12933 17
rect 12967 -17 13007 17
rect 13041 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13525 17
rect 13559 -17 13599 17
rect 13633 -17 13673 17
rect 13707 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13895 17
rect 13929 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14191 17
rect 14225 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14635 17
rect 14669 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14857 17
rect 14891 -17 14931 17
rect 14965 -17 15005 17
rect 15039 -17 15079 17
rect 15113 -17 15153 17
rect 15187 -17 15227 17
rect 15261 -17 15301 17
rect 15335 -17 15449 17
rect 15483 -17 15523 17
rect 15557 -17 15597 17
rect 15631 -17 15671 17
rect 15705 -17 15745 17
rect 15779 -17 15819 17
rect 15853 -17 15893 17
rect 15927 -17 15967 17
rect 16001 -17 16041 17
rect 16075 -17 16115 17
rect 16149 -17 16189 17
rect 16223 -17 16263 17
rect 16297 -17 16411 17
rect 16445 -17 16485 17
rect 16519 -17 16559 17
rect 16593 -17 16633 17
rect 16667 -17 16707 17
rect 16741 -17 16781 17
rect 16815 -17 16855 17
rect 16889 -17 16929 17
rect 16963 -17 17003 17
rect 17037 -17 17077 17
rect 17111 -17 17151 17
rect 17185 -17 17225 17
rect 17259 -17 17373 17
rect 17407 -17 17447 17
rect 17481 -17 17521 17
rect 17555 -17 17595 17
rect 17629 -17 17669 17
rect 17703 -17 17743 17
rect 17777 -17 17817 17
rect 17851 -17 17891 17
rect 17925 -17 18039 17
rect 18073 -17 18113 17
rect 18147 -17 18187 17
rect 18221 -17 18261 17
rect 18295 -17 18335 17
rect 18369 -17 18409 17
rect 18443 -17 18483 17
rect 18517 -17 18557 17
rect 18591 -17 18705 17
rect 18739 -17 18779 17
rect 18813 -17 18853 17
rect 18887 -17 18927 17
rect 18961 -17 19001 17
rect 19035 -17 19075 17
rect 19109 -17 19149 17
rect 19183 -17 19223 17
rect 19257 -17 19348 17
rect -34 -34 19348 -17
<< labels >>
rlabel metal1 2351 575 2385 609 1 SN
port 1 n
rlabel metal1 427 427 461 461 1 RN
port 2 n
rlabel metal1 427 501 461 535 1 RN
port 3 n
rlabel metal1 427 575 461 609 1 RN
port 4 n
rlabel metal1 427 649 461 683 1 RN
port 5 n
rlabel metal1 427 723 461 757 1 RN
port 6 n
rlabel metal1 427 871 461 905 1 RN
port 7 n
rlabel metal1 205 797 239 831 1 D
port 8 n
rlabel metal1 205 723 239 757 1 D
port 9 n
rlabel metal1 205 649 239 683 1 D
port 10 n
rlabel metal1 205 575 239 609 1 D
port 11 n
rlabel metal1 205 501 239 535 1 D
port 12 n
rlabel metal1 205 427 239 461 1 D
port 13 n
rlabel metal1 205 871 239 905 1 D
port 14 n
rlabel metal1 2351 501 2385 535 1 SN
port 15 n
rlabel metal1 5977 797 6011 831 1 D
port 16 n
rlabel metal1 11749 797 11783 831 1 D
port 17 n
rlabel metal1 11749 501 11783 535 1 D
port 18 n
rlabel metal1 5977 723 6011 757 1 D
port 19 n
rlabel metal1 5977 501 6011 535 1 D
port 20 n
rlabel metal1 3535 427 3569 461 1 RN
port 21 n
rlabel metal1 4275 427 4309 461 1 RN
port 22 n
rlabel metal1 3535 501 3569 535 1 RN
port 23 n
rlabel metal1 4275 501 4309 535 1 RN
port 24 n
rlabel metal1 4275 649 4309 683 1 RN
port 25 n
rlabel metal1 6199 427 6233 461 1 RN
port 26 n
rlabel metal1 6199 501 6233 535 1 RN
port 27 n
rlabel metal1 6199 723 6233 757 1 RN
port 28 n
rlabel metal1 9307 427 9341 461 1 RN
port 29 n
rlabel metal1 9307 501 9341 535 1 RN
port 30 n
rlabel metal1 10047 427 10081 461 1 RN
port 31 n
rlabel metal1 10047 501 10081 535 1 RN
port 32 n
rlabel metal1 11971 427 12005 461 1 RN
port 33 n
rlabel metal1 11971 501 12005 535 1 RN
port 34 n
rlabel metal1 11971 797 12005 831 1 RN
port 35 n
rlabel metal1 15079 427 15113 461 1 RN
port 36 n
rlabel metal1 15819 427 15853 461 1 RN
port 37 n
rlabel metal1 15819 501 15853 535 1 RN
port 38 n
rlabel metal1 15079 501 15113 535 1 RN
port 39 n
rlabel metal1 9085 871 9119 905 1 CLK
port 40 n
rlabel metal1 7161 871 7195 905 1 CLK
port 41 n
rlabel metal1 3313 871 3347 905 1 CLK
port 42 n
rlabel metal1 1389 871 1423 905 1 CLK
port 43 n
rlabel metal1 1389 723 1423 757 1 CLK
port 44 n
rlabel metal1 1389 575 1423 609 1 CLK
port 45 n
rlabel metal1 3313 501 3347 535 1 CLK
port 46 n
rlabel metal1 7161 723 7195 757 1 CLK
port 47 n
rlabel metal1 12933 871 12967 905 1 CLK
port 48 n
rlabel metal1 14857 871 14891 905 1 CLK
port 49 n
rlabel metal1 14857 501 14891 535 1 CLK
port 50 n
rlabel metal1 5237 575 5271 609 1 SN
port 51 n
rlabel metal1 5237 501 5271 535 1 SN
port 52 n
rlabel metal1 8123 575 8157 609 1 SN
port 53 n
rlabel metal1 5977 649 6011 683 1 D
port 54 n
rlabel metal1 6199 649 6233 683 1 RN
port 55 n
rlabel metal1 8123 501 8157 535 1 SN
port 56 n
rlabel metal1 11009 575 11043 609 1 SN
port 57 n
rlabel metal1 10047 649 10081 683 1 RN
port 58 n
rlabel metal1 13895 575 13929 609 1 SN
port 59 n
rlabel metal1 11971 649 12005 683 1 RN
port 60 n
rlabel metal1 11749 649 11783 683 1 D
port 61 n
rlabel metal1 15819 649 15853 683 1 RN
port 62 n
rlabel metal1 13895 501 13929 535 1 SN
port 63 n
rlabel metal1 9085 501 9119 535 1 CLK
port 64 n
rlabel metal1 19149 797 19183 831 1 Q
port 65 n
rlabel metal1 -34 1446 19348 1514 1 VPWR
port 66 n
rlabel metal1 -34 -34 19348 34 1 VGND
port 67 n
rlabel nwell 57 1463 91 1497 1 VPB
port 68 n
rlabel pwell 57 -17 91 17 1 VNB
port 69 n
<< end >>
