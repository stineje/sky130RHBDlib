magic
tech sky130A
magscale 1 2
timestamp 1652507010
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 427 871 461 905
rect 2647 871 2681 905
rect 4719 871 4753 905
rect 6939 871 6973 905
rect 9011 871 9045 905
rect 11231 871 11265 905
rect 15153 797 15187 831
rect 427 723 461 757
rect 4719 723 4753 757
rect 9011 723 9045 757
rect 15153 723 15187 757
rect 427 649 461 683
rect 2647 649 2681 683
rect 4719 649 4753 683
rect 6939 649 6973 683
rect 9011 649 9045 683
rect 11231 649 11265 683
rect 15153 649 15187 683
rect 427 575 461 609
rect 1315 575 1349 609
rect 2647 575 2681 609
rect 15153 575 15187 609
rect 427 501 461 535
rect 1315 501 1349 535
rect 5607 501 5641 535
rect 9899 501 9933 535
rect 15153 501 15187 535
rect 15153 427 15187 461
<< metal1 >>
rect -34 1446 15352 1514
rect 3349 904 4707 905
rect 479 873 2611 904
rect 2693 873 4707 904
rect 3349 871 4707 873
rect 4789 871 6903 905
rect 6985 871 8999 905
rect 9081 871 11195 905
rect 12079 871 12450 905
rect 3495 723 3827 757
rect 7741 723 8114 757
rect 11931 723 13041 757
rect 3348 575 14068 609
rect 1385 501 5595 535
rect 5677 501 9863 535
rect 7639 427 13263 461
rect -34 -34 15352 34
use li1_M1_contact  li1_M1_contact_14 pcells
timestamp 1648061256
transform -1 0 1332 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 4144 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 3330 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform -1 0 3478 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform 1 0 3848 0 1 740
box -53 -33 29 33
use dffx1_pcell  dffx1_pcell_0 pcells
timestamp 1652395794
transform 1 0 0 0 1 0
box -87 -34 4379 1550
use dffx1_pcell  dffx1_pcell_1
timestamp 1652395794
transform 1 0 4292 0 1 0
box -87 -34 4379 1550
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform -1 0 5624 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 8140 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform 1 0 8436 0 1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 7622 0 -1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 7770 0 -1 740
box -53 -33 29 33
use dffx1_pcell  dffx1_pcell_2
timestamp 1652395794
transform 1 0 8584 0 1 0
box -87 -34 4379 1550
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform 1 0 9916 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 13246 0 -1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 13024 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 12728 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 12432 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 11914 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 12062 0 -1 888
box -53 -33 29 33
use voter3x1_pcell  voter3x1_pcell_0 pcells
timestamp 1652393968
transform 1 0 12876 0 1 0
box -87 -34 2529 1550
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 14060 0 -1 592
box -53 -33 29 33
<< labels >>
rlabel locali 15153 797 15187 831 1 Q
port 1 nsew signal output
rlabel locali 15153 723 15187 757 1 Q
port 1 nsew signal output
rlabel locali 15153 649 15187 683 1 Q
port 1 nsew signal output
rlabel locali 15153 575 15187 609 1 Q
port 1 nsew signal output
rlabel locali 15153 501 15187 535 1 Q
port 1 nsew signal output
rlabel locali 15153 427 15187 461 1 Q
port 1 nsew signal output
rlabel locali 1315 501 1349 535 1 D
port 2 nsew signal input
rlabel locali 1315 575 1349 609 1 D
port 2 nsew signal input
rlabel locali 5607 501 5641 535 1 D
port 2 nsew signal input
rlabel locali 9899 501 9933 535 1 D
port 2 nsew signal input
rlabel locali 427 871 461 905 1 CLK
port 3 nsew signal input
rlabel locali 427 723 461 757 1 CLK
port 3 nsew signal input
rlabel locali 427 649 461 683 1 CLK
port 3 nsew signal input
rlabel locali 427 575 461 609 1 CLK
port 3 nsew signal input
rlabel locali 427 501 461 535 1 CLK
port 3 nsew signal input
rlabel locali 2647 649 2681 683 1 CLK
port 3 nsew signal input
rlabel locali 2647 575 2681 609 1 CLK
port 3 nsew signal input
rlabel locali 2647 871 2681 905 1 CLK
port 3 nsew signal input
rlabel locali 4719 649 4753 683 1 CLK
port 3 nsew signal input
rlabel locali 4719 723 4753 757 1 CLK
port 3 nsew signal input
rlabel locali 4719 871 4753 905 1 CLK
port 3 nsew signal input
rlabel locali 6939 649 6973 683 1 CLK
port 3 nsew signal input
rlabel locali 6939 871 6973 905 1 CLK
port 3 nsew signal input
rlabel locali 9011 649 9045 683 1 CLK
port 3 nsew signal input
rlabel locali 9011 723 9045 757 1 CLK
port 3 nsew signal input
rlabel locali 9011 871 9045 905 1 CLK
port 3 nsew signal input
rlabel locali 11231 649 11265 683 1 CLK
port 3 nsew signal input
rlabel locali 11231 871 11265 905 1 CLK
port 3 nsew signal input
rlabel metal1 -34 1446 15352 1514 1 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 -34 -34 15352 34 1 VGND
port 5 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
port 6 nsew power bidirectional
rlabel pwell 57 -17 91 17 1 VPB
port 7 nsew ground bidirectional
<< properties >>
string LEFclass CORE
string LEFsite unithd
string FIXED_BBOX 0 0 15318 1480
string LEFsymmetry X Y R90
<< end >>
