magic
tech sky130A
magscale 1 2
timestamp 1669200965
<< nwell >>
rect -87 786 1493 1550
<< pwell >>
rect -34 -34 1440 544
<< nmos >>
rect 147 290 177 351
tri 177 290 193 306 sw
rect 447 290 477 351
rect 147 260 253 290
tri 253 260 283 290 sw
rect 147 159 177 260
tri 177 244 193 260 nw
tri 237 244 253 260 ne
tri 177 159 193 175 sw
tri 237 159 253 175 se
rect 253 159 283 260
tri 342 260 372 290 se
rect 372 260 477 290
rect 342 166 372 260
tri 372 244 388 260 nw
tri 431 244 447 260 ne
tri 372 166 388 182 sw
tri 431 166 447 182 se
rect 447 166 477 260
tri 147 129 177 159 ne
rect 177 129 253 159
tri 253 129 283 159 nw
tri 342 136 372 166 ne
rect 372 136 447 166
tri 447 136 477 166 nw
rect 649 298 679 351
tri 679 298 695 314 sw
rect 649 268 755 298
tri 755 268 785 298 sw
rect 649 167 679 268
tri 679 252 695 268 nw
tri 739 252 755 268 ne
tri 679 167 695 183 sw
tri 739 167 755 183 se
rect 755 167 785 268
tri 649 137 679 167 ne
rect 679 137 755 167
tri 755 137 785 167 nw
rect 1117 297 1147 350
tri 1147 297 1163 313 sw
rect 1117 267 1223 297
tri 1223 267 1253 297 sw
rect 1117 166 1147 267
tri 1147 251 1163 267 nw
tri 1207 251 1223 267 ne
tri 1147 166 1163 182 sw
tri 1207 166 1223 182 se
rect 1223 166 1253 267
tri 1117 136 1147 166 ne
rect 1147 136 1223 166
tri 1223 136 1253 166 nw
<< pmos >>
rect 247 1004 277 1404
rect 335 1004 365 1404
rect 423 1004 453 1404
rect 511 1004 541 1404
rect 599 1004 629 1404
rect 687 1004 717 1404
rect 1126 1004 1156 1404
rect 1214 1004 1244 1404
<< ndiff >>
rect 91 335 147 351
rect 91 301 101 335
rect 135 301 147 335
rect 91 263 147 301
rect 177 335 447 351
rect 177 306 198 335
tri 177 290 193 306 ne
rect 193 301 198 306
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 447 335
rect 193 290 447 301
rect 477 335 533 351
rect 477 301 489 335
rect 523 301 533 335
rect 91 229 101 263
rect 135 229 147 263
tri 253 260 283 290 ne
rect 283 263 342 290
rect 91 195 147 229
rect 91 161 101 195
rect 135 161 147 195
rect 91 129 147 161
tri 177 244 193 260 se
rect 193 244 237 260
tri 237 244 253 260 sw
rect 177 210 253 244
rect 177 176 198 210
rect 232 176 253 210
rect 177 175 253 176
tri 177 159 193 175 ne
rect 193 159 237 175
tri 237 159 253 175 nw
rect 283 229 295 263
rect 329 229 342 263
tri 342 260 372 290 nw
rect 283 195 342 229
rect 283 161 295 195
rect 329 161 342 195
tri 372 244 388 260 se
rect 388 244 431 260
tri 431 244 447 260 sw
rect 372 216 447 244
rect 372 182 393 216
rect 427 182 447 216
tri 372 166 388 182 ne
rect 388 166 431 182
tri 431 166 447 182 nw
tri 147 129 177 159 sw
tri 253 129 283 159 se
rect 283 136 342 161
tri 342 136 372 166 sw
tri 447 136 477 166 se
rect 477 136 533 301
rect 283 129 533 136
rect 91 125 533 129
rect 91 91 101 125
rect 135 91 295 125
rect 329 91 392 125
rect 426 91 489 125
rect 523 91 533 125
rect 91 75 533 91
rect 593 335 649 351
rect 593 301 603 335
rect 637 301 649 335
rect 593 263 649 301
rect 679 314 841 351
tri 679 298 695 314 ne
rect 695 298 841 314
tri 755 268 785 298 ne
rect 593 229 603 263
rect 637 229 649 263
rect 593 195 649 229
rect 593 161 603 195
rect 637 161 649 195
tri 679 252 695 268 se
rect 695 252 739 268
tri 739 252 755 268 sw
rect 679 219 755 252
rect 679 185 700 219
rect 734 185 755 219
rect 679 183 755 185
tri 679 167 695 183 ne
rect 695 167 739 183
tri 739 167 755 183 nw
rect 785 263 841 298
rect 785 229 797 263
rect 831 229 841 263
rect 785 195 841 229
rect 593 137 649 161
tri 649 137 679 167 sw
tri 755 137 785 167 se
rect 785 161 797 195
rect 831 161 841 195
rect 785 137 841 161
rect 593 125 841 137
rect 593 91 603 125
rect 637 91 700 125
rect 734 91 797 125
rect 831 91 841 125
rect 593 75 841 91
rect 1061 334 1117 350
rect 1061 300 1071 334
rect 1105 300 1117 334
rect 1061 262 1117 300
rect 1147 334 1307 350
rect 1147 313 1265 334
tri 1147 297 1163 313 ne
rect 1163 300 1265 313
rect 1299 300 1307 334
rect 1163 297 1307 300
tri 1223 267 1253 297 ne
rect 1061 228 1071 262
rect 1105 228 1117 262
rect 1061 194 1117 228
rect 1061 160 1071 194
rect 1105 160 1117 194
tri 1147 251 1163 267 se
rect 1163 251 1207 267
tri 1207 251 1223 267 sw
rect 1147 218 1223 251
rect 1147 184 1167 218
rect 1201 184 1223 218
rect 1147 182 1223 184
tri 1147 166 1163 182 ne
rect 1163 166 1207 182
tri 1207 166 1223 182 nw
rect 1253 262 1307 297
rect 1253 228 1265 262
rect 1299 228 1307 262
rect 1253 194 1307 228
rect 1061 136 1117 160
tri 1117 136 1147 166 sw
tri 1223 136 1253 166 se
rect 1253 160 1265 194
rect 1299 160 1307 194
rect 1253 136 1307 160
rect 1061 124 1307 136
rect 1061 90 1071 124
rect 1105 90 1167 124
rect 1201 90 1265 124
rect 1299 90 1307 124
rect 1061 74 1307 90
<< pdiff >>
rect 191 1366 247 1404
rect 191 1332 201 1366
rect 235 1332 247 1366
rect 191 1298 247 1332
rect 191 1264 201 1298
rect 235 1264 247 1298
rect 191 1230 247 1264
rect 191 1196 201 1230
rect 235 1196 247 1230
rect 191 1162 247 1196
rect 191 1128 201 1162
rect 235 1128 247 1162
rect 191 1093 247 1128
rect 191 1059 201 1093
rect 235 1059 247 1093
rect 191 1004 247 1059
rect 277 1366 335 1404
rect 277 1332 289 1366
rect 323 1332 335 1366
rect 277 1298 335 1332
rect 277 1264 289 1298
rect 323 1264 335 1298
rect 277 1230 335 1264
rect 277 1196 289 1230
rect 323 1196 335 1230
rect 277 1162 335 1196
rect 277 1128 289 1162
rect 323 1128 335 1162
rect 277 1093 335 1128
rect 277 1059 289 1093
rect 323 1059 335 1093
rect 277 1004 335 1059
rect 365 1366 423 1404
rect 365 1332 377 1366
rect 411 1332 423 1366
rect 365 1298 423 1332
rect 365 1264 377 1298
rect 411 1264 423 1298
rect 365 1230 423 1264
rect 365 1196 377 1230
rect 411 1196 423 1230
rect 365 1162 423 1196
rect 365 1128 377 1162
rect 411 1128 423 1162
rect 365 1004 423 1128
rect 453 1366 511 1404
rect 453 1332 465 1366
rect 499 1332 511 1366
rect 453 1298 511 1332
rect 453 1264 465 1298
rect 499 1264 511 1298
rect 453 1230 511 1264
rect 453 1196 465 1230
rect 499 1196 511 1230
rect 453 1162 511 1196
rect 453 1128 465 1162
rect 499 1128 511 1162
rect 453 1093 511 1128
rect 453 1059 465 1093
rect 499 1059 511 1093
rect 453 1004 511 1059
rect 541 1366 599 1404
rect 541 1332 553 1366
rect 587 1332 599 1366
rect 541 1298 599 1332
rect 541 1264 553 1298
rect 587 1264 599 1298
rect 541 1230 599 1264
rect 541 1196 553 1230
rect 587 1196 599 1230
rect 541 1162 599 1196
rect 541 1128 553 1162
rect 587 1128 599 1162
rect 541 1004 599 1128
rect 629 1366 687 1404
rect 629 1332 641 1366
rect 675 1332 687 1366
rect 629 1298 687 1332
rect 629 1264 641 1298
rect 675 1264 687 1298
rect 629 1230 687 1264
rect 629 1196 641 1230
rect 675 1196 687 1230
rect 629 1162 687 1196
rect 629 1128 641 1162
rect 675 1128 687 1162
rect 629 1093 687 1128
rect 629 1059 641 1093
rect 675 1059 687 1093
rect 629 1004 687 1059
rect 717 1366 771 1404
rect 717 1332 729 1366
rect 763 1332 771 1366
rect 717 1298 771 1332
rect 717 1264 729 1298
rect 763 1264 771 1298
rect 717 1230 771 1264
rect 717 1196 729 1230
rect 763 1196 771 1230
rect 717 1162 771 1196
rect 717 1128 729 1162
rect 763 1128 771 1162
rect 717 1004 771 1128
rect 1070 1366 1126 1404
rect 1070 1332 1080 1366
rect 1114 1332 1126 1366
rect 1070 1298 1126 1332
rect 1070 1264 1080 1298
rect 1114 1264 1126 1298
rect 1070 1230 1126 1264
rect 1070 1196 1080 1230
rect 1114 1196 1126 1230
rect 1070 1162 1126 1196
rect 1070 1128 1080 1162
rect 1114 1128 1126 1162
rect 1070 1093 1126 1128
rect 1070 1059 1080 1093
rect 1114 1059 1126 1093
rect 1070 1004 1126 1059
rect 1156 1366 1214 1404
rect 1156 1332 1168 1366
rect 1202 1332 1214 1366
rect 1156 1298 1214 1332
rect 1156 1264 1168 1298
rect 1202 1264 1214 1298
rect 1156 1230 1214 1264
rect 1156 1196 1168 1230
rect 1202 1196 1214 1230
rect 1156 1162 1214 1196
rect 1156 1128 1168 1162
rect 1202 1128 1214 1162
rect 1156 1093 1214 1128
rect 1156 1059 1168 1093
rect 1202 1059 1214 1093
rect 1156 1004 1214 1059
rect 1244 1366 1298 1404
rect 1244 1332 1256 1366
rect 1290 1332 1298 1366
rect 1244 1298 1298 1332
rect 1244 1264 1256 1298
rect 1290 1264 1298 1298
rect 1244 1230 1298 1264
rect 1244 1196 1256 1230
rect 1290 1196 1298 1230
rect 1244 1162 1298 1196
rect 1244 1128 1256 1162
rect 1290 1128 1298 1162
rect 1244 1093 1298 1128
rect 1244 1059 1256 1093
rect 1290 1059 1298 1093
rect 1244 1004 1298 1059
<< ndiffc >>
rect 101 301 135 335
rect 198 301 232 335
rect 295 301 329 335
rect 392 301 426 335
rect 489 301 523 335
rect 101 229 135 263
rect 101 161 135 195
rect 198 176 232 210
rect 295 229 329 263
rect 295 161 329 195
rect 393 182 427 216
rect 101 91 135 125
rect 295 91 329 125
rect 392 91 426 125
rect 489 91 523 125
rect 603 301 637 335
rect 603 229 637 263
rect 603 161 637 195
rect 700 185 734 219
rect 797 229 831 263
rect 797 161 831 195
rect 603 91 637 125
rect 700 91 734 125
rect 797 91 831 125
rect 1071 300 1105 334
rect 1265 300 1299 334
rect 1071 228 1105 262
rect 1071 160 1105 194
rect 1167 184 1201 218
rect 1265 228 1299 262
rect 1265 160 1299 194
rect 1071 90 1105 124
rect 1167 90 1201 124
rect 1265 90 1299 124
<< pdiffc >>
rect 201 1332 235 1366
rect 201 1264 235 1298
rect 201 1196 235 1230
rect 201 1128 235 1162
rect 201 1059 235 1093
rect 289 1332 323 1366
rect 289 1264 323 1298
rect 289 1196 323 1230
rect 289 1128 323 1162
rect 289 1059 323 1093
rect 377 1332 411 1366
rect 377 1264 411 1298
rect 377 1196 411 1230
rect 377 1128 411 1162
rect 465 1332 499 1366
rect 465 1264 499 1298
rect 465 1196 499 1230
rect 465 1128 499 1162
rect 465 1059 499 1093
rect 553 1332 587 1366
rect 553 1264 587 1298
rect 553 1196 587 1230
rect 553 1128 587 1162
rect 641 1332 675 1366
rect 641 1264 675 1298
rect 641 1196 675 1230
rect 641 1128 675 1162
rect 641 1059 675 1093
rect 729 1332 763 1366
rect 729 1264 763 1298
rect 729 1196 763 1230
rect 729 1128 763 1162
rect 1080 1332 1114 1366
rect 1080 1264 1114 1298
rect 1080 1196 1114 1230
rect 1080 1128 1114 1162
rect 1080 1059 1114 1093
rect 1168 1332 1202 1366
rect 1168 1264 1202 1298
rect 1168 1196 1202 1230
rect 1168 1128 1202 1162
rect 1168 1059 1202 1093
rect 1256 1332 1290 1366
rect 1256 1264 1290 1298
rect 1256 1196 1290 1230
rect 1256 1128 1290 1162
rect 1256 1059 1290 1093
<< psubdiff >>
rect -34 482 1440 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 928 461 996 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 928 427 945 461
rect 979 427 996 461
rect 1372 461 1440 482
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect 1372 427 1389 461
rect 1423 427 1440 461
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 928 313 996 353
rect 1372 387 1440 427
rect 1372 353 1389 387
rect 1423 353 1440 387
rect 928 279 945 313
rect 979 279 996 313
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect -34 17 34 57
rect 928 57 945 91
rect 979 57 996 91
rect 1372 313 1440 353
rect 1372 279 1389 313
rect 1423 279 1440 313
rect 1372 239 1440 279
rect 1372 205 1389 239
rect 1423 205 1440 239
rect 1372 165 1440 205
rect 1372 131 1389 165
rect 1423 131 1440 165
rect 1372 91 1440 131
rect 928 17 996 57
rect 1372 57 1389 91
rect 1423 57 1440 91
rect 1372 17 1440 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1440 17
rect -34 -34 1440 -17
<< nsubdiff >>
rect -34 1497 1440 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1440 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 928 1423 996 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 1372 1423 1440 1463
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect 928 1019 945 1053
rect 979 1019 996 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 928 979 996 1019
rect 1372 1389 1389 1423
rect 1423 1389 1440 1423
rect 1372 1349 1440 1389
rect 1372 1315 1389 1349
rect 1423 1315 1440 1349
rect 1372 1275 1440 1315
rect 1372 1241 1389 1275
rect 1423 1241 1440 1275
rect 1372 1201 1440 1241
rect 1372 1167 1389 1201
rect 1423 1167 1440 1201
rect 1372 1127 1440 1167
rect 1372 1093 1389 1127
rect 1423 1093 1440 1127
rect 1372 1053 1440 1093
rect 1372 1019 1389 1053
rect 1423 1019 1440 1053
rect 928 945 945 979
rect 979 945 996 979
rect -34 871 -17 905
rect 17 884 34 905
rect 928 905 996 945
rect 1372 979 1440 1019
rect 1372 945 1389 979
rect 1423 945 1440 979
rect 928 884 945 905
rect 17 871 945 884
rect 979 884 996 905
rect 1372 905 1440 945
rect 1372 884 1389 905
rect 979 871 1389 884
rect 1423 871 1440 905
rect -34 822 1440 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 945 427 979 461
rect 945 353 979 387
rect 1389 427 1423 461
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1389 353 1423 387
rect 945 279 979 313
rect 945 205 979 239
rect 945 131 979 165
rect 945 57 979 91
rect 1389 279 1423 313
rect 1389 205 1423 239
rect 1389 131 1423 165
rect 1389 57 1423 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 945 1389 979 1423
rect 945 1315 979 1349
rect 945 1241 979 1275
rect 945 1167 979 1201
rect 945 1093 979 1127
rect 945 1019 979 1053
rect -17 945 17 979
rect 1389 1389 1423 1423
rect 1389 1315 1423 1349
rect 1389 1241 1423 1275
rect 1389 1167 1423 1201
rect 1389 1093 1423 1127
rect 1389 1019 1423 1053
rect 945 945 979 979
rect -17 871 17 905
rect 1389 945 1423 979
rect 945 871 979 905
rect 1389 871 1423 905
<< poly >>
rect 247 1404 277 1430
rect 335 1404 365 1430
rect 423 1404 453 1430
rect 511 1404 541 1430
rect 599 1404 629 1430
rect 687 1404 717 1430
rect 1126 1404 1156 1430
rect 1214 1404 1244 1430
rect 247 973 277 1004
rect 335 973 365 1004
rect 423 973 453 1004
rect 511 973 541 1004
rect 195 957 365 973
rect 195 923 205 957
rect 239 943 365 957
rect 417 957 541 973
rect 239 923 249 943
rect 195 907 249 923
rect 417 923 427 957
rect 461 943 541 957
rect 599 973 629 1004
rect 687 973 717 1004
rect 599 957 717 973
rect 599 943 649 957
rect 461 923 471 943
rect 417 907 471 923
rect 639 923 649 943
rect 683 943 717 957
rect 1126 973 1156 1004
rect 1214 973 1244 1004
rect 683 923 693 943
rect 639 907 693 923
rect 1083 957 1244 973
rect 1083 923 1093 957
rect 1127 943 1244 957
rect 1127 923 1137 943
rect 1083 907 1137 923
rect 195 433 249 449
rect 195 413 205 433
rect 147 399 205 413
rect 239 399 249 433
rect 147 383 249 399
rect 417 433 471 449
rect 417 399 427 433
rect 461 413 471 433
rect 639 433 693 449
rect 461 399 477 413
rect 417 383 477 399
rect 639 399 649 433
rect 683 399 693 433
rect 639 383 693 399
rect 147 351 177 383
rect 447 351 477 383
rect 649 351 679 383
rect 1083 434 1137 450
rect 1083 400 1093 434
rect 1127 413 1137 434
rect 1127 400 1147 413
rect 1083 384 1147 400
rect 1117 350 1147 384
<< polycont >>
rect 205 923 239 957
rect 427 923 461 957
rect 649 923 683 957
rect 1093 923 1127 957
rect 205 399 239 433
rect 427 399 461 433
rect 649 399 683 433
rect 1093 400 1127 434
<< locali >>
rect -34 1497 1440 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1440 1497
rect -34 1446 1440 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 201 1366 235 1446
rect 201 1298 235 1332
rect 201 1230 235 1264
rect 201 1162 235 1196
rect 201 1093 235 1128
rect 201 1043 235 1059
rect 289 1366 323 1404
rect 289 1298 323 1332
rect 289 1230 323 1264
rect 289 1162 323 1196
rect 289 1093 323 1128
rect 377 1366 411 1446
rect 377 1298 411 1332
rect 377 1230 411 1264
rect 377 1162 411 1196
rect 377 1111 411 1128
rect 465 1366 499 1404
rect 465 1298 499 1332
rect 465 1230 499 1264
rect 465 1162 499 1196
rect 289 1048 323 1059
rect 465 1093 499 1128
rect 553 1366 587 1446
rect 553 1298 587 1332
rect 553 1230 587 1264
rect 553 1162 587 1196
rect 553 1111 587 1128
rect 641 1366 675 1404
rect 641 1298 675 1332
rect 641 1230 675 1264
rect 641 1162 675 1196
rect 465 1048 499 1059
rect 641 1093 675 1128
rect 729 1366 763 1446
rect 729 1298 763 1332
rect 729 1230 763 1264
rect 729 1162 763 1196
rect 729 1111 763 1128
rect 928 1423 996 1446
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 641 1048 675 1059
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect -34 979 34 1019
rect 289 1014 831 1048
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 923
rect 205 383 239 399
rect 427 957 461 973
rect 427 433 461 923
rect 427 383 461 399
rect 649 957 683 973
rect 649 433 683 923
rect 649 383 683 399
rect 797 683 831 1014
rect 928 1019 945 1053
rect 979 1019 996 1053
rect 1080 1366 1114 1446
rect 1080 1298 1114 1332
rect 1080 1230 1114 1264
rect 1080 1162 1114 1196
rect 1080 1093 1114 1128
rect 1080 1037 1114 1059
rect 1168 1366 1202 1404
rect 1168 1298 1202 1332
rect 1168 1230 1202 1264
rect 1168 1162 1202 1196
rect 1168 1093 1202 1128
rect 928 979 996 1019
rect 928 945 945 979
rect 979 945 996 979
rect 928 905 996 945
rect 928 871 945 905
rect 979 871 996 905
rect 928 822 996 871
rect 1093 957 1127 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 101 335 135 351
rect 295 335 329 351
rect 489 335 523 351
rect 135 301 198 335
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 489 335
rect 101 263 135 301
rect 101 195 135 229
rect 295 263 329 301
rect 489 285 523 301
rect 603 335 637 351
rect 797 350 831 649
rect 1093 683 1127 923
rect 1168 933 1202 1059
rect 1256 1366 1290 1446
rect 1256 1298 1290 1332
rect 1256 1230 1290 1264
rect 1256 1162 1290 1196
rect 1256 1093 1290 1128
rect 1256 1037 1290 1059
rect 1372 1423 1440 1446
rect 1372 1389 1389 1423
rect 1423 1389 1440 1423
rect 1372 1349 1440 1389
rect 1372 1315 1389 1349
rect 1423 1315 1440 1349
rect 1372 1275 1440 1315
rect 1372 1241 1389 1275
rect 1423 1241 1440 1275
rect 1372 1201 1440 1241
rect 1372 1167 1389 1201
rect 1423 1167 1440 1201
rect 1372 1127 1440 1167
rect 1372 1093 1389 1127
rect 1423 1093 1440 1127
rect 1372 1053 1440 1093
rect 1372 1019 1389 1053
rect 1423 1019 1440 1053
rect 1372 979 1440 1019
rect 1372 945 1389 979
rect 1423 945 1440 979
rect 1168 899 1275 933
rect 603 263 637 301
rect 101 125 135 161
rect 101 75 135 91
rect 198 210 232 226
rect -34 34 34 57
rect 198 34 232 176
rect 295 195 329 229
rect 393 216 427 232
rect 603 216 637 229
rect 427 195 637 216
rect 427 182 603 195
rect 393 166 427 182
rect 295 125 329 161
rect 700 316 831 350
rect 928 461 996 544
rect 928 427 945 461
rect 979 427 996 461
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect 1093 434 1127 649
rect 1241 433 1275 899
rect 1372 905 1440 945
rect 1372 871 1389 905
rect 1423 871 1440 905
rect 1372 822 1440 871
rect 1093 384 1127 400
rect 1167 399 1275 433
rect 1372 461 1440 544
rect 1372 427 1389 461
rect 1423 427 1440 461
rect 700 219 734 316
rect 928 313 996 353
rect 928 279 945 313
rect 979 279 996 313
rect 700 169 734 185
rect 797 263 831 279
rect 797 195 831 229
rect 489 125 523 141
rect 329 91 392 125
rect 426 91 489 125
rect 295 75 329 91
rect 489 75 523 91
rect 603 125 637 161
rect 797 125 831 161
rect 637 91 700 125
rect 734 91 797 125
rect 603 75 637 91
rect 797 75 831 91
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect 928 57 945 91
rect 979 57 996 91
rect 928 34 996 57
rect 1071 334 1105 350
rect 1071 262 1105 300
rect 1071 194 1105 228
rect 1167 218 1201 399
rect 1372 387 1440 427
rect 1372 353 1389 387
rect 1423 353 1440 387
rect 1167 168 1201 184
rect 1265 334 1299 350
rect 1265 262 1299 300
rect 1265 194 1299 228
rect 1071 124 1105 160
rect 1265 124 1299 160
rect 1105 90 1167 124
rect 1201 90 1265 124
rect 1071 34 1105 90
rect 1168 34 1202 90
rect 1265 34 1299 90
rect 1372 313 1440 353
rect 1372 279 1389 313
rect 1423 279 1440 313
rect 1372 239 1440 279
rect 1372 205 1389 239
rect 1423 205 1440 239
rect 1372 165 1440 205
rect 1372 131 1389 165
rect 1423 131 1440 165
rect 1372 91 1440 131
rect 1372 57 1389 91
rect 1423 57 1440 91
rect 1372 34 1440 57
rect -34 17 1440 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1440 17
rect -34 -34 1440 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 797 649 831 683
rect 1093 649 1127 683
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
<< metal1 >>
rect -34 1497 1440 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1440 1497
rect -34 1446 1440 1463
rect 791 683 837 689
rect 1087 683 1133 689
rect 785 649 797 683
rect 831 649 1093 683
rect 1127 649 1139 683
rect 791 643 837 649
rect 1087 643 1133 649
rect -34 17 1440 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1440 17
rect -34 -34 1440 -17
<< labels >>
rlabel metal1 1241 427 1275 461 1 Y
port 1 n
rlabel metal1 1241 501 1275 535 1 Y
port 2 n
rlabel metal1 1241 575 1275 609 1 Y
port 3 n
rlabel metal1 1241 649 1275 683 1 Y
port 4 n
rlabel metal1 1241 723 1275 757 1 Y
port 5 n
rlabel metal1 1241 797 1275 831 1 Y
port 6 n
rlabel metal1 1241 871 1275 905 1 Y
port 7 n
rlabel metal1 205 871 239 905 1 A
port 8 n
rlabel metal1 205 797 239 831 1 A
port 9 n
rlabel metal1 205 723 239 757 1 A
port 10 n
rlabel metal1 205 649 239 683 1 A
port 11 n
rlabel metal1 205 575 239 609 1 A
port 12 n
rlabel metal1 205 501 239 535 1 A
port 13 n
rlabel metal1 205 427 239 461 1 A
port 14 n
rlabel metal1 427 871 461 905 1 B
port 15 n
rlabel metal1 427 797 461 831 1 B
port 16 n
rlabel metal1 427 723 461 757 1 B
port 17 n
rlabel metal1 427 649 461 683 1 B
port 18 n
rlabel metal1 427 575 461 609 1 B
port 19 n
rlabel metal1 427 501 461 535 1 B
port 20 n
rlabel metal1 427 427 461 461 1 B
port 21 n
rlabel metal1 649 871 683 905 1 C
port 22 n
rlabel metal1 649 797 683 831 1 C
port 23 n
rlabel metal1 649 723 683 757 1 C
port 24 n
rlabel metal1 649 649 683 683 1 C
port 25 n
rlabel metal1 649 575 683 609 1 C
port 26 n
rlabel metal1 649 501 683 535 1 C
port 27 n
rlabel metal1 649 427 683 461 1 C
port 28 n
rlabel metal1 -34 1446 1440 1514 1 VPWR
port 29 n
rlabel metal1 -34 -34 1440 34 1 VGND
port 30 n
rlabel nwell 57 1463 91 1497 1 VPB
port 31 n
rlabel pwell 57 -17 91 17 1 VNB
port 32 n
<< end >>
