* SPICE3 file created from DFFQNX1.ext - technology: sky130A

.subckt DFFQNX1 QN D CLK VDD GND
X0 VDD CLK a_277_1004 VDD pshort w=2 l=0.15 M=2
X1 QN a_3303_383 a_3072_73 GND nshort w=3 l=0.15
X2 VDD CLK a_147_159 VDD pshort w=2 l=0.15 M=2
X3 QN a_3303_383 VDD VDD pshort w=2 l=0.15 M=2
X4 GND a_147_159 a_91_75 GND nshort w=3 l=0.15
X5 VDD a_599_943 a_277_1004 VDD pshort w=2 l=0.15 M=2
X6 VDD a_277_1004 a_599_943 VDD pshort w=2 l=0.15 M=2
X7 a_3303_383 QN VDD VDD pshort w=2 l=0.15 M=2
X8 a_1845_1004 a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X9 VDD a_147_159 a_3303_383 VDD pshort w=2 l=0.15 M=2
X10 GND a_599_943 a_1740_73 GND nshort w=3 l=0.15
X11 a_372_182 CLK a_91_75 GND nshort w=3 l=0.15
X12 a_277_1004 a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X13 VDD D a_599_943 VDD pshort w=2 l=0.15 M=2
X14 a_147_159 CLK a_2406_73 GND nshort w=3 l=0.15
X15 VDD a_599_943 a_1845_1004 VDD pshort w=2 l=0.15 M=2
X16 GND QN a_3738_73 GND nshort w=3 l=0.15
X17 GND a_277_1004 a_1074_73 GND nshort w=3 l=0.15
X18 VDD a_277_1004 QN VDD pshort w=2 l=0.15 M=2
X19 a_1845_1004 a_147_159 a_1740_73 GND nshort w=3 l=0.15
X20 a_147_159 a_1845_1004 VDD VDD pshort w=2 l=0.15 M=2
X21 GND a_277_1004 a_3072_73 GND nshort w=3 l=0.15
X22 a_3303_383 a_147_159 a_3738_73 GND nshort w=3 l=0.15
X23 a_599_943 D a_1074_73 GND nshort w=3 l=0.15
X24 a_277_1004 a_599_943 a_372_182 GND nshort w=3 l=0.15
X25 GND a_1845_1004 a_2406_73 GND nshort w=3 l=0.15
C0 a_147_159 CLK 2.97fF
C1 a_277_1004 a_147_159 3.01fF
C2 a_277_1004 VDD 2.30fF
C3 a_147_159 VDD 3.14fF
C4 VDD GND 10.49fF
.ends
