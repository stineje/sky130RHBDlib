* SPICE3 file created from TMRDFFSNQX1.ext - technology: sky130A

.subckt TMRDFFSNQX1 Q D CLK SN VDD GND
M1000 a_8357_1050.t2 a_8483_411.t7 VDD.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_3599_411.t3 a_3473_1050.t5 VDD.t93 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t51 CLK.t0 a_6149_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t25 a_8483_411.t8 a_14869_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 GND a_11673_1050.t7 a_12470_101.t0 nshort w=-1.605u l=1.765u
+  ad=4.9019p pd=41.07u as=0p ps=0u
M1005 Q.t1 a_15044_209.t7 VDD.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_343_411.t3 a_1265_989.t5 VDD.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_13367_411.t3 a_11033_989.t5 VDD.t52 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t65 a_343_411.t7 a_3473_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_5227_411.t6 a_5101_1050.t5 VDD.t70 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VDD.t38 SN.t2 a_8483_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1265_989.t1 CLK.t1 VDD.t63 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 GND a_8483_411.t9 a_15430_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1013 VDD.t72 SN.t3 a_1905_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_11673_1050.t1 a_9985_1050.t6 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD.t81 CLK.t2 a_5227_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_15533_1051.t3 a_3599_411.t7 a_15044_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_3599_411.t6 SN.t4 VDD.t46 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 GND a_217_1050.t5 a_757_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 VDD.t9 CLK.t4 a_11033_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 GND D.t2 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t27 a_8357_1050.t5 a_8483_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_5227_411.t0 CLK.t5 VDD.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 GND a_343_411.t8 a_3368_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 VDD.t31 D.t0 a_5101_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_14869_1051.t0 a_3599_411.t8 a_15533_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VDD.t14 D.t1 a_217_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VDD.t67 a_1265_989.t7 a_1905_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_9985_1050.t4 a_10111_411.t7 VDD.t60 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 GND a_8357_1050.t6 a_8897_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1030 VDD.t16 a_5101_1050.t6 a_6789_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_15533_1051.t5 a_13367_411.t8 a_15044_209.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 VDD.t87 a_11033_989.t7 a_11673_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_3599_411.t4 a_1265_989.t9 VDD.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_6789_1050.t1 a_6149_989.t5 VDD.t95 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_13241_1050.t4 a_10111_411.t8 VDD.t89 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1905_1050.t6 a_217_1050.t6 VDD.t61 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VDD.t36 a_11673_1050.t8 a_11033_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_14869_1051.t4 a_8483_411.t10 a_15533_1051.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VDD.t29 a_343_411.t9 a_217_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 VDD.t88 a_5227_411.t8 a_5101_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 GND D.t3 a_9880_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1042 VDD.t55 a_217_1050.t7 a_343_411.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_11673_1050.t2 a_11033_989.t8 VDD.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 VDD.t33 a_13241_1050.t5 a_13367_411.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 GND a_217_1050.t8 a_1719_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_3473_1050.t4 a_3599_411.t9 VDD.t94 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_10111_411.t3 CLK.t7 VDD.t48 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_5227_411.t3 a_6149_989.t8 VDD.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_13241_1050.t2 a_13367_411.t10 VDD.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 VDD.t57 a_11033_989.t9 a_10111_411.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 VDD.t5 a_5227_411.t9 a_8357_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 a_6149_989.t0 CLK.t8 VDD.t86 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_14869_1051.t2 a_8483_411.t11 VDD.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 VDD.t62 a_6149_989.t9 a_8483_411.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_13367_411.t6 a_13241_1050.t6 VDD.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 VDD.t42 a_13367_411.t11 a_14869_1051.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 VDD.t17 CLK.t9 a_343_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 GND a_10111_411.t11 a_13136_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1059 GND a_1905_1050.t8 a_2702_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1060 a_3473_1050.t1 a_343_411.t10 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 VDD.t18 a_1905_1050.t7 a_1265_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_8483_411.t5 SN.t7 VDD.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 VDD.t47 SN.t8 a_13367_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_10111_411.t1 a_9985_1050.t7 VDD.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 GND a_13241_1050.t7 a_13781_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1066 GND a_5227_411.t10 a_8252_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_15533_1051.t6 a_8483_411.t12 a_14869_1051.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 VDD.t6 a_10111_411.t9 a_9985_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 Q a_15044_209.t9 GND.t5 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1070 VDD.t15 SN.t9 a_11673_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 GND a_5101_1050.t9 a_5641_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_6149_989.t4 a_6789_1050.t7 VDD.t90 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 VDD.t78 a_3473_1050.t6 a_3599_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 VDD.t10 a_1265_989.t10 a_3599_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 GND a_8483_411.t13 a_14764_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1076 VDD.t21 a_1265_989.t11 a_343_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 a_8483_411.t6 a_8357_1050.t7 VDD.t80 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 VDD.t3 a_15044_209.t8 Q.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VDD.t68 a_11033_989.t11 a_13367_411.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 VDD.t37 a_5101_1050.t7 a_5227_411.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 a_8483_411.t0 a_6149_989.t10 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 a_15533_1051.t0 a_3599_411.t11 a_14869_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_217_1050.t3 D.t4 VDD.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 VDD.t40 D.t5 a_9985_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_1905_1050.t0 a_1265_989.t12 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_6789_1050.t3 a_5101_1050.t8 VDD.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 VDD.t50 a_9985_1050.t8 a_11673_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 GND a_5101_1050.t10 a_6603_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_15044_209.t6 a_13367_411.t12 a_15533_1051.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 GND a_3473_1050.t7 a_4013_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1091 VDD.t77 SN.t12 a_3599_411.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 VDD.t79 SN.t13 a_6789_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_11033_989.t4 a_11673_1050.t9 VDD.t41 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 GND a_6789_1050.t9 a_7586_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1095 a_1905_1050.t3 SN.t14 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 a_217_1050.t0 a_343_411.t12 VDD.t64 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_5101_1050.t2 a_5227_411.t11 VDD.t58 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 GND a_9985_1050.t10 a_10525_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1099 GND a_3599_411.t14 a_16096_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1100 GND D.t7 a_4996_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1101 a_6789_1050.t5 SN.t15 VDD.t74 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_15044_209.t2 a_3599_411.t13 a_15533_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 VDD.t83 a_9985_1050.t9 a_10111_411.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_343_411.t5 a_217_1050.t9 VDD.t44 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 VDD.t26 a_8483_411.t14 a_8357_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VDD.t69 a_6149_989.t11 a_6789_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 a_10111_411.t4 a_11033_989.t13 VDD.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 VDD.t45 a_10111_411.t12 a_13241_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 VDD.t59 a_217_1050.t10 a_1905_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_8357_1050.t4 a_5227_411.t12 VDD.t43 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 VDD.t7 a_6789_1050.t8 a_6149_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1112 a_11033_989.t0 CLK.t13 VDD.t85 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 a_5101_1050.t1 D.t6 VDD.t32 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1114 a_14869_1051.t6 a_13367_411.t14 VDD.t39 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 a_343_411.t0 CLK.t14 VDD.t49 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 GND a_9985_1050.t5 a_11487_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_9985_1050.t0 D.t8 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_13367_411.t1 SN.t16 VDD.t92 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_1265_989.t4 a_1905_1050.t9 VDD.t53 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 VDD.t91 a_3599_411.t15 a_3473_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 VDD.t82 CLK.t15 a_10111_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 a_11673_1050.t5 SN.t17 VDD.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 VDD.t76 CLK.t17 a_1265_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1124 VDD.t34 a_6149_989.t13 a_5227_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1125 VDD.t54 a_13367_411.t15 a_13241_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 D SN 9.38fF
C1 VDD Q 0.76fF
C2 CLK SN 0.46fF
C3 VDD D 0.24fF
C4 VDD CLK 1.68fF
C5 D CLK 0.39fF
C6 VDD SN 0.30fF
R0 a_8483_411.n8 a_8483_411.t8 512.525
R1 a_8483_411.n6 a_8483_411.t10 477.179
R2 a_8483_411.n11 a_8483_411.t14 472.359
R3 a_8483_411.n6 a_8483_411.t12 406.485
R4 a_8483_411.n11 a_8483_411.t7 384.527
R5 a_8483_411.n8 a_8483_411.t11 371.139
R6 a_8483_411.n7 a_8483_411.t9 363.924
R7 a_8483_411.n10 a_8483_411.t13 277.053
R8 a_8483_411.n12 a_8483_411.t15 241.172
R9 a_8483_411.n16 a_8483_411.n14 213.104
R10 a_8483_411.n14 a_8483_411.n5 170.799
R11 a_8483_411.n12 a_8483_411.n11 110.06
R12 a_8483_411.n9 a_8483_411.n7 101.359
R13 a_8483_411.n13 a_8483_411.n10 94.999
R14 a_8483_411.n10 a_8483_411.n9 80.444
R15 a_8483_411.n13 a_8483_411.n12 80.035
R16 a_8483_411.n4 a_8483_411.n3 79.232
R17 a_8483_411.n14 a_8483_411.n13 76
R18 a_8483_411.n9 a_8483_411.n8 71.88
R19 a_8483_411.n5 a_8483_411.n4 63.152
R20 a_8483_411.n17 a_8483_411.n0 55.263
R21 a_8483_411.n16 a_8483_411.n15 30
R22 a_8483_411.n17 a_8483_411.n16 23.684
R23 a_8483_411.n5 a_8483_411.n1 16.08
R24 a_8483_411.n4 a_8483_411.n2 16.08
R25 a_8483_411.n7 a_8483_411.n6 15.776
R26 a_8483_411.n1 a_8483_411.t4 14.282
R27 a_8483_411.n1 a_8483_411.t0 14.282
R28 a_8483_411.n2 a_8483_411.t2 14.282
R29 a_8483_411.n2 a_8483_411.t5 14.282
R30 a_8483_411.n3 a_8483_411.t1 14.282
R31 a_8483_411.n3 a_8483_411.t6 14.282
R32 VDD.n839 VDD.n837 144.705
R33 VDD.n920 VDD.n918 144.705
R34 VDD.n1001 VDD.n999 144.705
R35 VDD.n1062 VDD.n1060 144.705
R36 VDD.n1123 VDD.n1121 144.705
R37 VDD.n1204 VDD.n1202 144.705
R38 VDD.n1265 VDD.n1263 144.705
R39 VDD.n1346 VDD.n1344 144.705
R40 VDD.n1427 VDD.n1425 144.705
R41 VDD.n744 VDD.n742 144.705
R42 VDD.n1488 VDD.n1486 144.705
R43 VDD.n663 VDD.n661 144.705
R44 VDD.n602 VDD.n600 144.705
R45 VDD.n521 VDD.n519 144.705
R46 VDD.n440 VDD.n438 144.705
R47 VDD.n379 VDD.n377 144.705
R48 VDD.n318 VDD.n316 144.705
R49 VDD.n237 VDD.n235 144.705
R50 VDD.n176 VDD.n174 144.705
R51 VDD.n122 VDD.n120 144.705
R52 VDD.n68 VDD.n66 144.705
R53 VDD.n26 VDD.n25 77.792
R54 VDD.n35 VDD.n34 77.792
R55 VDD.n29 VDD.n23 76.145
R56 VDD.n29 VDD.n28 76
R57 VDD.n33 VDD.n32 76
R58 VDD.n39 VDD.n38 76
R59 VDD.n43 VDD.n42 76
R60 VDD.n70 VDD.n69 76
R61 VDD.n74 VDD.n73 76
R62 VDD.n78 VDD.n77 76
R63 VDD.n82 VDD.n81 76
R64 VDD.n86 VDD.n85 76
R65 VDD.n90 VDD.n89 76
R66 VDD.n94 VDD.n93 76
R67 VDD.n98 VDD.n97 76
R68 VDD.n124 VDD.n123 76
R69 VDD.n128 VDD.n127 76
R70 VDD.n132 VDD.n131 76
R71 VDD.n136 VDD.n135 76
R72 VDD.n140 VDD.n139 76
R73 VDD.n144 VDD.n143 76
R74 VDD.n148 VDD.n147 76
R75 VDD.n152 VDD.n151 76
R76 VDD.n178 VDD.n177 76
R77 VDD.n183 VDD.n182 76
R78 VDD.n188 VDD.n187 76
R79 VDD.n194 VDD.n193 76
R80 VDD.n199 VDD.n198 76
R81 VDD.n204 VDD.n203 76
R82 VDD.n209 VDD.n208 76
R83 VDD.n213 VDD.n212 76
R84 VDD.n239 VDD.n238 76
R85 VDD.n243 VDD.n242 76
R86 VDD.n247 VDD.n246 76
R87 VDD.n252 VDD.n251 76
R88 VDD.n259 VDD.n258 76
R89 VDD.n264 VDD.n263 76
R90 VDD.n269 VDD.n268 76
R91 VDD.n276 VDD.n275 76
R92 VDD.n281 VDD.n280 76
R93 VDD.n286 VDD.n285 76
R94 VDD.n290 VDD.n289 76
R95 VDD.n294 VDD.n293 76
R96 VDD.n320 VDD.n319 76
R97 VDD.n325 VDD.n324 76
R98 VDD.n330 VDD.n329 76
R99 VDD.n336 VDD.n335 76
R100 VDD.n341 VDD.n340 76
R101 VDD.n346 VDD.n345 76
R102 VDD.n351 VDD.n350 76
R103 VDD.n355 VDD.n354 76
R104 VDD.n381 VDD.n380 76
R105 VDD.n386 VDD.n385 76
R106 VDD.n391 VDD.n390 76
R107 VDD.n397 VDD.n396 76
R108 VDD.n402 VDD.n401 76
R109 VDD.n407 VDD.n406 76
R110 VDD.n412 VDD.n411 76
R111 VDD.n416 VDD.n415 76
R112 VDD.n442 VDD.n441 76
R113 VDD.n446 VDD.n445 76
R114 VDD.n450 VDD.n449 76
R115 VDD.n455 VDD.n454 76
R116 VDD.n462 VDD.n461 76
R117 VDD.n467 VDD.n466 76
R118 VDD.n472 VDD.n471 76
R119 VDD.n479 VDD.n478 76
R120 VDD.n484 VDD.n483 76
R121 VDD.n489 VDD.n488 76
R122 VDD.n493 VDD.n492 76
R123 VDD.n497 VDD.n496 76
R124 VDD.n523 VDD.n522 76
R125 VDD.n527 VDD.n526 76
R126 VDD.n531 VDD.n530 76
R127 VDD.n536 VDD.n535 76
R128 VDD.n543 VDD.n542 76
R129 VDD.n548 VDD.n547 76
R130 VDD.n553 VDD.n552 76
R131 VDD.n560 VDD.n559 76
R132 VDD.n565 VDD.n564 76
R133 VDD.n570 VDD.n569 76
R134 VDD.n574 VDD.n573 76
R135 VDD.n578 VDD.n577 76
R136 VDD.n604 VDD.n603 76
R137 VDD.n609 VDD.n608 76
R138 VDD.n614 VDD.n613 76
R139 VDD.n620 VDD.n619 76
R140 VDD.n625 VDD.n624 76
R141 VDD.n630 VDD.n629 76
R142 VDD.n635 VDD.n634 76
R143 VDD.n639 VDD.n638 76
R144 VDD.n665 VDD.n664 76
R145 VDD.n669 VDD.n668 76
R146 VDD.n673 VDD.n672 76
R147 VDD.n678 VDD.n677 76
R148 VDD.n685 VDD.n684 76
R149 VDD.n690 VDD.n689 76
R150 VDD.n695 VDD.n694 76
R151 VDD.n702 VDD.n701 76
R152 VDD.n707 VDD.n706 76
R153 VDD.n712 VDD.n711 76
R154 VDD.n716 VDD.n715 76
R155 VDD.n720 VDD.n719 76
R156 VDD.n746 VDD.n745 76
R157 VDD.n751 VDD.n750 76
R158 VDD.n756 VDD.n755 76
R159 VDD.n1511 VDD.n1510 76
R160 VDD.n1505 VDD.n1504 76
R161 VDD.n1500 VDD.n1499 76
R162 VDD.n1495 VDD.n1494 76
R163 VDD.n1490 VDD.n1489 76
R164 VDD.n1464 VDD.n1463 76
R165 VDD.n1460 VDD.n1459 76
R166 VDD.n1455 VDD.n1454 76
R167 VDD.n1450 VDD.n1449 76
R168 VDD.n1444 VDD.n1443 76
R169 VDD.n1439 VDD.n1438 76
R170 VDD.n1434 VDD.n1433 76
R171 VDD.n1429 VDD.n1428 76
R172 VDD.n1403 VDD.n1402 76
R173 VDD.n1399 VDD.n1398 76
R174 VDD.n1395 VDD.n1394 76
R175 VDD.n1391 VDD.n1390 76
R176 VDD.n1386 VDD.n1385 76
R177 VDD.n1379 VDD.n1378 76
R178 VDD.n1374 VDD.n1373 76
R179 VDD.n1369 VDD.n1368 76
R180 VDD.n1362 VDD.n1361 76
R181 VDD.n1357 VDD.n1356 76
R182 VDD.n1352 VDD.n1351 76
R183 VDD.n1348 VDD.n1347 76
R184 VDD.n1322 VDD.n1321 76
R185 VDD.n1318 VDD.n1317 76
R186 VDD.n1314 VDD.n1313 76
R187 VDD.n1310 VDD.n1309 76
R188 VDD.n1305 VDD.n1304 76
R189 VDD.n1298 VDD.n1297 76
R190 VDD.n1293 VDD.n1292 76
R191 VDD.n1288 VDD.n1287 76
R192 VDD.n1281 VDD.n1280 76
R193 VDD.n1276 VDD.n1275 76
R194 VDD.n1271 VDD.n1270 76
R195 VDD.n1267 VDD.n1266 76
R196 VDD.n1241 VDD.n1240 76
R197 VDD.n1237 VDD.n1236 76
R198 VDD.n1232 VDD.n1231 76
R199 VDD.n1227 VDD.n1226 76
R200 VDD.n1221 VDD.n1220 76
R201 VDD.n1216 VDD.n1215 76
R202 VDD.n1211 VDD.n1210 76
R203 VDD.n1206 VDD.n1205 76
R204 VDD.n1180 VDD.n1179 76
R205 VDD.n1176 VDD.n1175 76
R206 VDD.n1172 VDD.n1171 76
R207 VDD.n1168 VDD.n1167 76
R208 VDD.n1163 VDD.n1162 76
R209 VDD.n1156 VDD.n1155 76
R210 VDD.n1151 VDD.n1150 76
R211 VDD.n1146 VDD.n1145 76
R212 VDD.n1139 VDD.n1138 76
R213 VDD.n1134 VDD.n1133 76
R214 VDD.n1129 VDD.n1128 76
R215 VDD.n1125 VDD.n1124 76
R216 VDD.n1099 VDD.n1098 76
R217 VDD.n1095 VDD.n1094 76
R218 VDD.n1090 VDD.n1089 76
R219 VDD.n1085 VDD.n1084 76
R220 VDD.n1079 VDD.n1078 76
R221 VDD.n1074 VDD.n1073 76
R222 VDD.n1069 VDD.n1068 76
R223 VDD.n1064 VDD.n1063 76
R224 VDD.n1038 VDD.n1037 76
R225 VDD.n1034 VDD.n1033 76
R226 VDD.n1029 VDD.n1028 76
R227 VDD.n1024 VDD.n1023 76
R228 VDD.n1018 VDD.n1017 76
R229 VDD.n1013 VDD.n1012 76
R230 VDD.n1008 VDD.n1007 76
R231 VDD.n1003 VDD.n1002 76
R232 VDD.n977 VDD.n976 76
R233 VDD.n973 VDD.n972 76
R234 VDD.n969 VDD.n968 76
R235 VDD.n965 VDD.n964 76
R236 VDD.n960 VDD.n959 76
R237 VDD.n953 VDD.n952 76
R238 VDD.n948 VDD.n947 76
R239 VDD.n943 VDD.n942 76
R240 VDD.n936 VDD.n935 76
R241 VDD.n931 VDD.n930 76
R242 VDD.n926 VDD.n925 76
R243 VDD.n922 VDD.n921 76
R244 VDD.n896 VDD.n895 76
R245 VDD.n892 VDD.n891 76
R246 VDD.n888 VDD.n887 76
R247 VDD.n884 VDD.n883 76
R248 VDD.n879 VDD.n878 76
R249 VDD.n872 VDD.n871 76
R250 VDD.n867 VDD.n866 76
R251 VDD.n862 VDD.n861 76
R252 VDD.n855 VDD.n854 76
R253 VDD.n850 VDD.n849 76
R254 VDD.n845 VDD.n844 76
R255 VDD.n841 VDD.n840 76
R256 VDD.n814 VDD.n813 76
R257 VDD.n810 VDD.n809 76
R258 VDD.n805 VDD.n804 76
R259 VDD.n800 VDD.n799 76
R260 VDD.n794 VDD.n793 76
R261 VDD.n789 VDD.n788 76
R262 VDD.n784 VDD.n783 76
R263 VDD.n779 VDD.n778 76
R264 VDD.n249 VDD.n248 64.064
R265 VDD.n452 VDD.n451 64.064
R266 VDD.n533 VDD.n532 64.064
R267 VDD.n675 VDD.n674 64.064
R268 VDD.n1388 VDD.n1387 64.064
R269 VDD.n1307 VDD.n1306 64.064
R270 VDD.n1165 VDD.n1164 64.064
R271 VDD.n962 VDD.n961 64.064
R272 VDD.n881 VDD.n880 64.064
R273 VDD.n278 VDD.n277 59.488
R274 VDD.n481 VDD.n480 59.488
R275 VDD.n562 VDD.n561 59.488
R276 VDD.n704 VDD.n703 59.488
R277 VDD.n1359 VDD.n1358 59.488
R278 VDD.n1278 VDD.n1277 59.488
R279 VDD.n1136 VDD.n1135 59.488
R280 VDD.n933 VDD.n932 59.488
R281 VDD.n852 VDD.n851 59.488
R282 VDD.n205 VDD.t23 55.465
R283 VDD.n179 VDD.t42 55.465
R284 VDD.n780 VDD.t35 55.106
R285 VDD.n846 VDD.t44 55.106
R286 VDD.n927 VDD.t61 55.106
R287 VDD.n1004 VDD.t53 55.106
R288 VDD.n1065 VDD.t12 55.106
R289 VDD.n1130 VDD.t93 55.106
R290 VDD.n1207 VDD.t32 55.106
R291 VDD.n1272 VDD.t70 55.106
R292 VDD.n1353 VDD.t22 55.106
R293 VDD.n1430 VDD.t90 55.106
R294 VDD.n1491 VDD.t43 55.106
R295 VDD.n708 VDD.t80 55.106
R296 VDD.n631 VDD.t0 55.106
R297 VDD.n566 VDD.t56 55.106
R298 VDD.n485 VDD.t2 55.106
R299 VDD.n408 VDD.t41 55.106
R300 VDD.n347 VDD.t89 55.106
R301 VDD.n282 VDD.t71 55.106
R302 VDD.n37 VDD.t20 55.106
R303 VDD.n24 VDD.t3 55.106
R304 VDD.n887 VDD.t21 55.106
R305 VDD.n968 VDD.t67 55.106
R306 VDD.n1171 VDD.t10 55.106
R307 VDD.n1313 VDD.t34 55.106
R308 VDD.n1394 VDD.t69 55.106
R309 VDD.n672 VDD.t62 55.106
R310 VDD.n530 VDD.t57 55.106
R311 VDD.n449 VDD.t87 55.106
R312 VDD.n246 VDD.t68 55.106
R313 VDD.n806 VDD.t29 55.106
R314 VDD.n1030 VDD.t76 55.106
R315 VDD.n1091 VDD.t91 55.106
R316 VDD.n1233 VDD.t88 55.106
R317 VDD.n1456 VDD.t51 55.106
R318 VDD.n747 VDD.t26 55.106
R319 VDD.n605 VDD.t6 55.106
R320 VDD.n382 VDD.t9 55.106
R321 VDD.n321 VDD.t54 55.106
R322 VDD.n190 VDD.n189 41.183
R323 VDD.n796 VDD.n795 40.824
R324 VDD.n857 VDD.n856 40.824
R325 VDD.n877 VDD.n876 40.824
R326 VDD.n938 VDD.n937 40.824
R327 VDD.n958 VDD.n957 40.824
R328 VDD.n1020 VDD.n1019 40.824
R329 VDD.n1081 VDD.n1080 40.824
R330 VDD.n1141 VDD.n1140 40.824
R331 VDD.n1161 VDD.n1160 40.824
R332 VDD.n1223 VDD.n1222 40.824
R333 VDD.n1283 VDD.n1282 40.824
R334 VDD.n1303 VDD.n1302 40.824
R335 VDD.n1364 VDD.n1363 40.824
R336 VDD.n1384 VDD.n1383 40.824
R337 VDD.n1446 VDD.n1445 40.824
R338 VDD.n1507 VDD.n1506 40.824
R339 VDD.n697 VDD.n696 40.824
R340 VDD.n683 VDD.n682 40.824
R341 VDD.n616 VDD.n615 40.824
R342 VDD.n555 VDD.n554 40.824
R343 VDD.n541 VDD.n540 40.824
R344 VDD.n474 VDD.n473 40.824
R345 VDD.n460 VDD.n459 40.824
R346 VDD.n393 VDD.n392 40.824
R347 VDD.n332 VDD.n331 40.824
R348 VDD.n271 VDD.n270 40.824
R349 VDD.n257 VDD.n256 40.824
R350 VDD.n901 VDD.n900 36.774
R351 VDD.n982 VDD.n981 36.774
R352 VDD.n1043 VDD.n1042 36.774
R353 VDD.n1104 VDD.n1103 36.774
R354 VDD.n1185 VDD.n1184 36.774
R355 VDD.n1246 VDD.n1245 36.774
R356 VDD.n1327 VDD.n1326 36.774
R357 VDD.n1408 VDD.n1407 36.774
R358 VDD.n1469 VDD.n1468 36.774
R359 VDD.n725 VDD.n724 36.774
R360 VDD.n644 VDD.n643 36.774
R361 VDD.n583 VDD.n582 36.774
R362 VDD.n502 VDD.n501 36.774
R363 VDD.n421 VDD.n420 36.774
R364 VDD.n360 VDD.n359 36.774
R365 VDD.n299 VDD.n298 36.774
R366 VDD.n218 VDD.n217 36.774
R367 VDD.n157 VDD.n156 36.774
R368 VDD.n103 VDD.n102 36.774
R369 VDD.n48 VDD.n47 36.774
R370 VDD.n830 VDD.n829 36.774
R371 VDD.n185 VDD.n184 36.608
R372 VDD.n327 VDD.n326 36.608
R373 VDD.n388 VDD.n387 36.608
R374 VDD.n611 VDD.n610 36.608
R375 VDD.n753 VDD.n752 36.608
R376 VDD.n1452 VDD.n1451 36.608
R377 VDD.n1229 VDD.n1228 36.608
R378 VDD.n1087 VDD.n1086 36.608
R379 VDD.n1026 VDD.n1025 36.608
R380 VDD.n802 VDD.n801 36.608
R381 VDD.n201 VDD.n200 32.032
R382 VDD.n343 VDD.n342 32.032
R383 VDD.n404 VDD.n403 32.032
R384 VDD.n627 VDD.n626 32.032
R385 VDD.n1497 VDD.n1496 32.032
R386 VDD.n1436 VDD.n1435 32.032
R387 VDD.n1213 VDD.n1212 32.032
R388 VDD.n1071 VDD.n1070 32.032
R389 VDD.n1010 VDD.n1009 32.032
R390 VDD.n786 VDD.n785 32.032
R391 VDD.n254 VDD.n253 27.456
R392 VDD.n457 VDD.n456 27.456
R393 VDD.n538 VDD.n537 27.456
R394 VDD.n680 VDD.n679 27.456
R395 VDD.n1381 VDD.n1380 27.456
R396 VDD.n1300 VDD.n1299 27.456
R397 VDD.n1158 VDD.n1157 27.456
R398 VDD.n955 VDD.n954 27.456
R399 VDD.n874 VDD.n873 27.456
R400 VDD.n273 VDD.n272 22.88
R401 VDD.n476 VDD.n475 22.88
R402 VDD.n557 VDD.n556 22.88
R403 VDD.n699 VDD.n698 22.88
R404 VDD.n1366 VDD.n1365 22.88
R405 VDD.n1285 VDD.n1284 22.88
R406 VDD.n1143 VDD.n1142 22.88
R407 VDD.n940 VDD.n939 22.88
R408 VDD.n859 VDD.n858 22.88
R409 VDD.n778 VDD.n775 21.841
R410 VDD.n23 VDD.n20 21.841
R411 VDD.n795 VDD.t64 14.282
R412 VDD.n795 VDD.t14 14.282
R413 VDD.n856 VDD.t49 14.282
R414 VDD.n856 VDD.t55 14.282
R415 VDD.n876 VDD.t11 14.282
R416 VDD.n876 VDD.t17 14.282
R417 VDD.n937 VDD.t8 14.282
R418 VDD.n937 VDD.t59 14.282
R419 VDD.n957 VDD.t4 14.282
R420 VDD.n957 VDD.t72 14.282
R421 VDD.n1019 VDD.t63 14.282
R422 VDD.n1019 VDD.t18 14.282
R423 VDD.n1080 VDD.t94 14.282
R424 VDD.n1080 VDD.t65 14.282
R425 VDD.n1140 VDD.t46 14.282
R426 VDD.n1140 VDD.t78 14.282
R427 VDD.n1160 VDD.t28 14.282
R428 VDD.n1160 VDD.t77 14.282
R429 VDD.n1222 VDD.t58 14.282
R430 VDD.n1222 VDD.t31 14.282
R431 VDD.n1282 VDD.t19 14.282
R432 VDD.n1282 VDD.t37 14.282
R433 VDD.n1302 VDD.t84 14.282
R434 VDD.n1302 VDD.t81 14.282
R435 VDD.n1363 VDD.t74 14.282
R436 VDD.n1363 VDD.t16 14.282
R437 VDD.n1383 VDD.t95 14.282
R438 VDD.n1383 VDD.t79 14.282
R439 VDD.n1445 VDD.t86 14.282
R440 VDD.n1445 VDD.t7 14.282
R441 VDD.n1506 VDD.t24 14.282
R442 VDD.n1506 VDD.t5 14.282
R443 VDD.n696 VDD.t73 14.282
R444 VDD.n696 VDD.t27 14.282
R445 VDD.n682 VDD.t1 14.282
R446 VDD.n682 VDD.t38 14.282
R447 VDD.n615 VDD.t60 14.282
R448 VDD.n615 VDD.t40 14.282
R449 VDD.n554 VDD.t48 14.282
R450 VDD.n554 VDD.t83 14.282
R451 VDD.n540 VDD.t30 14.282
R452 VDD.n540 VDD.t82 14.282
R453 VDD.n473 VDD.t75 14.282
R454 VDD.n473 VDD.t50 14.282
R455 VDD.n459 VDD.t13 14.282
R456 VDD.n459 VDD.t15 14.282
R457 VDD.n392 VDD.t85 14.282
R458 VDD.n392 VDD.t36 14.282
R459 VDD.n331 VDD.t66 14.282
R460 VDD.n331 VDD.t45 14.282
R461 VDD.n270 VDD.t92 14.282
R462 VDD.n270 VDD.t33 14.282
R463 VDD.n256 VDD.t52 14.282
R464 VDD.n256 VDD.t47 14.282
R465 VDD.n189 VDD.t39 14.282
R466 VDD.n189 VDD.t25 14.282
R467 VDD.n775 VDD.n758 14.167
R468 VDD.n758 VDD.n757 14.167
R469 VDD.n916 VDD.n898 14.167
R470 VDD.n898 VDD.n897 14.167
R471 VDD.n997 VDD.n979 14.167
R472 VDD.n979 VDD.n978 14.167
R473 VDD.n1058 VDD.n1040 14.167
R474 VDD.n1040 VDD.n1039 14.167
R475 VDD.n1119 VDD.n1101 14.167
R476 VDD.n1101 VDD.n1100 14.167
R477 VDD.n1200 VDD.n1182 14.167
R478 VDD.n1182 VDD.n1181 14.167
R479 VDD.n1261 VDD.n1243 14.167
R480 VDD.n1243 VDD.n1242 14.167
R481 VDD.n1342 VDD.n1324 14.167
R482 VDD.n1324 VDD.n1323 14.167
R483 VDD.n1423 VDD.n1405 14.167
R484 VDD.n1405 VDD.n1404 14.167
R485 VDD.n1484 VDD.n1466 14.167
R486 VDD.n1466 VDD.n1465 14.167
R487 VDD.n740 VDD.n722 14.167
R488 VDD.n722 VDD.n721 14.167
R489 VDD.n659 VDD.n641 14.167
R490 VDD.n641 VDD.n640 14.167
R491 VDD.n598 VDD.n580 14.167
R492 VDD.n580 VDD.n579 14.167
R493 VDD.n517 VDD.n499 14.167
R494 VDD.n499 VDD.n498 14.167
R495 VDD.n436 VDD.n418 14.167
R496 VDD.n418 VDD.n417 14.167
R497 VDD.n375 VDD.n357 14.167
R498 VDD.n357 VDD.n356 14.167
R499 VDD.n314 VDD.n296 14.167
R500 VDD.n296 VDD.n295 14.167
R501 VDD.n233 VDD.n215 14.167
R502 VDD.n215 VDD.n214 14.167
R503 VDD.n172 VDD.n154 14.167
R504 VDD.n154 VDD.n153 14.167
R505 VDD.n118 VDD.n100 14.167
R506 VDD.n100 VDD.n99 14.167
R507 VDD.n64 VDD.n45 14.167
R508 VDD.n45 VDD.n44 14.167
R509 VDD.n835 VDD.n816 14.167
R510 VDD.n816 VDD.n815 14.167
R511 VDD.n20 VDD.n19 14.167
R512 VDD.n19 VDD.n17 14.167
R513 VDD.n69 VDD.n65 14.167
R514 VDD.n123 VDD.n119 14.167
R515 VDD.n177 VDD.n173 14.167
R516 VDD.n238 VDD.n234 14.167
R517 VDD.n319 VDD.n315 14.167
R518 VDD.n380 VDD.n376 14.167
R519 VDD.n441 VDD.n437 14.167
R520 VDD.n522 VDD.n518 14.167
R521 VDD.n603 VDD.n599 14.167
R522 VDD.n664 VDD.n660 14.167
R523 VDD.n745 VDD.n741 14.167
R524 VDD.n1489 VDD.n1485 14.167
R525 VDD.n1428 VDD.n1424 14.167
R526 VDD.n1347 VDD.n1343 14.167
R527 VDD.n1266 VDD.n1262 14.167
R528 VDD.n1205 VDD.n1201 14.167
R529 VDD.n1124 VDD.n1120 14.167
R530 VDD.n1063 VDD.n1059 14.167
R531 VDD.n1002 VDD.n998 14.167
R532 VDD.n921 VDD.n917 14.167
R533 VDD.n840 VDD.n836 14.167
R534 VDD.n266 VDD.n265 13.728
R535 VDD.n469 VDD.n468 13.728
R536 VDD.n550 VDD.n549 13.728
R537 VDD.n692 VDD.n691 13.728
R538 VDD.n1371 VDD.n1370 13.728
R539 VDD.n1290 VDD.n1289 13.728
R540 VDD.n1148 VDD.n1147 13.728
R541 VDD.n945 VDD.n944 13.728
R542 VDD.n864 VDD.n863 13.728
R543 VDD.n23 VDD.n22 13.653
R544 VDD.n22 VDD.n21 13.653
R545 VDD.n28 VDD.n27 13.653
R546 VDD.n27 VDD.n26 13.653
R547 VDD.n32 VDD.n31 13.653
R548 VDD.n31 VDD.n30 13.653
R549 VDD.n38 VDD.n36 13.653
R550 VDD.n36 VDD.n35 13.653
R551 VDD.n42 VDD.n41 13.653
R552 VDD.n41 VDD.n40 13.653
R553 VDD.n69 VDD.n68 13.653
R554 VDD.n68 VDD.n67 13.653
R555 VDD.n73 VDD.n72 13.653
R556 VDD.n72 VDD.n71 13.653
R557 VDD.n77 VDD.n76 13.653
R558 VDD.n76 VDD.n75 13.653
R559 VDD.n81 VDD.n80 13.653
R560 VDD.n80 VDD.n79 13.653
R561 VDD.n85 VDD.n84 13.653
R562 VDD.n84 VDD.n83 13.653
R563 VDD.n89 VDD.n88 13.653
R564 VDD.n88 VDD.n87 13.653
R565 VDD.n93 VDD.n92 13.653
R566 VDD.n92 VDD.n91 13.653
R567 VDD.n97 VDD.n96 13.653
R568 VDD.n96 VDD.n95 13.653
R569 VDD.n123 VDD.n122 13.653
R570 VDD.n122 VDD.n121 13.653
R571 VDD.n127 VDD.n126 13.653
R572 VDD.n126 VDD.n125 13.653
R573 VDD.n131 VDD.n130 13.653
R574 VDD.n130 VDD.n129 13.653
R575 VDD.n135 VDD.n134 13.653
R576 VDD.n134 VDD.n133 13.653
R577 VDD.n139 VDD.n138 13.653
R578 VDD.n138 VDD.n137 13.653
R579 VDD.n143 VDD.n142 13.653
R580 VDD.n142 VDD.n141 13.653
R581 VDD.n147 VDD.n146 13.653
R582 VDD.n146 VDD.n145 13.653
R583 VDD.n151 VDD.n150 13.653
R584 VDD.n150 VDD.n149 13.653
R585 VDD.n177 VDD.n176 13.653
R586 VDD.n176 VDD.n175 13.653
R587 VDD.n182 VDD.n181 13.653
R588 VDD.n181 VDD.n180 13.653
R589 VDD.n187 VDD.n186 13.653
R590 VDD.n186 VDD.n185 13.653
R591 VDD.n193 VDD.n192 13.653
R592 VDD.n192 VDD.n191 13.653
R593 VDD.n198 VDD.n197 13.653
R594 VDD.n197 VDD.n196 13.653
R595 VDD.n203 VDD.n202 13.653
R596 VDD.n202 VDD.n201 13.653
R597 VDD.n208 VDD.n207 13.653
R598 VDD.n207 VDD.n206 13.653
R599 VDD.n212 VDD.n211 13.653
R600 VDD.n211 VDD.n210 13.653
R601 VDD.n238 VDD.n237 13.653
R602 VDD.n237 VDD.n236 13.653
R603 VDD.n242 VDD.n241 13.653
R604 VDD.n241 VDD.n240 13.653
R605 VDD.n246 VDD.n245 13.653
R606 VDD.n245 VDD.n244 13.653
R607 VDD.n251 VDD.n250 13.653
R608 VDD.n250 VDD.n249 13.653
R609 VDD.n258 VDD.n255 13.653
R610 VDD.n255 VDD.n254 13.653
R611 VDD.n263 VDD.n262 13.653
R612 VDD.n262 VDD.n261 13.653
R613 VDD.n268 VDD.n267 13.653
R614 VDD.n267 VDD.n266 13.653
R615 VDD.n275 VDD.n274 13.653
R616 VDD.n274 VDD.n273 13.653
R617 VDD.n280 VDD.n279 13.653
R618 VDD.n279 VDD.n278 13.653
R619 VDD.n285 VDD.n284 13.653
R620 VDD.n284 VDD.n283 13.653
R621 VDD.n289 VDD.n288 13.653
R622 VDD.n288 VDD.n287 13.653
R623 VDD.n293 VDD.n292 13.653
R624 VDD.n292 VDD.n291 13.653
R625 VDD.n319 VDD.n318 13.653
R626 VDD.n318 VDD.n317 13.653
R627 VDD.n324 VDD.n323 13.653
R628 VDD.n323 VDD.n322 13.653
R629 VDD.n329 VDD.n328 13.653
R630 VDD.n328 VDD.n327 13.653
R631 VDD.n335 VDD.n334 13.653
R632 VDD.n334 VDD.n333 13.653
R633 VDD.n340 VDD.n339 13.653
R634 VDD.n339 VDD.n338 13.653
R635 VDD.n345 VDD.n344 13.653
R636 VDD.n344 VDD.n343 13.653
R637 VDD.n350 VDD.n349 13.653
R638 VDD.n349 VDD.n348 13.653
R639 VDD.n354 VDD.n353 13.653
R640 VDD.n353 VDD.n352 13.653
R641 VDD.n380 VDD.n379 13.653
R642 VDD.n379 VDD.n378 13.653
R643 VDD.n385 VDD.n384 13.653
R644 VDD.n384 VDD.n383 13.653
R645 VDD.n390 VDD.n389 13.653
R646 VDD.n389 VDD.n388 13.653
R647 VDD.n396 VDD.n395 13.653
R648 VDD.n395 VDD.n394 13.653
R649 VDD.n401 VDD.n400 13.653
R650 VDD.n400 VDD.n399 13.653
R651 VDD.n406 VDD.n405 13.653
R652 VDD.n405 VDD.n404 13.653
R653 VDD.n411 VDD.n410 13.653
R654 VDD.n410 VDD.n409 13.653
R655 VDD.n415 VDD.n414 13.653
R656 VDD.n414 VDD.n413 13.653
R657 VDD.n441 VDD.n440 13.653
R658 VDD.n440 VDD.n439 13.653
R659 VDD.n445 VDD.n444 13.653
R660 VDD.n444 VDD.n443 13.653
R661 VDD.n449 VDD.n448 13.653
R662 VDD.n448 VDD.n447 13.653
R663 VDD.n454 VDD.n453 13.653
R664 VDD.n453 VDD.n452 13.653
R665 VDD.n461 VDD.n458 13.653
R666 VDD.n458 VDD.n457 13.653
R667 VDD.n466 VDD.n465 13.653
R668 VDD.n465 VDD.n464 13.653
R669 VDD.n471 VDD.n470 13.653
R670 VDD.n470 VDD.n469 13.653
R671 VDD.n478 VDD.n477 13.653
R672 VDD.n477 VDD.n476 13.653
R673 VDD.n483 VDD.n482 13.653
R674 VDD.n482 VDD.n481 13.653
R675 VDD.n488 VDD.n487 13.653
R676 VDD.n487 VDD.n486 13.653
R677 VDD.n492 VDD.n491 13.653
R678 VDD.n491 VDD.n490 13.653
R679 VDD.n496 VDD.n495 13.653
R680 VDD.n495 VDD.n494 13.653
R681 VDD.n522 VDD.n521 13.653
R682 VDD.n521 VDD.n520 13.653
R683 VDD.n526 VDD.n525 13.653
R684 VDD.n525 VDD.n524 13.653
R685 VDD.n530 VDD.n529 13.653
R686 VDD.n529 VDD.n528 13.653
R687 VDD.n535 VDD.n534 13.653
R688 VDD.n534 VDD.n533 13.653
R689 VDD.n542 VDD.n539 13.653
R690 VDD.n539 VDD.n538 13.653
R691 VDD.n547 VDD.n546 13.653
R692 VDD.n546 VDD.n545 13.653
R693 VDD.n552 VDD.n551 13.653
R694 VDD.n551 VDD.n550 13.653
R695 VDD.n559 VDD.n558 13.653
R696 VDD.n558 VDD.n557 13.653
R697 VDD.n564 VDD.n563 13.653
R698 VDD.n563 VDD.n562 13.653
R699 VDD.n569 VDD.n568 13.653
R700 VDD.n568 VDD.n567 13.653
R701 VDD.n573 VDD.n572 13.653
R702 VDD.n572 VDD.n571 13.653
R703 VDD.n577 VDD.n576 13.653
R704 VDD.n576 VDD.n575 13.653
R705 VDD.n603 VDD.n602 13.653
R706 VDD.n602 VDD.n601 13.653
R707 VDD.n608 VDD.n607 13.653
R708 VDD.n607 VDD.n606 13.653
R709 VDD.n613 VDD.n612 13.653
R710 VDD.n612 VDD.n611 13.653
R711 VDD.n619 VDD.n618 13.653
R712 VDD.n618 VDD.n617 13.653
R713 VDD.n624 VDD.n623 13.653
R714 VDD.n623 VDD.n622 13.653
R715 VDD.n629 VDD.n628 13.653
R716 VDD.n628 VDD.n627 13.653
R717 VDD.n634 VDD.n633 13.653
R718 VDD.n633 VDD.n632 13.653
R719 VDD.n638 VDD.n637 13.653
R720 VDD.n637 VDD.n636 13.653
R721 VDD.n664 VDD.n663 13.653
R722 VDD.n663 VDD.n662 13.653
R723 VDD.n668 VDD.n667 13.653
R724 VDD.n667 VDD.n666 13.653
R725 VDD.n672 VDD.n671 13.653
R726 VDD.n671 VDD.n670 13.653
R727 VDD.n677 VDD.n676 13.653
R728 VDD.n676 VDD.n675 13.653
R729 VDD.n684 VDD.n681 13.653
R730 VDD.n681 VDD.n680 13.653
R731 VDD.n689 VDD.n688 13.653
R732 VDD.n688 VDD.n687 13.653
R733 VDD.n694 VDD.n693 13.653
R734 VDD.n693 VDD.n692 13.653
R735 VDD.n701 VDD.n700 13.653
R736 VDD.n700 VDD.n699 13.653
R737 VDD.n706 VDD.n705 13.653
R738 VDD.n705 VDD.n704 13.653
R739 VDD.n711 VDD.n710 13.653
R740 VDD.n710 VDD.n709 13.653
R741 VDD.n715 VDD.n714 13.653
R742 VDD.n714 VDD.n713 13.653
R743 VDD.n719 VDD.n718 13.653
R744 VDD.n718 VDD.n717 13.653
R745 VDD.n745 VDD.n744 13.653
R746 VDD.n744 VDD.n743 13.653
R747 VDD.n750 VDD.n749 13.653
R748 VDD.n749 VDD.n748 13.653
R749 VDD.n755 VDD.n754 13.653
R750 VDD.n754 VDD.n753 13.653
R751 VDD.n1510 VDD.n1509 13.653
R752 VDD.n1509 VDD.n1508 13.653
R753 VDD.n1504 VDD.n1503 13.653
R754 VDD.n1503 VDD.n1502 13.653
R755 VDD.n1499 VDD.n1498 13.653
R756 VDD.n1498 VDD.n1497 13.653
R757 VDD.n1494 VDD.n1493 13.653
R758 VDD.n1493 VDD.n1492 13.653
R759 VDD.n1489 VDD.n1488 13.653
R760 VDD.n1488 VDD.n1487 13.653
R761 VDD.n1463 VDD.n1462 13.653
R762 VDD.n1462 VDD.n1461 13.653
R763 VDD.n1459 VDD.n1458 13.653
R764 VDD.n1458 VDD.n1457 13.653
R765 VDD.n1454 VDD.n1453 13.653
R766 VDD.n1453 VDD.n1452 13.653
R767 VDD.n1449 VDD.n1448 13.653
R768 VDD.n1448 VDD.n1447 13.653
R769 VDD.n1443 VDD.n1442 13.653
R770 VDD.n1442 VDD.n1441 13.653
R771 VDD.n1438 VDD.n1437 13.653
R772 VDD.n1437 VDD.n1436 13.653
R773 VDD.n1433 VDD.n1432 13.653
R774 VDD.n1432 VDD.n1431 13.653
R775 VDD.n1428 VDD.n1427 13.653
R776 VDD.n1427 VDD.n1426 13.653
R777 VDD.n1402 VDD.n1401 13.653
R778 VDD.n1401 VDD.n1400 13.653
R779 VDD.n1398 VDD.n1397 13.653
R780 VDD.n1397 VDD.n1396 13.653
R781 VDD.n1394 VDD.n1393 13.653
R782 VDD.n1393 VDD.n1392 13.653
R783 VDD.n1390 VDD.n1389 13.653
R784 VDD.n1389 VDD.n1388 13.653
R785 VDD.n1385 VDD.n1382 13.653
R786 VDD.n1382 VDD.n1381 13.653
R787 VDD.n1378 VDD.n1377 13.653
R788 VDD.n1377 VDD.n1376 13.653
R789 VDD.n1373 VDD.n1372 13.653
R790 VDD.n1372 VDD.n1371 13.653
R791 VDD.n1368 VDD.n1367 13.653
R792 VDD.n1367 VDD.n1366 13.653
R793 VDD.n1361 VDD.n1360 13.653
R794 VDD.n1360 VDD.n1359 13.653
R795 VDD.n1356 VDD.n1355 13.653
R796 VDD.n1355 VDD.n1354 13.653
R797 VDD.n1351 VDD.n1350 13.653
R798 VDD.n1350 VDD.n1349 13.653
R799 VDD.n1347 VDD.n1346 13.653
R800 VDD.n1346 VDD.n1345 13.653
R801 VDD.n1321 VDD.n1320 13.653
R802 VDD.n1320 VDD.n1319 13.653
R803 VDD.n1317 VDD.n1316 13.653
R804 VDD.n1316 VDD.n1315 13.653
R805 VDD.n1313 VDD.n1312 13.653
R806 VDD.n1312 VDD.n1311 13.653
R807 VDD.n1309 VDD.n1308 13.653
R808 VDD.n1308 VDD.n1307 13.653
R809 VDD.n1304 VDD.n1301 13.653
R810 VDD.n1301 VDD.n1300 13.653
R811 VDD.n1297 VDD.n1296 13.653
R812 VDD.n1296 VDD.n1295 13.653
R813 VDD.n1292 VDD.n1291 13.653
R814 VDD.n1291 VDD.n1290 13.653
R815 VDD.n1287 VDD.n1286 13.653
R816 VDD.n1286 VDD.n1285 13.653
R817 VDD.n1280 VDD.n1279 13.653
R818 VDD.n1279 VDD.n1278 13.653
R819 VDD.n1275 VDD.n1274 13.653
R820 VDD.n1274 VDD.n1273 13.653
R821 VDD.n1270 VDD.n1269 13.653
R822 VDD.n1269 VDD.n1268 13.653
R823 VDD.n1266 VDD.n1265 13.653
R824 VDD.n1265 VDD.n1264 13.653
R825 VDD.n1240 VDD.n1239 13.653
R826 VDD.n1239 VDD.n1238 13.653
R827 VDD.n1236 VDD.n1235 13.653
R828 VDD.n1235 VDD.n1234 13.653
R829 VDD.n1231 VDD.n1230 13.653
R830 VDD.n1230 VDD.n1229 13.653
R831 VDD.n1226 VDD.n1225 13.653
R832 VDD.n1225 VDD.n1224 13.653
R833 VDD.n1220 VDD.n1219 13.653
R834 VDD.n1219 VDD.n1218 13.653
R835 VDD.n1215 VDD.n1214 13.653
R836 VDD.n1214 VDD.n1213 13.653
R837 VDD.n1210 VDD.n1209 13.653
R838 VDD.n1209 VDD.n1208 13.653
R839 VDD.n1205 VDD.n1204 13.653
R840 VDD.n1204 VDD.n1203 13.653
R841 VDD.n1179 VDD.n1178 13.653
R842 VDD.n1178 VDD.n1177 13.653
R843 VDD.n1175 VDD.n1174 13.653
R844 VDD.n1174 VDD.n1173 13.653
R845 VDD.n1171 VDD.n1170 13.653
R846 VDD.n1170 VDD.n1169 13.653
R847 VDD.n1167 VDD.n1166 13.653
R848 VDD.n1166 VDD.n1165 13.653
R849 VDD.n1162 VDD.n1159 13.653
R850 VDD.n1159 VDD.n1158 13.653
R851 VDD.n1155 VDD.n1154 13.653
R852 VDD.n1154 VDD.n1153 13.653
R853 VDD.n1150 VDD.n1149 13.653
R854 VDD.n1149 VDD.n1148 13.653
R855 VDD.n1145 VDD.n1144 13.653
R856 VDD.n1144 VDD.n1143 13.653
R857 VDD.n1138 VDD.n1137 13.653
R858 VDD.n1137 VDD.n1136 13.653
R859 VDD.n1133 VDD.n1132 13.653
R860 VDD.n1132 VDD.n1131 13.653
R861 VDD.n1128 VDD.n1127 13.653
R862 VDD.n1127 VDD.n1126 13.653
R863 VDD.n1124 VDD.n1123 13.653
R864 VDD.n1123 VDD.n1122 13.653
R865 VDD.n1098 VDD.n1097 13.653
R866 VDD.n1097 VDD.n1096 13.653
R867 VDD.n1094 VDD.n1093 13.653
R868 VDD.n1093 VDD.n1092 13.653
R869 VDD.n1089 VDD.n1088 13.653
R870 VDD.n1088 VDD.n1087 13.653
R871 VDD.n1084 VDD.n1083 13.653
R872 VDD.n1083 VDD.n1082 13.653
R873 VDD.n1078 VDD.n1077 13.653
R874 VDD.n1077 VDD.n1076 13.653
R875 VDD.n1073 VDD.n1072 13.653
R876 VDD.n1072 VDD.n1071 13.653
R877 VDD.n1068 VDD.n1067 13.653
R878 VDD.n1067 VDD.n1066 13.653
R879 VDD.n1063 VDD.n1062 13.653
R880 VDD.n1062 VDD.n1061 13.653
R881 VDD.n1037 VDD.n1036 13.653
R882 VDD.n1036 VDD.n1035 13.653
R883 VDD.n1033 VDD.n1032 13.653
R884 VDD.n1032 VDD.n1031 13.653
R885 VDD.n1028 VDD.n1027 13.653
R886 VDD.n1027 VDD.n1026 13.653
R887 VDD.n1023 VDD.n1022 13.653
R888 VDD.n1022 VDD.n1021 13.653
R889 VDD.n1017 VDD.n1016 13.653
R890 VDD.n1016 VDD.n1015 13.653
R891 VDD.n1012 VDD.n1011 13.653
R892 VDD.n1011 VDD.n1010 13.653
R893 VDD.n1007 VDD.n1006 13.653
R894 VDD.n1006 VDD.n1005 13.653
R895 VDD.n1002 VDD.n1001 13.653
R896 VDD.n1001 VDD.n1000 13.653
R897 VDD.n976 VDD.n975 13.653
R898 VDD.n975 VDD.n974 13.653
R899 VDD.n972 VDD.n971 13.653
R900 VDD.n971 VDD.n970 13.653
R901 VDD.n968 VDD.n967 13.653
R902 VDD.n967 VDD.n966 13.653
R903 VDD.n964 VDD.n963 13.653
R904 VDD.n963 VDD.n962 13.653
R905 VDD.n959 VDD.n956 13.653
R906 VDD.n956 VDD.n955 13.653
R907 VDD.n952 VDD.n951 13.653
R908 VDD.n951 VDD.n950 13.653
R909 VDD.n947 VDD.n946 13.653
R910 VDD.n946 VDD.n945 13.653
R911 VDD.n942 VDD.n941 13.653
R912 VDD.n941 VDD.n940 13.653
R913 VDD.n935 VDD.n934 13.653
R914 VDD.n934 VDD.n933 13.653
R915 VDD.n930 VDD.n929 13.653
R916 VDD.n929 VDD.n928 13.653
R917 VDD.n925 VDD.n924 13.653
R918 VDD.n924 VDD.n923 13.653
R919 VDD.n921 VDD.n920 13.653
R920 VDD.n920 VDD.n919 13.653
R921 VDD.n895 VDD.n894 13.653
R922 VDD.n894 VDD.n893 13.653
R923 VDD.n891 VDD.n890 13.653
R924 VDD.n890 VDD.n889 13.653
R925 VDD.n887 VDD.n886 13.653
R926 VDD.n886 VDD.n885 13.653
R927 VDD.n883 VDD.n882 13.653
R928 VDD.n882 VDD.n881 13.653
R929 VDD.n878 VDD.n875 13.653
R930 VDD.n875 VDD.n874 13.653
R931 VDD.n871 VDD.n870 13.653
R932 VDD.n870 VDD.n869 13.653
R933 VDD.n866 VDD.n865 13.653
R934 VDD.n865 VDD.n864 13.653
R935 VDD.n861 VDD.n860 13.653
R936 VDD.n860 VDD.n859 13.653
R937 VDD.n854 VDD.n853 13.653
R938 VDD.n853 VDD.n852 13.653
R939 VDD.n849 VDD.n848 13.653
R940 VDD.n848 VDD.n847 13.653
R941 VDD.n844 VDD.n843 13.653
R942 VDD.n843 VDD.n842 13.653
R943 VDD.n840 VDD.n839 13.653
R944 VDD.n839 VDD.n838 13.653
R945 VDD.n813 VDD.n812 13.653
R946 VDD.n812 VDD.n811 13.653
R947 VDD.n809 VDD.n808 13.653
R948 VDD.n808 VDD.n807 13.653
R949 VDD.n804 VDD.n803 13.653
R950 VDD.n803 VDD.n802 13.653
R951 VDD.n799 VDD.n798 13.653
R952 VDD.n798 VDD.n797 13.653
R953 VDD.n793 VDD.n792 13.653
R954 VDD.n792 VDD.n791 13.653
R955 VDD.n788 VDD.n787 13.653
R956 VDD.n787 VDD.n786 13.653
R957 VDD.n783 VDD.n782 13.653
R958 VDD.n782 VDD.n781 13.653
R959 VDD.n778 VDD.n777 13.653
R960 VDD.n777 VDD.n776 13.653
R961 VDD.n4 VDD.n2 12.915
R962 VDD.n4 VDD.n3 12.66
R963 VDD.n10 VDD.n9 12.343
R964 VDD.n12 VDD.n11 12.343
R965 VDD.n10 VDD.n7 12.343
R966 VDD.n261 VDD.n260 9.152
R967 VDD.n464 VDD.n463 9.152
R968 VDD.n545 VDD.n544 9.152
R969 VDD.n687 VDD.n686 9.152
R970 VDD.n1376 VDD.n1375 9.152
R971 VDD.n1295 VDD.n1294 9.152
R972 VDD.n1153 VDD.n1152 9.152
R973 VDD.n950 VDD.n949 9.152
R974 VDD.n869 VDD.n868 9.152
R975 VDD.n193 VDD.n190 8.658
R976 VDD.n335 VDD.n332 8.658
R977 VDD.n396 VDD.n393 8.658
R978 VDD.n619 VDD.n616 8.658
R979 VDD.n1510 VDD.n1507 8.658
R980 VDD.n1449 VDD.n1446 8.658
R981 VDD.n1226 VDD.n1223 8.658
R982 VDD.n1084 VDD.n1081 8.658
R983 VDD.n1023 VDD.n1020 8.658
R984 VDD.n799 VDD.n796 8.658
R985 VDD.n917 VDD.n916 7.674
R986 VDD.n998 VDD.n997 7.674
R987 VDD.n1059 VDD.n1058 7.674
R988 VDD.n1120 VDD.n1119 7.674
R989 VDD.n1201 VDD.n1200 7.674
R990 VDD.n1262 VDD.n1261 7.674
R991 VDD.n1343 VDD.n1342 7.674
R992 VDD.n1424 VDD.n1423 7.674
R993 VDD.n1485 VDD.n1484 7.674
R994 VDD.n741 VDD.n740 7.674
R995 VDD.n660 VDD.n659 7.674
R996 VDD.n599 VDD.n598 7.674
R997 VDD.n518 VDD.n517 7.674
R998 VDD.n437 VDD.n436 7.674
R999 VDD.n376 VDD.n375 7.674
R1000 VDD.n315 VDD.n314 7.674
R1001 VDD.n234 VDD.n233 7.674
R1002 VDD.n173 VDD.n172 7.674
R1003 VDD.n119 VDD.n118 7.674
R1004 VDD.n65 VDD.n64 7.674
R1005 VDD.n836 VDD.n835 7.674
R1006 VDD.n59 VDD.n58 7.5
R1007 VDD.n53 VDD.n52 7.5
R1008 VDD.n55 VDD.n54 7.5
R1009 VDD.n50 VDD.n49 7.5
R1010 VDD.n64 VDD.n63 7.5
R1011 VDD.n113 VDD.n112 7.5
R1012 VDD.n107 VDD.n106 7.5
R1013 VDD.n109 VDD.n108 7.5
R1014 VDD.n115 VDD.n105 7.5
R1015 VDD.n115 VDD.n103 7.5
R1016 VDD.n118 VDD.n117 7.5
R1017 VDD.n167 VDD.n166 7.5
R1018 VDD.n161 VDD.n160 7.5
R1019 VDD.n163 VDD.n162 7.5
R1020 VDD.n169 VDD.n159 7.5
R1021 VDD.n169 VDD.n157 7.5
R1022 VDD.n172 VDD.n171 7.5
R1023 VDD.n228 VDD.n227 7.5
R1024 VDD.n222 VDD.n221 7.5
R1025 VDD.n224 VDD.n223 7.5
R1026 VDD.n230 VDD.n220 7.5
R1027 VDD.n230 VDD.n218 7.5
R1028 VDD.n233 VDD.n232 7.5
R1029 VDD.n309 VDD.n308 7.5
R1030 VDD.n303 VDD.n302 7.5
R1031 VDD.n305 VDD.n304 7.5
R1032 VDD.n311 VDD.n301 7.5
R1033 VDD.n311 VDD.n299 7.5
R1034 VDD.n314 VDD.n313 7.5
R1035 VDD.n370 VDD.n369 7.5
R1036 VDD.n364 VDD.n363 7.5
R1037 VDD.n366 VDD.n365 7.5
R1038 VDD.n372 VDD.n362 7.5
R1039 VDD.n372 VDD.n360 7.5
R1040 VDD.n375 VDD.n374 7.5
R1041 VDD.n431 VDD.n430 7.5
R1042 VDD.n425 VDD.n424 7.5
R1043 VDD.n427 VDD.n426 7.5
R1044 VDD.n433 VDD.n423 7.5
R1045 VDD.n433 VDD.n421 7.5
R1046 VDD.n436 VDD.n435 7.5
R1047 VDD.n512 VDD.n511 7.5
R1048 VDD.n506 VDD.n505 7.5
R1049 VDD.n508 VDD.n507 7.5
R1050 VDD.n514 VDD.n504 7.5
R1051 VDD.n514 VDD.n502 7.5
R1052 VDD.n517 VDD.n516 7.5
R1053 VDD.n593 VDD.n592 7.5
R1054 VDD.n587 VDD.n586 7.5
R1055 VDD.n589 VDD.n588 7.5
R1056 VDD.n595 VDD.n585 7.5
R1057 VDD.n595 VDD.n583 7.5
R1058 VDD.n598 VDD.n597 7.5
R1059 VDD.n654 VDD.n653 7.5
R1060 VDD.n648 VDD.n647 7.5
R1061 VDD.n650 VDD.n649 7.5
R1062 VDD.n656 VDD.n646 7.5
R1063 VDD.n656 VDD.n644 7.5
R1064 VDD.n659 VDD.n658 7.5
R1065 VDD.n735 VDD.n734 7.5
R1066 VDD.n729 VDD.n728 7.5
R1067 VDD.n731 VDD.n730 7.5
R1068 VDD.n737 VDD.n727 7.5
R1069 VDD.n737 VDD.n725 7.5
R1070 VDD.n740 VDD.n739 7.5
R1071 VDD.n1479 VDD.n1478 7.5
R1072 VDD.n1473 VDD.n1472 7.5
R1073 VDD.n1475 VDD.n1474 7.5
R1074 VDD.n1481 VDD.n1471 7.5
R1075 VDD.n1481 VDD.n1469 7.5
R1076 VDD.n1484 VDD.n1483 7.5
R1077 VDD.n1418 VDD.n1417 7.5
R1078 VDD.n1412 VDD.n1411 7.5
R1079 VDD.n1414 VDD.n1413 7.5
R1080 VDD.n1420 VDD.n1410 7.5
R1081 VDD.n1420 VDD.n1408 7.5
R1082 VDD.n1423 VDD.n1422 7.5
R1083 VDD.n1337 VDD.n1336 7.5
R1084 VDD.n1331 VDD.n1330 7.5
R1085 VDD.n1333 VDD.n1332 7.5
R1086 VDD.n1339 VDD.n1329 7.5
R1087 VDD.n1339 VDD.n1327 7.5
R1088 VDD.n1342 VDD.n1341 7.5
R1089 VDD.n1256 VDD.n1255 7.5
R1090 VDD.n1250 VDD.n1249 7.5
R1091 VDD.n1252 VDD.n1251 7.5
R1092 VDD.n1258 VDD.n1248 7.5
R1093 VDD.n1258 VDD.n1246 7.5
R1094 VDD.n1261 VDD.n1260 7.5
R1095 VDD.n1195 VDD.n1194 7.5
R1096 VDD.n1189 VDD.n1188 7.5
R1097 VDD.n1191 VDD.n1190 7.5
R1098 VDD.n1197 VDD.n1187 7.5
R1099 VDD.n1197 VDD.n1185 7.5
R1100 VDD.n1200 VDD.n1199 7.5
R1101 VDD.n1114 VDD.n1113 7.5
R1102 VDD.n1108 VDD.n1107 7.5
R1103 VDD.n1110 VDD.n1109 7.5
R1104 VDD.n1116 VDD.n1106 7.5
R1105 VDD.n1116 VDD.n1104 7.5
R1106 VDD.n1119 VDD.n1118 7.5
R1107 VDD.n1053 VDD.n1052 7.5
R1108 VDD.n1047 VDD.n1046 7.5
R1109 VDD.n1049 VDD.n1048 7.5
R1110 VDD.n1055 VDD.n1045 7.5
R1111 VDD.n1055 VDD.n1043 7.5
R1112 VDD.n1058 VDD.n1057 7.5
R1113 VDD.n992 VDD.n991 7.5
R1114 VDD.n986 VDD.n985 7.5
R1115 VDD.n988 VDD.n987 7.5
R1116 VDD.n994 VDD.n984 7.5
R1117 VDD.n994 VDD.n982 7.5
R1118 VDD.n997 VDD.n996 7.5
R1119 VDD.n911 VDD.n910 7.5
R1120 VDD.n905 VDD.n904 7.5
R1121 VDD.n907 VDD.n906 7.5
R1122 VDD.n913 VDD.n903 7.5
R1123 VDD.n913 VDD.n901 7.5
R1124 VDD.n916 VDD.n915 7.5
R1125 VDD.n820 VDD.n819 7.5
R1126 VDD.n823 VDD.n822 7.5
R1127 VDD.n825 VDD.n824 7.5
R1128 VDD.n828 VDD.n827 7.5
R1129 VDD.n835 VDD.n834 7.5
R1130 VDD.n770 VDD.n769 7.5
R1131 VDD.n764 VDD.n763 7.5
R1132 VDD.n766 VDD.n765 7.5
R1133 VDD.n772 VDD.n762 7.5
R1134 VDD.n772 VDD.n760 7.5
R1135 VDD.n775 VDD.n774 7.5
R1136 VDD.n20 VDD.n16 7.5
R1137 VDD.n2 VDD.n1 7.5
R1138 VDD.n9 VDD.n8 7.5
R1139 VDD.n7 VDD.n6 7.5
R1140 VDD.n19 VDD.n18 7.5
R1141 VDD.n14 VDD.n0 7.5
R1142 VDD.n51 VDD.n48 6.772
R1143 VDD.n62 VDD.n46 6.772
R1144 VDD.n60 VDD.n57 6.772
R1145 VDD.n56 VDD.n53 6.772
R1146 VDD.n116 VDD.n101 6.772
R1147 VDD.n114 VDD.n111 6.772
R1148 VDD.n110 VDD.n107 6.772
R1149 VDD.n170 VDD.n155 6.772
R1150 VDD.n168 VDD.n165 6.772
R1151 VDD.n164 VDD.n161 6.772
R1152 VDD.n231 VDD.n216 6.772
R1153 VDD.n229 VDD.n226 6.772
R1154 VDD.n225 VDD.n222 6.772
R1155 VDD.n312 VDD.n297 6.772
R1156 VDD.n310 VDD.n307 6.772
R1157 VDD.n306 VDD.n303 6.772
R1158 VDD.n373 VDD.n358 6.772
R1159 VDD.n371 VDD.n368 6.772
R1160 VDD.n367 VDD.n364 6.772
R1161 VDD.n434 VDD.n419 6.772
R1162 VDD.n432 VDD.n429 6.772
R1163 VDD.n428 VDD.n425 6.772
R1164 VDD.n515 VDD.n500 6.772
R1165 VDD.n513 VDD.n510 6.772
R1166 VDD.n509 VDD.n506 6.772
R1167 VDD.n596 VDD.n581 6.772
R1168 VDD.n594 VDD.n591 6.772
R1169 VDD.n590 VDD.n587 6.772
R1170 VDD.n657 VDD.n642 6.772
R1171 VDD.n655 VDD.n652 6.772
R1172 VDD.n651 VDD.n648 6.772
R1173 VDD.n738 VDD.n723 6.772
R1174 VDD.n736 VDD.n733 6.772
R1175 VDD.n732 VDD.n729 6.772
R1176 VDD.n1482 VDD.n1467 6.772
R1177 VDD.n1480 VDD.n1477 6.772
R1178 VDD.n1476 VDD.n1473 6.772
R1179 VDD.n1421 VDD.n1406 6.772
R1180 VDD.n1419 VDD.n1416 6.772
R1181 VDD.n1415 VDD.n1412 6.772
R1182 VDD.n1340 VDD.n1325 6.772
R1183 VDD.n1338 VDD.n1335 6.772
R1184 VDD.n1334 VDD.n1331 6.772
R1185 VDD.n1259 VDD.n1244 6.772
R1186 VDD.n1257 VDD.n1254 6.772
R1187 VDD.n1253 VDD.n1250 6.772
R1188 VDD.n1198 VDD.n1183 6.772
R1189 VDD.n1196 VDD.n1193 6.772
R1190 VDD.n1192 VDD.n1189 6.772
R1191 VDD.n1117 VDD.n1102 6.772
R1192 VDD.n1115 VDD.n1112 6.772
R1193 VDD.n1111 VDD.n1108 6.772
R1194 VDD.n1056 VDD.n1041 6.772
R1195 VDD.n1054 VDD.n1051 6.772
R1196 VDD.n1050 VDD.n1047 6.772
R1197 VDD.n995 VDD.n980 6.772
R1198 VDD.n993 VDD.n990 6.772
R1199 VDD.n989 VDD.n986 6.772
R1200 VDD.n914 VDD.n899 6.772
R1201 VDD.n912 VDD.n909 6.772
R1202 VDD.n908 VDD.n905 6.772
R1203 VDD.n773 VDD.n759 6.772
R1204 VDD.n771 VDD.n768 6.772
R1205 VDD.n767 VDD.n764 6.772
R1206 VDD.n51 VDD.n50 6.772
R1207 VDD.n56 VDD.n55 6.772
R1208 VDD.n60 VDD.n59 6.772
R1209 VDD.n63 VDD.n62 6.772
R1210 VDD.n110 VDD.n109 6.772
R1211 VDD.n114 VDD.n113 6.772
R1212 VDD.n117 VDD.n116 6.772
R1213 VDD.n164 VDD.n163 6.772
R1214 VDD.n168 VDD.n167 6.772
R1215 VDD.n171 VDD.n170 6.772
R1216 VDD.n225 VDD.n224 6.772
R1217 VDD.n229 VDD.n228 6.772
R1218 VDD.n232 VDD.n231 6.772
R1219 VDD.n306 VDD.n305 6.772
R1220 VDD.n310 VDD.n309 6.772
R1221 VDD.n313 VDD.n312 6.772
R1222 VDD.n367 VDD.n366 6.772
R1223 VDD.n371 VDD.n370 6.772
R1224 VDD.n374 VDD.n373 6.772
R1225 VDD.n428 VDD.n427 6.772
R1226 VDD.n432 VDD.n431 6.772
R1227 VDD.n435 VDD.n434 6.772
R1228 VDD.n509 VDD.n508 6.772
R1229 VDD.n513 VDD.n512 6.772
R1230 VDD.n516 VDD.n515 6.772
R1231 VDD.n590 VDD.n589 6.772
R1232 VDD.n594 VDD.n593 6.772
R1233 VDD.n597 VDD.n596 6.772
R1234 VDD.n651 VDD.n650 6.772
R1235 VDD.n655 VDD.n654 6.772
R1236 VDD.n658 VDD.n657 6.772
R1237 VDD.n732 VDD.n731 6.772
R1238 VDD.n736 VDD.n735 6.772
R1239 VDD.n739 VDD.n738 6.772
R1240 VDD.n1476 VDD.n1475 6.772
R1241 VDD.n1480 VDD.n1479 6.772
R1242 VDD.n1483 VDD.n1482 6.772
R1243 VDD.n1415 VDD.n1414 6.772
R1244 VDD.n1419 VDD.n1418 6.772
R1245 VDD.n1422 VDD.n1421 6.772
R1246 VDD.n1334 VDD.n1333 6.772
R1247 VDD.n1338 VDD.n1337 6.772
R1248 VDD.n1341 VDD.n1340 6.772
R1249 VDD.n1253 VDD.n1252 6.772
R1250 VDD.n1257 VDD.n1256 6.772
R1251 VDD.n1260 VDD.n1259 6.772
R1252 VDD.n1192 VDD.n1191 6.772
R1253 VDD.n1196 VDD.n1195 6.772
R1254 VDD.n1199 VDD.n1198 6.772
R1255 VDD.n1111 VDD.n1110 6.772
R1256 VDD.n1115 VDD.n1114 6.772
R1257 VDD.n1118 VDD.n1117 6.772
R1258 VDD.n1050 VDD.n1049 6.772
R1259 VDD.n1054 VDD.n1053 6.772
R1260 VDD.n1057 VDD.n1056 6.772
R1261 VDD.n989 VDD.n988 6.772
R1262 VDD.n993 VDD.n992 6.772
R1263 VDD.n996 VDD.n995 6.772
R1264 VDD.n908 VDD.n907 6.772
R1265 VDD.n912 VDD.n911 6.772
R1266 VDD.n915 VDD.n914 6.772
R1267 VDD.n767 VDD.n766 6.772
R1268 VDD.n771 VDD.n770 6.772
R1269 VDD.n774 VDD.n773 6.772
R1270 VDD.n834 VDD.n833 6.772
R1271 VDD.n821 VDD.n818 6.772
R1272 VDD.n826 VDD.n823 6.772
R1273 VDD.n831 VDD.n828 6.772
R1274 VDD.n831 VDD.n830 6.772
R1275 VDD.n826 VDD.n825 6.772
R1276 VDD.n821 VDD.n820 6.772
R1277 VDD.n833 VDD.n817 6.772
R1278 VDD.n275 VDD.n271 6.69
R1279 VDD.n478 VDD.n474 6.69
R1280 VDD.n559 VDD.n555 6.69
R1281 VDD.n701 VDD.n697 6.69
R1282 VDD.n1368 VDD.n1364 6.69
R1283 VDD.n1287 VDD.n1283 6.69
R1284 VDD.n1145 VDD.n1141 6.69
R1285 VDD.n942 VDD.n938 6.69
R1286 VDD.n861 VDD.n857 6.69
R1287 VDD.n16 VDD.n15 6.458
R1288 VDD.n258 VDD.n257 6.296
R1289 VDD.n461 VDD.n460 6.296
R1290 VDD.n542 VDD.n541 6.296
R1291 VDD.n684 VDD.n683 6.296
R1292 VDD.n1385 VDD.n1384 6.296
R1293 VDD.n1304 VDD.n1303 6.296
R1294 VDD.n1162 VDD.n1161 6.296
R1295 VDD.n959 VDD.n958 6.296
R1296 VDD.n878 VDD.n877 6.296
R1297 VDD.n105 VDD.n104 6.202
R1298 VDD.n159 VDD.n158 6.202
R1299 VDD.n220 VDD.n219 6.202
R1300 VDD.n301 VDD.n300 6.202
R1301 VDD.n362 VDD.n361 6.202
R1302 VDD.n423 VDD.n422 6.202
R1303 VDD.n504 VDD.n503 6.202
R1304 VDD.n585 VDD.n584 6.202
R1305 VDD.n646 VDD.n645 6.202
R1306 VDD.n727 VDD.n726 6.202
R1307 VDD.n1471 VDD.n1470 6.202
R1308 VDD.n1410 VDD.n1409 6.202
R1309 VDD.n1329 VDD.n1328 6.202
R1310 VDD.n1248 VDD.n1247 6.202
R1311 VDD.n1187 VDD.n1186 6.202
R1312 VDD.n1106 VDD.n1105 6.202
R1313 VDD.n1045 VDD.n1044 6.202
R1314 VDD.n984 VDD.n983 6.202
R1315 VDD.n903 VDD.n902 6.202
R1316 VDD.n762 VDD.n761 6.202
R1317 VDD.n196 VDD.n195 4.576
R1318 VDD.n338 VDD.n337 4.576
R1319 VDD.n399 VDD.n398 4.576
R1320 VDD.n622 VDD.n621 4.576
R1321 VDD.n1502 VDD.n1501 4.576
R1322 VDD.n1441 VDD.n1440 4.576
R1323 VDD.n1218 VDD.n1217 4.576
R1324 VDD.n1076 VDD.n1075 4.576
R1325 VDD.n1015 VDD.n1014 4.576
R1326 VDD.n791 VDD.n790 4.576
R1327 VDD.n208 VDD.n205 2.754
R1328 VDD.n350 VDD.n347 2.754
R1329 VDD.n411 VDD.n408 2.754
R1330 VDD.n634 VDD.n631 2.754
R1331 VDD.n1494 VDD.n1491 2.754
R1332 VDD.n1433 VDD.n1430 2.754
R1333 VDD.n1210 VDD.n1207 2.754
R1334 VDD.n1068 VDD.n1065 2.754
R1335 VDD.n1007 VDD.n1004 2.754
R1336 VDD.n783 VDD.n780 2.754
R1337 VDD.n182 VDD.n179 2.361
R1338 VDD.n324 VDD.n321 2.361
R1339 VDD.n385 VDD.n382 2.361
R1340 VDD.n608 VDD.n605 2.361
R1341 VDD.n750 VDD.n747 2.361
R1342 VDD.n1459 VDD.n1456 2.361
R1343 VDD.n1236 VDD.n1233 2.361
R1344 VDD.n1094 VDD.n1091 2.361
R1345 VDD.n1033 VDD.n1030 2.361
R1346 VDD.n809 VDD.n806 2.361
R1347 VDD.n28 VDD.n24 1.967
R1348 VDD.n38 VDD.n37 1.967
R1349 VDD.n14 VDD.n5 1.329
R1350 VDD.n14 VDD.n10 1.329
R1351 VDD.n14 VDD.n12 1.329
R1352 VDD.n14 VDD.n13 1.329
R1353 VDD.n15 VDD.n14 0.696
R1354 VDD.n14 VDD.n4 0.696
R1355 VDD.n285 VDD.n282 0.393
R1356 VDD.n488 VDD.n485 0.393
R1357 VDD.n569 VDD.n566 0.393
R1358 VDD.n711 VDD.n708 0.393
R1359 VDD.n1356 VDD.n1353 0.393
R1360 VDD.n1275 VDD.n1272 0.393
R1361 VDD.n1133 VDD.n1130 0.393
R1362 VDD.n930 VDD.n927 0.393
R1363 VDD.n849 VDD.n846 0.393
R1364 VDD.n61 VDD.n60 0.365
R1365 VDD.n61 VDD.n56 0.365
R1366 VDD.n61 VDD.n51 0.365
R1367 VDD.n62 VDD.n61 0.365
R1368 VDD.n115 VDD.n114 0.365
R1369 VDD.n115 VDD.n110 0.365
R1370 VDD.n116 VDD.n115 0.365
R1371 VDD.n169 VDD.n168 0.365
R1372 VDD.n169 VDD.n164 0.365
R1373 VDD.n170 VDD.n169 0.365
R1374 VDD.n230 VDD.n229 0.365
R1375 VDD.n230 VDD.n225 0.365
R1376 VDD.n231 VDD.n230 0.365
R1377 VDD.n311 VDD.n310 0.365
R1378 VDD.n311 VDD.n306 0.365
R1379 VDD.n312 VDD.n311 0.365
R1380 VDD.n372 VDD.n371 0.365
R1381 VDD.n372 VDD.n367 0.365
R1382 VDD.n373 VDD.n372 0.365
R1383 VDD.n433 VDD.n432 0.365
R1384 VDD.n433 VDD.n428 0.365
R1385 VDD.n434 VDD.n433 0.365
R1386 VDD.n514 VDD.n513 0.365
R1387 VDD.n514 VDD.n509 0.365
R1388 VDD.n515 VDD.n514 0.365
R1389 VDD.n595 VDD.n594 0.365
R1390 VDD.n595 VDD.n590 0.365
R1391 VDD.n596 VDD.n595 0.365
R1392 VDD.n656 VDD.n655 0.365
R1393 VDD.n656 VDD.n651 0.365
R1394 VDD.n657 VDD.n656 0.365
R1395 VDD.n737 VDD.n736 0.365
R1396 VDD.n737 VDD.n732 0.365
R1397 VDD.n738 VDD.n737 0.365
R1398 VDD.n1481 VDD.n1480 0.365
R1399 VDD.n1481 VDD.n1476 0.365
R1400 VDD.n1482 VDD.n1481 0.365
R1401 VDD.n1420 VDD.n1419 0.365
R1402 VDD.n1420 VDD.n1415 0.365
R1403 VDD.n1421 VDD.n1420 0.365
R1404 VDD.n1339 VDD.n1338 0.365
R1405 VDD.n1339 VDD.n1334 0.365
R1406 VDD.n1340 VDD.n1339 0.365
R1407 VDD.n1258 VDD.n1257 0.365
R1408 VDD.n1258 VDD.n1253 0.365
R1409 VDD.n1259 VDD.n1258 0.365
R1410 VDD.n1197 VDD.n1196 0.365
R1411 VDD.n1197 VDD.n1192 0.365
R1412 VDD.n1198 VDD.n1197 0.365
R1413 VDD.n1116 VDD.n1115 0.365
R1414 VDD.n1116 VDD.n1111 0.365
R1415 VDD.n1117 VDD.n1116 0.365
R1416 VDD.n1055 VDD.n1054 0.365
R1417 VDD.n1055 VDD.n1050 0.365
R1418 VDD.n1056 VDD.n1055 0.365
R1419 VDD.n994 VDD.n993 0.365
R1420 VDD.n994 VDD.n989 0.365
R1421 VDD.n995 VDD.n994 0.365
R1422 VDD.n913 VDD.n912 0.365
R1423 VDD.n913 VDD.n908 0.365
R1424 VDD.n914 VDD.n913 0.365
R1425 VDD.n772 VDD.n771 0.365
R1426 VDD.n772 VDD.n767 0.365
R1427 VDD.n773 VDD.n772 0.365
R1428 VDD.n832 VDD.n831 0.365
R1429 VDD.n832 VDD.n826 0.365
R1430 VDD.n832 VDD.n821 0.365
R1431 VDD.n833 VDD.n832 0.365
R1432 VDD.n70 VDD.n43 0.29
R1433 VDD.n124 VDD.n98 0.29
R1434 VDD.n178 VDD.n152 0.29
R1435 VDD.n239 VDD.n213 0.29
R1436 VDD.n320 VDD.n294 0.29
R1437 VDD.n381 VDD.n355 0.29
R1438 VDD.n442 VDD.n416 0.29
R1439 VDD.n523 VDD.n497 0.29
R1440 VDD.n604 VDD.n578 0.29
R1441 VDD.n665 VDD.n639 0.29
R1442 VDD.n746 VDD.n720 0.29
R1443 VDD.n1490 VDD.n1464 0.29
R1444 VDD.n1429 VDD.n1403 0.29
R1445 VDD.n1348 VDD.n1322 0.29
R1446 VDD.n1267 VDD.n1241 0.29
R1447 VDD.n1206 VDD.n1180 0.29
R1448 VDD.n1125 VDD.n1099 0.29
R1449 VDD.n1064 VDD.n1038 0.29
R1450 VDD.n1003 VDD.n977 0.29
R1451 VDD.n922 VDD.n896 0.29
R1452 VDD.n841 VDD.n814 0.29
R1453 VDD.n779 VDD 0.207
R1454 VDD.n269 VDD.n264 0.197
R1455 VDD.n472 VDD.n467 0.197
R1456 VDD.n553 VDD.n548 0.197
R1457 VDD.n695 VDD.n690 0.197
R1458 VDD.n1379 VDD.n1374 0.197
R1459 VDD.n1298 VDD.n1293 0.197
R1460 VDD.n1156 VDD.n1151 0.197
R1461 VDD.n953 VDD.n948 0.197
R1462 VDD.n872 VDD.n867 0.197
R1463 VDD.n86 VDD.n82 0.181
R1464 VDD.n140 VDD.n136 0.181
R1465 VDD.n199 VDD.n194 0.181
R1466 VDD.n341 VDD.n336 0.181
R1467 VDD.n402 VDD.n397 0.181
R1468 VDD.n625 VDD.n620 0.181
R1469 VDD.n1511 VDD.n1505 0.181
R1470 VDD.n1450 VDD.n1444 0.181
R1471 VDD.n1227 VDD.n1221 0.181
R1472 VDD.n1085 VDD.n1079 0.181
R1473 VDD.n1024 VDD.n1018 0.181
R1474 VDD.n800 VDD.n794 0.181
R1475 VDD.n33 VDD.n29 0.157
R1476 VDD.n39 VDD.n33 0.157
R1477 VDD.n43 VDD.n39 0.145
R1478 VDD.n74 VDD.n70 0.145
R1479 VDD.n78 VDD.n74 0.145
R1480 VDD.n82 VDD.n78 0.145
R1481 VDD.n90 VDD.n86 0.145
R1482 VDD.n94 VDD.n90 0.145
R1483 VDD.n98 VDD.n94 0.145
R1484 VDD.n128 VDD.n124 0.145
R1485 VDD.n132 VDD.n128 0.145
R1486 VDD.n136 VDD.n132 0.145
R1487 VDD.n144 VDD.n140 0.145
R1488 VDD.n148 VDD.n144 0.145
R1489 VDD.n152 VDD.n148 0.145
R1490 VDD.n183 VDD.n178 0.145
R1491 VDD.n188 VDD.n183 0.145
R1492 VDD.n194 VDD.n188 0.145
R1493 VDD.n204 VDD.n199 0.145
R1494 VDD.n209 VDD.n204 0.145
R1495 VDD.n213 VDD.n209 0.145
R1496 VDD.n243 VDD.n239 0.145
R1497 VDD.n247 VDD.n243 0.145
R1498 VDD.n252 VDD.n247 0.145
R1499 VDD.n259 VDD.n252 0.145
R1500 VDD.n264 VDD.n259 0.145
R1501 VDD.n276 VDD.n269 0.145
R1502 VDD.n281 VDD.n276 0.145
R1503 VDD.n286 VDD.n281 0.145
R1504 VDD.n290 VDD.n286 0.145
R1505 VDD.n294 VDD.n290 0.145
R1506 VDD.n325 VDD.n320 0.145
R1507 VDD.n330 VDD.n325 0.145
R1508 VDD.n336 VDD.n330 0.145
R1509 VDD.n346 VDD.n341 0.145
R1510 VDD.n351 VDD.n346 0.145
R1511 VDD.n355 VDD.n351 0.145
R1512 VDD.n386 VDD.n381 0.145
R1513 VDD.n391 VDD.n386 0.145
R1514 VDD.n397 VDD.n391 0.145
R1515 VDD.n407 VDD.n402 0.145
R1516 VDD.n412 VDD.n407 0.145
R1517 VDD.n416 VDD.n412 0.145
R1518 VDD.n446 VDD.n442 0.145
R1519 VDD.n450 VDD.n446 0.145
R1520 VDD.n455 VDD.n450 0.145
R1521 VDD.n462 VDD.n455 0.145
R1522 VDD.n467 VDD.n462 0.145
R1523 VDD.n479 VDD.n472 0.145
R1524 VDD.n484 VDD.n479 0.145
R1525 VDD.n489 VDD.n484 0.145
R1526 VDD.n493 VDD.n489 0.145
R1527 VDD.n497 VDD.n493 0.145
R1528 VDD.n527 VDD.n523 0.145
R1529 VDD.n531 VDD.n527 0.145
R1530 VDD.n536 VDD.n531 0.145
R1531 VDD.n543 VDD.n536 0.145
R1532 VDD.n548 VDD.n543 0.145
R1533 VDD.n560 VDD.n553 0.145
R1534 VDD.n565 VDD.n560 0.145
R1535 VDD.n570 VDD.n565 0.145
R1536 VDD.n574 VDD.n570 0.145
R1537 VDD.n578 VDD.n574 0.145
R1538 VDD.n609 VDD.n604 0.145
R1539 VDD.n614 VDD.n609 0.145
R1540 VDD.n620 VDD.n614 0.145
R1541 VDD.n630 VDD.n625 0.145
R1542 VDD.n635 VDD.n630 0.145
R1543 VDD.n639 VDD.n635 0.145
R1544 VDD.n669 VDD.n665 0.145
R1545 VDD.n673 VDD.n669 0.145
R1546 VDD.n678 VDD.n673 0.145
R1547 VDD.n685 VDD.n678 0.145
R1548 VDD.n690 VDD.n685 0.145
R1549 VDD.n702 VDD.n695 0.145
R1550 VDD.n707 VDD.n702 0.145
R1551 VDD.n712 VDD.n707 0.145
R1552 VDD.n716 VDD.n712 0.145
R1553 VDD.n720 VDD.n716 0.145
R1554 VDD.n751 VDD.n746 0.145
R1555 VDD.n756 VDD.n751 0.145
R1556 VDD.n1505 VDD.n1500 0.145
R1557 VDD.n1500 VDD.n1495 0.145
R1558 VDD.n1495 VDD.n1490 0.145
R1559 VDD.n1464 VDD.n1460 0.145
R1560 VDD.n1460 VDD.n1455 0.145
R1561 VDD.n1455 VDD.n1450 0.145
R1562 VDD.n1444 VDD.n1439 0.145
R1563 VDD.n1439 VDD.n1434 0.145
R1564 VDD.n1434 VDD.n1429 0.145
R1565 VDD.n1403 VDD.n1399 0.145
R1566 VDD.n1399 VDD.n1395 0.145
R1567 VDD.n1395 VDD.n1391 0.145
R1568 VDD.n1391 VDD.n1386 0.145
R1569 VDD.n1386 VDD.n1379 0.145
R1570 VDD.n1374 VDD.n1369 0.145
R1571 VDD.n1369 VDD.n1362 0.145
R1572 VDD.n1362 VDD.n1357 0.145
R1573 VDD.n1357 VDD.n1352 0.145
R1574 VDD.n1352 VDD.n1348 0.145
R1575 VDD.n1322 VDD.n1318 0.145
R1576 VDD.n1318 VDD.n1314 0.145
R1577 VDD.n1314 VDD.n1310 0.145
R1578 VDD.n1310 VDD.n1305 0.145
R1579 VDD.n1305 VDD.n1298 0.145
R1580 VDD.n1293 VDD.n1288 0.145
R1581 VDD.n1288 VDD.n1281 0.145
R1582 VDD.n1281 VDD.n1276 0.145
R1583 VDD.n1276 VDD.n1271 0.145
R1584 VDD.n1271 VDD.n1267 0.145
R1585 VDD.n1241 VDD.n1237 0.145
R1586 VDD.n1237 VDD.n1232 0.145
R1587 VDD.n1232 VDD.n1227 0.145
R1588 VDD.n1221 VDD.n1216 0.145
R1589 VDD.n1216 VDD.n1211 0.145
R1590 VDD.n1211 VDD.n1206 0.145
R1591 VDD.n1180 VDD.n1176 0.145
R1592 VDD.n1176 VDD.n1172 0.145
R1593 VDD.n1172 VDD.n1168 0.145
R1594 VDD.n1168 VDD.n1163 0.145
R1595 VDD.n1163 VDD.n1156 0.145
R1596 VDD.n1151 VDD.n1146 0.145
R1597 VDD.n1146 VDD.n1139 0.145
R1598 VDD.n1139 VDD.n1134 0.145
R1599 VDD.n1134 VDD.n1129 0.145
R1600 VDD.n1129 VDD.n1125 0.145
R1601 VDD.n1099 VDD.n1095 0.145
R1602 VDD.n1095 VDD.n1090 0.145
R1603 VDD.n1090 VDD.n1085 0.145
R1604 VDD.n1079 VDD.n1074 0.145
R1605 VDD.n1074 VDD.n1069 0.145
R1606 VDD.n1069 VDD.n1064 0.145
R1607 VDD.n1038 VDD.n1034 0.145
R1608 VDD.n1034 VDD.n1029 0.145
R1609 VDD.n1029 VDD.n1024 0.145
R1610 VDD.n1018 VDD.n1013 0.145
R1611 VDD.n1013 VDD.n1008 0.145
R1612 VDD.n1008 VDD.n1003 0.145
R1613 VDD.n977 VDD.n973 0.145
R1614 VDD.n973 VDD.n969 0.145
R1615 VDD.n969 VDD.n965 0.145
R1616 VDD.n965 VDD.n960 0.145
R1617 VDD.n960 VDD.n953 0.145
R1618 VDD.n948 VDD.n943 0.145
R1619 VDD.n943 VDD.n936 0.145
R1620 VDD.n936 VDD.n931 0.145
R1621 VDD.n931 VDD.n926 0.145
R1622 VDD.n926 VDD.n922 0.145
R1623 VDD.n896 VDD.n892 0.145
R1624 VDD.n892 VDD.n888 0.145
R1625 VDD.n888 VDD.n884 0.145
R1626 VDD.n884 VDD.n879 0.145
R1627 VDD.n879 VDD.n872 0.145
R1628 VDD.n867 VDD.n862 0.145
R1629 VDD.n862 VDD.n855 0.145
R1630 VDD.n855 VDD.n850 0.145
R1631 VDD.n850 VDD.n845 0.145
R1632 VDD.n845 VDD.n841 0.145
R1633 VDD.n814 VDD.n810 0.145
R1634 VDD.n810 VDD.n805 0.145
R1635 VDD.n805 VDD.n800 0.145
R1636 VDD.n794 VDD.n789 0.145
R1637 VDD.n789 VDD.n784 0.145
R1638 VDD.n784 VDD.n779 0.145
R1639 VDD VDD.n756 0.086
R1640 VDD VDD.n1511 0.058
R1641 a_8357_1050.n0 a_8357_1050.t5 512.525
R1642 a_8357_1050.n0 a_8357_1050.t7 371.139
R1643 a_8357_1050.n1 a_8357_1050.t6 340.774
R1644 a_8357_1050.n6 a_8357_1050.n5 263.698
R1645 a_8357_1050.n6 a_8357_1050.n1 153.315
R1646 a_8357_1050.n1 a_8357_1050.n0 109.607
R1647 a_8357_1050.n8 a_8357_1050.n6 99.394
R1648 a_8357_1050.n8 a_8357_1050.n7 76.002
R1649 a_8357_1050.n5 a_8357_1050.n4 30
R1650 a_8357_1050.n3 a_8357_1050.n2 24.383
R1651 a_8357_1050.n5 a_8357_1050.n3 23.684
R1652 a_8357_1050.n7 a_8357_1050.t0 14.282
R1653 a_8357_1050.n7 a_8357_1050.t4 14.282
R1654 a_8357_1050.n9 a_8357_1050.t1 14.282
R1655 a_8357_1050.t2 a_8357_1050.n9 14.282
R1656 a_8357_1050.n9 a_8357_1050.n8 12.848
R1657 SN.n14 SN.t3 479.223
R1658 SN.n11 SN.t12 479.223
R1659 SN.n8 SN.t13 479.223
R1660 SN.n5 SN.t2 479.223
R1661 SN.n2 SN.t9 479.223
R1662 SN.n0 SN.t8 479.223
R1663 SN.n14 SN.t14 375.52
R1664 SN.n11 SN.t4 375.52
R1665 SN.n8 SN.t15 375.52
R1666 SN.n5 SN.t7 375.52
R1667 SN.n2 SN.t17 375.52
R1668 SN.n0 SN.t16 375.52
R1669 SN.n15 SN.n14 175.429
R1670 SN.n12 SN.n11 175.429
R1671 SN.n9 SN.n8 175.429
R1672 SN.n6 SN.n5 175.429
R1673 SN.n3 SN.n2 175.429
R1674 SN.n1 SN.n0 175.429
R1675 SN.n15 SN.t11 162.048
R1676 SN.n12 SN.t1 162.048
R1677 SN.n9 SN.t0 162.048
R1678 SN.n6 SN.t6 162.048
R1679 SN.n3 SN.t5 162.048
R1680 SN.n1 SN.t10 162.048
R1681 SN.n4 SN.n1 84.388
R1682 SN.n4 SN.n3 76
R1683 SN.n7 SN.n6 76
R1684 SN.n10 SN.n9 76
R1685 SN.n13 SN.n12 76
R1686 SN.n16 SN.n15 76
R1687 SN.n7 SN.n4 9.476
R1688 SN.n13 SN.n10 9.476
R1689 SN.n10 SN.n7 8.388
R1690 SN.n16 SN.n13 8.388
R1691 SN.n16 SN 0.046
R1692 a_6603_103.t0 a_6603_103.n3 117.777
R1693 a_6603_103.n6 a_6603_103.n5 45.444
R1694 a_6603_103.t0 a_6603_103.n6 21.213
R1695 a_6603_103.t0 a_6603_103.n4 11.595
R1696 a_6603_103.n2 a_6603_103.n0 8.543
R1697 a_6603_103.t0 a_6603_103.n2 3.034
R1698 a_6603_103.n2 a_6603_103.n1 0.443
R1699 a_6884_210.n8 a_6884_210.n6 96.467
R1700 a_6884_210.n3 a_6884_210.n1 44.628
R1701 a_6884_210.t0 a_6884_210.n8 32.417
R1702 a_6884_210.n3 a_6884_210.n2 23.284
R1703 a_6884_210.n6 a_6884_210.n5 22.349
R1704 a_6884_210.t0 a_6884_210.n10 20.241
R1705 a_6884_210.n10 a_6884_210.n9 13.494
R1706 a_6884_210.n6 a_6884_210.n4 8.443
R1707 a_6884_210.t0 a_6884_210.n0 8.137
R1708 a_6884_210.t0 a_6884_210.n3 5.727
R1709 a_6884_210.n8 a_6884_210.n7 1.435
R1710 a_3473_1050.n3 a_3473_1050.t6 512.525
R1711 a_3473_1050.n3 a_3473_1050.t5 371.139
R1712 a_3473_1050.n4 a_3473_1050.t7 340.774
R1713 a_3473_1050.n7 a_3473_1050.n5 270.22
R1714 a_3473_1050.n5 a_3473_1050.n4 153.315
R1715 a_3473_1050.n4 a_3473_1050.n3 109.607
R1716 a_3473_1050.n5 a_3473_1050.n2 99.394
R1717 a_3473_1050.n2 a_3473_1050.n1 76.002
R1718 a_3473_1050.n7 a_3473_1050.n6 15.218
R1719 a_3473_1050.n0 a_3473_1050.t3 14.282
R1720 a_3473_1050.n0 a_3473_1050.t4 14.282
R1721 a_3473_1050.n1 a_3473_1050.t2 14.282
R1722 a_3473_1050.n1 a_3473_1050.t1 14.282
R1723 a_3473_1050.n2 a_3473_1050.n0 12.85
R1724 a_3473_1050.n8 a_3473_1050.n7 12.014
R1725 a_3599_411.n3 a_3599_411.t7 512.525
R1726 a_3599_411.n2 a_3599_411.t11 512.525
R1727 a_3599_411.n7 a_3599_411.t15 472.359
R1728 a_3599_411.n7 a_3599_411.t9 384.527
R1729 a_3599_411.n3 a_3599_411.t13 371.139
R1730 a_3599_411.n2 a_3599_411.t8 371.139
R1731 a_3599_411.n4 a_3599_411.n3 265.439
R1732 a_3599_411.n8 a_3599_411.t12 214.619
R1733 a_3599_411.n15 a_3599_411.n14 197.352
R1734 a_3599_411.n14 a_3599_411.n13 186.551
R1735 a_3599_411.n6 a_3599_411.n2 185.78
R1736 a_3599_411.n4 a_3599_411.t14 176.995
R1737 a_3599_411.n5 a_3599_411.t10 170.569
R1738 a_3599_411.n5 a_3599_411.n4 153.043
R1739 a_3599_411.n8 a_3599_411.n7 136.613
R1740 a_3599_411.n9 a_3599_411.n6 116.763
R1741 a_3599_411.n9 a_3599_411.n8 80.035
R1742 a_3599_411.n6 a_3599_411.n5 79.658
R1743 a_3599_411.n17 a_3599_411.n16 79.231
R1744 a_3599_411.n14 a_3599_411.n9 76
R1745 a_3599_411.n16 a_3599_411.n15 63.152
R1746 a_3599_411.n13 a_3599_411.n12 30
R1747 a_3599_411.n11 a_3599_411.n10 24.383
R1748 a_3599_411.n13 a_3599_411.n11 23.684
R1749 a_3599_411.n15 a_3599_411.n1 16.08
R1750 a_3599_411.n16 a_3599_411.n0 16.08
R1751 a_3599_411.n1 a_3599_411.t1 14.282
R1752 a_3599_411.n1 a_3599_411.t4 14.282
R1753 a_3599_411.n0 a_3599_411.t5 14.282
R1754 a_3599_411.n0 a_3599_411.t6 14.282
R1755 a_3599_411.n17 a_3599_411.t2 14.282
R1756 a_3599_411.t3 a_3599_411.n17 14.282
R1757 CLK.n15 CLK.t17 472.359
R1758 CLK.n6 CLK.t0 472.359
R1759 CLK.n0 CLK.t4 472.359
R1760 CLK.n20 CLK.t9 459.505
R1761 CLK.n11 CLK.t2 459.505
R1762 CLK.n2 CLK.t15 459.505
R1763 CLK.n20 CLK.t14 384.527
R1764 CLK.n15 CLK.t1 384.527
R1765 CLK.n11 CLK.t5 384.527
R1766 CLK.n6 CLK.t8 384.527
R1767 CLK.n2 CLK.t7 384.527
R1768 CLK.n0 CLK.t13 384.527
R1769 CLK.n21 CLK.t11 322.152
R1770 CLK.n12 CLK.t12 322.151
R1771 CLK.n3 CLK.t3 322.151
R1772 CLK.n1 CLK.t10 321.724
R1773 CLK.n17 CLK.t16 319.581
R1774 CLK.n8 CLK.t6 319.581
R1775 CLK.n9 CLK.n8 75.621
R1776 CLK.n18 CLK.n17 75.621
R1777 CLK.n22 CLK.n21 49.342
R1778 CLK.n4 CLK.n3 49.342
R1779 CLK.n13 CLK.n12 49.342
R1780 CLK.n4 CLK.n1 43.573
R1781 CLK.n21 CLK.n20 27.599
R1782 CLK.n3 CLK.n2 27.599
R1783 CLK.n12 CLK.n11 27.599
R1784 CLK.n1 CLK.n0 23.329
R1785 CLK.n16 CLK.n15 21.176
R1786 CLK.n7 CLK.n6 21.176
R1787 CLK.n5 CLK.n4 11.101
R1788 CLK.n14 CLK.n13 11.101
R1789 CLK.n13 CLK.n10 6.718
R1790 CLK.n22 CLK.n19 6.718
R1791 CLK.n17 CLK.n16 4.419
R1792 CLK.n8 CLK.n7 4.419
R1793 CLK.n22 CLK 0.046
R1794 CLK.n10 CLK.n9 0.038
R1795 CLK.n19 CLK.n18 0.038
R1796 CLK.n9 CLK.n5 0.008
R1797 CLK.n18 CLK.n14 0.008
R1798 a_6149_989.n2 a_6149_989.t5 454.685
R1799 a_6149_989.n4 a_6149_989.t8 454.685
R1800 a_6149_989.n0 a_6149_989.t10 454.685
R1801 a_6149_989.n2 a_6149_989.t11 428.979
R1802 a_6149_989.n4 a_6149_989.t13 428.979
R1803 a_6149_989.n0 a_6149_989.t9 428.979
R1804 a_6149_989.n3 a_6149_989.t7 264.512
R1805 a_6149_989.n5 a_6149_989.t6 264.512
R1806 a_6149_989.n1 a_6149_989.t12 264.512
R1807 a_6149_989.n12 a_6149_989.n11 237.145
R1808 a_6149_989.n14 a_6149_989.n12 125.947
R1809 a_6149_989.n7 a_6149_989.n1 81.396
R1810 a_6149_989.n6 a_6149_989.n5 79.491
R1811 a_6149_989.n14 a_6149_989.n13 76.002
R1812 a_6149_989.n6 a_6149_989.n3 76
R1813 a_6149_989.n12 a_6149_989.n7 76
R1814 a_6149_989.n3 a_6149_989.n2 71.894
R1815 a_6149_989.n5 a_6149_989.n4 71.894
R1816 a_6149_989.n1 a_6149_989.n0 71.894
R1817 a_6149_989.n11 a_6149_989.n10 30
R1818 a_6149_989.n9 a_6149_989.n8 24.383
R1819 a_6149_989.n11 a_6149_989.n9 23.684
R1820 a_6149_989.n13 a_6149_989.t3 14.282
R1821 a_6149_989.n13 a_6149_989.t4 14.282
R1822 a_6149_989.t1 a_6149_989.n15 14.282
R1823 a_6149_989.n15 a_6149_989.t0 14.282
R1824 a_6149_989.n15 a_6149_989.n14 12.848
R1825 a_6149_989.n7 a_6149_989.n6 2.947
R1826 a_14869_1051.n4 a_14869_1051.n3 195.987
R1827 a_14869_1051.n2 a_14869_1051.t0 89.553
R1828 a_14869_1051.n5 a_14869_1051.n4 75.27
R1829 a_14869_1051.n3 a_14869_1051.n2 75.214
R1830 a_14869_1051.n4 a_14869_1051.n0 36.519
R1831 a_14869_1051.n3 a_14869_1051.t5 14.338
R1832 a_14869_1051.n0 a_14869_1051.t7 14.282
R1833 a_14869_1051.n0 a_14869_1051.t6 14.282
R1834 a_14869_1051.n1 a_14869_1051.t1 14.282
R1835 a_14869_1051.n1 a_14869_1051.t4 14.282
R1836 a_14869_1051.t3 a_14869_1051.n5 14.282
R1837 a_14869_1051.n5 a_14869_1051.t2 14.282
R1838 a_14869_1051.n2 a_14869_1051.n1 12.119
R1839 a_13367_411.n1 a_13367_411.t8 475.572
R1840 a_13367_411.n6 a_13367_411.t15 472.359
R1841 a_13367_411.n3 a_13367_411.t11 469.145
R1842 a_13367_411.n6 a_13367_411.t10 384.527
R1843 a_13367_411.n3 a_13367_411.t14 384.527
R1844 a_13367_411.n1 a_13367_411.t12 384.527
R1845 a_13367_411.n7 a_13367_411.t7 294.278
R1846 a_13367_411.n4 a_13367_411.t13 294.278
R1847 a_13367_411.n2 a_13367_411.t9 294.278
R1848 a_13367_411.n12 a_13367_411.n11 281.733
R1849 a_13367_411.n13 a_13367_411.n12 117.693
R1850 a_13367_411.n5 a_13367_411.n2 80.851
R1851 a_13367_411.n8 a_13367_411.n7 80.035
R1852 a_13367_411.n15 a_13367_411.n14 79.232
R1853 a_13367_411.n5 a_13367_411.n4 76
R1854 a_13367_411.n12 a_13367_411.n8 76
R1855 a_13367_411.n15 a_13367_411.n13 63.152
R1856 a_13367_411.n2 a_13367_411.n1 57.842
R1857 a_13367_411.n7 a_13367_411.n6 56.954
R1858 a_13367_411.n4 a_13367_411.n3 56.833
R1859 a_13367_411.n11 a_13367_411.n10 22.578
R1860 a_13367_411.n13 a_13367_411.n0 16.08
R1861 a_13367_411.n16 a_13367_411.n15 16.078
R1862 a_13367_411.n0 a_13367_411.t4 14.282
R1863 a_13367_411.n0 a_13367_411.t3 14.282
R1864 a_13367_411.n14 a_13367_411.t0 14.282
R1865 a_13367_411.n14 a_13367_411.t6 14.282
R1866 a_13367_411.t2 a_13367_411.n16 14.282
R1867 a_13367_411.n16 a_13367_411.t1 14.282
R1868 a_13367_411.n11 a_13367_411.n9 8.58
R1869 a_13367_411.n8 a_13367_411.n5 1.859
R1870 a_13136_101.t0 a_13136_101.n1 93.333
R1871 a_13136_101.n4 a_13136_101.n2 55.07
R1872 a_13136_101.t0 a_13136_101.n0 8.137
R1873 a_13136_101.n4 a_13136_101.n3 4.619
R1874 a_13136_101.t0 a_13136_101.n4 0.071
R1875 a_13241_1050.n0 a_13241_1050.t5 512.525
R1876 a_13241_1050.n0 a_13241_1050.t6 371.139
R1877 a_13241_1050.n1 a_13241_1050.t7 368.112
R1878 a_13241_1050.n3 a_13241_1050.n2 311.99
R1879 a_13241_1050.n3 a_13241_1050.n1 126.657
R1880 a_13241_1050.n1 a_13241_1050.n0 79.811
R1881 a_13241_1050.n5 a_13241_1050.n4 76.002
R1882 a_13241_1050.n5 a_13241_1050.n3 72.841
R1883 a_13241_1050.n4 a_13241_1050.t3 14.282
R1884 a_13241_1050.n4 a_13241_1050.t4 14.282
R1885 a_13241_1050.n6 a_13241_1050.t1 14.282
R1886 a_13241_1050.t2 a_13241_1050.n6 14.282
R1887 a_13241_1050.n6 a_13241_1050.n5 12.848
R1888 a_4013_103.t0 a_4013_103.n3 117.777
R1889 a_4013_103.n6 a_4013_103.n5 45.444
R1890 a_4013_103.t0 a_4013_103.n6 21.213
R1891 a_4013_103.t0 a_4013_103.n4 11.595
R1892 a_4013_103.n2 a_4013_103.n0 8.543
R1893 a_4013_103.t0 a_4013_103.n2 3.034
R1894 a_4013_103.n2 a_4013_103.n1 0.443
R1895 a_4294_210.n8 a_4294_210.n6 96.467
R1896 a_4294_210.n3 a_4294_210.n1 44.628
R1897 a_4294_210.t0 a_4294_210.n8 32.417
R1898 a_4294_210.n3 a_4294_210.n2 23.284
R1899 a_4294_210.n6 a_4294_210.n5 22.349
R1900 a_4294_210.t0 a_4294_210.n10 20.241
R1901 a_4294_210.n10 a_4294_210.n9 13.494
R1902 a_4294_210.n6 a_4294_210.n4 8.443
R1903 a_4294_210.t0 a_4294_210.n0 8.137
R1904 a_4294_210.t0 a_4294_210.n3 5.727
R1905 a_4294_210.n8 a_4294_210.n7 1.435
R1906 a_9985_1050.n5 a_9985_1050.t9 512.525
R1907 a_9985_1050.n3 a_9985_1050.t8 512.525
R1908 a_9985_1050.n5 a_9985_1050.t7 371.139
R1909 a_9985_1050.n3 a_9985_1050.t6 371.139
R1910 a_9985_1050.n4 a_9985_1050.t5 234.562
R1911 a_9985_1050.n6 a_9985_1050.t10 234.204
R1912 a_9985_1050.n6 a_9985_1050.n5 216.178
R1913 a_9985_1050.n4 a_9985_1050.n3 215.819
R1914 a_9985_1050.n8 a_9985_1050.n2 205.605
R1915 a_9985_1050.n10 a_9985_1050.n8 164.008
R1916 a_9985_1050.n7 a_9985_1050.n4 79.488
R1917 a_9985_1050.n8 a_9985_1050.n7 77.314
R1918 a_9985_1050.n2 a_9985_1050.n1 76.002
R1919 a_9985_1050.n7 a_9985_1050.n6 76
R1920 a_9985_1050.n10 a_9985_1050.n9 15.218
R1921 a_9985_1050.n0 a_9985_1050.t1 14.282
R1922 a_9985_1050.n0 a_9985_1050.t4 14.282
R1923 a_9985_1050.n1 a_9985_1050.t3 14.282
R1924 a_9985_1050.n1 a_9985_1050.t0 14.282
R1925 a_9985_1050.n2 a_9985_1050.n0 12.85
R1926 a_9985_1050.n11 a_9985_1050.n10 12.014
R1927 a_11487_103.t0 a_11487_103.n3 117.777
R1928 a_11487_103.n6 a_11487_103.n5 45.444
R1929 a_11487_103.t0 a_11487_103.n6 21.213
R1930 a_11487_103.t0 a_11487_103.n4 11.595
R1931 a_11487_103.n2 a_11487_103.n0 8.543
R1932 a_11487_103.t0 a_11487_103.n2 3.034
R1933 a_11487_103.n2 a_11487_103.n1 0.443
R1934 GND.n30 GND.n29 219.745
R1935 GND.n63 GND.n61 219.745
R1936 GND.n96 GND.n94 219.745
R1937 GND.n436 GND.n435 219.745
R1938 GND.n478 GND.n476 219.745
R1939 GND.n520 GND.n518 219.745
R1940 GND.n550 GND.n548 219.745
R1941 GND.n580 GND.n578 219.745
R1942 GND.n622 GND.n620 219.745
R1943 GND.n652 GND.n650 219.745
R1944 GND.n694 GND.n692 219.745
R1945 GND.n736 GND.n734 219.745
R1946 GND.n766 GND.n764 219.745
R1947 GND.n396 GND.n394 219.745
R1948 GND.n351 GND.n349 219.745
R1949 GND.n321 GND.n319 219.745
R1950 GND.n276 GND.n274 219.745
R1951 GND.n234 GND.n232 219.745
R1952 GND.n204 GND.n202 219.745
R1953 GND.n174 GND.n172 219.745
R1954 GND.n129 GND.n128 219.745
R1955 GND.n265 GND.n264 85.559
R1956 GND.n703 GND.n702 85.559
R1957 GND.n661 GND.n660 85.559
R1958 GND.n589 GND.n588 85.559
R1959 GND.n487 GND.n486 85.559
R1960 GND.n445 GND.n444 85.559
R1961 GND.n30 GND.n28 85.529
R1962 GND.n63 GND.n62 85.529
R1963 GND.n96 GND.n95 85.529
R1964 GND.n436 GND.n434 85.529
R1965 GND.n478 GND.n477 85.529
R1966 GND.n520 GND.n519 85.529
R1967 GND.n550 GND.n549 85.529
R1968 GND.n580 GND.n579 85.529
R1969 GND.n622 GND.n621 85.529
R1970 GND.n652 GND.n651 85.529
R1971 GND.n694 GND.n693 85.529
R1972 GND.n736 GND.n735 85.529
R1973 GND.n766 GND.n765 85.529
R1974 GND.n396 GND.n395 85.529
R1975 GND.n351 GND.n350 85.529
R1976 GND.n321 GND.n320 85.529
R1977 GND.n276 GND.n275 85.529
R1978 GND.n234 GND.n233 85.529
R1979 GND.n204 GND.n203 85.529
R1980 GND.n174 GND.n173 85.529
R1981 GND.n129 GND.n127 85.529
R1982 GND.n192 GND.n191 84.842
R1983 GND.n222 GND.n221 84.842
R1984 GND.n339 GND.n338 84.842
R1985 GND.n774 GND.n773 84.842
R1986 GND.n744 GND.n743 84.842
R1987 GND.n630 GND.n629 84.842
R1988 GND.n558 GND.n557 84.842
R1989 GND.n528 GND.n527 84.842
R1990 GND.n414 GND.n413 84.842
R1991 GND.n9 GND.n1 76.145
R1992 GND.n409 GND.n408 76
R1993 GND.n76 GND.n75 76
R1994 GND.n79 GND.n78 76
R1995 GND.n87 GND.n86 76
R1996 GND.n90 GND.n89 76
R1997 GND.n93 GND.n92 76
R1998 GND.n100 GND.n99 76
R1999 GND.n103 GND.n102 76
R2000 GND.n106 GND.n105 76
R2001 GND.n109 GND.n108 76
R2002 GND.n112 GND.n111 76
R2003 GND.n120 GND.n119 76
R2004 GND.n123 GND.n122 76
R2005 GND.n126 GND.n125 76
R2006 GND.n133 GND.n132 76
R2007 GND.n136 GND.n135 76
R2008 GND.n139 GND.n138 76
R2009 GND.n142 GND.n141 76
R2010 GND.n145 GND.n144 76
R2011 GND.n148 GND.n147 76
R2012 GND.n151 GND.n150 76
R2013 GND.n154 GND.n153 76
R2014 GND.n157 GND.n156 76
R2015 GND.n165 GND.n164 76
R2016 GND.n168 GND.n167 76
R2017 GND.n171 GND.n170 76
R2018 GND.n178 GND.n177 76
R2019 GND.n181 GND.n180 76
R2020 GND.n184 GND.n183 76
R2021 GND.n187 GND.n186 76
R2022 GND.n190 GND.n189 76
R2023 GND.n195 GND.n194 76
R2024 GND.n198 GND.n197 76
R2025 GND.n201 GND.n200 76
R2026 GND.n208 GND.n207 76
R2027 GND.n211 GND.n210 76
R2028 GND.n214 GND.n213 76
R2029 GND.n217 GND.n216 76
R2030 GND.n220 GND.n219 76
R2031 GND.n225 GND.n224 76
R2032 GND.n228 GND.n227 76
R2033 GND.n231 GND.n230 76
R2034 GND.n238 GND.n237 76
R2035 GND.n241 GND.n240 76
R2036 GND.n244 GND.n243 76
R2037 GND.n247 GND.n246 76
R2038 GND.n250 GND.n249 76
R2039 GND.n253 GND.n252 76
R2040 GND.n256 GND.n255 76
R2041 GND.n259 GND.n258 76
R2042 GND.n262 GND.n261 76
R2043 GND.n267 GND.n266 76
R2044 GND.n270 GND.n269 76
R2045 GND.n273 GND.n272 76
R2046 GND.n280 GND.n279 76
R2047 GND.n283 GND.n282 76
R2048 GND.n286 GND.n285 76
R2049 GND.n289 GND.n288 76
R2050 GND.n292 GND.n291 76
R2051 GND.n295 GND.n294 76
R2052 GND.n298 GND.n297 76
R2053 GND.n301 GND.n300 76
R2054 GND.n304 GND.n303 76
R2055 GND.n312 GND.n311 76
R2056 GND.n315 GND.n314 76
R2057 GND.n318 GND.n317 76
R2058 GND.n325 GND.n324 76
R2059 GND.n328 GND.n327 76
R2060 GND.n331 GND.n330 76
R2061 GND.n334 GND.n333 76
R2062 GND.n337 GND.n336 76
R2063 GND.n342 GND.n341 76
R2064 GND.n345 GND.n344 76
R2065 GND.n348 GND.n347 76
R2066 GND.n355 GND.n354 76
R2067 GND.n358 GND.n357 76
R2068 GND.n361 GND.n360 76
R2069 GND.n364 GND.n363 76
R2070 GND.n367 GND.n366 76
R2071 GND.n370 GND.n369 76
R2072 GND.n373 GND.n372 76
R2073 GND.n376 GND.n375 76
R2074 GND.n379 GND.n378 76
R2075 GND.n387 GND.n386 76
R2076 GND.n390 GND.n389 76
R2077 GND.n393 GND.n392 76
R2078 GND.n400 GND.n399 76
R2079 GND.n403 GND.n402 76
R2080 GND.n406 GND.n405 76
R2081 GND.n783 GND.n782 76
R2082 GND.n780 GND.n779 76
R2083 GND.n777 GND.n776 76
R2084 GND.n772 GND.n771 76
R2085 GND.n769 GND.n768 76
R2086 GND.n762 GND.n761 76
R2087 GND.n759 GND.n758 76
R2088 GND.n756 GND.n755 76
R2089 GND.n753 GND.n752 76
R2090 GND.n750 GND.n749 76
R2091 GND.n747 GND.n746 76
R2092 GND.n742 GND.n741 76
R2093 GND.n739 GND.n738 76
R2094 GND.n732 GND.n731 76
R2095 GND.n729 GND.n728 76
R2096 GND.n726 GND.n725 76
R2097 GND.n723 GND.n722 76
R2098 GND.n720 GND.n719 76
R2099 GND.n717 GND.n716 76
R2100 GND.n714 GND.n713 76
R2101 GND.n711 GND.n710 76
R2102 GND.n708 GND.n707 76
R2103 GND.n705 GND.n704 76
R2104 GND.n700 GND.n699 76
R2105 GND.n697 GND.n696 76
R2106 GND.n690 GND.n689 76
R2107 GND.n687 GND.n686 76
R2108 GND.n684 GND.n683 76
R2109 GND.n681 GND.n680 76
R2110 GND.n678 GND.n677 76
R2111 GND.n675 GND.n674 76
R2112 GND.n672 GND.n671 76
R2113 GND.n669 GND.n668 76
R2114 GND.n666 GND.n665 76
R2115 GND.n663 GND.n662 76
R2116 GND.n658 GND.n657 76
R2117 GND.n655 GND.n654 76
R2118 GND.n648 GND.n647 76
R2119 GND.n645 GND.n644 76
R2120 GND.n642 GND.n641 76
R2121 GND.n639 GND.n638 76
R2122 GND.n636 GND.n635 76
R2123 GND.n633 GND.n632 76
R2124 GND.n628 GND.n627 76
R2125 GND.n625 GND.n624 76
R2126 GND.n618 GND.n617 76
R2127 GND.n615 GND.n614 76
R2128 GND.n612 GND.n611 76
R2129 GND.n609 GND.n608 76
R2130 GND.n606 GND.n605 76
R2131 GND.n603 GND.n602 76
R2132 GND.n600 GND.n599 76
R2133 GND.n597 GND.n596 76
R2134 GND.n594 GND.n593 76
R2135 GND.n591 GND.n590 76
R2136 GND.n586 GND.n585 76
R2137 GND.n583 GND.n582 76
R2138 GND.n576 GND.n575 76
R2139 GND.n573 GND.n572 76
R2140 GND.n570 GND.n569 76
R2141 GND.n567 GND.n566 76
R2142 GND.n564 GND.n563 76
R2143 GND.n561 GND.n560 76
R2144 GND.n556 GND.n555 76
R2145 GND.n553 GND.n552 76
R2146 GND.n546 GND.n545 76
R2147 GND.n543 GND.n542 76
R2148 GND.n540 GND.n539 76
R2149 GND.n537 GND.n536 76
R2150 GND.n534 GND.n533 76
R2151 GND.n531 GND.n530 76
R2152 GND.n526 GND.n525 76
R2153 GND.n523 GND.n522 76
R2154 GND.n516 GND.n515 76
R2155 GND.n513 GND.n512 76
R2156 GND.n510 GND.n509 76
R2157 GND.n507 GND.n506 76
R2158 GND.n504 GND.n503 76
R2159 GND.n501 GND.n500 76
R2160 GND.n498 GND.n497 76
R2161 GND.n495 GND.n494 76
R2162 GND.n492 GND.n491 76
R2163 GND.n489 GND.n488 76
R2164 GND.n484 GND.n483 76
R2165 GND.n481 GND.n480 76
R2166 GND.n474 GND.n473 76
R2167 GND.n471 GND.n470 76
R2168 GND.n468 GND.n467 76
R2169 GND.n465 GND.n464 76
R2170 GND.n462 GND.n461 76
R2171 GND.n459 GND.n458 76
R2172 GND.n456 GND.n455 76
R2173 GND.n453 GND.n452 76
R2174 GND.n450 GND.n449 76
R2175 GND.n447 GND.n446 76
R2176 GND.n442 GND.n441 76
R2177 GND.n439 GND.n438 76
R2178 GND.n432 GND.n431 76
R2179 GND.n429 GND.n428 76
R2180 GND.n426 GND.n425 76
R2181 GND.n423 GND.n422 76
R2182 GND.n420 GND.n419 76
R2183 GND.n417 GND.n416 76
R2184 GND.n412 GND.n411 76
R2185 GND.n9 GND.n8 76
R2186 GND.n17 GND.n16 76
R2187 GND.n24 GND.n23 76
R2188 GND.n27 GND.n26 76
R2189 GND.n34 GND.n33 76
R2190 GND.n37 GND.n36 76
R2191 GND.n40 GND.n39 76
R2192 GND.n43 GND.n42 76
R2193 GND.n46 GND.n45 76
R2194 GND.n54 GND.n53 76
R2195 GND.n57 GND.n56 76
R2196 GND.n60 GND.n59 76
R2197 GND.n67 GND.n66 76
R2198 GND.n70 GND.n69 76
R2199 GND.n73 GND.n72 76
R2200 GND.n163 GND.n162 64.552
R2201 GND.n310 GND.n309 64.552
R2202 GND.n385 GND.n384 64.552
R2203 GND.n84 GND.n83 63.835
R2204 GND.n117 GND.n116 63.835
R2205 GND.n51 GND.n50 63.835
R2206 GND.n5 GND.n4 35.01
R2207 GND.n3 GND.n2 29.127
R2208 GND.n83 GND.n82 28.421
R2209 GND.n116 GND.n115 28.421
R2210 GND.n162 GND.n161 28.421
R2211 GND.n309 GND.n308 28.421
R2212 GND.n384 GND.n383 28.421
R2213 GND.n50 GND.n49 28.421
R2214 GND.n83 GND.n81 25.263
R2215 GND.n116 GND.n114 25.263
R2216 GND.n162 GND.n160 25.263
R2217 GND.n309 GND.n307 25.263
R2218 GND.n384 GND.n382 25.263
R2219 GND.n50 GND.n48 25.263
R2220 GND.n81 GND.n80 24.383
R2221 GND.n114 GND.n113 24.383
R2222 GND.n160 GND.n159 24.383
R2223 GND.n307 GND.n306 24.383
R2224 GND.n382 GND.n381 24.383
R2225 GND.n48 GND.n47 24.383
R2226 GND.n12 GND.t5 20.794
R2227 GND.n6 GND.n5 19.735
R2228 GND.n14 GND.n13 19.735
R2229 GND.n21 GND.n20 19.735
R2230 GND.n5 GND.n3 19.017
R2231 GND.n33 GND.n31 14.167
R2232 GND.n66 GND.n64 14.167
R2233 GND.n99 GND.n97 14.167
R2234 GND.n132 GND.n130 14.167
R2235 GND.n177 GND.n175 14.167
R2236 GND.n207 GND.n205 14.167
R2237 GND.n237 GND.n235 14.167
R2238 GND.n279 GND.n277 14.167
R2239 GND.n324 GND.n322 14.167
R2240 GND.n354 GND.n352 14.167
R2241 GND.n399 GND.n397 14.167
R2242 GND.n768 GND.n767 14.167
R2243 GND.n738 GND.n737 14.167
R2244 GND.n696 GND.n695 14.167
R2245 GND.n654 GND.n653 14.167
R2246 GND.n624 GND.n623 14.167
R2247 GND.n582 GND.n581 14.167
R2248 GND.n552 GND.n551 14.167
R2249 GND.n522 GND.n521 14.167
R2250 GND.n480 GND.n479 14.167
R2251 GND.n438 GND.n437 14.167
R2252 GND.n411 GND.n410 13.653
R2253 GND.n416 GND.n415 13.653
R2254 GND.n419 GND.n418 13.653
R2255 GND.n422 GND.n421 13.653
R2256 GND.n425 GND.n424 13.653
R2257 GND.n428 GND.n427 13.653
R2258 GND.n431 GND.n430 13.653
R2259 GND.n438 GND.n433 13.653
R2260 GND.n441 GND.n440 13.653
R2261 GND.n446 GND.n443 13.653
R2262 GND.n449 GND.n448 13.653
R2263 GND.n452 GND.n451 13.653
R2264 GND.n455 GND.n454 13.653
R2265 GND.n458 GND.n457 13.653
R2266 GND.n461 GND.n460 13.653
R2267 GND.n464 GND.n463 13.653
R2268 GND.n467 GND.n466 13.653
R2269 GND.n470 GND.n469 13.653
R2270 GND.n473 GND.n472 13.653
R2271 GND.n480 GND.n475 13.653
R2272 GND.n483 GND.n482 13.653
R2273 GND.n488 GND.n485 13.653
R2274 GND.n491 GND.n490 13.653
R2275 GND.n494 GND.n493 13.653
R2276 GND.n497 GND.n496 13.653
R2277 GND.n500 GND.n499 13.653
R2278 GND.n503 GND.n502 13.653
R2279 GND.n506 GND.n505 13.653
R2280 GND.n509 GND.n508 13.653
R2281 GND.n512 GND.n511 13.653
R2282 GND.n515 GND.n514 13.653
R2283 GND.n522 GND.n517 13.653
R2284 GND.n525 GND.n524 13.653
R2285 GND.n530 GND.n529 13.653
R2286 GND.n533 GND.n532 13.653
R2287 GND.n536 GND.n535 13.653
R2288 GND.n539 GND.n538 13.653
R2289 GND.n542 GND.n541 13.653
R2290 GND.n545 GND.n544 13.653
R2291 GND.n552 GND.n547 13.653
R2292 GND.n555 GND.n554 13.653
R2293 GND.n560 GND.n559 13.653
R2294 GND.n563 GND.n562 13.653
R2295 GND.n566 GND.n565 13.653
R2296 GND.n569 GND.n568 13.653
R2297 GND.n572 GND.n571 13.653
R2298 GND.n575 GND.n574 13.653
R2299 GND.n582 GND.n577 13.653
R2300 GND.n585 GND.n584 13.653
R2301 GND.n590 GND.n587 13.653
R2302 GND.n593 GND.n592 13.653
R2303 GND.n596 GND.n595 13.653
R2304 GND.n599 GND.n598 13.653
R2305 GND.n602 GND.n601 13.653
R2306 GND.n605 GND.n604 13.653
R2307 GND.n608 GND.n607 13.653
R2308 GND.n611 GND.n610 13.653
R2309 GND.n614 GND.n613 13.653
R2310 GND.n617 GND.n616 13.653
R2311 GND.n624 GND.n619 13.653
R2312 GND.n627 GND.n626 13.653
R2313 GND.n632 GND.n631 13.653
R2314 GND.n635 GND.n634 13.653
R2315 GND.n638 GND.n637 13.653
R2316 GND.n641 GND.n640 13.653
R2317 GND.n644 GND.n643 13.653
R2318 GND.n647 GND.n646 13.653
R2319 GND.n654 GND.n649 13.653
R2320 GND.n657 GND.n656 13.653
R2321 GND.n662 GND.n659 13.653
R2322 GND.n665 GND.n664 13.653
R2323 GND.n668 GND.n667 13.653
R2324 GND.n671 GND.n670 13.653
R2325 GND.n674 GND.n673 13.653
R2326 GND.n677 GND.n676 13.653
R2327 GND.n680 GND.n679 13.653
R2328 GND.n683 GND.n682 13.653
R2329 GND.n686 GND.n685 13.653
R2330 GND.n689 GND.n688 13.653
R2331 GND.n696 GND.n691 13.653
R2332 GND.n699 GND.n698 13.653
R2333 GND.n704 GND.n701 13.653
R2334 GND.n707 GND.n706 13.653
R2335 GND.n710 GND.n709 13.653
R2336 GND.n713 GND.n712 13.653
R2337 GND.n716 GND.n715 13.653
R2338 GND.n719 GND.n718 13.653
R2339 GND.n722 GND.n721 13.653
R2340 GND.n725 GND.n724 13.653
R2341 GND.n728 GND.n727 13.653
R2342 GND.n731 GND.n730 13.653
R2343 GND.n738 GND.n733 13.653
R2344 GND.n741 GND.n740 13.653
R2345 GND.n746 GND.n745 13.653
R2346 GND.n749 GND.n748 13.653
R2347 GND.n752 GND.n751 13.653
R2348 GND.n755 GND.n754 13.653
R2349 GND.n758 GND.n757 13.653
R2350 GND.n761 GND.n760 13.653
R2351 GND.n768 GND.n763 13.653
R2352 GND.n771 GND.n770 13.653
R2353 GND.n776 GND.n775 13.653
R2354 GND.n779 GND.n778 13.653
R2355 GND.n782 GND.n781 13.653
R2356 GND.n405 GND.n404 13.653
R2357 GND.n402 GND.n401 13.653
R2358 GND.n399 GND.n398 13.653
R2359 GND.n392 GND.n391 13.653
R2360 GND.n389 GND.n388 13.653
R2361 GND.n386 GND.n380 13.653
R2362 GND.n378 GND.n377 13.653
R2363 GND.n375 GND.n374 13.653
R2364 GND.n372 GND.n371 13.653
R2365 GND.n369 GND.n368 13.653
R2366 GND.n366 GND.n365 13.653
R2367 GND.n363 GND.n362 13.653
R2368 GND.n360 GND.n359 13.653
R2369 GND.n357 GND.n356 13.653
R2370 GND.n354 GND.n353 13.653
R2371 GND.n347 GND.n346 13.653
R2372 GND.n344 GND.n343 13.653
R2373 GND.n341 GND.n340 13.653
R2374 GND.n336 GND.n335 13.653
R2375 GND.n333 GND.n332 13.653
R2376 GND.n330 GND.n329 13.653
R2377 GND.n327 GND.n326 13.653
R2378 GND.n324 GND.n323 13.653
R2379 GND.n317 GND.n316 13.653
R2380 GND.n314 GND.n313 13.653
R2381 GND.n311 GND.n305 13.653
R2382 GND.n303 GND.n302 13.653
R2383 GND.n300 GND.n299 13.653
R2384 GND.n297 GND.n296 13.653
R2385 GND.n294 GND.n293 13.653
R2386 GND.n291 GND.n290 13.653
R2387 GND.n288 GND.n287 13.653
R2388 GND.n285 GND.n284 13.653
R2389 GND.n282 GND.n281 13.653
R2390 GND.n279 GND.n278 13.653
R2391 GND.n272 GND.n271 13.653
R2392 GND.n269 GND.n268 13.653
R2393 GND.n266 GND.n263 13.653
R2394 GND.n261 GND.n260 13.653
R2395 GND.n258 GND.n257 13.653
R2396 GND.n255 GND.n254 13.653
R2397 GND.n252 GND.n251 13.653
R2398 GND.n249 GND.n248 13.653
R2399 GND.n246 GND.n245 13.653
R2400 GND.n243 GND.n242 13.653
R2401 GND.n240 GND.n239 13.653
R2402 GND.n237 GND.n236 13.653
R2403 GND.n230 GND.n229 13.653
R2404 GND.n227 GND.n226 13.653
R2405 GND.n224 GND.n223 13.653
R2406 GND.n219 GND.n218 13.653
R2407 GND.n216 GND.n215 13.653
R2408 GND.n213 GND.n212 13.653
R2409 GND.n210 GND.n209 13.653
R2410 GND.n207 GND.n206 13.653
R2411 GND.n200 GND.n199 13.653
R2412 GND.n197 GND.n196 13.653
R2413 GND.n194 GND.n193 13.653
R2414 GND.n189 GND.n188 13.653
R2415 GND.n186 GND.n185 13.653
R2416 GND.n183 GND.n182 13.653
R2417 GND.n180 GND.n179 13.653
R2418 GND.n177 GND.n176 13.653
R2419 GND.n170 GND.n169 13.653
R2420 GND.n167 GND.n166 13.653
R2421 GND.n164 GND.n158 13.653
R2422 GND.n156 GND.n155 13.653
R2423 GND.n153 GND.n152 13.653
R2424 GND.n150 GND.n149 13.653
R2425 GND.n147 GND.n146 13.653
R2426 GND.n144 GND.n143 13.653
R2427 GND.n141 GND.n140 13.653
R2428 GND.n138 GND.n137 13.653
R2429 GND.n135 GND.n134 13.653
R2430 GND.n132 GND.n131 13.653
R2431 GND.n125 GND.n124 13.653
R2432 GND.n122 GND.n121 13.653
R2433 GND.n119 GND.n118 13.653
R2434 GND.n111 GND.n110 13.653
R2435 GND.n108 GND.n107 13.653
R2436 GND.n105 GND.n104 13.653
R2437 GND.n102 GND.n101 13.653
R2438 GND.n99 GND.n98 13.653
R2439 GND.n92 GND.n91 13.653
R2440 GND.n89 GND.n88 13.653
R2441 GND.n86 GND.n85 13.653
R2442 GND.n78 GND.n77 13.653
R2443 GND.n75 GND.n74 13.653
R2444 GND.n8 GND.n7 13.653
R2445 GND.n16 GND.n15 13.653
R2446 GND.n23 GND.n22 13.653
R2447 GND.n26 GND.n25 13.653
R2448 GND.n33 GND.n32 13.653
R2449 GND.n36 GND.n35 13.653
R2450 GND.n39 GND.n38 13.653
R2451 GND.n42 GND.n41 13.653
R2452 GND.n45 GND.n44 13.653
R2453 GND.n53 GND.n52 13.653
R2454 GND.n56 GND.n55 13.653
R2455 GND.n59 GND.n58 13.653
R2456 GND.n66 GND.n65 13.653
R2457 GND.n69 GND.n68 13.653
R2458 GND.n72 GND.n71 13.653
R2459 GND.n20 GND.n19 12.837
R2460 GND.n19 GND.n18 7.566
R2461 GND.n31 GND.n30 7.312
R2462 GND.n64 GND.n63 7.312
R2463 GND.n97 GND.n96 7.312
R2464 GND.n437 GND.n436 7.312
R2465 GND.n479 GND.n478 7.312
R2466 GND.n521 GND.n520 7.312
R2467 GND.n551 GND.n550 7.312
R2468 GND.n581 GND.n580 7.312
R2469 GND.n623 GND.n622 7.312
R2470 GND.n653 GND.n652 7.312
R2471 GND.n695 GND.n694 7.312
R2472 GND.n737 GND.n736 7.312
R2473 GND.n767 GND.n766 7.312
R2474 GND.n397 GND.n396 7.312
R2475 GND.n352 GND.n351 7.312
R2476 GND.n322 GND.n321 7.312
R2477 GND.n277 GND.n276 7.312
R2478 GND.n235 GND.n234 7.312
R2479 GND.n205 GND.n204 7.312
R2480 GND.n175 GND.n174 7.312
R2481 GND.n130 GND.n129 7.312
R2482 GND.n11 GND.n10 4.551
R2483 GND.n8 GND.n6 3.935
R2484 GND.n53 GND.n51 3.935
R2485 GND.n86 GND.n84 3.935
R2486 GND.n119 GND.n117 3.935
R2487 GND.n194 GND.n192 3.935
R2488 GND.n224 GND.n222 3.935
R2489 GND.n341 GND.n339 3.935
R2490 GND.n776 GND.n774 3.935
R2491 GND.n746 GND.n744 3.935
R2492 GND.n632 GND.n630 3.935
R2493 GND.n560 GND.n558 3.935
R2494 GND.n530 GND.n528 3.935
R2495 GND.n416 GND.n414 3.935
R2496 GND.n23 GND.n21 3.541
R2497 GND.t5 GND.n11 2.238
R2498 GND.n408 GND.n407 0.596
R2499 GND.n1 GND.n0 0.596
R2500 GND.n13 GND.n12 0.358
R2501 GND.n34 GND.n27 0.29
R2502 GND.n67 GND.n60 0.29
R2503 GND.n100 GND.n93 0.29
R2504 GND.n133 GND.n126 0.29
R2505 GND.n178 GND.n171 0.29
R2506 GND.n208 GND.n201 0.29
R2507 GND.n238 GND.n231 0.29
R2508 GND.n280 GND.n273 0.29
R2509 GND.n325 GND.n318 0.29
R2510 GND.n355 GND.n348 0.29
R2511 GND.n400 GND.n393 0.29
R2512 GND.n769 GND.n762 0.29
R2513 GND.n739 GND.n732 0.29
R2514 GND.n697 GND.n690 0.29
R2515 GND.n655 GND.n648 0.29
R2516 GND.n625 GND.n618 0.29
R2517 GND.n583 GND.n576 0.29
R2518 GND.n553 GND.n546 0.29
R2519 GND.n523 GND.n516 0.29
R2520 GND.n481 GND.n474 0.29
R2521 GND.n439 GND.n432 0.29
R2522 GND.n409 GND 0.207
R2523 GND.n151 GND.n148 0.197
R2524 GND.n256 GND.n253 0.197
R2525 GND.n298 GND.n295 0.197
R2526 GND.n373 GND.n370 0.197
R2527 GND.n717 GND.n714 0.197
R2528 GND.n675 GND.n672 0.197
R2529 GND.n603 GND.n600 0.197
R2530 GND.n501 GND.n498 0.197
R2531 GND.n459 GND.n456 0.197
R2532 GND.n16 GND.n14 0.196
R2533 GND.n164 GND.n163 0.196
R2534 GND.n266 GND.n265 0.196
R2535 GND.n311 GND.n310 0.196
R2536 GND.n386 GND.n385 0.196
R2537 GND.n704 GND.n703 0.196
R2538 GND.n662 GND.n661 0.196
R2539 GND.n590 GND.n589 0.196
R2540 GND.n488 GND.n487 0.196
R2541 GND.n446 GND.n445 0.196
R2542 GND.n46 GND.n43 0.181
R2543 GND.n79 GND.n76 0.181
R2544 GND.n112 GND.n109 0.181
R2545 GND.n190 GND.n187 0.181
R2546 GND.n220 GND.n217 0.181
R2547 GND.n337 GND.n334 0.181
R2548 GND.n783 GND.n780 0.181
R2549 GND.n753 GND.n750 0.181
R2550 GND.n639 GND.n636 0.181
R2551 GND.n567 GND.n564 0.181
R2552 GND.n537 GND.n534 0.181
R2553 GND.n423 GND.n420 0.181
R2554 GND.n17 GND.n9 0.157
R2555 GND.n24 GND.n17 0.157
R2556 GND.n27 GND.n24 0.145
R2557 GND.n37 GND.n34 0.145
R2558 GND.n40 GND.n37 0.145
R2559 GND.n43 GND.n40 0.145
R2560 GND.n54 GND.n46 0.145
R2561 GND.n57 GND.n54 0.145
R2562 GND.n60 GND.n57 0.145
R2563 GND.n70 GND.n67 0.145
R2564 GND.n73 GND.n70 0.145
R2565 GND.n76 GND.n73 0.145
R2566 GND.n87 GND.n79 0.145
R2567 GND.n90 GND.n87 0.145
R2568 GND.n93 GND.n90 0.145
R2569 GND.n103 GND.n100 0.145
R2570 GND.n106 GND.n103 0.145
R2571 GND.n109 GND.n106 0.145
R2572 GND.n120 GND.n112 0.145
R2573 GND.n123 GND.n120 0.145
R2574 GND.n126 GND.n123 0.145
R2575 GND.n136 GND.n133 0.145
R2576 GND.n139 GND.n136 0.145
R2577 GND.n142 GND.n139 0.145
R2578 GND.n145 GND.n142 0.145
R2579 GND.n148 GND.n145 0.145
R2580 GND.n154 GND.n151 0.145
R2581 GND.n157 GND.n154 0.145
R2582 GND.n165 GND.n157 0.145
R2583 GND.n168 GND.n165 0.145
R2584 GND.n171 GND.n168 0.145
R2585 GND.n181 GND.n178 0.145
R2586 GND.n184 GND.n181 0.145
R2587 GND.n187 GND.n184 0.145
R2588 GND.n195 GND.n190 0.145
R2589 GND.n198 GND.n195 0.145
R2590 GND.n201 GND.n198 0.145
R2591 GND.n211 GND.n208 0.145
R2592 GND.n214 GND.n211 0.145
R2593 GND.n217 GND.n214 0.145
R2594 GND.n225 GND.n220 0.145
R2595 GND.n228 GND.n225 0.145
R2596 GND.n231 GND.n228 0.145
R2597 GND.n241 GND.n238 0.145
R2598 GND.n244 GND.n241 0.145
R2599 GND.n247 GND.n244 0.145
R2600 GND.n250 GND.n247 0.145
R2601 GND.n253 GND.n250 0.145
R2602 GND.n259 GND.n256 0.145
R2603 GND.n262 GND.n259 0.145
R2604 GND.n267 GND.n262 0.145
R2605 GND.n270 GND.n267 0.145
R2606 GND.n273 GND.n270 0.145
R2607 GND.n283 GND.n280 0.145
R2608 GND.n286 GND.n283 0.145
R2609 GND.n289 GND.n286 0.145
R2610 GND.n292 GND.n289 0.145
R2611 GND.n295 GND.n292 0.145
R2612 GND.n301 GND.n298 0.145
R2613 GND.n304 GND.n301 0.145
R2614 GND.n312 GND.n304 0.145
R2615 GND.n315 GND.n312 0.145
R2616 GND.n318 GND.n315 0.145
R2617 GND.n328 GND.n325 0.145
R2618 GND.n331 GND.n328 0.145
R2619 GND.n334 GND.n331 0.145
R2620 GND.n342 GND.n337 0.145
R2621 GND.n345 GND.n342 0.145
R2622 GND.n348 GND.n345 0.145
R2623 GND.n358 GND.n355 0.145
R2624 GND.n361 GND.n358 0.145
R2625 GND.n364 GND.n361 0.145
R2626 GND.n367 GND.n364 0.145
R2627 GND.n370 GND.n367 0.145
R2628 GND.n376 GND.n373 0.145
R2629 GND.n379 GND.n376 0.145
R2630 GND.n387 GND.n379 0.145
R2631 GND.n390 GND.n387 0.145
R2632 GND.n393 GND.n390 0.145
R2633 GND.n403 GND.n400 0.145
R2634 GND.n406 GND.n403 0.145
R2635 GND.n780 GND.n777 0.145
R2636 GND.n777 GND.n772 0.145
R2637 GND.n772 GND.n769 0.145
R2638 GND.n762 GND.n759 0.145
R2639 GND.n759 GND.n756 0.145
R2640 GND.n756 GND.n753 0.145
R2641 GND.n750 GND.n747 0.145
R2642 GND.n747 GND.n742 0.145
R2643 GND.n742 GND.n739 0.145
R2644 GND.n732 GND.n729 0.145
R2645 GND.n729 GND.n726 0.145
R2646 GND.n726 GND.n723 0.145
R2647 GND.n723 GND.n720 0.145
R2648 GND.n720 GND.n717 0.145
R2649 GND.n714 GND.n711 0.145
R2650 GND.n711 GND.n708 0.145
R2651 GND.n708 GND.n705 0.145
R2652 GND.n705 GND.n700 0.145
R2653 GND.n700 GND.n697 0.145
R2654 GND.n690 GND.n687 0.145
R2655 GND.n687 GND.n684 0.145
R2656 GND.n684 GND.n681 0.145
R2657 GND.n681 GND.n678 0.145
R2658 GND.n678 GND.n675 0.145
R2659 GND.n672 GND.n669 0.145
R2660 GND.n669 GND.n666 0.145
R2661 GND.n666 GND.n663 0.145
R2662 GND.n663 GND.n658 0.145
R2663 GND.n658 GND.n655 0.145
R2664 GND.n648 GND.n645 0.145
R2665 GND.n645 GND.n642 0.145
R2666 GND.n642 GND.n639 0.145
R2667 GND.n636 GND.n633 0.145
R2668 GND.n633 GND.n628 0.145
R2669 GND.n628 GND.n625 0.145
R2670 GND.n618 GND.n615 0.145
R2671 GND.n615 GND.n612 0.145
R2672 GND.n612 GND.n609 0.145
R2673 GND.n609 GND.n606 0.145
R2674 GND.n606 GND.n603 0.145
R2675 GND.n600 GND.n597 0.145
R2676 GND.n597 GND.n594 0.145
R2677 GND.n594 GND.n591 0.145
R2678 GND.n591 GND.n586 0.145
R2679 GND.n586 GND.n583 0.145
R2680 GND.n576 GND.n573 0.145
R2681 GND.n573 GND.n570 0.145
R2682 GND.n570 GND.n567 0.145
R2683 GND.n564 GND.n561 0.145
R2684 GND.n561 GND.n556 0.145
R2685 GND.n556 GND.n553 0.145
R2686 GND.n546 GND.n543 0.145
R2687 GND.n543 GND.n540 0.145
R2688 GND.n540 GND.n537 0.145
R2689 GND.n534 GND.n531 0.145
R2690 GND.n531 GND.n526 0.145
R2691 GND.n526 GND.n523 0.145
R2692 GND.n516 GND.n513 0.145
R2693 GND.n513 GND.n510 0.145
R2694 GND.n510 GND.n507 0.145
R2695 GND.n507 GND.n504 0.145
R2696 GND.n504 GND.n501 0.145
R2697 GND.n498 GND.n495 0.145
R2698 GND.n495 GND.n492 0.145
R2699 GND.n492 GND.n489 0.145
R2700 GND.n489 GND.n484 0.145
R2701 GND.n484 GND.n481 0.145
R2702 GND.n474 GND.n471 0.145
R2703 GND.n471 GND.n468 0.145
R2704 GND.n468 GND.n465 0.145
R2705 GND.n465 GND.n462 0.145
R2706 GND.n462 GND.n459 0.145
R2707 GND.n456 GND.n453 0.145
R2708 GND.n453 GND.n450 0.145
R2709 GND.n450 GND.n447 0.145
R2710 GND.n447 GND.n442 0.145
R2711 GND.n442 GND.n439 0.145
R2712 GND.n432 GND.n429 0.145
R2713 GND.n429 GND.n426 0.145
R2714 GND.n426 GND.n423 0.145
R2715 GND.n420 GND.n417 0.145
R2716 GND.n417 GND.n412 0.145
R2717 GND.n412 GND.n409 0.145
R2718 GND GND.n406 0.086
R2719 GND GND.n783 0.058
R2720 a_15044_209.n4 a_15044_209.t8 512.525
R2721 a_15044_209.n4 a_15044_209.t7 371.139
R2722 a_15044_209.n5 a_15044_209.t9 263.54
R2723 a_15044_209.n10 a_15044_209.n6 216.728
R2724 a_15044_209.n6 a_15044_209.n5 153.043
R2725 a_15044_209.n6 a_15044_209.n3 126.664
R2726 a_15044_209.n5 a_15044_209.n4 120.094
R2727 a_15044_209.n15 a_15044_209.n14 98.501
R2728 a_15044_209.n17 a_15044_209.n15 96.417
R2729 a_15044_209.n9 a_15044_209.n7 80.526
R2730 a_15044_209.n15 a_15044_209.n10 78.403
R2731 a_15044_209.n3 a_15044_209.n2 75.271
R2732 a_15044_209.n14 a_15044_209.n13 30
R2733 a_15044_209.n9 a_15044_209.n8 30
R2734 a_15044_209.n17 a_15044_209.n16 30
R2735 a_15044_209.n12 a_15044_209.n11 24.383
R2736 a_15044_209.n18 a_15044_209.n0 24.383
R2737 a_15044_209.n14 a_15044_209.n12 23.684
R2738 a_15044_209.n18 a_15044_209.n17 23.684
R2739 a_15044_209.n10 a_15044_209.n9 20.417
R2740 a_15044_209.n1 a_15044_209.t4 14.282
R2741 a_15044_209.n1 a_15044_209.t6 14.282
R2742 a_15044_209.n2 a_15044_209.t1 14.282
R2743 a_15044_209.n2 a_15044_209.t2 14.282
R2744 a_15044_209.n3 a_15044_209.n1 12.119
R2745 Q.n2 Q.n1 253.86
R2746 Q.n2 Q.n0 130.901
R2747 Q.n3 Q.n2 76
R2748 Q.n0 Q.t0 14.282
R2749 Q.n0 Q.t1 14.282
R2750 Q.n3 Q 0.046
R2751 a_1265_989.n2 a_1265_989.t12 454.685
R2752 a_1265_989.n4 a_1265_989.t5 454.685
R2753 a_1265_989.n0 a_1265_989.t9 454.685
R2754 a_1265_989.n2 a_1265_989.t7 428.979
R2755 a_1265_989.n4 a_1265_989.t11 428.979
R2756 a_1265_989.n0 a_1265_989.t10 428.979
R2757 a_1265_989.n3 a_1265_989.t6 264.512
R2758 a_1265_989.n5 a_1265_989.t8 264.512
R2759 a_1265_989.n1 a_1265_989.t13 264.512
R2760 a_1265_989.n12 a_1265_989.n11 237.145
R2761 a_1265_989.n14 a_1265_989.n12 125.947
R2762 a_1265_989.n7 a_1265_989.n1 81.396
R2763 a_1265_989.n6 a_1265_989.n5 79.491
R2764 a_1265_989.n14 a_1265_989.n13 76.002
R2765 a_1265_989.n6 a_1265_989.n3 76
R2766 a_1265_989.n12 a_1265_989.n7 76
R2767 a_1265_989.n3 a_1265_989.n2 71.894
R2768 a_1265_989.n5 a_1265_989.n4 71.894
R2769 a_1265_989.n1 a_1265_989.n0 71.894
R2770 a_1265_989.n11 a_1265_989.n10 30
R2771 a_1265_989.n9 a_1265_989.n8 24.383
R2772 a_1265_989.n11 a_1265_989.n9 23.684
R2773 a_1265_989.n13 a_1265_989.t3 14.282
R2774 a_1265_989.n13 a_1265_989.t4 14.282
R2775 a_1265_989.n15 a_1265_989.t0 14.282
R2776 a_1265_989.t1 a_1265_989.n15 14.282
R2777 a_1265_989.n15 a_1265_989.n14 12.848
R2778 a_1265_989.n7 a_1265_989.n6 2.947
R2779 a_343_411.n1 a_343_411.t7 480.392
R2780 a_343_411.n3 a_343_411.t9 472.359
R2781 a_343_411.n1 a_343_411.t10 403.272
R2782 a_343_411.n3 a_343_411.t12 384.527
R2783 a_343_411.n2 a_343_411.t8 336.586
R2784 a_343_411.n4 a_343_411.t11 294.278
R2785 a_343_411.n10 a_343_411.n9 265.87
R2786 a_343_411.n11 a_343_411.n10 117.354
R2787 a_343_411.n5 a_343_411.n2 83.304
R2788 a_343_411.n5 a_343_411.n4 80.032
R2789 a_343_411.n13 a_343_411.n12 79.232
R2790 a_343_411.n10 a_343_411.n5 76
R2791 a_343_411.n13 a_343_411.n11 63.152
R2792 a_343_411.n4 a_343_411.n3 56.954
R2793 a_343_411.n2 a_343_411.n1 45.341
R2794 a_343_411.n9 a_343_411.n8 30
R2795 a_343_411.n7 a_343_411.n6 24.383
R2796 a_343_411.n9 a_343_411.n7 23.684
R2797 a_343_411.n11 a_343_411.n0 16.08
R2798 a_343_411.n14 a_343_411.n13 16.078
R2799 a_343_411.n0 a_343_411.t2 14.282
R2800 a_343_411.n0 a_343_411.t3 14.282
R2801 a_343_411.n12 a_343_411.t6 14.282
R2802 a_343_411.n12 a_343_411.t5 14.282
R2803 a_343_411.t1 a_343_411.n14 14.282
R2804 a_343_411.n14 a_343_411.t0 14.282
R2805 a_11033_989.n2 a_11033_989.t8 454.685
R2806 a_11033_989.n4 a_11033_989.t13 454.685
R2807 a_11033_989.n0 a_11033_989.t5 454.685
R2808 a_11033_989.n2 a_11033_989.t7 428.979
R2809 a_11033_989.n4 a_11033_989.t9 428.979
R2810 a_11033_989.n0 a_11033_989.t11 428.979
R2811 a_11033_989.n3 a_11033_989.t12 264.512
R2812 a_11033_989.n5 a_11033_989.t10 264.512
R2813 a_11033_989.n1 a_11033_989.t6 264.512
R2814 a_11033_989.n12 a_11033_989.n11 237.145
R2815 a_11033_989.n14 a_11033_989.n12 125.947
R2816 a_11033_989.n7 a_11033_989.n1 81.396
R2817 a_11033_989.n6 a_11033_989.n5 79.491
R2818 a_11033_989.n14 a_11033_989.n13 76.002
R2819 a_11033_989.n6 a_11033_989.n3 76
R2820 a_11033_989.n12 a_11033_989.n7 76
R2821 a_11033_989.n3 a_11033_989.n2 71.894
R2822 a_11033_989.n5 a_11033_989.n4 71.894
R2823 a_11033_989.n1 a_11033_989.n0 71.894
R2824 a_11033_989.n11 a_11033_989.n10 30
R2825 a_11033_989.n9 a_11033_989.n8 24.383
R2826 a_11033_989.n11 a_11033_989.n9 23.684
R2827 a_11033_989.n13 a_11033_989.t3 14.282
R2828 a_11033_989.n13 a_11033_989.t4 14.282
R2829 a_11033_989.t1 a_11033_989.n15 14.282
R2830 a_11033_989.n15 a_11033_989.t0 14.282
R2831 a_11033_989.n15 a_11033_989.n14 12.848
R2832 a_11033_989.n7 a_11033_989.n6 2.947
R2833 a_5101_1050.n5 a_5101_1050.t7 512.525
R2834 a_5101_1050.n3 a_5101_1050.t6 512.525
R2835 a_5101_1050.n5 a_5101_1050.t5 371.139
R2836 a_5101_1050.n3 a_5101_1050.t8 371.139
R2837 a_5101_1050.n4 a_5101_1050.t10 234.562
R2838 a_5101_1050.n6 a_5101_1050.t9 234.204
R2839 a_5101_1050.n6 a_5101_1050.n5 216.178
R2840 a_5101_1050.n4 a_5101_1050.n3 215.819
R2841 a_5101_1050.n8 a_5101_1050.n2 205.605
R2842 a_5101_1050.n10 a_5101_1050.n8 164.008
R2843 a_5101_1050.n7 a_5101_1050.n4 79.488
R2844 a_5101_1050.n8 a_5101_1050.n7 77.314
R2845 a_5101_1050.n2 a_5101_1050.n1 76.002
R2846 a_5101_1050.n7 a_5101_1050.n6 76
R2847 a_5101_1050.n10 a_5101_1050.n9 15.218
R2848 a_5101_1050.n0 a_5101_1050.t4 14.282
R2849 a_5101_1050.n0 a_5101_1050.t2 14.282
R2850 a_5101_1050.n1 a_5101_1050.t0 14.282
R2851 a_5101_1050.n1 a_5101_1050.t1 14.282
R2852 a_5101_1050.n2 a_5101_1050.n0 12.85
R2853 a_5101_1050.n11 a_5101_1050.n10 12.014
R2854 a_5227_411.n1 a_5227_411.t9 480.392
R2855 a_5227_411.n3 a_5227_411.t8 472.359
R2856 a_5227_411.n1 a_5227_411.t12 403.272
R2857 a_5227_411.n3 a_5227_411.t11 384.527
R2858 a_5227_411.n2 a_5227_411.t10 336.586
R2859 a_5227_411.n4 a_5227_411.t7 294.278
R2860 a_5227_411.n10 a_5227_411.n9 265.87
R2861 a_5227_411.n11 a_5227_411.n10 117.354
R2862 a_5227_411.n5 a_5227_411.n2 83.304
R2863 a_5227_411.n5 a_5227_411.n4 80.032
R2864 a_5227_411.n13 a_5227_411.n12 79.232
R2865 a_5227_411.n10 a_5227_411.n5 76
R2866 a_5227_411.n13 a_5227_411.n11 63.152
R2867 a_5227_411.n4 a_5227_411.n3 56.954
R2868 a_5227_411.n2 a_5227_411.n1 45.341
R2869 a_5227_411.n9 a_5227_411.n8 30
R2870 a_5227_411.n7 a_5227_411.n6 24.383
R2871 a_5227_411.n9 a_5227_411.n7 23.684
R2872 a_5227_411.n11 a_5227_411.n0 16.08
R2873 a_5227_411.n14 a_5227_411.n13 16.078
R2874 a_5227_411.n0 a_5227_411.t2 14.282
R2875 a_5227_411.n0 a_5227_411.t3 14.282
R2876 a_5227_411.n12 a_5227_411.t5 14.282
R2877 a_5227_411.n12 a_5227_411.t6 14.282
R2878 a_5227_411.t1 a_5227_411.n14 14.282
R2879 a_5227_411.n14 a_5227_411.t0 14.282
R2880 a_1905_1050.n0 a_1905_1050.t7 480.392
R2881 a_1905_1050.n0 a_1905_1050.t9 403.272
R2882 a_1905_1050.n1 a_1905_1050.t8 230.374
R2883 a_1905_1050.n10 a_1905_1050.n6 223.905
R2884 a_1905_1050.n6 a_1905_1050.n5 159.998
R2885 a_1905_1050.n6 a_1905_1050.n1 153.315
R2886 a_1905_1050.n1 a_1905_1050.n0 151.553
R2887 a_1905_1050.n9 a_1905_1050.n8 79.232
R2888 a_1905_1050.n10 a_1905_1050.n9 63.152
R2889 a_1905_1050.n5 a_1905_1050.n4 30
R2890 a_1905_1050.n3 a_1905_1050.n2 24.383
R2891 a_1905_1050.n5 a_1905_1050.n3 23.684
R2892 a_1905_1050.n9 a_1905_1050.n7 16.08
R2893 a_1905_1050.n11 a_1905_1050.n10 16.078
R2894 a_1905_1050.n7 a_1905_1050.t4 14.282
R2895 a_1905_1050.n7 a_1905_1050.t3 14.282
R2896 a_1905_1050.n8 a_1905_1050.t5 14.282
R2897 a_1905_1050.n8 a_1905_1050.t6 14.282
R2898 a_1905_1050.t1 a_1905_1050.n11 14.282
R2899 a_1905_1050.n11 a_1905_1050.t0 14.282
R2900 a_11673_1050.n2 a_11673_1050.t8 480.392
R2901 a_11673_1050.n2 a_11673_1050.t9 403.272
R2902 a_11673_1050.n3 a_11673_1050.t7 230.374
R2903 a_11673_1050.n9 a_11673_1050.n8 223.905
R2904 a_11673_1050.n8 a_11673_1050.n7 159.998
R2905 a_11673_1050.n8 a_11673_1050.n3 153.315
R2906 a_11673_1050.n3 a_11673_1050.n2 151.553
R2907 a_11673_1050.n11 a_11673_1050.n10 79.231
R2908 a_11673_1050.n10 a_11673_1050.n9 63.152
R2909 a_11673_1050.n7 a_11673_1050.n6 30
R2910 a_11673_1050.n5 a_11673_1050.n4 24.383
R2911 a_11673_1050.n7 a_11673_1050.n5 23.684
R2912 a_11673_1050.n9 a_11673_1050.n1 16.08
R2913 a_11673_1050.n10 a_11673_1050.n0 16.08
R2914 a_11673_1050.n1 a_11673_1050.t3 14.282
R2915 a_11673_1050.n1 a_11673_1050.t2 14.282
R2916 a_11673_1050.n0 a_11673_1050.t6 14.282
R2917 a_11673_1050.n0 a_11673_1050.t5 14.282
R2918 a_11673_1050.n11 a_11673_1050.t0 14.282
R2919 a_11673_1050.t1 a_11673_1050.n11 14.282
R2920 a_15533_1051.n4 a_15533_1051.n3 196.002
R2921 a_15533_1051.n2 a_15533_1051.t5 89.553
R2922 a_15533_1051.n4 a_15533_1051.n0 75.271
R2923 a_15533_1051.n3 a_15533_1051.n2 75.214
R2924 a_15533_1051.n5 a_15533_1051.n4 36.519
R2925 a_15533_1051.n3 a_15533_1051.t2 14.338
R2926 a_15533_1051.n1 a_15533_1051.t4 14.282
R2927 a_15533_1051.n1 a_15533_1051.t3 14.282
R2928 a_15533_1051.n0 a_15533_1051.t7 14.282
R2929 a_15533_1051.n0 a_15533_1051.t6 14.282
R2930 a_15533_1051.t1 a_15533_1051.n5 14.282
R2931 a_15533_1051.n5 a_15533_1051.t0 14.282
R2932 a_15533_1051.n2 a_15533_1051.n1 12.119
R2933 a_2000_210.n9 a_2000_210.n7 82.852
R2934 a_2000_210.n3 a_2000_210.n1 44.628
R2935 a_2000_210.t0 a_2000_210.n9 32.417
R2936 a_2000_210.n7 a_2000_210.n6 27.2
R2937 a_2000_210.n5 a_2000_210.n4 23.498
R2938 a_2000_210.n3 a_2000_210.n2 23.284
R2939 a_2000_210.n7 a_2000_210.n5 22.4
R2940 a_2000_210.t0 a_2000_210.n11 20.241
R2941 a_2000_210.n11 a_2000_210.n10 13.494
R2942 a_2000_210.t0 a_2000_210.n0 8.137
R2943 a_2000_210.t0 a_2000_210.n3 5.727
R2944 a_2000_210.n9 a_2000_210.n8 1.435
R2945 a_10525_103.n4 a_10525_103.n3 19.724
R2946 a_10525_103.t0 a_10525_103.n5 11.595
R2947 a_10525_103.t0 a_10525_103.n4 9.207
R2948 a_10525_103.n2 a_10525_103.n0 8.543
R2949 a_10525_103.t0 a_10525_103.n2 3.034
R2950 a_10525_103.n2 a_10525_103.n1 0.443
R2951 a_10806_210.n12 a_10806_210.n10 82.852
R2952 a_10806_210.n13 a_10806_210.n0 49.6
R2953 a_10806_210.t1 a_10806_210.n2 46.91
R2954 a_10806_210.n7 a_10806_210.n5 34.805
R2955 a_10806_210.n7 a_10806_210.n6 32.622
R2956 a_10806_210.n10 a_10806_210.t1 32.416
R2957 a_10806_210.n12 a_10806_210.n11 27.2
R2958 a_10806_210.n13 a_10806_210.n12 22.4
R2959 a_10806_210.n9 a_10806_210.n7 19.017
R2960 a_10806_210.n2 a_10806_210.n1 17.006
R2961 a_10806_210.n5 a_10806_210.n4 7.5
R2962 a_10806_210.n9 a_10806_210.n8 7.5
R2963 a_10806_210.t1 a_10806_210.n3 7.04
R2964 a_10806_210.n10 a_10806_210.n9 1.435
R2965 a_12470_101.t0 a_12470_101.n1 34.62
R2966 a_12470_101.t0 a_12470_101.n0 8.137
R2967 a_12470_101.t0 a_12470_101.n2 4.69
R2968 D.n5 D.t1 480.392
R2969 D.n2 D.t0 480.392
R2970 D.n0 D.t5 480.392
R2971 D.n5 D.t4 403.272
R2972 D.n2 D.t6 403.272
R2973 D.n0 D.t8 403.272
R2974 D.n6 D.n5 204.659
R2975 D.n3 D.n2 204.659
R2976 D.n1 D.n0 204.659
R2977 D.n6 D.t2 183.422
R2978 D.n3 D.t7 183.422
R2979 D.n1 D.t3 183.422
R2980 D.n4 D.n1 93.91
R2981 D.n4 D.n3 76
R2982 D.n7 D.n6 76
R2983 D.n7 D.n4 17.91
R2984 D.n7 D 0.046
R2985 a_217_1050.n2 a_217_1050.t7 512.525
R2986 a_217_1050.n0 a_217_1050.t10 512.525
R2987 a_217_1050.n2 a_217_1050.t9 371.139
R2988 a_217_1050.n0 a_217_1050.t6 371.139
R2989 a_217_1050.n1 a_217_1050.t8 234.562
R2990 a_217_1050.n3 a_217_1050.t5 234.204
R2991 a_217_1050.n3 a_217_1050.n2 216.178
R2992 a_217_1050.n1 a_217_1050.n0 215.819
R2993 a_217_1050.n11 a_217_1050.n9 205.605
R2994 a_217_1050.n9 a_217_1050.n8 157.486
R2995 a_217_1050.n4 a_217_1050.n1 79.488
R2996 a_217_1050.n9 a_217_1050.n4 77.314
R2997 a_217_1050.n11 a_217_1050.n10 76.002
R2998 a_217_1050.n4 a_217_1050.n3 76
R2999 a_217_1050.n8 a_217_1050.n7 30
R3000 a_217_1050.n6 a_217_1050.n5 24.383
R3001 a_217_1050.n8 a_217_1050.n6 23.684
R3002 a_217_1050.n10 a_217_1050.t4 14.282
R3003 a_217_1050.n10 a_217_1050.t3 14.282
R3004 a_217_1050.t1 a_217_1050.n12 14.282
R3005 a_217_1050.n12 a_217_1050.t0 14.282
R3006 a_217_1050.n12 a_217_1050.n11 12.848
R3007 a_15430_101.t0 a_15430_101.n0 34.602
R3008 a_15430_101.t0 a_15430_101.n1 2.138
R3009 a_10111_411.n2 a_10111_411.t12 480.392
R3010 a_10111_411.n4 a_10111_411.t9 472.359
R3011 a_10111_411.n2 a_10111_411.t8 403.272
R3012 a_10111_411.n4 a_10111_411.t7 384.527
R3013 a_10111_411.n3 a_10111_411.t11 336.586
R3014 a_10111_411.n5 a_10111_411.t10 294.278
R3015 a_10111_411.n10 a_10111_411.n9 281.393
R3016 a_10111_411.n11 a_10111_411.n10 117.354
R3017 a_10111_411.n6 a_10111_411.n3 83.304
R3018 a_10111_411.n6 a_10111_411.n5 80.032
R3019 a_10111_411.n13 a_10111_411.n12 79.231
R3020 a_10111_411.n10 a_10111_411.n6 76
R3021 a_10111_411.n12 a_10111_411.n11 63.152
R3022 a_10111_411.n5 a_10111_411.n4 56.954
R3023 a_10111_411.n3 a_10111_411.n2 45.341
R3024 a_10111_411.n9 a_10111_411.n8 22.578
R3025 a_10111_411.n11 a_10111_411.n1 16.08
R3026 a_10111_411.n12 a_10111_411.n0 16.08
R3027 a_10111_411.n1 a_10111_411.t5 14.282
R3028 a_10111_411.n1 a_10111_411.t4 14.282
R3029 a_10111_411.n0 a_10111_411.t2 14.282
R3030 a_10111_411.n0 a_10111_411.t3 14.282
R3031 a_10111_411.n13 a_10111_411.t0 14.282
R3032 a_10111_411.t1 a_10111_411.n13 14.282
R3033 a_10111_411.n9 a_10111_411.n7 8.58
R3034 a_6789_1050.n0 a_6789_1050.t8 480.392
R3035 a_6789_1050.n0 a_6789_1050.t7 403.272
R3036 a_6789_1050.n1 a_6789_1050.t9 230.374
R3037 a_6789_1050.n7 a_6789_1050.n3 223.905
R3038 a_6789_1050.n3 a_6789_1050.n2 181.737
R3039 a_6789_1050.n3 a_6789_1050.n1 153.315
R3040 a_6789_1050.n1 a_6789_1050.n0 151.553
R3041 a_6789_1050.n6 a_6789_1050.n5 79.232
R3042 a_6789_1050.n7 a_6789_1050.n6 63.152
R3043 a_6789_1050.n6 a_6789_1050.n4 16.08
R3044 a_6789_1050.n8 a_6789_1050.n7 16.078
R3045 a_6789_1050.n4 a_6789_1050.t6 14.282
R3046 a_6789_1050.n4 a_6789_1050.t5 14.282
R3047 a_6789_1050.n5 a_6789_1050.t4 14.282
R3048 a_6789_1050.n5 a_6789_1050.t3 14.282
R3049 a_6789_1050.n8 a_6789_1050.t0 14.282
R3050 a_6789_1050.t1 a_6789_1050.n8 14.282
R3051 a_1038_210.n10 a_1038_210.n8 82.852
R3052 a_1038_210.n7 a_1038_210.n6 32.833
R3053 a_1038_210.n8 a_1038_210.t1 32.416
R3054 a_1038_210.n10 a_1038_210.n9 27.2
R3055 a_1038_210.n11 a_1038_210.n0 23.498
R3056 a_1038_210.n3 a_1038_210.n2 23.284
R3057 a_1038_210.n11 a_1038_210.n10 22.4
R3058 a_1038_210.n7 a_1038_210.n4 19.017
R3059 a_1038_210.n6 a_1038_210.n5 13.494
R3060 a_1038_210.t1 a_1038_210.n1 7.04
R3061 a_1038_210.t1 a_1038_210.n3 5.727
R3062 a_1038_210.n8 a_1038_210.n7 1.435
R3063 a_14062_210.n9 a_14062_210.n7 82.852
R3064 a_14062_210.n3 a_14062_210.n1 44.628
R3065 a_14062_210.t0 a_14062_210.n9 32.417
R3066 a_14062_210.n7 a_14062_210.n6 27.2
R3067 a_14062_210.n5 a_14062_210.n4 23.498
R3068 a_14062_210.n3 a_14062_210.n2 23.284
R3069 a_14062_210.n7 a_14062_210.n5 22.4
R3070 a_14062_210.t0 a_14062_210.n11 20.241
R3071 a_14062_210.n11 a_14062_210.n10 13.494
R3072 a_14062_210.t0 a_14062_210.n0 8.137
R3073 a_14062_210.t0 a_14062_210.n3 5.727
R3074 a_14062_210.n9 a_14062_210.n8 1.435
R3075 a_11768_210.n8 a_11768_210.n6 96.467
R3076 a_11768_210.n3 a_11768_210.n1 44.628
R3077 a_11768_210.t0 a_11768_210.n8 32.417
R3078 a_11768_210.n3 a_11768_210.n2 23.284
R3079 a_11768_210.n6 a_11768_210.n5 22.349
R3080 a_11768_210.t0 a_11768_210.n10 20.241
R3081 a_11768_210.n10 a_11768_210.n9 13.494
R3082 a_11768_210.n6 a_11768_210.n4 8.443
R3083 a_11768_210.t0 a_11768_210.n0 8.137
R3084 a_11768_210.t0 a_11768_210.n3 5.727
R3085 a_11768_210.n8 a_11768_210.n7 1.435
R3086 a_7586_101.t0 a_7586_101.n1 34.62
R3087 a_7586_101.t0 a_7586_101.n0 8.137
R3088 a_7586_101.t0 a_7586_101.n2 4.69
R3089 a_757_103.n1 a_757_103.n0 25.576
R3090 a_757_103.n3 a_757_103.n2 9.111
R3091 a_757_103.n7 a_757_103.n6 2.455
R3092 a_757_103.n5 a_757_103.n3 1.964
R3093 a_757_103.n5 a_757_103.n4 1.964
R3094 a_757_103.t0 a_757_103.n1 1.871
R3095 a_757_103.n7 a_757_103.n5 0.636
R3096 a_757_103.t0 a_757_103.n7 0.246
R3097 a_5922_210.n10 a_5922_210.n8 82.852
R3098 a_5922_210.n7 a_5922_210.n6 32.833
R3099 a_5922_210.n8 a_5922_210.t1 32.416
R3100 a_5922_210.n10 a_5922_210.n9 27.2
R3101 a_5922_210.n11 a_5922_210.n0 23.498
R3102 a_5922_210.n3 a_5922_210.n2 23.284
R3103 a_5922_210.n11 a_5922_210.n10 22.4
R3104 a_5922_210.n7 a_5922_210.n4 19.017
R3105 a_5922_210.n6 a_5922_210.n5 13.494
R3106 a_5922_210.t1 a_5922_210.n1 7.04
R3107 a_5922_210.t1 a_5922_210.n3 5.727
R3108 a_5922_210.n8 a_5922_210.n7 1.435
R3109 a_16096_101.t0 a_16096_101.n1 34.62
R3110 a_16096_101.t0 a_16096_101.n0 8.137
R3111 a_16096_101.t0 a_16096_101.n2 4.69
R3112 a_4996_101.t0 a_4996_101.n1 34.62
R3113 a_4996_101.t0 a_4996_101.n0 8.137
R3114 a_4996_101.t0 a_4996_101.n2 4.69
R3115 a_112_101.t0 a_112_101.n1 34.62
R3116 a_112_101.t0 a_112_101.n0 8.137
R3117 a_112_101.t0 a_112_101.n2 4.69
R3118 a_8897_103.n4 a_8897_103.n3 19.724
R3119 a_8897_103.t0 a_8897_103.n5 11.595
R3120 a_8897_103.t0 a_8897_103.n4 9.207
R3121 a_8897_103.n2 a_8897_103.n0 8.543
R3122 a_8897_103.t0 a_8897_103.n2 3.034
R3123 a_8897_103.n2 a_8897_103.n1 0.443
R3124 a_9178_210.n8 a_9178_210.n6 96.467
R3125 a_9178_210.n3 a_9178_210.n1 44.628
R3126 a_9178_210.t0 a_9178_210.n8 32.417
R3127 a_9178_210.n3 a_9178_210.n2 23.284
R3128 a_9178_210.n6 a_9178_210.n5 22.349
R3129 a_9178_210.t0 a_9178_210.n10 20.241
R3130 a_9178_210.n10 a_9178_210.n9 13.494
R3131 a_9178_210.n6 a_9178_210.n4 8.443
R3132 a_9178_210.t0 a_9178_210.n0 8.137
R3133 a_9178_210.t0 a_9178_210.n3 5.727
R3134 a_9178_210.n8 a_9178_210.n7 1.435
R3135 a_3368_101.t0 a_3368_101.n1 34.62
R3136 a_3368_101.t0 a_3368_101.n0 8.137
R3137 a_3368_101.t0 a_3368_101.n2 4.69
R3138 a_9880_101.n12 a_9880_101.n11 26.811
R3139 a_9880_101.n6 a_9880_101.n5 24.977
R3140 a_9880_101.n2 a_9880_101.n1 24.877
R3141 a_9880_101.t0 a_9880_101.n2 12.677
R3142 a_9880_101.t0 a_9880_101.n3 11.595
R3143 a_9880_101.t1 a_9880_101.n8 8.137
R3144 a_9880_101.t0 a_9880_101.n4 7.273
R3145 a_9880_101.t0 a_9880_101.n0 6.109
R3146 a_9880_101.t1 a_9880_101.n7 4.864
R3147 a_9880_101.t0 a_9880_101.n12 2.074
R3148 a_9880_101.n7 a_9880_101.n6 1.13
R3149 a_9880_101.n12 a_9880_101.t1 0.937
R3150 a_9880_101.t1 a_9880_101.n10 0.804
R3151 a_9880_101.n10 a_9880_101.n9 0.136
R3152 a_1719_103.n1 a_1719_103.n0 25.576
R3153 a_1719_103.n3 a_1719_103.n2 9.111
R3154 a_1719_103.n7 a_1719_103.n6 2.455
R3155 a_1719_103.n5 a_1719_103.n3 1.964
R3156 a_1719_103.n5 a_1719_103.n4 1.964
R3157 a_1719_103.t0 a_1719_103.n1 1.871
R3158 a_1719_103.n7 a_1719_103.n5 0.636
R3159 a_1719_103.t0 a_1719_103.n7 0.246
R3160 a_13781_103.n5 a_13781_103.n4 19.724
R3161 a_13781_103.t0 a_13781_103.n3 11.595
R3162 a_13781_103.t0 a_13781_103.n5 9.207
R3163 a_13781_103.n2 a_13781_103.n1 2.455
R3164 a_13781_103.n2 a_13781_103.n0 1.32
R3165 a_13781_103.t0 a_13781_103.n2 0.246
R3166 a_2702_101.t0 a_2702_101.n1 34.62
R3167 a_2702_101.t0 a_2702_101.n0 8.137
R3168 a_2702_101.t0 a_2702_101.n2 4.69
R3169 a_8252_101.n12 a_8252_101.n11 26.811
R3170 a_8252_101.n6 a_8252_101.n5 24.977
R3171 a_8252_101.n2 a_8252_101.n1 24.877
R3172 a_8252_101.t0 a_8252_101.n2 12.677
R3173 a_8252_101.t0 a_8252_101.n3 11.595
R3174 a_8252_101.t1 a_8252_101.n8 8.137
R3175 a_8252_101.t0 a_8252_101.n4 7.273
R3176 a_8252_101.t0 a_8252_101.n0 6.109
R3177 a_8252_101.t1 a_8252_101.n7 4.864
R3178 a_8252_101.t0 a_8252_101.n12 2.074
R3179 a_8252_101.n7 a_8252_101.n6 1.13
R3180 a_8252_101.n12 a_8252_101.t1 0.937
R3181 a_8252_101.t1 a_8252_101.n10 0.804
R3182 a_8252_101.n10 a_8252_101.n9 0.136
R3183 a_5641_103.n1 a_5641_103.n0 25.576
R3184 a_5641_103.n3 a_5641_103.n2 9.111
R3185 a_5641_103.n7 a_5641_103.n6 2.455
R3186 a_5641_103.n5 a_5641_103.n3 1.964
R3187 a_5641_103.n5 a_5641_103.n4 1.964
R3188 a_5641_103.t0 a_5641_103.n1 1.871
R3189 a_5641_103.n7 a_5641_103.n5 0.636
R3190 a_5641_103.t0 a_5641_103.n7 0.246
R3191 a_14764_101.n1 a_14764_101.n0 32.249
R3192 a_14764_101.t0 a_14764_101.n5 7.911
R3193 a_14764_101.n4 a_14764_101.n2 4.032
R3194 a_14764_101.n4 a_14764_101.n3 3.644
R3195 a_14764_101.t0 a_14764_101.n1 2.534
R3196 a_14764_101.t0 a_14764_101.n4 1.099
C7 SN GND 8.21fF
C8 VDD GND 62.21fF
C9 a_14764_101.n0 GND 0.11fF
C10 a_14764_101.n1 GND 0.09fF
C11 a_14764_101.n2 GND 0.08fF
C12 a_14764_101.n3 GND 0.02fF
C13 a_14764_101.n4 GND 0.01fF
C14 a_14764_101.n5 GND 0.06fF
C15 a_5641_103.n0 GND 0.09fF
C16 a_5641_103.n1 GND 0.10fF
C17 a_5641_103.n2 GND 0.05fF
C18 a_5641_103.n3 GND 0.03fF
C19 a_5641_103.n4 GND 0.04fF
C20 a_5641_103.n5 GND 0.03fF
C21 a_5641_103.n6 GND 0.04fF
C22 a_8252_101.n0 GND 0.02fF
C23 a_8252_101.n1 GND 0.10fF
C24 a_8252_101.n2 GND 0.06fF
C25 a_8252_101.n3 GND 0.06fF
C26 a_8252_101.n4 GND 0.00fF
C27 a_8252_101.n5 GND 0.04fF
C28 a_8252_101.n6 GND 0.05fF
C29 a_8252_101.n7 GND 0.02fF
C30 a_8252_101.n8 GND 0.05fF
C31 a_8252_101.n9 GND 0.08fF
C32 a_8252_101.n10 GND 0.17fF
C33 a_8252_101.t1 GND 0.23fF
C34 a_8252_101.n11 GND 0.09fF
C35 a_8252_101.n12 GND 0.00fF
C36 a_2702_101.n0 GND 0.05fF
C37 a_2702_101.n1 GND 0.12fF
C38 a_2702_101.n2 GND 0.04fF
C39 a_13781_103.n0 GND 0.10fF
C40 a_13781_103.n1 GND 0.04fF
C41 a_13781_103.n2 GND 0.03fF
C42 a_13781_103.n3 GND 0.07fF
C43 a_13781_103.n4 GND 0.08fF
C44 a_13781_103.n5 GND 0.06fF
C45 a_1719_103.n0 GND 0.09fF
C46 a_1719_103.n1 GND 0.10fF
C47 a_1719_103.n2 GND 0.05fF
C48 a_1719_103.n3 GND 0.03fF
C49 a_1719_103.n4 GND 0.04fF
C50 a_1719_103.n5 GND 0.03fF
C51 a_1719_103.n6 GND 0.04fF
C52 a_9880_101.n0 GND 0.02fF
C53 a_9880_101.n1 GND 0.10fF
C54 a_9880_101.n2 GND 0.06fF
C55 a_9880_101.n3 GND 0.06fF
C56 a_9880_101.n4 GND 0.00fF
C57 a_9880_101.n5 GND 0.04fF
C58 a_9880_101.n6 GND 0.05fF
C59 a_9880_101.n7 GND 0.02fF
C60 a_9880_101.n8 GND 0.05fF
C61 a_9880_101.n9 GND 0.08fF
C62 a_9880_101.n10 GND 0.17fF
C63 a_9880_101.t1 GND 0.23fF
C64 a_9880_101.n11 GND 0.09fF
C65 a_9880_101.n12 GND 0.00fF
C66 a_3368_101.n0 GND 0.05fF
C67 a_3368_101.n1 GND 0.12fF
C68 a_3368_101.n2 GND 0.04fF
C69 a_9178_210.n0 GND 0.07fF
C70 a_9178_210.n1 GND 0.09fF
C71 a_9178_210.n2 GND 0.13fF
C72 a_9178_210.n3 GND 0.11fF
C73 a_9178_210.n4 GND 0.02fF
C74 a_9178_210.n5 GND 0.03fF
C75 a_9178_210.n6 GND 0.06fF
C76 a_9178_210.n7 GND 0.03fF
C77 a_9178_210.n8 GND 0.12fF
C78 a_9178_210.n9 GND 0.06fF
C79 a_9178_210.n10 GND 0.01fF
C80 a_9178_210.t0 GND 0.33fF
C81 a_8897_103.n0 GND 0.20fF
C82 a_8897_103.n1 GND 0.04fF
C83 a_8897_103.n2 GND 0.01fF
C84 a_8897_103.n3 GND 0.08fF
C85 a_8897_103.n4 GND 0.06fF
C86 a_8897_103.n5 GND 0.07fF
C87 a_112_101.n0 GND 0.05fF
C88 a_112_101.n1 GND 0.12fF
C89 a_112_101.n2 GND 0.04fF
C90 a_4996_101.n0 GND 0.05fF
C91 a_4996_101.n1 GND 0.12fF
C92 a_4996_101.n2 GND 0.04fF
C93 a_16096_101.n0 GND 0.06fF
C94 a_16096_101.n1 GND 0.14fF
C95 a_16096_101.n2 GND 0.04fF
C96 a_5922_210.n0 GND 0.02fF
C97 a_5922_210.n1 GND 0.09fF
C98 a_5922_210.n2 GND 0.13fF
C99 a_5922_210.n3 GND 0.11fF
C100 a_5922_210.t1 GND 0.30fF
C101 a_5922_210.n4 GND 0.09fF
C102 a_5922_210.n5 GND 0.06fF
C103 a_5922_210.n6 GND 0.01fF
C104 a_5922_210.n7 GND 0.03fF
C105 a_5922_210.n8 GND 0.11fF
C106 a_5922_210.n9 GND 0.02fF
C107 a_5922_210.n10 GND 0.05fF
C108 a_5922_210.n11 GND 0.03fF
C109 a_757_103.n0 GND 0.09fF
C110 a_757_103.n1 GND 0.10fF
C111 a_757_103.n2 GND 0.05fF
C112 a_757_103.n3 GND 0.03fF
C113 a_757_103.n4 GND 0.04fF
C114 a_757_103.n5 GND 0.03fF
C115 a_757_103.n6 GND 0.04fF
C116 a_7586_101.n0 GND 0.05fF
C117 a_7586_101.n1 GND 0.12fF
C118 a_7586_101.n2 GND 0.04fF
C119 a_11768_210.n0 GND 0.07fF
C120 a_11768_210.n1 GND 0.09fF
C121 a_11768_210.n2 GND 0.13fF
C122 a_11768_210.n3 GND 0.11fF
C123 a_11768_210.n4 GND 0.02fF
C124 a_11768_210.n5 GND 0.03fF
C125 a_11768_210.n6 GND 0.06fF
C126 a_11768_210.n7 GND 0.03fF
C127 a_11768_210.n8 GND 0.12fF
C128 a_11768_210.n9 GND 0.06fF
C129 a_11768_210.n10 GND 0.01fF
C130 a_11768_210.t0 GND 0.33fF
C131 a_14062_210.n0 GND 0.07fF
C132 a_14062_210.n1 GND 0.09fF
C133 a_14062_210.n2 GND 0.13fF
C134 a_14062_210.n3 GND 0.11fF
C135 a_14062_210.n4 GND 0.02fF
C136 a_14062_210.n5 GND 0.03fF
C137 a_14062_210.n6 GND 0.02fF
C138 a_14062_210.n7 GND 0.05fF
C139 a_14062_210.n8 GND 0.03fF
C140 a_14062_210.n9 GND 0.11fF
C141 a_14062_210.n10 GND 0.06fF
C142 a_14062_210.n11 GND 0.01fF
C143 a_14062_210.t0 GND 0.33fF
C144 a_1038_210.n0 GND 0.02fF
C145 a_1038_210.n1 GND 0.09fF
C146 a_1038_210.n2 GND 0.13fF
C147 a_1038_210.n3 GND 0.11fF
C148 a_1038_210.t1 GND 0.30fF
C149 a_1038_210.n4 GND 0.09fF
C150 a_1038_210.n5 GND 0.06fF
C151 a_1038_210.n6 GND 0.01fF
C152 a_1038_210.n7 GND 0.03fF
C153 a_1038_210.n8 GND 0.11fF
C154 a_1038_210.n9 GND 0.02fF
C155 a_1038_210.n10 GND 0.05fF
C156 a_1038_210.n11 GND 0.03fF
C157 a_6789_1050.n0 GND 0.45fF
C158 a_6789_1050.n1 GND 0.58fF
C159 a_6789_1050.n2 GND 0.35fF
C160 a_6789_1050.n3 GND 0.68fF
C161 a_6789_1050.n4 GND 0.55fF
C162 a_6789_1050.n5 GND 0.65fF
C163 a_6789_1050.n6 GND 0.21fF
C164 a_6789_1050.n7 GND 0.38fF
C165 a_6789_1050.n8 GND 0.55fF
C166 a_10111_411.n0 GND 0.86fF
C167 a_10111_411.n1 GND 0.86fF
C168 a_10111_411.n2 GND 0.50fF
C169 a_10111_411.n3 GND 0.76fF
C170 a_10111_411.n4 GND 0.44fF
C171 a_10111_411.t10 GND 0.94fF
C172 a_10111_411.n5 GND 0.65fF
C173 a_10111_411.n6 GND 4.01fF
C174 a_10111_411.n7 GND 0.07fF
C175 a_10111_411.n8 GND 0.09fF
C176 a_10111_411.n9 GND 0.60fF
C177 a_10111_411.n10 GND 0.76fF
C178 a_10111_411.n11 GND 0.39fF
C179 a_10111_411.n12 GND 0.32fF
C180 a_10111_411.n13 GND 1.01fF
C181 a_15430_101.n0 GND 0.13fF
C182 a_15430_101.n1 GND 0.13fF
C183 a_217_1050.n0 GND 0.35fF
C184 a_217_1050.n1 GND 0.42fF
C185 a_217_1050.n2 GND 0.35fF
C186 a_217_1050.n3 GND 0.41fF
C187 a_217_1050.n4 GND 0.99fF
C188 a_217_1050.n5 GND 0.04fF
C189 a_217_1050.n6 GND 0.05fF
C190 a_217_1050.n7 GND 0.03fF
C191 a_217_1050.n8 GND 0.21fF
C192 a_217_1050.n9 GND 0.38fF
C193 a_217_1050.n10 GND 0.55fF
C194 a_217_1050.n11 GND 0.32fF
C195 a_217_1050.n12 GND 0.46fF
C196 a_12470_101.n0 GND 0.05fF
C197 a_12470_101.n1 GND 0.12fF
C198 a_12470_101.n2 GND 0.04fF
C199 a_10806_210.n0 GND 0.02fF
C200 a_10806_210.n1 GND 0.07fF
C201 a_10806_210.n2 GND 0.13fF
C202 a_10806_210.n3 GND 0.09fF
C203 a_10806_210.t1 GND 0.25fF
C204 a_10806_210.n4 GND 0.05fF
C205 a_10806_210.n5 GND 0.06fF
C206 a_10806_210.n6 GND 0.07fF
C207 a_10806_210.n7 GND 0.07fF
C208 a_10806_210.n8 GND 0.03fF
C209 a_10806_210.n9 GND 0.01fF
C210 a_10806_210.n10 GND 0.11fF
C211 a_10806_210.n11 GND 0.02fF
C212 a_10806_210.n12 GND 0.05fF
C213 a_10806_210.n13 GND 0.02fF
C214 a_10525_103.n0 GND 0.20fF
C215 a_10525_103.n1 GND 0.04fF
C216 a_10525_103.n2 GND 0.01fF
C217 a_10525_103.n3 GND 0.08fF
C218 a_10525_103.n4 GND 0.06fF
C219 a_10525_103.n5 GND 0.07fF
C220 a_2000_210.n0 GND 0.07fF
C221 a_2000_210.n1 GND 0.09fF
C222 a_2000_210.n2 GND 0.13fF
C223 a_2000_210.n3 GND 0.11fF
C224 a_2000_210.n4 GND 0.02fF
C225 a_2000_210.n5 GND 0.03fF
C226 a_2000_210.n6 GND 0.02fF
C227 a_2000_210.n7 GND 0.05fF
C228 a_2000_210.n8 GND 0.03fF
C229 a_2000_210.n9 GND 0.11fF
C230 a_2000_210.n10 GND 0.06fF
C231 a_2000_210.n11 GND 0.01fF
C232 a_2000_210.t0 GND 0.33fF
C233 a_15533_1051.n0 GND 0.36fF
C234 a_15533_1051.n1 GND 0.29fF
C235 a_15533_1051.n2 GND 0.20fF
C236 a_15533_1051.n3 GND 0.57fF
C237 a_15533_1051.n4 GND 0.25fF
C238 a_15533_1051.n5 GND 0.28fF
C239 a_11673_1050.n0 GND 0.55fF
C240 a_11673_1050.n1 GND 0.55fF
C241 a_11673_1050.n2 GND 0.45fF
C242 a_11673_1050.n3 GND 0.57fF
C243 a_11673_1050.n4 GND 0.04fF
C244 a_11673_1050.n5 GND 0.06fF
C245 a_11673_1050.n6 GND 0.04fF
C246 a_11673_1050.n7 GND 0.24fF
C247 a_11673_1050.n8 GND 0.65fF
C248 a_11673_1050.n9 GND 0.38fF
C249 a_11673_1050.n10 GND 0.20fF
C250 a_11673_1050.n11 GND 0.65fF
C251 a_1905_1050.n0 GND 0.41fF
C252 a_1905_1050.n1 GND 0.53fF
C253 a_1905_1050.n2 GND 0.04fF
C254 a_1905_1050.n3 GND 0.05fF
C255 a_1905_1050.n4 GND 0.03fF
C256 a_1905_1050.n5 GND 0.22fF
C257 a_1905_1050.n6 GND 0.59fF
C258 a_1905_1050.n7 GND 0.50fF
C259 a_1905_1050.n8 GND 0.59fF
C260 a_1905_1050.n9 GND 0.19fF
C261 a_1905_1050.n10 GND 0.35fF
C262 a_1905_1050.n11 GND 0.50fF
C263 a_5227_411.n0 GND 0.83fF
C264 a_5227_411.n1 GND 0.48fF
C265 a_5227_411.n2 GND 0.74fF
C266 a_5227_411.n3 GND 0.43fF
C267 a_5227_411.t7 GND 0.91fF
C268 a_5227_411.n4 GND 0.63fF
C269 a_5227_411.n5 GND 3.88fF
C270 a_5227_411.n6 GND 0.06fF
C271 a_5227_411.n7 GND 0.08fF
C272 a_5227_411.n8 GND 0.05fF
C273 a_5227_411.n9 GND 0.56fF
C274 a_5227_411.n10 GND 0.70fF
C275 a_5227_411.n11 GND 0.38fF
C276 a_5227_411.n12 GND 0.98fF
C277 a_5227_411.n13 GND 0.31fF
C278 a_5227_411.n14 GND 0.83fF
C279 a_5101_1050.n0 GND 0.71fF
C280 a_5101_1050.n1 GND 0.84fF
C281 a_5101_1050.n2 GND 0.49fF
C282 a_5101_1050.n3 GND 0.54fF
C283 a_5101_1050.n4 GND 0.65fF
C284 a_5101_1050.n5 GND 0.54fF
C285 a_5101_1050.n6 GND 0.63fF
C286 a_5101_1050.n7 GND 1.52fF
C287 a_5101_1050.n8 GND 0.59fF
C288 a_5101_1050.n9 GND 0.11fF
C289 a_5101_1050.n10 GND 0.30fF
C290 a_5101_1050.n11 GND 0.06fF
C291 a_11033_989.n0 GND 0.59fF
C292 a_11033_989.t6 GND 0.97fF
C293 a_11033_989.n1 GND 0.71fF
C294 a_11033_989.n2 GND 0.59fF
C295 a_11033_989.t12 GND 0.96fF
C296 a_11033_989.n3 GND 0.64fF
C297 a_11033_989.n4 GND 0.59fF
C298 a_11033_989.t10 GND 0.97fF
C299 a_11033_989.n5 GND 0.67fF
C300 a_11033_989.n6 GND 1.96fF
C301 a_11033_989.n7 GND 2.64fF
C302 a_11033_989.n8 GND 0.07fF
C303 a_11033_989.n9 GND 0.09fF
C304 a_11033_989.n10 GND 0.06fF
C305 a_11033_989.n11 GND 0.57fF
C306 a_11033_989.n12 GND 0.73fF
C307 a_11033_989.n13 GND 1.08fF
C308 a_11033_989.n14 GND 0.47fF
C309 a_11033_989.n15 GND 0.91fF
C310 a_343_411.n0 GND 0.72fF
C311 a_343_411.n1 GND 0.42fF
C312 a_343_411.n2 GND 0.64fF
C313 a_343_411.n3 GND 0.37fF
C314 a_343_411.t11 GND 0.79fF
C315 a_343_411.n4 GND 0.55fF
C316 a_343_411.n5 GND 3.36fF
C317 a_343_411.n6 GND 0.05fF
C318 a_343_411.n7 GND 0.07fF
C319 a_343_411.n8 GND 0.05fF
C320 a_343_411.n9 GND 0.49fF
C321 a_343_411.n10 GND 0.61fF
C322 a_343_411.n11 GND 0.33fF
C323 a_343_411.n12 GND 0.85fF
C324 a_343_411.n13 GND 0.27fF
C325 a_343_411.n14 GND 0.72fF
C326 a_1265_989.n0 GND 0.45fF
C327 a_1265_989.t13 GND 0.73fF
C328 a_1265_989.n1 GND 0.54fF
C329 a_1265_989.n2 GND 0.45fF
C330 a_1265_989.t6 GND 0.73fF
C331 a_1265_989.n3 GND 0.48fF
C332 a_1265_989.n4 GND 0.45fF
C333 a_1265_989.t8 GND 0.73fF
C334 a_1265_989.n5 GND 0.51fF
C335 a_1265_989.n6 GND 1.49fF
C336 a_1265_989.n7 GND 2.01fF
C337 a_1265_989.n8 GND 0.05fF
C338 a_1265_989.n9 GND 0.07fF
C339 a_1265_989.n10 GND 0.04fF
C340 a_1265_989.n11 GND 0.43fF
C341 a_1265_989.n12 GND 0.55fF
C342 a_1265_989.n13 GND 0.82fF
C343 a_1265_989.n14 GND 0.36fF
C344 a_1265_989.n15 GND 0.69fF
C345 Q.n0 GND 0.75fF
C346 Q.n1 GND 0.45fF
C347 Q.n2 GND 0.51fF
C348 Q.n3 GND 0.01fF
C349 a_15044_209.n0 GND 0.03fF
C350 a_15044_209.n1 GND 0.37fF
C351 a_15044_209.n2 GND 0.45fF
C352 a_15044_209.n3 GND 0.23fF
C353 a_15044_209.n4 GND 0.26fF
C354 a_15044_209.n5 GND 0.48fF
C355 a_15044_209.n6 GND 0.45fF
C356 a_15044_209.n7 GND 0.05fF
C357 a_15044_209.n8 GND 0.03fF
C358 a_15044_209.n9 GND 0.07fF
C359 a_15044_209.n10 GND 0.25fF
C360 a_15044_209.n11 GND 0.03fF
C361 a_15044_209.n12 GND 0.04fF
C362 a_15044_209.n13 GND 0.03fF
C363 a_15044_209.n14 GND 0.09fF
C364 a_15044_209.n15 GND 0.96fF
C365 a_15044_209.n16 GND 0.03fF
C366 a_15044_209.n17 GND 0.08fF
C367 a_15044_209.n18 GND 0.04fF
C368 a_11487_103.n0 GND 0.20fF
C369 a_11487_103.n1 GND 0.04fF
C370 a_11487_103.n2 GND 0.01fF
C371 a_11487_103.n3 GND 0.03fF
C372 a_11487_103.n4 GND 0.05fF
C373 a_11487_103.n5 GND 0.09fF
C374 a_11487_103.n6 GND 0.07fF
C375 a_9985_1050.n0 GND 0.71fF
C376 a_9985_1050.n1 GND 0.83fF
C377 a_9985_1050.n2 GND 0.49fF
C378 a_9985_1050.n3 GND 0.53fF
C379 a_9985_1050.n4 GND 0.65fF
C380 a_9985_1050.n5 GND 0.53fF
C381 a_9985_1050.n6 GND 0.62fF
C382 a_9985_1050.n7 GND 1.51fF
C383 a_9985_1050.n8 GND 0.58fF
C384 a_9985_1050.n9 GND 0.11fF
C385 a_9985_1050.n10 GND 0.30fF
C386 a_9985_1050.n11 GND 0.06fF
C387 a_4294_210.n0 GND 0.07fF
C388 a_4294_210.n1 GND 0.09fF
C389 a_4294_210.n2 GND 0.13fF
C390 a_4294_210.n3 GND 0.11fF
C391 a_4294_210.n4 GND 0.02fF
C392 a_4294_210.n5 GND 0.03fF
C393 a_4294_210.n6 GND 0.06fF
C394 a_4294_210.n7 GND 0.03fF
C395 a_4294_210.n8 GND 0.12fF
C396 a_4294_210.n9 GND 0.06fF
C397 a_4294_210.n10 GND 0.01fF
C398 a_4294_210.t0 GND 0.33fF
C399 a_4013_103.n0 GND 0.20fF
C400 a_4013_103.n1 GND 0.04fF
C401 a_4013_103.n2 GND 0.01fF
C402 a_4013_103.n3 GND 0.03fF
C403 a_4013_103.n4 GND 0.05fF
C404 a_4013_103.n5 GND 0.09fF
C405 a_4013_103.n6 GND 0.07fF
C406 a_13241_1050.n0 GND 0.24fF
C407 a_13241_1050.n1 GND 0.70fF
C408 a_13241_1050.n2 GND 0.48fF
C409 a_13241_1050.n3 GND 0.59fF
C410 a_13241_1050.n4 GND 0.62fF
C411 a_13241_1050.n5 GND 0.21fF
C412 a_13241_1050.n6 GND 0.52fF
C413 a_13136_101.n0 GND 0.05fF
C414 a_13136_101.n1 GND 0.02fF
C415 a_13136_101.n2 GND 0.12fF
C416 a_13136_101.n3 GND 0.04fF
C417 a_13136_101.n4 GND 0.17fF
C418 a_13367_411.n0 GND 0.58fF
C419 a_13367_411.n1 GND 0.33fF
C420 a_13367_411.t9 GND 0.63fF
C421 a_13367_411.n2 GND 0.47fF
C422 a_13367_411.n3 GND 0.30fF
C423 a_13367_411.t13 GND 0.63fF
C424 a_13367_411.n4 GND 0.41fF
C425 a_13367_411.n5 GND 1.40fF
C426 a_13367_411.n6 GND 0.30fF
C427 a_13367_411.t7 GND 0.63fF
C428 a_13367_411.n7 GND 0.44fF
C429 a_13367_411.n8 GND 1.22fF
C430 a_13367_411.n9 GND 0.05fF
C431 a_13367_411.n10 GND 0.06fF
C432 a_13367_411.n11 GND 0.40fF
C433 a_13367_411.n12 GND 0.51fF
C434 a_13367_411.n13 GND 0.26fF
C435 a_13367_411.n14 GND 0.68fF
C436 a_13367_411.n15 GND 0.21fF
C437 a_13367_411.n16 GND 0.58fF
C438 a_14869_1051.n0 GND 0.37fF
C439 a_14869_1051.n1 GND 0.33fF
C440 a_14869_1051.n2 GND 0.23fF
C441 a_14869_1051.n3 GND 0.63fF
C442 a_14869_1051.n4 GND 0.28fF
C443 a_14869_1051.n5 GND 0.41fF
C444 a_6149_989.n0 GND 0.53fF
C445 a_6149_989.t12 GND 0.86fF
C446 a_6149_989.n1 GND 0.63fF
C447 a_6149_989.n2 GND 0.53fF
C448 a_6149_989.t7 GND 0.85fF
C449 a_6149_989.n3 GND 0.56fF
C450 a_6149_989.n4 GND 0.53fF
C451 a_6149_989.t6 GND 0.86fF
C452 a_6149_989.n5 GND 0.59fF
C453 a_6149_989.n6 GND 1.74fF
C454 a_6149_989.n7 GND 2.34fF
C455 a_6149_989.n8 GND 0.06fF
C456 a_6149_989.n9 GND 0.08fF
C457 a_6149_989.n10 GND 0.05fF
C458 a_6149_989.n11 GND 0.50fF
C459 a_6149_989.n12 GND 0.65fF
C460 a_6149_989.n13 GND 0.96fF
C461 a_6149_989.n14 GND 0.42fF
C462 a_6149_989.n15 GND 0.81fF
C463 a_3599_411.n0 GND 1.04fF
C464 a_3599_411.n1 GND 1.04fF
C465 a_3599_411.n2 GND 0.73fF
C466 a_3599_411.n3 GND 0.91fF
C467 a_3599_411.n4 GND 1.13fF
C468 a_3599_411.t10 GND 0.85fF
C469 a_3599_411.n5 GND 0.70fF
C470 a_3599_411.n6 GND 3.68fF
C471 a_3599_411.n7 GND 0.71fF
C472 a_3599_411.t12 GND 0.98fF
C473 a_3599_411.n8 GND 0.78fF
C474 a_3599_411.n9 GND 16.28fF
C475 a_3599_411.n10 GND 0.08fF
C476 a_3599_411.n11 GND 0.10fF
C477 a_3599_411.n12 GND 0.07fF
C478 a_3599_411.n13 GND 0.52fF
C479 a_3599_411.n14 GND 0.87fF
C480 a_3599_411.n15 GND 0.65fF
C481 a_3599_411.n16 GND 0.38fF
C482 a_3599_411.n17 GND 1.22fF
C483 a_3473_1050.n0 GND 0.57fF
C484 a_3473_1050.n1 GND 0.67fF
C485 a_3473_1050.n2 GND 0.26fF
C486 a_3473_1050.n3 GND 0.29fF
C487 a_3473_1050.n4 GND 0.71fF
C488 a_3473_1050.n5 GND 0.65fF
C489 a_3473_1050.n6 GND 0.09fF
C490 a_3473_1050.n7 GND 0.38fF
C491 a_3473_1050.n8 GND 0.05fF
C492 a_6884_210.n0 GND 0.07fF
C493 a_6884_210.n1 GND 0.09fF
C494 a_6884_210.n2 GND 0.13fF
C495 a_6884_210.n3 GND 0.11fF
C496 a_6884_210.n4 GND 0.02fF
C497 a_6884_210.n5 GND 0.03fF
C498 a_6884_210.n6 GND 0.06fF
C499 a_6884_210.n7 GND 0.03fF
C500 a_6884_210.n8 GND 0.12fF
C501 a_6884_210.n9 GND 0.06fF
C502 a_6884_210.n10 GND 0.01fF
C503 a_6884_210.t0 GND 0.33fF
C504 a_6603_103.n0 GND 0.20fF
C505 a_6603_103.n1 GND 0.04fF
C506 a_6603_103.n2 GND 0.01fF
C507 a_6603_103.n3 GND 0.03fF
C508 a_6603_103.n4 GND 0.05fF
C509 a_6603_103.n5 GND 0.09fF
C510 a_6603_103.n6 GND 0.07fF
C511 SN.n0 GND 0.87fF
C512 SN.t10 GND 0.80fF
C513 SN.n1 GND 0.83fF
C514 SN.n2 GND 0.87fF
C515 SN.t5 GND 0.80fF
C516 SN.n3 GND 0.65fF
C517 SN.n4 GND 5.21fF
C518 SN.n5 GND 0.87fF
C519 SN.t6 GND 0.80fF
C520 SN.n6 GND 0.65fF
C521 SN.n7 GND 3.64fF
C522 SN.n8 GND 0.87fF
C523 SN.t0 GND 0.80fF
C524 SN.n9 GND 0.65fF
C525 SN.n10 GND 3.64fF
C526 SN.n11 GND 0.87fF
C527 SN.t1 GND 0.80fF
C528 SN.n12 GND 0.65fF
C529 SN.n13 GND 3.64fF
C530 SN.n14 GND 0.87fF
C531 SN.t11 GND 0.80fF
C532 SN.n15 GND 0.65fF
C533 SN.n16 GND 1.73fF
C534 a_8357_1050.n0 GND 0.31fF
C535 a_8357_1050.n1 GND 0.74fF
C536 a_8357_1050.n2 GND 0.05fF
C537 a_8357_1050.n3 GND 0.06fF
C538 a_8357_1050.n4 GND 0.04fF
C539 a_8357_1050.n5 GND 0.40fF
C540 a_8357_1050.n6 GND 0.67fF
C541 a_8357_1050.n7 GND 0.70fF
C542 a_8357_1050.n8 GND 0.27fF
C543 a_8357_1050.n9 GND 0.59fF
C544 VDD.n0 GND 0.12fF
C545 VDD.n1 GND 0.03fF
C546 VDD.n2 GND 0.02fF
C547 VDD.n3 GND 0.05fF
C548 VDD.n4 GND 0.01fF
C549 VDD.n6 GND 0.02fF
C550 VDD.n7 GND 0.02fF
C551 VDD.n8 GND 0.02fF
C552 VDD.n9 GND 0.02fF
C553 VDD.n11 GND 0.02fF
C554 VDD.n14 GND 0.46fF
C555 VDD.n16 GND 0.03fF
C556 VDD.n17 GND 0.02fF
C557 VDD.n18 GND 0.02fF
C558 VDD.n19 GND 0.02fF
C559 VDD.n20 GND 0.04fF
C560 VDD.n21 GND 0.27fF
C561 VDD.n22 GND 0.02fF
C562 VDD.n23 GND 0.03fF
C563 VDD.n24 GND 0.06fF
C564 VDD.n25 GND 0.15fF
C565 VDD.n26 GND 0.20fF
C566 VDD.n27 GND 0.01fF
C567 VDD.n28 GND 0.01fF
C568 VDD.n29 GND 0.07fF
C569 VDD.n30 GND 0.17fF
C570 VDD.n31 GND 0.01fF
C571 VDD.n32 GND 0.02fF
C572 VDD.n33 GND 0.02fF
C573 VDD.n34 GND 0.15fF
C574 VDD.n35 GND 0.20fF
C575 VDD.n36 GND 0.01fF
C576 VDD.n37 GND 0.06fF
C577 VDD.n38 GND 0.01fF
C578 VDD.n39 GND 0.02fF
C579 VDD.n40 GND 0.27fF
C580 VDD.n41 GND 0.01fF
C581 VDD.n42 GND 0.02fF
C582 VDD.n43 GND 0.03fF
C583 VDD.n44 GND 0.02fF
C584 VDD.n45 GND 0.02fF
C585 VDD.n46 GND 0.02fF
C586 VDD.n47 GND 0.18fF
C587 VDD.n48 GND 0.04fF
C588 VDD.n49 GND 0.04fF
C589 VDD.n50 GND 0.02fF
C590 VDD.n52 GND 0.02fF
C591 VDD.n53 GND 0.02fF
C592 VDD.n54 GND 0.02fF
C593 VDD.n55 GND 0.02fF
C594 VDD.n57 GND 0.02fF
C595 VDD.n58 GND 0.02fF
C596 VDD.n59 GND 0.02fF
C597 VDD.n61 GND 0.27fF
C598 VDD.n63 GND 0.02fF
C599 VDD.n64 GND 0.02fF
C600 VDD.n65 GND 0.03fF
C601 VDD.n66 GND 0.02fF
C602 VDD.n67 GND 0.27fF
C603 VDD.n68 GND 0.01fF
C604 VDD.n69 GND 0.02fF
C605 VDD.n70 GND 0.03fF
C606 VDD.n71 GND 0.27fF
C607 VDD.n72 GND 0.01fF
C608 VDD.n73 GND 0.02fF
C609 VDD.n74 GND 0.02fF
C610 VDD.n75 GND 0.27fF
C611 VDD.n76 GND 0.01fF
C612 VDD.n77 GND 0.02fF
C613 VDD.n78 GND 0.02fF
C614 VDD.n79 GND 0.31fF
C615 VDD.n80 GND 0.01fF
C616 VDD.n81 GND 0.03fF
C617 VDD.n82 GND 0.03fF
C618 VDD.n83 GND 0.31fF
C619 VDD.n84 GND 0.01fF
C620 VDD.n85 GND 0.03fF
C621 VDD.n86 GND 0.03fF
C622 VDD.n87 GND 0.27fF
C623 VDD.n88 GND 0.01fF
C624 VDD.n89 GND 0.02fF
C625 VDD.n90 GND 0.02fF
C626 VDD.n91 GND 0.27fF
C627 VDD.n92 GND 0.01fF
C628 VDD.n93 GND 0.02fF
C629 VDD.n94 GND 0.02fF
C630 VDD.n95 GND 0.27fF
C631 VDD.n96 GND 0.01fF
C632 VDD.n97 GND 0.02fF
C633 VDD.n98 GND 0.03fF
C634 VDD.n99 GND 0.02fF
C635 VDD.n100 GND 0.02fF
C636 VDD.n101 GND 0.02fF
C637 VDD.n102 GND 0.22fF
C638 VDD.n103 GND 0.04fF
C639 VDD.n104 GND 0.03fF
C640 VDD.n105 GND 0.02fF
C641 VDD.n106 GND 0.02fF
C642 VDD.n107 GND 0.02fF
C643 VDD.n108 GND 0.03fF
C644 VDD.n109 GND 0.02fF
C645 VDD.n111 GND 0.02fF
C646 VDD.n112 GND 0.02fF
C647 VDD.n113 GND 0.02fF
C648 VDD.n115 GND 0.27fF
C649 VDD.n117 GND 0.02fF
C650 VDD.n118 GND 0.02fF
C651 VDD.n119 GND 0.03fF
C652 VDD.n120 GND 0.02fF
C653 VDD.n121 GND 0.27fF
C654 VDD.n122 GND 0.01fF
C655 VDD.n123 GND 0.02fF
C656 VDD.n124 GND 0.03fF
C657 VDD.n125 GND 0.27fF
C658 VDD.n126 GND 0.01fF
C659 VDD.n127 GND 0.02fF
C660 VDD.n128 GND 0.02fF
C661 VDD.n129 GND 0.27fF
C662 VDD.n130 GND 0.01fF
C663 VDD.n131 GND 0.02fF
C664 VDD.n132 GND 0.02fF
C665 VDD.n133 GND 0.31fF
C666 VDD.n134 GND 0.01fF
C667 VDD.n135 GND 0.03fF
C668 VDD.n136 GND 0.03fF
C669 VDD.n137 GND 0.31fF
C670 VDD.n138 GND 0.01fF
C671 VDD.n139 GND 0.03fF
C672 VDD.n140 GND 0.03fF
C673 VDD.n141 GND 0.27fF
C674 VDD.n142 GND 0.01fF
C675 VDD.n143 GND 0.02fF
C676 VDD.n144 GND 0.02fF
C677 VDD.n145 GND 0.27fF
C678 VDD.n146 GND 0.01fF
C679 VDD.n147 GND 0.02fF
C680 VDD.n148 GND 0.02fF
C681 VDD.n149 GND 0.27fF
C682 VDD.n150 GND 0.01fF
C683 VDD.n151 GND 0.02fF
C684 VDD.n152 GND 0.03fF
C685 VDD.n153 GND 0.02fF
C686 VDD.n154 GND 0.02fF
C687 VDD.n155 GND 0.02fF
C688 VDD.n156 GND 0.22fF
C689 VDD.n157 GND 0.04fF
C690 VDD.n158 GND 0.03fF
C691 VDD.n159 GND 0.02fF
C692 VDD.n160 GND 0.02fF
C693 VDD.n161 GND 0.02fF
C694 VDD.n162 GND 0.03fF
C695 VDD.n163 GND 0.02fF
C696 VDD.n165 GND 0.02fF
C697 VDD.n166 GND 0.02fF
C698 VDD.n167 GND 0.02fF
C699 VDD.n169 GND 0.27fF
C700 VDD.n171 GND 0.02fF
C701 VDD.n172 GND 0.02fF
C702 VDD.n173 GND 0.03fF
C703 VDD.n174 GND 0.02fF
C704 VDD.n175 GND 0.27fF
C705 VDD.n176 GND 0.01fF
C706 VDD.n177 GND 0.02fF
C707 VDD.n178 GND 0.03fF
C708 VDD.n179 GND 0.06fF
C709 VDD.n180 GND 0.24fF
C710 VDD.n181 GND 0.01fF
C711 VDD.n182 GND 0.01fF
C712 VDD.n183 GND 0.02fF
C713 VDD.n184 GND 0.14fF
C714 VDD.n185 GND 0.17fF
C715 VDD.n186 GND 0.01fF
C716 VDD.n187 GND 0.02fF
C717 VDD.n188 GND 0.02fF
C718 VDD.n189 GND 0.11fF
C719 VDD.n190 GND 0.03fF
C720 VDD.n191 GND 0.31fF
C721 VDD.n192 GND 0.01fF
C722 VDD.n193 GND 0.02fF
C723 VDD.n194 GND 0.03fF
C724 VDD.n195 GND 0.17fF
C725 VDD.n196 GND 0.14fF
C726 VDD.n197 GND 0.01fF
C727 VDD.n198 GND 0.02fF
C728 VDD.n199 GND 0.03fF
C729 VDD.n200 GND 0.14fF
C730 VDD.n201 GND 0.16fF
C731 VDD.n202 GND 0.01fF
C732 VDD.n203 GND 0.02fF
C733 VDD.n204 GND 0.02fF
C734 VDD.n205 GND 0.06fF
C735 VDD.n206 GND 0.25fF
C736 VDD.n207 GND 0.01fF
C737 VDD.n208 GND 0.01fF
C738 VDD.n209 GND 0.02fF
C739 VDD.n210 GND 0.27fF
C740 VDD.n211 GND 0.01fF
C741 VDD.n212 GND 0.02fF
C742 VDD.n213 GND 0.03fF
C743 VDD.n214 GND 0.02fF
C744 VDD.n215 GND 0.02fF
C745 VDD.n216 GND 0.02fF
C746 VDD.n217 GND 0.26fF
C747 VDD.n218 GND 0.04fF
C748 VDD.n219 GND 0.03fF
C749 VDD.n220 GND 0.02fF
C750 VDD.n221 GND 0.02fF
C751 VDD.n222 GND 0.02fF
C752 VDD.n223 GND 0.03fF
C753 VDD.n224 GND 0.02fF
C754 VDD.n226 GND 0.02fF
C755 VDD.n227 GND 0.02fF
C756 VDD.n228 GND 0.02fF
C757 VDD.n230 GND 0.27fF
C758 VDD.n232 GND 0.02fF
C759 VDD.n233 GND 0.02fF
C760 VDD.n234 GND 0.03fF
C761 VDD.n235 GND 0.02fF
C762 VDD.n236 GND 0.27fF
C763 VDD.n237 GND 0.01fF
C764 VDD.n238 GND 0.02fF
C765 VDD.n239 GND 0.03fF
C766 VDD.n240 GND 0.27fF
C767 VDD.n241 GND 0.01fF
C768 VDD.n242 GND 0.02fF
C769 VDD.n243 GND 0.02fF
C770 VDD.n244 GND 0.22fF
C771 VDD.n245 GND 0.01fF
C772 VDD.n246 GND 0.07fF
C773 VDD.n247 GND 0.02fF
C774 VDD.n248 GND 0.14fF
C775 VDD.n249 GND 0.17fF
C776 VDD.n250 GND 0.01fF
C777 VDD.n251 GND 0.02fF
C778 VDD.n252 GND 0.02fF
C779 VDD.n253 GND 0.14fF
C780 VDD.n254 GND 0.16fF
C781 VDD.n255 GND 0.01fF
C782 VDD.n256 GND 0.11fF
C783 VDD.n257 GND 0.02fF
C784 VDD.n258 GND 0.02fF
C785 VDD.n259 GND 0.02fF
C786 VDD.n260 GND 0.18fF
C787 VDD.n261 GND 0.14fF
C788 VDD.n262 GND 0.01fF
C789 VDD.n263 GND 0.02fF
C790 VDD.n264 GND 0.03fF
C791 VDD.n265 GND 0.18fF
C792 VDD.n266 GND 0.15fF
C793 VDD.n267 GND 0.01fF
C794 VDD.n268 GND 0.02fF
C795 VDD.n269 GND 0.03fF
C796 VDD.n270 GND 0.11fF
C797 VDD.n271 GND 0.02fF
C798 VDD.n272 GND 0.14fF
C799 VDD.n273 GND 0.16fF
C800 VDD.n274 GND 0.01fF
C801 VDD.n275 GND 0.02fF
C802 VDD.n276 GND 0.02fF
C803 VDD.n277 GND 0.14fF
C804 VDD.n278 GND 0.17fF
C805 VDD.n279 GND 0.01fF
C806 VDD.n280 GND 0.02fF
C807 VDD.n281 GND 0.02fF
C808 VDD.n282 GND 0.06fF
C809 VDD.n283 GND 0.23fF
C810 VDD.n284 GND 0.01fF
C811 VDD.n285 GND 0.01fF
C812 VDD.n286 GND 0.02fF
C813 VDD.n287 GND 0.27fF
C814 VDD.n288 GND 0.01fF
C815 VDD.n289 GND 0.02fF
C816 VDD.n290 GND 0.02fF
C817 VDD.n291 GND 0.27fF
C818 VDD.n292 GND 0.01fF
C819 VDD.n293 GND 0.02fF
C820 VDD.n294 GND 0.03fF
C821 VDD.n295 GND 0.02fF
C822 VDD.n296 GND 0.02fF
C823 VDD.n297 GND 0.02fF
C824 VDD.n298 GND 0.26fF
C825 VDD.n299 GND 0.04fF
C826 VDD.n300 GND 0.03fF
C827 VDD.n301 GND 0.02fF
C828 VDD.n302 GND 0.02fF
C829 VDD.n303 GND 0.02fF
C830 VDD.n304 GND 0.03fF
C831 VDD.n305 GND 0.02fF
C832 VDD.n307 GND 0.02fF
C833 VDD.n308 GND 0.02fF
C834 VDD.n309 GND 0.02fF
C835 VDD.n311 GND 0.27fF
C836 VDD.n313 GND 0.02fF
C837 VDD.n314 GND 0.02fF
C838 VDD.n315 GND 0.03fF
C839 VDD.n316 GND 0.02fF
C840 VDD.n317 GND 0.27fF
C841 VDD.n318 GND 0.01fF
C842 VDD.n319 GND 0.02fF
C843 VDD.n320 GND 0.03fF
C844 VDD.n321 GND 0.06fF
C845 VDD.n322 GND 0.24fF
C846 VDD.n323 GND 0.01fF
C847 VDD.n324 GND 0.01fF
C848 VDD.n325 GND 0.02fF
C849 VDD.n326 GND 0.14fF
C850 VDD.n327 GND 0.17fF
C851 VDD.n328 GND 0.01fF
C852 VDD.n329 GND 0.02fF
C853 VDD.n330 GND 0.02fF
C854 VDD.n331 GND 0.11fF
C855 VDD.n332 GND 0.03fF
C856 VDD.n333 GND 0.31fF
C857 VDD.n334 GND 0.01fF
C858 VDD.n335 GND 0.02fF
C859 VDD.n336 GND 0.03fF
C860 VDD.n337 GND 0.17fF
C861 VDD.n338 GND 0.14fF
C862 VDD.n339 GND 0.01fF
C863 VDD.n340 GND 0.02fF
C864 VDD.n341 GND 0.03fF
C865 VDD.n342 GND 0.14fF
C866 VDD.n343 GND 0.16fF
C867 VDD.n344 GND 0.01fF
C868 VDD.n345 GND 0.02fF
C869 VDD.n346 GND 0.02fF
C870 VDD.n347 GND 0.06fF
C871 VDD.n348 GND 0.25fF
C872 VDD.n349 GND 0.01fF
C873 VDD.n350 GND 0.01fF
C874 VDD.n351 GND 0.02fF
C875 VDD.n352 GND 0.27fF
C876 VDD.n353 GND 0.01fF
C877 VDD.n354 GND 0.02fF
C878 VDD.n355 GND 0.03fF
C879 VDD.n356 GND 0.02fF
C880 VDD.n357 GND 0.02fF
C881 VDD.n358 GND 0.02fF
C882 VDD.n359 GND 0.22fF
C883 VDD.n360 GND 0.04fF
C884 VDD.n361 GND 0.03fF
C885 VDD.n362 GND 0.02fF
C886 VDD.n363 GND 0.02fF
C887 VDD.n364 GND 0.02fF
C888 VDD.n365 GND 0.03fF
C889 VDD.n366 GND 0.02fF
C890 VDD.n368 GND 0.02fF
C891 VDD.n369 GND 0.02fF
C892 VDD.n370 GND 0.02fF
C893 VDD.n372 GND 0.27fF
C894 VDD.n374 GND 0.02fF
C895 VDD.n375 GND 0.02fF
C896 VDD.n376 GND 0.03fF
C897 VDD.n377 GND 0.02fF
C898 VDD.n378 GND 0.27fF
C899 VDD.n379 GND 0.01fF
C900 VDD.n380 GND 0.02fF
C901 VDD.n381 GND 0.03fF
C902 VDD.n382 GND 0.06fF
C903 VDD.n383 GND 0.24fF
C904 VDD.n384 GND 0.01fF
C905 VDD.n385 GND 0.01fF
C906 VDD.n386 GND 0.02fF
C907 VDD.n387 GND 0.14fF
C908 VDD.n388 GND 0.17fF
C909 VDD.n389 GND 0.01fF
C910 VDD.n390 GND 0.02fF
C911 VDD.n391 GND 0.02fF
C912 VDD.n392 GND 0.11fF
C913 VDD.n393 GND 0.03fF
C914 VDD.n394 GND 0.31fF
C915 VDD.n395 GND 0.01fF
C916 VDD.n396 GND 0.02fF
C917 VDD.n397 GND 0.03fF
C918 VDD.n398 GND 0.17fF
C919 VDD.n399 GND 0.14fF
C920 VDD.n400 GND 0.01fF
C921 VDD.n401 GND 0.02fF
C922 VDD.n402 GND 0.03fF
C923 VDD.n403 GND 0.14fF
C924 VDD.n404 GND 0.16fF
C925 VDD.n405 GND 0.01fF
C926 VDD.n406 GND 0.02fF
C927 VDD.n407 GND 0.02fF
C928 VDD.n408 GND 0.06fF
C929 VDD.n409 GND 0.25fF
C930 VDD.n410 GND 0.01fF
C931 VDD.n411 GND 0.01fF
C932 VDD.n412 GND 0.02fF
C933 VDD.n413 GND 0.27fF
C934 VDD.n414 GND 0.01fF
C935 VDD.n415 GND 0.02fF
C936 VDD.n416 GND 0.03fF
C937 VDD.n417 GND 0.02fF
C938 VDD.n418 GND 0.02fF
C939 VDD.n419 GND 0.02fF
C940 VDD.n420 GND 0.26fF
C941 VDD.n421 GND 0.04fF
C942 VDD.n422 GND 0.03fF
C943 VDD.n423 GND 0.02fF
C944 VDD.n424 GND 0.02fF
C945 VDD.n425 GND 0.02fF
C946 VDD.n426 GND 0.03fF
C947 VDD.n427 GND 0.02fF
C948 VDD.n429 GND 0.02fF
C949 VDD.n430 GND 0.02fF
C950 VDD.n431 GND 0.02fF
C951 VDD.n433 GND 0.27fF
C952 VDD.n435 GND 0.02fF
C953 VDD.n436 GND 0.02fF
C954 VDD.n437 GND 0.03fF
C955 VDD.n438 GND 0.02fF
C956 VDD.n439 GND 0.27fF
C957 VDD.n440 GND 0.01fF
C958 VDD.n441 GND 0.02fF
C959 VDD.n442 GND 0.03fF
C960 VDD.n443 GND 0.27fF
C961 VDD.n444 GND 0.01fF
C962 VDD.n445 GND 0.02fF
C963 VDD.n446 GND 0.02fF
C964 VDD.n447 GND 0.22fF
C965 VDD.n448 GND 0.01fF
C966 VDD.n449 GND 0.07fF
C967 VDD.n450 GND 0.02fF
C968 VDD.n451 GND 0.14fF
C969 VDD.n452 GND 0.17fF
C970 VDD.n453 GND 0.01fF
C971 VDD.n454 GND 0.02fF
C972 VDD.n455 GND 0.02fF
C973 VDD.n456 GND 0.14fF
C974 VDD.n457 GND 0.16fF
C975 VDD.n458 GND 0.01fF
C976 VDD.n459 GND 0.11fF
C977 VDD.n460 GND 0.02fF
C978 VDD.n461 GND 0.02fF
C979 VDD.n462 GND 0.02fF
C980 VDD.n463 GND 0.18fF
C981 VDD.n464 GND 0.14fF
C982 VDD.n465 GND 0.01fF
C983 VDD.n466 GND 0.02fF
C984 VDD.n467 GND 0.03fF
C985 VDD.n468 GND 0.18fF
C986 VDD.n469 GND 0.15fF
C987 VDD.n470 GND 0.01fF
C988 VDD.n471 GND 0.02fF
C989 VDD.n472 GND 0.03fF
C990 VDD.n473 GND 0.11fF
C991 VDD.n474 GND 0.02fF
C992 VDD.n475 GND 0.14fF
C993 VDD.n476 GND 0.16fF
C994 VDD.n477 GND 0.01fF
C995 VDD.n478 GND 0.02fF
C996 VDD.n479 GND 0.02fF
C997 VDD.n480 GND 0.14fF
C998 VDD.n481 GND 0.17fF
C999 VDD.n482 GND 0.01fF
C1000 VDD.n483 GND 0.02fF
C1001 VDD.n484 GND 0.02fF
C1002 VDD.n485 GND 0.06fF
C1003 VDD.n486 GND 0.23fF
C1004 VDD.n487 GND 0.01fF
C1005 VDD.n488 GND 0.01fF
C1006 VDD.n489 GND 0.02fF
C1007 VDD.n490 GND 0.27fF
C1008 VDD.n491 GND 0.01fF
C1009 VDD.n492 GND 0.02fF
C1010 VDD.n493 GND 0.02fF
C1011 VDD.n494 GND 0.27fF
C1012 VDD.n495 GND 0.01fF
C1013 VDD.n496 GND 0.02fF
C1014 VDD.n497 GND 0.03fF
C1015 VDD.n498 GND 0.02fF
C1016 VDD.n499 GND 0.02fF
C1017 VDD.n500 GND 0.02fF
C1018 VDD.n501 GND 0.31fF
C1019 VDD.n502 GND 0.04fF
C1020 VDD.n503 GND 0.03fF
C1021 VDD.n504 GND 0.02fF
C1022 VDD.n505 GND 0.02fF
C1023 VDD.n506 GND 0.02fF
C1024 VDD.n507 GND 0.03fF
C1025 VDD.n508 GND 0.02fF
C1026 VDD.n510 GND 0.02fF
C1027 VDD.n511 GND 0.02fF
C1028 VDD.n512 GND 0.02fF
C1029 VDD.n514 GND 0.27fF
C1030 VDD.n516 GND 0.02fF
C1031 VDD.n517 GND 0.02fF
C1032 VDD.n518 GND 0.03fF
C1033 VDD.n519 GND 0.02fF
C1034 VDD.n520 GND 0.27fF
C1035 VDD.n521 GND 0.01fF
C1036 VDD.n522 GND 0.02fF
C1037 VDD.n523 GND 0.03fF
C1038 VDD.n524 GND 0.27fF
C1039 VDD.n525 GND 0.01fF
C1040 VDD.n526 GND 0.02fF
C1041 VDD.n527 GND 0.02fF
C1042 VDD.n528 GND 0.22fF
C1043 VDD.n529 GND 0.01fF
C1044 VDD.n530 GND 0.07fF
C1045 VDD.n531 GND 0.02fF
C1046 VDD.n532 GND 0.14fF
C1047 VDD.n533 GND 0.17fF
C1048 VDD.n534 GND 0.01fF
C1049 VDD.n535 GND 0.02fF
C1050 VDD.n536 GND 0.02fF
C1051 VDD.n537 GND 0.14fF
C1052 VDD.n538 GND 0.16fF
C1053 VDD.n539 GND 0.01fF
C1054 VDD.n540 GND 0.11fF
C1055 VDD.n541 GND 0.02fF
C1056 VDD.n542 GND 0.02fF
C1057 VDD.n543 GND 0.02fF
C1058 VDD.n544 GND 0.18fF
C1059 VDD.n545 GND 0.14fF
C1060 VDD.n546 GND 0.01fF
C1061 VDD.n547 GND 0.02fF
C1062 VDD.n548 GND 0.03fF
C1063 VDD.n549 GND 0.18fF
C1064 VDD.n550 GND 0.15fF
C1065 VDD.n551 GND 0.01fF
C1066 VDD.n552 GND 0.02fF
C1067 VDD.n553 GND 0.03fF
C1068 VDD.n554 GND 0.11fF
C1069 VDD.n555 GND 0.02fF
C1070 VDD.n556 GND 0.14fF
C1071 VDD.n557 GND 0.16fF
C1072 VDD.n558 GND 0.01fF
C1073 VDD.n559 GND 0.02fF
C1074 VDD.n560 GND 0.02fF
C1075 VDD.n561 GND 0.14fF
C1076 VDD.n562 GND 0.17fF
C1077 VDD.n563 GND 0.01fF
C1078 VDD.n564 GND 0.02fF
C1079 VDD.n565 GND 0.02fF
C1080 VDD.n566 GND 0.06fF
C1081 VDD.n567 GND 0.23fF
C1082 VDD.n568 GND 0.01fF
C1083 VDD.n569 GND 0.01fF
C1084 VDD.n570 GND 0.02fF
C1085 VDD.n571 GND 0.27fF
C1086 VDD.n572 GND 0.01fF
C1087 VDD.n573 GND 0.02fF
C1088 VDD.n574 GND 0.02fF
C1089 VDD.n575 GND 0.27fF
C1090 VDD.n576 GND 0.01fF
C1091 VDD.n577 GND 0.02fF
C1092 VDD.n578 GND 0.03fF
C1093 VDD.n579 GND 0.02fF
C1094 VDD.n580 GND 0.02fF
C1095 VDD.n581 GND 0.02fF
C1096 VDD.n582 GND 0.26fF
C1097 VDD.n583 GND 0.04fF
C1098 VDD.n584 GND 0.03fF
C1099 VDD.n585 GND 0.02fF
C1100 VDD.n586 GND 0.02fF
C1101 VDD.n587 GND 0.02fF
C1102 VDD.n588 GND 0.03fF
C1103 VDD.n589 GND 0.02fF
C1104 VDD.n591 GND 0.02fF
C1105 VDD.n592 GND 0.02fF
C1106 VDD.n593 GND 0.02fF
C1107 VDD.n595 GND 0.27fF
C1108 VDD.n597 GND 0.02fF
C1109 VDD.n598 GND 0.02fF
C1110 VDD.n599 GND 0.03fF
C1111 VDD.n600 GND 0.02fF
C1112 VDD.n601 GND 0.27fF
C1113 VDD.n602 GND 0.01fF
C1114 VDD.n603 GND 0.02fF
C1115 VDD.n604 GND 0.03fF
C1116 VDD.n605 GND 0.06fF
C1117 VDD.n606 GND 0.24fF
C1118 VDD.n607 GND 0.01fF
C1119 VDD.n608 GND 0.01fF
C1120 VDD.n609 GND 0.02fF
C1121 VDD.n610 GND 0.14fF
C1122 VDD.n611 GND 0.17fF
C1123 VDD.n612 GND 0.01fF
C1124 VDD.n613 GND 0.02fF
C1125 VDD.n614 GND 0.02fF
C1126 VDD.n615 GND 0.11fF
C1127 VDD.n616 GND 0.03fF
C1128 VDD.n617 GND 0.31fF
C1129 VDD.n618 GND 0.01fF
C1130 VDD.n619 GND 0.02fF
C1131 VDD.n620 GND 0.03fF
C1132 VDD.n621 GND 0.17fF
C1133 VDD.n622 GND 0.14fF
C1134 VDD.n623 GND 0.01fF
C1135 VDD.n624 GND 0.02fF
C1136 VDD.n625 GND 0.03fF
C1137 VDD.n626 GND 0.14fF
C1138 VDD.n627 GND 0.16fF
C1139 VDD.n628 GND 0.01fF
C1140 VDD.n629 GND 0.02fF
C1141 VDD.n630 GND 0.02fF
C1142 VDD.n631 GND 0.06fF
C1143 VDD.n632 GND 0.25fF
C1144 VDD.n633 GND 0.01fF
C1145 VDD.n634 GND 0.01fF
C1146 VDD.n635 GND 0.02fF
C1147 VDD.n636 GND 0.27fF
C1148 VDD.n637 GND 0.01fF
C1149 VDD.n638 GND 0.02fF
C1150 VDD.n639 GND 0.03fF
C1151 VDD.n640 GND 0.02fF
C1152 VDD.n641 GND 0.02fF
C1153 VDD.n642 GND 0.02fF
C1154 VDD.n643 GND 0.26fF
C1155 VDD.n644 GND 0.04fF
C1156 VDD.n645 GND 0.03fF
C1157 VDD.n646 GND 0.02fF
C1158 VDD.n647 GND 0.02fF
C1159 VDD.n648 GND 0.02fF
C1160 VDD.n649 GND 0.03fF
C1161 VDD.n650 GND 0.02fF
C1162 VDD.n652 GND 0.02fF
C1163 VDD.n653 GND 0.02fF
C1164 VDD.n654 GND 0.02fF
C1165 VDD.n656 GND 0.27fF
C1166 VDD.n658 GND 0.02fF
C1167 VDD.n659 GND 0.02fF
C1168 VDD.n660 GND 0.03fF
C1169 VDD.n661 GND 0.02fF
C1170 VDD.n662 GND 0.27fF
C1171 VDD.n663 GND 0.01fF
C1172 VDD.n664 GND 0.02fF
C1173 VDD.n665 GND 0.03fF
C1174 VDD.n666 GND 0.27fF
C1175 VDD.n667 GND 0.01fF
C1176 VDD.n668 GND 0.02fF
C1177 VDD.n669 GND 0.02fF
C1178 VDD.n670 GND 0.22fF
C1179 VDD.n671 GND 0.01fF
C1180 VDD.n672 GND 0.07fF
C1181 VDD.n673 GND 0.02fF
C1182 VDD.n674 GND 0.14fF
C1183 VDD.n675 GND 0.17fF
C1184 VDD.n676 GND 0.01fF
C1185 VDD.n677 GND 0.02fF
C1186 VDD.n678 GND 0.02fF
C1187 VDD.n679 GND 0.14fF
C1188 VDD.n680 GND 0.16fF
C1189 VDD.n681 GND 0.01fF
C1190 VDD.n682 GND 0.11fF
C1191 VDD.n683 GND 0.02fF
C1192 VDD.n684 GND 0.02fF
C1193 VDD.n685 GND 0.02fF
C1194 VDD.n686 GND 0.18fF
C1195 VDD.n687 GND 0.14fF
C1196 VDD.n688 GND 0.01fF
C1197 VDD.n689 GND 0.02fF
C1198 VDD.n690 GND 0.03fF
C1199 VDD.n691 GND 0.18fF
C1200 VDD.n692 GND 0.15fF
C1201 VDD.n693 GND 0.01fF
C1202 VDD.n694 GND 0.02fF
C1203 VDD.n695 GND 0.03fF
C1204 VDD.n696 GND 0.11fF
C1205 VDD.n697 GND 0.02fF
C1206 VDD.n698 GND 0.14fF
C1207 VDD.n699 GND 0.16fF
C1208 VDD.n700 GND 0.01fF
C1209 VDD.n701 GND 0.02fF
C1210 VDD.n702 GND 0.02fF
C1211 VDD.n703 GND 0.14fF
C1212 VDD.n704 GND 0.17fF
C1213 VDD.n705 GND 0.01fF
C1214 VDD.n706 GND 0.02fF
C1215 VDD.n707 GND 0.02fF
C1216 VDD.n708 GND 0.06fF
C1217 VDD.n709 GND 0.23fF
C1218 VDD.n710 GND 0.01fF
C1219 VDD.n711 GND 0.01fF
C1220 VDD.n712 GND 0.02fF
C1221 VDD.n713 GND 0.27fF
C1222 VDD.n714 GND 0.01fF
C1223 VDD.n715 GND 0.02fF
C1224 VDD.n716 GND 0.02fF
C1225 VDD.n717 GND 0.27fF
C1226 VDD.n718 GND 0.01fF
C1227 VDD.n719 GND 0.02fF
C1228 VDD.n720 GND 0.03fF
C1229 VDD.n721 GND 0.02fF
C1230 VDD.n722 GND 0.02fF
C1231 VDD.n723 GND 0.02fF
C1232 VDD.n724 GND 0.26fF
C1233 VDD.n725 GND 0.04fF
C1234 VDD.n726 GND 0.03fF
C1235 VDD.n727 GND 0.02fF
C1236 VDD.n728 GND 0.02fF
C1237 VDD.n729 GND 0.02fF
C1238 VDD.n730 GND 0.03fF
C1239 VDD.n731 GND 0.02fF
C1240 VDD.n733 GND 0.02fF
C1241 VDD.n734 GND 0.02fF
C1242 VDD.n735 GND 0.02fF
C1243 VDD.n737 GND 0.27fF
C1244 VDD.n739 GND 0.02fF
C1245 VDD.n740 GND 0.02fF
C1246 VDD.n741 GND 0.03fF
C1247 VDD.n742 GND 0.02fF
C1248 VDD.n743 GND 0.27fF
C1249 VDD.n744 GND 0.01fF
C1250 VDD.n745 GND 0.02fF
C1251 VDD.n746 GND 0.03fF
C1252 VDD.n747 GND 0.06fF
C1253 VDD.n748 GND 0.24fF
C1254 VDD.n749 GND 0.01fF
C1255 VDD.n750 GND 0.01fF
C1256 VDD.n751 GND 0.02fF
C1257 VDD.n752 GND 0.14fF
C1258 VDD.n753 GND 0.17fF
C1259 VDD.n754 GND 0.01fF
C1260 VDD.n755 GND 0.02fF
C1261 VDD.n756 GND 0.02fF
C1262 VDD.n757 GND 0.02fF
C1263 VDD.n758 GND 0.02fF
C1264 VDD.n759 GND 0.02fF
C1265 VDD.n760 GND 0.15fF
C1266 VDD.n761 GND 0.03fF
C1267 VDD.n762 GND 0.02fF
C1268 VDD.n763 GND 0.02fF
C1269 VDD.n764 GND 0.02fF
C1270 VDD.n765 GND 0.03fF
C1271 VDD.n766 GND 0.02fF
C1272 VDD.n768 GND 0.02fF
C1273 VDD.n769 GND 0.02fF
C1274 VDD.n770 GND 0.02fF
C1275 VDD.n772 GND 0.46fF
C1276 VDD.n774 GND 0.03fF
C1277 VDD.n775 GND 0.04fF
C1278 VDD.n776 GND 0.27fF
C1279 VDD.n777 GND 0.02fF
C1280 VDD.n778 GND 0.03fF
C1281 VDD.n779 GND 0.03fF
C1282 VDD.n780 GND 0.06fF
C1283 VDD.n781 GND 0.25fF
C1284 VDD.n782 GND 0.01fF
C1285 VDD.n783 GND 0.01fF
C1286 VDD.n784 GND 0.02fF
C1287 VDD.n785 GND 0.14fF
C1288 VDD.n786 GND 0.16fF
C1289 VDD.n787 GND 0.01fF
C1290 VDD.n788 GND 0.02fF
C1291 VDD.n789 GND 0.02fF
C1292 VDD.n790 GND 0.17fF
C1293 VDD.n791 GND 0.14fF
C1294 VDD.n792 GND 0.01fF
C1295 VDD.n793 GND 0.02fF
C1296 VDD.n794 GND 0.03fF
C1297 VDD.n795 GND 0.11fF
C1298 VDD.n796 GND 0.03fF
C1299 VDD.n797 GND 0.31fF
C1300 VDD.n798 GND 0.01fF
C1301 VDD.n799 GND 0.02fF
C1302 VDD.n800 GND 0.03fF
C1303 VDD.n801 GND 0.14fF
C1304 VDD.n802 GND 0.17fF
C1305 VDD.n803 GND 0.01fF
C1306 VDD.n804 GND 0.02fF
C1307 VDD.n805 GND 0.02fF
C1308 VDD.n806 GND 0.06fF
C1309 VDD.n807 GND 0.24fF
C1310 VDD.n808 GND 0.01fF
C1311 VDD.n809 GND 0.01fF
C1312 VDD.n810 GND 0.02fF
C1313 VDD.n811 GND 0.27fF
C1314 VDD.n812 GND 0.01fF
C1315 VDD.n813 GND 0.02fF
C1316 VDD.n814 GND 0.03fF
C1317 VDD.n815 GND 0.02fF
C1318 VDD.n816 GND 0.02fF
C1319 VDD.n817 GND 0.02fF
C1320 VDD.n818 GND 0.02fF
C1321 VDD.n819 GND 0.02fF
C1322 VDD.n820 GND 0.02fF
C1323 VDD.n822 GND 0.02fF
C1324 VDD.n823 GND 0.02fF
C1325 VDD.n824 GND 0.02fF
C1326 VDD.n825 GND 0.02fF
C1327 VDD.n827 GND 0.04fF
C1328 VDD.n828 GND 0.02fF
C1329 VDD.n829 GND 0.27fF
C1330 VDD.n830 GND 0.04fF
C1331 VDD.n832 GND 0.27fF
C1332 VDD.n834 GND 0.02fF
C1333 VDD.n835 GND 0.02fF
C1334 VDD.n836 GND 0.03fF
C1335 VDD.n837 GND 0.02fF
C1336 VDD.n838 GND 0.27fF
C1337 VDD.n839 GND 0.01fF
C1338 VDD.n840 GND 0.02fF
C1339 VDD.n841 GND 0.03fF
C1340 VDD.n842 GND 0.27fF
C1341 VDD.n843 GND 0.01fF
C1342 VDD.n844 GND 0.02fF
C1343 VDD.n845 GND 0.02fF
C1344 VDD.n846 GND 0.06fF
C1345 VDD.n847 GND 0.23fF
C1346 VDD.n848 GND 0.01fF
C1347 VDD.n849 GND 0.01fF
C1348 VDD.n850 GND 0.02fF
C1349 VDD.n851 GND 0.14fF
C1350 VDD.n852 GND 0.17fF
C1351 VDD.n853 GND 0.01fF
C1352 VDD.n854 GND 0.02fF
C1353 VDD.n855 GND 0.02fF
C1354 VDD.n856 GND 0.11fF
C1355 VDD.n857 GND 0.02fF
C1356 VDD.n858 GND 0.14fF
C1357 VDD.n859 GND 0.16fF
C1358 VDD.n860 GND 0.01fF
C1359 VDD.n861 GND 0.02fF
C1360 VDD.n862 GND 0.02fF
C1361 VDD.n863 GND 0.18fF
C1362 VDD.n864 GND 0.15fF
C1363 VDD.n865 GND 0.01fF
C1364 VDD.n866 GND 0.02fF
C1365 VDD.n867 GND 0.03fF
C1366 VDD.n868 GND 0.18fF
C1367 VDD.n869 GND 0.14fF
C1368 VDD.n870 GND 0.01fF
C1369 VDD.n871 GND 0.02fF
C1370 VDD.n872 GND 0.03fF
C1371 VDD.n873 GND 0.14fF
C1372 VDD.n874 GND 0.16fF
C1373 VDD.n875 GND 0.01fF
C1374 VDD.n876 GND 0.11fF
C1375 VDD.n877 GND 0.02fF
C1376 VDD.n878 GND 0.02fF
C1377 VDD.n879 GND 0.02fF
C1378 VDD.n880 GND 0.14fF
C1379 VDD.n881 GND 0.17fF
C1380 VDD.n882 GND 0.01fF
C1381 VDD.n883 GND 0.02fF
C1382 VDD.n884 GND 0.02fF
C1383 VDD.n885 GND 0.22fF
C1384 VDD.n886 GND 0.01fF
C1385 VDD.n887 GND 0.07fF
C1386 VDD.n888 GND 0.02fF
C1387 VDD.n889 GND 0.27fF
C1388 VDD.n890 GND 0.01fF
C1389 VDD.n891 GND 0.02fF
C1390 VDD.n892 GND 0.02fF
C1391 VDD.n893 GND 0.27fF
C1392 VDD.n894 GND 0.01fF
C1393 VDD.n895 GND 0.02fF
C1394 VDD.n896 GND 0.03fF
C1395 VDD.n897 GND 0.02fF
C1396 VDD.n898 GND 0.02fF
C1397 VDD.n899 GND 0.02fF
C1398 VDD.n900 GND 0.31fF
C1399 VDD.n901 GND 0.04fF
C1400 VDD.n902 GND 0.03fF
C1401 VDD.n903 GND 0.02fF
C1402 VDD.n904 GND 0.02fF
C1403 VDD.n905 GND 0.02fF
C1404 VDD.n906 GND 0.03fF
C1405 VDD.n907 GND 0.02fF
C1406 VDD.n909 GND 0.02fF
C1407 VDD.n910 GND 0.02fF
C1408 VDD.n911 GND 0.02fF
C1409 VDD.n913 GND 0.27fF
C1410 VDD.n915 GND 0.02fF
C1411 VDD.n916 GND 0.02fF
C1412 VDD.n917 GND 0.03fF
C1413 VDD.n918 GND 0.02fF
C1414 VDD.n919 GND 0.27fF
C1415 VDD.n920 GND 0.01fF
C1416 VDD.n921 GND 0.02fF
C1417 VDD.n922 GND 0.03fF
C1418 VDD.n923 GND 0.27fF
C1419 VDD.n924 GND 0.01fF
C1420 VDD.n925 GND 0.02fF
C1421 VDD.n926 GND 0.02fF
C1422 VDD.n927 GND 0.06fF
C1423 VDD.n928 GND 0.23fF
C1424 VDD.n929 GND 0.01fF
C1425 VDD.n930 GND 0.01fF
C1426 VDD.n931 GND 0.02fF
C1427 VDD.n932 GND 0.14fF
C1428 VDD.n933 GND 0.17fF
C1429 VDD.n934 GND 0.01fF
C1430 VDD.n935 GND 0.02fF
C1431 VDD.n936 GND 0.02fF
C1432 VDD.n937 GND 0.11fF
C1433 VDD.n938 GND 0.02fF
C1434 VDD.n939 GND 0.14fF
C1435 VDD.n940 GND 0.16fF
C1436 VDD.n941 GND 0.01fF
C1437 VDD.n942 GND 0.02fF
C1438 VDD.n943 GND 0.02fF
C1439 VDD.n944 GND 0.18fF
C1440 VDD.n945 GND 0.15fF
C1441 VDD.n946 GND 0.01fF
C1442 VDD.n947 GND 0.02fF
C1443 VDD.n948 GND 0.03fF
C1444 VDD.n949 GND 0.18fF
C1445 VDD.n950 GND 0.14fF
C1446 VDD.n951 GND 0.01fF
C1447 VDD.n952 GND 0.02fF
C1448 VDD.n953 GND 0.03fF
C1449 VDD.n954 GND 0.14fF
C1450 VDD.n955 GND 0.16fF
C1451 VDD.n956 GND 0.01fF
C1452 VDD.n957 GND 0.11fF
C1453 VDD.n958 GND 0.02fF
C1454 VDD.n959 GND 0.02fF
C1455 VDD.n960 GND 0.02fF
C1456 VDD.n961 GND 0.14fF
C1457 VDD.n962 GND 0.17fF
C1458 VDD.n963 GND 0.01fF
C1459 VDD.n964 GND 0.02fF
C1460 VDD.n965 GND 0.02fF
C1461 VDD.n966 GND 0.22fF
C1462 VDD.n967 GND 0.01fF
C1463 VDD.n968 GND 0.07fF
C1464 VDD.n969 GND 0.02fF
C1465 VDD.n970 GND 0.27fF
C1466 VDD.n971 GND 0.01fF
C1467 VDD.n972 GND 0.02fF
C1468 VDD.n973 GND 0.02fF
C1469 VDD.n974 GND 0.27fF
C1470 VDD.n975 GND 0.01fF
C1471 VDD.n976 GND 0.02fF
C1472 VDD.n977 GND 0.03fF
C1473 VDD.n978 GND 0.02fF
C1474 VDD.n979 GND 0.02fF
C1475 VDD.n980 GND 0.02fF
C1476 VDD.n981 GND 0.26fF
C1477 VDD.n982 GND 0.04fF
C1478 VDD.n983 GND 0.03fF
C1479 VDD.n984 GND 0.02fF
C1480 VDD.n985 GND 0.02fF
C1481 VDD.n986 GND 0.02fF
C1482 VDD.n987 GND 0.03fF
C1483 VDD.n988 GND 0.02fF
C1484 VDD.n990 GND 0.02fF
C1485 VDD.n991 GND 0.02fF
C1486 VDD.n992 GND 0.02fF
C1487 VDD.n994 GND 0.27fF
C1488 VDD.n996 GND 0.02fF
C1489 VDD.n997 GND 0.02fF
C1490 VDD.n998 GND 0.03fF
C1491 VDD.n999 GND 0.02fF
C1492 VDD.n1000 GND 0.27fF
C1493 VDD.n1001 GND 0.01fF
C1494 VDD.n1002 GND 0.02fF
C1495 VDD.n1003 GND 0.03fF
C1496 VDD.n1004 GND 0.06fF
C1497 VDD.n1005 GND 0.25fF
C1498 VDD.n1006 GND 0.01fF
C1499 VDD.n1007 GND 0.01fF
C1500 VDD.n1008 GND 0.02fF
C1501 VDD.n1009 GND 0.14fF
C1502 VDD.n1010 GND 0.16fF
C1503 VDD.n1011 GND 0.01fF
C1504 VDD.n1012 GND 0.02fF
C1505 VDD.n1013 GND 0.02fF
C1506 VDD.n1014 GND 0.17fF
C1507 VDD.n1015 GND 0.14fF
C1508 VDD.n1016 GND 0.01fF
C1509 VDD.n1017 GND 0.02fF
C1510 VDD.n1018 GND 0.03fF
C1511 VDD.n1019 GND 0.11fF
C1512 VDD.n1020 GND 0.03fF
C1513 VDD.n1021 GND 0.31fF
C1514 VDD.n1022 GND 0.01fF
C1515 VDD.n1023 GND 0.02fF
C1516 VDD.n1024 GND 0.03fF
C1517 VDD.n1025 GND 0.14fF
C1518 VDD.n1026 GND 0.17fF
C1519 VDD.n1027 GND 0.01fF
C1520 VDD.n1028 GND 0.02fF
C1521 VDD.n1029 GND 0.02fF
C1522 VDD.n1030 GND 0.06fF
C1523 VDD.n1031 GND 0.24fF
C1524 VDD.n1032 GND 0.01fF
C1525 VDD.n1033 GND 0.01fF
C1526 VDD.n1034 GND 0.02fF
C1527 VDD.n1035 GND 0.27fF
C1528 VDD.n1036 GND 0.01fF
C1529 VDD.n1037 GND 0.02fF
C1530 VDD.n1038 GND 0.03fF
C1531 VDD.n1039 GND 0.02fF
C1532 VDD.n1040 GND 0.02fF
C1533 VDD.n1041 GND 0.02fF
C1534 VDD.n1042 GND 0.22fF
C1535 VDD.n1043 GND 0.04fF
C1536 VDD.n1044 GND 0.03fF
C1537 VDD.n1045 GND 0.02fF
C1538 VDD.n1046 GND 0.02fF
C1539 VDD.n1047 GND 0.02fF
C1540 VDD.n1048 GND 0.03fF
C1541 VDD.n1049 GND 0.02fF
C1542 VDD.n1051 GND 0.02fF
C1543 VDD.n1052 GND 0.02fF
C1544 VDD.n1053 GND 0.02fF
C1545 VDD.n1055 GND 0.27fF
C1546 VDD.n1057 GND 0.02fF
C1547 VDD.n1058 GND 0.02fF
C1548 VDD.n1059 GND 0.03fF
C1549 VDD.n1060 GND 0.02fF
C1550 VDD.n1061 GND 0.27fF
C1551 VDD.n1062 GND 0.01fF
C1552 VDD.n1063 GND 0.02fF
C1553 VDD.n1064 GND 0.03fF
C1554 VDD.n1065 GND 0.06fF
C1555 VDD.n1066 GND 0.25fF
C1556 VDD.n1067 GND 0.01fF
C1557 VDD.n1068 GND 0.01fF
C1558 VDD.n1069 GND 0.02fF
C1559 VDD.n1070 GND 0.14fF
C1560 VDD.n1071 GND 0.16fF
C1561 VDD.n1072 GND 0.01fF
C1562 VDD.n1073 GND 0.02fF
C1563 VDD.n1074 GND 0.02fF
C1564 VDD.n1075 GND 0.17fF
C1565 VDD.n1076 GND 0.14fF
C1566 VDD.n1077 GND 0.01fF
C1567 VDD.n1078 GND 0.02fF
C1568 VDD.n1079 GND 0.03fF
C1569 VDD.n1080 GND 0.11fF
C1570 VDD.n1081 GND 0.03fF
C1571 VDD.n1082 GND 0.31fF
C1572 VDD.n1083 GND 0.01fF
C1573 VDD.n1084 GND 0.02fF
C1574 VDD.n1085 GND 0.03fF
C1575 VDD.n1086 GND 0.14fF
C1576 VDD.n1087 GND 0.17fF
C1577 VDD.n1088 GND 0.01fF
C1578 VDD.n1089 GND 0.02fF
C1579 VDD.n1090 GND 0.02fF
C1580 VDD.n1091 GND 0.06fF
C1581 VDD.n1092 GND 0.24fF
C1582 VDD.n1093 GND 0.01fF
C1583 VDD.n1094 GND 0.01fF
C1584 VDD.n1095 GND 0.02fF
C1585 VDD.n1096 GND 0.27fF
C1586 VDD.n1097 GND 0.01fF
C1587 VDD.n1098 GND 0.02fF
C1588 VDD.n1099 GND 0.03fF
C1589 VDD.n1100 GND 0.02fF
C1590 VDD.n1101 GND 0.02fF
C1591 VDD.n1102 GND 0.02fF
C1592 VDD.n1103 GND 0.26fF
C1593 VDD.n1104 GND 0.04fF
C1594 VDD.n1105 GND 0.03fF
C1595 VDD.n1106 GND 0.02fF
C1596 VDD.n1107 GND 0.02fF
C1597 VDD.n1108 GND 0.02fF
C1598 VDD.n1109 GND 0.03fF
C1599 VDD.n1110 GND 0.02fF
C1600 VDD.n1112 GND 0.02fF
C1601 VDD.n1113 GND 0.02fF
C1602 VDD.n1114 GND 0.02fF
C1603 VDD.n1116 GND 0.27fF
C1604 VDD.n1118 GND 0.02fF
C1605 VDD.n1119 GND 0.02fF
C1606 VDD.n1120 GND 0.03fF
C1607 VDD.n1121 GND 0.02fF
C1608 VDD.n1122 GND 0.27fF
C1609 VDD.n1123 GND 0.01fF
C1610 VDD.n1124 GND 0.02fF
C1611 VDD.n1125 GND 0.03fF
C1612 VDD.n1126 GND 0.27fF
C1613 VDD.n1127 GND 0.01fF
C1614 VDD.n1128 GND 0.02fF
C1615 VDD.n1129 GND 0.02fF
C1616 VDD.n1130 GND 0.06fF
C1617 VDD.n1131 GND 0.23fF
C1618 VDD.n1132 GND 0.01fF
C1619 VDD.n1133 GND 0.01fF
C1620 VDD.n1134 GND 0.02fF
C1621 VDD.n1135 GND 0.14fF
C1622 VDD.n1136 GND 0.17fF
C1623 VDD.n1137 GND 0.01fF
C1624 VDD.n1138 GND 0.02fF
C1625 VDD.n1139 GND 0.02fF
C1626 VDD.n1140 GND 0.11fF
C1627 VDD.n1141 GND 0.02fF
C1628 VDD.n1142 GND 0.14fF
C1629 VDD.n1143 GND 0.16fF
C1630 VDD.n1144 GND 0.01fF
C1631 VDD.n1145 GND 0.02fF
C1632 VDD.n1146 GND 0.02fF
C1633 VDD.n1147 GND 0.18fF
C1634 VDD.n1148 GND 0.15fF
C1635 VDD.n1149 GND 0.01fF
C1636 VDD.n1150 GND 0.02fF
C1637 VDD.n1151 GND 0.03fF
C1638 VDD.n1152 GND 0.18fF
C1639 VDD.n1153 GND 0.14fF
C1640 VDD.n1154 GND 0.01fF
C1641 VDD.n1155 GND 0.02fF
C1642 VDD.n1156 GND 0.03fF
C1643 VDD.n1157 GND 0.14fF
C1644 VDD.n1158 GND 0.16fF
C1645 VDD.n1159 GND 0.01fF
C1646 VDD.n1160 GND 0.11fF
C1647 VDD.n1161 GND 0.02fF
C1648 VDD.n1162 GND 0.02fF
C1649 VDD.n1163 GND 0.02fF
C1650 VDD.n1164 GND 0.14fF
C1651 VDD.n1165 GND 0.17fF
C1652 VDD.n1166 GND 0.01fF
C1653 VDD.n1167 GND 0.02fF
C1654 VDD.n1168 GND 0.02fF
C1655 VDD.n1169 GND 0.22fF
C1656 VDD.n1170 GND 0.01fF
C1657 VDD.n1171 GND 0.07fF
C1658 VDD.n1172 GND 0.02fF
C1659 VDD.n1173 GND 0.27fF
C1660 VDD.n1174 GND 0.01fF
C1661 VDD.n1175 GND 0.02fF
C1662 VDD.n1176 GND 0.02fF
C1663 VDD.n1177 GND 0.27fF
C1664 VDD.n1178 GND 0.01fF
C1665 VDD.n1179 GND 0.02fF
C1666 VDD.n1180 GND 0.03fF
C1667 VDD.n1181 GND 0.02fF
C1668 VDD.n1182 GND 0.02fF
C1669 VDD.n1183 GND 0.02fF
C1670 VDD.n1184 GND 0.26fF
C1671 VDD.n1185 GND 0.04fF
C1672 VDD.n1186 GND 0.03fF
C1673 VDD.n1187 GND 0.02fF
C1674 VDD.n1188 GND 0.02fF
C1675 VDD.n1189 GND 0.02fF
C1676 VDD.n1190 GND 0.03fF
C1677 VDD.n1191 GND 0.02fF
C1678 VDD.n1193 GND 0.02fF
C1679 VDD.n1194 GND 0.02fF
C1680 VDD.n1195 GND 0.02fF
C1681 VDD.n1197 GND 0.27fF
C1682 VDD.n1199 GND 0.02fF
C1683 VDD.n1200 GND 0.02fF
C1684 VDD.n1201 GND 0.03fF
C1685 VDD.n1202 GND 0.02fF
C1686 VDD.n1203 GND 0.27fF
C1687 VDD.n1204 GND 0.01fF
C1688 VDD.n1205 GND 0.02fF
C1689 VDD.n1206 GND 0.03fF
C1690 VDD.n1207 GND 0.06fF
C1691 VDD.n1208 GND 0.25fF
C1692 VDD.n1209 GND 0.01fF
C1693 VDD.n1210 GND 0.01fF
C1694 VDD.n1211 GND 0.02fF
C1695 VDD.n1212 GND 0.14fF
C1696 VDD.n1213 GND 0.16fF
C1697 VDD.n1214 GND 0.01fF
C1698 VDD.n1215 GND 0.02fF
C1699 VDD.n1216 GND 0.02fF
C1700 VDD.n1217 GND 0.17fF
C1701 VDD.n1218 GND 0.14fF
C1702 VDD.n1219 GND 0.01fF
C1703 VDD.n1220 GND 0.02fF
C1704 VDD.n1221 GND 0.03fF
C1705 VDD.n1222 GND 0.11fF
C1706 VDD.n1223 GND 0.03fF
C1707 VDD.n1224 GND 0.31fF
C1708 VDD.n1225 GND 0.01fF
C1709 VDD.n1226 GND 0.02fF
C1710 VDD.n1227 GND 0.03fF
C1711 VDD.n1228 GND 0.14fF
C1712 VDD.n1229 GND 0.17fF
C1713 VDD.n1230 GND 0.01fF
C1714 VDD.n1231 GND 0.02fF
C1715 VDD.n1232 GND 0.02fF
C1716 VDD.n1233 GND 0.06fF
C1717 VDD.n1234 GND 0.24fF
C1718 VDD.n1235 GND 0.01fF
C1719 VDD.n1236 GND 0.01fF
C1720 VDD.n1237 GND 0.02fF
C1721 VDD.n1238 GND 0.27fF
C1722 VDD.n1239 GND 0.01fF
C1723 VDD.n1240 GND 0.02fF
C1724 VDD.n1241 GND 0.03fF
C1725 VDD.n1242 GND 0.02fF
C1726 VDD.n1243 GND 0.02fF
C1727 VDD.n1244 GND 0.02fF
C1728 VDD.n1245 GND 0.26fF
C1729 VDD.n1246 GND 0.04fF
C1730 VDD.n1247 GND 0.03fF
C1731 VDD.n1248 GND 0.02fF
C1732 VDD.n1249 GND 0.02fF
C1733 VDD.n1250 GND 0.02fF
C1734 VDD.n1251 GND 0.03fF
C1735 VDD.n1252 GND 0.02fF
C1736 VDD.n1254 GND 0.02fF
C1737 VDD.n1255 GND 0.02fF
C1738 VDD.n1256 GND 0.02fF
C1739 VDD.n1258 GND 0.27fF
C1740 VDD.n1260 GND 0.02fF
C1741 VDD.n1261 GND 0.02fF
C1742 VDD.n1262 GND 0.03fF
C1743 VDD.n1263 GND 0.02fF
C1744 VDD.n1264 GND 0.27fF
C1745 VDD.n1265 GND 0.01fF
C1746 VDD.n1266 GND 0.02fF
C1747 VDD.n1267 GND 0.03fF
C1748 VDD.n1268 GND 0.27fF
C1749 VDD.n1269 GND 0.01fF
C1750 VDD.n1270 GND 0.02fF
C1751 VDD.n1271 GND 0.02fF
C1752 VDD.n1272 GND 0.06fF
C1753 VDD.n1273 GND 0.23fF
C1754 VDD.n1274 GND 0.01fF
C1755 VDD.n1275 GND 0.01fF
C1756 VDD.n1276 GND 0.02fF
C1757 VDD.n1277 GND 0.14fF
C1758 VDD.n1278 GND 0.17fF
C1759 VDD.n1279 GND 0.01fF
C1760 VDD.n1280 GND 0.02fF
C1761 VDD.n1281 GND 0.02fF
C1762 VDD.n1282 GND 0.11fF
C1763 VDD.n1283 GND 0.02fF
C1764 VDD.n1284 GND 0.14fF
C1765 VDD.n1285 GND 0.16fF
C1766 VDD.n1286 GND 0.01fF
C1767 VDD.n1287 GND 0.02fF
C1768 VDD.n1288 GND 0.02fF
C1769 VDD.n1289 GND 0.18fF
C1770 VDD.n1290 GND 0.15fF
C1771 VDD.n1291 GND 0.01fF
C1772 VDD.n1292 GND 0.02fF
C1773 VDD.n1293 GND 0.03fF
C1774 VDD.n1294 GND 0.18fF
C1775 VDD.n1295 GND 0.14fF
C1776 VDD.n1296 GND 0.01fF
C1777 VDD.n1297 GND 0.02fF
C1778 VDD.n1298 GND 0.03fF
C1779 VDD.n1299 GND 0.14fF
C1780 VDD.n1300 GND 0.16fF
C1781 VDD.n1301 GND 0.01fF
C1782 VDD.n1302 GND 0.11fF
C1783 VDD.n1303 GND 0.02fF
C1784 VDD.n1304 GND 0.02fF
C1785 VDD.n1305 GND 0.02fF
C1786 VDD.n1306 GND 0.14fF
C1787 VDD.n1307 GND 0.17fF
C1788 VDD.n1308 GND 0.01fF
C1789 VDD.n1309 GND 0.02fF
C1790 VDD.n1310 GND 0.02fF
C1791 VDD.n1311 GND 0.22fF
C1792 VDD.n1312 GND 0.01fF
C1793 VDD.n1313 GND 0.07fF
C1794 VDD.n1314 GND 0.02fF
C1795 VDD.n1315 GND 0.27fF
C1796 VDD.n1316 GND 0.01fF
C1797 VDD.n1317 GND 0.02fF
C1798 VDD.n1318 GND 0.02fF
C1799 VDD.n1319 GND 0.27fF
C1800 VDD.n1320 GND 0.01fF
C1801 VDD.n1321 GND 0.02fF
C1802 VDD.n1322 GND 0.03fF
C1803 VDD.n1323 GND 0.02fF
C1804 VDD.n1324 GND 0.02fF
C1805 VDD.n1325 GND 0.02fF
C1806 VDD.n1326 GND 0.31fF
C1807 VDD.n1327 GND 0.04fF
C1808 VDD.n1328 GND 0.03fF
C1809 VDD.n1329 GND 0.02fF
C1810 VDD.n1330 GND 0.02fF
C1811 VDD.n1331 GND 0.02fF
C1812 VDD.n1332 GND 0.03fF
C1813 VDD.n1333 GND 0.02fF
C1814 VDD.n1335 GND 0.02fF
C1815 VDD.n1336 GND 0.02fF
C1816 VDD.n1337 GND 0.02fF
C1817 VDD.n1339 GND 0.27fF
C1818 VDD.n1341 GND 0.02fF
C1819 VDD.n1342 GND 0.02fF
C1820 VDD.n1343 GND 0.03fF
C1821 VDD.n1344 GND 0.02fF
C1822 VDD.n1345 GND 0.27fF
C1823 VDD.n1346 GND 0.01fF
C1824 VDD.n1347 GND 0.02fF
C1825 VDD.n1348 GND 0.03fF
C1826 VDD.n1349 GND 0.27fF
C1827 VDD.n1350 GND 0.01fF
C1828 VDD.n1351 GND 0.02fF
C1829 VDD.n1352 GND 0.02fF
C1830 VDD.n1353 GND 0.06fF
C1831 VDD.n1354 GND 0.23fF
C1832 VDD.n1355 GND 0.01fF
C1833 VDD.n1356 GND 0.01fF
C1834 VDD.n1357 GND 0.02fF
C1835 VDD.n1358 GND 0.14fF
C1836 VDD.n1359 GND 0.17fF
C1837 VDD.n1360 GND 0.01fF
C1838 VDD.n1361 GND 0.02fF
C1839 VDD.n1362 GND 0.02fF
C1840 VDD.n1363 GND 0.11fF
C1841 VDD.n1364 GND 0.02fF
C1842 VDD.n1365 GND 0.14fF
C1843 VDD.n1366 GND 0.16fF
C1844 VDD.n1367 GND 0.01fF
C1845 VDD.n1368 GND 0.02fF
C1846 VDD.n1369 GND 0.02fF
C1847 VDD.n1370 GND 0.18fF
C1848 VDD.n1371 GND 0.15fF
C1849 VDD.n1372 GND 0.01fF
C1850 VDD.n1373 GND 0.02fF
C1851 VDD.n1374 GND 0.03fF
C1852 VDD.n1375 GND 0.18fF
C1853 VDD.n1376 GND 0.14fF
C1854 VDD.n1377 GND 0.01fF
C1855 VDD.n1378 GND 0.02fF
C1856 VDD.n1379 GND 0.03fF
C1857 VDD.n1380 GND 0.14fF
C1858 VDD.n1381 GND 0.16fF
C1859 VDD.n1382 GND 0.01fF
C1860 VDD.n1383 GND 0.11fF
C1861 VDD.n1384 GND 0.02fF
C1862 VDD.n1385 GND 0.02fF
C1863 VDD.n1386 GND 0.02fF
C1864 VDD.n1387 GND 0.14fF
C1865 VDD.n1388 GND 0.17fF
C1866 VDD.n1389 GND 0.01fF
C1867 VDD.n1390 GND 0.02fF
C1868 VDD.n1391 GND 0.02fF
C1869 VDD.n1392 GND 0.22fF
C1870 VDD.n1393 GND 0.01fF
C1871 VDD.n1394 GND 0.07fF
C1872 VDD.n1395 GND 0.02fF
C1873 VDD.n1396 GND 0.27fF
C1874 VDD.n1397 GND 0.01fF
C1875 VDD.n1398 GND 0.02fF
C1876 VDD.n1399 GND 0.02fF
C1877 VDD.n1400 GND 0.27fF
C1878 VDD.n1401 GND 0.01fF
C1879 VDD.n1402 GND 0.02fF
C1880 VDD.n1403 GND 0.03fF
C1881 VDD.n1404 GND 0.02fF
C1882 VDD.n1405 GND 0.02fF
C1883 VDD.n1406 GND 0.02fF
C1884 VDD.n1407 GND 0.26fF
C1885 VDD.n1408 GND 0.04fF
C1886 VDD.n1409 GND 0.03fF
C1887 VDD.n1410 GND 0.02fF
C1888 VDD.n1411 GND 0.02fF
C1889 VDD.n1412 GND 0.02fF
C1890 VDD.n1413 GND 0.03fF
C1891 VDD.n1414 GND 0.02fF
C1892 VDD.n1416 GND 0.02fF
C1893 VDD.n1417 GND 0.02fF
C1894 VDD.n1418 GND 0.02fF
C1895 VDD.n1420 GND 0.27fF
C1896 VDD.n1422 GND 0.02fF
C1897 VDD.n1423 GND 0.02fF
C1898 VDD.n1424 GND 0.03fF
C1899 VDD.n1425 GND 0.02fF
C1900 VDD.n1426 GND 0.27fF
C1901 VDD.n1427 GND 0.01fF
C1902 VDD.n1428 GND 0.02fF
C1903 VDD.n1429 GND 0.03fF
C1904 VDD.n1430 GND 0.06fF
C1905 VDD.n1431 GND 0.25fF
C1906 VDD.n1432 GND 0.01fF
C1907 VDD.n1433 GND 0.01fF
C1908 VDD.n1434 GND 0.02fF
C1909 VDD.n1435 GND 0.14fF
C1910 VDD.n1436 GND 0.16fF
C1911 VDD.n1437 GND 0.01fF
C1912 VDD.n1438 GND 0.02fF
C1913 VDD.n1439 GND 0.02fF
C1914 VDD.n1440 GND 0.17fF
C1915 VDD.n1441 GND 0.14fF
C1916 VDD.n1442 GND 0.01fF
C1917 VDD.n1443 GND 0.02fF
C1918 VDD.n1444 GND 0.03fF
C1919 VDD.n1445 GND 0.11fF
C1920 VDD.n1446 GND 0.03fF
C1921 VDD.n1447 GND 0.31fF
C1922 VDD.n1448 GND 0.01fF
C1923 VDD.n1449 GND 0.02fF
C1924 VDD.n1450 GND 0.03fF
C1925 VDD.n1451 GND 0.14fF
C1926 VDD.n1452 GND 0.17fF
C1927 VDD.n1453 GND 0.01fF
C1928 VDD.n1454 GND 0.02fF
C1929 VDD.n1455 GND 0.02fF
C1930 VDD.n1456 GND 0.06fF
C1931 VDD.n1457 GND 0.24fF
C1932 VDD.n1458 GND 0.01fF
C1933 VDD.n1459 GND 0.01fF
C1934 VDD.n1460 GND 0.02fF
C1935 VDD.n1461 GND 0.27fF
C1936 VDD.n1462 GND 0.01fF
C1937 VDD.n1463 GND 0.02fF
C1938 VDD.n1464 GND 0.03fF
C1939 VDD.n1465 GND 0.02fF
C1940 VDD.n1466 GND 0.02fF
C1941 VDD.n1467 GND 0.02fF
C1942 VDD.n1468 GND 0.22fF
C1943 VDD.n1469 GND 0.04fF
C1944 VDD.n1470 GND 0.03fF
C1945 VDD.n1471 GND 0.02fF
C1946 VDD.n1472 GND 0.02fF
C1947 VDD.n1473 GND 0.02fF
C1948 VDD.n1474 GND 0.03fF
C1949 VDD.n1475 GND 0.02fF
C1950 VDD.n1477 GND 0.02fF
C1951 VDD.n1478 GND 0.02fF
C1952 VDD.n1479 GND 0.02fF
C1953 VDD.n1481 GND 0.27fF
C1954 VDD.n1483 GND 0.02fF
C1955 VDD.n1484 GND 0.02fF
C1956 VDD.n1485 GND 0.03fF
C1957 VDD.n1486 GND 0.02fF
C1958 VDD.n1487 GND 0.27fF
C1959 VDD.n1488 GND 0.01fF
C1960 VDD.n1489 GND 0.02fF
C1961 VDD.n1490 GND 0.03fF
C1962 VDD.n1491 GND 0.06fF
C1963 VDD.n1492 GND 0.25fF
C1964 VDD.n1493 GND 0.01fF
C1965 VDD.n1494 GND 0.01fF
C1966 VDD.n1495 GND 0.02fF
C1967 VDD.n1496 GND 0.14fF
C1968 VDD.n1497 GND 0.16fF
C1969 VDD.n1498 GND 0.01fF
C1970 VDD.n1499 GND 0.02fF
C1971 VDD.n1500 GND 0.02fF
C1972 VDD.n1501 GND 0.17fF
C1973 VDD.n1502 GND 0.14fF
C1974 VDD.n1503 GND 0.01fF
C1975 VDD.n1504 GND 0.02fF
C1976 VDD.n1505 GND 0.03fF
C1977 VDD.n1506 GND 0.11fF
C1978 VDD.n1507 GND 0.03fF
C1979 VDD.n1508 GND 0.31fF
C1980 VDD.n1509 GND 0.01fF
C1981 VDD.n1510 GND 0.02fF
C1982 VDD.n1511 GND 0.02fF
C1983 a_8483_411.n0 GND 0.08fF
C1984 a_8483_411.n1 GND 1.05fF
C1985 a_8483_411.n2 GND 1.05fF
C1986 a_8483_411.n3 GND 1.23fF
C1987 a_8483_411.n4 GND 0.39fF
C1988 a_8483_411.n5 GND 0.60fF
C1989 a_8483_411.n6 GND 0.54fF
C1990 a_8483_411.n7 GND 1.45fF
C1991 a_8483_411.n8 GND 0.48fF
C1992 a_8483_411.n9 GND 1.04fF
C1993 a_8483_411.n10 GND 1.55fF
C1994 a_8483_411.n11 GND 0.66fF
C1995 a_8483_411.t15 GND 1.04fF
C1996 a_8483_411.n12 GND 0.79fF
C1997 a_8483_411.n13 GND 9.28fF
C1998 a_8483_411.n14 GND 0.88fF
C1999 a_8483_411.n15 GND 0.08fF
C2000 a_8483_411.n16 GND 0.59fF
C2001 a_8483_411.n17 GND 0.09fF
.ends
