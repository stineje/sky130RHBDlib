// File: TMRDFFSNQNX1.spi.pex
// Created: Tue Oct 15 15:52:31 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_TMRDFFSNQNX1\%GND ( 1 139 143 146 151 159 165 175 181 191 197 203 \
 211 219 227 237 245 253 259 269 275 285 291 297 305 313 321 331 339 347 353 \
 363 369 379 385 391 399 407 415 425 433 441 447 453 466 470 473 476 479 481 \
 483 485 488 491 494 496 498 500 503 506 509 511 513 515 518 520 521 522 523 \
 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 )
c976 ( 540 0 ) capacitor c=0.0215012f //x=80.91 //y=0.865
c977 ( 539 0 ) capacitor c=0.0215012f //x=77.58 //y=0.865
c978 ( 538 0 ) capacitor c=0.0207524f //x=74.25 //y=0.865
c979 ( 537 0 ) capacitor c=0.0226075f //x=69.335 //y=0.875
c980 ( 536 0 ) capacitor c=0.0207407f //x=66.11 //y=0.865
c981 ( 535 0 ) capacitor c=0.0207407f //x=62.78 //y=0.865
c982 ( 534 0 ) capacitor c=0.0225954f //x=57.865 //y=0.875
c983 ( 533 0 ) capacitor c=0.0226075f //x=53.055 //y=0.875
c984 ( 532 0 ) capacitor c=0.0207407f //x=49.83 //y=0.865
c985 ( 531 0 ) capacitor c=0.0226075f //x=44.915 //y=0.875
c986 ( 530 0 ) capacitor c=0.0207407f //x=41.69 //y=0.865
c987 ( 529 0 ) capacitor c=0.0207407f //x=38.36 //y=0.865
c988 ( 528 0 ) capacitor c=0.0225954f //x=33.445 //y=0.875
c989 ( 527 0 ) capacitor c=0.0226075f //x=28.635 //y=0.875
c990 ( 526 0 ) capacitor c=0.0207407f //x=25.41 //y=0.865
c991 ( 525 0 ) capacitor c=0.0226075f //x=20.495 //y=0.875
c992 ( 524 0 ) capacitor c=0.0207407f //x=17.27 //y=0.865
c993 ( 523 0 ) capacitor c=0.0207407f //x=13.94 //y=0.865
c994 ( 522 0 ) capacitor c=0.0226205f //x=9.025 //y=0.875
c995 ( 521 0 ) capacitor c=0.0226323f //x=4.215 //y=0.875
c996 ( 520 0 ) capacitor c=0.0207863f //x=0.99 //y=0.865
c997 ( 519 0 ) capacitor c=0.00440095f //x=81.1 //y=0
c998 ( 518 0 ) capacitor c=0.101477f //x=79.92 //y=0
c999 ( 517 0 ) capacitor c=0.00440095f //x=77.7 //y=0
c1000 ( 515 0 ) capacitor c=0.116995f //x=76.59 //y=0
c1001 ( 514 0 ) capacitor c=0.00440095f //x=74.44 //y=0
c1002 ( 513 0 ) capacitor c=0.106826f //x=73.26 //y=0
c1003 ( 512 0 ) capacitor c=0.00440144f //x=69.525 //y=0
c1004 ( 511 0 ) capacitor c=0.104091f //x=68.45 //y=0
c1005 ( 510 0 ) capacitor c=0.00440095f //x=66.3 //y=0
c1006 ( 509 0 ) capacitor c=0.105123f //x=65.12 //y=0
c1007 ( 508 0 ) capacitor c=0.00440095f //x=62.9 //y=0
c1008 ( 506 0 ) capacitor c=0.108248f //x=61.79 //y=0
c1009 ( 505 0 ) capacitor c=0.00440144f //x=58.09 //y=0
c1010 ( 503 0 ) capacitor c=0.107229f //x=56.98 //y=0
c1011 ( 502 0 ) capacitor c=0.00440144f //x=53.28 //y=0
c1012 ( 500 0 ) capacitor c=0.104113f //x=52.17 //y=0
c1013 ( 499 0 ) capacitor c=0.00440095f //x=50.02 //y=0
c1014 ( 498 0 ) capacitor c=0.108568f //x=48.84 //y=0
c1015 ( 497 0 ) capacitor c=0.00440144f //x=45.105 //y=0
c1016 ( 496 0 ) capacitor c=0.10408f //x=44.03 //y=0
c1017 ( 495 0 ) capacitor c=0.00440095f //x=41.88 //y=0
c1018 ( 494 0 ) capacitor c=0.104882f //x=40.7 //y=0
c1019 ( 493 0 ) capacitor c=0.00440095f //x=38.48 //y=0
c1020 ( 491 0 ) capacitor c=0.108248f //x=37.37 //y=0
c1021 ( 490 0 ) capacitor c=0.00440144f //x=33.67 //y=0
c1022 ( 488 0 ) capacitor c=0.107229f //x=32.56 //y=0
c1023 ( 487 0 ) capacitor c=0.00440144f //x=28.86 //y=0
c1024 ( 485 0 ) capacitor c=0.104143f //x=27.75 //y=0
c1025 ( 484 0 ) capacitor c=0.00440095f //x=25.6 //y=0
c1026 ( 483 0 ) capacitor c=0.108018f //x=24.42 //y=0
c1027 ( 482 0 ) capacitor c=0.00440144f //x=20.685 //y=0
c1028 ( 481 0 ) capacitor c=0.104091f //x=19.61 //y=0
c1029 ( 480 0 ) capacitor c=0.00440095f //x=17.46 //y=0
c1030 ( 479 0 ) capacitor c=0.105123f //x=16.28 //y=0
c1031 ( 478 0 ) capacitor c=0.00440095f //x=14.06 //y=0
c1032 ( 476 0 ) capacitor c=0.108248f //x=12.95 //y=0
c1033 ( 475 0 ) capacitor c=0.00440144f //x=9.25 //y=0
c1034 ( 473 0 ) capacitor c=0.108235f //x=8.14 //y=0
c1035 ( 472 0 ) capacitor c=0.00440144f //x=4.44 //y=0
c1036 ( 470 0 ) capacitor c=0.105313f //x=3.33 //y=0
c1037 ( 469 0 ) capacitor c=0.00440095f //x=1.18 //y=0
c1038 ( 466 0 ) capacitor c=0.258637f //x=82.51 //y=0
c1039 ( 453 0 ) capacitor c=0.0389876f //x=81.015 //y=0
c1040 ( 447 0 ) capacitor c=0.0716428f //x=79.75 //y=0
c1041 ( 441 0 ) capacitor c=0.0388276f //x=77.685 //y=0
c1042 ( 433 0 ) capacitor c=0.071962f //x=76.42 //y=0
c1043 ( 425 0 ) capacitor c=0.0391432f //x=74.355 //y=0
c1044 ( 415 0 ) capacitor c=0.133607f //x=73.09 //y=0
c1045 ( 407 0 ) capacitor c=0.0339325f //x=69.44 //y=0
c1046 ( 399 0 ) capacitor c=0.0718026f //x=68.28 //y=0
c1047 ( 391 0 ) capacitor c=0.0388888f //x=66.215 //y=0
c1048 ( 385 0 ) capacitor c=0.0718026f //x=64.95 //y=0
c1049 ( 379 0 ) capacitor c=0.0388888f //x=62.885 //y=0
c1050 ( 369 0 ) capacitor c=0.133362f //x=61.62 //y=0
c1051 ( 363 0 ) capacitor c=0.0339325f //x=57.97 //y=0
c1052 ( 353 0 ) capacitor c=0.133362f //x=56.81 //y=0
c1053 ( 347 0 ) capacitor c=0.0339325f //x=53.16 //y=0
c1054 ( 339 0 ) capacitor c=0.0718026f //x=52 //y=0
c1055 ( 331 0 ) capacitor c=0.0388888f //x=49.935 //y=0
c1056 ( 321 0 ) capacitor c=0.133362f //x=48.67 //y=0
c1057 ( 313 0 ) capacitor c=0.0339325f //x=45.02 //y=0
c1058 ( 305 0 ) capacitor c=0.0718026f //x=43.86 //y=0
c1059 ( 297 0 ) capacitor c=0.0388888f //x=41.795 //y=0
c1060 ( 291 0 ) capacitor c=0.0718026f //x=40.53 //y=0
c1061 ( 285 0 ) capacitor c=0.0388888f //x=38.465 //y=0
c1062 ( 275 0 ) capacitor c=0.133362f //x=37.2 //y=0
c1063 ( 269 0 ) capacitor c=0.0339325f //x=33.55 //y=0
c1064 ( 259 0 ) capacitor c=0.133362f //x=32.39 //y=0
c1065 ( 253 0 ) capacitor c=0.0339325f //x=28.74 //y=0
c1066 ( 245 0 ) capacitor c=0.0718026f //x=27.58 //y=0
c1067 ( 237 0 ) capacitor c=0.0388888f //x=25.515 //y=0
c1068 ( 227 0 ) capacitor c=0.133362f //x=24.25 //y=0
c1069 ( 219 0 ) capacitor c=0.0339325f //x=20.6 //y=0
c1070 ( 211 0 ) capacitor c=0.0718026f //x=19.44 //y=0
c1071 ( 203 0 ) capacitor c=0.0388888f //x=17.375 //y=0
c1072 ( 197 0 ) capacitor c=0.0718026f //x=16.11 //y=0
c1073 ( 191 0 ) capacitor c=0.0388888f //x=14.045 //y=0
c1074 ( 181 0 ) capacitor c=0.133404f //x=12.78 //y=0
c1075 ( 175 0 ) capacitor c=0.0339482f //x=9.13 //y=0
c1076 ( 165 0 ) capacitor c=0.133515f //x=7.97 //y=0
c1077 ( 159 0 ) capacitor c=0.0339482f //x=4.32 //y=0
c1078 ( 151 0 ) capacitor c=0.0720441f //x=3.16 //y=0
c1079 ( 146 0 ) capacitor c=0.179262f //x=0.74 //y=0
c1080 ( 143 0 ) capacitor c=0.0426751f //x=1.095 //y=0
c1081 ( 139 0 ) capacitor c=2.51766f //x=82.51 //y=0
r1082 (  464 466 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=81.4 //y=0 //x2=82.51 //y2=0
r1083 (  462 519 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.185 //y=0 //x2=81.1 //y2=0
r1084 (  462 464 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=81.185 //y=0 //x2=81.4 //y2=0
r1085 (  457 519 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.1 //y=0.17 //x2=81.1 //y2=0
r1086 (  457 540 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=81.1 //y=0.17 //x2=81.1 //y2=0.955
r1087 (  454 518 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=80.09 //y=0 //x2=79.92 //y2=0
r1088 (  454 456 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=80.09 //y=0 //x2=80.29 //y2=0
r1089 (  453 519 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.015 //y=0 //x2=81.1 //y2=0
r1090 (  453 456 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=81.015 //y=0 //x2=80.29 //y2=0
r1091 (  448 517 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.855 //y=0 //x2=77.77 //y2=0
r1092 (  448 450 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=77.855 //y=0 //x2=78.81 //y2=0
r1093 (  447 518 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=79.75 //y=0 //x2=79.92 //y2=0
r1094 (  447 450 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=79.75 //y=0 //x2=78.81 //y2=0
r1095 (  443 517 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.77 //y=0.17 //x2=77.77 //y2=0
r1096 (  443 539 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=77.77 //y=0.17 //x2=77.77 //y2=0.955
r1097 (  442 515 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.76 //y=0 //x2=76.59 //y2=0
r1098 (  441 517 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.685 //y=0 //x2=77.77 //y2=0
r1099 (  441 442 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=77.685 //y=0 //x2=76.76 //y2=0
r1100 (  436 438 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=75.11 //y=0 //x2=76.22 //y2=0
r1101 (  434 514 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.525 //y=0 //x2=74.44 //y2=0
r1102 (  434 436 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=74.525 //y=0 //x2=75.11 //y2=0
r1103 (  433 515 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.42 //y=0 //x2=76.59 //y2=0
r1104 (  433 438 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=76.42 //y=0 //x2=76.22 //y2=0
r1105 (  429 514 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.44 //y=0.17 //x2=74.44 //y2=0
r1106 (  429 538 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=74.44 //y=0.17 //x2=74.44 //y2=0.955
r1107 (  426 513 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.43 //y=0 //x2=73.26 //y2=0
r1108 (  426 428 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=73.43 //y=0 //x2=74 //y2=0
r1109 (  425 514 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.355 //y=0 //x2=74.44 //y2=0
r1110 (  425 428 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=74.355 //y=0 //x2=74 //y2=0
r1111 (  420 422 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=71.41 //y=0 //x2=72.52 //y2=0
r1112 (  418 420 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=70.3 //y=0 //x2=71.41 //y2=0
r1113 (  416 512 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.61 //y=0 //x2=69.525 //y2=0
r1114 (  416 418 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=69.61 //y=0 //x2=70.3 //y2=0
r1115 (  415 513 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.09 //y=0 //x2=73.26 //y2=0
r1116 (  415 422 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=73.09 //y=0 //x2=72.52 //y2=0
r1117 (  411 512 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.525 //y=0.17 //x2=69.525 //y2=0
r1118 (  411 537 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=69.525 //y=0.17 //x2=69.525 //y2=0.965
r1119 (  408 511 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.62 //y=0 //x2=68.45 //y2=0
r1120 (  408 410 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=68.62 //y=0 //x2=69.19 //y2=0
r1121 (  407 512 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.44 //y=0 //x2=69.525 //y2=0
r1122 (  407 410 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=69.44 //y=0 //x2=69.19 //y2=0
r1123 (  402 404 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=66.6 //y=0 //x2=67.71 //y2=0
r1124 (  400 510 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.385 //y=0 //x2=66.3 //y2=0
r1125 (  400 402 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=66.385 //y=0 //x2=66.6 //y2=0
r1126 (  399 511 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.28 //y=0 //x2=68.45 //y2=0
r1127 (  399 404 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=68.28 //y=0 //x2=67.71 //y2=0
r1128 (  395 510 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=66.3 //y=0.17 //x2=66.3 //y2=0
r1129 (  395 536 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=66.3 //y=0.17 //x2=66.3 //y2=0.955
r1130 (  392 509 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.29 //y=0 //x2=65.12 //y2=0
r1131 (  392 394 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=65.29 //y=0 //x2=65.49 //y2=0
r1132 (  391 510 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.215 //y=0 //x2=66.3 //y2=0
r1133 (  391 394 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=66.215 //y=0 //x2=65.49 //y2=0
r1134 (  386 508 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.055 //y=0 //x2=62.97 //y2=0
r1135 (  386 388 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=63.055 //y=0 //x2=64.01 //y2=0
r1136 (  385 509 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.95 //y=0 //x2=65.12 //y2=0
r1137 (  385 388 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=64.95 //y=0 //x2=64.01 //y2=0
r1138 (  381 508 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.97 //y=0.17 //x2=62.97 //y2=0
r1139 (  381 535 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=62.97 //y=0.17 //x2=62.97 //y2=0.955
r1140 (  380 506 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.96 //y=0 //x2=61.79 //y2=0
r1141 (  379 508 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.885 //y=0 //x2=62.97 //y2=0
r1142 (  379 380 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=62.885 //y=0 //x2=61.96 //y2=0
r1143 (  374 376 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=60.31 //y=0 //x2=61.42 //y2=0
r1144 (  372 374 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=59.2 //y=0 //x2=60.31 //y2=0
r1145 (  370 505 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.14 //y=0 //x2=58.055 //y2=0
r1146 (  370 372 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=58.14 //y=0 //x2=59.2 //y2=0
r1147 (  369 506 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.62 //y=0 //x2=61.79 //y2=0
r1148 (  369 376 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=61.62 //y=0 //x2=61.42 //y2=0
r1149 (  365 505 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.055 //y=0.17 //x2=58.055 //y2=0
r1150 (  365 534 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=58.055 //y=0.17 //x2=58.055 //y2=0.965
r1151 (  364 503 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.15 //y=0 //x2=56.98 //y2=0
r1152 (  363 505 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=57.97 //y=0 //x2=58.055 //y2=0
r1153 (  363 364 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=57.97 //y=0 //x2=57.15 //y2=0
r1154 (  358 360 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=55.5 //y=0 //x2=56.61 //y2=0
r1155 (  356 358 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=54.39 //y=0 //x2=55.5 //y2=0
r1156 (  354 502 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.33 //y=0 //x2=53.245 //y2=0
r1157 (  354 356 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=53.33 //y=0 //x2=54.39 //y2=0
r1158 (  353 503 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.81 //y=0 //x2=56.98 //y2=0
r1159 (  353 360 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=56.81 //y=0 //x2=56.61 //y2=0
r1160 (  349 502 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.245 //y=0.17 //x2=53.245 //y2=0
r1161 (  349 533 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=53.245 //y=0.17 //x2=53.245 //y2=0.965
r1162 (  348 500 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.34 //y=0 //x2=52.17 //y2=0
r1163 (  347 502 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.16 //y=0 //x2=53.245 //y2=0
r1164 (  347 348 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=53.16 //y=0 //x2=52.34 //y2=0
r1165 (  342 344 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=50.69 //y=0 //x2=51.8 //y2=0
r1166 (  340 499 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.105 //y=0 //x2=50.02 //y2=0
r1167 (  340 342 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=50.105 //y=0 //x2=50.69 //y2=0
r1168 (  339 500 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52 //y=0 //x2=52.17 //y2=0
r1169 (  339 344 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=52 //y=0 //x2=51.8 //y2=0
r1170 (  335 499 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.02 //y=0.17 //x2=50.02 //y2=0
r1171 (  335 532 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=50.02 //y=0.17 //x2=50.02 //y2=0.955
r1172 (  332 498 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.01 //y=0 //x2=48.84 //y2=0
r1173 (  332 334 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=49.01 //y=0 //x2=49.58 //y2=0
r1174 (  331 499 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.935 //y=0 //x2=50.02 //y2=0
r1175 (  331 334 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=49.935 //y=0 //x2=49.58 //y2=0
r1176 (  326 328 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=46.99 //y=0 //x2=48.1 //y2=0
r1177 (  324 326 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=45.88 //y=0 //x2=46.99 //y2=0
r1178 (  322 497 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.19 //y=0 //x2=45.105 //y2=0
r1179 (  322 324 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=45.19 //y=0 //x2=45.88 //y2=0
r1180 (  321 498 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.67 //y=0 //x2=48.84 //y2=0
r1181 (  321 328 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.67 //y=0 //x2=48.1 //y2=0
r1182 (  317 497 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=45.105 //y=0.17 //x2=45.105 //y2=0
r1183 (  317 531 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=45.105 //y=0.17 //x2=45.105 //y2=0.965
r1184 (  314 496 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.2 //y=0 //x2=44.03 //y2=0
r1185 (  314 316 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=44.2 //y=0 //x2=44.77 //y2=0
r1186 (  313 497 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.02 //y=0 //x2=45.105 //y2=0
r1187 (  313 316 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=45.02 //y=0 //x2=44.77 //y2=0
r1188 (  308 310 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=42.18 //y=0 //x2=43.29 //y2=0
r1189 (  306 495 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.965 //y=0 //x2=41.88 //y2=0
r1190 (  306 308 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=41.965 //y=0 //x2=42.18 //y2=0
r1191 (  305 496 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.86 //y=0 //x2=44.03 //y2=0
r1192 (  305 310 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.86 //y=0 //x2=43.29 //y2=0
r1193 (  301 495 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=41.88 //y=0.17 //x2=41.88 //y2=0
r1194 (  301 530 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=41.88 //y=0.17 //x2=41.88 //y2=0.955
r1195 (  298 494 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.87 //y=0 //x2=40.7 //y2=0
r1196 (  298 300 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=40.87 //y=0 //x2=41.07 //y2=0
r1197 (  297 495 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.795 //y=0 //x2=41.88 //y2=0
r1198 (  297 300 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=41.795 //y=0 //x2=41.07 //y2=0
r1199 (  292 493 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.635 //y=0 //x2=38.55 //y2=0
r1200 (  292 294 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=38.635 //y=0 //x2=39.59 //y2=0
r1201 (  291 494 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.53 //y=0 //x2=40.7 //y2=0
r1202 (  291 294 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=40.53 //y=0 //x2=39.59 //y2=0
r1203 (  287 493 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.55 //y=0.17 //x2=38.55 //y2=0
r1204 (  287 529 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=38.55 //y=0.17 //x2=38.55 //y2=0.955
r1205 (  286 491 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.54 //y=0 //x2=37.37 //y2=0
r1206 (  285 493 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.465 //y=0 //x2=38.55 //y2=0
r1207 (  285 286 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=38.465 //y=0 //x2=37.54 //y2=0
r1208 (  280 282 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=35.89 //y=0 //x2=37 //y2=0
r1209 (  278 280 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=34.78 //y=0 //x2=35.89 //y2=0
r1210 (  276 490 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.72 //y=0 //x2=33.635 //y2=0
r1211 (  276 278 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=33.72 //y=0 //x2=34.78 //y2=0
r1212 (  275 491 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.2 //y=0 //x2=37.37 //y2=0
r1213 (  275 282 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=37.2 //y=0 //x2=37 //y2=0
r1214 (  271 490 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.635 //y=0.17 //x2=33.635 //y2=0
r1215 (  271 528 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=33.635 //y=0.17 //x2=33.635 //y2=0.965
r1216 (  270 488 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.73 //y=0 //x2=32.56 //y2=0
r1217 (  269 490 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.55 //y=0 //x2=33.635 //y2=0
r1218 (  269 270 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=33.55 //y=0 //x2=32.73 //y2=0
r1219 (  264 266 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=31.08 //y=0 //x2=32.19 //y2=0
r1220 (  262 264 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=29.97 //y=0 //x2=31.08 //y2=0
r1221 (  260 487 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.91 //y=0 //x2=28.825 //y2=0
r1222 (  260 262 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=28.91 //y=0 //x2=29.97 //y2=0
r1223 (  259 488 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.39 //y=0 //x2=32.56 //y2=0
r1224 (  259 266 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=32.39 //y=0 //x2=32.19 //y2=0
r1225 (  255 487 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.825 //y=0.17 //x2=28.825 //y2=0
r1226 (  255 527 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=28.825 //y=0.17 //x2=28.825 //y2=0.965
r1227 (  254 485 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.92 //y=0 //x2=27.75 //y2=0
r1228 (  253 487 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.74 //y=0 //x2=28.825 //y2=0
r1229 (  253 254 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=28.74 //y=0 //x2=27.92 //y2=0
r1230 (  248 250 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=26.27 //y=0 //x2=27.38 //y2=0
r1231 (  246 484 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.685 //y=0 //x2=25.6 //y2=0
r1232 (  246 248 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=25.685 //y=0 //x2=26.27 //y2=0
r1233 (  245 485 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.58 //y=0 //x2=27.75 //y2=0
r1234 (  245 250 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=27.58 //y=0 //x2=27.38 //y2=0
r1235 (  241 484 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.6 //y=0.17 //x2=25.6 //y2=0
r1236 (  241 526 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=25.6 //y=0.17 //x2=25.6 //y2=0.955
r1237 (  238 483 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.59 //y=0 //x2=24.42 //y2=0
r1238 (  238 240 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.59 //y=0 //x2=25.16 //y2=0
r1239 (  237 484 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.515 //y=0 //x2=25.6 //y2=0
r1240 (  237 240 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=25.515 //y=0 //x2=25.16 //y2=0
r1241 (  232 234 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=22.57 //y=0 //x2=23.68 //y2=0
r1242 (  230 232 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.46 //y=0 //x2=22.57 //y2=0
r1243 (  228 482 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.77 //y=0 //x2=20.685 //y2=0
r1244 (  228 230 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=20.77 //y=0 //x2=21.46 //y2=0
r1245 (  227 483 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.25 //y=0 //x2=24.42 //y2=0
r1246 (  227 234 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.25 //y=0 //x2=23.68 //y2=0
r1247 (  223 482 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.685 //y=0.17 //x2=20.685 //y2=0
r1248 (  223 525 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=20.685 //y=0.17 //x2=20.685 //y2=0.965
r1249 (  220 481 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.78 //y=0 //x2=19.61 //y2=0
r1250 (  220 222 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.78 //y=0 //x2=20.35 //y2=0
r1251 (  219 482 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.6 //y=0 //x2=20.685 //y2=0
r1252 (  219 222 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=20.6 //y=0 //x2=20.35 //y2=0
r1253 (  214 216 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.76 //y=0 //x2=18.87 //y2=0
r1254 (  212 480 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.545 //y=0 //x2=17.46 //y2=0
r1255 (  212 214 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=17.545 //y=0 //x2=17.76 //y2=0
r1256 (  211 481 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.44 //y=0 //x2=19.61 //y2=0
r1257 (  211 216 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.44 //y=0 //x2=18.87 //y2=0
r1258 (  207 480 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.46 //y=0.17 //x2=17.46 //y2=0
r1259 (  207 524 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=17.46 //y=0.17 //x2=17.46 //y2=0.955
r1260 (  204 479 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.45 //y=0 //x2=16.28 //y2=0
r1261 (  204 206 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=16.45 //y=0 //x2=16.65 //y2=0
r1262 (  203 480 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.375 //y=0 //x2=17.46 //y2=0
r1263 (  203 206 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=17.375 //y=0 //x2=16.65 //y2=0
r1264 (  198 478 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.215 //y=0 //x2=14.13 //y2=0
r1265 (  198 200 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=14.215 //y=0 //x2=15.17 //y2=0
r1266 (  197 479 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.11 //y=0 //x2=16.28 //y2=0
r1267 (  197 200 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=16.11 //y=0 //x2=15.17 //y2=0
r1268 (  193 478 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.13 //y=0.17 //x2=14.13 //y2=0
r1269 (  193 523 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=14.13 //y=0.17 //x2=14.13 //y2=0.955
r1270 (  192 476 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=0 //x2=12.95 //y2=0
r1271 (  191 478 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.045 //y=0 //x2=14.13 //y2=0
r1272 (  191 192 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=14.045 //y=0 //x2=13.12 //y2=0
r1273 (  186 188 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r1274 (  184 186 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=10.36 //y=0 //x2=11.47 //y2=0
r1275 (  182 475 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.3 //y=0 //x2=9.215 //y2=0
r1276 (  182 184 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=9.3 //y=0 //x2=10.36 //y2=0
r1277 (  181 476 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.95 //y2=0
r1278 (  181 188 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.58 //y2=0
r1279 (  177 475 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.215 //y=0.17 //x2=9.215 //y2=0
r1280 (  177 522 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=9.215 //y=0.17 //x2=9.215 //y2=0.965
r1281 (  176 473 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=0 //x2=8.14 //y2=0
r1282 (  175 475 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.13 //y=0 //x2=9.215 //y2=0
r1283 (  175 176 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=9.13 //y=0 //x2=8.31 //y2=0
r1284 (  170 172 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r1285 (  168 170 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=5.55 //y=0 //x2=6.66 //y2=0
r1286 (  166 472 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.49 //y=0 //x2=4.405 //y2=0
r1287 (  166 168 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=4.49 //y=0 //x2=5.55 //y2=0
r1288 (  165 473 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=8.14 //y2=0
r1289 (  165 172 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=7.77 //y2=0
r1290 (  161 472 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.405 //y=0.17 //x2=4.405 //y2=0
r1291 (  161 521 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=4.405 //y=0.17 //x2=4.405 //y2=0.965
r1292 (  160 470 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=0 //x2=3.33 //y2=0
r1293 (  159 472 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.32 //y=0 //x2=4.405 //y2=0
r1294 (  159 160 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=4.32 //y=0 //x2=3.5 //y2=0
r1295 (  154 156 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r1296 (  152 469 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.18 //y2=0
r1297 (  152 154 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.85 //y2=0
r1298 (  151 470 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=3.33 //y2=0
r1299 (  151 156 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r1300 (  147 469 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r1301 (  147 520 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.955
r1302 (  143 469 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=1.18 //y2=0
r1303 (  143 146 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=0.74 //y2=0
r1304 (  139 466 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.51 //y=0 //x2=82.51 //y2=0
r1305 (  137 464 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=81.4 //y=0 //x2=81.4 //y2=0
r1306 (  137 139 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=81.4 //y=0 //x2=82.51 //y2=0
r1307 (  135 456 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=80.29 //y=0 //x2=80.29 //y2=0
r1308 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=80.29 //y=0 //x2=81.4 //y2=0
r1309 (  133 450 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.81 //y=0 //x2=78.81 //y2=0
r1310 (  133 135 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=78.81 //y=0 //x2=80.29 //y2=0
r1311 (  131 517 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=77.7 //y=0 //x2=77.7 //y2=0
r1312 (  131 133 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=77.7 //y=0 //x2=78.81 //y2=0
r1313 (  129 438 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.22 //y=0 //x2=76.22 //y2=0
r1314 (  129 131 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.22 //y=0 //x2=77.7 //y2=0
r1315 (  127 436 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.11 //y=0 //x2=75.11 //y2=0
r1316 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=0 //x2=76.22 //y2=0
r1317 (  125 428 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74 //y=0 //x2=74 //y2=0
r1318 (  125 127 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74 //y=0 //x2=75.11 //y2=0
r1319 (  123 422 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.52 //y=0 //x2=72.52 //y2=0
r1320 (  123 125 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=72.52 //y=0 //x2=74 //y2=0
r1321 (  121 420 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=0 //x2=71.41 //y2=0
r1322 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=0 //x2=72.52 //y2=0
r1323 (  119 418 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=70.3 //y=0 //x2=70.3 //y2=0
r1324 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=70.3 //y=0 //x2=71.41 //y2=0
r1325 (  117 410 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.19 //y=0 //x2=69.19 //y2=0
r1326 (  117 119 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.19 //y=0 //x2=70.3 //y2=0
r1327 (  115 404 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=67.71 //y=0 //x2=67.71 //y2=0
r1328 (  115 117 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=67.71 //y=0 //x2=69.19 //y2=0
r1329 (  113 402 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.6 //y=0 //x2=66.6 //y2=0
r1330 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=66.6 //y=0 //x2=67.71 //y2=0
r1331 (  111 394 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.49 //y=0 //x2=65.49 //y2=0
r1332 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.49 //y=0 //x2=66.6 //y2=0
r1333 (  109 388 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=64.01 //y=0 //x2=64.01 //y2=0
r1334 (  109 111 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=64.01 //y=0 //x2=65.49 //y2=0
r1335 (  107 508 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=62.9 //y=0 //x2=62.9 //y2=0
r1336 (  107 109 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=62.9 //y=0 //x2=64.01 //y2=0
r1337 (  105 376 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.42 //y=0 //x2=61.42 //y2=0
r1338 (  105 107 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.42 //y=0 //x2=62.9 //y2=0
r1339 (  103 374 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=60.31 //y=0 //x2=60.31 //y2=0
r1340 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=60.31 //y=0 //x2=61.42 //y2=0
r1341 (  101 372 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.2 //y=0 //x2=59.2 //y2=0
r1342 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.2 //y=0 //x2=60.31 //y2=0
r1343 (  99 505 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.09 //y=0 //x2=58.09 //y2=0
r1344 (  99 101 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.09 //y=0 //x2=59.2 //y2=0
r1345 (  97 360 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.61 //y=0 //x2=56.61 //y2=0
r1346 (  97 99 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.61 //y=0 //x2=58.09 //y2=0
r1347 (  95 358 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.5 //y=0 //x2=55.5 //y2=0
r1348 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.5 //y=0 //x2=56.61 //y2=0
r1349 (  93 356 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.39 //y=0 //x2=54.39 //y2=0
r1350 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.39 //y=0 //x2=55.5 //y2=0
r1351 (  91 502 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.28 //y=0 //x2=53.28 //y2=0
r1352 (  91 93 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=53.28 //y=0 //x2=54.39 //y2=0
r1353 (  89 344 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.8 //y=0 //x2=51.8 //y2=0
r1354 (  89 91 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=51.8 //y=0 //x2=53.28 //y2=0
r1355 (  87 342 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=50.69 //y=0 //x2=50.69 //y2=0
r1356 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=50.69 //y=0 //x2=51.8 //y2=0
r1357 (  85 334 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.58 //y=0 //x2=49.58 //y2=0
r1358 (  85 87 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.58 //y=0 //x2=50.69 //y2=0
r1359 (  83 328 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.1 //y=0 //x2=48.1 //y2=0
r1360 (  83 85 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=48.1 //y=0 //x2=49.58 //y2=0
r1361 (  81 326 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.99 //y=0 //x2=46.99 //y2=0
r1362 (  81 83 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.99 //y=0 //x2=48.1 //y2=0
r1363 (  79 324 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.88 //y=0 //x2=45.88 //y2=0
r1364 (  79 81 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.88 //y=0 //x2=46.99 //y2=0
r1365 (  77 316 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.77 //y=0 //x2=44.77 //y2=0
r1366 (  77 79 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.77 //y=0 //x2=45.88 //y2=0
r1367 (  75 310 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=43.29 //y=0 //x2=43.29 //y2=0
r1368 (  75 77 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=43.29 //y=0 //x2=44.77 //y2=0
r1369 (  73 308 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.18 //y=0 //x2=42.18 //y2=0
r1370 (  73 75 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=42.18 //y=0 //x2=43.29 //y2=0
r1371 (  70 300 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.07 //y=0 //x2=41.07 //y2=0
r1372 (  68 294 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.59 //y=0 //x2=39.59 //y2=0
r1373 (  68 70 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=39.59 //y=0 //x2=41.07 //y2=0
r1374 (  66 493 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=38.48 //y=0 //x2=38.48 //y2=0
r1375 (  66 68 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=38.48 //y=0 //x2=39.59 //y2=0
r1376 (  64 282 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37 //y=0 //x2=37 //y2=0
r1377 (  64 66 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=37 //y=0 //x2=38.48 //y2=0
r1378 (  62 280 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.89 //y=0 //x2=35.89 //y2=0
r1379 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.89 //y=0 //x2=37 //y2=0
r1380 (  60 278 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.78 //y=0 //x2=34.78 //y2=0
r1381 (  60 62 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.78 //y=0 //x2=35.89 //y2=0
r1382 (  58 490 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=33.67 //y=0 //x2=33.67 //y2=0
r1383 (  58 60 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=33.67 //y=0 //x2=34.78 //y2=0
r1384 (  56 266 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.19 //y=0 //x2=32.19 //y2=0
r1385 (  56 58 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.19 //y=0 //x2=33.67 //y2=0
r1386 (  54 264 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.08 //y=0 //x2=31.08 //y2=0
r1387 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.08 //y=0 //x2=32.19 //y2=0
r1388 (  52 262 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.97 //y=0 //x2=29.97 //y2=0
r1389 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=29.97 //y=0 //x2=31.08 //y2=0
r1390 (  50 487 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.86 //y=0 //x2=28.86 //y2=0
r1391 (  50 52 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=28.86 //y=0 //x2=29.97 //y2=0
r1392 (  48 250 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.38 //y=0 //x2=27.38 //y2=0
r1393 (  48 50 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=27.38 //y=0 //x2=28.86 //y2=0
r1394 (  46 248 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.27 //y=0 //x2=26.27 //y2=0
r1395 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.27 //y=0 //x2=27.38 //y2=0
r1396 (  44 240 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.16 //y=0 //x2=25.16 //y2=0
r1397 (  44 46 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.16 //y=0 //x2=26.27 //y2=0
r1398 (  42 234 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=0 //x2=23.68 //y2=0
r1399 (  42 44 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=0 //x2=25.16 //y2=0
r1400 (  40 232 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=0 //x2=22.57 //y2=0
r1401 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=0 //x2=23.68 //y2=0
r1402 (  38 230 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.46 //y=0 //x2=21.46 //y2=0
r1403 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.46 //y=0 //x2=22.57 //y2=0
r1404 (  36 222 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=0 //x2=20.35 //y2=0
r1405 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=0 //x2=21.46 //y2=0
r1406 (  34 216 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=0 //x2=18.87 //y2=0
r1407 (  34 36 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=0 //x2=20.35 //y2=0
r1408 (  32 214 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=0 //x2=17.76 //y2=0
r1409 (  32 34 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=0 //x2=18.87 //y2=0
r1410 (  30 206 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=0 //x2=16.65 //y2=0
r1411 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=0 //x2=17.76 //y2=0
r1412 (  28 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r1413 (  28 30 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.65 //y2=0
r1414 (  26 478 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=0 //x2=14.06 //y2=0
r1415 (  26 28 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=0 //x2=15.17 //y2=0
r1416 (  24 188 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r1417 (  24 26 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=0 //x2=14.06 //y2=0
r1418 (  22 186 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r1419 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=0 //x2=12.58 //y2=0
r1420 (  20 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r1421 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r1422 (  18 475 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=0 //x2=9.25 //y2=0
r1423 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=0 //x2=10.36 //y2=0
r1424 (  16 172 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r1425 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=9.25 //y2=0
r1426 (  14 170 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r1427 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r1428 (  12 168 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r1429 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r1430 (  10 472 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r1431 (  10 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.55 //y2=0
r1432 (  8 156 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r1433 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r1434 (  6 154 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r1435 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r1436 (  3 146 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r1437 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r1438 (  1 73 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=41.625 //y=0 //x2=42.18 //y2=0
r1439 (  1 70 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=41.625 //y=0 //x2=41.07 //y2=0
ends PM_TMRDFFSNQNX1\%GND

subckt PM_TMRDFFSNQNX1\%VDD ( 1 139 151 159 169 175 183 191 201 211 217 225 \
 233 243 253 259 267 277 287 291 301 311 319 323 333 343 351 361 367 375 383 \
 393 399 407 415 425 435 441 449 457 467 477 483 491 501 511 515 525 535 543 \
 547 557 567 575 585 591 599 607 617 623 631 639 649 659 665 673 681 691 701 \
 707 715 725 735 739 749 759 767 771 781 791 799 809 815 823 831 841 847 862 \
 866 869 875 881 885 890 895 900 906 912 916 921 926 931 937 943 947 952 957 \
 962 963 964 965 966 967 968 969 970 971 972 973 974 975 976 977 978 979 980 \
 981 982 983 984 985 986 987 988 989 990 991 992 993 994 995 996 997 998 999 \
 1000 1001 1002 1003 1004 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 \
 1015 1016 1017 1018 1019 1020 1021 1022 1023 1024 1025 1026 1027 1028 1029 )
c1064 ( 1029 0 ) capacitor c=0.0476806f //x=75.665 //y=5.025
c1065 ( 1028 0 ) capacitor c=0.0241714f //x=74.785 //y=5.025
c1066 ( 1027 0 ) capacitor c=0.0467094f //x=73.915 //y=5.025
c1067 ( 1026 0 ) capacitor c=0.0452179f //x=72.035 //y=5.02
c1068 ( 1025 0 ) capacitor c=0.024152f //x=71.155 //y=5.02
c1069 ( 1024 0 ) capacitor c=0.024152f //x=70.275 //y=5.02
c1070 ( 1023 0 ) capacitor c=0.0531852f //x=69.405 //y=5.02
c1071 ( 1022 0 ) capacitor c=0.0381674f //x=67.525 //y=5.02
c1072 ( 1021 0 ) capacitor c=0.0241306f //x=66.645 //y=5.02
c1073 ( 1020 0 ) capacitor c=0.0493657f //x=65.775 //y=5.02
c1074 ( 1019 0 ) capacitor c=0.0381505f //x=64.195 //y=5.02
c1075 ( 1018 0 ) capacitor c=0.0240074f //x=63.315 //y=5.02
c1076 ( 1017 0 ) capacitor c=0.049209f //x=62.445 //y=5.02
c1077 ( 1016 0 ) capacitor c=0.0452179f //x=60.565 //y=5.02
c1078 ( 1015 0 ) capacitor c=0.024152f //x=59.685 //y=5.02
c1079 ( 1014 0 ) capacitor c=0.024152f //x=58.805 //y=5.02
c1080 ( 1013 0 ) capacitor c=0.053132f //x=57.935 //y=5.02
c1081 ( 1012 0 ) capacitor c=0.0452179f //x=55.755 //y=5.02
c1082 ( 1011 0 ) capacitor c=0.024152f //x=54.875 //y=5.02
c1083 ( 1010 0 ) capacitor c=0.024152f //x=53.995 //y=5.02
c1084 ( 1009 0 ) capacitor c=0.0531894f //x=53.125 //y=5.02
c1085 ( 1008 0 ) capacitor c=0.0380679f //x=51.245 //y=5.02
c1086 ( 1007 0 ) capacitor c=0.024008f //x=50.365 //y=5.02
c1087 ( 1006 0 ) capacitor c=0.049209f //x=49.495 //y=5.02
c1088 ( 1005 0 ) capacitor c=0.0452179f //x=47.615 //y=5.02
c1089 ( 1004 0 ) capacitor c=0.024152f //x=46.735 //y=5.02
c1090 ( 1003 0 ) capacitor c=0.024152f //x=45.855 //y=5.02
c1091 ( 1002 0 ) capacitor c=0.0531894f //x=44.985 //y=5.02
c1092 ( 1001 0 ) capacitor c=0.0380679f //x=43.105 //y=5.02
c1093 ( 1000 0 ) capacitor c=0.024008f //x=42.225 //y=5.02
c1094 ( 999 0 ) capacitor c=0.0490303f //x=41.355 //y=5.02
c1095 ( 998 0 ) capacitor c=0.0380679f //x=39.775 //y=5.02
c1096 ( 997 0 ) capacitor c=0.0240074f //x=38.895 //y=5.02
c1097 ( 996 0 ) capacitor c=0.049209f //x=38.025 //y=5.02
c1098 ( 995 0 ) capacitor c=0.0452179f //x=36.145 //y=5.02
c1099 ( 994 0 ) capacitor c=0.024152f //x=35.265 //y=5.02
c1100 ( 993 0 ) capacitor c=0.024152f //x=34.385 //y=5.02
c1101 ( 992 0 ) capacitor c=0.053132f //x=33.515 //y=5.02
c1102 ( 991 0 ) capacitor c=0.0452179f //x=31.335 //y=5.02
c1103 ( 990 0 ) capacitor c=0.024152f //x=30.455 //y=5.02
c1104 ( 989 0 ) capacitor c=0.024152f //x=29.575 //y=5.02
c1105 ( 988 0 ) capacitor c=0.0531894f //x=28.705 //y=5.02
c1106 ( 987 0 ) capacitor c=0.0380679f //x=26.825 //y=5.02
c1107 ( 986 0 ) capacitor c=0.024008f //x=25.945 //y=5.02
c1108 ( 985 0 ) capacitor c=0.049209f //x=25.075 //y=5.02
c1109 ( 984 0 ) capacitor c=0.0452179f //x=23.195 //y=5.02
c1110 ( 983 0 ) capacitor c=0.024152f //x=22.315 //y=5.02
c1111 ( 982 0 ) capacitor c=0.024152f //x=21.435 //y=5.02
c1112 ( 981 0 ) capacitor c=0.0531894f //x=20.565 //y=5.02
c1113 ( 980 0 ) capacitor c=0.0380679f //x=18.685 //y=5.02
c1114 ( 979 0 ) capacitor c=0.024008f //x=17.805 //y=5.02
c1115 ( 978 0 ) capacitor c=0.0490303f //x=16.935 //y=5.02
c1116 ( 977 0 ) capacitor c=0.0380679f //x=15.355 //y=5.02
c1117 ( 976 0 ) capacitor c=0.0240074f //x=14.475 //y=5.02
c1118 ( 975 0 ) capacitor c=0.049209f //x=13.605 //y=5.02
c1119 ( 974 0 ) capacitor c=0.0452179f //x=11.725 //y=5.02
c1120 ( 973 0 ) capacitor c=0.024152f //x=10.845 //y=5.02
c1121 ( 972 0 ) capacitor c=0.024152f //x=9.965 //y=5.02
c1122 ( 971 0 ) capacitor c=0.053132f //x=9.095 //y=5.02
c1123 ( 970 0 ) capacitor c=0.0452179f //x=6.915 //y=5.02
c1124 ( 969 0 ) capacitor c=0.024152f //x=6.035 //y=5.02
c1125 ( 968 0 ) capacitor c=0.02424f //x=5.155 //y=5.02
c1126 ( 967 0 ) capacitor c=0.0532367f //x=4.285 //y=5.02
c1127 ( 966 0 ) capacitor c=0.0381505f //x=2.405 //y=5.02
c1128 ( 965 0 ) capacitor c=0.0241853f //x=1.525 //y=5.02
c1129 ( 964 0 ) capacitor c=0.053196f //x=0.655 //y=5.02
c1130 ( 963 0 ) capacitor c=0.113329f //x=79.92 //y=7.4
c1131 ( 962 0 ) capacitor c=0.121062f //x=76.59 //y=7.4
c1132 ( 961 0 ) capacitor c=0.00591168f //x=75.81 //y=7.4
c1133 ( 960 0 ) capacitor c=0.00591168f //x=74.93 //y=7.4
c1134 ( 959 0 ) capacitor c=0.00591168f //x=74 //y=7.4
c1135 ( 957 0 ) capacitor c=0.136602f //x=73.26 //y=7.4
c1136 ( 956 0 ) capacitor c=0.00591168f //x=72.18 //y=7.4
c1137 ( 955 0 ) capacitor c=0.00591168f //x=71.3 //y=7.4
c1138 ( 954 0 ) capacitor c=0.00591168f //x=70.42 //y=7.4
c1139 ( 953 0 ) capacitor c=0.00591168f //x=69.54 //y=7.4
c1140 ( 952 0 ) capacitor c=0.13471f //x=68.45 //y=7.4
c1141 ( 951 0 ) capacitor c=0.00591168f //x=67.71 //y=7.4
c1142 ( 949 0 ) capacitor c=0.00591168f //x=66.79 //y=7.4
c1143 ( 948 0 ) capacitor c=0.00591168f //x=65.91 //y=7.4
c1144 ( 947 0 ) capacitor c=0.115932f //x=65.12 //y=7.4
c1145 ( 946 0 ) capacitor c=0.00591168f //x=64.34 //y=7.4
c1146 ( 945 0 ) capacitor c=0.00591168f //x=63.46 //y=7.4
c1147 ( 944 0 ) capacitor c=0.00591168f //x=62.58 //y=7.4
c1148 ( 943 0 ) capacitor c=0.13452f //x=61.79 //y=7.4
c1149 ( 942 0 ) capacitor c=0.00591168f //x=60.71 //y=7.4
c1150 ( 941 0 ) capacitor c=0.00591168f //x=59.83 //y=7.4
c1151 ( 940 0 ) capacitor c=0.00591168f //x=58.95 //y=7.4
c1152 ( 939 0 ) capacitor c=0.00591168f //x=58.09 //y=7.4
c1153 ( 937 0 ) capacitor c=0.155082f //x=56.98 //y=7.4
c1154 ( 936 0 ) capacitor c=0.00591168f //x=55.9 //y=7.4
c1155 ( 935 0 ) capacitor c=0.00591168f //x=55.02 //y=7.4
c1156 ( 934 0 ) capacitor c=0.00591168f //x=54.14 //y=7.4
c1157 ( 933 0 ) capacitor c=0.00591168f //x=53.28 //y=7.4
c1158 ( 931 0 ) capacitor c=0.135216f //x=52.17 //y=7.4
c1159 ( 930 0 ) capacitor c=0.00591168f //x=51.39 //y=7.4
c1160 ( 929 0 ) capacitor c=0.00591168f //x=50.51 //y=7.4
c1161 ( 928 0 ) capacitor c=0.00591168f //x=49.58 //y=7.4
c1162 ( 926 0 ) capacitor c=0.138747f //x=48.84 //y=7.4
c1163 ( 925 0 ) capacitor c=0.00591168f //x=47.76 //y=7.4
c1164 ( 924 0 ) capacitor c=0.00591168f //x=46.88 //y=7.4
c1165 ( 923 0 ) capacitor c=0.00591168f //x=46 //y=7.4
c1166 ( 922 0 ) capacitor c=0.00591168f //x=45.12 //y=7.4
c1167 ( 921 0 ) capacitor c=0.135109f //x=44.03 //y=7.4
c1168 ( 920 0 ) capacitor c=0.00591168f //x=43.29 //y=7.4
c1169 ( 918 0 ) capacitor c=0.00591168f //x=42.37 //y=7.4
c1170 ( 917 0 ) capacitor c=0.00591168f //x=41.49 //y=7.4
c1171 ( 916 0 ) capacitor c=0.11432f //x=40.7 //y=7.4
c1172 ( 915 0 ) capacitor c=0.00591168f //x=39.92 //y=7.4
c1173 ( 914 0 ) capacitor c=0.00591168f //x=39.04 //y=7.4
c1174 ( 913 0 ) capacitor c=0.00591168f //x=38.16 //y=7.4
c1175 ( 912 0 ) capacitor c=0.13452f //x=37.37 //y=7.4
c1176 ( 911 0 ) capacitor c=0.00591168f //x=36.29 //y=7.4
c1177 ( 910 0 ) capacitor c=0.00591168f //x=35.41 //y=7.4
c1178 ( 909 0 ) capacitor c=0.00591168f //x=34.53 //y=7.4
c1179 ( 908 0 ) capacitor c=0.00591168f //x=33.67 //y=7.4
c1180 ( 906 0 ) capacitor c=0.155082f //x=32.56 //y=7.4
c1181 ( 905 0 ) capacitor c=0.00591168f //x=31.48 //y=7.4
c1182 ( 904 0 ) capacitor c=0.00591168f //x=30.6 //y=7.4
c1183 ( 903 0 ) capacitor c=0.00591168f //x=29.72 //y=7.4
c1184 ( 902 0 ) capacitor c=0.00591168f //x=28.86 //y=7.4
c1185 ( 900 0 ) capacitor c=0.135216f //x=27.75 //y=7.4
c1186 ( 899 0 ) capacitor c=0.00591168f //x=26.97 //y=7.4
c1187 ( 898 0 ) capacitor c=0.00591168f //x=26.09 //y=7.4
c1188 ( 897 0 ) capacitor c=0.00591168f //x=25.16 //y=7.4
c1189 ( 895 0 ) capacitor c=0.138734f //x=24.42 //y=7.4
c1190 ( 894 0 ) capacitor c=0.00591168f //x=23.34 //y=7.4
c1191 ( 893 0 ) capacitor c=0.00591168f //x=22.46 //y=7.4
c1192 ( 892 0 ) capacitor c=0.00591168f //x=21.58 //y=7.4
c1193 ( 891 0 ) capacitor c=0.00591168f //x=20.7 //y=7.4
c1194 ( 890 0 ) capacitor c=0.135109f //x=19.61 //y=7.4
c1195 ( 889 0 ) capacitor c=0.00591168f //x=18.87 //y=7.4
c1196 ( 887 0 ) capacitor c=0.00591168f //x=17.95 //y=7.4
c1197 ( 886 0 ) capacitor c=0.00591168f //x=17.07 //y=7.4
c1198 ( 885 0 ) capacitor c=0.11432f //x=16.28 //y=7.4
c1199 ( 884 0 ) capacitor c=0.00591168f //x=15.5 //y=7.4
c1200 ( 883 0 ) capacitor c=0.00591168f //x=14.62 //y=7.4
c1201 ( 882 0 ) capacitor c=0.00591168f //x=13.74 //y=7.4
c1202 ( 881 0 ) capacitor c=0.13452f //x=12.95 //y=7.4
c1203 ( 880 0 ) capacitor c=0.00591168f //x=11.87 //y=7.4
c1204 ( 879 0 ) capacitor c=0.00591168f //x=10.99 //y=7.4
c1205 ( 878 0 ) capacitor c=0.00591168f //x=10.11 //y=7.4
c1206 ( 877 0 ) capacitor c=0.00591168f //x=9.25 //y=7.4
c1207 ( 875 0 ) capacitor c=0.155082f //x=8.14 //y=7.4
c1208 ( 874 0 ) capacitor c=0.00591168f //x=7.06 //y=7.4
c1209 ( 873 0 ) capacitor c=0.00591168f //x=6.18 //y=7.4
c1210 ( 872 0 ) capacitor c=0.00591168f //x=5.3 //y=7.4
c1211 ( 871 0 ) capacitor c=0.00591168f //x=4.44 //y=7.4
c1212 ( 869 0 ) capacitor c=0.137297f //x=3.33 //y=7.4
c1213 ( 868 0 ) capacitor c=0.00591168f //x=2.55 //y=7.4
c1214 ( 867 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c1215 ( 866 0 ) capacitor c=0.248311f //x=0.74 //y=7.4
c1216 ( 862 0 ) capacitor c=0.334471f //x=82.51 //y=7.4
c1217 ( 847 0 ) capacitor c=0.120978f //x=79.75 //y=7.4
c1218 ( 841 0 ) capacitor c=0.0236224f //x=76.42 //y=7.4
c1219 ( 831 0 ) capacitor c=0.028539f //x=75.725 //y=7.4
c1220 ( 823 0 ) capacitor c=0.0285075f //x=74.845 //y=7.4
c1221 ( 815 0 ) capacitor c=0.0240981f //x=73.965 //y=7.4
c1222 ( 809 0 ) capacitor c=0.0394667f //x=73.09 //y=7.4
c1223 ( 799 0 ) capacitor c=0.0288488f //x=72.095 //y=7.4
c1224 ( 791 0 ) capacitor c=0.0287514f //x=71.215 //y=7.4
c1225 ( 781 0 ) capacitor c=0.0284966f //x=70.335 //y=7.4
c1226 ( 771 0 ) capacitor c=0.0383672f //x=69.455 //y=7.4
c1227 ( 767 0 ) capacitor c=0.0237088f //x=68.28 //y=7.4
c1228 ( 759 0 ) capacitor c=0.0288637f //x=67.585 //y=7.4
c1229 ( 749 0 ) capacitor c=0.0291038f //x=66.705 //y=7.4
c1230 ( 739 0 ) capacitor c=0.0240981f //x=65.825 //y=7.4
c1231 ( 735 0 ) capacitor c=0.0236224f //x=64.95 //y=7.4
c1232 ( 725 0 ) capacitor c=0.0288598f //x=64.255 //y=7.4
c1233 ( 715 0 ) capacitor c=0.0288369f //x=63.375 //y=7.4
c1234 ( 707 0 ) capacitor c=0.0240981f //x=62.495 //y=7.4
c1235 ( 701 0 ) capacitor c=0.0394667f //x=61.62 //y=7.4
c1236 ( 691 0 ) capacitor c=0.0288488f //x=60.625 //y=7.4
c1237 ( 681 0 ) capacitor c=0.0287514f //x=59.745 //y=7.4
c1238 ( 673 0 ) capacitor c=0.0284966f //x=58.865 //y=7.4
c1239 ( 665 0 ) capacitor c=0.0383672f //x=57.985 //y=7.4
c1240 ( 659 0 ) capacitor c=0.0394667f //x=56.81 //y=7.4
c1241 ( 649 0 ) capacitor c=0.0288488f //x=55.815 //y=7.4
c1242 ( 639 0 ) capacitor c=0.0287505f //x=54.935 //y=7.4
c1243 ( 631 0 ) capacitor c=0.0284966f //x=54.055 //y=7.4
c1244 ( 623 0 ) capacitor c=0.0383672f //x=53.175 //y=7.4
c1245 ( 617 0 ) capacitor c=0.0236224f //x=52 //y=7.4
c1246 ( 607 0 ) capacitor c=0.0288359f //x=51.305 //y=7.4
c1247 ( 599 0 ) capacitor c=0.0288369f //x=50.425 //y=7.4
c1248 ( 591 0 ) capacitor c=0.0240981f //x=49.545 //y=7.4
c1249 ( 585 0 ) capacitor c=0.0394667f //x=48.67 //y=7.4
c1250 ( 575 0 ) capacitor c=0.0288488f //x=47.675 //y=7.4
c1251 ( 567 0 ) capacitor c=0.0287514f //x=46.795 //y=7.4
c1252 ( 557 0 ) capacitor c=0.0284966f //x=45.915 //y=7.4
c1253 ( 547 0 ) capacitor c=0.0383672f //x=45.035 //y=7.4
c1254 ( 543 0 ) capacitor c=0.0236224f //x=43.86 //y=7.4
c1255 ( 535 0 ) capacitor c=0.0288359f //x=43.165 //y=7.4
c1256 ( 525 0 ) capacitor c=0.0288369f //x=42.285 //y=7.4
c1257 ( 515 0 ) capacitor c=0.0240981f //x=41.405 //y=7.4
c1258 ( 511 0 ) capacitor c=0.0236224f //x=40.53 //y=7.4
c1259 ( 501 0 ) capacitor c=0.0288357f //x=39.835 //y=7.4
c1260 ( 491 0 ) capacitor c=0.0288369f //x=38.955 //y=7.4
c1261 ( 483 0 ) capacitor c=0.0240981f //x=38.075 //y=7.4
c1262 ( 477 0 ) capacitor c=0.0394667f //x=37.2 //y=7.4
c1263 ( 467 0 ) capacitor c=0.0288488f //x=36.205 //y=7.4
c1264 ( 457 0 ) capacitor c=0.0287514f //x=35.325 //y=7.4
c1265 ( 449 0 ) capacitor c=0.0284966f //x=34.445 //y=7.4
c1266 ( 441 0 ) capacitor c=0.0383672f //x=33.565 //y=7.4
c1267 ( 435 0 ) capacitor c=0.0394667f //x=32.39 //y=7.4
c1268 ( 425 0 ) capacitor c=0.0288488f //x=31.395 //y=7.4
c1269 ( 415 0 ) capacitor c=0.0287505f //x=30.515 //y=7.4
c1270 ( 407 0 ) capacitor c=0.0284966f //x=29.635 //y=7.4
c1271 ( 399 0 ) capacitor c=0.0383672f //x=28.755 //y=7.4
c1272 ( 393 0 ) capacitor c=0.0236224f //x=27.58 //y=7.4
c1273 ( 383 0 ) capacitor c=0.0288359f //x=26.885 //y=7.4
c1274 ( 375 0 ) capacitor c=0.0288369f //x=26.005 //y=7.4
c1275 ( 367 0 ) capacitor c=0.0240981f //x=25.125 //y=7.4
c1276 ( 361 0 ) capacitor c=0.0394667f //x=24.25 //y=7.4
c1277 ( 351 0 ) capacitor c=0.0288488f //x=23.255 //y=7.4
c1278 ( 343 0 ) capacitor c=0.0287514f //x=22.375 //y=7.4
c1279 ( 333 0 ) capacitor c=0.0284966f //x=21.495 //y=7.4
c1280 ( 323 0 ) capacitor c=0.0383672f //x=20.615 //y=7.4
c1281 ( 319 0 ) capacitor c=0.0236224f //x=19.44 //y=7.4
c1282 ( 311 0 ) capacitor c=0.0288359f //x=18.745 //y=7.4
c1283 ( 301 0 ) capacitor c=0.0288369f //x=17.865 //y=7.4
c1284 ( 291 0 ) capacitor c=0.0240981f //x=16.985 //y=7.4
c1285 ( 287 0 ) capacitor c=0.0236224f //x=16.11 //y=7.4
c1286 ( 277 0 ) capacitor c=0.0288357f //x=15.415 //y=7.4
c1287 ( 267 0 ) capacitor c=0.0288369f //x=14.535 //y=7.4
c1288 ( 259 0 ) capacitor c=0.0240981f //x=13.655 //y=7.4
c1289 ( 253 0 ) capacitor c=0.0394667f //x=12.78 //y=7.4
c1290 ( 243 0 ) capacitor c=0.0288488f //x=11.785 //y=7.4
c1291 ( 233 0 ) capacitor c=0.0287514f //x=10.905 //y=7.4
c1292 ( 225 0 ) capacitor c=0.0284966f //x=10.025 //y=7.4
c1293 ( 217 0 ) capacitor c=0.0383672f //x=9.145 //y=7.4
c1294 ( 211 0 ) capacitor c=0.0394667f //x=7.97 //y=7.4
c1295 ( 201 0 ) capacitor c=0.0288488f //x=6.975 //y=7.4
c1296 ( 191 0 ) capacitor c=0.0287505f //x=6.095 //y=7.4
c1297 ( 183 0 ) capacitor c=0.028511f //x=5.215 //y=7.4
c1298 ( 175 0 ) capacitor c=0.0383672f //x=4.335 //y=7.4
c1299 ( 169 0 ) capacitor c=0.0236224f //x=3.16 //y=7.4
c1300 ( 159 0 ) capacitor c=0.0288637f //x=2.465 //y=7.4
c1301 ( 151 0 ) capacitor c=0.0286367f //x=1.585 //y=7.4
c1302 ( 139 0 ) capacitor c=2.74745f //x=82.51 //y=7.4
r1303 (  860 862 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=81.4 //y=7.4 //x2=82.51 //y2=7.4
r1304 (  858 860 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=80.29 //y=7.4 //x2=81.4 //y2=7.4
r1305 (  856 963 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=80.09 //y=7.4 //x2=79.92 //y2=7.4
r1306 (  856 858 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=80.09 //y=7.4 //x2=80.29 //y2=7.4
r1307 (  850 852 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=77.7 //y=7.4 //x2=78.81 //y2=7.4
r1308 (  848 962 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.76 //y=7.4 //x2=76.59 //y2=7.4
r1309 (  848 850 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=76.76 //y=7.4 //x2=77.7 //y2=7.4
r1310 (  847 963 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=79.75 //y=7.4 //x2=79.92 //y2=7.4
r1311 (  847 852 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=79.75 //y=7.4 //x2=78.81 //y2=7.4
r1312 (  842 961 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.895 //y=7.4 //x2=75.81 //y2=7.4
r1313 (  842 844 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=75.895 //y=7.4 //x2=76.22 //y2=7.4
r1314 (  841 962 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.42 //y=7.4 //x2=76.59 //y2=7.4
r1315 (  841 844 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=76.42 //y=7.4 //x2=76.22 //y2=7.4
r1316 (  835 961 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=75.81 //y=7.23 //x2=75.81 //y2=7.4
r1317 (  835 1029 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=75.81 //y=7.23 //x2=75.81 //y2=6.4
r1318 (  832 960 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.015 //y=7.4 //x2=74.93 //y2=7.4
r1319 (  832 834 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=75.015 //y=7.4 //x2=75.11 //y2=7.4
r1320 (  831 961 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.725 //y=7.4 //x2=75.81 //y2=7.4
r1321 (  831 834 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=75.725 //y=7.4 //x2=75.11 //y2=7.4
r1322 (  825 960 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.93 //y=7.23 //x2=74.93 //y2=7.4
r1323 (  825 1028 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=74.93 //y=7.23 //x2=74.93 //y2=6.74
r1324 (  824 959 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.135 //y=7.4 //x2=74.05 //y2=7.4
r1325 (  823 960 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.845 //y=7.4 //x2=74.93 //y2=7.4
r1326 (  823 824 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=74.845 //y=7.4 //x2=74.135 //y2=7.4
r1327 (  817 959 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.05 //y=7.23 //x2=74.05 //y2=7.4
r1328 (  817 1027 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=74.05 //y=7.23 //x2=74.05 //y2=6.4
r1329 (  816 957 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.43 //y=7.4 //x2=73.26 //y2=7.4
r1330 (  815 959 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.965 //y=7.4 //x2=74.05 //y2=7.4
r1331 (  815 816 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=73.965 //y=7.4 //x2=73.43 //y2=7.4
r1332 (  810 956 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.265 //y=7.4 //x2=72.18 //y2=7.4
r1333 (  810 812 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=72.265 //y=7.4 //x2=72.52 //y2=7.4
r1334 (  809 957 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.09 //y=7.4 //x2=73.26 //y2=7.4
r1335 (  809 812 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=73.09 //y=7.4 //x2=72.52 //y2=7.4
r1336 (  803 956 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=72.18 //y=7.23 //x2=72.18 //y2=7.4
r1337 (  803 1026 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=72.18 //y=7.23 //x2=72.18 //y2=6.745
r1338 (  800 955 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.385 //y=7.4 //x2=71.3 //y2=7.4
r1339 (  800 802 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=71.385 //y=7.4 //x2=71.41 //y2=7.4
r1340 (  799 956 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.095 //y=7.4 //x2=72.18 //y2=7.4
r1341 (  799 802 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=72.095 //y=7.4 //x2=71.41 //y2=7.4
r1342 (  793 955 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.3 //y=7.23 //x2=71.3 //y2=7.4
r1343 (  793 1025 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=71.3 //y=7.23 //x2=71.3 //y2=6.745
r1344 (  792 954 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.505 //y=7.4 //x2=70.42 //y2=7.4
r1345 (  791 955 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.215 //y=7.4 //x2=71.3 //y2=7.4
r1346 (  791 792 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=71.215 //y=7.4 //x2=70.505 //y2=7.4
r1347 (  785 954 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=70.42 //y=7.23 //x2=70.42 //y2=7.4
r1348 (  785 1024 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=70.42 //y=7.23 //x2=70.42 //y2=6.745
r1349 (  782 953 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.625 //y=7.4 //x2=69.54 //y2=7.4
r1350 (  782 784 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=69.625 //y=7.4 //x2=70.3 //y2=7.4
r1351 (  781 954 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.335 //y=7.4 //x2=70.42 //y2=7.4
r1352 (  781 784 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=70.335 //y=7.4 //x2=70.3 //y2=7.4
r1353 (  775 953 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.54 //y=7.23 //x2=69.54 //y2=7.4
r1354 (  775 1023 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=69.54 //y=7.23 //x2=69.54 //y2=6.405
r1355 (  772 952 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.62 //y=7.4 //x2=68.45 //y2=7.4
r1356 (  772 774 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=68.62 //y=7.4 //x2=69.19 //y2=7.4
r1357 (  771 953 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.455 //y=7.4 //x2=69.54 //y2=7.4
r1358 (  771 774 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=69.455 //y=7.4 //x2=69.19 //y2=7.4
r1359 (  768 951 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.755 //y=7.4 //x2=67.67 //y2=7.4
r1360 (  767 952 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.28 //y=7.4 //x2=68.45 //y2=7.4
r1361 (  767 768 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=68.28 //y=7.4 //x2=67.755 //y2=7.4
r1362 (  761 951 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.67 //y=7.23 //x2=67.67 //y2=7.4
r1363 (  761 1022 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=67.67 //y=7.23 //x2=67.67 //y2=6.745
r1364 (  760 949 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.875 //y=7.4 //x2=66.79 //y2=7.4
r1365 (  759 951 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.585 //y=7.4 //x2=67.67 //y2=7.4
r1366 (  759 760 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=67.585 //y=7.4 //x2=66.875 //y2=7.4
r1367 (  753 949 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=66.79 //y=7.23 //x2=66.79 //y2=7.4
r1368 (  753 1021 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=66.79 //y=7.23 //x2=66.79 //y2=6.745
r1369 (  750 948 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.995 //y=7.4 //x2=65.91 //y2=7.4
r1370 (  750 752 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=65.995 //y=7.4 //x2=66.6 //y2=7.4
r1371 (  749 949 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.705 //y=7.4 //x2=66.79 //y2=7.4
r1372 (  749 752 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=66.705 //y=7.4 //x2=66.6 //y2=7.4
r1373 (  743 948 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.91 //y=7.23 //x2=65.91 //y2=7.4
r1374 (  743 1020 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=65.91 //y=7.23 //x2=65.91 //y2=6.405
r1375 (  740 947 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.29 //y=7.4 //x2=65.12 //y2=7.4
r1376 (  740 742 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=65.29 //y=7.4 //x2=65.49 //y2=7.4
r1377 (  739 948 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.825 //y=7.4 //x2=65.91 //y2=7.4
r1378 (  739 742 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=65.825 //y=7.4 //x2=65.49 //y2=7.4
r1379 (  736 946 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.425 //y=7.4 //x2=64.34 //y2=7.4
r1380 (  735 947 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.95 //y=7.4 //x2=65.12 //y2=7.4
r1381 (  735 736 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=64.95 //y=7.4 //x2=64.425 //y2=7.4
r1382 (  729 946 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.34 //y=7.23 //x2=64.34 //y2=7.4
r1383 (  729 1019 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=64.34 //y=7.23 //x2=64.34 //y2=6.745
r1384 (  726 945 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.545 //y=7.4 //x2=63.46 //y2=7.4
r1385 (  726 728 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=63.545 //y=7.4 //x2=64.01 //y2=7.4
r1386 (  725 946 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.255 //y=7.4 //x2=64.34 //y2=7.4
r1387 (  725 728 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=64.255 //y=7.4 //x2=64.01 //y2=7.4
r1388 (  719 945 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=63.46 //y=7.23 //x2=63.46 //y2=7.4
r1389 (  719 1018 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=63.46 //y=7.23 //x2=63.46 //y2=6.745
r1390 (  716 944 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.665 //y=7.4 //x2=62.58 //y2=7.4
r1391 (  716 718 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=62.665 //y=7.4 //x2=62.9 //y2=7.4
r1392 (  715 945 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.375 //y=7.4 //x2=63.46 //y2=7.4
r1393 (  715 718 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=63.375 //y=7.4 //x2=62.9 //y2=7.4
r1394 (  709 944 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.58 //y=7.23 //x2=62.58 //y2=7.4
r1395 (  709 1017 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=62.58 //y=7.23 //x2=62.58 //y2=6.405
r1396 (  708 943 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.96 //y=7.4 //x2=61.79 //y2=7.4
r1397 (  707 944 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.495 //y=7.4 //x2=62.58 //y2=7.4
r1398 (  707 708 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=62.495 //y=7.4 //x2=61.96 //y2=7.4
r1399 (  702 942 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.795 //y=7.4 //x2=60.71 //y2=7.4
r1400 (  702 704 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=60.795 //y=7.4 //x2=61.42 //y2=7.4
r1401 (  701 943 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.62 //y=7.4 //x2=61.79 //y2=7.4
r1402 (  701 704 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=61.62 //y=7.4 //x2=61.42 //y2=7.4
r1403 (  695 942 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=60.71 //y=7.23 //x2=60.71 //y2=7.4
r1404 (  695 1016 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.71 //y=7.23 //x2=60.71 //y2=6.745
r1405 (  692 941 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.915 //y=7.4 //x2=59.83 //y2=7.4
r1406 (  692 694 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=59.915 //y=7.4 //x2=60.31 //y2=7.4
r1407 (  691 942 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.625 //y=7.4 //x2=60.71 //y2=7.4
r1408 (  691 694 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=60.625 //y=7.4 //x2=60.31 //y2=7.4
r1409 (  685 941 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=59.83 //y=7.23 //x2=59.83 //y2=7.4
r1410 (  685 1015 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.83 //y=7.23 //x2=59.83 //y2=6.745
r1411 (  682 940 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.035 //y=7.4 //x2=58.95 //y2=7.4
r1412 (  682 684 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=59.035 //y=7.4 //x2=59.2 //y2=7.4
r1413 (  681 941 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.745 //y=7.4 //x2=59.83 //y2=7.4
r1414 (  681 684 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=59.745 //y=7.4 //x2=59.2 //y2=7.4
r1415 (  675 940 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.95 //y=7.23 //x2=58.95 //y2=7.4
r1416 (  675 1014 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=58.95 //y=7.23 //x2=58.95 //y2=6.745
r1417 (  674 939 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.155 //y=7.4 //x2=58.07 //y2=7.4
r1418 (  673 940 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.865 //y=7.4 //x2=58.95 //y2=7.4
r1419 (  673 674 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=58.865 //y=7.4 //x2=58.155 //y2=7.4
r1420 (  667 939 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.07 //y=7.23 //x2=58.07 //y2=7.4
r1421 (  667 1013 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=58.07 //y=7.23 //x2=58.07 //y2=6.405
r1422 (  666 937 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.15 //y=7.4 //x2=56.98 //y2=7.4
r1423 (  665 939 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=57.985 //y=7.4 //x2=58.07 //y2=7.4
r1424 (  665 666 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=57.985 //y=7.4 //x2=57.15 //y2=7.4
r1425 (  660 936 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.985 //y=7.4 //x2=55.9 //y2=7.4
r1426 (  660 662 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=55.985 //y=7.4 //x2=56.61 //y2=7.4
r1427 (  659 937 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.81 //y=7.4 //x2=56.98 //y2=7.4
r1428 (  659 662 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=56.81 //y=7.4 //x2=56.61 //y2=7.4
r1429 (  653 936 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=55.9 //y=7.23 //x2=55.9 //y2=7.4
r1430 (  653 1012 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.9 //y=7.23 //x2=55.9 //y2=6.745
r1431 (  650 935 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.105 //y=7.4 //x2=55.02 //y2=7.4
r1432 (  650 652 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=55.105 //y=7.4 //x2=55.5 //y2=7.4
r1433 (  649 936 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.815 //y=7.4 //x2=55.9 //y2=7.4
r1434 (  649 652 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=55.815 //y=7.4 //x2=55.5 //y2=7.4
r1435 (  643 935 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=55.02 //y=7.23 //x2=55.02 //y2=7.4
r1436 (  643 1011 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.02 //y=7.23 //x2=55.02 //y2=6.745
r1437 (  640 934 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.225 //y=7.4 //x2=54.14 //y2=7.4
r1438 (  640 642 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=54.225 //y=7.4 //x2=54.39 //y2=7.4
r1439 (  639 935 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.935 //y=7.4 //x2=55.02 //y2=7.4
r1440 (  639 642 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=54.935 //y=7.4 //x2=54.39 //y2=7.4
r1441 (  633 934 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=54.14 //y=7.23 //x2=54.14 //y2=7.4
r1442 (  633 1010 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.14 //y=7.23 //x2=54.14 //y2=6.745
r1443 (  632 933 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.345 //y=7.4 //x2=53.26 //y2=7.4
r1444 (  631 934 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.055 //y=7.4 //x2=54.14 //y2=7.4
r1445 (  631 632 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=54.055 //y=7.4 //x2=53.345 //y2=7.4
r1446 (  625 933 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.26 //y=7.23 //x2=53.26 //y2=7.4
r1447 (  625 1009 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=53.26 //y=7.23 //x2=53.26 //y2=6.405
r1448 (  624 931 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.34 //y=7.4 //x2=52.17 //y2=7.4
r1449 (  623 933 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.175 //y=7.4 //x2=53.26 //y2=7.4
r1450 (  623 624 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=53.175 //y=7.4 //x2=52.34 //y2=7.4
r1451 (  618 930 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.475 //y=7.4 //x2=51.39 //y2=7.4
r1452 (  618 620 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=51.475 //y=7.4 //x2=51.8 //y2=7.4
r1453 (  617 931 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52 //y=7.4 //x2=52.17 //y2=7.4
r1454 (  617 620 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=52 //y=7.4 //x2=51.8 //y2=7.4
r1455 (  611 930 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.39 //y=7.23 //x2=51.39 //y2=7.4
r1456 (  611 1008 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=51.39 //y=7.23 //x2=51.39 //y2=6.745
r1457 (  608 929 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.595 //y=7.4 //x2=50.51 //y2=7.4
r1458 (  608 610 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=50.595 //y=7.4 //x2=50.69 //y2=7.4
r1459 (  607 930 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.305 //y=7.4 //x2=51.39 //y2=7.4
r1460 (  607 610 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=51.305 //y=7.4 //x2=50.69 //y2=7.4
r1461 (  601 929 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.51 //y=7.23 //x2=50.51 //y2=7.4
r1462 (  601 1007 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.51 //y=7.23 //x2=50.51 //y2=6.745
r1463 (  600 928 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.715 //y=7.4 //x2=49.63 //y2=7.4
r1464 (  599 929 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.425 //y=7.4 //x2=50.51 //y2=7.4
r1465 (  599 600 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.425 //y=7.4 //x2=49.715 //y2=7.4
r1466 (  593 928 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.63 //y=7.23 //x2=49.63 //y2=7.4
r1467 (  593 1006 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=49.63 //y=7.23 //x2=49.63 //y2=6.405
r1468 (  592 926 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.01 //y=7.4 //x2=48.84 //y2=7.4
r1469 (  591 928 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.545 //y=7.4 //x2=49.63 //y2=7.4
r1470 (  591 592 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=49.545 //y=7.4 //x2=49.01 //y2=7.4
r1471 (  586 925 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.845 //y=7.4 //x2=47.76 //y2=7.4
r1472 (  586 588 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=47.845 //y=7.4 //x2=48.1 //y2=7.4
r1473 (  585 926 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.67 //y=7.4 //x2=48.84 //y2=7.4
r1474 (  585 588 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.67 //y=7.4 //x2=48.1 //y2=7.4
r1475 (  579 925 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.76 //y=7.23 //x2=47.76 //y2=7.4
r1476 (  579 1005 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=47.76 //y=7.23 //x2=47.76 //y2=6.745
r1477 (  576 924 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.965 //y=7.4 //x2=46.88 //y2=7.4
r1478 (  576 578 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=46.965 //y=7.4 //x2=46.99 //y2=7.4
r1479 (  575 925 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.675 //y=7.4 //x2=47.76 //y2=7.4
r1480 (  575 578 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=47.675 //y=7.4 //x2=46.99 //y2=7.4
r1481 (  569 924 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=46.88 //y=7.23 //x2=46.88 //y2=7.4
r1482 (  569 1004 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.88 //y=7.23 //x2=46.88 //y2=6.745
r1483 (  568 923 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.085 //y=7.4 //x2=46 //y2=7.4
r1484 (  567 924 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.795 //y=7.4 //x2=46.88 //y2=7.4
r1485 (  567 568 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.795 //y=7.4 //x2=46.085 //y2=7.4
r1486 (  561 923 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=46 //y=7.23 //x2=46 //y2=7.4
r1487 (  561 1003 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46 //y=7.23 //x2=46 //y2=6.745
r1488 (  558 922 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.205 //y=7.4 //x2=45.12 //y2=7.4
r1489 (  558 560 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=45.205 //y=7.4 //x2=45.88 //y2=7.4
r1490 (  557 923 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.915 //y=7.4 //x2=46 //y2=7.4
r1491 (  557 560 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=45.915 //y=7.4 //x2=45.88 //y2=7.4
r1492 (  551 922 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=45.12 //y=7.23 //x2=45.12 //y2=7.4
r1493 (  551 1002 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=45.12 //y=7.23 //x2=45.12 //y2=6.405
r1494 (  548 921 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.2 //y=7.4 //x2=44.03 //y2=7.4
r1495 (  548 550 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=44.2 //y=7.4 //x2=44.77 //y2=7.4
r1496 (  547 922 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.035 //y=7.4 //x2=45.12 //y2=7.4
r1497 (  547 550 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=45.035 //y=7.4 //x2=44.77 //y2=7.4
r1498 (  544 920 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=43.335 //y=7.4 //x2=43.25 //y2=7.4
r1499 (  543 921 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.86 //y=7.4 //x2=44.03 //y2=7.4
r1500 (  543 544 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=43.86 //y=7.4 //x2=43.335 //y2=7.4
r1501 (  537 920 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.25 //y=7.23 //x2=43.25 //y2=7.4
r1502 (  537 1001 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=43.25 //y=7.23 //x2=43.25 //y2=6.745
r1503 (  536 918 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.455 //y=7.4 //x2=42.37 //y2=7.4
r1504 (  535 920 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=43.165 //y=7.4 //x2=43.25 //y2=7.4
r1505 (  535 536 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=43.165 //y=7.4 //x2=42.455 //y2=7.4
r1506 (  529 918 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=42.37 //y=7.23 //x2=42.37 //y2=7.4
r1507 (  529 1000 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=42.37 //y=7.23 //x2=42.37 //y2=6.745
r1508 (  526 917 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.575 //y=7.4 //x2=41.49 //y2=7.4
r1509 (  526 528 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=41.575 //y=7.4 //x2=42.18 //y2=7.4
r1510 (  525 918 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.285 //y=7.4 //x2=42.37 //y2=7.4
r1511 (  525 528 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=42.285 //y=7.4 //x2=42.18 //y2=7.4
r1512 (  519 917 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=41.49 //y=7.23 //x2=41.49 //y2=7.4
r1513 (  519 999 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=41.49 //y=7.23 //x2=41.49 //y2=6.405
r1514 (  516 916 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.87 //y=7.4 //x2=40.7 //y2=7.4
r1515 (  516 518 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=40.87 //y=7.4 //x2=41.07 //y2=7.4
r1516 (  515 917 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.405 //y=7.4 //x2=41.49 //y2=7.4
r1517 (  515 518 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=41.405 //y=7.4 //x2=41.07 //y2=7.4
r1518 (  512 915 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.005 //y=7.4 //x2=39.92 //y2=7.4
r1519 (  511 916 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.53 //y=7.4 //x2=40.7 //y2=7.4
r1520 (  511 512 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=40.53 //y=7.4 //x2=40.005 //y2=7.4
r1521 (  505 915 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.92 //y=7.23 //x2=39.92 //y2=7.4
r1522 (  505 998 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=39.92 //y=7.23 //x2=39.92 //y2=6.745
r1523 (  502 914 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.125 //y=7.4 //x2=39.04 //y2=7.4
r1524 (  502 504 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=39.125 //y=7.4 //x2=39.59 //y2=7.4
r1525 (  501 915 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.835 //y=7.4 //x2=39.92 //y2=7.4
r1526 (  501 504 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=39.835 //y=7.4 //x2=39.59 //y2=7.4
r1527 (  495 914 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.04 //y=7.23 //x2=39.04 //y2=7.4
r1528 (  495 997 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=39.04 //y=7.23 //x2=39.04 //y2=6.745
r1529 (  492 913 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.245 //y=7.4 //x2=38.16 //y2=7.4
r1530 (  492 494 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=38.245 //y=7.4 //x2=38.48 //y2=7.4
r1531 (  491 914 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.955 //y=7.4 //x2=39.04 //y2=7.4
r1532 (  491 494 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=38.955 //y=7.4 //x2=38.48 //y2=7.4
r1533 (  485 913 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.16 //y=7.23 //x2=38.16 //y2=7.4
r1534 (  485 996 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=38.16 //y=7.23 //x2=38.16 //y2=6.405
r1535 (  484 912 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.54 //y=7.4 //x2=37.37 //y2=7.4
r1536 (  483 913 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.075 //y=7.4 //x2=38.16 //y2=7.4
r1537 (  483 484 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=38.075 //y=7.4 //x2=37.54 //y2=7.4
r1538 (  478 911 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.375 //y=7.4 //x2=36.29 //y2=7.4
r1539 (  478 480 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=36.375 //y=7.4 //x2=37 //y2=7.4
r1540 (  477 912 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.2 //y=7.4 //x2=37.37 //y2=7.4
r1541 (  477 480 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=37.2 //y=7.4 //x2=37 //y2=7.4
r1542 (  471 911 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.29 //y=7.23 //x2=36.29 //y2=7.4
r1543 (  471 995 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=36.29 //y=7.23 //x2=36.29 //y2=6.745
r1544 (  468 910 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.495 //y=7.4 //x2=35.41 //y2=7.4
r1545 (  468 470 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=35.495 //y=7.4 //x2=35.89 //y2=7.4
r1546 (  467 911 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.205 //y=7.4 //x2=36.29 //y2=7.4
r1547 (  467 470 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=36.205 //y=7.4 //x2=35.89 //y2=7.4
r1548 (  461 910 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.41 //y=7.23 //x2=35.41 //y2=7.4
r1549 (  461 994 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.41 //y=7.23 //x2=35.41 //y2=6.745
r1550 (  458 909 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.615 //y=7.4 //x2=34.53 //y2=7.4
r1551 (  458 460 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=34.615 //y=7.4 //x2=34.78 //y2=7.4
r1552 (  457 910 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.325 //y=7.4 //x2=35.41 //y2=7.4
r1553 (  457 460 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=35.325 //y=7.4 //x2=34.78 //y2=7.4
r1554 (  451 909 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.53 //y=7.23 //x2=34.53 //y2=7.4
r1555 (  451 993 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=34.53 //y=7.23 //x2=34.53 //y2=6.745
r1556 (  450 908 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.735 //y=7.4 //x2=33.65 //y2=7.4
r1557 (  449 909 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.445 //y=7.4 //x2=34.53 //y2=7.4
r1558 (  449 450 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=34.445 //y=7.4 //x2=33.735 //y2=7.4
r1559 (  443 908 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.65 //y=7.23 //x2=33.65 //y2=7.4
r1560 (  443 992 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=33.65 //y=7.23 //x2=33.65 //y2=6.405
r1561 (  442 906 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.73 //y=7.4 //x2=32.56 //y2=7.4
r1562 (  441 908 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.565 //y=7.4 //x2=33.65 //y2=7.4
r1563 (  441 442 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=33.565 //y=7.4 //x2=32.73 //y2=7.4
r1564 (  436 905 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.565 //y=7.4 //x2=31.48 //y2=7.4
r1565 (  436 438 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=31.565 //y=7.4 //x2=32.19 //y2=7.4
r1566 (  435 906 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.39 //y=7.4 //x2=32.56 //y2=7.4
r1567 (  435 438 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=32.39 //y=7.4 //x2=32.19 //y2=7.4
r1568 (  429 905 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.48 //y=7.23 //x2=31.48 //y2=7.4
r1569 (  429 991 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.48 //y=7.23 //x2=31.48 //y2=6.745
r1570 (  426 904 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.685 //y=7.4 //x2=30.6 //y2=7.4
r1571 (  426 428 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=30.685 //y=7.4 //x2=31.08 //y2=7.4
r1572 (  425 905 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.395 //y=7.4 //x2=31.48 //y2=7.4
r1573 (  425 428 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=31.395 //y=7.4 //x2=31.08 //y2=7.4
r1574 (  419 904 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.6 //y=7.23 //x2=30.6 //y2=7.4
r1575 (  419 990 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=30.6 //y=7.23 //x2=30.6 //y2=6.745
r1576 (  416 903 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.805 //y=7.4 //x2=29.72 //y2=7.4
r1577 (  416 418 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=29.805 //y=7.4 //x2=29.97 //y2=7.4
r1578 (  415 904 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.515 //y=7.4 //x2=30.6 //y2=7.4
r1579 (  415 418 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=30.515 //y=7.4 //x2=29.97 //y2=7.4
r1580 (  409 903 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.72 //y=7.23 //x2=29.72 //y2=7.4
r1581 (  409 989 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=29.72 //y=7.23 //x2=29.72 //y2=6.745
r1582 (  408 902 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.925 //y=7.4 //x2=28.84 //y2=7.4
r1583 (  407 903 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.635 //y=7.4 //x2=29.72 //y2=7.4
r1584 (  407 408 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=29.635 //y=7.4 //x2=28.925 //y2=7.4
r1585 (  401 902 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.84 //y=7.23 //x2=28.84 //y2=7.4
r1586 (  401 988 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=28.84 //y=7.23 //x2=28.84 //y2=6.405
r1587 (  400 900 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.92 //y=7.4 //x2=27.75 //y2=7.4
r1588 (  399 902 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.755 //y=7.4 //x2=28.84 //y2=7.4
r1589 (  399 400 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=28.755 //y=7.4 //x2=27.92 //y2=7.4
r1590 (  394 899 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.055 //y=7.4 //x2=26.97 //y2=7.4
r1591 (  394 396 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=27.055 //y=7.4 //x2=27.38 //y2=7.4
r1592 (  393 900 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.58 //y=7.4 //x2=27.75 //y2=7.4
r1593 (  393 396 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=27.58 //y=7.4 //x2=27.38 //y2=7.4
r1594 (  387 899 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.97 //y=7.23 //x2=26.97 //y2=7.4
r1595 (  387 987 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.97 //y=7.23 //x2=26.97 //y2=6.745
r1596 (  384 898 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.175 //y=7.4 //x2=26.09 //y2=7.4
r1597 (  384 386 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=26.175 //y=7.4 //x2=26.27 //y2=7.4
r1598 (  383 899 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.885 //y=7.4 //x2=26.97 //y2=7.4
r1599 (  383 386 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=26.885 //y=7.4 //x2=26.27 //y2=7.4
r1600 (  377 898 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.09 //y=7.23 //x2=26.09 //y2=7.4
r1601 (  377 986 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.09 //y=7.23 //x2=26.09 //y2=6.745
r1602 (  376 897 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.295 //y=7.4 //x2=25.21 //y2=7.4
r1603 (  375 898 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.005 //y=7.4 //x2=26.09 //y2=7.4
r1604 (  375 376 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.005 //y=7.4 //x2=25.295 //y2=7.4
r1605 (  369 897 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.21 //y=7.23 //x2=25.21 //y2=7.4
r1606 (  369 985 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=25.21 //y=7.23 //x2=25.21 //y2=6.405
r1607 (  368 895 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.59 //y=7.4 //x2=24.42 //y2=7.4
r1608 (  367 897 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.125 //y=7.4 //x2=25.21 //y2=7.4
r1609 (  367 368 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=25.125 //y=7.4 //x2=24.59 //y2=7.4
r1610 (  362 894 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.425 //y=7.4 //x2=23.34 //y2=7.4
r1611 (  362 364 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=23.425 //y=7.4 //x2=23.68 //y2=7.4
r1612 (  361 895 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.25 //y=7.4 //x2=24.42 //y2=7.4
r1613 (  361 364 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.25 //y=7.4 //x2=23.68 //y2=7.4
r1614 (  355 894 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.34 //y=7.23 //x2=23.34 //y2=7.4
r1615 (  355 984 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=23.34 //y=7.23 //x2=23.34 //y2=6.745
r1616 (  352 893 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.545 //y=7.4 //x2=22.46 //y2=7.4
r1617 (  352 354 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=22.545 //y=7.4 //x2=22.57 //y2=7.4
r1618 (  351 894 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.255 //y=7.4 //x2=23.34 //y2=7.4
r1619 (  351 354 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=23.255 //y=7.4 //x2=22.57 //y2=7.4
r1620 (  345 893 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.46 //y=7.23 //x2=22.46 //y2=7.4
r1621 (  345 983 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.46 //y=7.23 //x2=22.46 //y2=6.745
r1622 (  344 892 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.665 //y=7.4 //x2=21.58 //y2=7.4
r1623 (  343 893 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.375 //y=7.4 //x2=22.46 //y2=7.4
r1624 (  343 344 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.375 //y=7.4 //x2=21.665 //y2=7.4
r1625 (  337 892 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.58 //y=7.23 //x2=21.58 //y2=7.4
r1626 (  337 982 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.58 //y=7.23 //x2=21.58 //y2=6.745
r1627 (  334 891 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.785 //y=7.4 //x2=20.7 //y2=7.4
r1628 (  334 336 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=20.785 //y=7.4 //x2=21.46 //y2=7.4
r1629 (  333 892 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.495 //y=7.4 //x2=21.58 //y2=7.4
r1630 (  333 336 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=21.495 //y=7.4 //x2=21.46 //y2=7.4
r1631 (  327 891 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.7 //y=7.23 //x2=20.7 //y2=7.4
r1632 (  327 981 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=20.7 //y=7.23 //x2=20.7 //y2=6.405
r1633 (  324 890 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.78 //y=7.4 //x2=19.61 //y2=7.4
r1634 (  324 326 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.78 //y=7.4 //x2=20.35 //y2=7.4
r1635 (  323 891 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.615 //y=7.4 //x2=20.7 //y2=7.4
r1636 (  323 326 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.615 //y=7.4 //x2=20.35 //y2=7.4
r1637 (  320 889 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.915 //y=7.4 //x2=18.83 //y2=7.4
r1638 (  319 890 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.44 //y=7.4 //x2=19.61 //y2=7.4
r1639 (  319 320 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=19.44 //y=7.4 //x2=18.915 //y2=7.4
r1640 (  313 889 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.83 //y=7.23 //x2=18.83 //y2=7.4
r1641 (  313 980 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=18.83 //y=7.23 //x2=18.83 //y2=6.745
r1642 (  312 887 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.035 //y=7.4 //x2=17.95 //y2=7.4
r1643 (  311 889 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.745 //y=7.4 //x2=18.83 //y2=7.4
r1644 (  311 312 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=18.745 //y=7.4 //x2=18.035 //y2=7.4
r1645 (  305 887 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.95 //y=7.23 //x2=17.95 //y2=7.4
r1646 (  305 979 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.95 //y=7.23 //x2=17.95 //y2=6.745
r1647 (  302 886 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.155 //y=7.4 //x2=17.07 //y2=7.4
r1648 (  302 304 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=17.155 //y=7.4 //x2=17.76 //y2=7.4
r1649 (  301 887 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.865 //y=7.4 //x2=17.95 //y2=7.4
r1650 (  301 304 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=17.865 //y=7.4 //x2=17.76 //y2=7.4
r1651 (  295 886 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.07 //y=7.23 //x2=17.07 //y2=7.4
r1652 (  295 978 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=17.07 //y=7.23 //x2=17.07 //y2=6.405
r1653 (  292 885 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.45 //y=7.4 //x2=16.28 //y2=7.4
r1654 (  292 294 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=16.45 //y=7.4 //x2=16.65 //y2=7.4
r1655 (  291 886 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.985 //y=7.4 //x2=17.07 //y2=7.4
r1656 (  291 294 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=16.985 //y=7.4 //x2=16.65 //y2=7.4
r1657 (  288 884 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.585 //y=7.4 //x2=15.5 //y2=7.4
r1658 (  287 885 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.11 //y=7.4 //x2=16.28 //y2=7.4
r1659 (  287 288 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=16.11 //y=7.4 //x2=15.585 //y2=7.4
r1660 (  281 884 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.5 //y=7.23 //x2=15.5 //y2=7.4
r1661 (  281 977 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.5 //y=7.23 //x2=15.5 //y2=6.745
r1662 (  278 883 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.705 //y=7.4 //x2=14.62 //y2=7.4
r1663 (  278 280 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=14.705 //y=7.4 //x2=15.17 //y2=7.4
r1664 (  277 884 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.415 //y=7.4 //x2=15.5 //y2=7.4
r1665 (  277 280 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=15.415 //y=7.4 //x2=15.17 //y2=7.4
r1666 (  271 883 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.62 //y=7.23 //x2=14.62 //y2=7.4
r1667 (  271 976 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.62 //y=7.23 //x2=14.62 //y2=6.745
r1668 (  268 882 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.825 //y=7.4 //x2=13.74 //y2=7.4
r1669 (  268 270 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=13.825 //y=7.4 //x2=14.06 //y2=7.4
r1670 (  267 883 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.535 //y=7.4 //x2=14.62 //y2=7.4
r1671 (  267 270 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=14.535 //y=7.4 //x2=14.06 //y2=7.4
r1672 (  261 882 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.74 //y=7.23 //x2=13.74 //y2=7.4
r1673 (  261 975 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=13.74 //y=7.23 //x2=13.74 //y2=6.405
r1674 (  260 881 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=7.4 //x2=12.95 //y2=7.4
r1675 (  259 882 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.655 //y=7.4 //x2=13.74 //y2=7.4
r1676 (  259 260 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=13.655 //y=7.4 //x2=13.12 //y2=7.4
r1677 (  254 880 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.955 //y=7.4 //x2=11.87 //y2=7.4
r1678 (  254 256 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=11.955 //y=7.4 //x2=12.58 //y2=7.4
r1679 (  253 881 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.95 //y2=7.4
r1680 (  253 256 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.58 //y2=7.4
r1681 (  247 880 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.87 //y=7.23 //x2=11.87 //y2=7.4
r1682 (  247 974 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.87 //y=7.23 //x2=11.87 //y2=6.745
r1683 (  244 879 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.075 //y=7.4 //x2=10.99 //y2=7.4
r1684 (  244 246 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=11.075 //y=7.4 //x2=11.47 //y2=7.4
r1685 (  243 880 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.785 //y=7.4 //x2=11.87 //y2=7.4
r1686 (  243 246 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=11.785 //y=7.4 //x2=11.47 //y2=7.4
r1687 (  237 879 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.99 //y=7.23 //x2=10.99 //y2=7.4
r1688 (  237 973 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.99 //y=7.23 //x2=10.99 //y2=6.745
r1689 (  234 878 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.195 //y=7.4 //x2=10.11 //y2=7.4
r1690 (  234 236 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=10.195 //y=7.4 //x2=10.36 //y2=7.4
r1691 (  233 879 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.905 //y=7.4 //x2=10.99 //y2=7.4
r1692 (  233 236 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=10.905 //y=7.4 //x2=10.36 //y2=7.4
r1693 (  227 878 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.11 //y=7.23 //x2=10.11 //y2=7.4
r1694 (  227 972 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.11 //y=7.23 //x2=10.11 //y2=6.745
r1695 (  226 877 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.315 //y=7.4 //x2=9.23 //y2=7.4
r1696 (  225 878 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.025 //y=7.4 //x2=10.11 //y2=7.4
r1697 (  225 226 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.025 //y=7.4 //x2=9.315 //y2=7.4
r1698 (  219 877 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.23 //y=7.23 //x2=9.23 //y2=7.4
r1699 (  219 971 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=9.23 //y=7.23 //x2=9.23 //y2=6.405
r1700 (  218 875 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=7.4 //x2=8.14 //y2=7.4
r1701 (  217 877 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.145 //y=7.4 //x2=9.23 //y2=7.4
r1702 (  217 218 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=9.145 //y=7.4 //x2=8.31 //y2=7.4
r1703 (  212 874 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.145 //y=7.4 //x2=7.06 //y2=7.4
r1704 (  212 214 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=7.145 //y=7.4 //x2=7.77 //y2=7.4
r1705 (  211 875 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=8.14 //y2=7.4
r1706 (  211 214 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=7.77 //y2=7.4
r1707 (  205 874 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.06 //y=7.23 //x2=7.06 //y2=7.4
r1708 (  205 970 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.06 //y=7.23 //x2=7.06 //y2=6.745
r1709 (  202 873 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.265 //y=7.4 //x2=6.18 //y2=7.4
r1710 (  202 204 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=6.265 //y=7.4 //x2=6.66 //y2=7.4
r1711 (  201 874 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.975 //y=7.4 //x2=7.06 //y2=7.4
r1712 (  201 204 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=6.975 //y=7.4 //x2=6.66 //y2=7.4
r1713 (  195 873 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.18 //y=7.23 //x2=6.18 //y2=7.4
r1714 (  195 969 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.18 //y=7.23 //x2=6.18 //y2=6.745
r1715 (  192 872 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.385 //y=7.4 //x2=5.3 //y2=7.4
r1716 (  192 194 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=5.385 //y=7.4 //x2=5.55 //y2=7.4
r1717 (  191 873 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.095 //y=7.4 //x2=6.18 //y2=7.4
r1718 (  191 194 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=6.095 //y=7.4 //x2=5.55 //y2=7.4
r1719 (  185 872 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.3 //y=7.23 //x2=5.3 //y2=7.4
r1720 (  185 968 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=5.3 //y=7.23 //x2=5.3 //y2=6.745
r1721 (  184 871 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.505 //y=7.4 //x2=4.42 //y2=7.4
r1722 (  183 872 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.215 //y=7.4 //x2=5.3 //y2=7.4
r1723 (  183 184 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.215 //y=7.4 //x2=4.505 //y2=7.4
r1724 (  177 871 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.42 //y=7.23 //x2=4.42 //y2=7.4
r1725 (  177 967 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.42 //y=7.23 //x2=4.42 //y2=6.405
r1726 (  176 869 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r1727 (  175 871 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.335 //y=7.4 //x2=4.42 //y2=7.4
r1728 (  175 176 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=4.335 //y=7.4 //x2=3.5 //y2=7.4
r1729 (  170 868 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.55 //y2=7.4
r1730 (  170 172 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.96 //y2=7.4
r1731 (  169 869 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r1732 (  169 172 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r1733 (  163 868 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r1734 (  163 966 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.745
r1735 (  160 867 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r1736 (  160 162 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r1737 (  159 868 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r1738 (  159 162 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r1739 (  153 867 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r1740 (  153 965 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.745
r1741 (  152 866 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r1742 (  151 867 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r1743 (  151 152 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r1744 (  145 866 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r1745 (  145 964 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.405
r1746 (  139 862 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.51 //y=7.4 //x2=82.51 //y2=7.4
r1747 (  137 860 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=81.4 //y=7.4 //x2=81.4 //y2=7.4
r1748 (  137 139 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=81.4 //y=7.4 //x2=82.51 //y2=7.4
r1749 (  135 858 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=80.29 //y=7.4 //x2=80.29 //y2=7.4
r1750 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=80.29 //y=7.4 //x2=81.4 //y2=7.4
r1751 (  133 852 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.81 //y=7.4 //x2=78.81 //y2=7.4
r1752 (  133 135 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=78.81 //y=7.4 //x2=80.29 //y2=7.4
r1753 (  131 850 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=77.7 //y=7.4 //x2=77.7 //y2=7.4
r1754 (  131 133 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=77.7 //y=7.4 //x2=78.81 //y2=7.4
r1755 (  129 844 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.22 //y=7.4 //x2=76.22 //y2=7.4
r1756 (  129 131 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.22 //y=7.4 //x2=77.7 //y2=7.4
r1757 (  127 834 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.11 //y=7.4 //x2=75.11 //y2=7.4
r1758 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=7.4 //x2=76.22 //y2=7.4
r1759 (  125 959 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74 //y=7.4 //x2=74 //y2=7.4
r1760 (  125 127 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74 //y=7.4 //x2=75.11 //y2=7.4
r1761 (  123 812 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.52 //y=7.4 //x2=72.52 //y2=7.4
r1762 (  123 125 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=72.52 //y=7.4 //x2=74 //y2=7.4
r1763 (  121 802 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=7.4 //x2=71.41 //y2=7.4
r1764 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=7.4 //x2=72.52 //y2=7.4
r1765 (  119 784 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=70.3 //y=7.4 //x2=70.3 //y2=7.4
r1766 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=70.3 //y=7.4 //x2=71.41 //y2=7.4
r1767 (  117 774 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.19 //y=7.4 //x2=69.19 //y2=7.4
r1768 (  117 119 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.19 //y=7.4 //x2=70.3 //y2=7.4
r1769 (  115 951 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=67.71 //y=7.4 //x2=67.71 //y2=7.4
r1770 (  115 117 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=67.71 //y=7.4 //x2=69.19 //y2=7.4
r1771 (  113 752 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.6 //y=7.4 //x2=66.6 //y2=7.4
r1772 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=66.6 //y=7.4 //x2=67.71 //y2=7.4
r1773 (  111 742 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.49 //y=7.4 //x2=65.49 //y2=7.4
r1774 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.49 //y=7.4 //x2=66.6 //y2=7.4
r1775 (  109 728 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=64.01 //y=7.4 //x2=64.01 //y2=7.4
r1776 (  109 111 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=64.01 //y=7.4 //x2=65.49 //y2=7.4
r1777 (  107 718 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=62.9 //y=7.4 //x2=62.9 //y2=7.4
r1778 (  107 109 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=62.9 //y=7.4 //x2=64.01 //y2=7.4
r1779 (  105 704 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.42 //y=7.4 //x2=61.42 //y2=7.4
r1780 (  105 107 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.42 //y=7.4 //x2=62.9 //y2=7.4
r1781 (  103 694 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=60.31 //y=7.4 //x2=60.31 //y2=7.4
r1782 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=60.31 //y=7.4 //x2=61.42 //y2=7.4
r1783 (  101 684 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.2 //y=7.4 //x2=59.2 //y2=7.4
r1784 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.2 //y=7.4 //x2=60.31 //y2=7.4
r1785 (  99 939 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.09 //y=7.4 //x2=58.09 //y2=7.4
r1786 (  99 101 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.09 //y=7.4 //x2=59.2 //y2=7.4
r1787 (  97 662 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.61 //y=7.4 //x2=56.61 //y2=7.4
r1788 (  97 99 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.61 //y=7.4 //x2=58.09 //y2=7.4
r1789 (  95 652 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.5 //y=7.4 //x2=55.5 //y2=7.4
r1790 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.5 //y=7.4 //x2=56.61 //y2=7.4
r1791 (  93 642 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.39 //y=7.4 //x2=54.39 //y2=7.4
r1792 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.39 //y=7.4 //x2=55.5 //y2=7.4
r1793 (  91 933 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.28 //y=7.4 //x2=53.28 //y2=7.4
r1794 (  91 93 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=53.28 //y=7.4 //x2=54.39 //y2=7.4
r1795 (  89 620 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.8 //y=7.4 //x2=51.8 //y2=7.4
r1796 (  89 91 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=51.8 //y=7.4 //x2=53.28 //y2=7.4
r1797 (  87 610 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=50.69 //y=7.4 //x2=50.69 //y2=7.4
r1798 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=50.69 //y=7.4 //x2=51.8 //y2=7.4
r1799 (  85 928 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.58 //y=7.4 //x2=49.58 //y2=7.4
r1800 (  85 87 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.58 //y=7.4 //x2=50.69 //y2=7.4
r1801 (  83 588 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.1 //y=7.4 //x2=48.1 //y2=7.4
r1802 (  83 85 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=48.1 //y=7.4 //x2=49.58 //y2=7.4
r1803 (  81 578 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.99 //y=7.4 //x2=46.99 //y2=7.4
r1804 (  81 83 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.99 //y=7.4 //x2=48.1 //y2=7.4
r1805 (  79 560 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.88 //y=7.4 //x2=45.88 //y2=7.4
r1806 (  79 81 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.88 //y=7.4 //x2=46.99 //y2=7.4
r1807 (  77 550 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.77 //y=7.4 //x2=44.77 //y2=7.4
r1808 (  77 79 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.77 //y=7.4 //x2=45.88 //y2=7.4
r1809 (  75 920 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=43.29 //y=7.4 //x2=43.29 //y2=7.4
r1810 (  75 77 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=43.29 //y=7.4 //x2=44.77 //y2=7.4
r1811 (  73 528 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.18 //y=7.4 //x2=42.18 //y2=7.4
r1812 (  73 75 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=42.18 //y=7.4 //x2=43.29 //y2=7.4
r1813 (  70 518 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.07 //y=7.4 //x2=41.07 //y2=7.4
r1814 (  68 504 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.59 //y=7.4 //x2=39.59 //y2=7.4
r1815 (  68 70 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=39.59 //y=7.4 //x2=41.07 //y2=7.4
r1816 (  66 494 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=38.48 //y=7.4 //x2=38.48 //y2=7.4
r1817 (  66 68 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=38.48 //y=7.4 //x2=39.59 //y2=7.4
r1818 (  64 480 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37 //y=7.4 //x2=37 //y2=7.4
r1819 (  64 66 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=37 //y=7.4 //x2=38.48 //y2=7.4
r1820 (  62 470 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.89 //y=7.4 //x2=35.89 //y2=7.4
r1821 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.89 //y=7.4 //x2=37 //y2=7.4
r1822 (  60 460 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.78 //y=7.4 //x2=34.78 //y2=7.4
r1823 (  60 62 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.78 //y=7.4 //x2=35.89 //y2=7.4
r1824 (  58 908 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=33.67 //y=7.4 //x2=33.67 //y2=7.4
r1825 (  58 60 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=33.67 //y=7.4 //x2=34.78 //y2=7.4
r1826 (  56 438 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.19 //y=7.4 //x2=32.19 //y2=7.4
r1827 (  56 58 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.19 //y=7.4 //x2=33.67 //y2=7.4
r1828 (  54 428 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.08 //y=7.4 //x2=31.08 //y2=7.4
r1829 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.08 //y=7.4 //x2=32.19 //y2=7.4
r1830 (  52 418 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.97 //y=7.4 //x2=29.97 //y2=7.4
r1831 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=29.97 //y=7.4 //x2=31.08 //y2=7.4
r1832 (  50 902 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.86 //y=7.4 //x2=28.86 //y2=7.4
r1833 (  50 52 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=28.86 //y=7.4 //x2=29.97 //y2=7.4
r1834 (  48 396 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.38 //y=7.4 //x2=27.38 //y2=7.4
r1835 (  48 50 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=27.38 //y=7.4 //x2=28.86 //y2=7.4
r1836 (  46 386 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.27 //y=7.4 //x2=26.27 //y2=7.4
r1837 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.27 //y=7.4 //x2=27.38 //y2=7.4
r1838 (  44 897 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.16 //y=7.4 //x2=25.16 //y2=7.4
r1839 (  44 46 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.16 //y=7.4 //x2=26.27 //y2=7.4
r1840 (  42 364 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=7.4 //x2=23.68 //y2=7.4
r1841 (  42 44 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=7.4 //x2=25.16 //y2=7.4
r1842 (  40 354 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=7.4 //x2=22.57 //y2=7.4
r1843 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=7.4 //x2=23.68 //y2=7.4
r1844 (  38 336 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.46 //y=7.4 //x2=21.46 //y2=7.4
r1845 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.46 //y=7.4 //x2=22.57 //y2=7.4
r1846 (  36 326 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=7.4 //x2=20.35 //y2=7.4
r1847 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=7.4 //x2=21.46 //y2=7.4
r1848 (  34 889 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=7.4 //x2=18.87 //y2=7.4
r1849 (  34 36 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=7.4 //x2=20.35 //y2=7.4
r1850 (  32 304 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=7.4 //x2=17.76 //y2=7.4
r1851 (  32 34 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=7.4 //x2=18.87 //y2=7.4
r1852 (  30 294 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=7.4 //x2=16.65 //y2=7.4
r1853 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=7.4 //x2=17.76 //y2=7.4
r1854 (  28 280 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r1855 (  28 30 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.65 //y2=7.4
r1856 (  26 270 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=7.4 //x2=14.06 //y2=7.4
r1857 (  26 28 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=7.4 //x2=15.17 //y2=7.4
r1858 (  24 256 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r1859 (  24 26 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.4 //x2=14.06 //y2=7.4
r1860 (  22 246 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r1861 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=7.4 //x2=12.58 //y2=7.4
r1862 (  20 236 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r1863 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r1864 (  18 877 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=7.4 //x2=9.25 //y2=7.4
r1865 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=7.4 //x2=10.36 //y2=7.4
r1866 (  16 214 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r1867 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=9.25 //y2=7.4
r1868 (  14 204 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r1869 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r1870 (  12 194 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r1871 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r1872 (  10 871 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r1873 (  10 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.55 //y2=7.4
r1874 (  8 172 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r1875 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r1876 (  6 162 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r1877 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r1878 (  3 866 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r1879 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r1880 (  1 73 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=41.625 //y=7.4 //x2=42.18 //y2=7.4
r1881 (  1 70 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=41.625 //y=7.4 //x2=41.07 //y2=7.4
ends PM_TMRDFFSNQNX1\%VDD

subckt PM_TMRDFFSNQNX1\%noxref_3 ( 1 2 3 4 17 18 29 31 32 36 38 46 53 54 55 56 \
 57 58 59 60 61 62 63 64 66 72 73 74 75 79 80 81 82 83 85 91 92 93 94 114 116 \
 117 )
c244 ( 117 0 ) capacitor c=0.0220291f //x=1.965 //y=5.02
c245 ( 116 0 ) capacitor c=0.0217503f //x=1.085 //y=5.02
c246 ( 114 0 ) capacitor c=0.0084702f //x=1.96 //y=0.905
c247 ( 94 0 ) capacitor c=0.0556143f //x=9.525 //y=4.79
c248 ( 93 0 ) capacitor c=0.0293157f //x=9.815 //y=4.79
c249 ( 92 0 ) capacitor c=0.0347816f //x=9.48 //y=1.22
c250 ( 91 0 ) capacitor c=0.0187487f //x=9.48 //y=0.875
c251 ( 85 0 ) capacitor c=0.0137055f //x=9.325 //y=1.375
c252 ( 83 0 ) capacitor c=0.0149861f //x=9.325 //y=0.72
c253 ( 82 0 ) capacitor c=0.0965257f //x=8.95 //y=1.915
c254 ( 81 0 ) capacitor c=0.0229444f //x=8.95 //y=1.53
c255 ( 80 0 ) capacitor c=0.0234352f //x=8.95 //y=1.22
c256 ( 79 0 ) capacitor c=0.0198724f //x=8.95 //y=0.875
c257 ( 75 0 ) capacitor c=0.055995f //x=4.715 //y=4.79
c258 ( 74 0 ) capacitor c=0.0298189f //x=5.005 //y=4.79
c259 ( 73 0 ) capacitor c=0.0347816f //x=4.67 //y=1.22
c260 ( 72 0 ) capacitor c=0.0187487f //x=4.67 //y=0.875
c261 ( 66 0 ) capacitor c=0.0137055f //x=4.515 //y=1.375
c262 ( 64 0 ) capacitor c=0.0149861f //x=4.515 //y=0.72
c263 ( 63 0 ) capacitor c=0.0965245f //x=4.14 //y=1.915
c264 ( 62 0 ) capacitor c=0.0229444f //x=4.14 //y=1.53
c265 ( 61 0 ) capacitor c=0.0234352f //x=4.14 //y=1.22
c266 ( 60 0 ) capacitor c=0.0198724f //x=4.14 //y=0.875
c267 ( 59 0 ) capacitor c=0.110114f //x=9.89 //y=6.02
c268 ( 58 0 ) capacitor c=0.158956f //x=9.45 //y=6.02
c269 ( 57 0 ) capacitor c=0.110114f //x=5.08 //y=6.02
c270 ( 56 0 ) capacitor c=0.158956f //x=4.64 //y=6.02
c271 ( 53 0 ) capacitor c=0.0023043f //x=2.11 //y=5.2
c272 ( 46 0 ) capacitor c=0.100197f //x=9.25 //y=2.08
c273 ( 38 0 ) capacitor c=0.104868f //x=4.44 //y=2.08
c274 ( 36 0 ) capacitor c=0.110973f //x=2.59 //y=2.59
c275 ( 32 0 ) capacitor c=0.00468667f //x=2.235 //y=1.655
c276 ( 31 0 ) capacitor c=0.013082f //x=2.505 //y=1.655
c277 ( 29 0 ) capacitor c=0.0140934f //x=2.505 //y=5.2
c278 ( 18 0 ) capacitor c=0.00295092f //x=1.315 //y=5.2
c279 ( 17 0 ) capacitor c=0.0162034f //x=2.025 //y=5.2
c280 ( 4 0 ) capacitor c=0.00988709f //x=4.705 //y=2.59
c281 ( 3 0 ) capacitor c=0.110983f //x=9.135 //y=2.59
c282 ( 2 0 ) capacitor c=0.0138866f //x=2.705 //y=2.59
c283 ( 1 0 ) capacitor c=0.0386784f //x=4.295 //y=2.59
r284 (  93 95 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.815 //y=4.79 //x2=9.89 //y2=4.865
r285 (  93 94 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=9.815 //y=4.79 //x2=9.525 //y2=4.79
r286 (  92 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.48 //y=1.22 //x2=9.44 //y2=1.375
r287 (  91 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.48 //y=0.875 //x2=9.44 //y2=0.72
r288 (  91 92 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.48 //y=0.875 //x2=9.48 //y2=1.22
r289 (  88 94 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.45 //y=4.865 //x2=9.525 //y2=4.79
r290 (  88 111 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=9.45 //y=4.865 //x2=9.25 //y2=4.7
r291 (  86 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.105 //y=1.375 //x2=8.99 //y2=1.375
r292 (  85 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.325 //y=1.375 //x2=9.44 //y2=1.375
r293 (  84 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.105 //y=0.72 //x2=8.99 //y2=0.72
r294 (  83 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.325 //y=0.72 //x2=9.44 //y2=0.72
r295 (  83 84 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=9.325 //y=0.72 //x2=9.105 //y2=0.72
r296 (  82 109 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.915 //x2=9.25 //y2=2.08
r297 (  81 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.53 //x2=8.99 //y2=1.375
r298 (  81 82 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.53 //x2=8.95 //y2=1.915
r299 (  80 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.22 //x2=8.99 //y2=1.375
r300 (  79 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=0.875 //x2=8.99 //y2=0.72
r301 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.95 //y=0.875 //x2=8.95 //y2=1.22
r302 (  74 76 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.005 //y=4.79 //x2=5.08 //y2=4.865
r303 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=5.005 //y=4.79 //x2=4.715 //y2=4.79
r304 (  73 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.67 //y=1.22 //x2=4.63 //y2=1.375
r305 (  72 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.67 //y=0.875 //x2=4.63 //y2=0.72
r306 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.67 //y=0.875 //x2=4.67 //y2=1.22
r307 (  69 75 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.64 //y=4.865 //x2=4.715 //y2=4.79
r308 (  69 103 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=4.64 //y=4.865 //x2=4.44 //y2=4.7
r309 (  67 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.295 //y=1.375 //x2=4.18 //y2=1.375
r310 (  66 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.515 //y=1.375 //x2=4.63 //y2=1.375
r311 (  65 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.295 //y=0.72 //x2=4.18 //y2=0.72
r312 (  64 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.515 //y=0.72 //x2=4.63 //y2=0.72
r313 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.515 //y=0.72 //x2=4.295 //y2=0.72
r314 (  63 101 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.915 //x2=4.44 //y2=2.08
r315 (  62 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.53 //x2=4.18 //y2=1.375
r316 (  62 63 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.53 //x2=4.14 //y2=1.915
r317 (  61 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.22 //x2=4.18 //y2=1.375
r318 (  60 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=0.875 //x2=4.18 //y2=0.72
r319 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.14 //y=0.875 //x2=4.14 //y2=1.22
r320 (  59 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.89 //y=6.02 //x2=9.89 //y2=4.865
r321 (  58 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.45 //y=6.02 //x2=9.45 //y2=4.865
r322 (  57 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.08 //y=6.02 //x2=5.08 //y2=4.865
r323 (  56 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.64 //y=6.02 //x2=4.64 //y2=4.865
r324 (  55 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.375 //x2=9.325 //y2=1.375
r325 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.375 //x2=9.105 //y2=1.375
r326 (  54 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.405 //y=1.375 //x2=4.515 //y2=1.375
r327 (  54 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.405 //y=1.375 //x2=4.295 //y2=1.375
r328 (  51 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=4.7 //x2=9.25 //y2=4.7
r329 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.59 //x2=9.25 //y2=4.7
r330 (  46 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=2.08 //x2=9.25 //y2=2.08
r331 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.08 //x2=9.25 //y2=2.59
r332 (  43 103 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=4.7 //x2=4.44 //y2=4.7
r333 (  41 43 ) resistor r=144.77 //w=0.187 //l=2.115 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.585 //x2=4.44 //y2=4.7
r334 (  38 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=2.08 //x2=4.44 //y2=2.08
r335 (  38 41 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.08 //x2=4.44 //y2=2.585
r336 (  34 36 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.115 //x2=2.59 //y2=2.59
r337 (  33 36 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=2.59
r338 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r339 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r340 (  30 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.195 //y=5.2 //x2=2.11 //y2=5.2
r341 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.59 //y2=5.115
r342 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.195 //y2=5.2
r343 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.235 //y2=1.655
r344 (  25 114 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r345 (  19 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.2
r346 (  19 117 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.725
r347 (  17 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=2.11 //y2=5.2
r348 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=1.315 //y2=5.2
r349 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.315 //y2=5.2
r350 (  11 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.23 //y2=5.725
r351 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.25 //y=2.59 //x2=9.25 //y2=2.59
r352 (  8 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=2.585 //x2=4.44 //y2=2.585
r353 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=2.59 //x2=2.59 //y2=2.59
r354 (  4 8 ) resistor r=0.164988 //w=0.206 //l=0.267488 //layer=m1 \
 //thickness=0.36 //x=4.705 //y=2.59 //x2=4.44 //y2=2.585
r355 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.135 //y=2.59 //x2=9.25 //y2=2.59
r356 (  3 4 ) resistor r=4.2271 //w=0.131 //l=4.43 //layer=m1 //thickness=0.36 \
 //x=9.135 //y=2.59 //x2=4.705 //y2=2.59
r357 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=2.59 //x2=2.59 //y2=2.59
r358 (  1 8 ) resistor r=0.0921728 //w=0.206 //l=0.147479 //layer=m1 \
 //thickness=0.36 //x=4.295 //y=2.59 //x2=4.44 //y2=2.585
r359 (  1 2 ) resistor r=1.51718 //w=0.131 //l=1.59 //layer=m1 \
 //thickness=0.36 //x=4.295 //y=2.59 //x2=2.705 //y2=2.59
ends PM_TMRDFFSNQNX1\%noxref_3

subckt PM_TMRDFFSNQNX1\%noxref_4 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 61 63 66 67 77 80 82 83 84 )
c164 ( 84 0 ) capacitor c=0.023087f //x=11.285 //y=5.02
c165 ( 83 0 ) capacitor c=0.023519f //x=10.405 //y=5.02
c166 ( 82 0 ) capacitor c=0.0224735f //x=9.525 //y=5.02
c167 ( 80 0 ) capacitor c=0.00872971f //x=11.535 //y=0.915
c168 ( 77 0 ) capacitor c=0.0588816f //x=14.06 //y=4.7
c169 ( 67 0 ) capacitor c=0.0318948f //x=14.395 //y=1.21
c170 ( 66 0 ) capacitor c=0.0187384f //x=14.395 //y=0.865
c171 ( 63 0 ) capacitor c=0.0141798f //x=14.24 //y=1.365
c172 ( 61 0 ) capacitor c=0.0149844f //x=14.24 //y=0.71
c173 ( 57 0 ) capacitor c=0.0813322f //x=13.865 //y=1.915
c174 ( 56 0 ) capacitor c=0.0229267f //x=13.865 //y=1.52
c175 ( 55 0 ) capacitor c=0.0234352f //x=13.865 //y=1.21
c176 ( 54 0 ) capacitor c=0.0199343f //x=13.865 //y=0.865
c177 ( 53 0 ) capacitor c=0.110275f //x=14.4 //y=6.02
c178 ( 52 0 ) capacitor c=0.154305f //x=13.96 //y=6.02
c179 ( 50 0 ) capacitor c=0.00106608f //x=11.43 //y=5.155
c180 ( 49 0 ) capacitor c=0.00207319f //x=10.55 //y=5.155
c181 ( 42 0 ) capacitor c=0.0869732f //x=14.06 //y=2.08
c182 ( 40 0 ) capacitor c=0.107064f //x=12.21 //y=2.59
c183 ( 36 0 ) capacitor c=0.00398962f //x=11.81 //y=1.665
c184 ( 35 0 ) capacitor c=0.0137288f //x=12.125 //y=1.665
c185 ( 29 0 ) capacitor c=0.0284988f //x=12.125 //y=5.155
c186 ( 21 0 ) capacitor c=0.0176454f //x=11.345 //y=5.155
c187 ( 14 0 ) capacitor c=0.00332903f //x=9.755 //y=5.155
c188 ( 13 0 ) capacitor c=0.0148427f //x=10.465 //y=5.155
c189 ( 2 0 ) capacitor c=0.00808366f //x=12.325 //y=2.59
c190 ( 1 0 ) capacitor c=0.0353429f //x=13.945 //y=2.59
r191 (  75 77 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=13.96 //y=4.7 //x2=14.06 //y2=4.7
r192 (  68 77 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=14.4 //y=4.865 //x2=14.06 //y2=4.7
r193 (  67 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.395 //y=1.21 //x2=14.355 //y2=1.365
r194 (  66 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.395 //y=0.865 //x2=14.355 //y2=0.71
r195 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.395 //y=0.865 //x2=14.395 //y2=1.21
r196 (  64 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.02 //y=1.365 //x2=13.905 //y2=1.365
r197 (  63 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.24 //y=1.365 //x2=14.355 //y2=1.365
r198 (  62 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.02 //y=0.71 //x2=13.905 //y2=0.71
r199 (  61 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.24 //y=0.71 //x2=14.355 //y2=0.71
r200 (  61 62 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=14.24 //y=0.71 //x2=14.02 //y2=0.71
r201 (  58 75 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=13.96 //y=4.865 //x2=13.96 //y2=4.7
r202 (  57 72 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.915 //x2=14.06 //y2=2.08
r203 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.52 //x2=13.905 //y2=1.365
r204 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.52 //x2=13.865 //y2=1.915
r205 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.21 //x2=13.905 //y2=1.365
r206 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=0.865 //x2=13.905 //y2=0.71
r207 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.865 //y=0.865 //x2=13.865 //y2=1.21
r208 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.4 //y=6.02 //x2=14.4 //y2=4.865
r209 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.96 //y=6.02 //x2=13.96 //y2=4.865
r210 (  51 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.13 //y=1.365 //x2=14.24 //y2=1.365
r211 (  51 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.13 //y=1.365 //x2=14.02 //y2=1.365
r212 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=4.7 //x2=14.06 //y2=4.7
r213 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.59 //x2=14.06 //y2=4.7
r214 (  42 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=2.08 //x2=14.06 //y2=2.08
r215 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.08 //x2=14.06 //y2=2.59
r216 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=12.21 //y=5.07 //x2=12.21 //y2=2.59
r217 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.75 //x2=12.21 //y2=2.59
r218 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.665 //x2=12.21 //y2=1.75
r219 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.665 //x2=11.81 //y2=1.665
r220 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.725 //y=1.58 //x2=11.81 //y2=1.665
r221 (  31 80 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=11.725 //y=1.58 //x2=11.725 //y2=1.01
r222 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.515 //y=5.155 //x2=11.43 //y2=5.155
r223 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.155 //x2=12.21 //y2=5.07
r224 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.155 //x2=11.515 //y2=5.155
r225 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.43 //y=5.24 //x2=11.43 //y2=5.155
r226 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.43 //y=5.24 //x2=11.43 //y2=5.725
r227 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.635 //y=5.155 //x2=10.55 //y2=5.155
r228 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.345 //y=5.155 //x2=11.43 //y2=5.155
r229 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.345 //y=5.155 //x2=10.635 //y2=5.155
r230 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.55 //y=5.24 //x2=10.55 //y2=5.155
r231 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.55 //y=5.24 //x2=10.55 //y2=5.725
r232 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.465 //y=5.155 //x2=10.55 //y2=5.155
r233 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.465 //y=5.155 //x2=9.755 //y2=5.155
r234 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.67 //y=5.24 //x2=9.755 //y2=5.155
r235 (  7 82 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.67 //y=5.24 //x2=9.67 //y2=5.725
r236 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=2.59 //x2=14.06 //y2=2.59
r237 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.21 //y=2.59 //x2=12.21 //y2=2.59
r238 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.325 //y=2.59 //x2=12.21 //y2=2.59
r239 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=2.59 //x2=14.06 //y2=2.59
r240 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=13.945 //y=2.59 //x2=12.325 //y2=2.59
ends PM_TMRDFFSNQNX1\%noxref_4

subckt PM_TMRDFFSNQNX1\%noxref_5 ( 1 2 3 4 11 13 23 24 31 39 45 46 50 52 61 62 \
 64 65 67 68 69 70 71 72 73 74 75 80 82 84 90 91 92 93 94 95 99 101 104 105 \
 110 111 114 128 131 133 134 135 )
c278 ( 135 0 ) capacitor c=0.023087f //x=6.475 //y=5.02
c279 ( 134 0 ) capacitor c=0.023519f //x=5.595 //y=5.02
c280 ( 133 0 ) capacitor c=0.0224735f //x=4.715 //y=5.02
c281 ( 131 0 ) capacitor c=0.00853354f //x=6.725 //y=0.915
c282 ( 128 0 ) capacitor c=0.0588816f //x=17.39 //y=4.7
c283 ( 114 0 ) capacitor c=0.0331534f //x=1.88 //y=4.7
c284 ( 111 0 ) capacitor c=0.0279499f //x=1.85 //y=1.915
c285 ( 110 0 ) capacitor c=0.0422587f //x=1.85 //y=2.08
c286 ( 105 0 ) capacitor c=0.0318948f //x=17.725 //y=1.21
c287 ( 104 0 ) capacitor c=0.0187384f //x=17.725 //y=0.865
c288 ( 101 0 ) capacitor c=0.0141798f //x=17.57 //y=1.365
c289 ( 99 0 ) capacitor c=0.0149844f //x=17.57 //y=0.71
c290 ( 95 0 ) capacitor c=0.0813322f //x=17.195 //y=1.915
c291 ( 94 0 ) capacitor c=0.0229267f //x=17.195 //y=1.52
c292 ( 93 0 ) capacitor c=0.0234352f //x=17.195 //y=1.21
c293 ( 92 0 ) capacitor c=0.0199343f //x=17.195 //y=0.865
c294 ( 91 0 ) capacitor c=0.0429696f //x=2.415 //y=1.25
c295 ( 90 0 ) capacitor c=0.0192208f //x=2.415 //y=0.905
c296 ( 84 0 ) capacitor c=0.0158629f //x=2.26 //y=1.405
c297 ( 82 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c298 ( 80 0 ) capacitor c=0.0299681f //x=2.255 //y=4.79
c299 ( 75 0 ) capacitor c=0.0205163f //x=1.885 //y=1.56
c300 ( 74 0 ) capacitor c=0.0168481f //x=1.885 //y=1.25
c301 ( 73 0 ) capacitor c=0.0174783f //x=1.885 //y=0.905
c302 ( 72 0 ) capacitor c=0.110275f //x=17.73 //y=6.02
c303 ( 71 0 ) capacitor c=0.154305f //x=17.29 //y=6.02
c304 ( 70 0 ) capacitor c=0.15358f //x=2.33 //y=6.02
c305 ( 69 0 ) capacitor c=0.110281f //x=1.89 //y=6.02
c306 ( 65 0 ) capacitor c=0.0755336f //x=7.397 //y=3.905
c307 ( 64 0 ) capacitor c=0.0101843f //x=7.395 //y=4.07
c308 ( 62 0 ) capacitor c=0.00106608f //x=6.62 //y=5.155
c309 ( 61 0 ) capacitor c=0.00207162f //x=5.74 //y=5.155
c310 ( 52 0 ) capacitor c=0.0888543f //x=17.39 //y=2.08
c311 ( 50 0 ) capacitor c=0.0236247f //x=7.4 //y=5.07
c312 ( 46 0 ) capacitor c=0.00431225f //x=7 //y=1.665
c313 ( 45 0 ) capacitor c=0.0141453f //x=7.315 //y=1.665
c314 ( 39 0 ) capacitor c=0.0281378f //x=7.315 //y=5.155
c315 ( 31 0 ) capacitor c=0.0176454f //x=6.535 //y=5.155
c316 ( 24 0 ) capacitor c=0.00351598f //x=4.945 //y=5.155
c317 ( 23 0 ) capacitor c=0.0154196f //x=5.655 //y=5.155
c318 ( 13 0 ) capacitor c=0.0765924f //x=1.85 //y=2.08
c319 ( 11 0 ) capacitor c=0.00453889f //x=1.85 //y=4.535
c320 ( 4 0 ) capacitor c=0.00551102f //x=7.51 //y=4.07
c321 ( 3 0 ) capacitor c=0.141703f //x=17.275 //y=4.07
c322 ( 2 0 ) capacitor c=0.0165998f //x=1.965 //y=4.07
c323 ( 1 0 ) capacitor c=0.143583f //x=7.28 //y=4.07
r324 (  126 128 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=17.29 //y=4.7 //x2=17.39 //y2=4.7
r325 (  116 117 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.79 //x2=1.88 //y2=4.865
r326 (  114 116 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.7 //x2=1.88 //y2=4.79
r327 (  110 111 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r328 (  106 128 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=17.73 //y=4.865 //x2=17.39 //y2=4.7
r329 (  105 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.725 //y=1.21 //x2=17.685 //y2=1.365
r330 (  104 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.725 //y=0.865 //x2=17.685 //y2=0.71
r331 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.725 //y=0.865 //x2=17.725 //y2=1.21
r332 (  102 125 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.35 //y=1.365 //x2=17.235 //y2=1.365
r333 (  101 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.57 //y=1.365 //x2=17.685 //y2=1.365
r334 (  100 124 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.35 //y=0.71 //x2=17.235 //y2=0.71
r335 (  99 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.57 //y=0.71 //x2=17.685 //y2=0.71
r336 (  99 100 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.57 //y=0.71 //x2=17.35 //y2=0.71
r337 (  96 126 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.29 //y=4.865 //x2=17.29 //y2=4.7
r338 (  95 123 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.915 //x2=17.39 //y2=2.08
r339 (  94 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.52 //x2=17.235 //y2=1.365
r340 (  94 95 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.52 //x2=17.195 //y2=1.915
r341 (  93 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.21 //x2=17.235 //y2=1.365
r342 (  92 124 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=0.865 //x2=17.235 //y2=0.71
r343 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.195 //y=0.865 //x2=17.195 //y2=1.21
r344 (  91 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r345 (  90 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r346 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r347 (  85 119 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r348 (  84 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r349 (  83 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r350 (  82 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r351 (  82 83 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r352 (  81 116 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.015 //y=4.79 //x2=1.88 //y2=4.79
r353 (  80 87 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.33 //y2=4.865
r354 (  80 81 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.015 //y2=4.79
r355 (  75 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r356 (  75 111 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r357 (  74 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r358 (  73 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r359 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r360 (  72 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.73 //y=6.02 //x2=17.73 //y2=4.865
r361 (  71 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.29 //y=6.02 //x2=17.29 //y2=4.865
r362 (  70 87 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.02 //x2=2.33 //y2=4.865
r363 (  69 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.02 //x2=1.89 //y2=4.865
r364 (  68 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.46 //y=1.365 //x2=17.57 //y2=1.365
r365 (  68 102 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.46 //y=1.365 //x2=17.35 //y2=1.365
r366 (  67 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r367 (  67 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r368 (  64 66 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=7.397 //y=4.07 //x2=7.397 //y2=4.235
r369 (  64 65 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=7.397 //y=4.07 //x2=7.397 //y2=3.905
r370 (  60 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.88 //y=4.7 //x2=1.88 //y2=4.7
r371 (  57 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.39 //y=4.7 //x2=17.39 //y2=4.7
r372 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=17.39 //y=4.07 //x2=17.39 //y2=4.7
r373 (  52 123 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.39 //y=2.08 //x2=17.39 //y2=2.08
r374 (  52 55 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=17.39 //y=2.08 //x2=17.39 //y2=4.07
r375 (  50 66 ) resistor r=57.1551 //w=0.187 //l=0.835 //layer=li \
 //thickness=0.1 //x=7.4 //y=5.07 //x2=7.4 //y2=4.235
r376 (  47 65 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=7.4 //y=1.75 //x2=7.4 //y2=3.905
r377 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.665 //x2=7.4 //y2=1.75
r378 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.665 //x2=7 //y2=1.665
r379 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.915 //y=1.58 //x2=7 //y2=1.665
r380 (  41 131 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=6.915 //y=1.58 //x2=6.915 //y2=1.01
r381 (  40 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.705 //y=5.155 //x2=6.62 //y2=5.155
r382 (  39 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.155 //x2=7.4 //y2=5.07
r383 (  39 40 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.155 //x2=6.705 //y2=5.155
r384 (  33 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.62 //y=5.24 //x2=6.62 //y2=5.155
r385 (  33 135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.62 //y=5.24 //x2=6.62 //y2=5.725
r386 (  32 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.825 //y=5.155 //x2=5.74 //y2=5.155
r387 (  31 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.535 //y=5.155 //x2=6.62 //y2=5.155
r388 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.535 //y=5.155 //x2=5.825 //y2=5.155
r389 (  25 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.74 //y=5.24 //x2=5.74 //y2=5.155
r390 (  25 134 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=5.74 //y=5.24 //x2=5.74 //y2=5.725
r391 (  23 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.655 //y=5.155 //x2=5.74 //y2=5.155
r392 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.655 //y=5.155 //x2=4.945 //y2=5.155
r393 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.86 //y=5.24 //x2=4.945 //y2=5.155
r394 (  17 133 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.86 //y=5.24 //x2=4.86 //y2=5.725
r395 (  13 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r396 (  13 16 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.08 //x2=1.85 //y2=4.07
r397 (  11 60 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.865 //y2=4.7
r398 (  11 16 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.85 //y2=4.07
r399 (  10 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.39 //y=4.07 //x2=17.39 //y2=4.07
r400 (  8 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.395 //y=4.07 //x2=7.395 //y2=4.07
r401 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.85 //y=4.07 //x2=1.85 //y2=4.07
r402 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.51 //y=4.07 //x2=7.395 //y2=4.07
r403 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.275 //y=4.07 //x2=17.39 //y2=4.07
r404 (  3 4 ) resistor r=9.31775 //w=0.131 //l=9.765 //layer=m1 \
 //thickness=0.36 //x=17.275 //y=4.07 //x2=7.51 //y2=4.07
r405 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.965 //y=4.07 //x2=1.85 //y2=4.07
r406 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.28 //y=4.07 //x2=7.395 //y2=4.07
r407 (  1 2 ) resistor r=5.07156 //w=0.131 //l=5.315 //layer=m1 \
 //thickness=0.36 //x=7.28 //y=4.07 //x2=1.965 //y2=4.07
ends PM_TMRDFFSNQNX1\%noxref_5

subckt PM_TMRDFFSNQNX1\%noxref_6 ( 1 2 3 4 5 6 16 24 37 38 49 51 52 56 58 65 \
 66 67 68 69 70 71 72 73 74 78 79 80 85 87 90 91 95 96 97 102 104 107 108 112 \
 113 114 119 121 124 125 127 128 133 137 138 143 147 148 153 156 158 159 )
c324 ( 159 0 ) capacitor c=0.0220291f //x=14.915 //y=5.02
c325 ( 158 0 ) capacitor c=0.0217503f //x=14.035 //y=5.02
c326 ( 156 0 ) capacitor c=0.00866655f //x=14.91 //y=0.905
c327 ( 153 0 ) capacitor c=0.0587755f //x=22.94 //y=4.7
c328 ( 148 0 ) capacitor c=0.0273931f //x=22.94 //y=1.915
c329 ( 147 0 ) capacitor c=0.0456313f //x=22.94 //y=2.08
c330 ( 143 0 ) capacitor c=0.0587755f //x=11.47 //y=4.7
c331 ( 138 0 ) capacitor c=0.0273931f //x=11.47 //y=1.915
c332 ( 137 0 ) capacitor c=0.0456313f //x=11.47 //y=2.08
c333 ( 133 0 ) capacitor c=0.058931f //x=6.66 //y=4.7
c334 ( 128 0 ) capacitor c=0.0267105f //x=6.66 //y=1.915
c335 ( 127 0 ) capacitor c=0.0457054f //x=6.66 //y=2.08
c336 ( 125 0 ) capacitor c=0.0432517f //x=23.46 //y=1.26
c337 ( 124 0 ) capacitor c=0.0200379f //x=23.46 //y=0.915
c338 ( 121 0 ) capacitor c=0.0148873f //x=23.305 //y=1.415
c339 ( 119 0 ) capacitor c=0.0157803f //x=23.305 //y=0.76
c340 ( 114 0 ) capacitor c=0.0218028f //x=22.93 //y=1.57
c341 ( 113 0 ) capacitor c=0.0207459f //x=22.93 //y=1.26
c342 ( 112 0 ) capacitor c=0.0194308f //x=22.93 //y=0.915
c343 ( 108 0 ) capacitor c=0.0432517f //x=11.99 //y=1.26
c344 ( 107 0 ) capacitor c=0.0200379f //x=11.99 //y=0.915
c345 ( 104 0 ) capacitor c=0.0148873f //x=11.835 //y=1.415
c346 ( 102 0 ) capacitor c=0.0157803f //x=11.835 //y=0.76
c347 ( 97 0 ) capacitor c=0.0218028f //x=11.46 //y=1.57
c348 ( 96 0 ) capacitor c=0.0207459f //x=11.46 //y=1.26
c349 ( 95 0 ) capacitor c=0.0194308f //x=11.46 //y=0.915
c350 ( 91 0 ) capacitor c=0.0432517f //x=7.18 //y=1.26
c351 ( 90 0 ) capacitor c=0.0200379f //x=7.18 //y=0.915
c352 ( 87 0 ) capacitor c=0.0158629f //x=7.025 //y=1.415
c353 ( 85 0 ) capacitor c=0.0157803f //x=7.025 //y=0.76
c354 ( 80 0 ) capacitor c=0.0218028f //x=6.65 //y=1.57
c355 ( 79 0 ) capacitor c=0.0207459f //x=6.65 //y=1.26
c356 ( 78 0 ) capacitor c=0.0194308f //x=6.65 //y=0.915
c357 ( 74 0 ) capacitor c=0.158794f //x=23.12 //y=6.02
c358 ( 73 0 ) capacitor c=0.110114f //x=22.68 //y=6.02
c359 ( 72 0 ) capacitor c=0.158794f //x=11.65 //y=6.02
c360 ( 71 0 ) capacitor c=0.110114f //x=11.21 //y=6.02
c361 ( 70 0 ) capacitor c=0.158048f //x=6.84 //y=6.02
c362 ( 69 0 ) capacitor c=0.110114f //x=6.4 //y=6.02
c363 ( 65 0 ) capacitor c=0.00211606f //x=15.06 //y=5.2
c364 ( 58 0 ) capacitor c=0.0820102f //x=22.94 //y=2.08
c365 ( 56 0 ) capacitor c=0.106638f //x=15.54 //y=3.7
c366 ( 52 0 ) capacitor c=0.00404073f //x=15.185 //y=1.655
c367 ( 51 0 ) capacitor c=0.0122201f //x=15.455 //y=1.655
c368 ( 49 0 ) capacitor c=0.0137522f //x=15.455 //y=5.2
c369 ( 38 0 ) capacitor c=0.00251635f //x=14.265 //y=5.2
c370 ( 37 0 ) capacitor c=0.0142529f //x=14.975 //y=5.2
c371 ( 24 0 ) capacitor c=0.0834768f //x=11.47 //y=2.08
c372 ( 16 0 ) capacitor c=0.0842778f //x=6.66 //y=2.08
c373 ( 6 0 ) capacitor c=0.0043044f //x=15.655 //y=3.7
c374 ( 5 0 ) capacitor c=0.130401f //x=22.825 //y=3.7
c375 ( 4 0 ) capacitor c=0.00443912f //x=11.585 //y=3.7
c376 ( 3 0 ) capacitor c=0.0668348f //x=15.425 //y=3.7
c377 ( 2 0 ) capacitor c=0.0143354f //x=6.775 //y=3.7
c378 ( 1 0 ) capacitor c=0.0815699f //x=11.355 //y=3.7
r379 (  147 148 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=22.94 //y=2.08 //x2=22.94 //y2=1.915
r380 (  137 138 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11.47 //y=2.08 //x2=11.47 //y2=1.915
r381 (  127 128 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.66 //y=2.08 //x2=6.66 //y2=1.915
r382 (  125 155 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.46 //y=1.26 //x2=23.42 //y2=1.415
r383 (  124 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.46 //y=0.915 //x2=23.42 //y2=0.76
r384 (  124 125 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.46 //y=0.915 //x2=23.46 //y2=1.26
r385 (  122 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.085 //y=1.415 //x2=22.97 //y2=1.415
r386 (  121 155 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.305 //y=1.415 //x2=23.42 //y2=1.415
r387 (  120 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.085 //y=0.76 //x2=22.97 //y2=0.76
r388 (  119 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.305 //y=0.76 //x2=23.42 //y2=0.76
r389 (  119 120 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=23.305 //y=0.76 //x2=23.085 //y2=0.76
r390 (  116 153 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=23.12 //y=4.865 //x2=22.94 //y2=4.7
r391 (  114 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.57 //x2=22.97 //y2=1.415
r392 (  114 148 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.57 //x2=22.93 //y2=1.915
r393 (  113 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.26 //x2=22.97 //y2=1.415
r394 (  112 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=0.915 //x2=22.97 //y2=0.76
r395 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.93 //y=0.915 //x2=22.93 //y2=1.26
r396 (  109 153 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=22.68 //y=4.865 //x2=22.94 //y2=4.7
r397 (  108 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.99 //y=1.26 //x2=11.95 //y2=1.415
r398 (  107 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.99 //y=0.915 //x2=11.95 //y2=0.76
r399 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.99 //y=0.915 //x2=11.99 //y2=1.26
r400 (  105 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.615 //y=1.415 //x2=11.5 //y2=1.415
r401 (  104 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.835 //y=1.415 //x2=11.95 //y2=1.415
r402 (  103 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.615 //y=0.76 //x2=11.5 //y2=0.76
r403 (  102 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.835 //y=0.76 //x2=11.95 //y2=0.76
r404 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=11.835 //y=0.76 //x2=11.615 //y2=0.76
r405 (  99 143 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=11.65 //y=4.865 //x2=11.47 //y2=4.7
r406 (  97 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.57 //x2=11.5 //y2=1.415
r407 (  97 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.57 //x2=11.46 //y2=1.915
r408 (  96 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.26 //x2=11.5 //y2=1.415
r409 (  95 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=0.915 //x2=11.5 //y2=0.76
r410 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.46 //y=0.915 //x2=11.46 //y2=1.26
r411 (  92 143 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=11.21 //y=4.865 //x2=11.47 //y2=4.7
r412 (  91 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.18 //y=1.26 //x2=7.14 //y2=1.415
r413 (  90 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.18 //y=0.915 //x2=7.14 //y2=0.76
r414 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.18 //y=0.915 //x2=7.18 //y2=1.26
r415 (  88 131 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.805 //y=1.415 //x2=6.69 //y2=1.415
r416 (  87 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.025 //y=1.415 //x2=7.14 //y2=1.415
r417 (  86 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.805 //y=0.76 //x2=6.69 //y2=0.76
r418 (  85 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.025 //y=0.76 //x2=7.14 //y2=0.76
r419 (  85 86 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.025 //y=0.76 //x2=6.805 //y2=0.76
r420 (  82 133 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=6.84 //y=4.865 //x2=6.66 //y2=4.7
r421 (  80 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.57 //x2=6.69 //y2=1.415
r422 (  80 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.57 //x2=6.65 //y2=1.915
r423 (  79 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.26 //x2=6.69 //y2=1.415
r424 (  78 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=0.915 //x2=6.69 //y2=0.76
r425 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.65 //y=0.915 //x2=6.65 //y2=1.26
r426 (  75 133 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=6.4 //y=4.865 //x2=6.66 //y2=4.7
r427 (  74 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.12 //y=6.02 //x2=23.12 //y2=4.865
r428 (  73 109 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.68 //y=6.02 //x2=22.68 //y2=4.865
r429 (  72 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.65 //y=6.02 //x2=11.65 //y2=4.865
r430 (  71 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.21 //y=6.02 //x2=11.21 //y2=4.865
r431 (  70 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.84 //y=6.02 //x2=6.84 //y2=4.865
r432 (  69 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.4 //y=6.02 //x2=6.4 //y2=4.865
r433 (  68 121 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.195 //y=1.415 //x2=23.305 //y2=1.415
r434 (  68 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.195 //y=1.415 //x2=23.085 //y2=1.415
r435 (  67 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.725 //y=1.415 //x2=11.835 //y2=1.415
r436 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.725 //y=1.415 //x2=11.615 //y2=1.415
r437 (  66 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.915 //y=1.415 //x2=7.025 //y2=1.415
r438 (  66 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.915 //y=1.415 //x2=6.805 //y2=1.415
r439 (  63 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.94 //y=4.7 //x2=22.94 //y2=4.7
r440 (  61 63 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=22.94 //y=3.7 //x2=22.94 //y2=4.7
r441 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.94 //y=2.08 //x2=22.94 //y2=2.08
r442 (  58 61 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=22.94 //y=2.08 //x2=22.94 //y2=3.7
r443 (  54 56 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=15.54 //y=5.115 //x2=15.54 //y2=3.7
r444 (  53 56 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=15.54 //y=1.74 //x2=15.54 //y2=3.7
r445 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.455 //y=1.655 //x2=15.54 //y2=1.74
r446 (  51 52 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=15.455 //y=1.655 //x2=15.185 //y2=1.655
r447 (  50 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.145 //y=5.2 //x2=15.06 //y2=5.2
r448 (  49 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.455 //y=5.2 //x2=15.54 //y2=5.115
r449 (  49 50 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=15.455 //y=5.2 //x2=15.145 //y2=5.2
r450 (  45 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.1 //y=1.57 //x2=15.185 //y2=1.655
r451 (  45 156 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=15.1 //y=1.57 //x2=15.1 //y2=1
r452 (  39 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.06 //y=5.285 //x2=15.06 //y2=5.2
r453 (  39 159 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=15.06 //y=5.285 //x2=15.06 //y2=5.725
r454 (  37 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.975 //y=5.2 //x2=15.06 //y2=5.2
r455 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=14.975 //y=5.2 //x2=14.265 //y2=5.2
r456 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.18 //y=5.285 //x2=14.265 //y2=5.2
r457 (  31 158 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=14.18 //y=5.285 //x2=14.18 //y2=5.725
r458 (  29 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=4.7 //x2=11.47 //y2=4.7
r459 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=11.47 //y=3.7 //x2=11.47 //y2=4.7
r460 (  24 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=2.08 //x2=11.47 //y2=2.08
r461 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=11.47 //y=2.08 //x2=11.47 //y2=3.7
r462 (  21 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=4.7 //x2=6.66 //y2=4.7
r463 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=6.66 //y=3.7 //x2=6.66 //y2=4.7
r464 (  16 127 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.08 //x2=6.66 //y2=2.08
r465 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.08 //x2=6.66 //y2=3.7
r466 (  14 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=22.94 //y=3.7 //x2=22.94 //y2=3.7
r467 (  12 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=3.7 //x2=15.54 //y2=3.7
r468 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.47 //y=3.7 //x2=11.47 //y2=3.7
r469 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=3.7 //x2=6.66 //y2=3.7
r470 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.655 //y=3.7 //x2=15.54 //y2=3.7
r471 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=22.825 //y=3.7 //x2=22.94 //y2=3.7
r472 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=22.825 //y=3.7 //x2=15.655 //y2=3.7
r473 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.585 //y=3.7 //x2=11.47 //y2=3.7
r474 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=3.7 //x2=15.54 //y2=3.7
r475 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=3.7 //x2=11.585 //y2=3.7
r476 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.775 //y=3.7 //x2=6.66 //y2=3.7
r477 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=3.7 //x2=11.47 //y2=3.7
r478 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=3.7 //x2=6.775 //y2=3.7
ends PM_TMRDFFSNQNX1\%noxref_6

subckt PM_TMRDFFSNQNX1\%noxref_7 ( 1 2 7 9 19 20 27 35 41 42 46 49 50 51 52 53 \
 54 55 56 61 63 65 71 72 74 75 78 86 88 89 90 )
c183 ( 90 0 ) capacitor c=0.023087f //x=22.755 //y=5.02
c184 ( 89 0 ) capacitor c=0.023519f //x=21.875 //y=5.02
c185 ( 88 0 ) capacitor c=0.0224735f //x=20.995 //y=5.02
c186 ( 86 0 ) capacitor c=0.00872971f //x=23.005 //y=0.915
c187 ( 78 0 ) capacitor c=0.0331095f //x=18.16 //y=4.7
c188 ( 75 0 ) capacitor c=0.0279499f //x=18.13 //y=1.915
c189 ( 74 0 ) capacitor c=0.0421676f //x=18.13 //y=2.08
c190 ( 72 0 ) capacitor c=0.0429696f //x=18.695 //y=1.25
c191 ( 71 0 ) capacitor c=0.0192208f //x=18.695 //y=0.905
c192 ( 65 0 ) capacitor c=0.0148884f //x=18.54 //y=1.405
c193 ( 63 0 ) capacitor c=0.0157803f //x=18.54 //y=0.75
c194 ( 61 0 ) capacitor c=0.0295235f //x=18.535 //y=4.79
c195 ( 56 0 ) capacitor c=0.0205163f //x=18.165 //y=1.56
c196 ( 55 0 ) capacitor c=0.0168481f //x=18.165 //y=1.25
c197 ( 54 0 ) capacitor c=0.0174783f //x=18.165 //y=0.905
c198 ( 53 0 ) capacitor c=0.15358f //x=18.61 //y=6.02
c199 ( 52 0 ) capacitor c=0.110281f //x=18.17 //y=6.02
c200 ( 50 0 ) capacitor c=0.00106608f //x=22.9 //y=5.155
c201 ( 49 0 ) capacitor c=0.00207319f //x=22.02 //y=5.155
c202 ( 46 0 ) capacitor c=0.108218f //x=23.68 //y=4.07
c203 ( 42 0 ) capacitor c=0.00398962f //x=23.28 //y=1.665
c204 ( 41 0 ) capacitor c=0.0137288f //x=23.595 //y=1.665
c205 ( 35 0 ) capacitor c=0.0284988f //x=23.595 //y=5.155
c206 ( 27 0 ) capacitor c=0.0176454f //x=22.815 //y=5.155
c207 ( 20 0 ) capacitor c=0.00332903f //x=21.225 //y=5.155
c208 ( 19 0 ) capacitor c=0.0148427f //x=21.935 //y=5.155
c209 ( 9 0 ) capacitor c=0.0709461f //x=18.13 //y=2.08
c210 ( 7 0 ) capacitor c=0.00453889f //x=18.13 //y=4.535
c211 ( 2 0 ) capacitor c=0.00621861f //x=18.245 //y=4.07
c212 ( 1 0 ) capacitor c=0.0857087f //x=23.565 //y=4.07
r213 (  80 81 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=18.16 //y=4.79 //x2=18.16 //y2=4.865
r214 (  78 80 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=18.16 //y=4.7 //x2=18.16 //y2=4.79
r215 (  74 75 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=18.13 //y=2.08 //x2=18.13 //y2=1.915
r216 (  72 85 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.695 //y=1.25 //x2=18.655 //y2=1.405
r217 (  71 84 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.695 //y=0.905 //x2=18.655 //y2=0.75
r218 (  71 72 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.695 //y=0.905 //x2=18.695 //y2=1.25
r219 (  66 83 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.32 //y=1.405 //x2=18.205 //y2=1.405
r220 (  65 85 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.54 //y=1.405 //x2=18.655 //y2=1.405
r221 (  64 82 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.32 //y=0.75 //x2=18.205 //y2=0.75
r222 (  63 84 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.54 //y=0.75 //x2=18.655 //y2=0.75
r223 (  63 64 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.54 //y=0.75 //x2=18.32 //y2=0.75
r224 (  62 80 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=18.295 //y=4.79 //x2=18.16 //y2=4.79
r225 (  61 68 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.79 //x2=18.61 //y2=4.865
r226 (  61 62 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.79 //x2=18.295 //y2=4.79
r227 (  56 83 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.56 //x2=18.205 //y2=1.405
r228 (  56 75 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.56 //x2=18.165 //y2=1.915
r229 (  55 83 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.25 //x2=18.205 //y2=1.405
r230 (  54 82 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=0.905 //x2=18.205 //y2=0.75
r231 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.165 //y=0.905 //x2=18.165 //y2=1.25
r232 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.61 //y=6.02 //x2=18.61 //y2=4.865
r233 (  52 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.17 //y=6.02 //x2=18.17 //y2=4.865
r234 (  51 65 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.43 //y=1.405 //x2=18.54 //y2=1.405
r235 (  51 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.43 //y=1.405 //x2=18.32 //y2=1.405
r236 (  48 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.16 //y=4.7 //x2=18.16 //y2=4.7
r237 (  44 46 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=23.68 //y=5.07 //x2=23.68 //y2=4.07
r238 (  43 46 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=23.68 //y=1.75 //x2=23.68 //y2=4.07
r239 (  41 43 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.595 //y=1.665 //x2=23.68 //y2=1.75
r240 (  41 42 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=23.595 //y=1.665 //x2=23.28 //y2=1.665
r241 (  37 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.195 //y=1.58 //x2=23.28 //y2=1.665
r242 (  37 86 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.195 //y=1.58 //x2=23.195 //y2=1.01
r243 (  36 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.985 //y=5.155 //x2=22.9 //y2=5.155
r244 (  35 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.595 //y=5.155 //x2=23.68 //y2=5.07
r245 (  35 36 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=23.595 //y=5.155 //x2=22.985 //y2=5.155
r246 (  29 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.9 //y=5.24 //x2=22.9 //y2=5.155
r247 (  29 90 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.9 //y=5.24 //x2=22.9 //y2=5.725
r248 (  28 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.105 //y=5.155 //x2=22.02 //y2=5.155
r249 (  27 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.815 //y=5.155 //x2=22.9 //y2=5.155
r250 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.815 //y=5.155 //x2=22.105 //y2=5.155
r251 (  21 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.02 //y=5.24 //x2=22.02 //y2=5.155
r252 (  21 89 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.02 //y=5.24 //x2=22.02 //y2=5.725
r253 (  19 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.935 //y=5.155 //x2=22.02 //y2=5.155
r254 (  19 20 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=21.935 //y=5.155 //x2=21.225 //y2=5.155
r255 (  13 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.14 //y=5.24 //x2=21.225 //y2=5.155
r256 (  13 88 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.14 //y=5.24 //x2=21.14 //y2=5.725
r257 (  9 74 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.13 //y=2.08 //x2=18.13 //y2=2.08
r258 (  9 12 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=18.13 //y=2.08 //x2=18.13 //y2=4.07
r259 (  7 48 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.535 //x2=18.145 //y2=4.7
r260 (  7 12 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.535 //x2=18.13 //y2=4.07
r261 (  6 46 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.68 //y=4.07 //x2=23.68 //y2=4.07
r262 (  4 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.13 //y=4.07 //x2=18.13 //y2=4.07
r263 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.245 //y=4.07 //x2=18.13 //y2=4.07
r264 (  1 6 ) resistor r=0.0738079 //w=0.207 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.565 //y=4.07 //x2=23.68 //y2=4.07
r265 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=23.565 //y=4.07 //x2=18.245 //y2=4.07
ends PM_TMRDFFSNQNX1\%noxref_7

subckt PM_TMRDFFSNQNX1\%noxref_8 ( 1 2 3 4 17 18 29 31 32 36 38 46 53 54 55 56 \
 57 58 59 60 61 62 63 64 66 72 73 74 75 79 80 81 82 83 85 91 92 93 94 114 116 \
 117 )
c232 ( 117 0 ) capacitor c=0.0220291f //x=26.385 //y=5.02
c233 ( 116 0 ) capacitor c=0.0217503f //x=25.505 //y=5.02
c234 ( 114 0 ) capacitor c=0.0084702f //x=26.38 //y=0.905
c235 ( 94 0 ) capacitor c=0.0556143f //x=33.945 //y=4.79
c236 ( 93 0 ) capacitor c=0.0293157f //x=34.235 //y=4.79
c237 ( 92 0 ) capacitor c=0.0347816f //x=33.9 //y=1.22
c238 ( 91 0 ) capacitor c=0.0187487f //x=33.9 //y=0.875
c239 ( 85 0 ) capacitor c=0.0137055f //x=33.745 //y=1.375
c240 ( 83 0 ) capacitor c=0.0149861f //x=33.745 //y=0.72
c241 ( 82 0 ) capacitor c=0.096037f //x=33.37 //y=1.915
c242 ( 81 0 ) capacitor c=0.0228993f //x=33.37 //y=1.53
c243 ( 80 0 ) capacitor c=0.0234352f //x=33.37 //y=1.22
c244 ( 79 0 ) capacitor c=0.0198724f //x=33.37 //y=0.875
c245 ( 75 0 ) capacitor c=0.0557698f //x=29.135 //y=4.79
c246 ( 74 0 ) capacitor c=0.0293157f //x=29.425 //y=4.79
c247 ( 73 0 ) capacitor c=0.0347816f //x=29.09 //y=1.22
c248 ( 72 0 ) capacitor c=0.0187487f //x=29.09 //y=0.875
c249 ( 66 0 ) capacitor c=0.0137055f //x=28.935 //y=1.375
c250 ( 64 0 ) capacitor c=0.0149861f //x=28.935 //y=0.72
c251 ( 63 0 ) capacitor c=0.096037f //x=28.56 //y=1.915
c252 ( 62 0 ) capacitor c=0.0228993f //x=28.56 //y=1.53
c253 ( 61 0 ) capacitor c=0.0234352f //x=28.56 //y=1.22
c254 ( 60 0 ) capacitor c=0.0198724f //x=28.56 //y=0.875
c255 ( 59 0 ) capacitor c=0.110114f //x=34.31 //y=6.02
c256 ( 58 0 ) capacitor c=0.158956f //x=33.87 //y=6.02
c257 ( 57 0 ) capacitor c=0.110114f //x=29.5 //y=6.02
c258 ( 56 0 ) capacitor c=0.158956f //x=29.06 //y=6.02
c259 ( 53 0 ) capacitor c=0.00211606f //x=26.53 //y=5.2
c260 ( 46 0 ) capacitor c=0.0943831f //x=33.67 //y=2.08
c261 ( 38 0 ) capacitor c=0.0969522f //x=28.86 //y=2.08
c262 ( 36 0 ) capacitor c=0.105125f //x=27.01 //y=2.59
c263 ( 32 0 ) capacitor c=0.00404073f //x=26.655 //y=1.655
c264 ( 31 0 ) capacitor c=0.0122201f //x=26.925 //y=1.655
c265 ( 29 0 ) capacitor c=0.0137995f //x=26.925 //y=5.2
c266 ( 18 0 ) capacitor c=0.00251635f //x=25.735 //y=5.2
c267 ( 17 0 ) capacitor c=0.0143649f //x=26.445 //y=5.2
c268 ( 4 0 ) capacitor c=0.00673266f //x=29.125 //y=2.59
c269 ( 3 0 ) capacitor c=0.0686809f //x=33.555 //y=2.59
c270 ( 2 0 ) capacitor c=0.0121637f //x=27.125 //y=2.59
c271 ( 1 0 ) capacitor c=0.0230071f //x=28.715 //y=2.59
r272 (  93 95 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=34.235 //y=4.79 //x2=34.31 //y2=4.865
r273 (  93 94 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=34.235 //y=4.79 //x2=33.945 //y2=4.79
r274 (  92 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.9 //y=1.22 //x2=33.86 //y2=1.375
r275 (  91 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.9 //y=0.875 //x2=33.86 //y2=0.72
r276 (  91 92 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=33.9 //y=0.875 //x2=33.9 //y2=1.22
r277 (  88 94 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=33.87 //y=4.865 //x2=33.945 //y2=4.79
r278 (  88 111 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=33.87 //y=4.865 //x2=33.67 //y2=4.7
r279 (  86 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=33.525 //y=1.375 //x2=33.41 //y2=1.375
r280 (  85 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=33.745 //y=1.375 //x2=33.86 //y2=1.375
r281 (  84 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=33.525 //y=0.72 //x2=33.41 //y2=0.72
r282 (  83 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=33.745 //y=0.72 //x2=33.86 //y2=0.72
r283 (  83 84 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=33.745 //y=0.72 //x2=33.525 //y2=0.72
r284 (  82 109 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=33.37 //y=1.915 //x2=33.67 //y2=2.08
r285 (  81 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.37 //y=1.53 //x2=33.41 //y2=1.375
r286 (  81 82 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=33.37 //y=1.53 //x2=33.37 //y2=1.915
r287 (  80 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.37 //y=1.22 //x2=33.41 //y2=1.375
r288 (  79 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.37 //y=0.875 //x2=33.41 //y2=0.72
r289 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=33.37 //y=0.875 //x2=33.37 //y2=1.22
r290 (  74 76 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=29.425 //y=4.79 //x2=29.5 //y2=4.865
r291 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=29.425 //y=4.79 //x2=29.135 //y2=4.79
r292 (  73 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.09 //y=1.22 //x2=29.05 //y2=1.375
r293 (  72 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.09 //y=0.875 //x2=29.05 //y2=0.72
r294 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=29.09 //y=0.875 //x2=29.09 //y2=1.22
r295 (  69 75 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=29.06 //y=4.865 //x2=29.135 //y2=4.79
r296 (  69 103 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=29.06 //y=4.865 //x2=28.86 //y2=4.7
r297 (  67 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.715 //y=1.375 //x2=28.6 //y2=1.375
r298 (  66 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.935 //y=1.375 //x2=29.05 //y2=1.375
r299 (  65 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.715 //y=0.72 //x2=28.6 //y2=0.72
r300 (  64 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.935 //y=0.72 //x2=29.05 //y2=0.72
r301 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=28.935 //y=0.72 //x2=28.715 //y2=0.72
r302 (  63 101 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=28.56 //y=1.915 //x2=28.86 //y2=2.08
r303 (  62 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.56 //y=1.53 //x2=28.6 //y2=1.375
r304 (  62 63 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=28.56 //y=1.53 //x2=28.56 //y2=1.915
r305 (  61 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.56 //y=1.22 //x2=28.6 //y2=1.375
r306 (  60 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.56 //y=0.875 //x2=28.6 //y2=0.72
r307 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=28.56 //y=0.875 //x2=28.56 //y2=1.22
r308 (  59 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.31 //y=6.02 //x2=34.31 //y2=4.865
r309 (  58 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=33.87 //y=6.02 //x2=33.87 //y2=4.865
r310 (  57 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=29.5 //y=6.02 //x2=29.5 //y2=4.865
r311 (  56 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=29.06 //y=6.02 //x2=29.06 //y2=4.865
r312 (  55 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=33.635 //y=1.375 //x2=33.745 //y2=1.375
r313 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=33.635 //y=1.375 //x2=33.525 //y2=1.375
r314 (  54 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=28.825 //y=1.375 //x2=28.935 //y2=1.375
r315 (  54 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=28.825 //y=1.375 //x2=28.715 //y2=1.375
r316 (  51 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=33.67 //y=4.7 //x2=33.67 //y2=4.7
r317 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=33.67 //y=2.59 //x2=33.67 //y2=4.7
r318 (  46 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=33.67 //y=2.08 //x2=33.67 //y2=2.08
r319 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=33.67 //y=2.08 //x2=33.67 //y2=2.59
r320 (  43 103 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.86 //y=4.7 //x2=28.86 //y2=4.7
r321 (  41 43 ) resistor r=144.77 //w=0.187 //l=2.115 //layer=li \
 //thickness=0.1 //x=28.86 //y=2.585 //x2=28.86 //y2=4.7
r322 (  38 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.86 //y=2.08 //x2=28.86 //y2=2.08
r323 (  38 41 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=28.86 //y=2.08 //x2=28.86 //y2=2.585
r324 (  34 36 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=27.01 //y=5.115 //x2=27.01 //y2=2.59
r325 (  33 36 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=27.01 //y=1.74 //x2=27.01 //y2=2.59
r326 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.925 //y=1.655 //x2=27.01 //y2=1.74
r327 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=26.925 //y=1.655 //x2=26.655 //y2=1.655
r328 (  30 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.615 //y=5.2 //x2=26.53 //y2=5.2
r329 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.925 //y=5.2 //x2=27.01 //y2=5.115
r330 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=26.925 //y=5.2 //x2=26.615 //y2=5.2
r331 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.57 //y=1.57 //x2=26.655 //y2=1.655
r332 (  25 114 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=26.57 //y=1.57 //x2=26.57 //y2=1
r333 (  19 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.53 //y=5.285 //x2=26.53 //y2=5.2
r334 (  19 117 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=26.53 //y=5.285 //x2=26.53 //y2=5.725
r335 (  17 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.445 //y=5.2 //x2=26.53 //y2=5.2
r336 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.445 //y=5.2 //x2=25.735 //y2=5.2
r337 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.65 //y=5.285 //x2=25.735 //y2=5.2
r338 (  11 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=25.65 //y=5.285 //x2=25.65 //y2=5.725
r339 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=33.67 //y=2.59 //x2=33.67 //y2=2.59
r340 (  8 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.86 //y=2.585 //x2=28.86 //y2=2.585
r341 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=27.01 //y=2.59 //x2=27.01 //y2=2.59
r342 (  4 8 ) resistor r=0.164988 //w=0.206 //l=0.267488 //layer=m1 \
 //thickness=0.36 //x=29.125 //y=2.59 //x2=28.86 //y2=2.585
r343 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=33.555 //y=2.59 //x2=33.67 //y2=2.59
r344 (  3 4 ) resistor r=4.2271 //w=0.131 //l=4.43 //layer=m1 //thickness=0.36 \
 //x=33.555 //y=2.59 //x2=29.125 //y2=2.59
r345 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.125 //y=2.59 //x2=27.01 //y2=2.59
r346 (  1 8 ) resistor r=0.0921728 //w=0.206 //l=0.147479 //layer=m1 \
 //thickness=0.36 //x=28.715 //y=2.59 //x2=28.86 //y2=2.585
r347 (  1 2 ) resistor r=1.51718 //w=0.131 //l=1.59 //layer=m1 \
 //thickness=0.36 //x=28.715 //y=2.59 //x2=27.125 //y2=2.59
ends PM_TMRDFFSNQNX1\%noxref_8

subckt PM_TMRDFFSNQNX1\%noxref_9 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 61 63 66 67 77 80 82 83 84 )
c166 ( 84 0 ) capacitor c=0.023087f //x=35.705 //y=5.02
c167 ( 83 0 ) capacitor c=0.023519f //x=34.825 //y=5.02
c168 ( 82 0 ) capacitor c=0.0224735f //x=33.945 //y=5.02
c169 ( 80 0 ) capacitor c=0.00872971f //x=35.955 //y=0.915
c170 ( 77 0 ) capacitor c=0.0588816f //x=38.48 //y=4.7
c171 ( 67 0 ) capacitor c=0.0318948f //x=38.815 //y=1.21
c172 ( 66 0 ) capacitor c=0.0187384f //x=38.815 //y=0.865
c173 ( 63 0 ) capacitor c=0.0141798f //x=38.66 //y=1.365
c174 ( 61 0 ) capacitor c=0.0149844f //x=38.66 //y=0.71
c175 ( 57 0 ) capacitor c=0.0813322f //x=38.285 //y=1.915
c176 ( 56 0 ) capacitor c=0.0229267f //x=38.285 //y=1.52
c177 ( 55 0 ) capacitor c=0.0234352f //x=38.285 //y=1.21
c178 ( 54 0 ) capacitor c=0.0199343f //x=38.285 //y=0.865
c179 ( 53 0 ) capacitor c=0.110275f //x=38.82 //y=6.02
c180 ( 52 0 ) capacitor c=0.154305f //x=38.38 //y=6.02
c181 ( 50 0 ) capacitor c=0.00106608f //x=35.85 //y=5.155
c182 ( 49 0 ) capacitor c=0.00207319f //x=34.97 //y=5.155
c183 ( 42 0 ) capacitor c=0.0839295f //x=38.48 //y=2.08
c184 ( 40 0 ) capacitor c=0.10402f //x=36.63 //y=2.59
c185 ( 36 0 ) capacitor c=0.00398962f //x=36.23 //y=1.665
c186 ( 35 0 ) capacitor c=0.0137288f //x=36.545 //y=1.665
c187 ( 29 0 ) capacitor c=0.0284988f //x=36.545 //y=5.155
c188 ( 21 0 ) capacitor c=0.0176454f //x=35.765 //y=5.155
c189 ( 14 0 ) capacitor c=0.00332903f //x=34.175 //y=5.155
c190 ( 13 0 ) capacitor c=0.0148427f //x=34.885 //y=5.155
c191 ( 2 0 ) capacitor c=0.00808366f //x=36.745 //y=2.59
c192 ( 1 0 ) capacitor c=0.0353429f //x=38.365 //y=2.59
r193 (  75 77 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=38.38 //y=4.7 //x2=38.48 //y2=4.7
r194 (  68 77 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=38.82 //y=4.865 //x2=38.48 //y2=4.7
r195 (  67 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.815 //y=1.21 //x2=38.775 //y2=1.365
r196 (  66 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.815 //y=0.865 //x2=38.775 //y2=0.71
r197 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=38.815 //y=0.865 //x2=38.815 //y2=1.21
r198 (  64 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.44 //y=1.365 //x2=38.325 //y2=1.365
r199 (  63 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.66 //y=1.365 //x2=38.775 //y2=1.365
r200 (  62 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.44 //y=0.71 //x2=38.325 //y2=0.71
r201 (  61 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.66 //y=0.71 //x2=38.775 //y2=0.71
r202 (  61 62 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=38.66 //y=0.71 //x2=38.44 //y2=0.71
r203 (  58 75 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=38.38 //y=4.865 //x2=38.38 //y2=4.7
r204 (  57 72 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=38.285 //y=1.915 //x2=38.48 //y2=2.08
r205 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.285 //y=1.52 //x2=38.325 //y2=1.365
r206 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=38.285 //y=1.52 //x2=38.285 //y2=1.915
r207 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.285 //y=1.21 //x2=38.325 //y2=1.365
r208 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.285 //y=0.865 //x2=38.325 //y2=0.71
r209 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=38.285 //y=0.865 //x2=38.285 //y2=1.21
r210 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=38.82 //y=6.02 //x2=38.82 //y2=4.865
r211 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=38.38 //y=6.02 //x2=38.38 //y2=4.865
r212 (  51 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=38.55 //y=1.365 //x2=38.66 //y2=1.365
r213 (  51 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=38.55 //y=1.365 //x2=38.44 //y2=1.365
r214 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=38.48 //y=4.7 //x2=38.48 //y2=4.7
r215 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=38.48 //y=2.59 //x2=38.48 //y2=4.7
r216 (  42 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=38.48 //y=2.08 //x2=38.48 //y2=2.08
r217 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=38.48 //y=2.08 //x2=38.48 //y2=2.59
r218 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=36.63 //y=5.07 //x2=36.63 //y2=2.59
r219 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=36.63 //y=1.75 //x2=36.63 //y2=2.59
r220 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=36.545 //y=1.665 //x2=36.63 //y2=1.75
r221 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=36.545 //y=1.665 //x2=36.23 //y2=1.665
r222 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=36.145 //y=1.58 //x2=36.23 //y2=1.665
r223 (  31 80 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=36.145 //y=1.58 //x2=36.145 //y2=1.01
r224 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.935 //y=5.155 //x2=35.85 //y2=5.155
r225 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=36.545 //y=5.155 //x2=36.63 //y2=5.07
r226 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=36.545 //y=5.155 //x2=35.935 //y2=5.155
r227 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.85 //y=5.24 //x2=35.85 //y2=5.155
r228 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.85 //y=5.24 //x2=35.85 //y2=5.725
r229 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.055 //y=5.155 //x2=34.97 //y2=5.155
r230 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.765 //y=5.155 //x2=35.85 //y2=5.155
r231 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=35.765 //y=5.155 //x2=35.055 //y2=5.155
r232 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.97 //y=5.24 //x2=34.97 //y2=5.155
r233 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=34.97 //y=5.24 //x2=34.97 //y2=5.725
r234 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.885 //y=5.155 //x2=34.97 //y2=5.155
r235 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=34.885 //y=5.155 //x2=34.175 //y2=5.155
r236 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.09 //y=5.24 //x2=34.175 //y2=5.155
r237 (  7 82 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=34.09 //y=5.24 //x2=34.09 //y2=5.725
r238 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=38.48 //y=2.59 //x2=38.48 //y2=2.59
r239 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=36.63 //y=2.59 //x2=36.63 //y2=2.59
r240 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=36.745 //y=2.59 //x2=36.63 //y2=2.59
r241 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=38.365 //y=2.59 //x2=38.48 //y2=2.59
r242 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=38.365 //y=2.59 //x2=36.745 //y2=2.59
ends PM_TMRDFFSNQNX1\%noxref_9

subckt PM_TMRDFFSNQNX1\%noxref_10 ( 1 2 3 4 11 13 23 24 31 39 45 46 50 52 61 \
 62 64 65 67 68 69 70 71 72 73 74 75 80 82 84 90 91 92 93 94 95 99 101 104 105 \
 110 111 114 128 131 133 134 135 )
c282 ( 135 0 ) capacitor c=0.023087f //x=30.895 //y=5.02
c283 ( 134 0 ) capacitor c=0.023519f //x=30.015 //y=5.02
c284 ( 133 0 ) capacitor c=0.0224735f //x=29.135 //y=5.02
c285 ( 131 0 ) capacitor c=0.00853354f //x=31.145 //y=0.915
c286 ( 128 0 ) capacitor c=0.0588816f //x=41.81 //y=4.7
c287 ( 114 0 ) capacitor c=0.0331095f //x=26.3 //y=4.7
c288 ( 111 0 ) capacitor c=0.0279499f //x=26.27 //y=1.915
c289 ( 110 0 ) capacitor c=0.0421676f //x=26.27 //y=2.08
c290 ( 105 0 ) capacitor c=0.0318948f //x=42.145 //y=1.21
c291 ( 104 0 ) capacitor c=0.0187384f //x=42.145 //y=0.865
c292 ( 101 0 ) capacitor c=0.0141798f //x=41.99 //y=1.365
c293 ( 99 0 ) capacitor c=0.0149844f //x=41.99 //y=0.71
c294 ( 95 0 ) capacitor c=0.0813322f //x=41.615 //y=1.915
c295 ( 94 0 ) capacitor c=0.0229267f //x=41.615 //y=1.52
c296 ( 93 0 ) capacitor c=0.0234352f //x=41.615 //y=1.21
c297 ( 92 0 ) capacitor c=0.0199343f //x=41.615 //y=0.865
c298 ( 91 0 ) capacitor c=0.0429696f //x=26.835 //y=1.25
c299 ( 90 0 ) capacitor c=0.0192208f //x=26.835 //y=0.905
c300 ( 84 0 ) capacitor c=0.0148884f //x=26.68 //y=1.405
c301 ( 82 0 ) capacitor c=0.0157803f //x=26.68 //y=0.75
c302 ( 80 0 ) capacitor c=0.0295235f //x=26.675 //y=4.79
c303 ( 75 0 ) capacitor c=0.0205163f //x=26.305 //y=1.56
c304 ( 74 0 ) capacitor c=0.0168481f //x=26.305 //y=1.25
c305 ( 73 0 ) capacitor c=0.0174783f //x=26.305 //y=0.905
c306 ( 72 0 ) capacitor c=0.110275f //x=42.15 //y=6.02
c307 ( 71 0 ) capacitor c=0.154305f //x=41.71 //y=6.02
c308 ( 70 0 ) capacitor c=0.15358f //x=26.75 //y=6.02
c309 ( 69 0 ) capacitor c=0.110281f //x=26.31 //y=6.02
c310 ( 65 0 ) capacitor c=0.0715637f //x=31.817 //y=3.905
c311 ( 64 0 ) capacitor c=0.0101843f //x=31.815 //y=4.07
c312 ( 62 0 ) capacitor c=0.00106608f //x=31.04 //y=5.155
c313 ( 61 0 ) capacitor c=0.00207162f //x=30.16 //y=5.155
c314 ( 52 0 ) capacitor c=0.0857541f //x=41.81 //y=2.08
c315 ( 50 0 ) capacitor c=0.0236247f //x=31.82 //y=5.07
c316 ( 46 0 ) capacitor c=0.00398962f //x=31.42 //y=1.665
c317 ( 45 0 ) capacitor c=0.0135805f //x=31.735 //y=1.665
c318 ( 39 0 ) capacitor c=0.0281378f //x=31.735 //y=5.155
c319 ( 31 0 ) capacitor c=0.0176454f //x=30.955 //y=5.155
c320 ( 24 0 ) capacitor c=0.00332903f //x=29.365 //y=5.155
c321 ( 23 0 ) capacitor c=0.014837f //x=30.075 //y=5.155
c322 ( 13 0 ) capacitor c=0.0709324f //x=26.27 //y=2.08
c323 ( 11 0 ) capacitor c=0.00453889f //x=26.27 //y=4.535
c324 ( 4 0 ) capacitor c=0.00551102f //x=31.93 //y=4.07
c325 ( 3 0 ) capacitor c=0.141703f //x=41.695 //y=4.07
c326 ( 2 0 ) capacitor c=0.00979524f //x=26.385 //y=4.07
c327 ( 1 0 ) capacitor c=0.0882171f //x=31.7 //y=4.07
r328 (  126 128 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=41.71 //y=4.7 //x2=41.81 //y2=4.7
r329 (  116 117 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=26.3 //y=4.79 //x2=26.3 //y2=4.865
r330 (  114 116 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=26.3 //y=4.7 //x2=26.3 //y2=4.79
r331 (  110 111 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=26.27 //y=2.08 //x2=26.27 //y2=1.915
r332 (  106 128 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=42.15 //y=4.865 //x2=41.81 //y2=4.7
r333 (  105 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.145 //y=1.21 //x2=42.105 //y2=1.365
r334 (  104 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.145 //y=0.865 //x2=42.105 //y2=0.71
r335 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.145 //y=0.865 //x2=42.145 //y2=1.21
r336 (  102 125 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.77 //y=1.365 //x2=41.655 //y2=1.365
r337 (  101 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.99 //y=1.365 //x2=42.105 //y2=1.365
r338 (  100 124 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.77 //y=0.71 //x2=41.655 //y2=0.71
r339 (  99 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.99 //y=0.71 //x2=42.105 //y2=0.71
r340 (  99 100 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=41.99 //y=0.71 //x2=41.77 //y2=0.71
r341 (  96 126 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=41.71 //y=4.865 //x2=41.71 //y2=4.7
r342 (  95 123 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=41.615 //y=1.915 //x2=41.81 //y2=2.08
r343 (  94 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.615 //y=1.52 //x2=41.655 //y2=1.365
r344 (  94 95 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=41.615 //y=1.52 //x2=41.615 //y2=1.915
r345 (  93 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.615 //y=1.21 //x2=41.655 //y2=1.365
r346 (  92 124 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.615 //y=0.865 //x2=41.655 //y2=0.71
r347 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=41.615 //y=0.865 //x2=41.615 //y2=1.21
r348 (  91 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.835 //y=1.25 //x2=26.795 //y2=1.405
r349 (  90 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.835 //y=0.905 //x2=26.795 //y2=0.75
r350 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=26.835 //y=0.905 //x2=26.835 //y2=1.25
r351 (  85 119 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.46 //y=1.405 //x2=26.345 //y2=1.405
r352 (  84 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.68 //y=1.405 //x2=26.795 //y2=1.405
r353 (  83 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.46 //y=0.75 //x2=26.345 //y2=0.75
r354 (  82 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.68 //y=0.75 //x2=26.795 //y2=0.75
r355 (  82 83 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=26.68 //y=0.75 //x2=26.46 //y2=0.75
r356 (  81 116 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=26.435 //y=4.79 //x2=26.3 //y2=4.79
r357 (  80 87 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=26.675 //y=4.79 //x2=26.75 //y2=4.865
r358 (  80 81 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=26.675 //y=4.79 //x2=26.435 //y2=4.79
r359 (  75 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.305 //y=1.56 //x2=26.345 //y2=1.405
r360 (  75 111 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=26.305 //y=1.56 //x2=26.305 //y2=1.915
r361 (  74 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.305 //y=1.25 //x2=26.345 //y2=1.405
r362 (  73 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.305 //y=0.905 //x2=26.345 //y2=0.75
r363 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=26.305 //y=0.905 //x2=26.305 //y2=1.25
r364 (  72 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=42.15 //y=6.02 //x2=42.15 //y2=4.865
r365 (  71 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.71 //y=6.02 //x2=41.71 //y2=4.865
r366 (  70 87 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.75 //y=6.02 //x2=26.75 //y2=4.865
r367 (  69 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.31 //y=6.02 //x2=26.31 //y2=4.865
r368 (  68 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=41.88 //y=1.365 //x2=41.99 //y2=1.365
r369 (  68 102 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=41.88 //y=1.365 //x2=41.77 //y2=1.365
r370 (  67 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=26.57 //y=1.405 //x2=26.68 //y2=1.405
r371 (  67 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=26.57 //y=1.405 //x2=26.46 //y2=1.405
r372 (  64 66 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=31.817 //y=4.07 //x2=31.817 //y2=4.235
r373 (  64 65 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=31.817 //y=4.07 //x2=31.817 //y2=3.905
r374 (  60 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.3 //y=4.7 //x2=26.3 //y2=4.7
r375 (  57 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.81 //y=4.7 //x2=41.81 //y2=4.7
r376 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=41.81 //y=4.07 //x2=41.81 //y2=4.7
r377 (  52 123 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.81 //y=2.08 //x2=41.81 //y2=2.08
r378 (  52 55 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=41.81 //y=2.08 //x2=41.81 //y2=4.07
r379 (  50 66 ) resistor r=57.1551 //w=0.187 //l=0.835 //layer=li \
 //thickness=0.1 //x=31.82 //y=5.07 //x2=31.82 //y2=4.235
r380 (  47 65 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=31.82 //y=1.75 //x2=31.82 //y2=3.905
r381 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=31.735 //y=1.665 //x2=31.82 //y2=1.75
r382 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=31.735 //y=1.665 //x2=31.42 //y2=1.665
r383 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=31.335 //y=1.58 //x2=31.42 //y2=1.665
r384 (  41 131 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=31.335 //y=1.58 //x2=31.335 //y2=1.01
r385 (  40 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.125 //y=5.155 //x2=31.04 //y2=5.155
r386 (  39 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=31.735 //y=5.155 //x2=31.82 //y2=5.07
r387 (  39 40 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=31.735 //y=5.155 //x2=31.125 //y2=5.155
r388 (  33 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.04 //y=5.24 //x2=31.04 //y2=5.155
r389 (  33 135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.04 //y=5.24 //x2=31.04 //y2=5.725
r390 (  32 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.245 //y=5.155 //x2=30.16 //y2=5.155
r391 (  31 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.955 //y=5.155 //x2=31.04 //y2=5.155
r392 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=30.955 //y=5.155 //x2=30.245 //y2=5.155
r393 (  25 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.16 //y=5.24 //x2=30.16 //y2=5.155
r394 (  25 134 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=30.16 //y=5.24 //x2=30.16 //y2=5.725
r395 (  23 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.075 //y=5.155 //x2=30.16 //y2=5.155
r396 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=30.075 //y=5.155 //x2=29.365 //y2=5.155
r397 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=29.28 //y=5.24 //x2=29.365 //y2=5.155
r398 (  17 133 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=29.28 //y=5.24 //x2=29.28 //y2=5.725
r399 (  13 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=2.08 //x2=26.27 //y2=2.08
r400 (  13 16 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.08 //x2=26.27 //y2=4.07
r401 (  11 60 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=26.27 //y=4.535 //x2=26.285 //y2=4.7
r402 (  11 16 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=26.27 //y=4.535 //x2=26.27 //y2=4.07
r403 (  10 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=41.81 //y=4.07 //x2=41.81 //y2=4.07
r404 (  8 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=31.815 //y=4.07 //x2=31.815 //y2=4.07
r405 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=26.27 //y=4.07 //x2=26.27 //y2=4.07
r406 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.93 //y=4.07 //x2=31.815 //y2=4.07
r407 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=41.695 //y=4.07 //x2=41.81 //y2=4.07
r408 (  3 4 ) resistor r=9.31775 //w=0.131 //l=9.765 //layer=m1 \
 //thickness=0.36 //x=41.695 //y=4.07 //x2=31.93 //y2=4.07
r409 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=26.385 //y=4.07 //x2=26.27 //y2=4.07
r410 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.7 //y=4.07 //x2=31.815 //y2=4.07
r411 (  1 2 ) resistor r=5.07156 //w=0.131 //l=5.315 //layer=m1 \
 //thickness=0.36 //x=31.7 //y=4.07 //x2=26.385 //y2=4.07
ends PM_TMRDFFSNQNX1\%noxref_10

subckt PM_TMRDFFSNQNX1\%noxref_11 ( 1 2 3 4 5 6 16 24 37 38 49 51 52 56 58 65 \
 66 67 68 69 70 71 72 73 74 78 79 80 85 87 90 91 95 96 97 102 104 107 108 112 \
 113 114 119 121 124 125 127 128 133 137 138 143 147 148 153 156 158 159 )
c322 ( 159 0 ) capacitor c=0.0220291f //x=39.335 //y=5.02
c323 ( 158 0 ) capacitor c=0.0217503f //x=38.455 //y=5.02
c324 ( 156 0 ) capacitor c=0.00866655f //x=39.33 //y=0.905
c325 ( 153 0 ) capacitor c=0.0587755f //x=47.36 //y=4.7
c326 ( 148 0 ) capacitor c=0.0273931f //x=47.36 //y=1.915
c327 ( 147 0 ) capacitor c=0.0456313f //x=47.36 //y=2.08
c328 ( 143 0 ) capacitor c=0.0587755f //x=35.89 //y=4.7
c329 ( 138 0 ) capacitor c=0.0273931f //x=35.89 //y=1.915
c330 ( 137 0 ) capacitor c=0.0456313f //x=35.89 //y=2.08
c331 ( 133 0 ) capacitor c=0.058931f //x=31.08 //y=4.7
c332 ( 128 0 ) capacitor c=0.0267105f //x=31.08 //y=1.915
c333 ( 127 0 ) capacitor c=0.0456313f //x=31.08 //y=2.08
c334 ( 125 0 ) capacitor c=0.0432517f //x=47.88 //y=1.26
c335 ( 124 0 ) capacitor c=0.0200379f //x=47.88 //y=0.915
c336 ( 121 0 ) capacitor c=0.0148873f //x=47.725 //y=1.415
c337 ( 119 0 ) capacitor c=0.0157803f //x=47.725 //y=0.76
c338 ( 114 0 ) capacitor c=0.0218028f //x=47.35 //y=1.57
c339 ( 113 0 ) capacitor c=0.0207459f //x=47.35 //y=1.26
c340 ( 112 0 ) capacitor c=0.0194308f //x=47.35 //y=0.915
c341 ( 108 0 ) capacitor c=0.0432517f //x=36.41 //y=1.26
c342 ( 107 0 ) capacitor c=0.0200379f //x=36.41 //y=0.915
c343 ( 104 0 ) capacitor c=0.0148873f //x=36.255 //y=1.415
c344 ( 102 0 ) capacitor c=0.0157803f //x=36.255 //y=0.76
c345 ( 97 0 ) capacitor c=0.0218028f //x=35.88 //y=1.57
c346 ( 96 0 ) capacitor c=0.0207459f //x=35.88 //y=1.26
c347 ( 95 0 ) capacitor c=0.0194308f //x=35.88 //y=0.915
c348 ( 91 0 ) capacitor c=0.0432517f //x=31.6 //y=1.26
c349 ( 90 0 ) capacitor c=0.0200379f //x=31.6 //y=0.915
c350 ( 87 0 ) capacitor c=0.0148873f //x=31.445 //y=1.415
c351 ( 85 0 ) capacitor c=0.0157803f //x=31.445 //y=0.76
c352 ( 80 0 ) capacitor c=0.0218028f //x=31.07 //y=1.57
c353 ( 79 0 ) capacitor c=0.0207459f //x=31.07 //y=1.26
c354 ( 78 0 ) capacitor c=0.0194308f //x=31.07 //y=0.915
c355 ( 74 0 ) capacitor c=0.158794f //x=47.54 //y=6.02
c356 ( 73 0 ) capacitor c=0.110114f //x=47.1 //y=6.02
c357 ( 72 0 ) capacitor c=0.158794f //x=36.07 //y=6.02
c358 ( 71 0 ) capacitor c=0.110114f //x=35.63 //y=6.02
c359 ( 70 0 ) capacitor c=0.158048f //x=31.26 //y=6.02
c360 ( 69 0 ) capacitor c=0.110114f //x=30.82 //y=6.02
c361 ( 65 0 ) capacitor c=0.00211606f //x=39.48 //y=5.2
c362 ( 58 0 ) capacitor c=0.0796302f //x=47.36 //y=2.08
c363 ( 56 0 ) capacitor c=0.103614f //x=39.96 //y=3.7
c364 ( 52 0 ) capacitor c=0.00404073f //x=39.605 //y=1.655
c365 ( 51 0 ) capacitor c=0.0122201f //x=39.875 //y=1.655
c366 ( 49 0 ) capacitor c=0.0137522f //x=39.875 //y=5.2
c367 ( 38 0 ) capacitor c=0.00251635f //x=38.685 //y=5.2
c368 ( 37 0 ) capacitor c=0.0142529f //x=39.395 //y=5.2
c369 ( 24 0 ) capacitor c=0.0811636f //x=35.89 //y=2.08
c370 ( 16 0 ) capacitor c=0.0796434f //x=31.08 //y=2.08
c371 ( 6 0 ) capacitor c=0.00405261f //x=40.075 //y=3.7
c372 ( 5 0 ) capacitor c=0.120326f //x=47.245 //y=3.7
c373 ( 4 0 ) capacitor c=0.00412452f //x=36.005 //y=3.7
c374 ( 3 0 ) capacitor c=0.0546427f //x=39.845 //y=3.7
c375 ( 2 0 ) capacitor c=0.0138772f //x=31.195 //y=3.7
c376 ( 1 0 ) capacitor c=0.0670382f //x=35.775 //y=3.7
r377 (  147 148 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=47.36 //y=2.08 //x2=47.36 //y2=1.915
r378 (  137 138 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=35.89 //y=2.08 //x2=35.89 //y2=1.915
r379 (  127 128 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=31.08 //y=2.08 //x2=31.08 //y2=1.915
r380 (  125 155 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.88 //y=1.26 //x2=47.84 //y2=1.415
r381 (  124 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.88 //y=0.915 //x2=47.84 //y2=0.76
r382 (  124 125 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=47.88 //y=0.915 //x2=47.88 //y2=1.26
r383 (  122 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.505 //y=1.415 //x2=47.39 //y2=1.415
r384 (  121 155 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.725 //y=1.415 //x2=47.84 //y2=1.415
r385 (  120 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.505 //y=0.76 //x2=47.39 //y2=0.76
r386 (  119 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.725 //y=0.76 //x2=47.84 //y2=0.76
r387 (  119 120 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=47.725 //y=0.76 //x2=47.505 //y2=0.76
r388 (  116 153 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=47.54 //y=4.865 //x2=47.36 //y2=4.7
r389 (  114 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.35 //y=1.57 //x2=47.39 //y2=1.415
r390 (  114 148 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=47.35 //y=1.57 //x2=47.35 //y2=1.915
r391 (  113 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.35 //y=1.26 //x2=47.39 //y2=1.415
r392 (  112 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.35 //y=0.915 //x2=47.39 //y2=0.76
r393 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=47.35 //y=0.915 //x2=47.35 //y2=1.26
r394 (  109 153 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=47.1 //y=4.865 //x2=47.36 //y2=4.7
r395 (  108 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.41 //y=1.26 //x2=36.37 //y2=1.415
r396 (  107 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.41 //y=0.915 //x2=36.37 //y2=0.76
r397 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=36.41 //y=0.915 //x2=36.41 //y2=1.26
r398 (  105 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.035 //y=1.415 //x2=35.92 //y2=1.415
r399 (  104 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.255 //y=1.415 //x2=36.37 //y2=1.415
r400 (  103 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.035 //y=0.76 //x2=35.92 //y2=0.76
r401 (  102 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.255 //y=0.76 //x2=36.37 //y2=0.76
r402 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=36.255 //y=0.76 //x2=36.035 //y2=0.76
r403 (  99 143 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=36.07 //y=4.865 //x2=35.89 //y2=4.7
r404 (  97 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.88 //y=1.57 //x2=35.92 //y2=1.415
r405 (  97 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=35.88 //y=1.57 //x2=35.88 //y2=1.915
r406 (  96 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.88 //y=1.26 //x2=35.92 //y2=1.415
r407 (  95 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.88 //y=0.915 //x2=35.92 //y2=0.76
r408 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=35.88 //y=0.915 //x2=35.88 //y2=1.26
r409 (  92 143 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=35.63 //y=4.865 //x2=35.89 //y2=4.7
r410 (  91 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.6 //y=1.26 //x2=31.56 //y2=1.415
r411 (  90 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.6 //y=0.915 //x2=31.56 //y2=0.76
r412 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.6 //y=0.915 //x2=31.6 //y2=1.26
r413 (  88 131 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.225 //y=1.415 //x2=31.11 //y2=1.415
r414 (  87 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.445 //y=1.415 //x2=31.56 //y2=1.415
r415 (  86 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.225 //y=0.76 //x2=31.11 //y2=0.76
r416 (  85 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.445 //y=0.76 //x2=31.56 //y2=0.76
r417 (  85 86 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=31.445 //y=0.76 //x2=31.225 //y2=0.76
r418 (  82 133 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=31.26 //y=4.865 //x2=31.08 //y2=4.7
r419 (  80 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.07 //y=1.57 //x2=31.11 //y2=1.415
r420 (  80 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.07 //y=1.57 //x2=31.07 //y2=1.915
r421 (  79 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.07 //y=1.26 //x2=31.11 //y2=1.415
r422 (  78 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.07 //y=0.915 //x2=31.11 //y2=0.76
r423 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.07 //y=0.915 //x2=31.07 //y2=1.26
r424 (  75 133 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=30.82 //y=4.865 //x2=31.08 //y2=4.7
r425 (  74 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=47.54 //y=6.02 //x2=47.54 //y2=4.865
r426 (  73 109 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=47.1 //y=6.02 //x2=47.1 //y2=4.865
r427 (  72 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=36.07 //y=6.02 //x2=36.07 //y2=4.865
r428 (  71 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.63 //y=6.02 //x2=35.63 //y2=4.865
r429 (  70 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.26 //y=6.02 //x2=31.26 //y2=4.865
r430 (  69 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.82 //y=6.02 //x2=30.82 //y2=4.865
r431 (  68 121 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=47.615 //y=1.415 //x2=47.725 //y2=1.415
r432 (  68 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=47.615 //y=1.415 //x2=47.505 //y2=1.415
r433 (  67 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=36.145 //y=1.415 //x2=36.255 //y2=1.415
r434 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=36.145 //y=1.415 //x2=36.035 //y2=1.415
r435 (  66 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=31.335 //y=1.415 //x2=31.445 //y2=1.415
r436 (  66 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=31.335 //y=1.415 //x2=31.225 //y2=1.415
r437 (  63 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=47.36 //y=4.7 //x2=47.36 //y2=4.7
r438 (  61 63 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=47.36 //y=3.7 //x2=47.36 //y2=4.7
r439 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=47.36 //y=2.08 //x2=47.36 //y2=2.08
r440 (  58 61 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=47.36 //y=2.08 //x2=47.36 //y2=3.7
r441 (  54 56 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=39.96 //y=5.115 //x2=39.96 //y2=3.7
r442 (  53 56 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=39.96 //y=1.74 //x2=39.96 //y2=3.7
r443 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=39.875 //y=1.655 //x2=39.96 //y2=1.74
r444 (  51 52 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=39.875 //y=1.655 //x2=39.605 //y2=1.655
r445 (  50 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.565 //y=5.2 //x2=39.48 //y2=5.2
r446 (  49 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=39.875 //y=5.2 //x2=39.96 //y2=5.115
r447 (  49 50 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=39.875 //y=5.2 //x2=39.565 //y2=5.2
r448 (  45 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=39.52 //y=1.57 //x2=39.605 //y2=1.655
r449 (  45 156 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=39.52 //y=1.57 //x2=39.52 //y2=1
r450 (  39 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.48 //y=5.285 //x2=39.48 //y2=5.2
r451 (  39 159 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=39.48 //y=5.285 //x2=39.48 //y2=5.725
r452 (  37 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.395 //y=5.2 //x2=39.48 //y2=5.2
r453 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=39.395 //y=5.2 //x2=38.685 //y2=5.2
r454 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=38.6 //y=5.285 //x2=38.685 //y2=5.2
r455 (  31 158 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=38.6 //y=5.285 //x2=38.6 //y2=5.725
r456 (  29 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.89 //y=4.7 //x2=35.89 //y2=4.7
r457 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=35.89 //y=3.7 //x2=35.89 //y2=4.7
r458 (  24 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.89 //y=2.08 //x2=35.89 //y2=2.08
r459 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=35.89 //y=2.08 //x2=35.89 //y2=3.7
r460 (  21 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.08 //y=4.7 //x2=31.08 //y2=4.7
r461 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=31.08 //y=3.7 //x2=31.08 //y2=4.7
r462 (  16 127 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.08 //y=2.08 //x2=31.08 //y2=2.08
r463 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=31.08 //y=2.08 //x2=31.08 //y2=3.7
r464 (  14 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=47.36 //y=3.7 //x2=47.36 //y2=3.7
r465 (  12 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=39.96 //y=3.7 //x2=39.96 //y2=3.7
r466 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=35.89 //y=3.7 //x2=35.89 //y2=3.7
r467 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=31.08 //y=3.7 //x2=31.08 //y2=3.7
r468 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=40.075 //y=3.7 //x2=39.96 //y2=3.7
r469 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.245 //y=3.7 //x2=47.36 //y2=3.7
r470 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=47.245 //y=3.7 //x2=40.075 //y2=3.7
r471 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=36.005 //y=3.7 //x2=35.89 //y2=3.7
r472 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=39.845 //y=3.7 //x2=39.96 //y2=3.7
r473 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=39.845 //y=3.7 //x2=36.005 //y2=3.7
r474 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.195 //y=3.7 //x2=31.08 //y2=3.7
r475 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=35.775 //y=3.7 //x2=35.89 //y2=3.7
r476 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=35.775 //y=3.7 //x2=31.195 //y2=3.7
ends PM_TMRDFFSNQNX1\%noxref_11

subckt PM_TMRDFFSNQNX1\%noxref_12 ( 1 2 7 9 19 20 27 35 41 42 46 49 50 51 52 \
 53 54 55 56 61 63 65 71 72 74 75 78 86 88 89 90 )
c181 ( 90 0 ) capacitor c=0.023087f //x=47.175 //y=5.02
c182 ( 89 0 ) capacitor c=0.023519f //x=46.295 //y=5.02
c183 ( 88 0 ) capacitor c=0.0224735f //x=45.415 //y=5.02
c184 ( 86 0 ) capacitor c=0.00872971f //x=47.425 //y=0.915
c185 ( 78 0 ) capacitor c=0.0331095f //x=42.58 //y=4.7
c186 ( 75 0 ) capacitor c=0.0279499f //x=42.55 //y=1.915
c187 ( 74 0 ) capacitor c=0.0421676f //x=42.55 //y=2.08
c188 ( 72 0 ) capacitor c=0.0429696f //x=43.115 //y=1.25
c189 ( 71 0 ) capacitor c=0.0192208f //x=43.115 //y=0.905
c190 ( 65 0 ) capacitor c=0.0148884f //x=42.96 //y=1.405
c191 ( 63 0 ) capacitor c=0.0157803f //x=42.96 //y=0.75
c192 ( 61 0 ) capacitor c=0.0295235f //x=42.955 //y=4.79
c193 ( 56 0 ) capacitor c=0.0205163f //x=42.585 //y=1.56
c194 ( 55 0 ) capacitor c=0.0168481f //x=42.585 //y=1.25
c195 ( 54 0 ) capacitor c=0.0174783f //x=42.585 //y=0.905
c196 ( 53 0 ) capacitor c=0.15358f //x=43.03 //y=6.02
c197 ( 52 0 ) capacitor c=0.110281f //x=42.59 //y=6.02
c198 ( 50 0 ) capacitor c=0.00106608f //x=47.32 //y=5.155
c199 ( 49 0 ) capacitor c=0.00207319f //x=46.44 //y=5.155
c200 ( 46 0 ) capacitor c=0.106168f //x=48.1 //y=4.07
c201 ( 42 0 ) capacitor c=0.00398962f //x=47.7 //y=1.665
c202 ( 41 0 ) capacitor c=0.0137288f //x=48.015 //y=1.665
c203 ( 35 0 ) capacitor c=0.0284988f //x=48.015 //y=5.155
c204 ( 27 0 ) capacitor c=0.0176454f //x=47.235 //y=5.155
c205 ( 20 0 ) capacitor c=0.00332903f //x=45.645 //y=5.155
c206 ( 19 0 ) capacitor c=0.0148427f //x=46.355 //y=5.155
c207 ( 9 0 ) capacitor c=0.0689632f //x=42.55 //y=2.08
c208 ( 7 0 ) capacitor c=0.00453889f //x=42.55 //y=4.535
c209 ( 2 0 ) capacitor c=0.00621861f //x=42.665 //y=4.07
c210 ( 1 0 ) capacitor c=0.0841928f //x=47.985 //y=4.07
r211 (  80 81 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=42.58 //y=4.79 //x2=42.58 //y2=4.865
r212 (  78 80 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=42.58 //y=4.7 //x2=42.58 //y2=4.79
r213 (  74 75 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=42.55 //y=2.08 //x2=42.55 //y2=1.915
r214 (  72 85 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=43.115 //y=1.25 //x2=43.075 //y2=1.405
r215 (  71 84 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=43.115 //y=0.905 //x2=43.075 //y2=0.75
r216 (  71 72 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=43.115 //y=0.905 //x2=43.115 //y2=1.25
r217 (  66 83 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.74 //y=1.405 //x2=42.625 //y2=1.405
r218 (  65 85 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.96 //y=1.405 //x2=43.075 //y2=1.405
r219 (  64 82 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.74 //y=0.75 //x2=42.625 //y2=0.75
r220 (  63 84 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.96 //y=0.75 //x2=43.075 //y2=0.75
r221 (  63 64 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=42.96 //y=0.75 //x2=42.74 //y2=0.75
r222 (  62 80 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=42.715 //y=4.79 //x2=42.58 //y2=4.79
r223 (  61 68 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=42.955 //y=4.79 //x2=43.03 //y2=4.865
r224 (  61 62 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=42.955 //y=4.79 //x2=42.715 //y2=4.79
r225 (  56 83 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.585 //y=1.56 //x2=42.625 //y2=1.405
r226 (  56 75 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=42.585 //y=1.56 //x2=42.585 //y2=1.915
r227 (  55 83 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.585 //y=1.25 //x2=42.625 //y2=1.405
r228 (  54 82 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.585 //y=0.905 //x2=42.625 //y2=0.75
r229 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.585 //y=0.905 //x2=42.585 //y2=1.25
r230 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=43.03 //y=6.02 //x2=43.03 //y2=4.865
r231 (  52 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=42.59 //y=6.02 //x2=42.59 //y2=4.865
r232 (  51 65 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.85 //y=1.405 //x2=42.96 //y2=1.405
r233 (  51 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.85 //y=1.405 //x2=42.74 //y2=1.405
r234 (  48 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=42.58 //y=4.7 //x2=42.58 //y2=4.7
r235 (  44 46 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=48.1 //y=5.07 //x2=48.1 //y2=4.07
r236 (  43 46 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=48.1 //y=1.75 //x2=48.1 //y2=4.07
r237 (  41 43 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=48.015 //y=1.665 //x2=48.1 //y2=1.75
r238 (  41 42 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=48.015 //y=1.665 //x2=47.7 //y2=1.665
r239 (  37 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=47.615 //y=1.58 //x2=47.7 //y2=1.665
r240 (  37 86 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=47.615 //y=1.58 //x2=47.615 //y2=1.01
r241 (  36 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.405 //y=5.155 //x2=47.32 //y2=5.155
r242 (  35 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=48.015 //y=5.155 //x2=48.1 //y2=5.07
r243 (  35 36 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=48.015 //y=5.155 //x2=47.405 //y2=5.155
r244 (  29 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.32 //y=5.24 //x2=47.32 //y2=5.155
r245 (  29 90 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=47.32 //y=5.24 //x2=47.32 //y2=5.725
r246 (  28 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.525 //y=5.155 //x2=46.44 //y2=5.155
r247 (  27 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.235 //y=5.155 //x2=47.32 //y2=5.155
r248 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=47.235 //y=5.155 //x2=46.525 //y2=5.155
r249 (  21 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.44 //y=5.24 //x2=46.44 //y2=5.155
r250 (  21 89 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.44 //y=5.24 //x2=46.44 //y2=5.725
r251 (  19 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.355 //y=5.155 //x2=46.44 //y2=5.155
r252 (  19 20 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.355 //y=5.155 //x2=45.645 //y2=5.155
r253 (  13 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=45.56 //y=5.24 //x2=45.645 //y2=5.155
r254 (  13 88 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.56 //y=5.24 //x2=45.56 //y2=5.725
r255 (  9 74 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=42.55 //y=2.08 //x2=42.55 //y2=2.08
r256 (  9 12 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=42.55 //y=2.08 //x2=42.55 //y2=4.07
r257 (  7 48 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=42.55 //y=4.535 //x2=42.565 //y2=4.7
r258 (  7 12 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=42.55 //y=4.535 //x2=42.55 //y2=4.07
r259 (  6 46 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=48.1 //y=4.07 //x2=48.1 //y2=4.07
r260 (  4 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=42.55 //y=4.07 //x2=42.55 //y2=4.07
r261 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=42.665 //y=4.07 //x2=42.55 //y2=4.07
r262 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.985 //y=4.07 //x2=48.1 //y2=4.07
r263 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=47.985 //y=4.07 //x2=42.665 //y2=4.07
ends PM_TMRDFFSNQNX1\%noxref_12

subckt PM_TMRDFFSNQNX1\%D ( 1 2 3 4 11 12 13 14 15 16 17 18 19 20 21 22 23 25 \
 38 49 58 59 60 61 62 63 64 65 66 67 68 69 70 74 76 79 80 84 85 86 87 91 93 96 \
 97 101 102 103 104 108 110 113 114 124 133 142 )
c323 ( 142 0 ) capacitor c=0.0588816f //x=49.95 //y=4.7
c324 ( 133 0 ) capacitor c=0.0588816f //x=25.53 //y=4.7
c325 ( 124 0 ) capacitor c=0.0667949f //x=1.11 //y=4.7
c326 ( 114 0 ) capacitor c=0.0318948f //x=50.285 //y=1.21
c327 ( 113 0 ) capacitor c=0.0187384f //x=50.285 //y=0.865
c328 ( 110 0 ) capacitor c=0.0141798f //x=50.13 //y=1.365
c329 ( 108 0 ) capacitor c=0.0149844f //x=50.13 //y=0.71
c330 ( 104 0 ) capacitor c=0.0813322f //x=49.755 //y=1.915
c331 ( 103 0 ) capacitor c=0.0229267f //x=49.755 //y=1.52
c332 ( 102 0 ) capacitor c=0.0234352f //x=49.755 //y=1.21
c333 ( 101 0 ) capacitor c=0.0199343f //x=49.755 //y=0.865
c334 ( 97 0 ) capacitor c=0.0318948f //x=25.865 //y=1.21
c335 ( 96 0 ) capacitor c=0.0187384f //x=25.865 //y=0.865
c336 ( 93 0 ) capacitor c=0.0141798f //x=25.71 //y=1.365
c337 ( 91 0 ) capacitor c=0.0149844f //x=25.71 //y=0.71
c338 ( 87 0 ) capacitor c=0.0813322f //x=25.335 //y=1.915
c339 ( 86 0 ) capacitor c=0.0229267f //x=25.335 //y=1.52
c340 ( 85 0 ) capacitor c=0.0234352f //x=25.335 //y=1.21
c341 ( 84 0 ) capacitor c=0.0199343f //x=25.335 //y=0.865
c342 ( 80 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c343 ( 79 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c344 ( 76 0 ) capacitor c=0.0141798f //x=1.29 //y=1.365
c345 ( 74 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c346 ( 70 0 ) capacitor c=0.0844059f //x=0.915 //y=1.915
c347 ( 69 0 ) capacitor c=0.0229722f //x=0.915 //y=1.52
c348 ( 68 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c349 ( 67 0 ) capacitor c=0.0199343f //x=0.915 //y=0.865
c350 ( 66 0 ) capacitor c=0.110275f //x=50.29 //y=6.02
c351 ( 65 0 ) capacitor c=0.154305f //x=49.85 //y=6.02
c352 ( 64 0 ) capacitor c=0.110275f //x=25.87 //y=6.02
c353 ( 63 0 ) capacitor c=0.154305f //x=25.43 //y=6.02
c354 ( 62 0 ) capacitor c=0.110275f //x=1.45 //y=6.02
c355 ( 61 0 ) capacitor c=0.154305f //x=1.01 //y=6.02
c356 ( 49 0 ) capacitor c=0.0877439f //x=49.95 //y=2.08
c357 ( 38 0 ) capacitor c=0.0899325f //x=25.53 //y=2.08
c358 ( 25 0 ) capacitor c=0.111725f //x=1.11 //y=2.08
c359 ( 4 0 ) capacitor c=0.00583987f //x=25.645 //y=2.96
c360 ( 3 0 ) capacitor c=0.366619f //x=49.835 //y=2.96
c361 ( 2 0 ) capacitor c=0.0150814f //x=1.225 //y=2.96
c362 ( 1 0 ) capacitor c=0.47261f //x=25.415 //y=2.96
r363 (  140 142 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=49.85 //y=4.7 //x2=49.95 //y2=4.7
r364 (  131 133 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=25.43 //y=4.7 //x2=25.53 //y2=4.7
r365 (  122 124 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.7 //x2=1.11 //y2=4.7
r366 (  115 142 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=50.29 //y=4.865 //x2=49.95 //y2=4.7
r367 (  114 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.285 //y=1.21 //x2=50.245 //y2=1.365
r368 (  113 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.285 //y=0.865 //x2=50.245 //y2=0.71
r369 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=50.285 //y=0.865 //x2=50.285 //y2=1.21
r370 (  111 139 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.91 //y=1.365 //x2=49.795 //y2=1.365
r371 (  110 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.13 //y=1.365 //x2=50.245 //y2=1.365
r372 (  109 138 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.91 //y=0.71 //x2=49.795 //y2=0.71
r373 (  108 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.13 //y=0.71 //x2=50.245 //y2=0.71
r374 (  108 109 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=50.13 //y=0.71 //x2=49.91 //y2=0.71
r375 (  105 140 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=49.85 //y=4.865 //x2=49.85 //y2=4.7
r376 (  104 137 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=49.755 //y=1.915 //x2=49.95 //y2=2.08
r377 (  103 139 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.755 //y=1.52 //x2=49.795 //y2=1.365
r378 (  103 104 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=49.755 //y=1.52 //x2=49.755 //y2=1.915
r379 (  102 139 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.755 //y=1.21 //x2=49.795 //y2=1.365
r380 (  101 138 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.755 //y=0.865 //x2=49.795 //y2=0.71
r381 (  101 102 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=49.755 //y=0.865 //x2=49.755 //y2=1.21
r382 (  98 133 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=25.87 //y=4.865 //x2=25.53 //y2=4.7
r383 (  97 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.865 //y=1.21 //x2=25.825 //y2=1.365
r384 (  96 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.865 //y=0.865 //x2=25.825 //y2=0.71
r385 (  96 97 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=25.865 //y=0.865 //x2=25.865 //y2=1.21
r386 (  94 130 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.49 //y=1.365 //x2=25.375 //y2=1.365
r387 (  93 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.71 //y=1.365 //x2=25.825 //y2=1.365
r388 (  92 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.49 //y=0.71 //x2=25.375 //y2=0.71
r389 (  91 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.71 //y=0.71 //x2=25.825 //y2=0.71
r390 (  91 92 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=25.71 //y=0.71 //x2=25.49 //y2=0.71
r391 (  88 131 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=25.43 //y=4.865 //x2=25.43 //y2=4.7
r392 (  87 128 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=25.335 //y=1.915 //x2=25.53 //y2=2.08
r393 (  86 130 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.335 //y=1.52 //x2=25.375 //y2=1.365
r394 (  86 87 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=25.335 //y=1.52 //x2=25.335 //y2=1.915
r395 (  85 130 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.335 //y=1.21 //x2=25.375 //y2=1.365
r396 (  84 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.335 //y=0.865 //x2=25.375 //y2=0.71
r397 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=25.335 //y=0.865 //x2=25.335 //y2=1.21
r398 (  81 124 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=1.45 //y=4.865 //x2=1.11 //y2=4.7
r399 (  80 126 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r400 (  79 125 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r401 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r402 (  77 121 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r403 (  76 126 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r404 (  75 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r405 (  74 125 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r406 (  74 75 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r407 (  71 122 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.865 //x2=1.01 //y2=4.7
r408 (  70 119 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r409 (  69 121 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r410 (  69 70 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r411 (  68 121 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r412 (  67 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r413 (  67 68 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r414 (  66 115 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.29 //y=6.02 //x2=50.29 //y2=4.865
r415 (  65 105 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.85 //y=6.02 //x2=49.85 //y2=4.865
r416 (  64 98 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.87 //y=6.02 //x2=25.87 //y2=4.865
r417 (  63 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.43 //y=6.02 //x2=25.43 //y2=4.865
r418 (  62 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.02 //x2=1.45 //y2=4.865
r419 (  61 71 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.02 //x2=1.01 //y2=4.865
r420 (  60 110 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.02 //y=1.365 //x2=50.13 //y2=1.365
r421 (  60 111 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.02 //y=1.365 //x2=49.91 //y2=1.365
r422 (  59 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.6 //y=1.365 //x2=25.71 //y2=1.365
r423 (  59 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.6 //y=1.365 //x2=25.49 //y2=1.365
r424 (  58 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r425 (  58 77 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r426 (  56 142 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.95 //y=4.7 //x2=49.95 //y2=4.7
r427 (  49 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.95 //y=2.08 //x2=49.95 //y2=2.08
r428 (  46 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.53 //y=4.7 //x2=25.53 //y2=4.7
r429 (  38 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.53 //y=2.08 //x2=25.53 //y2=2.08
r430 (  35 124 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r431 (  25 119 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r432 (  23 56 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=49.95 //y=4.07 //x2=49.95 //y2=4.7
r433 (  22 23 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=49.95 //y=3.7 //x2=49.95 //y2=4.07
r434 (  21 22 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=49.95 //y=2.96 //x2=49.95 //y2=3.7
r435 (  21 49 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=49.95 //y=2.96 //x2=49.95 //y2=2.08
r436 (  20 46 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=25.53 //y=4.07 //x2=25.53 //y2=4.7
r437 (  19 20 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.53 //y=3.7 //x2=25.53 //y2=4.07
r438 (  18 19 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=25.53 //y=2.96 //x2=25.53 //y2=3.7
r439 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.53 //y=2.59 //x2=25.53 //y2=2.96
r440 (  17 38 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=25.53 //y=2.59 //x2=25.53 //y2=2.08
r441 (  16 35 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.44 //x2=1.11 //y2=4.7
r442 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r443 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r444 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r445 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r446 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r447 (  11 25 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.59 //x2=1.11 //y2=2.08
r448 (  10 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=49.95 //y=2.96 //x2=49.95 //y2=2.96
r449 (  8 18 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.53 //y=2.96 //x2=25.53 //y2=2.96
r450 (  6 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=2.96 //x2=1.11 //y2=2.96
r451 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.645 //y=2.96 //x2=25.53 //y2=2.96
r452 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=49.835 //y=2.96 //x2=49.95 //y2=2.96
r453 (  3 4 ) resistor r=23.0821 //w=0.131 //l=24.19 //layer=m1 \
 //thickness=0.36 //x=49.835 //y=2.96 //x2=25.645 //y2=2.96
r454 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=2.96 //x2=1.11 //y2=2.96
r455 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.415 //y=2.96 //x2=25.53 //y2=2.96
r456 (  1 2 ) resistor r=23.0821 //w=0.131 //l=24.19 //layer=m1 \
 //thickness=0.36 //x=25.415 //y=2.96 //x2=1.225 //y2=2.96
ends PM_TMRDFFSNQNX1\%D

subckt PM_TMRDFFSNQNX1\%noxref_14 ( 1 2 3 4 17 18 29 31 32 36 38 46 53 54 55 \
 56 57 58 59 60 61 62 63 64 66 72 73 74 75 79 80 81 82 83 85 91 92 93 94 114 \
 116 117 )
c236 ( 117 0 ) capacitor c=0.0220291f //x=50.805 //y=5.02
c237 ( 116 0 ) capacitor c=0.0217503f //x=49.925 //y=5.02
c238 ( 114 0 ) capacitor c=0.0084702f //x=50.8 //y=0.905
c239 ( 94 0 ) capacitor c=0.0556143f //x=58.365 //y=4.79
c240 ( 93 0 ) capacitor c=0.0293157f //x=58.655 //y=4.79
c241 ( 92 0 ) capacitor c=0.0347816f //x=58.32 //y=1.22
c242 ( 91 0 ) capacitor c=0.0187487f //x=58.32 //y=0.875
c243 ( 85 0 ) capacitor c=0.0137055f //x=58.165 //y=1.375
c244 ( 83 0 ) capacitor c=0.0149861f //x=58.165 //y=0.72
c245 ( 82 0 ) capacitor c=0.096037f //x=57.79 //y=1.915
c246 ( 81 0 ) capacitor c=0.0228993f //x=57.79 //y=1.53
c247 ( 80 0 ) capacitor c=0.0234352f //x=57.79 //y=1.22
c248 ( 79 0 ) capacitor c=0.0198724f //x=57.79 //y=0.875
c249 ( 75 0 ) capacitor c=0.0557698f //x=53.555 //y=4.79
c250 ( 74 0 ) capacitor c=0.0293157f //x=53.845 //y=4.79
c251 ( 73 0 ) capacitor c=0.0347816f //x=53.51 //y=1.22
c252 ( 72 0 ) capacitor c=0.0187487f //x=53.51 //y=0.875
c253 ( 66 0 ) capacitor c=0.0137055f //x=53.355 //y=1.375
c254 ( 64 0 ) capacitor c=0.0149861f //x=53.355 //y=0.72
c255 ( 63 0 ) capacitor c=0.096037f //x=52.98 //y=1.915
c256 ( 62 0 ) capacitor c=0.0228993f //x=52.98 //y=1.53
c257 ( 61 0 ) capacitor c=0.0234352f //x=52.98 //y=1.22
c258 ( 60 0 ) capacitor c=0.0198724f //x=52.98 //y=0.875
c259 ( 59 0 ) capacitor c=0.110114f //x=58.73 //y=6.02
c260 ( 58 0 ) capacitor c=0.158956f //x=58.29 //y=6.02
c261 ( 57 0 ) capacitor c=0.110114f //x=53.92 //y=6.02
c262 ( 56 0 ) capacitor c=0.158956f //x=53.48 //y=6.02
c263 ( 53 0 ) capacitor c=0.00211606f //x=50.95 //y=5.2
c264 ( 46 0 ) capacitor c=0.0943831f //x=58.09 //y=2.08
c265 ( 38 0 ) capacitor c=0.0969368f //x=53.28 //y=2.08
c266 ( 36 0 ) capacitor c=0.104691f //x=51.43 //y=2.59
c267 ( 32 0 ) capacitor c=0.00404073f //x=51.075 //y=1.655
c268 ( 31 0 ) capacitor c=0.0122201f //x=51.345 //y=1.655
c269 ( 29 0 ) capacitor c=0.0137995f //x=51.345 //y=5.2
c270 ( 18 0 ) capacitor c=0.00251635f //x=50.155 //y=5.2
c271 ( 17 0 ) capacitor c=0.0143649f //x=50.865 //y=5.2
c272 ( 4 0 ) capacitor c=0.00673266f //x=53.545 //y=2.59
c273 ( 3 0 ) capacitor c=0.0686809f //x=57.975 //y=2.59
c274 ( 2 0 ) capacitor c=0.00544459f //x=51.545 //y=2.59
c275 ( 1 0 ) capacitor c=0.0230071f //x=53.135 //y=2.59
r276 (  93 95 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=58.655 //y=4.79 //x2=58.73 //y2=4.865
r277 (  93 94 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=58.655 //y=4.79 //x2=58.365 //y2=4.79
r278 (  92 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.32 //y=1.22 //x2=58.28 //y2=1.375
r279 (  91 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.32 //y=0.875 //x2=58.28 //y2=0.72
r280 (  91 92 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=58.32 //y=0.875 //x2=58.32 //y2=1.22
r281 (  88 94 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=58.29 //y=4.865 //x2=58.365 //y2=4.79
r282 (  88 111 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=58.29 //y=4.865 //x2=58.09 //y2=4.7
r283 (  86 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=57.945 //y=1.375 //x2=57.83 //y2=1.375
r284 (  85 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.165 //y=1.375 //x2=58.28 //y2=1.375
r285 (  84 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=57.945 //y=0.72 //x2=57.83 //y2=0.72
r286 (  83 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.165 //y=0.72 //x2=58.28 //y2=0.72
r287 (  83 84 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=58.165 //y=0.72 //x2=57.945 //y2=0.72
r288 (  82 109 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=57.79 //y=1.915 //x2=58.09 //y2=2.08
r289 (  81 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.79 //y=1.53 //x2=57.83 //y2=1.375
r290 (  81 82 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=57.79 //y=1.53 //x2=57.79 //y2=1.915
r291 (  80 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.79 //y=1.22 //x2=57.83 //y2=1.375
r292 (  79 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.79 //y=0.875 //x2=57.83 //y2=0.72
r293 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=57.79 //y=0.875 //x2=57.79 //y2=1.22
r294 (  74 76 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=53.845 //y=4.79 //x2=53.92 //y2=4.865
r295 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=53.845 //y=4.79 //x2=53.555 //y2=4.79
r296 (  73 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.51 //y=1.22 //x2=53.47 //y2=1.375
r297 (  72 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.51 //y=0.875 //x2=53.47 //y2=0.72
r298 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=53.51 //y=0.875 //x2=53.51 //y2=1.22
r299 (  69 75 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=53.48 //y=4.865 //x2=53.555 //y2=4.79
r300 (  69 103 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=53.48 //y=4.865 //x2=53.28 //y2=4.7
r301 (  67 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.135 //y=1.375 //x2=53.02 //y2=1.375
r302 (  66 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.355 //y=1.375 //x2=53.47 //y2=1.375
r303 (  65 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.135 //y=0.72 //x2=53.02 //y2=0.72
r304 (  64 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.355 //y=0.72 //x2=53.47 //y2=0.72
r305 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=53.355 //y=0.72 //x2=53.135 //y2=0.72
r306 (  63 101 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=52.98 //y=1.915 //x2=53.28 //y2=2.08
r307 (  62 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.98 //y=1.53 //x2=53.02 //y2=1.375
r308 (  62 63 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=52.98 //y=1.53 //x2=52.98 //y2=1.915
r309 (  61 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.98 //y=1.22 //x2=53.02 //y2=1.375
r310 (  60 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.98 //y=0.875 //x2=53.02 //y2=0.72
r311 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=52.98 //y=0.875 //x2=52.98 //y2=1.22
r312 (  59 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=58.73 //y=6.02 //x2=58.73 //y2=4.865
r313 (  58 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=58.29 //y=6.02 //x2=58.29 //y2=4.865
r314 (  57 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=53.92 //y=6.02 //x2=53.92 //y2=4.865
r315 (  56 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=53.48 //y=6.02 //x2=53.48 //y2=4.865
r316 (  55 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.055 //y=1.375 //x2=58.165 //y2=1.375
r317 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.055 //y=1.375 //x2=57.945 //y2=1.375
r318 (  54 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.245 //y=1.375 //x2=53.355 //y2=1.375
r319 (  54 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.245 //y=1.375 //x2=53.135 //y2=1.375
r320 (  51 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.09 //y=4.7 //x2=58.09 //y2=4.7
r321 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=58.09 //y=2.59 //x2=58.09 //y2=4.7
r322 (  46 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.09 //y=2.08 //x2=58.09 //y2=2.08
r323 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=58.09 //y=2.08 //x2=58.09 //y2=2.59
r324 (  43 103 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=53.28 //y=4.7 //x2=53.28 //y2=4.7
r325 (  41 43 ) resistor r=144.77 //w=0.187 //l=2.115 //layer=li \
 //thickness=0.1 //x=53.28 //y=2.585 //x2=53.28 //y2=4.7
r326 (  38 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=53.28 //y=2.08 //x2=53.28 //y2=2.08
r327 (  38 41 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=53.28 //y=2.08 //x2=53.28 //y2=2.585
r328 (  34 36 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=51.43 //y=5.115 //x2=51.43 //y2=2.59
r329 (  33 36 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=51.43 //y=1.74 //x2=51.43 //y2=2.59
r330 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=51.345 //y=1.655 //x2=51.43 //y2=1.74
r331 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=51.345 //y=1.655 //x2=51.075 //y2=1.655
r332 (  30 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.035 //y=5.2 //x2=50.95 //y2=5.2
r333 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=51.345 //y=5.2 //x2=51.43 //y2=5.115
r334 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=51.345 //y=5.2 //x2=51.035 //y2=5.2
r335 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=50.99 //y=1.57 //x2=51.075 //y2=1.655
r336 (  25 114 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=50.99 //y=1.57 //x2=50.99 //y2=1
r337 (  19 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.95 //y=5.285 //x2=50.95 //y2=5.2
r338 (  19 117 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=50.95 //y=5.285 //x2=50.95 //y2=5.725
r339 (  17 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.865 //y=5.2 //x2=50.95 //y2=5.2
r340 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.865 //y=5.2 //x2=50.155 //y2=5.2
r341 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=50.07 //y=5.285 //x2=50.155 //y2=5.2
r342 (  11 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=50.07 //y=5.285 //x2=50.07 //y2=5.725
r343 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=58.09 //y=2.59 //x2=58.09 //y2=2.59
r344 (  8 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=53.28 //y=2.585 //x2=53.28 //y2=2.585
r345 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=51.43 //y=2.59 //x2=51.43 //y2=2.59
r346 (  4 8 ) resistor r=0.164988 //w=0.206 //l=0.267488 //layer=m1 \
 //thickness=0.36 //x=53.545 //y=2.59 //x2=53.28 //y2=2.585
r347 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=57.975 //y=2.59 //x2=58.09 //y2=2.59
r348 (  3 4 ) resistor r=4.2271 //w=0.131 //l=4.43 //layer=m1 //thickness=0.36 \
 //x=57.975 //y=2.59 //x2=53.545 //y2=2.59
r349 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=51.545 //y=2.59 //x2=51.43 //y2=2.59
r350 (  1 8 ) resistor r=0.0921728 //w=0.206 //l=0.147479 //layer=m1 \
 //thickness=0.36 //x=53.135 //y=2.59 //x2=53.28 //y2=2.585
r351 (  1 2 ) resistor r=1.51718 //w=0.131 //l=1.59 //layer=m1 \
 //thickness=0.36 //x=53.135 //y=2.59 //x2=51.545 //y2=2.59
ends PM_TMRDFFSNQNX1\%noxref_14

subckt PM_TMRDFFSNQNX1\%noxref_15 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 61 63 66 67 77 80 82 83 84 )
c164 ( 84 0 ) capacitor c=0.023087f //x=60.125 //y=5.02
c165 ( 83 0 ) capacitor c=0.023519f //x=59.245 //y=5.02
c166 ( 82 0 ) capacitor c=0.0224735f //x=58.365 //y=5.02
c167 ( 80 0 ) capacitor c=0.00872971f //x=60.375 //y=0.915
c168 ( 77 0 ) capacitor c=0.0588816f //x=62.9 //y=4.7
c169 ( 67 0 ) capacitor c=0.0318948f //x=63.235 //y=1.21
c170 ( 66 0 ) capacitor c=0.0187384f //x=63.235 //y=0.865
c171 ( 63 0 ) capacitor c=0.0141798f //x=63.08 //y=1.365
c172 ( 61 0 ) capacitor c=0.0149844f //x=63.08 //y=0.71
c173 ( 57 0 ) capacitor c=0.0813322f //x=62.705 //y=1.915
c174 ( 56 0 ) capacitor c=0.0229267f //x=62.705 //y=1.52
c175 ( 55 0 ) capacitor c=0.0234352f //x=62.705 //y=1.21
c176 ( 54 0 ) capacitor c=0.0199343f //x=62.705 //y=0.865
c177 ( 53 0 ) capacitor c=0.110275f //x=63.24 //y=6.02
c178 ( 52 0 ) capacitor c=0.154305f //x=62.8 //y=6.02
c179 ( 50 0 ) capacitor c=0.00106608f //x=60.27 //y=5.155
c180 ( 49 0 ) capacitor c=0.00207319f //x=59.39 //y=5.155
c181 ( 42 0 ) capacitor c=0.0839295f //x=62.9 //y=2.08
c182 ( 40 0 ) capacitor c=0.10402f //x=61.05 //y=2.59
c183 ( 36 0 ) capacitor c=0.00398962f //x=60.65 //y=1.665
c184 ( 35 0 ) capacitor c=0.0137288f //x=60.965 //y=1.665
c185 ( 29 0 ) capacitor c=0.0284988f //x=60.965 //y=5.155
c186 ( 21 0 ) capacitor c=0.0176454f //x=60.185 //y=5.155
c187 ( 14 0 ) capacitor c=0.00332903f //x=58.595 //y=5.155
c188 ( 13 0 ) capacitor c=0.0148427f //x=59.305 //y=5.155
c189 ( 2 0 ) capacitor c=0.00808366f //x=61.165 //y=2.59
c190 ( 1 0 ) capacitor c=0.0353429f //x=62.785 //y=2.59
r191 (  75 77 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=62.8 //y=4.7 //x2=62.9 //y2=4.7
r192 (  68 77 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=63.24 //y=4.865 //x2=62.9 //y2=4.7
r193 (  67 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.235 //y=1.21 //x2=63.195 //y2=1.365
r194 (  66 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.235 //y=0.865 //x2=63.195 //y2=0.71
r195 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.235 //y=0.865 //x2=63.235 //y2=1.21
r196 (  64 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.86 //y=1.365 //x2=62.745 //y2=1.365
r197 (  63 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.08 //y=1.365 //x2=63.195 //y2=1.365
r198 (  62 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.86 //y=0.71 //x2=62.745 //y2=0.71
r199 (  61 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.08 //y=0.71 //x2=63.195 //y2=0.71
r200 (  61 62 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=63.08 //y=0.71 //x2=62.86 //y2=0.71
r201 (  58 75 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=62.8 //y=4.865 //x2=62.8 //y2=4.7
r202 (  57 72 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=62.705 //y=1.915 //x2=62.9 //y2=2.08
r203 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.705 //y=1.52 //x2=62.745 //y2=1.365
r204 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=62.705 //y=1.52 //x2=62.705 //y2=1.915
r205 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.705 //y=1.21 //x2=62.745 //y2=1.365
r206 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.705 //y=0.865 //x2=62.745 //y2=0.71
r207 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=62.705 //y=0.865 //x2=62.705 //y2=1.21
r208 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=63.24 //y=6.02 //x2=63.24 //y2=4.865
r209 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=62.8 //y=6.02 //x2=62.8 //y2=4.865
r210 (  51 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=62.97 //y=1.365 //x2=63.08 //y2=1.365
r211 (  51 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=62.97 //y=1.365 //x2=62.86 //y2=1.365
r212 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.9 //y=4.7 //x2=62.9 //y2=4.7
r213 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=62.9 //y=2.59 //x2=62.9 //y2=4.7
r214 (  42 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.9 //y=2.08 //x2=62.9 //y2=2.08
r215 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=62.9 //y=2.08 //x2=62.9 //y2=2.59
r216 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=61.05 //y=5.07 //x2=61.05 //y2=2.59
r217 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=61.05 //y=1.75 //x2=61.05 //y2=2.59
r218 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.965 //y=1.665 //x2=61.05 //y2=1.75
r219 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=60.965 //y=1.665 //x2=60.65 //y2=1.665
r220 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.565 //y=1.58 //x2=60.65 //y2=1.665
r221 (  31 80 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=60.565 //y=1.58 //x2=60.565 //y2=1.01
r222 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.355 //y=5.155 //x2=60.27 //y2=5.155
r223 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.965 //y=5.155 //x2=61.05 //y2=5.07
r224 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=60.965 //y=5.155 //x2=60.355 //y2=5.155
r225 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.27 //y=5.24 //x2=60.27 //y2=5.155
r226 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.27 //y=5.24 //x2=60.27 //y2=5.725
r227 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.475 //y=5.155 //x2=59.39 //y2=5.155
r228 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.185 //y=5.155 //x2=60.27 //y2=5.155
r229 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=60.185 //y=5.155 //x2=59.475 //y2=5.155
r230 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.39 //y=5.24 //x2=59.39 //y2=5.155
r231 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.39 //y=5.24 //x2=59.39 //y2=5.725
r232 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.305 //y=5.155 //x2=59.39 //y2=5.155
r233 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=59.305 //y=5.155 //x2=58.595 //y2=5.155
r234 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=58.51 //y=5.24 //x2=58.595 //y2=5.155
r235 (  7 82 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=58.51 //y=5.24 //x2=58.51 //y2=5.725
r236 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=62.9 //y=2.59 //x2=62.9 //y2=2.59
r237 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=61.05 //y=2.59 //x2=61.05 //y2=2.59
r238 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=61.165 //y=2.59 //x2=61.05 //y2=2.59
r239 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=62.785 //y=2.59 //x2=62.9 //y2=2.59
r240 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=62.785 //y=2.59 //x2=61.165 //y2=2.59
ends PM_TMRDFFSNQNX1\%noxref_15

subckt PM_TMRDFFSNQNX1\%CLK ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 31 \
 32 33 34 35 36 37 39 49 51 58 66 68 74 82 84 95 96 97 98 99 100 101 102 103 \
 104 105 106 107 108 109 110 111 112 113 114 115 117 123 124 125 126 127 132 \
 133 134 139 141 143 149 150 151 152 153 155 161 162 163 164 165 170 171 172 \
 177 179 181 187 188 189 190 191 193 199 200 201 202 203 208 209 210 215 217 \
 219 225 226 230 239 240 243 254 263 264 267 278 287 288 291 )
c752 ( 291 0 ) capacitor c=0.0331838f //x=63.67 //y=4.7
c753 ( 288 0 ) capacitor c=0.0279499f //x=63.64 //y=1.915
c754 ( 287 0 ) capacitor c=0.0421676f //x=63.64 //y=2.08
c755 ( 278 0 ) capacitor c=0.0334842f //x=54.39 //y=4.7
c756 ( 267 0 ) capacitor c=0.0331706f //x=39.25 //y=4.7
c757 ( 264 0 ) capacitor c=0.0279499f //x=39.22 //y=1.915
c758 ( 263 0 ) capacitor c=0.0421676f //x=39.22 //y=2.08
c759 ( 254 0 ) capacitor c=0.0334842f //x=29.97 //y=4.7
c760 ( 243 0 ) capacitor c=0.0331706f //x=14.83 //y=4.7
c761 ( 240 0 ) capacitor c=0.0279499f //x=14.8 //y=1.915
c762 ( 239 0 ) capacitor c=0.0421676f //x=14.8 //y=2.08
c763 ( 230 0 ) capacitor c=0.0334842f //x=5.55 //y=4.7
c764 ( 226 0 ) capacitor c=0.0429696f //x=64.205 //y=1.25
c765 ( 225 0 ) capacitor c=0.0192208f //x=64.205 //y=0.905
c766 ( 219 0 ) capacitor c=0.0148884f //x=64.05 //y=1.405
c767 ( 217 0 ) capacitor c=0.0157803f //x=64.05 //y=0.75
c768 ( 215 0 ) capacitor c=0.0299681f //x=64.045 //y=4.79
c769 ( 210 0 ) capacitor c=0.0205163f //x=63.675 //y=1.56
c770 ( 209 0 ) capacitor c=0.0168481f //x=63.675 //y=1.25
c771 ( 208 0 ) capacitor c=0.0174783f //x=63.675 //y=0.905
c772 ( 203 0 ) capacitor c=0.0245352f //x=54.725 //y=4.79
c773 ( 202 0 ) capacitor c=0.0825763f //x=54.48 //y=1.915
c774 ( 201 0 ) capacitor c=0.0170266f //x=54.48 //y=1.45
c775 ( 200 0 ) capacitor c=0.018609f //x=54.48 //y=1.22
c776 ( 199 0 ) capacitor c=0.0187309f //x=54.48 //y=0.91
c777 ( 193 0 ) capacitor c=0.014725f //x=54.325 //y=1.375
c778 ( 191 0 ) capacitor c=0.0146567f //x=54.325 //y=0.755
c779 ( 190 0 ) capacitor c=0.0335408f //x=53.955 //y=1.22
c780 ( 189 0 ) capacitor c=0.0173761f //x=53.955 //y=0.91
c781 ( 188 0 ) capacitor c=0.0429696f //x=39.785 //y=1.25
c782 ( 187 0 ) capacitor c=0.0192208f //x=39.785 //y=0.905
c783 ( 181 0 ) capacitor c=0.0148884f //x=39.63 //y=1.405
c784 ( 179 0 ) capacitor c=0.0157803f //x=39.63 //y=0.75
c785 ( 177 0 ) capacitor c=0.0295235f //x=39.625 //y=4.79
c786 ( 172 0 ) capacitor c=0.0205163f //x=39.255 //y=1.56
c787 ( 171 0 ) capacitor c=0.0168481f //x=39.255 //y=1.25
c788 ( 170 0 ) capacitor c=0.0174783f //x=39.255 //y=0.905
c789 ( 165 0 ) capacitor c=0.0245352f //x=30.305 //y=4.79
c790 ( 164 0 ) capacitor c=0.0825763f //x=30.06 //y=1.915
c791 ( 163 0 ) capacitor c=0.0170266f //x=30.06 //y=1.45
c792 ( 162 0 ) capacitor c=0.018609f //x=30.06 //y=1.22
c793 ( 161 0 ) capacitor c=0.0187309f //x=30.06 //y=0.91
c794 ( 155 0 ) capacitor c=0.014725f //x=29.905 //y=1.375
c795 ( 153 0 ) capacitor c=0.0146567f //x=29.905 //y=0.755
c796 ( 152 0 ) capacitor c=0.0335408f //x=29.535 //y=1.22
c797 ( 151 0 ) capacitor c=0.0173761f //x=29.535 //y=0.91
c798 ( 150 0 ) capacitor c=0.0429696f //x=15.365 //y=1.25
c799 ( 149 0 ) capacitor c=0.0192208f //x=15.365 //y=0.905
c800 ( 143 0 ) capacitor c=0.0148884f //x=15.21 //y=1.405
c801 ( 141 0 ) capacitor c=0.0157803f //x=15.21 //y=0.75
c802 ( 139 0 ) capacitor c=0.0295235f //x=15.205 //y=4.79
c803 ( 134 0 ) capacitor c=0.0205163f //x=14.835 //y=1.56
c804 ( 133 0 ) capacitor c=0.0168481f //x=14.835 //y=1.25
c805 ( 132 0 ) capacitor c=0.0174783f //x=14.835 //y=0.905
c806 ( 127 0 ) capacitor c=0.0245352f //x=5.885 //y=4.79
c807 ( 126 0 ) capacitor c=0.0826403f //x=5.64 //y=1.915
c808 ( 125 0 ) capacitor c=0.0170266f //x=5.64 //y=1.45
c809 ( 124 0 ) capacitor c=0.018609f //x=5.64 //y=1.22
c810 ( 123 0 ) capacitor c=0.0187309f //x=5.64 //y=0.91
c811 ( 117 0 ) capacitor c=0.014725f //x=5.485 //y=1.375
c812 ( 115 0 ) capacitor c=0.0146567f //x=5.485 //y=0.755
c813 ( 114 0 ) capacitor c=0.0335408f //x=5.115 //y=1.22
c814 ( 113 0 ) capacitor c=0.0173761f //x=5.115 //y=0.91
c815 ( 112 0 ) capacitor c=0.15358f //x=64.12 //y=6.02
c816 ( 111 0 ) capacitor c=0.110281f //x=63.68 //y=6.02
c817 ( 110 0 ) capacitor c=0.110114f //x=54.8 //y=6.02
c818 ( 109 0 ) capacitor c=0.11012f //x=54.36 //y=6.02
c819 ( 108 0 ) capacitor c=0.15358f //x=39.7 //y=6.02
c820 ( 107 0 ) capacitor c=0.110281f //x=39.26 //y=6.02
c821 ( 106 0 ) capacitor c=0.110114f //x=30.38 //y=6.02
c822 ( 105 0 ) capacitor c=0.11012f //x=29.94 //y=6.02
c823 ( 104 0 ) capacitor c=0.15358f //x=15.28 //y=6.02
c824 ( 103 0 ) capacitor c=0.110281f //x=14.84 //y=6.02
c825 ( 102 0 ) capacitor c=0.110114f //x=5.96 //y=6.02
c826 ( 101 0 ) capacitor c=0.11012f //x=5.52 //y=6.02
c827 ( 84 0 ) capacitor c=0.0687295f //x=63.64 //y=2.08
c828 ( 82 0 ) capacitor c=0.00369614f //x=63.64 //y=4.535
c829 ( 74 0 ) capacitor c=0.0900341f //x=54.39 //y=2.08
c830 ( 68 0 ) capacitor c=0.0687295f //x=39.22 //y=2.08
c831 ( 66 0 ) capacitor c=0.00369614f //x=39.22 //y=4.535
c832 ( 58 0 ) capacitor c=0.0900341f //x=29.97 //y=2.08
c833 ( 51 0 ) capacitor c=0.0707124f //x=14.8 //y=2.08
c834 ( 49 0 ) capacitor c=0.00369614f //x=14.8 //y=4.535
c835 ( 39 0 ) capacitor c=0.0953538f //x=5.55 //y=2.08
c836 ( 10 0 ) capacitor c=0.00697397f //x=54.505 //y=4.44
c837 ( 9 0 ) capacitor c=0.213744f //x=63.525 //y=4.44
c838 ( 8 0 ) capacitor c=0.00680508f //x=39.335 //y=4.44
c839 ( 7 0 ) capacitor c=0.354845f //x=54.275 //y=4.44
c840 ( 6 0 ) capacitor c=0.00697397f //x=30.085 //y=4.44
c841 ( 5 0 ) capacitor c=0.201328f //x=39.105 //y=4.44
c842 ( 4 0 ) capacitor c=0.00680508f //x=14.915 //y=4.44
c843 ( 3 0 ) capacitor c=0.353849f //x=29.855 //y=4.44
c844 ( 2 0 ) capacitor c=0.0154455f //x=5.665 //y=4.44
c845 ( 1 0 ) capacitor c=0.201328f //x=14.685 //y=4.44
r846 (  293 294 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=63.67 //y=4.79 //x2=63.67 //y2=4.865
r847 (  291 293 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=63.67 //y=4.7 //x2=63.67 //y2=4.79
r848 (  287 288 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=63.64 //y=2.08 //x2=63.64 //y2=1.915
r849 (  280 281 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=54.39 //y=4.79 //x2=54.39 //y2=4.865
r850 (  278 280 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=54.39 //y=4.7 //x2=54.39 //y2=4.79
r851 (  269 270 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=39.25 //y=4.79 //x2=39.25 //y2=4.865
r852 (  267 269 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=39.25 //y=4.7 //x2=39.25 //y2=4.79
r853 (  263 264 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=39.22 //y=2.08 //x2=39.22 //y2=1.915
r854 (  256 257 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=29.97 //y=4.79 //x2=29.97 //y2=4.865
r855 (  254 256 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=29.97 //y=4.7 //x2=29.97 //y2=4.79
r856 (  245 246 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=14.83 //y=4.79 //x2=14.83 //y2=4.865
r857 (  243 245 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=14.83 //y=4.7 //x2=14.83 //y2=4.79
r858 (  239 240 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=14.8 //y=2.08 //x2=14.8 //y2=1.915
r859 (  232 233 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=5.55 //y=4.79 //x2=5.55 //y2=4.865
r860 (  230 232 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=5.55 //y=4.7 //x2=5.55 //y2=4.79
r861 (  226 298 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.205 //y=1.25 //x2=64.165 //y2=1.405
r862 (  225 297 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.205 //y=0.905 //x2=64.165 //y2=0.75
r863 (  225 226 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=64.205 //y=0.905 //x2=64.205 //y2=1.25
r864 (  220 296 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.83 //y=1.405 //x2=63.715 //y2=1.405
r865 (  219 298 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.05 //y=1.405 //x2=64.165 //y2=1.405
r866 (  218 295 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.83 //y=0.75 //x2=63.715 //y2=0.75
r867 (  217 297 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.05 //y=0.75 //x2=64.165 //y2=0.75
r868 (  217 218 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=64.05 //y=0.75 //x2=63.83 //y2=0.75
r869 (  216 293 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=63.805 //y=4.79 //x2=63.67 //y2=4.79
r870 (  215 222 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=64.045 //y=4.79 //x2=64.12 //y2=4.865
r871 (  215 216 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=64.045 //y=4.79 //x2=63.805 //y2=4.79
r872 (  210 296 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.675 //y=1.56 //x2=63.715 //y2=1.405
r873 (  210 288 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=63.675 //y=1.56 //x2=63.675 //y2=1.915
r874 (  209 296 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.675 //y=1.25 //x2=63.715 //y2=1.405
r875 (  208 295 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.675 //y=0.905 //x2=63.715 //y2=0.75
r876 (  208 209 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.675 //y=0.905 //x2=63.675 //y2=1.25
r877 (  204 280 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=54.525 //y=4.79 //x2=54.39 //y2=4.79
r878 (  203 205 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=54.725 //y=4.79 //x2=54.8 //y2=4.865
r879 (  203 204 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=54.725 //y=4.79 //x2=54.525 //y2=4.79
r880 (  202 285 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=54.48 //y=1.915 //x2=54.405 //y2=2.08
r881 (  201 283 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=54.48 //y=1.45 //x2=54.44 //y2=1.375
r882 (  201 202 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=54.48 //y=1.45 //x2=54.48 //y2=1.915
r883 (  200 283 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.48 //y=1.22 //x2=54.44 //y2=1.375
r884 (  199 282 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.48 //y=0.91 //x2=54.44 //y2=0.755
r885 (  199 200 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=54.48 //y=0.91 //x2=54.48 //y2=1.22
r886 (  194 276 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.11 //y=1.375 //x2=53.995 //y2=1.375
r887 (  193 283 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.325 //y=1.375 //x2=54.44 //y2=1.375
r888 (  192 275 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.11 //y=0.755 //x2=53.995 //y2=0.755
r889 (  191 282 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.325 //y=0.755 //x2=54.44 //y2=0.755
r890 (  191 192 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=54.325 //y=0.755 //x2=54.11 //y2=0.755
r891 (  190 276 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.955 //y=1.22 //x2=53.995 //y2=1.375
r892 (  189 275 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.955 //y=0.91 //x2=53.995 //y2=0.755
r893 (  189 190 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=53.955 //y=0.91 //x2=53.955 //y2=1.22
r894 (  188 274 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.785 //y=1.25 //x2=39.745 //y2=1.405
r895 (  187 273 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.785 //y=0.905 //x2=39.745 //y2=0.75
r896 (  187 188 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=39.785 //y=0.905 //x2=39.785 //y2=1.25
r897 (  182 272 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.41 //y=1.405 //x2=39.295 //y2=1.405
r898 (  181 274 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.63 //y=1.405 //x2=39.745 //y2=1.405
r899 (  180 271 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.41 //y=0.75 //x2=39.295 //y2=0.75
r900 (  179 273 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.63 //y=0.75 //x2=39.745 //y2=0.75
r901 (  179 180 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=39.63 //y=0.75 //x2=39.41 //y2=0.75
r902 (  178 269 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=39.385 //y=4.79 //x2=39.25 //y2=4.79
r903 (  177 184 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=39.625 //y=4.79 //x2=39.7 //y2=4.865
r904 (  177 178 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=39.625 //y=4.79 //x2=39.385 //y2=4.79
r905 (  172 272 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.255 //y=1.56 //x2=39.295 //y2=1.405
r906 (  172 264 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=39.255 //y=1.56 //x2=39.255 //y2=1.915
r907 (  171 272 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.255 //y=1.25 //x2=39.295 //y2=1.405
r908 (  170 271 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.255 //y=0.905 //x2=39.295 //y2=0.75
r909 (  170 171 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=39.255 //y=0.905 //x2=39.255 //y2=1.25
r910 (  166 256 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=30.105 //y=4.79 //x2=29.97 //y2=4.79
r911 (  165 167 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=30.305 //y=4.79 //x2=30.38 //y2=4.865
r912 (  165 166 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=30.305 //y=4.79 //x2=30.105 //y2=4.79
r913 (  164 261 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=30.06 //y=1.915 //x2=29.985 //y2=2.08
r914 (  163 259 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=30.06 //y=1.45 //x2=30.02 //y2=1.375
r915 (  163 164 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=30.06 //y=1.45 //x2=30.06 //y2=1.915
r916 (  162 259 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.06 //y=1.22 //x2=30.02 //y2=1.375
r917 (  161 258 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.06 //y=0.91 //x2=30.02 //y2=0.755
r918 (  161 162 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=30.06 //y=0.91 //x2=30.06 //y2=1.22
r919 (  156 252 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.69 //y=1.375 //x2=29.575 //y2=1.375
r920 (  155 259 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.905 //y=1.375 //x2=30.02 //y2=1.375
r921 (  154 251 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.69 //y=0.755 //x2=29.575 //y2=0.755
r922 (  153 258 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.905 //y=0.755 //x2=30.02 //y2=0.755
r923 (  153 154 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=29.905 //y=0.755 //x2=29.69 //y2=0.755
r924 (  152 252 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.535 //y=1.22 //x2=29.575 //y2=1.375
r925 (  151 251 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.535 //y=0.91 //x2=29.575 //y2=0.755
r926 (  151 152 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=29.535 //y=0.91 //x2=29.535 //y2=1.22
r927 (  150 250 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.365 //y=1.25 //x2=15.325 //y2=1.405
r928 (  149 249 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.365 //y=0.905 //x2=15.325 //y2=0.75
r929 (  149 150 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.365 //y=0.905 //x2=15.365 //y2=1.25
r930 (  144 248 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.99 //y=1.405 //x2=14.875 //y2=1.405
r931 (  143 250 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.21 //y=1.405 //x2=15.325 //y2=1.405
r932 (  142 247 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.99 //y=0.75 //x2=14.875 //y2=0.75
r933 (  141 249 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.21 //y=0.75 //x2=15.325 //y2=0.75
r934 (  141 142 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.21 //y=0.75 //x2=14.99 //y2=0.75
r935 (  140 245 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=14.965 //y=4.79 //x2=14.83 //y2=4.79
r936 (  139 146 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.79 //x2=15.28 //y2=4.865
r937 (  139 140 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.79 //x2=14.965 //y2=4.79
r938 (  134 248 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.56 //x2=14.875 //y2=1.405
r939 (  134 240 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.56 //x2=14.835 //y2=1.915
r940 (  133 248 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.25 //x2=14.875 //y2=1.405
r941 (  132 247 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=0.905 //x2=14.875 //y2=0.75
r942 (  132 133 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.835 //y=0.905 //x2=14.835 //y2=1.25
r943 (  128 232 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=5.685 //y=4.79 //x2=5.55 //y2=4.79
r944 (  127 129 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.885 //y=4.79 //x2=5.96 //y2=4.865
r945 (  127 128 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=5.885 //y=4.79 //x2=5.685 //y2=4.79
r946 (  126 237 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.915 //x2=5.565 //y2=2.08
r947 (  125 235 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.45 //x2=5.6 //y2=1.375
r948 (  125 126 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.45 //x2=5.64 //y2=1.915
r949 (  124 235 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.22 //x2=5.6 //y2=1.375
r950 (  123 234 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.64 //y=0.91 //x2=5.6 //y2=0.755
r951 (  123 124 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=5.64 //y=0.91 //x2=5.64 //y2=1.22
r952 (  118 228 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.27 //y=1.375 //x2=5.155 //y2=1.375
r953 (  117 235 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.485 //y=1.375 //x2=5.6 //y2=1.375
r954 (  116 227 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.27 //y=0.755 //x2=5.155 //y2=0.755
r955 (  115 234 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.485 //y=0.755 //x2=5.6 //y2=0.755
r956 (  115 116 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=5.485 //y=0.755 //x2=5.27 //y2=0.755
r957 (  114 228 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.115 //y=1.22 //x2=5.155 //y2=1.375
r958 (  113 227 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.115 //y=0.91 //x2=5.155 //y2=0.755
r959 (  113 114 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=5.115 //y=0.91 //x2=5.115 //y2=1.22
r960 (  112 222 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=64.12 //y=6.02 //x2=64.12 //y2=4.865
r961 (  111 294 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=63.68 //y=6.02 //x2=63.68 //y2=4.865
r962 (  110 205 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.8 //y=6.02 //x2=54.8 //y2=4.865
r963 (  109 281 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.36 //y=6.02 //x2=54.36 //y2=4.865
r964 (  108 184 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=39.7 //y=6.02 //x2=39.7 //y2=4.865
r965 (  107 270 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=39.26 //y=6.02 //x2=39.26 //y2=4.865
r966 (  106 167 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.38 //y=6.02 //x2=30.38 //y2=4.865
r967 (  105 257 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=29.94 //y=6.02 //x2=29.94 //y2=4.865
r968 (  104 146 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.28 //y=6.02 //x2=15.28 //y2=4.865
r969 (  103 246 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.84 //y=6.02 //x2=14.84 //y2=4.865
r970 (  102 129 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.96 //y=6.02 //x2=5.96 //y2=4.865
r971 (  101 233 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.52 //y=6.02 //x2=5.52 //y2=4.865
r972 (  100 219 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.94 //y=1.405 //x2=64.05 //y2=1.405
r973 (  100 220 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.94 //y=1.405 //x2=63.83 //y2=1.405
r974 (  99 193 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=54.217 //y=1.375 //x2=54.325 //y2=1.375
r975 (  99 194 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=54.217 //y=1.375 //x2=54.11 //y2=1.375
r976 (  98 181 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.52 //y=1.405 //x2=39.63 //y2=1.405
r977 (  98 182 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.52 //y=1.405 //x2=39.41 //y2=1.405
r978 (  97 155 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=29.797 //y=1.375 //x2=29.905 //y2=1.375
r979 (  97 156 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=29.797 //y=1.375 //x2=29.69 //y2=1.375
r980 (  96 143 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.1 //y=1.405 //x2=15.21 //y2=1.405
r981 (  96 144 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.1 //y=1.405 //x2=14.99 //y2=1.405
r982 (  95 117 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=5.377 //y=1.375 //x2=5.485 //y2=1.375
r983 (  95 118 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=5.377 //y=1.375 //x2=5.27 //y2=1.375
r984 (  94 291 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.67 //y=4.7 //x2=63.67 //y2=4.7
r985 (  92 267 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.25 //y=4.7 //x2=39.25 //y2=4.7
r986 (  90 243 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.83 //y=4.7 //x2=14.83 //y2=4.7
r987 (  84 287 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.64 //y=2.08 //x2=63.64 //y2=2.08
r988 (  82 94 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=63.64 //y=4.535 //x2=63.655 //y2=4.7
r989 (  80 278 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.39 //y=4.7 //x2=54.39 //y2=4.7
r990 (  74 285 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.39 //y=2.08 //x2=54.39 //y2=2.08
r991 (  68 263 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.22 //y=2.08 //x2=39.22 //y2=2.08
r992 (  66 92 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=39.22 //y=4.535 //x2=39.235 //y2=4.7
r993 (  64 254 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.97 //y=4.7 //x2=29.97 //y2=4.7
r994 (  58 261 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.97 //y=2.08 //x2=29.97 //y2=2.08
r995 (  51 239 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.8 //y=2.08 //x2=14.8 //y2=2.08
r996 (  49 90 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=14.8 //y=4.535 //x2=14.815 //y2=4.7
r997 (  47 230 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=4.7 //x2=5.55 //y2=4.7
r998 (  39 237 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=2.08 //x2=5.55 //y2=2.08
r999 (  37 82 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=63.64 //y=4.44 //x2=63.64 //y2=4.535
r1000 (  36 37 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=63.64 //y=2.59 //x2=63.64 //y2=4.44
r1001 (  36 84 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=63.64 //y=2.59 //x2=63.64 //y2=2.08
r1002 (  35 80 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=54.39 //y=4.44 //x2=54.39 //y2=4.7
r1003 (  34 35 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=54.39 //y=3.7 //x2=54.39 //y2=4.44
r1004 (  34 74 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=54.39 //y=3.7 //x2=54.39 //y2=2.08
r1005 (  33 66 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=39.22 //y=4.44 //x2=39.22 //y2=4.535
r1006 (  32 33 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=39.22 //y=2.59 //x2=39.22 //y2=4.44
r1007 (  32 68 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=39.22 //y=2.59 //x2=39.22 //y2=2.08
r1008 (  31 64 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=29.97 //y=4.44 //x2=29.97 //y2=4.7
r1009 (  30 31 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=29.97 //y=3.7 //x2=29.97 //y2=4.44
r1010 (  30 58 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=29.97 //y=3.7 //x2=29.97 //y2=2.08
r1011 (  29 49 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=14.8 //y=4.44 //x2=14.8 //y2=4.535
r1012 (  28 29 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=14.8 //y=3.33 //x2=14.8 //y2=4.44
r1013 (  27 28 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=14.8 //y=2.59 //x2=14.8 //y2=3.33
r1014 (  27 51 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=14.8 //y=2.59 //x2=14.8 //y2=2.08
r1015 (  26 47 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=5.55 //y=4.44 //x2=5.55 //y2=4.7
r1016 (  25 26 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=5.55 //y=3.7 //x2=5.55 //y2=4.44
r1017 (  24 25 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=5.55 //y=3.33 //x2=5.55 //y2=3.7
r1018 (  23 24 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=5.55 //y=2.22 //x2=5.55 //y2=3.33
r1019 (  23 39 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=5.55 //y=2.22 //x2=5.55 //y2=2.08
r1020 (  22 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=63.64 //y=4.44 //x2=63.64 //y2=4.44
r1021 (  20 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=54.39 //y=4.44 //x2=54.39 //y2=4.44
r1022 (  18 33 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=39.22 //y=4.44 //x2=39.22 //y2=4.44
r1023 (  16 31 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=29.97 //y=4.44 //x2=29.97 //y2=4.44
r1024 (  14 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.8 //y=4.44 //x2=14.8 //y2=4.44
r1025 (  12 26 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.55 //y=4.44 //x2=5.55 //y2=4.44
r1026 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=54.505 //y=4.44 //x2=54.39 //y2=4.44
r1027 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.525 //y=4.44 //x2=63.64 //y2=4.44
r1028 (  9 10 ) resistor r=8.60687 //w=0.131 //l=9.02 //layer=m1 \
 //thickness=0.36 //x=63.525 //y=4.44 //x2=54.505 //y2=4.44
r1029 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=39.335 //y=4.44 //x2=39.22 //y2=4.44
r1030 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=54.275 //y=4.44 //x2=54.39 //y2=4.44
r1031 (  7 8 ) resistor r=14.2557 //w=0.131 //l=14.94 //layer=m1 \
 //thickness=0.36 //x=54.275 //y=4.44 //x2=39.335 //y2=4.44
r1032 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=30.085 //y=4.44 //x2=29.97 //y2=4.44
r1033 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=39.105 //y=4.44 //x2=39.22 //y2=4.44
r1034 (  5 6 ) resistor r=8.60687 //w=0.131 //l=9.02 //layer=m1 \
 //thickness=0.36 //x=39.105 //y=4.44 //x2=30.085 //y2=4.44
r1035 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.915 //y=4.44 //x2=14.8 //y2=4.44
r1036 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=29.855 //y=4.44 //x2=29.97 //y2=4.44
r1037 (  3 4 ) resistor r=14.2557 //w=0.131 //l=14.94 //layer=m1 \
 //thickness=0.36 //x=29.855 //y=4.44 //x2=14.915 //y2=4.44
r1038 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.665 //y=4.44 //x2=5.55 //y2=4.44
r1039 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.685 //y=4.44 //x2=14.8 //y2=4.44
r1040 (  1 2 ) resistor r=8.60687 //w=0.131 //l=9.02 //layer=m1 \
 //thickness=0.36 //x=14.685 //y=4.44 //x2=5.665 //y2=4.44
ends PM_TMRDFFSNQNX1\%CLK

subckt PM_TMRDFFSNQNX1\%noxref_17 ( 1 2 3 4 11 13 23 24 31 39 45 46 50 52 61 \
 62 64 65 67 68 69 70 71 72 73 74 75 80 82 84 90 91 92 93 94 95 99 101 104 105 \
 110 111 114 128 131 133 134 135 )
c291 ( 135 0 ) capacitor c=0.023087f //x=55.315 //y=5.02
c292 ( 134 0 ) capacitor c=0.023519f //x=54.435 //y=5.02
c293 ( 133 0 ) capacitor c=0.0224735f //x=53.555 //y=5.02
c294 ( 131 0 ) capacitor c=0.00853354f //x=55.565 //y=0.915
c295 ( 128 0 ) capacitor c=0.0597793f //x=66.23 //y=4.7
c296 ( 114 0 ) capacitor c=0.0331095f //x=50.72 //y=4.7
c297 ( 111 0 ) capacitor c=0.0279499f //x=50.69 //y=1.915
c298 ( 110 0 ) capacitor c=0.0421676f //x=50.69 //y=2.08
c299 ( 105 0 ) capacitor c=0.0318948f //x=66.565 //y=1.21
c300 ( 104 0 ) capacitor c=0.0187384f //x=66.565 //y=0.865
c301 ( 101 0 ) capacitor c=0.0141798f //x=66.41 //y=1.365
c302 ( 99 0 ) capacitor c=0.0149844f //x=66.41 //y=0.71
c303 ( 95 0 ) capacitor c=0.0813322f //x=66.035 //y=1.915
c304 ( 94 0 ) capacitor c=0.0229267f //x=66.035 //y=1.52
c305 ( 93 0 ) capacitor c=0.0234352f //x=66.035 //y=1.21
c306 ( 92 0 ) capacitor c=0.0199343f //x=66.035 //y=0.865
c307 ( 91 0 ) capacitor c=0.0429696f //x=51.255 //y=1.25
c308 ( 90 0 ) capacitor c=0.0192208f //x=51.255 //y=0.905
c309 ( 84 0 ) capacitor c=0.0148884f //x=51.1 //y=1.405
c310 ( 82 0 ) capacitor c=0.0157803f //x=51.1 //y=0.75
c311 ( 80 0 ) capacitor c=0.0295235f //x=51.095 //y=4.79
c312 ( 75 0 ) capacitor c=0.0205163f //x=50.725 //y=1.56
c313 ( 74 0 ) capacitor c=0.0168481f //x=50.725 //y=1.25
c314 ( 73 0 ) capacitor c=0.0174783f //x=50.725 //y=0.905
c315 ( 72 0 ) capacitor c=0.110275f //x=66.57 //y=6.02
c316 ( 71 0 ) capacitor c=0.154305f //x=66.13 //y=6.02
c317 ( 70 0 ) capacitor c=0.15358f //x=51.17 //y=6.02
c318 ( 69 0 ) capacitor c=0.110281f //x=50.73 //y=6.02
c319 ( 65 0 ) capacitor c=0.0715637f //x=56.237 //y=3.905
c320 ( 64 0 ) capacitor c=0.0101843f //x=56.235 //y=4.07
c321 ( 62 0 ) capacitor c=0.00106608f //x=55.46 //y=5.155
c322 ( 61 0 ) capacitor c=0.00207162f //x=54.58 //y=5.155
c323 ( 52 0 ) capacitor c=0.0878627f //x=66.23 //y=2.08
c324 ( 50 0 ) capacitor c=0.0236247f //x=56.24 //y=5.07
c325 ( 46 0 ) capacitor c=0.00398962f //x=55.84 //y=1.665
c326 ( 45 0 ) capacitor c=0.0135805f //x=56.155 //y=1.665
c327 ( 39 0 ) capacitor c=0.0281378f //x=56.155 //y=5.155
c328 ( 31 0 ) capacitor c=0.0176454f //x=55.375 //y=5.155
c329 ( 24 0 ) capacitor c=0.00332903f //x=53.785 //y=5.155
c330 ( 23 0 ) capacitor c=0.014837f //x=54.495 //y=5.155
c331 ( 13 0 ) capacitor c=0.0676664f //x=50.69 //y=2.08
c332 ( 11 0 ) capacitor c=0.00453889f //x=50.69 //y=4.535
c333 ( 4 0 ) capacitor c=0.00551102f //x=56.35 //y=4.07
c334 ( 3 0 ) capacitor c=0.173174f //x=66.115 //y=4.07
c335 ( 2 0 ) capacitor c=0.0100678f //x=50.805 //y=4.07
c336 ( 1 0 ) capacitor c=0.0882171f //x=56.12 //y=4.07
r337 (  126 128 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=66.13 //y=4.7 //x2=66.23 //y2=4.7
r338 (  116 117 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=50.72 //y=4.79 //x2=50.72 //y2=4.865
r339 (  114 116 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=50.72 //y=4.7 //x2=50.72 //y2=4.79
r340 (  110 111 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=50.69 //y=2.08 //x2=50.69 //y2=1.915
r341 (  106 128 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=66.57 //y=4.865 //x2=66.23 //y2=4.7
r342 (  105 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.565 //y=1.21 //x2=66.525 //y2=1.365
r343 (  104 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.565 //y=0.865 //x2=66.525 //y2=0.71
r344 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=66.565 //y=0.865 //x2=66.565 //y2=1.21
r345 (  102 125 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.19 //y=1.365 //x2=66.075 //y2=1.365
r346 (  101 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.41 //y=1.365 //x2=66.525 //y2=1.365
r347 (  100 124 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.19 //y=0.71 //x2=66.075 //y2=0.71
r348 (  99 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.41 //y=0.71 //x2=66.525 //y2=0.71
r349 (  99 100 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=66.41 //y=0.71 //x2=66.19 //y2=0.71
r350 (  96 126 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=66.13 //y=4.865 //x2=66.13 //y2=4.7
r351 (  95 123 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=66.035 //y=1.915 //x2=66.23 //y2=2.08
r352 (  94 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.035 //y=1.52 //x2=66.075 //y2=1.365
r353 (  94 95 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=66.035 //y=1.52 //x2=66.035 //y2=1.915
r354 (  93 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.035 //y=1.21 //x2=66.075 //y2=1.365
r355 (  92 124 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.035 //y=0.865 //x2=66.075 //y2=0.71
r356 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=66.035 //y=0.865 //x2=66.035 //y2=1.21
r357 (  91 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.255 //y=1.25 //x2=51.215 //y2=1.405
r358 (  90 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.255 //y=0.905 //x2=51.215 //y2=0.75
r359 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=51.255 //y=0.905 //x2=51.255 //y2=1.25
r360 (  85 119 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.88 //y=1.405 //x2=50.765 //y2=1.405
r361 (  84 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.1 //y=1.405 //x2=51.215 //y2=1.405
r362 (  83 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.88 //y=0.75 //x2=50.765 //y2=0.75
r363 (  82 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.1 //y=0.75 //x2=51.215 //y2=0.75
r364 (  82 83 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=51.1 //y=0.75 //x2=50.88 //y2=0.75
r365 (  81 116 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=50.855 //y=4.79 //x2=50.72 //y2=4.79
r366 (  80 87 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=51.095 //y=4.79 //x2=51.17 //y2=4.865
r367 (  80 81 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=51.095 //y=4.79 //x2=50.855 //y2=4.79
r368 (  75 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.725 //y=1.56 //x2=50.765 //y2=1.405
r369 (  75 111 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=50.725 //y=1.56 //x2=50.725 //y2=1.915
r370 (  74 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.725 //y=1.25 //x2=50.765 //y2=1.405
r371 (  73 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.725 //y=0.905 //x2=50.765 //y2=0.75
r372 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=50.725 //y=0.905 //x2=50.725 //y2=1.25
r373 (  72 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.57 //y=6.02 //x2=66.57 //y2=4.865
r374 (  71 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.13 //y=6.02 //x2=66.13 //y2=4.865
r375 (  70 87 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=51.17 //y=6.02 //x2=51.17 //y2=4.865
r376 (  69 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.73 //y=6.02 //x2=50.73 //y2=4.865
r377 (  68 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.3 //y=1.365 //x2=66.41 //y2=1.365
r378 (  68 102 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.3 //y=1.365 //x2=66.19 //y2=1.365
r379 (  67 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.99 //y=1.405 //x2=51.1 //y2=1.405
r380 (  67 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.99 //y=1.405 //x2=50.88 //y2=1.405
r381 (  64 66 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=56.237 //y=4.07 //x2=56.237 //y2=4.235
r382 (  64 65 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=56.237 //y=4.07 //x2=56.237 //y2=3.905
r383 (  60 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.72 //y=4.7 //x2=50.72 //y2=4.7
r384 (  57 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.23 //y=4.7 //x2=66.23 //y2=4.7
r385 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=66.23 //y=4.07 //x2=66.23 //y2=4.7
r386 (  52 123 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.23 //y=2.08 //x2=66.23 //y2=2.08
r387 (  52 55 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=66.23 //y=2.08 //x2=66.23 //y2=4.07
r388 (  50 66 ) resistor r=57.1551 //w=0.187 //l=0.835 //layer=li \
 //thickness=0.1 //x=56.24 //y=5.07 //x2=56.24 //y2=4.235
r389 (  47 65 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=56.24 //y=1.75 //x2=56.24 //y2=3.905
r390 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.155 //y=1.665 //x2=56.24 //y2=1.75
r391 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=56.155 //y=1.665 //x2=55.84 //y2=1.665
r392 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=55.755 //y=1.58 //x2=55.84 //y2=1.665
r393 (  41 131 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=55.755 //y=1.58 //x2=55.755 //y2=1.01
r394 (  40 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.545 //y=5.155 //x2=55.46 //y2=5.155
r395 (  39 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.155 //y=5.155 //x2=56.24 //y2=5.07
r396 (  39 40 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=56.155 //y=5.155 //x2=55.545 //y2=5.155
r397 (  33 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.46 //y=5.24 //x2=55.46 //y2=5.155
r398 (  33 135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.46 //y=5.24 //x2=55.46 //y2=5.725
r399 (  32 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.665 //y=5.155 //x2=54.58 //y2=5.155
r400 (  31 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.375 //y=5.155 //x2=55.46 //y2=5.155
r401 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=55.375 //y=5.155 //x2=54.665 //y2=5.155
r402 (  25 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.58 //y=5.24 //x2=54.58 //y2=5.155
r403 (  25 134 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.58 //y=5.24 //x2=54.58 //y2=5.725
r404 (  23 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.495 //y=5.155 //x2=54.58 //y2=5.155
r405 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=54.495 //y=5.155 //x2=53.785 //y2=5.155
r406 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=53.7 //y=5.24 //x2=53.785 //y2=5.155
r407 (  17 133 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=53.7 //y=5.24 //x2=53.7 //y2=5.725
r408 (  13 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.69 //y=2.08 //x2=50.69 //y2=2.08
r409 (  13 16 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=50.69 //y=2.08 //x2=50.69 //y2=4.07
r410 (  11 60 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=50.69 //y=4.535 //x2=50.705 //y2=4.7
r411 (  11 16 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=50.69 //y=4.535 //x2=50.69 //y2=4.07
r412 (  10 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.23 //y=4.07 //x2=66.23 //y2=4.07
r413 (  8 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=56.235 //y=4.07 //x2=56.235 //y2=4.07
r414 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=50.69 //y=4.07 //x2=50.69 //y2=4.07
r415 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.35 //y=4.07 //x2=56.235 //y2=4.07
r416 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.115 //y=4.07 //x2=66.23 //y2=4.07
r417 (  3 4 ) resistor r=9.31775 //w=0.131 //l=9.765 //layer=m1 \
 //thickness=0.36 //x=66.115 //y=4.07 //x2=56.35 //y2=4.07
r418 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.805 //y=4.07 //x2=50.69 //y2=4.07
r419 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.12 //y=4.07 //x2=56.235 //y2=4.07
r420 (  1 2 ) resistor r=5.07156 //w=0.131 //l=5.315 //layer=m1 \
 //thickness=0.36 //x=56.12 //y=4.07 //x2=50.805 //y2=4.07
ends PM_TMRDFFSNQNX1\%noxref_17

subckt PM_TMRDFFSNQNX1\%SN ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 31 \
 33 43 52 60 68 77 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 \
 103 104 106 112 113 114 115 116 121 122 123 125 131 132 133 134 135 140 141 \
 142 144 150 151 152 153 154 159 160 161 163 169 170 171 172 173 178 179 180 \
 182 188 189 190 191 192 197 198 199 201 207 208 209 210 211 219 230 241 252 \
 263 274 )
c818 ( 274 0 ) capacitor c=0.0337007f //x=70.67 //y=4.7
c819 ( 263 0 ) capacitor c=0.0335551f //x=59.2 //y=4.7
c820 ( 252 0 ) capacitor c=0.0335551f //x=46.25 //y=4.7
c821 ( 241 0 ) capacitor c=0.0335551f //x=34.78 //y=4.7
c822 ( 230 0 ) capacitor c=0.0335551f //x=21.83 //y=4.7
c823 ( 219 0 ) capacitor c=0.0335551f //x=10.36 //y=4.7
c824 ( 211 0 ) capacitor c=0.0245352f //x=71.005 //y=4.79
c825 ( 210 0 ) capacitor c=0.0827272f //x=70.76 //y=1.915
c826 ( 209 0 ) capacitor c=0.0170266f //x=70.76 //y=1.45
c827 ( 208 0 ) capacitor c=0.018609f //x=70.76 //y=1.22
c828 ( 207 0 ) capacitor c=0.0187309f //x=70.76 //y=0.91
c829 ( 201 0 ) capacitor c=0.014725f //x=70.605 //y=1.375
c830 ( 199 0 ) capacitor c=0.0146567f //x=70.605 //y=0.755
c831 ( 198 0 ) capacitor c=0.0335408f //x=70.235 //y=1.22
c832 ( 197 0 ) capacitor c=0.0173761f //x=70.235 //y=0.91
c833 ( 192 0 ) capacitor c=0.0245352f //x=59.535 //y=4.79
c834 ( 191 0 ) capacitor c=0.0825033f //x=59.29 //y=1.915
c835 ( 190 0 ) capacitor c=0.0170266f //x=59.29 //y=1.45
c836 ( 189 0 ) capacitor c=0.018609f //x=59.29 //y=1.22
c837 ( 188 0 ) capacitor c=0.0187309f //x=59.29 //y=0.91
c838 ( 182 0 ) capacitor c=0.014725f //x=59.135 //y=1.375
c839 ( 180 0 ) capacitor c=0.0146567f //x=59.135 //y=0.755
c840 ( 179 0 ) capacitor c=0.0335408f //x=58.765 //y=1.22
c841 ( 178 0 ) capacitor c=0.0173761f //x=58.765 //y=0.91
c842 ( 173 0 ) capacitor c=0.0245352f //x=46.585 //y=4.79
c843 ( 172 0 ) capacitor c=0.0825033f //x=46.34 //y=1.915
c844 ( 171 0 ) capacitor c=0.0170266f //x=46.34 //y=1.45
c845 ( 170 0 ) capacitor c=0.018609f //x=46.34 //y=1.22
c846 ( 169 0 ) capacitor c=0.0187309f //x=46.34 //y=0.91
c847 ( 163 0 ) capacitor c=0.014725f //x=46.185 //y=1.375
c848 ( 161 0 ) capacitor c=0.0146567f //x=46.185 //y=0.755
c849 ( 160 0 ) capacitor c=0.0335408f //x=45.815 //y=1.22
c850 ( 159 0 ) capacitor c=0.0173761f //x=45.815 //y=0.91
c851 ( 154 0 ) capacitor c=0.0245352f //x=35.115 //y=4.79
c852 ( 153 0 ) capacitor c=0.0825033f //x=34.87 //y=1.915
c853 ( 152 0 ) capacitor c=0.0170266f //x=34.87 //y=1.45
c854 ( 151 0 ) capacitor c=0.018609f //x=34.87 //y=1.22
c855 ( 150 0 ) capacitor c=0.0187309f //x=34.87 //y=0.91
c856 ( 144 0 ) capacitor c=0.014725f //x=34.715 //y=1.375
c857 ( 142 0 ) capacitor c=0.0146567f //x=34.715 //y=0.755
c858 ( 141 0 ) capacitor c=0.0335408f //x=34.345 //y=1.22
c859 ( 140 0 ) capacitor c=0.0173761f //x=34.345 //y=0.91
c860 ( 135 0 ) capacitor c=0.0245352f //x=22.165 //y=4.79
c861 ( 134 0 ) capacitor c=0.0825033f //x=21.92 //y=1.915
c862 ( 133 0 ) capacitor c=0.0170266f //x=21.92 //y=1.45
c863 ( 132 0 ) capacitor c=0.018609f //x=21.92 //y=1.22
c864 ( 131 0 ) capacitor c=0.0187309f //x=21.92 //y=0.91
c865 ( 125 0 ) capacitor c=0.014725f //x=21.765 //y=1.375
c866 ( 123 0 ) capacitor c=0.0146567f //x=21.765 //y=0.755
c867 ( 122 0 ) capacitor c=0.0335408f //x=21.395 //y=1.22
c868 ( 121 0 ) capacitor c=0.0173761f //x=21.395 //y=0.91
c869 ( 116 0 ) capacitor c=0.0245352f //x=10.695 //y=4.79
c870 ( 115 0 ) capacitor c=0.0826756f //x=10.45 //y=1.915
c871 ( 114 0 ) capacitor c=0.0170266f //x=10.45 //y=1.45
c872 ( 113 0 ) capacitor c=0.018609f //x=10.45 //y=1.22
c873 ( 112 0 ) capacitor c=0.0187309f //x=10.45 //y=0.91
c874 ( 106 0 ) capacitor c=0.014725f //x=10.295 //y=1.375
c875 ( 104 0 ) capacitor c=0.0146567f //x=10.295 //y=0.755
c876 ( 103 0 ) capacitor c=0.0335408f //x=9.925 //y=1.22
c877 ( 102 0 ) capacitor c=0.0173761f //x=9.925 //y=0.91
c878 ( 101 0 ) capacitor c=0.110114f //x=71.08 //y=6.02
c879 ( 100 0 ) capacitor c=0.11012f //x=70.64 //y=6.02
c880 ( 99 0 ) capacitor c=0.110114f //x=59.61 //y=6.02
c881 ( 98 0 ) capacitor c=0.11012f //x=59.17 //y=6.02
c882 ( 97 0 ) capacitor c=0.110114f //x=46.66 //y=6.02
c883 ( 96 0 ) capacitor c=0.11012f //x=46.22 //y=6.02
c884 ( 95 0 ) capacitor c=0.110114f //x=35.19 //y=6.02
c885 ( 94 0 ) capacitor c=0.11012f //x=34.75 //y=6.02
c886 ( 93 0 ) capacitor c=0.110114f //x=22.24 //y=6.02
c887 ( 92 0 ) capacitor c=0.11012f //x=21.8 //y=6.02
c888 ( 91 0 ) capacitor c=0.110114f //x=10.77 //y=6.02
c889 ( 90 0 ) capacitor c=0.11012f //x=10.33 //y=6.02
c890 ( 77 0 ) capacitor c=0.0905446f //x=70.67 //y=2.08
c891 ( 68 0 ) capacitor c=0.0895052f //x=59.2 //y=2.08
c892 ( 60 0 ) capacitor c=0.0878512f //x=46.25 //y=2.08
c893 ( 52 0 ) capacitor c=0.0895052f //x=34.78 //y=2.08
c894 ( 43 0 ) capacitor c=0.0904947f //x=21.83 //y=2.08
c895 ( 33 0 ) capacitor c=0.0921487f //x=10.36 //y=2.08
c896 ( 10 0 ) capacitor c=0.00692137f //x=59.315 //y=2.22
c897 ( 9 0 ) capacitor c=0.263633f //x=70.555 //y=2.22
c898 ( 8 0 ) capacitor c=0.00666809f //x=46.365 //y=2.22
c899 ( 7 0 ) capacitor c=0.252177f //x=59.085 //y=2.22
c900 ( 6 0 ) capacitor c=0.00692137f //x=34.895 //y=2.22
c901 ( 5 0 ) capacitor c=0.237521f //x=46.135 //y=2.22
c902 ( 4 0 ) capacitor c=0.00692137f //x=21.945 //y=2.22
c903 ( 3 0 ) capacitor c=0.266406f //x=34.665 //y=2.22
c904 ( 2 0 ) capacitor c=0.0154797f //x=10.475 //y=2.22
c905 ( 1 0 ) capacitor c=0.248273f //x=21.715 //y=2.22
r906 (  276 277 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=70.67 //y=4.79 //x2=70.67 //y2=4.865
r907 (  274 276 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=70.67 //y=4.7 //x2=70.67 //y2=4.79
r908 (  265 266 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=59.2 //y=4.79 //x2=59.2 //y2=4.865
r909 (  263 265 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=59.2 //y=4.7 //x2=59.2 //y2=4.79
r910 (  254 255 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=46.25 //y=4.79 //x2=46.25 //y2=4.865
r911 (  252 254 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=46.25 //y=4.7 //x2=46.25 //y2=4.79
r912 (  243 244 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=34.78 //y=4.79 //x2=34.78 //y2=4.865
r913 (  241 243 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=34.78 //y=4.7 //x2=34.78 //y2=4.79
r914 (  232 233 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=21.83 //y=4.79 //x2=21.83 //y2=4.865
r915 (  230 232 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=21.83 //y=4.7 //x2=21.83 //y2=4.79
r916 (  221 222 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=10.36 //y=4.79 //x2=10.36 //y2=4.865
r917 (  219 221 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=10.36 //y=4.7 //x2=10.36 //y2=4.79
r918 (  212 276 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=70.805 //y=4.79 //x2=70.67 //y2=4.79
r919 (  211 213 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=71.005 //y=4.79 //x2=71.08 //y2=4.865
r920 (  211 212 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=71.005 //y=4.79 //x2=70.805 //y2=4.79
r921 (  210 281 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=70.76 //y=1.915 //x2=70.685 //y2=2.08
r922 (  209 279 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=70.76 //y=1.45 //x2=70.72 //y2=1.375
r923 (  209 210 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=70.76 //y=1.45 //x2=70.76 //y2=1.915
r924 (  208 279 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.76 //y=1.22 //x2=70.72 //y2=1.375
r925 (  207 278 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.76 //y=0.91 //x2=70.72 //y2=0.755
r926 (  207 208 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=70.76 //y=0.91 //x2=70.76 //y2=1.22
r927 (  202 272 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.39 //y=1.375 //x2=70.275 //y2=1.375
r928 (  201 279 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.605 //y=1.375 //x2=70.72 //y2=1.375
r929 (  200 271 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.39 //y=0.755 //x2=70.275 //y2=0.755
r930 (  199 278 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.605 //y=0.755 //x2=70.72 //y2=0.755
r931 (  199 200 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=70.605 //y=0.755 //x2=70.39 //y2=0.755
r932 (  198 272 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.235 //y=1.22 //x2=70.275 //y2=1.375
r933 (  197 271 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.235 //y=0.91 //x2=70.275 //y2=0.755
r934 (  197 198 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=70.235 //y=0.91 //x2=70.235 //y2=1.22
r935 (  193 265 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=59.335 //y=4.79 //x2=59.2 //y2=4.79
r936 (  192 194 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=59.535 //y=4.79 //x2=59.61 //y2=4.865
r937 (  192 193 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=59.535 //y=4.79 //x2=59.335 //y2=4.79
r938 (  191 270 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=59.29 //y=1.915 //x2=59.215 //y2=2.08
r939 (  190 268 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=59.29 //y=1.45 //x2=59.25 //y2=1.375
r940 (  190 191 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=59.29 //y=1.45 //x2=59.29 //y2=1.915
r941 (  189 268 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.29 //y=1.22 //x2=59.25 //y2=1.375
r942 (  188 267 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.29 //y=0.91 //x2=59.25 //y2=0.755
r943 (  188 189 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=59.29 //y=0.91 //x2=59.29 //y2=1.22
r944 (  183 261 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.92 //y=1.375 //x2=58.805 //y2=1.375
r945 (  182 268 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.135 //y=1.375 //x2=59.25 //y2=1.375
r946 (  181 260 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.92 //y=0.755 //x2=58.805 //y2=0.755
r947 (  180 267 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.135 //y=0.755 //x2=59.25 //y2=0.755
r948 (  180 181 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=59.135 //y=0.755 //x2=58.92 //y2=0.755
r949 (  179 261 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.765 //y=1.22 //x2=58.805 //y2=1.375
r950 (  178 260 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.765 //y=0.91 //x2=58.805 //y2=0.755
r951 (  178 179 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=58.765 //y=0.91 //x2=58.765 //y2=1.22
r952 (  174 254 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=46.385 //y=4.79 //x2=46.25 //y2=4.79
r953 (  173 175 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=46.585 //y=4.79 //x2=46.66 //y2=4.865
r954 (  173 174 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=46.585 //y=4.79 //x2=46.385 //y2=4.79
r955 (  172 259 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=46.34 //y=1.915 //x2=46.265 //y2=2.08
r956 (  171 257 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=46.34 //y=1.45 //x2=46.3 //y2=1.375
r957 (  171 172 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=46.34 //y=1.45 //x2=46.34 //y2=1.915
r958 (  170 257 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.34 //y=1.22 //x2=46.3 //y2=1.375
r959 (  169 256 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.34 //y=0.91 //x2=46.3 //y2=0.755
r960 (  169 170 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=46.34 //y=0.91 //x2=46.34 //y2=1.22
r961 (  164 250 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.97 //y=1.375 //x2=45.855 //y2=1.375
r962 (  163 257 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.185 //y=1.375 //x2=46.3 //y2=1.375
r963 (  162 249 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.97 //y=0.755 //x2=45.855 //y2=0.755
r964 (  161 256 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.185 //y=0.755 //x2=46.3 //y2=0.755
r965 (  161 162 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=46.185 //y=0.755 //x2=45.97 //y2=0.755
r966 (  160 250 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.815 //y=1.22 //x2=45.855 //y2=1.375
r967 (  159 249 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.815 //y=0.91 //x2=45.855 //y2=0.755
r968 (  159 160 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=45.815 //y=0.91 //x2=45.815 //y2=1.22
r969 (  155 243 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=34.915 //y=4.79 //x2=34.78 //y2=4.79
r970 (  154 156 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=35.115 //y=4.79 //x2=35.19 //y2=4.865
r971 (  154 155 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=35.115 //y=4.79 //x2=34.915 //y2=4.79
r972 (  153 248 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=34.87 //y=1.915 //x2=34.795 //y2=2.08
r973 (  152 246 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=34.87 //y=1.45 //x2=34.83 //y2=1.375
r974 (  152 153 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=34.87 //y=1.45 //x2=34.87 //y2=1.915
r975 (  151 246 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.87 //y=1.22 //x2=34.83 //y2=1.375
r976 (  150 245 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.87 //y=0.91 //x2=34.83 //y2=0.755
r977 (  150 151 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=34.87 //y=0.91 //x2=34.87 //y2=1.22
r978 (  145 239 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.5 //y=1.375 //x2=34.385 //y2=1.375
r979 (  144 246 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.715 //y=1.375 //x2=34.83 //y2=1.375
r980 (  143 238 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.5 //y=0.755 //x2=34.385 //y2=0.755
r981 (  142 245 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.715 //y=0.755 //x2=34.83 //y2=0.755
r982 (  142 143 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=34.715 //y=0.755 //x2=34.5 //y2=0.755
r983 (  141 239 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.345 //y=1.22 //x2=34.385 //y2=1.375
r984 (  140 238 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.345 //y=0.91 //x2=34.385 //y2=0.755
r985 (  140 141 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=34.345 //y=0.91 //x2=34.345 //y2=1.22
r986 (  136 232 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=21.965 //y=4.79 //x2=21.83 //y2=4.79
r987 (  135 137 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=22.165 //y=4.79 //x2=22.24 //y2=4.865
r988 (  135 136 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=22.165 //y=4.79 //x2=21.965 //y2=4.79
r989 (  134 237 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.915 //x2=21.845 //y2=2.08
r990 (  133 235 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.45 //x2=21.88 //y2=1.375
r991 (  133 134 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.45 //x2=21.92 //y2=1.915
r992 (  132 235 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.22 //x2=21.88 //y2=1.375
r993 (  131 234 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.92 //y=0.91 //x2=21.88 //y2=0.755
r994 (  131 132 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.92 //y=0.91 //x2=21.92 //y2=1.22
r995 (  126 228 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.375 //x2=21.435 //y2=1.375
r996 (  125 235 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.765 //y=1.375 //x2=21.88 //y2=1.375
r997 (  124 227 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.755 //x2=21.435 //y2=0.755
r998 (  123 234 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.765 //y=0.755 //x2=21.88 //y2=0.755
r999 (  123 124 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=21.765 //y=0.755 //x2=21.55 //y2=0.755
r1000 (  122 228 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.395 //y=1.22 //x2=21.435 //y2=1.375
r1001 (  121 227 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.91 //x2=21.435 //y2=0.755
r1002 (  121 122 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.91 //x2=21.395 //y2=1.22
r1003 (  117 221 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=10.495 //y=4.79 //x2=10.36 //y2=4.79
r1004 (  116 118 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.695 //y=4.79 //x2=10.77 //y2=4.865
r1005 (  116 117 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=10.695 //y=4.79 //x2=10.495 //y2=4.79
r1006 (  115 226 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.915 //x2=10.375 //y2=2.08
r1007 (  114 224 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.45 //x2=10.41 //y2=1.375
r1008 (  114 115 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.45 //x2=10.45 //y2=1.915
r1009 (  113 224 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.22 //x2=10.41 //y2=1.375
r1010 (  112 223 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.45 //y=0.91 //x2=10.41 //y2=0.755
r1011 (  112 113 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=10.45 //y=0.91 //x2=10.45 //y2=1.22
r1012 (  107 217 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.08 //y=1.375 //x2=9.965 //y2=1.375
r1013 (  106 224 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.295 //y=1.375 //x2=10.41 //y2=1.375
r1014 (  105 216 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.08 //y=0.755 //x2=9.965 //y2=0.755
r1015 (  104 223 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.295 //y=0.755 //x2=10.41 //y2=0.755
r1016 (  104 105 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=10.295 //y=0.755 //x2=10.08 //y2=0.755
r1017 (  103 217 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.925 //y=1.22 //x2=9.965 //y2=1.375
r1018 (  102 216 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.925 //y=0.91 //x2=9.965 //y2=0.755
r1019 (  102 103 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=9.925 //y=0.91 //x2=9.925 //y2=1.22
r1020 (  101 213 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=71.08 //y=6.02 //x2=71.08 //y2=4.865
r1021 (  100 277 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.64 //y=6.02 //x2=70.64 //y2=4.865
r1022 (  99 194 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.61 //y=6.02 //x2=59.61 //y2=4.865
r1023 (  98 266 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.17 //y=6.02 //x2=59.17 //y2=4.865
r1024 (  97 175 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.66 //y=6.02 //x2=46.66 //y2=4.865
r1025 (  96 255 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.22 //y=6.02 //x2=46.22 //y2=4.865
r1026 (  95 156 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.19 //y=6.02 //x2=35.19 //y2=4.865
r1027 (  94 244 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.75 //y=6.02 //x2=34.75 //y2=4.865
r1028 (  93 137 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.24 //y=6.02 //x2=22.24 //y2=4.865
r1029 (  92 233 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.8 //y=6.02 //x2=21.8 //y2=4.865
r1030 (  91 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.77 //y=6.02 //x2=10.77 //y2=4.865
r1031 (  90 222 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.33 //y=6.02 //x2=10.33 //y2=4.865
r1032 (  89 201 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=70.497 //y=1.375 //x2=70.605 //y2=1.375
r1033 (  89 202 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=70.497 //y=1.375 //x2=70.39 //y2=1.375
r1034 (  88 182 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=59.027 //y=1.375 //x2=59.135 //y2=1.375
r1035 (  88 183 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=59.027 //y=1.375 //x2=58.92 //y2=1.375
r1036 (  87 163 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=46.077 //y=1.375 //x2=46.185 //y2=1.375
r1037 (  87 164 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=46.077 //y=1.375 //x2=45.97 //y2=1.375
r1038 (  86 144 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=34.607 //y=1.375 //x2=34.715 //y2=1.375
r1039 (  86 145 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=34.607 //y=1.375 //x2=34.5 //y2=1.375
r1040 (  85 125 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=21.657 //y=1.375 //x2=21.765 //y2=1.375
r1041 (  85 126 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=21.657 //y=1.375 //x2=21.55 //y2=1.375
r1042 (  84 106 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=10.187 //y=1.375 //x2=10.295 //y2=1.375
r1043 (  84 107 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=10.187 //y=1.375 //x2=10.08 //y2=1.375
r1044 (  82 274 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=4.7 //x2=70.67 //y2=4.7
r1045 (  77 281 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=2.08 //x2=70.67 //y2=2.08
r1046 (  74 263 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.2 //y=4.7 //x2=59.2 //y2=4.7
r1047 (  68 270 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.2 //y=2.08 //x2=59.2 //y2=2.08
r1048 (  65 252 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.25 //y=4.7 //x2=46.25 //y2=4.7
r1049 (  63 65 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=46.25 //y=2.22 //x2=46.25 //y2=4.7
r1050 (  60 259 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.25 //y=2.08 //x2=46.25 //y2=2.08
r1051 (  60 63 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=46.25 //y=2.08 //x2=46.25 //y2=2.22
r1052 (  57 241 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.78 //y=4.7 //x2=34.78 //y2=4.7
r1053 (  52 248 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.78 //y=2.08 //x2=34.78 //y2=2.08
r1054 (  49 230 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.83 //y=4.7 //x2=21.83 //y2=4.7
r1055 (  43 237 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.83 //y=2.08 //x2=21.83 //y2=2.08
r1056 (  40 219 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=4.7 //x2=10.36 //y2=4.7
r1057 (  33 226 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=2.08 //x2=10.36 //y2=2.08
r1058 (  31 82 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=70.67 //y=2.22 //x2=70.67 //y2=4.7
r1059 (  31 77 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=70.67 //y=2.22 //x2=70.67 //y2=2.08
r1060 (  30 74 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=59.2 //y=2.59 //x2=59.2 //y2=4.7
r1061 (  29 30 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=59.2 //y=2.22 //x2=59.2 //y2=2.59
r1062 (  29 68 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=59.2 //y=2.22 //x2=59.2 //y2=2.08
r1063 (  28 57 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=34.78 //y=2.22 //x2=34.78 //y2=4.7
r1064 (  28 52 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=34.78 //y=2.22 //x2=34.78 //y2=2.08
r1065 (  27 49 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.59 //x2=21.83 //y2=4.7
r1066 (  26 27 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.22 //x2=21.83 //y2=2.59
r1067 (  26 43 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.22 //x2=21.83 //y2=2.08
r1068 (  25 40 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=10.36 //y=3.33 //x2=10.36 //y2=4.7
r1069 (  24 25 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.59 //x2=10.36 //y2=3.33
r1070 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.22 //x2=10.36 //y2=2.59
r1071 (  23 33 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.22 //x2=10.36 //y2=2.08
r1072 (  22 31 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=70.67 //y=2.22 //x2=70.67 //y2=2.22
r1073 (  20 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=59.2 //y=2.22 //x2=59.2 //y2=2.22
r1074 (  18 63 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=46.25 //y=2.22 //x2=46.25 //y2=2.22
r1075 (  16 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=34.78 //y=2.22 //x2=34.78 //y2=2.22
r1076 (  14 26 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.83 //y=2.22 //x2=21.83 //y2=2.22
r1077 (  12 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=2.22 //x2=10.36 //y2=2.22
r1078 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=59.315 //y=2.22 //x2=59.2 //y2=2.22
r1079 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=2.22 //x2=70.67 //y2=2.22
r1080 (  9 10 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=2.22 //x2=59.315 //y2=2.22
r1081 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=46.365 //y=2.22 //x2=46.25 //y2=2.22
r1082 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=59.085 //y=2.22 //x2=59.2 //y2=2.22
r1083 (  7 8 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=59.085 //y=2.22 //x2=46.365 //y2=2.22
r1084 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.895 //y=2.22 //x2=34.78 //y2=2.22
r1085 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=46.135 //y=2.22 //x2=46.25 //y2=2.22
r1086 (  5 6 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=46.135 //y=2.22 //x2=34.895 //y2=2.22
r1087 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.945 //y=2.22 //x2=21.83 //y2=2.22
r1088 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=2.22 //x2=34.78 //y2=2.22
r1089 (  3 4 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=2.22 //x2=21.945 //y2=2.22
r1090 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.475 //y=2.22 //x2=10.36 //y2=2.22
r1091 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=2.22 //x2=21.83 //y2=2.22
r1092 (  1 2 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=2.22 //x2=10.475 //y2=2.22
ends PM_TMRDFFSNQNX1\%SN

subckt PM_TMRDFFSNQNX1\%noxref_19 ( 1 2 3 4 5 6 16 24 37 38 49 51 52 56 58 65 \
 66 67 68 69 70 71 72 73 74 78 79 80 85 87 90 91 95 96 97 102 104 107 108 112 \
 113 114 119 121 124 125 127 128 133 137 138 143 147 148 153 156 158 159 )
c321 ( 159 0 ) capacitor c=0.0220291f //x=63.755 //y=5.02
c322 ( 158 0 ) capacitor c=0.0217503f //x=62.875 //y=5.02
c323 ( 156 0 ) capacitor c=0.00866655f //x=63.75 //y=0.905
c324 ( 153 0 ) capacitor c=0.0587755f //x=71.78 //y=4.7
c325 ( 148 0 ) capacitor c=0.0273931f //x=71.78 //y=1.915
c326 ( 147 0 ) capacitor c=0.0458323f //x=71.78 //y=2.08
c327 ( 143 0 ) capacitor c=0.0587755f //x=60.31 //y=4.7
c328 ( 138 0 ) capacitor c=0.0273931f //x=60.31 //y=1.915
c329 ( 137 0 ) capacitor c=0.0456313f //x=60.31 //y=2.08
c330 ( 133 0 ) capacitor c=0.058931f //x=55.5 //y=4.7
c331 ( 128 0 ) capacitor c=0.0267105f //x=55.5 //y=1.915
c332 ( 127 0 ) capacitor c=0.0456313f //x=55.5 //y=2.08
c333 ( 125 0 ) capacitor c=0.0432517f //x=72.3 //y=1.26
c334 ( 124 0 ) capacitor c=0.0200379f //x=72.3 //y=0.915
c335 ( 121 0 ) capacitor c=0.0158629f //x=72.145 //y=1.415
c336 ( 119 0 ) capacitor c=0.0157803f //x=72.145 //y=0.76
c337 ( 114 0 ) capacitor c=0.0218028f //x=71.77 //y=1.57
c338 ( 113 0 ) capacitor c=0.0207459f //x=71.77 //y=1.26
c339 ( 112 0 ) capacitor c=0.0194308f //x=71.77 //y=0.915
c340 ( 108 0 ) capacitor c=0.0432517f //x=60.83 //y=1.26
c341 ( 107 0 ) capacitor c=0.0200379f //x=60.83 //y=0.915
c342 ( 104 0 ) capacitor c=0.0148873f //x=60.675 //y=1.415
c343 ( 102 0 ) capacitor c=0.0157803f //x=60.675 //y=0.76
c344 ( 97 0 ) capacitor c=0.0218028f //x=60.3 //y=1.57
c345 ( 96 0 ) capacitor c=0.0207459f //x=60.3 //y=1.26
c346 ( 95 0 ) capacitor c=0.0194308f //x=60.3 //y=0.915
c347 ( 91 0 ) capacitor c=0.0432517f //x=56.02 //y=1.26
c348 ( 90 0 ) capacitor c=0.0200379f //x=56.02 //y=0.915
c349 ( 87 0 ) capacitor c=0.0148873f //x=55.865 //y=1.415
c350 ( 85 0 ) capacitor c=0.0157803f //x=55.865 //y=0.76
c351 ( 80 0 ) capacitor c=0.0218028f //x=55.49 //y=1.57
c352 ( 79 0 ) capacitor c=0.0207459f //x=55.49 //y=1.26
c353 ( 78 0 ) capacitor c=0.0194308f //x=55.49 //y=0.915
c354 ( 74 0 ) capacitor c=0.158794f //x=71.96 //y=6.02
c355 ( 73 0 ) capacitor c=0.110114f //x=71.52 //y=6.02
c356 ( 72 0 ) capacitor c=0.158794f //x=60.49 //y=6.02
c357 ( 71 0 ) capacitor c=0.110114f //x=60.05 //y=6.02
c358 ( 70 0 ) capacitor c=0.158048f //x=55.68 //y=6.02
c359 ( 69 0 ) capacitor c=0.110114f //x=55.24 //y=6.02
c360 ( 65 0 ) capacitor c=0.0023043f //x=63.9 //y=5.2
c361 ( 58 0 ) capacitor c=0.0841207f //x=71.78 //y=2.08
c362 ( 56 0 ) capacitor c=0.10491f //x=64.38 //y=3.7
c363 ( 52 0 ) capacitor c=0.00404073f //x=64.025 //y=1.655
c364 ( 51 0 ) capacitor c=0.0122201f //x=64.295 //y=1.655
c365 ( 49 0 ) capacitor c=0.0140462f //x=64.295 //y=5.2
c366 ( 38 0 ) capacitor c=0.00251635f //x=63.105 //y=5.2
c367 ( 37 0 ) capacitor c=0.0143111f //x=63.815 //y=5.2
c368 ( 24 0 ) capacitor c=0.0811636f //x=60.31 //y=2.08
c369 ( 16 0 ) capacitor c=0.0796434f //x=55.5 //y=2.08
c370 ( 6 0 ) capacitor c=0.00405261f //x=64.495 //y=3.7
c371 ( 5 0 ) capacitor c=0.125528f //x=71.665 //y=3.7
c372 ( 4 0 ) capacitor c=0.00412452f //x=60.425 //y=3.7
c373 ( 3 0 ) capacitor c=0.0546427f //x=64.265 //y=3.7
c374 ( 2 0 ) capacitor c=0.0138772f //x=55.615 //y=3.7
c375 ( 1 0 ) capacitor c=0.0670382f //x=60.195 //y=3.7
r376 (  147 148 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=71.78 //y=2.08 //x2=71.78 //y2=1.915
r377 (  137 138 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=60.31 //y=2.08 //x2=60.31 //y2=1.915
r378 (  127 128 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=55.5 //y=2.08 //x2=55.5 //y2=1.915
r379 (  125 155 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.3 //y=1.26 //x2=72.26 //y2=1.415
r380 (  124 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.3 //y=0.915 //x2=72.26 //y2=0.76
r381 (  124 125 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=72.3 //y=0.915 //x2=72.3 //y2=1.26
r382 (  122 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.925 //y=1.415 //x2=71.81 //y2=1.415
r383 (  121 155 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=72.145 //y=1.415 //x2=72.26 //y2=1.415
r384 (  120 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.925 //y=0.76 //x2=71.81 //y2=0.76
r385 (  119 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=72.145 //y=0.76 //x2=72.26 //y2=0.76
r386 (  119 120 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=72.145 //y=0.76 //x2=71.925 //y2=0.76
r387 (  116 153 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=71.96 //y=4.865 //x2=71.78 //y2=4.7
r388 (  114 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.77 //y=1.57 //x2=71.81 //y2=1.415
r389 (  114 148 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=71.77 //y=1.57 //x2=71.77 //y2=1.915
r390 (  113 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.77 //y=1.26 //x2=71.81 //y2=1.415
r391 (  112 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.77 //y=0.915 //x2=71.81 //y2=0.76
r392 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=71.77 //y=0.915 //x2=71.77 //y2=1.26
r393 (  109 153 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=71.52 //y=4.865 //x2=71.78 //y2=4.7
r394 (  108 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.83 //y=1.26 //x2=60.79 //y2=1.415
r395 (  107 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.83 //y=0.915 //x2=60.79 //y2=0.76
r396 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=60.83 //y=0.915 //x2=60.83 //y2=1.26
r397 (  105 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.455 //y=1.415 //x2=60.34 //y2=1.415
r398 (  104 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.675 //y=1.415 //x2=60.79 //y2=1.415
r399 (  103 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.455 //y=0.76 //x2=60.34 //y2=0.76
r400 (  102 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.675 //y=0.76 //x2=60.79 //y2=0.76
r401 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=60.675 //y=0.76 //x2=60.455 //y2=0.76
r402 (  99 143 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=60.49 //y=4.865 //x2=60.31 //y2=4.7
r403 (  97 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.3 //y=1.57 //x2=60.34 //y2=1.415
r404 (  97 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=60.3 //y=1.57 //x2=60.3 //y2=1.915
r405 (  96 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.3 //y=1.26 //x2=60.34 //y2=1.415
r406 (  95 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.3 //y=0.915 //x2=60.34 //y2=0.76
r407 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=60.3 //y=0.915 //x2=60.3 //y2=1.26
r408 (  92 143 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=60.05 //y=4.865 //x2=60.31 //y2=4.7
r409 (  91 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.02 //y=1.26 //x2=55.98 //y2=1.415
r410 (  90 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.02 //y=0.915 //x2=55.98 //y2=0.76
r411 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.02 //y=0.915 //x2=56.02 //y2=1.26
r412 (  88 131 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.645 //y=1.415 //x2=55.53 //y2=1.415
r413 (  87 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.865 //y=1.415 //x2=55.98 //y2=1.415
r414 (  86 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.645 //y=0.76 //x2=55.53 //y2=0.76
r415 (  85 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.865 //y=0.76 //x2=55.98 //y2=0.76
r416 (  85 86 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=55.865 //y=0.76 //x2=55.645 //y2=0.76
r417 (  82 133 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=55.68 //y=4.865 //x2=55.5 //y2=4.7
r418 (  80 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.49 //y=1.57 //x2=55.53 //y2=1.415
r419 (  80 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=55.49 //y=1.57 //x2=55.49 //y2=1.915
r420 (  79 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.49 //y=1.26 //x2=55.53 //y2=1.415
r421 (  78 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.49 //y=0.915 //x2=55.53 //y2=0.76
r422 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=55.49 //y=0.915 //x2=55.49 //y2=1.26
r423 (  75 133 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=55.24 //y=4.865 //x2=55.5 //y2=4.7
r424 (  74 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=71.96 //y=6.02 //x2=71.96 //y2=4.865
r425 (  73 109 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=71.52 //y=6.02 //x2=71.52 //y2=4.865
r426 (  72 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.49 //y=6.02 //x2=60.49 //y2=4.865
r427 (  71 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.05 //y=6.02 //x2=60.05 //y2=4.865
r428 (  70 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.68 //y=6.02 //x2=55.68 //y2=4.865
r429 (  69 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.24 //y=6.02 //x2=55.24 //y2=4.865
r430 (  68 121 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=72.035 //y=1.415 //x2=72.145 //y2=1.415
r431 (  68 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=72.035 //y=1.415 //x2=71.925 //y2=1.415
r432 (  67 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=60.565 //y=1.415 //x2=60.675 //y2=1.415
r433 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=60.565 //y=1.415 //x2=60.455 //y2=1.415
r434 (  66 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=55.755 //y=1.415 //x2=55.865 //y2=1.415
r435 (  66 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=55.755 //y=1.415 //x2=55.645 //y2=1.415
r436 (  63 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=71.78 //y=4.7 //x2=71.78 //y2=4.7
r437 (  61 63 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=71.78 //y=3.7 //x2=71.78 //y2=4.7
r438 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=71.78 //y=2.08 //x2=71.78 //y2=2.08
r439 (  58 61 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=71.78 //y=2.08 //x2=71.78 //y2=3.7
r440 (  54 56 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=64.38 //y=5.115 //x2=64.38 //y2=3.7
r441 (  53 56 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=64.38 //y=1.74 //x2=64.38 //y2=3.7
r442 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=64.295 //y=1.655 //x2=64.38 //y2=1.74
r443 (  51 52 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=64.295 //y=1.655 //x2=64.025 //y2=1.655
r444 (  50 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.985 //y=5.2 //x2=63.9 //y2=5.2
r445 (  49 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=64.295 //y=5.2 //x2=64.38 //y2=5.115
r446 (  49 50 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=64.295 //y=5.2 //x2=63.985 //y2=5.2
r447 (  45 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.94 //y=1.57 //x2=64.025 //y2=1.655
r448 (  45 156 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=63.94 //y=1.57 //x2=63.94 //y2=1
r449 (  39 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.9 //y=5.285 //x2=63.9 //y2=5.2
r450 (  39 159 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=63.9 //y=5.285 //x2=63.9 //y2=5.725
r451 (  37 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.815 //y=5.2 //x2=63.9 //y2=5.2
r452 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=63.815 //y=5.2 //x2=63.105 //y2=5.2
r453 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.02 //y=5.285 //x2=63.105 //y2=5.2
r454 (  31 158 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=63.02 //y=5.285 //x2=63.02 //y2=5.725
r455 (  29 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=60.31 //y=4.7 //x2=60.31 //y2=4.7
r456 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=60.31 //y=3.7 //x2=60.31 //y2=4.7
r457 (  24 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=60.31 //y=2.08 //x2=60.31 //y2=2.08
r458 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=60.31 //y=2.08 //x2=60.31 //y2=3.7
r459 (  21 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.5 //y=4.7 //x2=55.5 //y2=4.7
r460 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=55.5 //y=3.7 //x2=55.5 //y2=4.7
r461 (  16 127 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.5 //y=2.08 //x2=55.5 //y2=2.08
r462 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=55.5 //y=2.08 //x2=55.5 //y2=3.7
r463 (  14 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=71.78 //y=3.7 //x2=71.78 //y2=3.7
r464 (  12 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=64.38 //y=3.7 //x2=64.38 //y2=3.7
r465 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=60.31 //y=3.7 //x2=60.31 //y2=3.7
r466 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=55.5 //y=3.7 //x2=55.5 //y2=3.7
r467 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=64.495 //y=3.7 //x2=64.38 //y2=3.7
r468 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=71.665 //y=3.7 //x2=71.78 //y2=3.7
r469 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=71.665 //y=3.7 //x2=64.495 //y2=3.7
r470 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.425 //y=3.7 //x2=60.31 //y2=3.7
r471 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=64.265 //y=3.7 //x2=64.38 //y2=3.7
r472 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=64.265 //y=3.7 //x2=60.425 //y2=3.7
r473 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.615 //y=3.7 //x2=55.5 //y2=3.7
r474 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.195 //y=3.7 //x2=60.31 //y2=3.7
r475 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=60.195 //y=3.7 //x2=55.615 //y2=3.7
ends PM_TMRDFFSNQNX1\%noxref_19

subckt PM_TMRDFFSNQNX1\%noxref_20 ( 1 2 7 9 19 20 27 35 41 42 46 49 50 51 52 \
 53 54 55 56 61 63 65 71 72 74 75 78 86 88 89 90 )
c183 ( 90 0 ) capacitor c=0.023087f //x=71.595 //y=5.02
c184 ( 89 0 ) capacitor c=0.023519f //x=70.715 //y=5.02
c185 ( 88 0 ) capacitor c=0.0224735f //x=69.835 //y=5.02
c186 ( 86 0 ) capacitor c=0.0087111f //x=71.845 //y=0.915
c187 ( 78 0 ) capacitor c=0.0331534f //x=67 //y=4.7
c188 ( 75 0 ) capacitor c=0.0279499f //x=66.97 //y=1.915
c189 ( 74 0 ) capacitor c=0.0421676f //x=66.97 //y=2.08
c190 ( 72 0 ) capacitor c=0.0429696f //x=67.535 //y=1.25
c191 ( 71 0 ) capacitor c=0.0192208f //x=67.535 //y=0.905
c192 ( 65 0 ) capacitor c=0.0148884f //x=67.38 //y=1.405
c193 ( 63 0 ) capacitor c=0.0157803f //x=67.38 //y=0.75
c194 ( 61 0 ) capacitor c=0.0299681f //x=67.375 //y=4.79
c195 ( 56 0 ) capacitor c=0.0205163f //x=67.005 //y=1.56
c196 ( 55 0 ) capacitor c=0.0168481f //x=67.005 //y=1.25
c197 ( 54 0 ) capacitor c=0.0174783f //x=67.005 //y=0.905
c198 ( 53 0 ) capacitor c=0.15358f //x=67.45 //y=6.02
c199 ( 52 0 ) capacitor c=0.110281f //x=67.01 //y=6.02
c200 ( 50 0 ) capacitor c=0.00106608f //x=71.74 //y=5.155
c201 ( 49 0 ) capacitor c=0.00207319f //x=70.86 //y=5.155
c202 ( 46 0 ) capacitor c=0.106476f //x=72.52 //y=4.07
c203 ( 42 0 ) capacitor c=0.00463522f //x=72.12 //y=1.665
c204 ( 41 0 ) capacitor c=0.0148737f //x=72.435 //y=1.665
c205 ( 35 0 ) capacitor c=0.0281866f //x=72.435 //y=5.155
c206 ( 27 0 ) capacitor c=0.0176454f //x=71.655 //y=5.155
c207 ( 20 0 ) capacitor c=0.00332903f //x=70.065 //y=5.155
c208 ( 19 0 ) capacitor c=0.0148427f //x=70.775 //y=5.155
c209 ( 9 0 ) capacitor c=0.070954f //x=66.97 //y=2.08
c210 ( 7 0 ) capacitor c=0.00453889f //x=66.97 //y=4.535
c211 ( 2 0 ) capacitor c=0.00822824f //x=67.085 //y=4.07
c212 ( 1 0 ) capacitor c=0.0897196f //x=72.405 //y=4.07
r213 (  80 81 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=67 //y=4.79 //x2=67 //y2=4.865
r214 (  78 80 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=67 //y=4.7 //x2=67 //y2=4.79
r215 (  74 75 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=66.97 //y=2.08 //x2=66.97 //y2=1.915
r216 (  72 85 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.535 //y=1.25 //x2=67.495 //y2=1.405
r217 (  71 84 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.535 //y=0.905 //x2=67.495 //y2=0.75
r218 (  71 72 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=67.535 //y=0.905 //x2=67.535 //y2=1.25
r219 (  66 83 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=67.16 //y=1.405 //x2=67.045 //y2=1.405
r220 (  65 85 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=67.38 //y=1.405 //x2=67.495 //y2=1.405
r221 (  64 82 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=67.16 //y=0.75 //x2=67.045 //y2=0.75
r222 (  63 84 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=67.38 //y=0.75 //x2=67.495 //y2=0.75
r223 (  63 64 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=67.38 //y=0.75 //x2=67.16 //y2=0.75
r224 (  62 80 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=67.135 //y=4.79 //x2=67 //y2=4.79
r225 (  61 68 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=67.375 //y=4.79 //x2=67.45 //y2=4.865
r226 (  61 62 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=67.375 //y=4.79 //x2=67.135 //y2=4.79
r227 (  56 83 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.005 //y=1.56 //x2=67.045 //y2=1.405
r228 (  56 75 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=67.005 //y=1.56 //x2=67.005 //y2=1.915
r229 (  55 83 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.005 //y=1.25 //x2=67.045 //y2=1.405
r230 (  54 82 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.005 //y=0.905 //x2=67.045 //y2=0.75
r231 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=67.005 //y=0.905 //x2=67.005 //y2=1.25
r232 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=67.45 //y=6.02 //x2=67.45 //y2=4.865
r233 (  52 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=67.01 //y=6.02 //x2=67.01 //y2=4.865
r234 (  51 65 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=67.27 //y=1.405 //x2=67.38 //y2=1.405
r235 (  51 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=67.27 //y=1.405 //x2=67.16 //y2=1.405
r236 (  48 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=67 //y=4.7 //x2=67 //y2=4.7
r237 (  44 46 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=72.52 //y=5.07 //x2=72.52 //y2=4.07
r238 (  43 46 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=72.52 //y=1.75 //x2=72.52 //y2=4.07
r239 (  41 43 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=72.435 //y=1.665 //x2=72.52 //y2=1.75
r240 (  41 42 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=72.435 //y=1.665 //x2=72.12 //y2=1.665
r241 (  37 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=72.035 //y=1.58 //x2=72.12 //y2=1.665
r242 (  37 86 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=72.035 //y=1.58 //x2=72.035 //y2=1.01
r243 (  36 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.825 //y=5.155 //x2=71.74 //y2=5.155
r244 (  35 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=72.435 //y=5.155 //x2=72.52 //y2=5.07
r245 (  35 36 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=72.435 //y=5.155 //x2=71.825 //y2=5.155
r246 (  29 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.74 //y=5.24 //x2=71.74 //y2=5.155
r247 (  29 90 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=71.74 //y=5.24 //x2=71.74 //y2=5.725
r248 (  28 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.945 //y=5.155 //x2=70.86 //y2=5.155
r249 (  27 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.655 //y=5.155 //x2=71.74 //y2=5.155
r250 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=71.655 //y=5.155 //x2=70.945 //y2=5.155
r251 (  21 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.86 //y=5.24 //x2=70.86 //y2=5.155
r252 (  21 89 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=70.86 //y=5.24 //x2=70.86 //y2=5.725
r253 (  19 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.775 //y=5.155 //x2=70.86 //y2=5.155
r254 (  19 20 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=70.775 //y=5.155 //x2=70.065 //y2=5.155
r255 (  13 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=69.98 //y=5.24 //x2=70.065 //y2=5.155
r256 (  13 88 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=69.98 //y=5.24 //x2=69.98 //y2=5.725
r257 (  9 74 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.97 //y=2.08 //x2=66.97 //y2=2.08
r258 (  9 12 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=66.97 //y=2.08 //x2=66.97 //y2=4.07
r259 (  7 48 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=66.97 //y=4.535 //x2=66.985 //y2=4.7
r260 (  7 12 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=66.97 //y=4.535 //x2=66.97 //y2=4.07
r261 (  6 46 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=72.52 //y=4.07 //x2=72.52 //y2=4.07
r262 (  4 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.97 //y=4.07 //x2=66.97 //y2=4.07
r263 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=67.085 //y=4.07 //x2=66.97 //y2=4.07
r264 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=72.405 //y=4.07 //x2=72.52 //y2=4.07
r265 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=72.405 //y=4.07 //x2=67.085 //y2=4.07
ends PM_TMRDFFSNQNX1\%noxref_20

subckt PM_TMRDFFSNQNX1\%noxref_21 ( 1 2 3 4 6 7 8 9 10 27 28 39 41 42 46 48 55 \
 57 65 69 73 76 77 78 79 80 81 82 83 84 85 86 87 88 89 91 97 98 99 100 104 105 \
 106 111 113 115 121 122 123 124 125 130 132 134 140 141 151 152 155 163 164 \
 167 175 177 178 )
c438 ( 178 0 ) capacitor c=0.0220291f //x=42.665 //y=5.02
c439 ( 177 0 ) capacitor c=0.0217503f //x=41.785 //y=5.02
c440 ( 175 0 ) capacitor c=0.0084702f //x=42.66 //y=0.905
c441 ( 167 0 ) capacitor c=0.0352016f //x=81.79 //y=4.705
c442 ( 164 0 ) capacitor c=0.0279733f //x=81.77 //y=1.915
c443 ( 163 0 ) capacitor c=0.0467621f //x=81.77 //y=2.08
c444 ( 155 0 ) capacitor c=0.03845f //x=75.15 //y=4.705
c445 ( 152 0 ) capacitor c=0.0300885f //x=75.11 //y=1.915
c446 ( 151 0 ) capacitor c=0.0520257f //x=75.11 //y=2.08
c447 ( 141 0 ) capacitor c=0.0237734f //x=82.335 //y=1.255
c448 ( 140 0 ) capacitor c=0.0191782f //x=82.335 //y=0.905
c449 ( 134 0 ) capacitor c=0.0351663f //x=82.18 //y=1.405
c450 ( 132 0 ) capacitor c=0.0157803f //x=82.18 //y=0.75
c451 ( 130 0 ) capacitor c=0.0373879f //x=82.175 //y=4.795
c452 ( 125 0 ) capacitor c=0.0200628f //x=81.805 //y=1.56
c453 ( 124 0 ) capacitor c=0.0168575f //x=81.805 //y=1.255
c454 ( 123 0 ) capacitor c=0.0174993f //x=81.805 //y=0.905
c455 ( 122 0 ) capacitor c=0.0447087f //x=75.675 //y=1.25
c456 ( 121 0 ) capacitor c=0.019286f //x=75.675 //y=0.905
c457 ( 115 0 ) capacitor c=0.0187932f //x=75.52 //y=1.405
c458 ( 113 0 ) capacitor c=0.0157795f //x=75.52 //y=0.75
c459 ( 111 0 ) capacitor c=0.029531f //x=75.515 //y=4.795
c460 ( 106 0 ) capacitor c=0.0206178f //x=75.145 //y=1.56
c461 ( 105 0 ) capacitor c=0.016848f //x=75.145 //y=1.25
c462 ( 104 0 ) capacitor c=0.0174777f //x=75.145 //y=0.905
c463 ( 100 0 ) capacitor c=0.0556143f //x=45.415 //y=4.79
c464 ( 99 0 ) capacitor c=0.0293157f //x=45.705 //y=4.79
c465 ( 98 0 ) capacitor c=0.0347816f //x=45.37 //y=1.22
c466 ( 97 0 ) capacitor c=0.0187487f //x=45.37 //y=0.875
c467 ( 91 0 ) capacitor c=0.0137055f //x=45.215 //y=1.375
c468 ( 89 0 ) capacitor c=0.0149861f //x=45.215 //y=0.72
c469 ( 88 0 ) capacitor c=0.096037f //x=44.84 //y=1.915
c470 ( 87 0 ) capacitor c=0.0228993f //x=44.84 //y=1.53
c471 ( 86 0 ) capacitor c=0.0234352f //x=44.84 //y=1.22
c472 ( 85 0 ) capacitor c=0.0198724f //x=44.84 //y=0.875
c473 ( 84 0 ) capacitor c=0.15325f //x=82.25 //y=6.025
c474 ( 83 0 ) capacitor c=0.110411f //x=81.81 //y=6.025
c475 ( 82 0 ) capacitor c=0.154236f //x=75.59 //y=6.025
c476 ( 81 0 ) capacitor c=0.110294f //x=75.15 //y=6.025
c477 ( 80 0 ) capacitor c=0.110114f //x=45.78 //y=6.02
c478 ( 79 0 ) capacitor c=0.158956f //x=45.34 //y=6.02
c479 ( 73 0 ) capacitor c=0.00501304f //x=81.79 //y=4.705
c480 ( 69 0 ) capacitor c=0.00211606f //x=42.81 //y=5.2
c481 ( 65 0 ) capacitor c=0.0899745f //x=81.77 //y=2.08
c482 ( 57 0 ) capacitor c=0.105317f //x=75.11 //y=2.08
c483 ( 55 0 ) capacitor c=0.00669947f //x=75.11 //y=4.54
c484 ( 48 0 ) capacitor c=0.0938724f //x=45.14 //y=2.08
c485 ( 46 0 ) capacitor c=0.10219f //x=43.29 //y=2.59
c486 ( 42 0 ) capacitor c=0.00404073f //x=42.935 //y=1.655
c487 ( 41 0 ) capacitor c=0.0122201f //x=43.205 //y=1.655
c488 ( 39 0 ) capacitor c=0.0137995f //x=43.205 //y=5.2
c489 ( 28 0 ) capacitor c=0.00251459f //x=42.015 //y=5.2
c490 ( 27 0 ) capacitor c=0.0143649f //x=42.725 //y=5.2
c491 ( 10 0 ) capacitor c=0.0100708f //x=75.225 //y=4.07
c492 ( 9 0 ) capacitor c=0.189034f //x=81.655 //y=4.07
c493 ( 8 0 ) capacitor c=1.21334e-19 //x=50.775 //y=2.96
c494 ( 7 0 ) capacitor c=0.431449f //x=74.995 //y=2.96
c495 ( 4 0 ) capacitor c=0.00409365f //x=45.255 //y=2.59
c496 ( 3 0 ) capacitor c=0.0720829f //x=50.605 //y=2.59
c497 ( 2 0 ) capacitor c=0.0120208f //x=43.405 //y=2.59
c498 ( 1 0 ) capacitor c=0.0233304f //x=45.025 //y=2.59
r499 (  169 170 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=81.79 //y=4.795 //x2=81.79 //y2=4.87
r500 (  167 169 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=81.79 //y=4.705 //x2=81.79 //y2=4.795
r501 (  163 164 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=81.77 //y=2.08 //x2=81.77 //y2=1.915
r502 (  155 157 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=75.15 //y=4.705 //x2=75.15 //y2=4.795
r503 (  151 152 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=75.11 //y=2.08 //x2=75.11 //y2=1.915
r504 (  141 174 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=82.335 //y=1.255 //x2=82.335 //y2=1.367
r505 (  140 173 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.335 //y=0.905 //x2=82.295 //y2=0.75
r506 (  140 141 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=82.335 //y=0.905 //x2=82.335 //y2=1.255
r507 (  135 172 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=81.96 //y=1.405 //x2=81.845 //y2=1.405
r508 (  134 174 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=82.18 //y=1.405 //x2=82.335 //y2=1.367
r509 (  133 171 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=81.96 //y=0.75 //x2=81.845 //y2=0.75
r510 (  132 173 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.18 //y=0.75 //x2=82.295 //y2=0.75
r511 (  132 133 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=82.18 //y=0.75 //x2=81.96 //y2=0.75
r512 (  131 169 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=81.925 //y=4.795 //x2=81.79 //y2=4.795
r513 (  130 137 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=82.175 //y=4.795 //x2=82.25 //y2=4.87
r514 (  130 131 ) resistor r=128.191 //w=0.094 //l=0.25 //layer=ply \
 //thickness=0.18 //x=82.175 //y=4.795 //x2=81.925 //y2=4.795
r515 (  125 172 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.805 //y=1.56 //x2=81.845 //y2=1.405
r516 (  125 164 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=81.805 //y=1.56 //x2=81.805 //y2=1.915
r517 (  124 172 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=81.805 //y=1.255 //x2=81.845 //y2=1.405
r518 (  123 171 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.805 //y=0.905 //x2=81.845 //y2=0.75
r519 (  123 124 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=81.805 //y=0.905 //x2=81.805 //y2=1.255
r520 (  122 161 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.675 //y=1.25 //x2=75.635 //y2=1.405
r521 (  121 160 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.675 //y=0.905 //x2=75.635 //y2=0.75
r522 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.675 //y=0.905 //x2=75.675 //y2=1.25
r523 (  116 159 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.3 //y=1.405 //x2=75.185 //y2=1.405
r524 (  115 161 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.52 //y=1.405 //x2=75.635 //y2=1.405
r525 (  114 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.3 //y=0.75 //x2=75.185 //y2=0.75
r526 (  113 160 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.52 //y=0.75 //x2=75.635 //y2=0.75
r527 (  113 114 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=75.52 //y=0.75 //x2=75.3 //y2=0.75
r528 (  112 157 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=75.285 //y=4.795 //x2=75.15 //y2=4.795
r529 (  111 118 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=75.515 //y=4.795 //x2=75.59 //y2=4.87
r530 (  111 112 ) resistor r=117.936 //w=0.094 //l=0.23 //layer=ply \
 //thickness=0.18 //x=75.515 //y=4.795 //x2=75.285 //y2=4.795
r531 (  108 157 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=75.15 //y=4.87 //x2=75.15 //y2=4.795
r532 (  106 159 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.145 //y=1.56 //x2=75.185 //y2=1.405
r533 (  106 152 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=75.145 //y=1.56 //x2=75.145 //y2=1.915
r534 (  105 159 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.145 //y=1.25 //x2=75.185 //y2=1.405
r535 (  104 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.145 //y=0.905 //x2=75.185 //y2=0.75
r536 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.145 //y=0.905 //x2=75.145 //y2=1.25
r537 (  99 101 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=45.705 //y=4.79 //x2=45.78 //y2=4.865
r538 (  99 100 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=45.705 //y=4.79 //x2=45.415 //y2=4.79
r539 (  98 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.37 //y=1.22 //x2=45.33 //y2=1.375
r540 (  97 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.37 //y=0.875 //x2=45.33 //y2=0.72
r541 (  97 98 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=45.37 //y=0.875 //x2=45.37 //y2=1.22
r542 (  94 100 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=45.34 //y=4.865 //x2=45.415 //y2=4.79
r543 (  94 147 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=45.34 //y=4.865 //x2=45.14 //y2=4.7
r544 (  92 143 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.995 //y=1.375 //x2=44.88 //y2=1.375
r545 (  91 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.215 //y=1.375 //x2=45.33 //y2=1.375
r546 (  90 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.995 //y=0.72 //x2=44.88 //y2=0.72
r547 (  89 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.215 //y=0.72 //x2=45.33 //y2=0.72
r548 (  89 90 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=45.215 //y=0.72 //x2=44.995 //y2=0.72
r549 (  88 145 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=44.84 //y=1.915 //x2=45.14 //y2=2.08
r550 (  87 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.84 //y=1.53 //x2=44.88 //y2=1.375
r551 (  87 88 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=44.84 //y=1.53 //x2=44.84 //y2=1.915
r552 (  86 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.84 //y=1.22 //x2=44.88 //y2=1.375
r553 (  85 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.84 //y=0.875 //x2=44.88 //y2=0.72
r554 (  85 86 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=44.84 //y=0.875 //x2=44.84 //y2=1.22
r555 (  84 137 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=82.25 //y=6.025 //x2=82.25 //y2=4.87
r556 (  83 170 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=81.81 //y=6.025 //x2=81.81 //y2=4.87
r557 (  82 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.59 //y=6.025 //x2=75.59 //y2=4.87
r558 (  81 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.15 //y=6.025 //x2=75.15 //y2=4.87
r559 (  80 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.78 //y=6.02 //x2=45.78 //y2=4.865
r560 (  79 94 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.34 //y=6.02 //x2=45.34 //y2=4.865
r561 (  78 134 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.07 //y=1.405 //x2=82.18 //y2=1.405
r562 (  78 135 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.07 //y=1.405 //x2=81.96 //y2=1.405
r563 (  77 115 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.41 //y=1.405 //x2=75.52 //y2=1.405
r564 (  77 116 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.41 //y=1.405 //x2=75.3 //y2=1.405
r565 (  76 91 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=45.105 //y=1.375 //x2=45.215 //y2=1.375
r566 (  76 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=45.105 //y=1.375 //x2=44.995 //y2=1.375
r567 (  73 167 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=81.79 //y=4.705 //x2=81.79 //y2=4.705
r568 (  73 74 ) resistor r=10.3507 //w=0.207 //l=0.165 //layer=li \
 //thickness=0.1 //x=81.78 //y=4.705 //x2=81.78 //y2=4.54
r569 (  71 155 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.15 //y=4.705 //x2=75.15 //y2=4.705
r570 (  68 74 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=81.77 //y=4.07 //x2=81.77 //y2=4.54
r571 (  65 163 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=81.77 //y=2.08 //x2=81.77 //y2=2.08
r572 (  65 68 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=81.77 //y=2.08 //x2=81.77 //y2=4.07
r573 (  60 62 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=75.11 //y=2.96 //x2=75.11 //y2=4.07
r574 (  57 151 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.11 //y=2.08 //x2=75.11 //y2=2.08
r575 (  57 60 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=75.11 //y=2.08 //x2=75.11 //y2=2.96
r576 (  55 71 ) resistor r=11.2426 //w=0.191 //l=0.174714 //layer=li \
 //thickness=0.1 //x=75.11 //y=4.54 //x2=75.13 //y2=4.705
r577 (  55 62 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=75.11 //y=4.54 //x2=75.11 //y2=4.07
r578 (  53 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.14 //y=4.7 //x2=45.14 //y2=4.7
r579 (  51 53 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=45.14 //y=2.59 //x2=45.14 //y2=4.7
r580 (  48 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.14 //y=2.08 //x2=45.14 //y2=2.08
r581 (  48 51 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=45.14 //y=2.08 //x2=45.14 //y2=2.59
r582 (  44 46 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=43.29 //y=5.115 //x2=43.29 //y2=2.59
r583 (  43 46 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=43.29 //y=1.74 //x2=43.29 //y2=2.59
r584 (  41 43 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=43.205 //y=1.655 //x2=43.29 //y2=1.74
r585 (  41 42 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=43.205 //y=1.655 //x2=42.935 //y2=1.655
r586 (  40 69 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.895 //y=5.2 //x2=42.81 //y2=5.2
r587 (  39 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=43.205 //y=5.2 //x2=43.29 //y2=5.115
r588 (  39 40 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=43.205 //y=5.2 //x2=42.895 //y2=5.2
r589 (  35 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.85 //y=1.57 //x2=42.935 //y2=1.655
r590 (  35 175 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=42.85 //y=1.57 //x2=42.85 //y2=1
r591 (  29 69 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.81 //y=5.285 //x2=42.81 //y2=5.2
r592 (  29 178 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=42.81 //y=5.285 //x2=42.81 //y2=5.725
r593 (  27 69 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.725 //y=5.2 //x2=42.81 //y2=5.2
r594 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=42.725 //y=5.2 //x2=42.015 //y2=5.2
r595 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=41.93 //y=5.285 //x2=42.015 //y2=5.2
r596 (  21 177 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=41.93 //y=5.285 //x2=41.93 //y2=5.725
r597 (  20 68 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=81.77 //y=4.07 //x2=81.77 //y2=4.07
r598 (  18 60 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.11 //y=2.96 //x2=75.11 //y2=2.96
r599 (  16 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.11 //y=4.07 //x2=75.11 //y2=4.07
r600 (  14 51 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=45.14 //y=2.59 //x2=45.14 //y2=2.59
r601 (  12 46 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=43.29 //y=2.59 //x2=43.29 //y2=2.59
r602 (  10 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.225 //y=4.07 //x2=75.11 //y2=4.07
r603 (  9 20 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=81.655 //y=4.07 //x2=81.77 //y2=4.07
r604 (  9 10 ) resistor r=6.1355 //w=0.131 //l=6.43 //layer=m1 \
 //thickness=0.36 //x=81.655 //y=4.07 //x2=75.225 //y2=4.07
r605 (  7 18 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=74.995 //y=2.96 //x2=75.11 //y2=2.96
r606 (  7 8 ) resistor r=23.1107 //w=0.131 //l=24.22 //layer=m1 \
 //thickness=0.36 //x=74.995 //y=2.96 //x2=50.775 //y2=2.96
r607 (  6 8 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=50.69 //y=2.875 //x2=50.775 //y2=2.96
r608 (  5 6 ) resistor r=0.19084 //w=0.131 //l=0.2 //layer=m1 //thickness=0.36 \
 //x=50.69 //y=2.675 //x2=50.69 //y2=2.875
r609 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.255 //y=2.59 //x2=45.14 //y2=2.59
r610 (  3 5 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=50.605 //y=2.59 //x2=50.69 //y2=2.675
r611 (  3 4 ) resistor r=5.10496 //w=0.131 //l=5.35 //layer=m1 \
 //thickness=0.36 //x=50.605 //y=2.59 //x2=45.255 //y2=2.59
r612 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=43.405 //y=2.59 //x2=43.29 //y2=2.59
r613 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.025 //y=2.59 //x2=45.14 //y2=2.59
r614 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=45.025 //y=2.59 //x2=43.405 //y2=2.59
ends PM_TMRDFFSNQNX1\%noxref_21

subckt PM_TMRDFFSNQNX1\%noxref_22 ( 1 2 13 14 15 23 29 30 37 50 51 52 53 54 )
c91 ( 54 0 ) capacitor c=0.034295f //x=78.985 //y=5.025
c92 ( 53 0 ) capacitor c=0.0174957f //x=78.105 //y=5.025
c93 ( 51 0 ) capacitor c=0.0214849f //x=75.225 //y=5.025
c94 ( 50 0 ) capacitor c=0.0217161f //x=74.345 //y=5.025
c95 ( 49 0 ) capacitor c=0.00115294f //x=78.25 //y=6.91
c96 ( 37 0 ) capacitor c=0.0131238f //x=79.045 //y=6.91
c97 ( 30 0 ) capacitor c=0.00386507f //x=77.455 //y=6.91
c98 ( 29 0 ) capacitor c=0.00951687f //x=78.165 //y=6.91
c99 ( 23 0 ) capacitor c=0.0455351f //x=77.37 //y=5.21
c100 ( 15 0 ) capacitor c=0.00871244f //x=75.37 //y=5.295
c101 ( 14 0 ) capacitor c=0.00290434f //x=74.575 //y=5.21
c102 ( 13 0 ) capacitor c=0.0139202f //x=75.285 //y=5.21
c103 ( 2 0 ) capacitor c=0.0091252f //x=75.485 //y=5.21
c104 ( 1 0 ) capacitor c=0.0484159f //x=77.255 //y=5.21
r105 (  39 54 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.13 //y=6.825 //x2=79.13 //y2=6.74
r106 (  38 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.335 //y=6.91 //x2=78.25 //y2=6.91
r107 (  37 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=79.045 //y=6.91 //x2=79.13 //y2=6.825
r108 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=79.045 //y=6.91 //x2=78.335 //y2=6.91
r109 (  31 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.25 //y=6.825 //x2=78.25 //y2=6.91
r110 (  31 53 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.25 //y=6.825 //x2=78.25 //y2=6.74
r111 (  29 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.165 //y=6.91 //x2=78.25 //y2=6.91
r112 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=78.165 //y=6.91 //x2=77.455 //y2=6.91
r113 (  23 52 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=77.37 //y=5.21 //x2=77.37 //y2=6.06
r114 (  21 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=77.37 //y=6.825 //x2=77.455 //y2=6.91
r115 (  21 52 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.37 //y=6.825 //x2=77.37 //y2=6.74
r116 (  15 48 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=75.37 //y=5.295 //x2=75.37 //y2=5.17
r117 (  15 51 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=75.37 //y=5.295 //x2=75.37 //y2=6.06
r118 (  13 48 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.285 //y=5.21 //x2=75.37 //y2=5.17
r119 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=75.285 //y=5.21 //x2=74.575 //y2=5.21
r120 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=74.49 //y=5.295 //x2=74.575 //y2=5.21
r121 (  7 50 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=74.49 //y=5.295 //x2=74.49 //y2=5.72
r122 (  6 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=77.37 //y=5.21 //x2=77.37 //y2=5.21
r123 (  4 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.37 //y=5.21 //x2=75.37 //y2=5.21
r124 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.485 //y=5.21 //x2=75.37 //y2=5.21
r125 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=77.255 //y=5.21 //x2=77.37 //y2=5.21
r126 (  1 2 ) resistor r=1.68893 //w=0.131 //l=1.77 //layer=m1 \
 //thickness=0.36 //x=77.255 //y=5.21 //x2=75.485 //y2=5.21
ends PM_TMRDFFSNQNX1\%noxref_22

subckt PM_TMRDFFSNQNX1\%noxref_23 ( 1 2 3 4 5 6 21 22 33 35 36 40 42 50 58 65 \
 66 67 68 69 70 71 72 73 74 75 76 77 78 79 81 87 88 89 90 94 95 96 97 101 103 \
 106 107 108 109 113 114 115 116 120 122 128 129 139 152 155 157 158 )
c349 ( 158 0 ) capacitor c=0.0220291f //x=67.085 //y=5.02
c350 ( 157 0 ) capacitor c=0.0217503f //x=66.205 //y=5.02
c351 ( 155 0 ) capacitor c=0.0084702f //x=67.08 //y=0.905
c352 ( 152 0 ) capacitor c=0.0655948f //x=77.7 //y=4.705
c353 ( 139 0 ) capacitor c=0.0545009f //x=74 //y=2.08
c354 ( 129 0 ) capacitor c=0.0342409f //x=78.035 //y=1.21
c355 ( 128 0 ) capacitor c=0.0187384f //x=78.035 //y=0.865
c356 ( 122 0 ) capacitor c=0.0141797f //x=77.88 //y=1.365
c357 ( 120 0 ) capacitor c=0.0149844f //x=77.88 //y=0.71
c358 ( 116 0 ) capacitor c=0.10193f //x=77.505 //y=1.915
c359 ( 115 0 ) capacitor c=0.0225105f //x=77.505 //y=1.52
c360 ( 114 0 ) capacitor c=0.0234376f //x=77.505 //y=1.21
c361 ( 113 0 ) capacitor c=0.0199343f //x=77.505 //y=0.865
c362 ( 109 0 ) capacitor c=0.0318948f //x=74.705 //y=1.21
c363 ( 108 0 ) capacitor c=0.0187384f //x=74.705 //y=0.865
c364 ( 107 0 ) capacitor c=0.0607141f //x=74.345 //y=4.795
c365 ( 106 0 ) capacitor c=0.0292043f //x=74.635 //y=4.795
c366 ( 103 0 ) capacitor c=0.0157913f //x=74.55 //y=1.365
c367 ( 101 0 ) capacitor c=0.0149844f //x=74.55 //y=0.71
c368 ( 97 0 ) capacitor c=0.0302441f //x=74.175 //y=1.915
c369 ( 96 0 ) capacitor c=0.0238107f //x=74.175 //y=1.52
c370 ( 95 0 ) capacitor c=0.0234352f //x=74.175 //y=1.21
c371 ( 94 0 ) capacitor c=0.0199931f //x=74.175 //y=0.865
c372 ( 90 0 ) capacitor c=0.0555336f //x=69.835 //y=4.79
c373 ( 89 0 ) capacitor c=0.0293157f //x=70.125 //y=4.79
c374 ( 88 0 ) capacitor c=0.0347816f //x=69.79 //y=1.22
c375 ( 87 0 ) capacitor c=0.0187487f //x=69.79 //y=0.875
c376 ( 81 0 ) capacitor c=0.0137055f //x=69.635 //y=1.375
c377 ( 79 0 ) capacitor c=0.0149861f //x=69.635 //y=0.72
c378 ( 78 0 ) capacitor c=0.096037f //x=69.26 //y=1.915
c379 ( 77 0 ) capacitor c=0.0228993f //x=69.26 //y=1.53
c380 ( 76 0 ) capacitor c=0.0234352f //x=69.26 //y=1.22
c381 ( 75 0 ) capacitor c=0.0198724f //x=69.26 //y=0.875
c382 ( 74 0 ) capacitor c=0.110336f //x=78.03 //y=6.025
c383 ( 73 0 ) capacitor c=0.154049f //x=77.59 //y=6.025
c384 ( 72 0 ) capacitor c=0.110003f //x=74.71 //y=6.025
c385 ( 71 0 ) capacitor c=0.15424f //x=74.27 //y=6.025
c386 ( 70 0 ) capacitor c=0.110114f //x=70.2 //y=6.02
c387 ( 69 0 ) capacitor c=0.158956f //x=69.76 //y=6.02
c388 ( 65 0 ) capacitor c=0.0023043f //x=67.23 //y=5.2
c389 ( 58 0 ) capacitor c=0.117496f //x=77.7 //y=2.08
c390 ( 50 0 ) capacitor c=0.0971978f //x=74 //y=2.08
c391 ( 42 0 ) capacitor c=0.0964287f //x=69.56 //y=2.08
c392 ( 40 0 ) capacitor c=0.104451f //x=67.71 //y=4.44
c393 ( 36 0 ) capacitor c=0.00404073f //x=67.355 //y=1.655
c394 ( 35 0 ) capacitor c=0.0122201f //x=67.625 //y=1.655
c395 ( 33 0 ) capacitor c=0.0139793f //x=67.625 //y=5.2
c396 ( 22 0 ) capacitor c=0.00272496f //x=66.435 //y=5.2
c397 ( 21 0 ) capacitor c=0.0154563f //x=67.145 //y=5.2
c398 ( 6 0 ) capacitor c=0.00561501f //x=74.115 //y=4.44
c399 ( 5 0 ) capacitor c=0.085624f //x=77.585 //y=4.44
c400 ( 4 0 ) capacitor c=0.00510592f //x=69.675 //y=4.44
c401 ( 3 0 ) capacitor c=0.100896f //x=73.885 //y=4.44
c402 ( 2 0 ) capacitor c=0.0110675f //x=67.825 //y=4.44
c403 ( 1 0 ) capacitor c=0.0443366f //x=69.445 //y=4.44
r404 (  150 152 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=77.59 //y=4.705 //x2=77.7 //y2=4.705
r405 (  129 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.035 //y=1.21 //x2=77.995 //y2=1.365
r406 (  128 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.035 //y=0.865 //x2=77.995 //y2=0.71
r407 (  128 129 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=78.035 //y=0.865 //x2=78.035 //y2=1.21
r408 (  125 152 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=78.03 //y=4.87 //x2=77.7 //y2=4.705
r409 (  123 149 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.66 //y=1.365 //x2=77.545 //y2=1.365
r410 (  122 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.88 //y=1.365 //x2=77.995 //y2=1.365
r411 (  121 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.66 //y=0.71 //x2=77.545 //y2=0.71
r412 (  120 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.88 //y=0.71 //x2=77.995 //y2=0.71
r413 (  120 121 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=77.88 //y=0.71 //x2=77.66 //y2=0.71
r414 (  117 150 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=77.59 //y=4.87 //x2=77.59 //y2=4.705
r415 (  116 147 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=77.505 //y=1.915 //x2=77.7 //y2=2.08
r416 (  115 149 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.505 //y=1.52 //x2=77.545 //y2=1.365
r417 (  115 116 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=77.505 //y=1.52 //x2=77.505 //y2=1.915
r418 (  114 149 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.505 //y=1.21 //x2=77.545 //y2=1.365
r419 (  113 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.505 //y=0.865 //x2=77.545 //y2=0.71
r420 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=77.505 //y=0.865 //x2=77.505 //y2=1.21
r421 (  109 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.705 //y=1.21 //x2=74.665 //y2=1.365
r422 (  108 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.705 //y=0.865 //x2=74.665 //y2=0.71
r423 (  108 109 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=74.705 //y=0.865 //x2=74.705 //y2=1.21
r424 (  106 110 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=74.635 //y=4.795 //x2=74.71 //y2=4.87
r425 (  106 107 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=74.635 //y=4.795 //x2=74.345 //y2=4.795
r426 (  104 143 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.33 //y=1.365 //x2=74.215 //y2=1.365
r427 (  103 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.55 //y=1.365 //x2=74.665 //y2=1.365
r428 (  102 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.33 //y=0.71 //x2=74.215 //y2=0.71
r429 (  101 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.55 //y=0.71 //x2=74.665 //y2=0.71
r430 (  101 102 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=74.55 //y=0.71 //x2=74.33 //y2=0.71
r431 (  98 107 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=74.27 //y=4.87 //x2=74.345 //y2=4.795
r432 (  98 141 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=74.27 //y=4.87 //x2=74 //y2=4.705
r433 (  97 139 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=74.175 //y=1.915 //x2=74 //y2=2.08
r434 (  96 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.175 //y=1.52 //x2=74.215 //y2=1.365
r435 (  96 97 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=74.175 //y=1.52 //x2=74.175 //y2=1.915
r436 (  95 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.175 //y=1.21 //x2=74.215 //y2=1.365
r437 (  94 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.175 //y=0.865 //x2=74.215 //y2=0.71
r438 (  94 95 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=74.175 //y=0.865 //x2=74.175 //y2=1.21
r439 (  89 91 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=70.125 //y=4.79 //x2=70.2 //y2=4.865
r440 (  89 90 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=70.125 //y=4.79 //x2=69.835 //y2=4.79
r441 (  88 137 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.79 //y=1.22 //x2=69.75 //y2=1.375
r442 (  87 136 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.79 //y=0.875 //x2=69.75 //y2=0.72
r443 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=69.79 //y=0.875 //x2=69.79 //y2=1.22
r444 (  84 90 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=69.76 //y=4.865 //x2=69.835 //y2=4.79
r445 (  84 135 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=69.76 //y=4.865 //x2=69.56 //y2=4.7
r446 (  82 131 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.415 //y=1.375 //x2=69.3 //y2=1.375
r447 (  81 137 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.635 //y=1.375 //x2=69.75 //y2=1.375
r448 (  80 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.415 //y=0.72 //x2=69.3 //y2=0.72
r449 (  79 136 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.635 //y=0.72 //x2=69.75 //y2=0.72
r450 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=69.635 //y=0.72 //x2=69.415 //y2=0.72
r451 (  78 133 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=69.26 //y=1.915 //x2=69.56 //y2=2.08
r452 (  77 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.26 //y=1.53 //x2=69.3 //y2=1.375
r453 (  77 78 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=69.26 //y=1.53 //x2=69.26 //y2=1.915
r454 (  76 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.26 //y=1.22 //x2=69.3 //y2=1.375
r455 (  75 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.26 //y=0.875 //x2=69.3 //y2=0.72
r456 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=69.26 //y=0.875 //x2=69.26 //y2=1.22
r457 (  74 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.03 //y=6.025 //x2=78.03 //y2=4.87
r458 (  73 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=77.59 //y=6.025 //x2=77.59 //y2=4.87
r459 (  72 110 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=74.71 //y=6.025 //x2=74.71 //y2=4.87
r460 (  71 98 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=74.27 //y=6.025 //x2=74.27 //y2=4.87
r461 (  70 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.2 //y=6.02 //x2=70.2 //y2=4.865
r462 (  69 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.76 //y=6.02 //x2=69.76 //y2=4.865
r463 (  68 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.365 //x2=77.88 //y2=1.365
r464 (  68 123 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.365 //x2=77.66 //y2=1.365
r465 (  67 103 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=74.44 //y=1.365 //x2=74.55 //y2=1.365
r466 (  67 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=74.44 //y=1.365 //x2=74.33 //y2=1.365
r467 (  66 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=69.525 //y=1.375 //x2=69.635 //y2=1.375
r468 (  66 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=69.525 //y=1.375 //x2=69.415 //y2=1.375
r469 (  63 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=77.7 //y=4.705 //x2=77.7 //y2=4.705
r470 (  61 63 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=77.7 //y=4.44 //x2=77.7 //y2=4.705
r471 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=77.7 //y=2.08 //x2=77.7 //y2=2.08
r472 (  58 61 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=77.7 //y=2.08 //x2=77.7 //y2=4.44
r473 (  55 141 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=74 //y=4.705 //x2=74 //y2=4.705
r474 (  53 55 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=74 //y=4.44 //x2=74 //y2=4.705
r475 (  50 139 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=74 //y=2.08 //x2=74 //y2=2.08
r476 (  50 53 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=74 //y=2.08 //x2=74 //y2=4.44
r477 (  47 135 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=69.56 //y=4.7 //x2=69.56 //y2=4.7
r478 (  45 47 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=69.56 //y=4.44 //x2=69.56 //y2=4.7
r479 (  42 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=69.56 //y=2.08 //x2=69.56 //y2=2.08
r480 (  42 45 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=69.56 //y=2.08 //x2=69.56 //y2=4.44
r481 (  38 40 ) resistor r=46.2032 //w=0.187 //l=0.675 //layer=li \
 //thickness=0.1 //x=67.71 //y=5.115 //x2=67.71 //y2=4.44
r482 (  37 40 ) resistor r=184.813 //w=0.187 //l=2.7 //layer=li \
 //thickness=0.1 //x=67.71 //y=1.74 //x2=67.71 //y2=4.44
r483 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=67.625 //y=1.655 //x2=67.71 //y2=1.74
r484 (  35 36 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=67.625 //y=1.655 //x2=67.355 //y2=1.655
r485 (  34 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.315 //y=5.2 //x2=67.23 //y2=5.2
r486 (  33 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=67.625 //y=5.2 //x2=67.71 //y2=5.115
r487 (  33 34 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=67.625 //y=5.2 //x2=67.315 //y2=5.2
r488 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=67.27 //y=1.57 //x2=67.355 //y2=1.655
r489 (  29 155 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.27 //y=1.57 //x2=67.27 //y2=1
r490 (  23 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.23 //y=5.285 //x2=67.23 //y2=5.2
r491 (  23 158 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=67.23 //y=5.285 //x2=67.23 //y2=5.725
r492 (  21 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.145 //y=5.2 //x2=67.23 //y2=5.2
r493 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=67.145 //y=5.2 //x2=66.435 //y2=5.2
r494 (  15 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=66.35 //y=5.285 //x2=66.435 //y2=5.2
r495 (  15 157 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=66.35 //y=5.285 //x2=66.35 //y2=5.725
r496 (  14 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=77.7 //y=4.44 //x2=77.7 //y2=4.44
r497 (  12 53 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=74 \
 //y=4.44 //x2=74 //y2=4.44
r498 (  10 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=69.56 //y=4.44 //x2=69.56 //y2=4.44
r499 (  8 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=67.71 //y=4.44 //x2=67.71 //y2=4.44
r500 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=74.115 //y=4.44 //x2=74 //y2=4.44
r501 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=77.585 //y=4.44 //x2=77.7 //y2=4.44
r502 (  5 6 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=77.585 //y=4.44 //x2=74.115 //y2=4.44
r503 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.675 //y=4.44 //x2=69.56 //y2=4.44
r504 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=73.885 //y=4.44 //x2=74 //y2=4.44
r505 (  3 4 ) resistor r=4.01718 //w=0.131 //l=4.21 //layer=m1 \
 //thickness=0.36 //x=73.885 //y=4.44 //x2=69.675 //y2=4.44
r506 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=67.825 //y=4.44 //x2=67.71 //y2=4.44
r507 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.445 //y=4.44 //x2=69.56 //y2=4.44
r508 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=69.445 //y=4.44 //x2=67.825 //y2=4.44
ends PM_TMRDFFSNQNX1\%noxref_23

subckt PM_TMRDFFSNQNX1\%noxref_24 ( 1 2 3 4 5 6 23 24 35 37 38 42 44 52 61 67 \
 68 69 70 71 72 73 74 75 76 77 78 79 80 81 83 89 90 91 92 99 100 101 102 103 \
 105 108 111 112 113 114 115 116 117 118 122 124 127 128 129 130 151 158 160 \
 161 )
c450 ( 161 0 ) capacitor c=0.0220291f //x=18.245 //y=5.02
c451 ( 160 0 ) capacitor c=0.0217503f //x=17.365 //y=5.02
c452 ( 158 0 ) capacitor c=0.0084702f //x=18.24 //y=0.905
c453 ( 151 0 ) capacitor c=0.0583848f //x=80.66 //y=2.08
c454 ( 130 0 ) capacitor c=0.0316774f //x=81.365 //y=1.21
c455 ( 129 0 ) capacitor c=0.0187384f //x=81.365 //y=0.865
c456 ( 128 0 ) capacitor c=0.0590362f //x=81.005 //y=4.795
c457 ( 127 0 ) capacitor c=0.0296075f //x=81.295 //y=4.795
c458 ( 124 0 ) capacitor c=0.0157912f //x=81.21 //y=1.365
c459 ( 122 0 ) capacitor c=0.0149844f //x=81.21 //y=0.71
c460 ( 118 0 ) capacitor c=0.0302441f //x=80.835 //y=1.915
c461 ( 117 0 ) capacitor c=0.0234157f //x=80.835 //y=1.52
c462 ( 116 0 ) capacitor c=0.0234376f //x=80.835 //y=1.21
c463 ( 115 0 ) capacitor c=0.0199931f //x=80.835 //y=0.865
c464 ( 114 0 ) capacitor c=0.0962905f //x=79.005 //y=1.915
c465 ( 113 0 ) capacitor c=0.0249466f //x=79.005 //y=1.56
c466 ( 112 0 ) capacitor c=0.0234397f //x=79.005 //y=1.25
c467 ( 111 0 ) capacitor c=0.0193195f //x=79.005 //y=0.905
c468 ( 108 0 ) capacitor c=0.0631944f //x=78.91 //y=4.87
c469 ( 105 0 ) capacitor c=0.0187941f //x=78.85 //y=1.405
c470 ( 103 0 ) capacitor c=0.0157803f //x=78.85 //y=0.75
c471 ( 102 0 ) capacitor c=0.010629f //x=78.545 //y=4.795
c472 ( 101 0 ) capacitor c=0.0194269f //x=78.835 //y=4.795
c473 ( 100 0 ) capacitor c=0.0365717f //x=78.475 //y=1.25
c474 ( 99 0 ) capacitor c=0.0175988f //x=78.475 //y=0.905
c475 ( 92 0 ) capacitor c=0.0556143f //x=20.995 //y=4.79
c476 ( 91 0 ) capacitor c=0.0293157f //x=21.285 //y=4.79
c477 ( 90 0 ) capacitor c=0.0347816f //x=20.95 //y=1.22
c478 ( 89 0 ) capacitor c=0.0187487f //x=20.95 //y=0.875
c479 ( 83 0 ) capacitor c=0.0137055f //x=20.795 //y=1.375
c480 ( 81 0 ) capacitor c=0.0149861f //x=20.795 //y=0.72
c481 ( 80 0 ) capacitor c=0.096037f //x=20.42 //y=1.915
c482 ( 79 0 ) capacitor c=0.0228993f //x=20.42 //y=1.53
c483 ( 78 0 ) capacitor c=0.0234352f //x=20.42 //y=1.22
c484 ( 77 0 ) capacitor c=0.0198724f //x=20.42 //y=0.875
c485 ( 76 0 ) capacitor c=0.110622f //x=81.37 //y=6.025
c486 ( 75 0 ) capacitor c=0.154068f //x=80.93 //y=6.025
c487 ( 74 0 ) capacitor c=0.154291f //x=78.91 //y=6.025
c488 ( 73 0 ) capacitor c=0.110404f //x=78.47 //y=6.025
c489 ( 72 0 ) capacitor c=0.110114f //x=21.36 //y=6.02
c490 ( 71 0 ) capacitor c=0.158956f //x=20.92 //y=6.02
c491 ( 67 0 ) capacitor c=0.00211606f //x=18.39 //y=5.2
c492 ( 61 0 ) capacitor c=0.100881f //x=80.66 //y=2.08
c493 ( 52 0 ) capacitor c=0.105667f //x=79.18 //y=2.08
c494 ( 44 0 ) capacitor c=0.0962061f //x=20.72 //y=2.08
c495 ( 42 0 ) capacitor c=0.104221f //x=18.87 //y=3.33
c496 ( 38 0 ) capacitor c=0.00404073f //x=18.515 //y=1.655
c497 ( 37 0 ) capacitor c=0.0122201f //x=18.785 //y=1.655
c498 ( 35 0 ) capacitor c=0.0137995f //x=18.785 //y=5.2
c499 ( 24 0 ) capacitor c=0.00251459f //x=17.595 //y=5.2
c500 ( 23 0 ) capacitor c=0.0143649f //x=18.305 //y=5.2
c501 ( 6 0 ) capacitor c=0.0112698f //x=79.295 //y=2.08
c502 ( 5 0 ) capacitor c=0.0463273f //x=80.545 //y=2.08
c503 ( 4 0 ) capacitor c=0.004304f //x=20.835 //y=3.33
c504 ( 3 0 ) capacitor c=0.987666f //x=79.065 //y=3.33
c505 ( 2 0 ) capacitor c=0.0124845f //x=18.985 //y=3.33
c506 ( 1 0 ) capacitor c=0.0280612f //x=20.605 //y=3.33
r507 (  130 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.365 //y=1.21 //x2=81.325 //y2=1.365
r508 (  129 156 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.365 //y=0.865 //x2=81.325 //y2=0.71
r509 (  129 130 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=81.365 //y=0.865 //x2=81.365 //y2=1.21
r510 (  127 131 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=81.295 //y=4.795 //x2=81.37 //y2=4.87
r511 (  127 128 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=81.295 //y=4.795 //x2=81.005 //y2=4.795
r512 (  125 155 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.99 //y=1.365 //x2=80.875 //y2=1.365
r513 (  124 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=81.21 //y=1.365 //x2=81.325 //y2=1.365
r514 (  123 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.99 //y=0.71 //x2=80.875 //y2=0.71
r515 (  122 156 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=81.21 //y=0.71 //x2=81.325 //y2=0.71
r516 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=81.21 //y=0.71 //x2=80.99 //y2=0.71
r517 (  119 128 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=80.93 //y=4.87 //x2=81.005 //y2=4.795
r518 (  119 153 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=80.93 //y=4.87 //x2=80.66 //y2=4.705
r519 (  118 151 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=80.835 //y=1.915 //x2=80.66 //y2=2.08
r520 (  117 155 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.835 //y=1.52 //x2=80.875 //y2=1.365
r521 (  117 118 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=80.835 //y=1.52 //x2=80.835 //y2=1.915
r522 (  116 155 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.835 //y=1.21 //x2=80.875 //y2=1.365
r523 (  115 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.835 //y=0.865 //x2=80.875 //y2=0.71
r524 (  115 116 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=80.835 //y=0.865 //x2=80.835 //y2=1.21
r525 (  114 147 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=79.005 //y=1.915 //x2=79.18 //y2=2.08
r526 (  113 145 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.005 //y=1.56 //x2=78.965 //y2=1.405
r527 (  113 114 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=79.005 //y=1.56 //x2=79.005 //y2=1.915
r528 (  112 145 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.005 //y=1.25 //x2=78.965 //y2=1.405
r529 (  111 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.005 //y=0.905 //x2=78.965 //y2=0.75
r530 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=79.005 //y=0.905 //x2=79.005 //y2=1.25
r531 (  108 149 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=78.91 //y=4.87 //x2=79.18 //y2=4.705
r532 (  106 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.63 //y=1.405 //x2=78.515 //y2=1.405
r533 (  105 145 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.85 //y=1.405 //x2=78.965 //y2=1.405
r534 (  104 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.63 //y=0.75 //x2=78.515 //y2=0.75
r535 (  103 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.85 //y=0.75 //x2=78.965 //y2=0.75
r536 (  103 104 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=78.85 //y=0.75 //x2=78.63 //y2=0.75
r537 (  101 108 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=78.835 //y=4.795 //x2=78.91 //y2=4.87
r538 (  101 102 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=78.835 //y=4.795 //x2=78.545 //y2=4.795
r539 (  100 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.475 //y=1.25 //x2=78.515 //y2=1.405
r540 (  99 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.475 //y=0.905 //x2=78.515 //y2=0.75
r541 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=78.475 //y=0.905 //x2=78.475 //y2=1.25
r542 (  96 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=78.47 //y=4.87 //x2=78.545 //y2=4.795
r543 (  91 93 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.285 //y=4.79 //x2=21.36 //y2=4.865
r544 (  91 92 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=21.285 //y=4.79 //x2=20.995 //y2=4.79
r545 (  90 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.95 //y=1.22 //x2=20.91 //y2=1.375
r546 (  89 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.95 //y=0.875 //x2=20.91 //y2=0.72
r547 (  89 90 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.95 //y=0.875 //x2=20.95 //y2=1.22
r548 (  86 92 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.92 //y=4.865 //x2=20.995 //y2=4.79
r549 (  86 139 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=20.92 //y=4.865 //x2=20.72 //y2=4.7
r550 (  84 135 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.575 //y=1.375 //x2=20.46 //y2=1.375
r551 (  83 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.795 //y=1.375 //x2=20.91 //y2=1.375
r552 (  82 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.575 //y=0.72 //x2=20.46 //y2=0.72
r553 (  81 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.795 //y=0.72 //x2=20.91 //y2=0.72
r554 (  81 82 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.795 //y=0.72 //x2=20.575 //y2=0.72
r555 (  80 137 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.915 //x2=20.72 //y2=2.08
r556 (  79 135 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.53 //x2=20.46 //y2=1.375
r557 (  79 80 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.53 //x2=20.42 //y2=1.915
r558 (  78 135 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.22 //x2=20.46 //y2=1.375
r559 (  77 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=0.875 //x2=20.46 //y2=0.72
r560 (  77 78 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.42 //y=0.875 //x2=20.42 //y2=1.22
r561 (  76 131 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=81.37 //y=6.025 //x2=81.37 //y2=4.87
r562 (  75 119 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=80.93 //y=6.025 //x2=80.93 //y2=4.87
r563 (  74 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.91 //y=6.025 //x2=78.91 //y2=4.87
r564 (  73 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.47 //y=6.025 //x2=78.47 //y2=4.87
r565 (  72 93 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.36 //y=6.02 //x2=21.36 //y2=4.865
r566 (  71 86 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.92 //y=6.02 //x2=20.92 //y2=4.865
r567 (  70 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=81.1 //y=1.365 //x2=81.21 //y2=1.365
r568 (  70 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=81.1 //y=1.365 //x2=80.99 //y2=1.365
r569 (  69 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.74 //y=1.405 //x2=78.85 //y2=1.405
r570 (  69 106 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.74 //y=1.405 //x2=78.63 //y2=1.405
r571 (  68 83 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.685 //y=1.375 //x2=20.795 //y2=1.375
r572 (  68 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.685 //y=1.375 //x2=20.575 //y2=1.375
r573 (  65 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=80.66 //y=4.705 //x2=80.66 //y2=4.705
r574 (  61 151 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=80.66 //y=2.08 //x2=80.66 //y2=2.08
r575 (  61 65 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=80.66 //y=2.08 //x2=80.66 //y2=4.705
r576 (  58 149 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.18 //y=4.705 //x2=79.18 //y2=4.705
r577 (  56 58 ) resistor r=94.1176 //w=0.187 //l=1.375 //layer=li \
 //thickness=0.1 //x=79.18 //y=3.33 //x2=79.18 //y2=4.705
r578 (  52 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.18 //y=2.08 //x2=79.18 //y2=2.08
r579 (  52 56 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=79.18 //y=2.08 //x2=79.18 //y2=3.33
r580 (  49 139 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.72 //y=4.7 //x2=20.72 //y2=4.7
r581 (  47 49 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=20.72 //y=3.33 //x2=20.72 //y2=4.7
r582 (  44 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.72 //y=2.08 //x2=20.72 //y2=2.08
r583 (  44 47 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.08 //x2=20.72 //y2=3.33
r584 (  40 42 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=18.87 //y=5.115 //x2=18.87 //y2=3.33
r585 (  39 42 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=18.87 //y=1.74 //x2=18.87 //y2=3.33
r586 (  37 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.785 //y=1.655 //x2=18.87 //y2=1.74
r587 (  37 38 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=18.785 //y=1.655 //x2=18.515 //y2=1.655
r588 (  36 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.475 //y=5.2 //x2=18.39 //y2=5.2
r589 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.785 //y=5.2 //x2=18.87 //y2=5.115
r590 (  35 36 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=18.785 //y=5.2 //x2=18.475 //y2=5.2
r591 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.43 //y=1.57 //x2=18.515 //y2=1.655
r592 (  31 158 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=18.43 //y=1.57 //x2=18.43 //y2=1
r593 (  25 67 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.39 //y=5.285 //x2=18.39 //y2=5.2
r594 (  25 161 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=18.39 //y=5.285 //x2=18.39 //y2=5.725
r595 (  23 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.305 //y=5.2 //x2=18.39 //y2=5.2
r596 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=18.305 //y=5.2 //x2=17.595 //y2=5.2
r597 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.51 //y=5.285 //x2=17.595 //y2=5.2
r598 (  17 160 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=17.51 //y=5.285 //x2=17.51 //y2=5.725
r599 (  16 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=80.66 //y=2.08 //x2=80.66 //y2=2.08
r600 (  14 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.18 //y=3.33 //x2=79.18 //y2=3.33
r601 (  12 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.18 //y=2.08 //x2=79.18 //y2=2.08
r602 (  10 47 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.72 //y=3.33 //x2=20.72 //y2=3.33
r603 (  8 42 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.87 //y=3.33 //x2=18.87 //y2=3.33
r604 (  6 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.295 //y=2.08 //x2=79.18 //y2=2.08
r605 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=80.545 //y=2.08 //x2=80.66 //y2=2.08
r606 (  5 6 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=80.545 //y=2.08 //x2=79.295 //y2=2.08
r607 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.835 //y=3.33 //x2=20.72 //y2=3.33
r608 (  3 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.065 //y=3.33 //x2=79.18 //y2=3.33
r609 (  3 4 ) resistor r=55.563 //w=0.131 //l=58.23 //layer=m1 \
 //thickness=0.36 //x=79.065 //y=3.33 //x2=20.835 //y2=3.33
r610 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.985 //y=3.33 //x2=18.87 //y2=3.33
r611 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=3.33 //x2=20.72 //y2=3.33
r612 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=20.605 //y=3.33 //x2=18.985 //y2=3.33
ends PM_TMRDFFSNQNX1\%noxref_24

subckt PM_TMRDFFSNQNX1\%noxref_25 ( 1 2 13 14 15 21 27 28 35 46 47 48 49 50 )
c89 ( 50 0 ) capacitor c=0.0308836f //x=82.325 //y=5.025
c90 ( 49 0 ) capacitor c=0.0173945f //x=81.445 //y=5.025
c91 ( 47 0 ) capacitor c=0.0169278f //x=78.545 //y=5.025
c92 ( 46 0 ) capacitor c=0.0166762f //x=77.665 //y=5.025
c93 ( 45 0 ) capacitor c=0.00115294f //x=81.59 //y=6.91
c94 ( 35 0 ) capacitor c=0.0132983f //x=82.385 //y=6.91
c95 ( 28 0 ) capacitor c=0.00388794f //x=80.795 //y=6.91
c96 ( 27 0 ) capacitor c=0.00985708f //x=81.505 //y=6.91
c97 ( 21 0 ) capacitor c=0.0442221f //x=80.71 //y=5.21
c98 ( 15 0 ) capacitor c=0.0105083f //x=78.69 //y=5.295
c99 ( 14 0 ) capacitor c=0.00227812f //x=77.895 //y=5.21
c100 ( 13 0 ) capacitor c=0.0174384f //x=78.605 //y=5.21
c101 ( 2 0 ) capacitor c=0.00682032f //x=78.805 //y=5.21
c102 ( 1 0 ) capacitor c=0.0574911f //x=80.595 //y=5.21
r103 (  37 50 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.47 //y=6.825 //x2=82.47 //y2=6.74
r104 (  36 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.675 //y=6.91 //x2=81.59 //y2=6.91
r105 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=82.385 //y=6.91 //x2=82.47 //y2=6.825
r106 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=82.385 //y=6.91 //x2=81.675 //y2=6.91
r107 (  29 45 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.59 //y=6.825 //x2=81.59 //y2=6.91
r108 (  29 49 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.59 //y=6.825 //x2=81.59 //y2=6.74
r109 (  27 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.505 //y=6.91 //x2=81.59 //y2=6.91
r110 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=81.505 //y=6.91 //x2=80.795 //y2=6.91
r111 (  21 48 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=80.71 //y=5.21 //x2=80.71 //y2=6.06
r112 (  19 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=80.71 //y=6.825 //x2=80.795 //y2=6.91
r113 (  19 48 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.71 //y=6.825 //x2=80.71 //y2=6.74
r114 (  15 44 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=78.69 //y=5.295 //x2=78.69 //y2=5.17
r115 (  15 47 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=78.69 //y=5.295 //x2=78.69 //y2=6.06
r116 (  13 44 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.605 //y=5.21 //x2=78.69 //y2=5.17
r117 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=78.605 //y=5.21 //x2=77.895 //y2=5.21
r118 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=77.81 //y=5.295 //x2=77.895 //y2=5.21
r119 (  7 46 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=77.81 //y=5.295 //x2=77.81 //y2=5.72
r120 (  6 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=80.71 //y=5.21 //x2=80.71 //y2=5.21
r121 (  4 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=78.69 //y=5.21 //x2=78.69 //y2=5.21
r122 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=78.805 //y=5.21 //x2=78.69 //y2=5.21
r123 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=80.595 //y=5.21 //x2=80.71 //y2=5.21
r124 (  1 2 ) resistor r=1.70802 //w=0.131 //l=1.79 //layer=m1 \
 //thickness=0.36 //x=80.595 //y=5.21 //x2=78.805 //y2=5.21
ends PM_TMRDFFSNQNX1\%noxref_25

subckt PM_TMRDFFSNQNX1\%QN ( 1 2 3 4 11 12 13 14 15 16 17 30 31 44 46 47 61 62 \
 63 64 68 69 )
c169 ( 69 0 ) capacitor c=0.0167617f //x=81.885 //y=5.025
c170 ( 68 0 ) capacitor c=0.0164812f //x=81.005 //y=5.025
c171 ( 64 0 ) capacitor c=0.0108176f //x=81.88 //y=0.905
c172 ( 63 0 ) capacitor c=0.0131637f //x=78.55 //y=0.905
c173 ( 62 0 ) capacitor c=0.0131367f //x=75.22 //y=0.905
c174 ( 61 0 ) capacitor c=0.00421476f //x=82.03 //y=5.21
c175 ( 47 0 ) capacitor c=0.00775877f //x=82.155 //y=1.645
c176 ( 46 0 ) capacitor c=0.0165978f //x=82.425 //y=1.645
c177 ( 44 0 ) capacitor c=0.0160142f //x=82.425 //y=5.21
c178 ( 31 0 ) capacitor c=0.0029383f //x=81.235 //y=5.21
c179 ( 30 0 ) capacitor c=0.0155464f //x=81.945 //y=5.21
c180 ( 11 0 ) capacitor c=0.133166f //x=82.51 //y=2.22
c181 ( 4 0 ) capacitor c=0.0054338f //x=78.855 //y=1.18
c182 ( 3 0 ) capacitor c=0.0704773f //x=81.955 //y=1.18
c183 ( 2 0 ) capacitor c=0.0153777f //x=75.525 //y=1.18
c184 ( 1 0 ) capacitor c=0.0651236f //x=78.625 //y=1.18
r185 (  60 62 ) resistor r=13.3953 //w=0.172 //l=0.18 //layer=li \
 //thickness=0.1 //x=75.407 //y=1.18 //x2=75.407 //y2=1
r186 (  46 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=82.425 //y=1.645 //x2=82.51 //y2=1.73
r187 (  46 47 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=82.425 //y=1.645 //x2=82.155 //y2=1.645
r188 (  45 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.115 //y=5.21 //x2=82.03 //y2=5.21
r189 (  44 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=82.425 //y=5.21 //x2=82.51 //y2=5.125
r190 (  44 45 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=82.425 //y=5.21 //x2=82.115 //y2=5.21
r191 (  43 64 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=82.07 //y=1.18 //x2=82.07 //y2=1
r192 (  38 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=82.07 //y=1.56 //x2=82.155 //y2=1.645
r193 (  38 43 ) resistor r=26.0107 //w=0.187 //l=0.38 //layer=li \
 //thickness=0.1 //x=82.07 //y=1.56 //x2=82.07 //y2=1.18
r194 (  32 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.03 //y=5.295 //x2=82.03 //y2=5.21
r195 (  32 69 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=82.03 //y=5.295 //x2=82.03 //y2=5.72
r196 (  30 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.945 //y=5.21 //x2=82.03 //y2=5.21
r197 (  30 31 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=81.945 //y=5.21 //x2=81.235 //y2=5.21
r198 (  24 31 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=81.15 //y=5.295 //x2=81.235 //y2=5.21
r199 (  24 68 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=81.15 //y=5.295 //x2=81.15 //y2=5.72
r200 (  22 63 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=78.74 //y=1.18 //x2=78.74 //y2=1
r201 (  17 49 ) resistor r=46.8877 //w=0.187 //l=0.685 //layer=li \
 //thickness=0.1 //x=82.51 //y=4.44 //x2=82.51 //y2=5.125
r202 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=82.51 //y=4.07 //x2=82.51 //y2=4.44
r203 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=82.51 //y=3.7 //x2=82.51 //y2=4.07
r204 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=82.51 //y=3.33 //x2=82.51 //y2=3.7
r205 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=82.51 //y=2.96 //x2=82.51 //y2=3.33
r206 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=82.51 //y=2.59 //x2=82.51 //y2=2.96
r207 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=82.51 //y=2.22 //x2=82.51 //y2=2.59
r208 (  11 48 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=82.51 //y=2.22 //x2=82.51 //y2=1.73
r209 (  10 43 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=82.07 //y=1.18 //x2=82.07 //y2=1.18
r210 (  8 22 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=78.74 //y=1.18 //x2=78.74 //y2=1.18
r211 (  6 60 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.41 //y=1.18 //x2=75.41 //y2=1.18
r212 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=78.855 //y=1.18 //x2=78.74 //y2=1.18
r213 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=81.955 //y=1.18 //x2=82.07 //y2=1.18
r214 (  3 4 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=81.955 //y=1.18 //x2=78.855 //y2=1.18
r215 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.525 //y=1.18 //x2=75.41 //y2=1.18
r216 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=78.625 //y=1.18 //x2=78.74 //y2=1.18
r217 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=78.625 //y=1.18 //x2=75.525 //y2=1.18
ends PM_TMRDFFSNQNX1\%QN

subckt PM_TMRDFFSNQNX1\%noxref_27 ( 1 5 9 10 13 17 29 )
c50 ( 29 0 ) capacitor c=0.0632971f //x=0.56 //y=0.365
c51 ( 17 0 ) capacitor c=0.0072343f //x=2.635 //y=0.615
c52 ( 13 0 ) capacitor c=0.0147753f //x=2.55 //y=0.53
c53 ( 10 0 ) capacitor c=0.00638095f //x=1.665 //y=1.495
c54 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c55 ( 5 0 ) capacitor c=0.02021f //x=1.58 //y=1.58
c56 ( 1 0 ) capacitor c=0.0113547f //x=0.695 //y=1.495
r57 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r58 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r59 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r60 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=2.15 //y2=0.53
r61 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r62 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.15 //y2=0.53
r63 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r64 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r65 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r66 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r67 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r68 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r69 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r70 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r71 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r72 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_27

subckt PM_TMRDFFSNQNX1\%noxref_28 ( 1 5 9 13 17 35 )
c51 ( 35 0 ) capacitor c=0.0680128f //x=3.785 //y=0.375
c52 ( 17 0 ) capacitor c=0.018806f //x=5.775 //y=1.59
c53 ( 13 0 ) capacitor c=0.0155484f //x=5.775 //y=0.54
c54 ( 9 0 ) capacitor c=0.00678203f //x=4.89 //y=0.625
c55 ( 5 0 ) capacitor c=0.017077f //x=4.805 //y=1.59
c56 ( 1 0 ) capacitor c=0.00729042f //x=3.92 //y=1.505
r57 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.975 //y=1.59 //x2=4.89 //y2=1.63
r58 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.975 //y=1.59 //x2=5.375 //y2=1.59
r59 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.775 //y=1.59 //x2=5.86 //y2=1.59
r60 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.775 //y=1.59 //x2=5.375 //y2=1.59
r61 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.975 //y=0.54 //x2=4.89 //y2=0.5
r62 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.975 //y=0.54 //x2=5.375 //y2=0.54
r63 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.775 //y=0.54 //x2=5.86 //y2=0.54
r64 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.775 //y=0.54 //x2=5.375 //y2=0.54
r65 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.89 //y=1.505 //x2=4.89 //y2=1.63
r66 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=4.89 //y=1.505 //x2=4.89 //y2=0.89
r67 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=4.89 //y=0.625 //x2=4.89 //y2=0.5
r68 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=4.89 //y=0.625 //x2=4.89 //y2=0.89
r69 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.005 //y=1.59 //x2=3.92 //y2=1.63
r70 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.005 //y=1.59 //x2=4.405 //y2=1.59
r71 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.805 //y=1.59 //x2=4.89 //y2=1.63
r72 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.805 //y=1.59 //x2=4.405 //y2=1.59
r73 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.92 //y=1.505 //x2=3.92 //y2=1.63
r74 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=3.92 //y=1.505 //x2=3.92 //y2=0.89
ends PM_TMRDFFSNQNX1\%noxref_28

subckt PM_TMRDFFSNQNX1\%noxref_29 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.041888f //x=6.295 //y=0.375
c53 ( 28 0 ) capacitor c=0.00460056f //x=5.19 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=6.43 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=7.4 //y=0.625
c56 ( 11 0 ) capacitor c=0.0145763f //x=7.315 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=6.43 //y=0.625
c58 ( 1 0 ) capacitor c=0.022715f //x=6.345 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.4 //y=0.625 //x2=7.4 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=7.4 //y=0.625 //x2=7.4 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.515 //y=0.54 //x2=6.43 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.515 //y=0.54 //x2=6.915 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.315 //y=0.54 //x2=7.4 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.315 //y=0.54 //x2=6.915 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.43 //y=1.08 //x2=6.43 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=6.43 //y=1.08 //x2=6.43 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.91 //x2=6.43 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.91 //x2=6.43 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.625 //x2=6.43 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.625 //x2=6.43 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.465 //y=0.995 //x2=5.38 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.345 //y=0.995 //x2=6.43 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=6.345 //y=0.995 //x2=5.465 //y2=0.995
ends PM_TMRDFFSNQNX1\%noxref_29

subckt PM_TMRDFFSNQNX1\%noxref_30 ( 1 5 9 13 17 35 )
c53 ( 35 0 ) capacitor c=0.0679545f //x=8.595 //y=0.375
c54 ( 17 0 ) capacitor c=0.0193993f //x=10.585 //y=1.59
c55 ( 13 0 ) capacitor c=0.0155066f //x=10.585 //y=0.54
c56 ( 9 0 ) capacitor c=0.00678203f //x=9.7 //y=0.625
c57 ( 5 0 ) capacitor c=0.0174845f //x=9.615 //y=1.59
c58 ( 1 0 ) capacitor c=0.00729042f //x=8.73 //y=1.505
r59 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.785 //y=1.59 //x2=9.7 //y2=1.63
r60 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.785 //y=1.59 //x2=10.185 //y2=1.59
r61 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.585 //y=1.59 //x2=10.67 //y2=1.59
r62 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.585 //y=1.59 //x2=10.185 //y2=1.59
r63 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.785 //y=0.54 //x2=9.7 //y2=0.5
r64 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.785 //y=0.54 //x2=10.185 //y2=0.54
r65 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.585 //y=0.54 //x2=10.67 //y2=0.54
r66 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.585 //y=0.54 //x2=10.185 //y2=0.54
r67 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.7 //y=1.505 //x2=9.7 //y2=1.63
r68 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.7 //y=1.505 //x2=9.7 //y2=0.89
r69 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.7 //y=0.625 //x2=9.7 //y2=0.5
r70 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=9.7 //y=0.625 //x2=9.7 //y2=0.89
r71 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.815 //y=1.59 //x2=8.73 //y2=1.63
r72 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.815 //y=1.59 //x2=9.215 //y2=1.59
r73 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.615 //y=1.59 //x2=9.7 //y2=1.63
r74 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.615 //y=1.59 //x2=9.215 //y2=1.59
r75 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.73 //y=1.505 //x2=8.73 //y2=1.63
r76 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.73 //y=1.505 //x2=8.73 //y2=0.89
ends PM_TMRDFFSNQNX1\%noxref_30

subckt PM_TMRDFFSNQNX1\%noxref_31 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=11.105 //y=0.375
c53 ( 28 0 ) capacitor c=0.00460343f //x=10 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=11.24 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=12.21 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=12.125 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=11.24 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=11.155 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=12.21 //y=0.625 //x2=12.21 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=12.21 //y=0.625 //x2=12.21 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.325 //y=0.54 //x2=11.24 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.325 //y=0.54 //x2=11.725 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.125 //y=0.54 //x2=12.21 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.125 //y=0.54 //x2=11.725 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.24 //y=1.08 //x2=11.24 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=11.24 //y=1.08 //x2=11.24 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.91 //x2=11.24 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.91 //x2=11.24 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.625 //x2=11.24 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.625 //x2=11.24 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.275 //y=0.995 //x2=10.19 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.155 //y=0.995 //x2=11.24 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=11.155 //y=0.995 //x2=10.275 //y2=0.995
ends PM_TMRDFFSNQNX1\%noxref_31

subckt PM_TMRDFFSNQNX1\%noxref_32 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=13.51 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722223f //x=15.585 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=15.5 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=14.615 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=14.615 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=14.53 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=13.645 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=15.585 //y=0.615 //x2=15.585 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.585 //y=0.615 //x2=15.585 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.7 //y=0.53 //x2=14.615 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.7 //y=0.53 //x2=15.1 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.5 //y=0.53 //x2=15.585 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.5 //y=0.53 //x2=15.1 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.615 //y=1.495 //x2=14.615 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=14.615 //y=1.495 //x2=14.615 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=14.615 //y=0.615 //x2=14.615 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=14.615 //y=0.615 //x2=14.615 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.73 //y=1.58 //x2=13.645 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.73 //y=1.58 //x2=14.13 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.53 //y=1.58 //x2=14.615 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.53 //y=1.58 //x2=14.13 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=13.645 //y=1.495 //x2=13.645 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.645 //y=1.495 //x2=13.645 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_32

subckt PM_TMRDFFSNQNX1\%noxref_33 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632684f //x=16.84 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=18.915 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=18.83 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=17.945 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=17.945 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=17.86 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=16.975 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=18.915 //y=0.615 //x2=18.915 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.915 //y=0.615 //x2=18.915 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.03 //y=0.53 //x2=17.945 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.03 //y=0.53 //x2=18.43 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.83 //y=0.53 //x2=18.915 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.83 //y=0.53 //x2=18.43 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=17.945 //y=1.495 //x2=17.945 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=17.945 //y=1.495 //x2=17.945 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=17.945 //y=0.615 //x2=17.945 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=17.945 //y=0.615 //x2=17.945 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.06 //y=1.58 //x2=16.975 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.06 //y=1.58 //x2=17.46 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.86 //y=1.58 //x2=17.945 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.86 //y=1.58 //x2=17.46 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=16.975 //y=1.495 //x2=16.975 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=16.975 //y=1.495 //x2=16.975 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_33

subckt PM_TMRDFFSNQNX1\%noxref_34 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=20.065 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=22.055 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=22.055 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=21.17 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=21.085 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=20.2 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.255 //y=1.59 //x2=21.17 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.255 //y=1.59 //x2=21.655 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.055 //y=1.59 //x2=22.14 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.055 //y=1.59 //x2=21.655 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.255 //y=0.54 //x2=21.17 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.255 //y=0.54 //x2=21.655 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.055 //y=0.54 //x2=22.14 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.055 //y=0.54 //x2=21.655 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=21.17 //y=1.505 //x2=21.17 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=21.17 //y=1.505 //x2=21.17 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=21.17 //y=0.625 //x2=21.17 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=21.17 //y=0.625 //x2=21.17 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.285 //y=1.59 //x2=20.2 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.285 //y=1.59 //x2=20.685 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.085 //y=1.59 //x2=21.17 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.085 //y=1.59 //x2=20.685 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.2 //y=1.505 //x2=20.2 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=20.2 //y=1.505 //x2=20.2 //y2=0.89
ends PM_TMRDFFSNQNX1\%noxref_34

subckt PM_TMRDFFSNQNX1\%noxref_35 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=22.575 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=21.47 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=22.71 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=23.68 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=23.595 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=22.71 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=22.625 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.68 //y=0.625 //x2=23.68 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=23.68 //y=0.625 //x2=23.68 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.795 //y=0.54 //x2=22.71 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.795 //y=0.54 //x2=23.195 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.595 //y=0.54 //x2=23.68 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.595 //y=0.54 //x2=23.195 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.71 //y=1.08 //x2=22.71 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=22.71 //y=1.08 //x2=22.71 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.91 //x2=22.71 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.91 //x2=22.71 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.625 //x2=22.71 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.625 //x2=22.71 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.745 //y=0.995 //x2=21.66 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.625 //y=0.995 //x2=22.71 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=22.625 //y=0.995 //x2=21.745 //y2=0.995
ends PM_TMRDFFSNQNX1\%noxref_35

subckt PM_TMRDFFSNQNX1\%noxref_36 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0633518f //x=24.98 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=27.055 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=26.97 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=26.085 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=26.085 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=26 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=25.115 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=27.055 //y=0.615 //x2=27.055 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=27.055 //y=0.615 //x2=27.055 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=26.17 //y=0.53 //x2=26.085 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.17 //y=0.53 //x2=26.57 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=26.97 //y=0.53 //x2=27.055 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.97 //y=0.53 //x2=26.57 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=26.085 //y=1.495 //x2=26.085 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=26.085 //y=1.495 //x2=26.085 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=26.085 //y=0.615 //x2=26.085 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=26.085 //y=0.615 //x2=26.085 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.2 //y=1.58 //x2=25.115 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.2 //y=1.58 //x2=25.6 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=26 //y=1.58 //x2=26.085 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26 //y=1.58 //x2=25.6 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=25.115 //y=1.495 //x2=25.115 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=25.115 //y=1.495 //x2=25.115 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_36

subckt PM_TMRDFFSNQNX1\%noxref_37 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673195f //x=28.205 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=30.195 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=30.195 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=29.31 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=29.225 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=28.34 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.395 //y=1.59 //x2=29.31 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.395 //y=1.59 //x2=29.795 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.195 //y=1.59 //x2=30.28 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.195 //y=1.59 //x2=29.795 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.395 //y=0.54 //x2=29.31 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.395 //y=0.54 //x2=29.795 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.195 //y=0.54 //x2=30.28 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.195 //y=0.54 //x2=29.795 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=29.31 //y=1.505 //x2=29.31 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=29.31 //y=1.505 //x2=29.31 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=29.31 //y=0.625 //x2=29.31 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=29.31 //y=0.625 //x2=29.31 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=28.425 //y=1.59 //x2=28.34 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.425 //y=1.59 //x2=28.825 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.225 //y=1.59 //x2=29.31 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.225 //y=1.59 //x2=28.825 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=28.34 //y=1.505 //x2=28.34 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=28.34 //y=1.505 //x2=28.34 //y2=0.89
ends PM_TMRDFFSNQNX1\%noxref_37

subckt PM_TMRDFFSNQNX1\%noxref_38 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414739f //x=30.715 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=29.61 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=30.85 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=31.82 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=31.735 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=30.85 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=30.765 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=31.82 //y=0.625 //x2=31.82 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=31.82 //y=0.625 //x2=31.82 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.935 //y=0.54 //x2=30.85 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.935 //y=0.54 //x2=31.335 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=31.735 //y=0.54 //x2=31.82 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=31.735 //y=0.54 //x2=31.335 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=30.85 //y=1.08 //x2=30.85 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=30.85 //y=1.08 //x2=30.85 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=30.85 //y=0.91 //x2=30.85 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=30.85 //y=0.91 //x2=30.85 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=30.85 //y=0.625 //x2=30.85 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=30.85 //y=0.625 //x2=30.85 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.885 //y=0.995 //x2=29.8 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=30.765 //y=0.995 //x2=30.85 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=30.765 //y=0.995 //x2=29.885 //y2=0.995
ends PM_TMRDFFSNQNX1\%noxref_38

subckt PM_TMRDFFSNQNX1\%noxref_39 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=33.015 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=35.005 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=35.005 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=34.12 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=34.035 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=33.15 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.205 //y=1.59 //x2=34.12 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.205 //y=1.59 //x2=34.605 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.005 //y=1.59 //x2=35.09 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.005 //y=1.59 //x2=34.605 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.205 //y=0.54 //x2=34.12 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.205 //y=0.54 //x2=34.605 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.005 //y=0.54 //x2=35.09 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.005 //y=0.54 //x2=34.605 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=34.12 //y=1.505 //x2=34.12 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=34.12 //y=1.505 //x2=34.12 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=34.12 //y=0.625 //x2=34.12 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=34.12 //y=0.625 //x2=34.12 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=33.235 //y=1.59 //x2=33.15 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=33.235 //y=1.59 //x2=33.635 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.035 //y=1.59 //x2=34.12 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.035 //y=1.59 //x2=33.635 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=33.15 //y=1.505 //x2=33.15 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=33.15 //y=1.505 //x2=33.15 //y2=0.89
ends PM_TMRDFFSNQNX1\%noxref_39

subckt PM_TMRDFFSNQNX1\%noxref_40 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=35.525 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=34.42 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=35.66 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=36.63 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=36.545 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=35.66 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=35.575 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=36.63 //y=0.625 //x2=36.63 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=36.63 //y=0.625 //x2=36.63 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=35.745 //y=0.54 //x2=35.66 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.745 //y=0.54 //x2=36.145 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=36.545 //y=0.54 //x2=36.63 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=36.545 //y=0.54 //x2=36.145 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=35.66 //y=1.08 //x2=35.66 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=35.66 //y=1.08 //x2=35.66 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=35.66 //y=0.91 //x2=35.66 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=35.66 //y=0.91 //x2=35.66 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=35.66 //y=0.625 //x2=35.66 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=35.66 //y=0.625 //x2=35.66 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.695 //y=0.995 //x2=34.61 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=35.575 //y=0.995 //x2=35.66 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=35.575 //y=0.995 //x2=34.695 //y2=0.995
ends PM_TMRDFFSNQNX1\%noxref_40

subckt PM_TMRDFFSNQNX1\%noxref_41 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=37.93 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722223f //x=40.005 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=39.92 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=39.035 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=39.035 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=38.95 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=38.065 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=40.005 //y=0.615 //x2=40.005 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=40.005 //y=0.615 //x2=40.005 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=39.12 //y=0.53 //x2=39.035 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=39.12 //y=0.53 //x2=39.52 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=39.92 //y=0.53 //x2=40.005 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=39.92 //y=0.53 //x2=39.52 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=39.035 //y=1.495 //x2=39.035 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=39.035 //y=1.495 //x2=39.035 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=39.035 //y=0.615 //x2=39.035 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=39.035 //y=0.615 //x2=39.035 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=38.15 //y=1.58 //x2=38.065 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=38.15 //y=1.58 //x2=38.55 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=38.95 //y=1.58 //x2=39.035 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=38.95 //y=1.58 //x2=38.55 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=38.065 //y=1.495 //x2=38.065 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=38.065 //y=1.495 //x2=38.065 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_41

subckt PM_TMRDFFSNQNX1\%noxref_42 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.063352f //x=41.26 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=43.335 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=43.25 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=42.365 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=42.365 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=42.28 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=41.395 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=43.335 //y=0.615 //x2=43.335 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=43.335 //y=0.615 //x2=43.335 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=42.45 //y=0.53 //x2=42.365 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=42.45 //y=0.53 //x2=42.85 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=43.25 //y=0.53 //x2=43.335 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=43.25 //y=0.53 //x2=42.85 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=42.365 //y=1.495 //x2=42.365 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=42.365 //y=1.495 //x2=42.365 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=42.365 //y=0.615 //x2=42.365 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=42.365 //y=0.615 //x2=42.365 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=41.48 //y=1.58 //x2=41.395 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=41.48 //y=1.58 //x2=41.88 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=42.28 //y=1.58 //x2=42.365 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=42.28 //y=1.58 //x2=41.88 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=41.395 //y=1.495 //x2=41.395 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=41.395 //y=1.495 //x2=41.395 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_42

subckt PM_TMRDFFSNQNX1\%noxref_43 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=44.485 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=46.475 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=46.475 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=45.59 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=45.505 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=44.62 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=45.675 //y=1.59 //x2=45.59 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.675 //y=1.59 //x2=46.075 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.475 //y=1.59 //x2=46.56 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.475 //y=1.59 //x2=46.075 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=45.675 //y=0.54 //x2=45.59 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.675 //y=0.54 //x2=46.075 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.475 //y=0.54 //x2=46.56 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.475 //y=0.54 //x2=46.075 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=45.59 //y=1.505 //x2=45.59 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=45.59 //y=1.505 //x2=45.59 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=45.59 //y=0.625 //x2=45.59 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=45.59 //y=0.625 //x2=45.59 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.705 //y=1.59 //x2=44.62 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.705 //y=1.59 //x2=45.105 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=45.505 //y=1.59 //x2=45.59 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.505 //y=1.59 //x2=45.105 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=44.62 //y=1.505 //x2=44.62 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=44.62 //y=1.505 //x2=44.62 //y2=0.89
ends PM_TMRDFFSNQNX1\%noxref_43

subckt PM_TMRDFFSNQNX1\%noxref_44 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=46.995 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=45.89 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=47.13 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=48.1 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=48.015 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=47.13 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=47.045 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=48.1 //y=0.625 //x2=48.1 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=48.1 //y=0.625 //x2=48.1 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=47.215 //y=0.54 //x2=47.13 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=47.215 //y=0.54 //x2=47.615 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=48.015 //y=0.54 //x2=48.1 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=48.015 //y=0.54 //x2=47.615 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=47.13 //y=1.08 //x2=47.13 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=47.13 //y=1.08 //x2=47.13 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=47.13 //y=0.91 //x2=47.13 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=47.13 //y=0.91 //x2=47.13 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=47.13 //y=0.625 //x2=47.13 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=47.13 //y=0.625 //x2=47.13 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.165 //y=0.995 //x2=46.08 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=47.045 //y=0.995 //x2=47.13 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=47.045 //y=0.995 //x2=46.165 //y2=0.995
ends PM_TMRDFFSNQNX1\%noxref_44

subckt PM_TMRDFFSNQNX1\%noxref_45 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0633518f //x=49.4 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=51.475 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=51.39 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=50.505 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=50.505 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=50.42 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=49.535 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=51.475 //y=0.615 //x2=51.475 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=51.475 //y=0.615 //x2=51.475 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=50.59 //y=0.53 //x2=50.505 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.59 //y=0.53 //x2=50.99 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=51.39 //y=0.53 //x2=51.475 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=51.39 //y=0.53 //x2=50.99 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=50.505 //y=1.495 //x2=50.505 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=50.505 //y=1.495 //x2=50.505 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=50.505 //y=0.615 //x2=50.505 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=50.505 //y=0.615 //x2=50.505 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.62 //y=1.58 //x2=49.535 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.62 //y=1.58 //x2=50.02 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=50.42 //y=1.58 //x2=50.505 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.42 //y=1.58 //x2=50.02 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=49.535 //y=1.495 //x2=49.535 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=49.535 //y=1.495 //x2=49.535 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_45

subckt PM_TMRDFFSNQNX1\%noxref_46 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673195f //x=52.625 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=54.615 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=54.615 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=53.73 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=53.645 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=52.76 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.815 //y=1.59 //x2=53.73 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.815 //y=1.59 //x2=54.215 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.615 //y=1.59 //x2=54.7 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.615 //y=1.59 //x2=54.215 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.815 //y=0.54 //x2=53.73 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.815 //y=0.54 //x2=54.215 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.615 //y=0.54 //x2=54.7 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.615 //y=0.54 //x2=54.215 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=53.73 //y=1.505 //x2=53.73 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=53.73 //y=1.505 //x2=53.73 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=53.73 //y=0.625 //x2=53.73 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=53.73 //y=0.625 //x2=53.73 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=52.845 //y=1.59 //x2=52.76 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=52.845 //y=1.59 //x2=53.245 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.645 //y=1.59 //x2=53.73 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.645 //y=1.59 //x2=53.245 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=52.76 //y=1.505 //x2=52.76 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=52.76 //y=1.505 //x2=52.76 //y2=0.89
ends PM_TMRDFFSNQNX1\%noxref_46

subckt PM_TMRDFFSNQNX1\%noxref_47 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414739f //x=55.135 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=54.03 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=55.27 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=56.24 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=56.155 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=55.27 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=55.185 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=56.24 //y=0.625 //x2=56.24 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=56.24 //y=0.625 //x2=56.24 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=55.355 //y=0.54 //x2=55.27 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=55.355 //y=0.54 //x2=55.755 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=56.155 //y=0.54 //x2=56.24 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=56.155 //y=0.54 //x2=55.755 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=55.27 //y=1.08 //x2=55.27 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=55.27 //y=1.08 //x2=55.27 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=55.27 //y=0.91 //x2=55.27 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=55.27 //y=0.91 //x2=55.27 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=55.27 //y=0.625 //x2=55.27 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=55.27 //y=0.625 //x2=55.27 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.305 //y=0.995 //x2=54.22 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=55.185 //y=0.995 //x2=55.27 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=55.185 //y=0.995 //x2=54.305 //y2=0.995
ends PM_TMRDFFSNQNX1\%noxref_47

subckt PM_TMRDFFSNQNX1\%noxref_48 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=57.435 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=59.425 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=59.425 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=58.54 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=58.455 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=57.57 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.625 //y=1.59 //x2=58.54 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.625 //y=1.59 //x2=59.025 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.425 //y=1.59 //x2=59.51 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.425 //y=1.59 //x2=59.025 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.625 //y=0.54 //x2=58.54 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.625 //y=0.54 //x2=59.025 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.425 //y=0.54 //x2=59.51 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.425 //y=0.54 //x2=59.025 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=58.54 //y=1.505 //x2=58.54 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=58.54 //y=1.505 //x2=58.54 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=58.54 //y=0.625 //x2=58.54 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=58.54 //y=0.625 //x2=58.54 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=57.655 //y=1.59 //x2=57.57 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=57.655 //y=1.59 //x2=58.055 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.455 //y=1.59 //x2=58.54 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.455 //y=1.59 //x2=58.055 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=57.57 //y=1.505 //x2=57.57 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=57.57 //y=1.505 //x2=57.57 //y2=0.89
ends PM_TMRDFFSNQNX1\%noxref_48

subckt PM_TMRDFFSNQNX1\%noxref_49 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=59.945 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=58.84 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=60.08 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=61.05 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=60.965 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=60.08 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=59.995 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=61.05 //y=0.625 //x2=61.05 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=61.05 //y=0.625 //x2=61.05 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=60.165 //y=0.54 //x2=60.08 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.165 //y=0.54 //x2=60.565 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=60.965 //y=0.54 //x2=61.05 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.965 //y=0.54 //x2=60.565 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.08 //y=1.08 //x2=60.08 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=60.08 //y=1.08 //x2=60.08 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.08 //y=0.91 //x2=60.08 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=60.08 //y=0.91 //x2=60.08 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=60.08 //y=0.625 //x2=60.08 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=60.08 //y=0.625 //x2=60.08 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.115 //y=0.995 //x2=59.03 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=59.995 //y=0.995 //x2=60.08 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=59.995 //y=0.995 //x2=59.115 //y2=0.995
ends PM_TMRDFFSNQNX1\%noxref_49

subckt PM_TMRDFFSNQNX1\%noxref_50 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=62.35 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722223f //x=64.425 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=64.34 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=63.455 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=63.455 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=63.37 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=62.485 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=64.425 //y=0.615 //x2=64.425 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=64.425 //y=0.615 //x2=64.425 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63.54 //y=0.53 //x2=63.455 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63.54 //y=0.53 //x2=63.94 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=64.34 //y=0.53 //x2=64.425 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.34 //y=0.53 //x2=63.94 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=63.455 //y=1.495 //x2=63.455 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=63.455 //y=1.495 //x2=63.455 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=63.455 //y=0.615 //x2=63.455 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=63.455 //y=0.615 //x2=63.455 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=62.57 //y=1.58 //x2=62.485 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=62.57 //y=1.58 //x2=62.97 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63.37 //y=1.58 //x2=63.455 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63.37 //y=1.58 //x2=62.97 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=62.485 //y=1.495 //x2=62.485 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=62.485 //y=1.495 //x2=62.485 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_50

subckt PM_TMRDFFSNQNX1\%noxref_51 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632684f //x=65.68 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=67.755 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=67.67 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=66.785 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=66.785 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=66.7 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=65.815 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=67.755 //y=0.615 //x2=67.755 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=67.755 //y=0.615 //x2=67.755 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.87 //y=0.53 //x2=66.785 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=66.87 //y=0.53 //x2=67.27 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=67.67 //y=0.53 //x2=67.755 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=67.67 //y=0.53 //x2=67.27 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=66.785 //y=1.495 //x2=66.785 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=66.785 //y=1.495 //x2=66.785 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=66.785 //y=0.615 //x2=66.785 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=66.785 //y=0.615 //x2=66.785 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=65.9 //y=1.58 //x2=65.815 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=65.9 //y=1.58 //x2=66.3 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.7 //y=1.58 //x2=66.785 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=66.7 //y=1.58 //x2=66.3 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=65.815 //y=1.495 //x2=65.815 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=65.815 //y=1.495 //x2=65.815 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_51

subckt PM_TMRDFFSNQNX1\%noxref_52 ( 1 5 9 13 17 35 )
c51 ( 35 0 ) capacitor c=0.0680259f //x=68.905 //y=0.375
c52 ( 17 0 ) capacitor c=0.0180446f //x=70.895 //y=1.59
c53 ( 13 0 ) capacitor c=0.0155283f //x=70.895 //y=0.54
c54 ( 9 0 ) capacitor c=0.00678203f //x=70.01 //y=0.625
c55 ( 5 0 ) capacitor c=0.0164013f //x=69.925 //y=1.59
c56 ( 1 0 ) capacitor c=0.00696517f //x=69.04 //y=1.505
r57 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=70.095 //y=1.59 //x2=70.01 //y2=1.63
r58 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.095 //y=1.59 //x2=70.495 //y2=1.59
r59 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.895 //y=1.59 //x2=70.98 //y2=1.59
r60 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.895 //y=1.59 //x2=70.495 //y2=1.59
r61 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=70.095 //y=0.54 //x2=70.01 //y2=0.5
r62 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.095 //y=0.54 //x2=70.495 //y2=0.54
r63 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.895 //y=0.54 //x2=70.98 //y2=0.54
r64 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.895 //y=0.54 //x2=70.495 //y2=0.54
r65 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=70.01 //y=1.505 //x2=70.01 //y2=1.63
r66 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=70.01 //y=1.505 //x2=70.01 //y2=0.89
r67 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=70.01 //y=0.625 //x2=70.01 //y2=0.5
r68 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=70.01 //y=0.625 //x2=70.01 //y2=0.89
r69 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=69.125 //y=1.59 //x2=69.04 //y2=1.63
r70 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.125 //y=1.59 //x2=69.525 //y2=1.59
r71 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=69.925 //y=1.59 //x2=70.01 //y2=1.63
r72 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.925 //y=1.59 //x2=69.525 //y2=1.59
r73 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=69.04 //y=1.505 //x2=69.04 //y2=1.63
r74 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=69.04 //y=1.505 //x2=69.04 //y2=0.89
ends PM_TMRDFFSNQNX1\%noxref_52

subckt PM_TMRDFFSNQNX1\%noxref_53 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.042068f //x=71.415 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=70.31 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=71.55 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=72.52 //y=0.625
c56 ( 11 0 ) capacitor c=0.014695f //x=72.435 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=71.55 //y=0.625
c58 ( 1 0 ) capacitor c=0.0234159f //x=71.465 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=72.52 //y=0.625 //x2=72.52 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=72.52 //y=0.625 //x2=72.52 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=71.635 //y=0.54 //x2=71.55 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=71.635 //y=0.54 //x2=72.035 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=72.435 //y=0.54 //x2=72.52 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=72.435 //y=0.54 //x2=72.035 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=71.55 //y=1.08 //x2=71.55 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=71.55 //y=1.08 //x2=71.55 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=71.55 //y=0.91 //x2=71.55 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=71.55 //y=0.91 //x2=71.55 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=71.55 //y=0.625 //x2=71.55 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=71.55 //y=0.625 //x2=71.55 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.585 //y=0.995 //x2=70.5 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=71.465 //y=0.995 //x2=71.55 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=71.465 //y=0.995 //x2=70.585 //y2=0.995
ends PM_TMRDFFSNQNX1\%noxref_53

subckt PM_TMRDFFSNQNX1\%noxref_54 ( 1 5 9 10 13 17 29 )
c57 ( 29 0 ) capacitor c=0.0761166f //x=73.82 //y=0.365
c58 ( 17 0 ) capacitor c=0.0072249f //x=75.895 //y=0.615
c59 ( 13 0 ) capacitor c=0.0154142f //x=75.81 //y=0.53
c60 ( 10 0 ) capacitor c=0.00754234f //x=74.925 //y=1.495
c61 ( 9 0 ) capacitor c=0.006761f //x=74.925 //y=0.615
c62 ( 5 0 ) capacitor c=0.0213241f //x=74.84 //y=1.58
c63 ( 1 0 ) capacitor c=0.00492513f //x=73.955 //y=1.495
r64 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=75.895 //y=0.615 //x2=75.895 //y2=0.49
r65 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=75.895 //y=0.615 //x2=75.895 //y2=1.22
r66 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.01 //y=0.53 //x2=74.925 //y2=0.49
r67 (  14 29 ) resistor r=27.0374 //w=0.187 //l=0.395 //layer=li \
 //thickness=0.1 //x=75.01 //y=0.53 //x2=75.405 //y2=0.53
r68 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.81 //y=0.53 //x2=75.895 //y2=0.49
r69 (  13 29 ) resistor r=27.7219 //w=0.187 //l=0.405 //layer=li \
 //thickness=0.1 //x=75.81 //y=0.53 //x2=75.405 //y2=0.53
r70 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=74.925 //y=1.495 //x2=74.925 //y2=1.62
r71 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=74.925 //y=1.495 //x2=74.925 //y2=0.88
r72 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=74.925 //y=0.615 //x2=74.925 //y2=0.49
r73 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=74.925 //y=0.615 //x2=74.925 //y2=0.88
r74 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=74.04 //y=1.58 //x2=73.955 //y2=1.62
r75 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=74.04 //y=1.58 //x2=74.44 //y2=1.58
r76 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=74.84 //y=1.58 //x2=74.925 //y2=1.62
r77 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=74.84 //y=1.58 //x2=74.44 //y2=1.58
r78 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=73.955 //y=1.495 //x2=73.955 //y2=1.62
r79 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=73.955 //y=1.495 //x2=73.955 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_54

subckt PM_TMRDFFSNQNX1\%noxref_55 ( 1 5 9 10 13 17 29 )
c55 ( 29 0 ) capacitor c=0.0723103f //x=77.15 //y=0.365
c56 ( 17 0 ) capacitor c=0.0072249f //x=79.225 //y=0.615
c57 ( 13 0 ) capacitor c=0.0155051f //x=79.14 //y=0.53
c58 ( 10 0 ) capacitor c=0.00907139f //x=78.255 //y=1.495
c59 ( 9 0 ) capacitor c=0.006761f //x=78.255 //y=0.615
c60 ( 5 0 ) capacitor c=0.019003f //x=78.17 //y=1.58
c61 ( 1 0 ) capacitor c=0.00885385f //x=77.285 //y=1.495
r62 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=79.225 //y=0.615 //x2=79.225 //y2=0.49
r63 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=79.225 //y=0.615 //x2=79.225 //y2=1.22
r64 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.34 //y=0.53 //x2=78.255 //y2=0.49
r65 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.34 //y=0.53 //x2=78.74 //y2=0.53
r66 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=79.14 //y=0.53 //x2=79.225 //y2=0.49
r67 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=79.14 //y=0.53 //x2=78.74 //y2=0.53
r68 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=78.255 //y=1.495 //x2=78.255 //y2=1.62
r69 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=78.255 //y=1.495 //x2=78.255 //y2=0.88
r70 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=78.255 //y=0.615 //x2=78.255 //y2=0.49
r71 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=78.255 //y=0.615 //x2=78.255 //y2=0.88
r72 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=77.37 //y=1.58 //x2=77.285 //y2=1.62
r73 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=77.37 //y=1.58 //x2=77.77 //y2=1.58
r74 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.17 //y=1.58 //x2=78.255 //y2=1.62
r75 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.17 //y=1.58 //x2=77.77 //y2=1.58
r76 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=77.285 //y=1.495 //x2=77.285 //y2=1.62
r77 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=77.285 //y=1.495 //x2=77.285 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_55

subckt PM_TMRDFFSNQNX1\%noxref_56 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.0643725f //x=80.48 //y=0.365
c54 ( 17 0 ) capacitor c=0.00722228f //x=82.555 //y=0.615
c55 ( 13 0 ) capacitor c=0.0141607f //x=82.47 //y=0.53
c56 ( 10 0 ) capacitor c=0.00712138f //x=81.585 //y=1.495
c57 ( 9 0 ) capacitor c=0.006761f //x=81.585 //y=0.615
c58 ( 5 0 ) capacitor c=0.0233454f //x=81.5 //y=1.58
c59 ( 1 0 ) capacitor c=0.00481264f //x=80.615 //y=1.495
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=82.555 //y=0.615 //x2=82.555 //y2=0.49
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=82.555 //y=0.615 //x2=82.555 //y2=0.88
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=81.67 //y=0.53 //x2=81.585 //y2=0.49
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=81.67 //y=0.53 //x2=82.07 //y2=0.53
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=82.47 //y=0.53 //x2=82.555 //y2=0.49
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=82.47 //y=0.53 //x2=82.07 //y2=0.53
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=81.585 //y=1.495 //x2=81.585 //y2=1.62
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=81.585 //y=1.495 //x2=81.585 //y2=0.88
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=81.585 //y=0.615 //x2=81.585 //y2=0.49
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=81.585 //y=0.615 //x2=81.585 //y2=0.88
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=80.7 //y=1.58 //x2=80.615 //y2=1.62
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=80.7 //y=1.58 //x2=81.1 //y2=1.58
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=81.5 //y=1.58 //x2=81.585 //y2=1.62
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=81.5 //y=1.58 //x2=81.1 //y2=1.58
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=80.615 //y=1.495 //x2=80.615 //y2=1.62
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=80.615 //y=1.495 //x2=80.615 //y2=0.88
ends PM_TMRDFFSNQNX1\%noxref_56

