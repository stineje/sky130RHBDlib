* SPICE3 file created from XOR2X1.ext - technology: sky130A

.subckt XOR2X1 Y A B VDD VSS
X0 a_807_990 B VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.00336 ps=2.736 w=2 l=0.15 M=2
X1 a_185_209 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X2 VSS A a_556_101 VSS sky130_fd_pr__nfet_01v8 ad=0.0026398 pd=1.934 as=0 ps=0 w=3 l=0.15
X3 a_185_209 A VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X4 a_575_1051 a_807_990 Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.00116 ps=9.16 w=2 l=0.15 M=2
X5 Y a_185_209 a_1222_101 VSS sky130_fd_pr__nfet_01v8 ad=0.003582 pd=3.14 as=0 ps=0 w=3 l=0.15
X6 a_1241_1051 B VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X7 a_807_990 B VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X8 a_1241_1051 a_185_209 Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X9 Y B a_556_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X10 VDD A a_575_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X11 VSS a_807_990 a_1222_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 a_807_990 B 2.21f
C1 VDD VSS 4.20f
.ends
