** sch_path: /home/rjridle/OpenRadHardSCL/sky130A/libs.tech/xschem/sky130_stdcells/nand2_1.sym
.subckt nand2_1

.ends
.end
