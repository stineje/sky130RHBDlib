magic
tech sky130A
magscale 1 2
timestamp 1648062678
<< nmos >>
rect 162 215 192 276
tri 57 185 87 215 se
rect 87 185 192 215
rect 57 91 87 185
tri 87 169 103 185 nw
tri 146 169 162 185 ne
tri 87 91 103 107 sw
tri 146 91 162 107 se
rect 162 91 192 185
tri 57 61 87 91 ne
rect 87 61 162 91
tri 162 61 192 91 nw
<< ndiff >>
rect 0 260 162 276
rect 0 226 10 260
rect 44 226 107 260
rect 141 226 162 260
rect 0 215 162 226
rect 192 260 248 276
rect 192 226 204 260
rect 238 226 248 260
rect 0 188 57 215
rect 0 154 10 188
rect 44 154 57 188
tri 57 185 87 215 nw
rect 0 120 57 154
rect 0 86 10 120
rect 44 86 57 120
tri 87 169 103 185 se
rect 103 169 146 185
tri 146 169 162 185 sw
rect 87 141 162 169
rect 87 107 108 141
rect 142 107 162 141
tri 87 91 103 107 ne
rect 103 91 146 107
tri 146 91 162 107 nw
rect 0 61 57 86
tri 57 61 87 91 sw
tri 162 61 192 91 se
rect 192 61 248 226
rect 0 50 248 61
rect 0 16 10 50
rect 44 16 107 50
rect 141 16 204 50
rect 238 16 248 50
rect 0 0 248 16
<< ndiffc >>
rect 10 226 44 260
rect 107 226 141 260
rect 204 226 238 260
rect 10 154 44 188
rect 10 86 44 120
rect 108 107 142 141
rect 10 16 44 50
rect 107 16 141 50
rect 204 16 238 50
<< poly >>
rect 162 276 192 302
<< locali >>
rect 10 260 44 276
rect 204 260 238 276
rect 44 226 107 260
rect 141 226 204 260
rect 10 188 44 226
rect 204 210 238 226
rect 10 120 44 154
rect 108 141 142 157
rect 108 91 142 107
rect 10 50 44 86
rect 204 50 238 66
rect 44 16 107 50
rect 141 16 204 50
rect 10 0 44 16
rect 204 0 238 16
<< end >>
