* SPICE3 file created from XNOR2X1.ext - technology: sky130A

.subckt XNOR2X1 Y A B VDD GND
X0 GND A xnor2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 GND B xnor2x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X2 VDD A xnor2x1_pcell_0/a_761_1330# VDD pshort w=2 l=0.15
X3 Y xnor2x1_pcell_0/m1_315_501# xnor2x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X4 Y B xnor2x1_pcell_0/a_761_1330# VDD pshort w=2 l=0.15
X5 Y xnor2x1_pcell_0/a_806_382# xnor2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X6 VDD xnor2x1_pcell_0/a_806_382# xnor2x1_pcell_0/a_1427_1330# VDD pshort w=2 l=0.15
X7 Y xnor2x1_pcell_0/m1_315_501# xnor2x1_pcell_0/a_1427_1330# VDD pshort w=2 l=0.15
X8 xnor2x1_pcell_0/m1_315_501# A GND GND nshort w=3 l=0.15
X9 VDD A xnor2x1_pcell_0/m1_315_501# VDD pshort w=2 l=0.15
X10 xnor2x1_pcell_0/a_806_382# B xnor2x1_pcell_0/li1_M1_contact_2/VSUBS xnor2x1_pcell_0/li1_M1_contact_2/VSUBS nshort w=3 l=0.15
X11 VDD B xnor2x1_pcell_0/a_806_382# VDD pshort w=2 l=0.15
C0 xnor2x1_pcell_0/a_806_382# B 2.06fF
C1 VDD xnor2x1_pcell_0/li1_M1_contact_2/VSUBS 14.21fF
.ends
