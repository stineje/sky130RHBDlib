// File: TMRDFFRNQNX1.spi.TMRDFFRNQNX1.pxi
// Created: Tue Oct 15 15:52:03 2024
// 
simulator lang=spectre
x_PM_TMRDFFRNQNX1\%GND ( GND N_GND_c_23_p N_GND_c_95_p N_GND_c_1_p \
 N_GND_c_24_p N_GND_c_25_p N_GND_c_71_p N_GND_c_32_p N_GND_c_39_p N_GND_c_47_p \
 N_GND_c_54_p N_GND_c_74_p N_GND_c_81_p N_GND_c_105_p N_GND_c_112_p \
 N_GND_c_190_p N_GND_c_197_p N_GND_c_150_p N_GND_c_157_p N_GND_c_120_p \
 N_GND_c_127_p N_GND_c_134_p N_GND_c_141_p N_GND_c_160_p N_GND_c_167_p \
 N_GND_c_173_p N_GND_c_180_p N_GND_c_293_p N_GND_c_294_p N_GND_c_227_p \
 N_GND_c_234_p N_GND_c_303_p N_GND_c_304_p N_GND_c_305_p N_GND_c_306_p \
 N_GND_c_237_p N_GND_c_244_p N_GND_c_342_p N_GND_c_349_p N_GND_c_388_p \
 N_GND_c_395_p N_GND_c_398_p N_GND_c_404_p N_GND_c_457_p N_GND_c_2_p \
 N_GND_c_3_p N_GND_c_4_p N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p N_GND_c_8_p \
 N_GND_c_9_p N_GND_c_10_p N_GND_c_11_p N_GND_c_12_p N_GND_c_13_p N_GND_c_14_p \
 N_GND_c_15_p N_GND_c_16_p N_GND_c_17_p N_GND_c_18_p N_GND_c_19_p N_GND_c_20_p \
 N_GND_c_21_p N_GND_c_22_p N_GND_M0_noxref_d N_GND_M3_noxref_d \
 N_GND_M6_noxref_d N_GND_M8_noxref_d N_GND_M11_noxref_d N_GND_M14_noxref_d \
 N_GND_M16_noxref_d N_GND_M19_noxref_d N_GND_M22_noxref_d N_GND_M24_noxref_d \
 N_GND_M27_noxref_d N_GND_M30_noxref_d N_GND_M32_noxref_d N_GND_M35_noxref_d \
 N_GND_M38_noxref_d N_GND_M40_noxref_d N_GND_M43_noxref_d N_GND_M46_noxref_d \
 N_GND_M48_noxref_d N_GND_M50_noxref_d N_GND_M52_noxref_d )  \
 PM_TMRDFFRNQNX1\%GND
x_PM_TMRDFFRNQNX1\%VDD ( VDD N_VDD_c_1015_p N_VDD_c_992_n N_VDD_c_1089_p \
 N_VDD_c_1090_p N_VDD_c_1033_p N_VDD_c_1100_p N_VDD_c_1480_p N_VDD_c_1016_p \
 N_VDD_c_1017_p N_VDD_c_1023_p N_VDD_c_1027_p N_VDD_c_1483_p N_VDD_c_1031_p \
 N_VDD_c_1059_p N_VDD_c_1485_p N_VDD_c_1486_p N_VDD_c_1071_p N_VDD_c_1156_p \
 N_VDD_c_1162_p N_VDD_c_1166_p N_VDD_c_1498_p N_VDD_c_1113_p N_VDD_c_1171_p \
 N_VDD_c_1177_p N_VDD_c_1181_p N_VDD_c_1501_p N_VDD_c_1185_p N_VDD_c_1202_p \
 N_VDD_c_1503_p N_VDD_c_1504_p N_VDD_c_1315_p N_VDD_c_1316_p N_VDD_c_1259_p \
 N_VDD_c_1326_p N_VDD_c_1516_p N_VDD_c_1242_p N_VDD_c_1243_p N_VDD_c_1249_p \
 N_VDD_c_1253_p N_VDD_c_1519_p N_VDD_c_1257_p N_VDD_c_1285_p N_VDD_c_1521_p \
 N_VDD_c_1522_p N_VDD_c_1297_p N_VDD_c_1414_p N_VDD_c_1420_p N_VDD_c_1424_p \
 N_VDD_c_1534_p N_VDD_c_1339_p N_VDD_c_1364_p N_VDD_c_1370_p N_VDD_c_1374_p \
 N_VDD_c_1537_p N_VDD_c_1378_p N_VDD_c_1438_p N_VDD_c_1539_p N_VDD_c_1540_p \
 N_VDD_c_1541_p N_VDD_c_1596_p N_VDD_c_1612_p N_VDD_c_1551_p N_VDD_c_1552_p \
 N_VDD_c_1553_p N_VDD_c_1474_p N_VDD_c_1688_p N_VDD_c_1554_p N_VDD_c_1555_p \
 N_VDD_c_1556_p N_VDD_c_1771_p N_VDD_c_1557_p N_VDD_c_1558_p N_VDD_c_1559_p \
 N_VDD_c_1600_p N_VDD_c_1692_p N_VDD_c_1706_p N_VDD_c_1707_p N_VDD_c_1629_p \
 N_VDD_c_1696_p N_VDD_c_1755_p N_VDD_c_1715_p N_VDD_c_1716_p N_VDD_c_1717_p \
 N_VDD_c_1780_p N_VDD_c_1825_p N_VDD_c_1820_p N_VDD_c_1978_p N_VDD_c_1999_p \
 N_VDD_c_1900_p N_VDD_c_993_n N_VDD_c_994_n N_VDD_c_995_n N_VDD_c_996_n \
 N_VDD_c_997_n N_VDD_c_998_n N_VDD_c_999_n N_VDD_c_1000_n N_VDD_c_1001_n \
 N_VDD_c_1002_n N_VDD_c_1003_n N_VDD_c_1004_n N_VDD_c_1005_n N_VDD_c_1006_n \
 N_VDD_c_1007_n N_VDD_c_1008_n N_VDD_c_1009_n N_VDD_c_1010_n N_VDD_c_1011_n \
 N_VDD_c_1012_n N_VDD_c_1013_n N_VDD_M54_noxref_s N_VDD_M55_noxref_d \
 N_VDD_M57_noxref_d N_VDD_M59_noxref_d N_VDD_M60_noxref_s N_VDD_M61_noxref_d \
 N_VDD_M63_noxref_d N_VDD_M65_noxref_d N_VDD_M66_noxref_s N_VDD_M67_noxref_d \
 N_VDD_M69_noxref_d N_VDD_M70_noxref_s N_VDD_M71_noxref_d N_VDD_M73_noxref_d \
 N_VDD_M75_noxref_d N_VDD_M76_noxref_s N_VDD_M77_noxref_d N_VDD_M79_noxref_d \
 N_VDD_M81_noxref_d N_VDD_M82_noxref_s N_VDD_M83_noxref_d N_VDD_M85_noxref_d \
 N_VDD_M86_noxref_s N_VDD_M87_noxref_d N_VDD_M89_noxref_d N_VDD_M91_noxref_d \
 N_VDD_M92_noxref_s N_VDD_M93_noxref_d N_VDD_M95_noxref_d N_VDD_M97_noxref_d \
 N_VDD_M98_noxref_s N_VDD_M99_noxref_d N_VDD_M101_noxref_d N_VDD_M102_noxref_s \
 N_VDD_M103_noxref_d N_VDD_M105_noxref_d N_VDD_M107_noxref_d \
 N_VDD_M108_noxref_s N_VDD_M109_noxref_d N_VDD_M111_noxref_d \
 N_VDD_M113_noxref_d N_VDD_M114_noxref_s N_VDD_M115_noxref_d \
 N_VDD_M117_noxref_d N_VDD_M118_noxref_s N_VDD_M119_noxref_d \
 N_VDD_M121_noxref_d N_VDD_M123_noxref_d N_VDD_M124_noxref_s \
 N_VDD_M125_noxref_d N_VDD_M127_noxref_d N_VDD_M129_noxref_d \
 N_VDD_M130_noxref_s N_VDD_M131_noxref_d N_VDD_M133_noxref_d \
 N_VDD_M134_noxref_s N_VDD_M135_noxref_d N_VDD_M137_noxref_d \
 N_VDD_M139_noxref_d N_VDD_M140_noxref_s N_VDD_M141_noxref_d \
 N_VDD_M143_noxref_d N_VDD_M145_noxref_d N_VDD_M146_noxref_s \
 N_VDD_M147_noxref_d N_VDD_M149_noxref_d N_VDD_M150_noxref_s \
 N_VDD_M151_noxref_d N_VDD_M153_noxref_d )  PM_TMRDFFRNQNX1\%VDD
x_PM_TMRDFFRNQNX1\%noxref_3 ( N_noxref_3_c_2093_n N_noxref_3_c_2097_n \
 N_noxref_3_c_2098_n N_noxref_3_c_2169_p N_noxref_3_c_2099_n \
 N_noxref_3_c_2114_n N_noxref_3_c_2118_n N_noxref_3_c_2120_n \
 N_noxref_3_c_2124_n N_noxref_3_c_2100_n N_noxref_3_c_2281_p \
 N_noxref_3_c_2128_n N_noxref_3_c_2101_n N_noxref_3_c_2249_p \
 N_noxref_3_c_2291_p N_noxref_3_M2_noxref_g N_noxref_3_M6_noxref_g \
 N_noxref_3_M58_noxref_g N_noxref_3_M59_noxref_g N_noxref_3_M66_noxref_g \
 N_noxref_3_M67_noxref_g N_noxref_3_c_2194_p N_noxref_3_c_2195_p \
 N_noxref_3_c_2196_p N_noxref_3_c_2197_p N_noxref_3_c_2177_p \
 N_noxref_3_c_2199_p N_noxref_3_c_2178_p N_noxref_3_c_2102_n \
 N_noxref_3_c_2104_n N_noxref_3_c_2105_n N_noxref_3_c_2106_n \
 N_noxref_3_c_2107_n N_noxref_3_c_2108_n N_noxref_3_c_2109_n \
 N_noxref_3_c_2111_n N_noxref_3_c_2183_p N_noxref_3_c_2184_p \
 N_noxref_3_c_2176_p N_noxref_3_c_2140_n N_noxref_3_M5_noxref_d \
 N_noxref_3_M60_noxref_d N_noxref_3_M62_noxref_d N_noxref_3_M64_noxref_d )  \
 PM_TMRDFFRNQNX1\%noxref_3
x_PM_TMRDFFRNQNX1\%noxref_4 ( N_noxref_4_c_2343_n N_noxref_4_c_2391_n \
 N_noxref_4_c_2360_n N_noxref_4_c_2364_n N_noxref_4_c_2366_n \
 N_noxref_4_c_2344_n N_noxref_4_c_2472_p N_noxref_4_c_2345_n \
 N_noxref_4_c_2346_n N_noxref_4_c_2425_p N_noxref_4_M8_noxref_g \
 N_noxref_4_M70_noxref_g N_noxref_4_M71_noxref_g N_noxref_4_c_2347_n \
 N_noxref_4_c_2349_n N_noxref_4_c_2350_n N_noxref_4_c_2351_n \
 N_noxref_4_c_2352_n N_noxref_4_c_2353_n N_noxref_4_c_2354_n \
 N_noxref_4_c_2356_n N_noxref_4_c_2416_p N_noxref_4_c_2378_n \
 N_noxref_4_M7_noxref_d N_noxref_4_M66_noxref_d N_noxref_4_M68_noxref_d )  \
 PM_TMRDFFRNQNX1\%noxref_4
x_PM_TMRDFFRNQNX1\%noxref_5 ( N_noxref_5_c_2568_n N_noxref_5_c_2569_n \
 N_noxref_5_c_2495_n N_noxref_5_c_2576_n N_noxref_5_c_2520_n \
 N_noxref_5_c_2524_n N_noxref_5_c_2526_n N_noxref_5_c_2530_n \
 N_noxref_5_c_2496_n N_noxref_5_c_2583_n N_noxref_5_c_2534_n \
 N_noxref_5_c_2497_n N_noxref_5_c_2498_n N_noxref_5_c_2670_p \
 N_noxref_5_c_2592_n N_noxref_5_M3_noxref_g N_noxref_5_M11_noxref_g \
 N_noxref_5_M60_noxref_g N_noxref_5_M61_noxref_g N_noxref_5_M76_noxref_g \
 N_noxref_5_M77_noxref_g N_noxref_5_c_2499_n N_noxref_5_c_2501_n \
 N_noxref_5_c_2502_n N_noxref_5_c_2503_n N_noxref_5_c_2504_n \
 N_noxref_5_c_2505_n N_noxref_5_c_2506_n N_noxref_5_c_2508_n \
 N_noxref_5_c_2597_n N_noxref_5_c_2549_n N_noxref_5_c_2509_n \
 N_noxref_5_c_2511_n N_noxref_5_c_2512_n N_noxref_5_c_2513_n \
 N_noxref_5_c_2514_n N_noxref_5_c_2515_n N_noxref_5_c_2516_n \
 N_noxref_5_c_2518_n N_noxref_5_c_2630_p N_noxref_5_c_2551_n \
 N_noxref_5_M2_noxref_d N_noxref_5_M54_noxref_d N_noxref_5_M56_noxref_d \
 N_noxref_5_M58_noxref_d )  PM_TMRDFFRNQNX1\%noxref_5
x_PM_TMRDFFRNQNX1\%noxref_6 ( N_noxref_6_c_2748_n N_noxref_6_c_2749_n \
 N_noxref_6_c_2787_n N_noxref_6_c_2891_n N_noxref_6_c_2788_n \
 N_noxref_6_c_2789_n N_noxref_6_c_2790_n N_noxref_6_c_2791_n \
 N_noxref_6_c_2975_p N_noxref_6_c_2792_n N_noxref_6_c_2750_n \
 N_noxref_6_c_2893_n N_noxref_6_c_2751_n N_noxref_6_c_2798_n \
 N_noxref_6_c_2802_n N_noxref_6_c_2804_n N_noxref_6_c_2808_n \
 N_noxref_6_c_2753_n N_noxref_6_c_3060_p N_noxref_6_c_2812_n \
 N_noxref_6_c_2813_n N_noxref_6_c_2817_n N_noxref_6_c_2819_n \
 N_noxref_6_c_2823_n N_noxref_6_c_2754_n N_noxref_6_c_3064_p \
 N_noxref_6_c_2827_n N_noxref_6_c_2755_n N_noxref_6_c_3016_p \
 N_noxref_6_c_2756_n N_noxref_6_c_3018_p N_noxref_6_c_3076_p \
 N_noxref_6_c_3098_p N_noxref_6_c_3121_p N_noxref_6_M0_noxref_g \
 N_noxref_6_M7_noxref_g N_noxref_6_M14_noxref_g N_noxref_6_M15_noxref_g \
 N_noxref_6_M54_noxref_g N_noxref_6_M55_noxref_g N_noxref_6_M68_noxref_g \
 N_noxref_6_M69_noxref_g N_noxref_6_M82_noxref_g N_noxref_6_M83_noxref_g \
 N_noxref_6_M84_noxref_g N_noxref_6_M85_noxref_g N_noxref_6_c_2758_n \
 N_noxref_6_c_2760_n N_noxref_6_c_2761_n N_noxref_6_c_2762_n \
 N_noxref_6_c_2763_n N_noxref_6_c_2764_n N_noxref_6_c_2765_n \
 N_noxref_6_c_2767_n N_noxref_6_c_2973_n N_noxref_6_c_2851_n \
 N_noxref_6_c_2902_n N_noxref_6_c_2905_n N_noxref_6_c_2907_n \
 N_noxref_6_c_2937_n N_noxref_6_c_2939_n N_noxref_6_c_2940_n \
 N_noxref_6_c_2910_n N_noxref_6_c_2911_n N_noxref_6_c_2768_n \
 N_noxref_6_c_2770_n N_noxref_6_c_2771_n N_noxref_6_c_2772_n \
 N_noxref_6_c_2773_n N_noxref_6_c_2774_n N_noxref_6_c_2775_n \
 N_noxref_6_c_2777_n N_noxref_6_c_3161_p N_noxref_6_c_3162_p \
 N_noxref_6_c_3163_p N_noxref_6_c_3019_p N_noxref_6_c_3164_p \
 N_noxref_6_c_3069_p N_noxref_6_c_3166_p N_noxref_6_c_3131_p \
 N_noxref_6_c_2912_n N_noxref_6_c_2946_n N_noxref_6_c_2914_n \
 N_noxref_6_c_2853_n N_noxref_6_c_3070_p N_noxref_6_c_3139_p \
 N_noxref_6_c_3021_p N_noxref_6_M10_noxref_d N_noxref_6_M13_noxref_d \
 N_noxref_6_M70_noxref_d N_noxref_6_M72_noxref_d N_noxref_6_M74_noxref_d \
 N_noxref_6_M76_noxref_d N_noxref_6_M78_noxref_d N_noxref_6_M80_noxref_d )  \
 PM_TMRDFFRNQNX1\%noxref_6
x_PM_TMRDFFRNQNX1\%noxref_7 ( N_noxref_7_c_3298_p N_noxref_7_c_3314_p \
 N_noxref_7_c_3290_p N_noxref_7_c_3303_p N_noxref_7_c_3233_n \
 N_noxref_7_c_3248_n N_noxref_7_c_3252_n N_noxref_7_c_3254_n \
 N_noxref_7_c_3258_n N_noxref_7_c_3234_n N_noxref_7_c_3417_p \
 N_noxref_7_c_3262_n N_noxref_7_c_3235_n N_noxref_7_c_3385_p \
 N_noxref_7_c_3426_p N_noxref_7_M18_noxref_g N_noxref_7_M22_noxref_g \
 N_noxref_7_M90_noxref_g N_noxref_7_M91_noxref_g N_noxref_7_M98_noxref_g \
 N_noxref_7_M99_noxref_g N_noxref_7_c_3327_p N_noxref_7_c_3328_p \
 N_noxref_7_c_3329_p N_noxref_7_c_3330_p N_noxref_7_c_3311_p \
 N_noxref_7_c_3332_p N_noxref_7_c_3312_p N_noxref_7_c_3236_n \
 N_noxref_7_c_3238_n N_noxref_7_c_3239_n N_noxref_7_c_3240_n \
 N_noxref_7_c_3241_n N_noxref_7_c_3242_n N_noxref_7_c_3243_n \
 N_noxref_7_c_3245_n N_noxref_7_c_3316_p N_noxref_7_c_3317_p \
 N_noxref_7_c_3310_p N_noxref_7_c_3274_n N_noxref_7_M21_noxref_d \
 N_noxref_7_M92_noxref_d N_noxref_7_M94_noxref_d N_noxref_7_M96_noxref_d )  \
 PM_TMRDFFRNQNX1\%noxref_7
x_PM_TMRDFFRNQNX1\%noxref_8 ( N_noxref_8_c_3535_p N_noxref_8_c_3527_n \
 N_noxref_8_c_3496_n N_noxref_8_c_3500_n N_noxref_8_c_3502_n \
 N_noxref_8_c_3480_n N_noxref_8_c_3606_p N_noxref_8_c_3481_n \
 N_noxref_8_c_3482_n N_noxref_8_c_3561_p N_noxref_8_M24_noxref_g \
 N_noxref_8_M102_noxref_g N_noxref_8_M103_noxref_g N_noxref_8_c_3483_n \
 N_noxref_8_c_3485_n N_noxref_8_c_3486_n N_noxref_8_c_3487_n \
 N_noxref_8_c_3488_n N_noxref_8_c_3489_n N_noxref_8_c_3490_n \
 N_noxref_8_c_3492_n N_noxref_8_c_3552_p N_noxref_8_c_3514_n \
 N_noxref_8_M23_noxref_d N_noxref_8_M98_noxref_d N_noxref_8_M100_noxref_d )  \
 PM_TMRDFFRNQNX1\%noxref_8
x_PM_TMRDFFRNQNX1\%noxref_9 ( N_noxref_9_c_3705_n N_noxref_9_c_3706_n \
 N_noxref_9_c_3708_n N_noxref_9_c_3713_n N_noxref_9_c_3657_n \
 N_noxref_9_c_3661_n N_noxref_9_c_3663_n N_noxref_9_c_3667_n \
 N_noxref_9_c_3633_n N_noxref_9_c_3824_p N_noxref_9_c_3671_n \
 N_noxref_9_c_3634_n N_noxref_9_c_3635_n N_noxref_9_c_3808_p \
 N_noxref_9_c_3728_n N_noxref_9_M19_noxref_g N_noxref_9_M27_noxref_g \
 N_noxref_9_M92_noxref_g N_noxref_9_M93_noxref_g N_noxref_9_M108_noxref_g \
 N_noxref_9_M109_noxref_g N_noxref_9_c_3636_n N_noxref_9_c_3638_n \
 N_noxref_9_c_3639_n N_noxref_9_c_3640_n N_noxref_9_c_3641_n \
 N_noxref_9_c_3642_n N_noxref_9_c_3643_n N_noxref_9_c_3645_n \
 N_noxref_9_c_3733_n N_noxref_9_c_3686_n N_noxref_9_c_3646_n \
 N_noxref_9_c_3648_n N_noxref_9_c_3649_n N_noxref_9_c_3650_n \
 N_noxref_9_c_3651_n N_noxref_9_c_3652_n N_noxref_9_c_3653_n \
 N_noxref_9_c_3655_n N_noxref_9_c_3751_p N_noxref_9_c_3688_n \
 N_noxref_9_M18_noxref_d N_noxref_9_M86_noxref_d N_noxref_9_M88_noxref_d \
 N_noxref_9_M90_noxref_d )  PM_TMRDFFRNQNX1\%noxref_9
x_PM_TMRDFFRNQNX1\%noxref_10 ( N_noxref_10_c_3951_p N_noxref_10_c_3946_n \
 N_noxref_10_c_3908_n N_noxref_10_c_3912_n N_noxref_10_c_3914_n \
 N_noxref_10_c_3918_n N_noxref_10_c_3895_n N_noxref_10_c_3989_p \
 N_noxref_10_c_3922_n N_noxref_10_c_3896_n N_noxref_10_c_3999_p \
 N_noxref_10_c_4009_p N_noxref_10_M30_noxref_g N_noxref_10_M114_noxref_g \
 N_noxref_10_M115_noxref_g N_noxref_10_c_3897_n N_noxref_10_c_3899_n \
 N_noxref_10_c_3900_n N_noxref_10_c_3901_n N_noxref_10_c_3902_n \
 N_noxref_10_c_3903_n N_noxref_10_c_3904_n N_noxref_10_c_3906_n \
 N_noxref_10_c_3930_n N_noxref_10_M29_noxref_d N_noxref_10_M108_noxref_d \
 N_noxref_10_M110_noxref_d N_noxref_10_M112_noxref_d )  \
 PM_TMRDFFRNQNX1\%noxref_10
x_PM_TMRDFFRNQNX1\%noxref_11 ( N_noxref_11_c_4075_n N_noxref_11_c_4077_n \
 N_noxref_11_c_4078_n N_noxref_11_c_4144_n N_noxref_11_c_4079_n \
 N_noxref_11_c_4081_n N_noxref_11_c_4058_n N_noxref_11_c_4146_n \
 N_noxref_11_c_4059_n N_noxref_11_c_4087_n N_noxref_11_c_4091_n \
 N_noxref_11_c_4093_n N_noxref_11_c_4097_n N_noxref_11_c_4061_n \
 N_noxref_11_c_4321_p N_noxref_11_c_4101_n N_noxref_11_c_4228_n \
 N_noxref_11_c_4062_n N_noxref_11_c_4280_p N_noxref_11_c_4331_p \
 N_noxref_11_M16_noxref_g N_noxref_11_M23_noxref_g N_noxref_11_M31_noxref_g \
 N_noxref_11_M86_noxref_g N_noxref_11_M87_noxref_g N_noxref_11_M100_noxref_g \
 N_noxref_11_M101_noxref_g N_noxref_11_M116_noxref_g N_noxref_11_M117_noxref_g \
 N_noxref_11_c_4064_n N_noxref_11_c_4066_n N_noxref_11_c_4067_n \
 N_noxref_11_c_4068_n N_noxref_11_c_4069_n N_noxref_11_c_4070_n \
 N_noxref_11_c_4071_n N_noxref_11_c_4073_n N_noxref_11_c_4222_n \
 N_noxref_11_c_4118_n N_noxref_11_c_4155_n N_noxref_11_c_4158_n \
 N_noxref_11_c_4160_n N_noxref_11_c_4190_n N_noxref_11_c_4192_n \
 N_noxref_11_c_4193_n N_noxref_11_c_4163_n N_noxref_11_c_4164_n \
 N_noxref_11_c_4237_n N_noxref_11_c_4240_n N_noxref_11_c_4242_n \
 N_noxref_11_c_4281_p N_noxref_11_c_4377_p N_noxref_11_c_4325_p \
 N_noxref_11_c_4245_n N_noxref_11_c_4246_n N_noxref_11_c_4165_n \
 N_noxref_11_c_4199_n N_noxref_11_c_4167_n N_noxref_11_c_4247_n \
 N_noxref_11_c_4371_p N_noxref_11_c_4249_n N_noxref_11_M26_noxref_d \
 N_noxref_11_M102_noxref_d N_noxref_11_M104_noxref_d N_noxref_11_M106_noxref_d \
 )  PM_TMRDFFRNQNX1\%noxref_11
x_PM_TMRDFFRNQNX1\%D ( N_D_c_4434_n N_D_c_4441_n N_D_c_4442_n N_D_c_4538_n D D \
 N_D_c_4448_n N_D_c_4449_n N_D_c_4450_n N_D_M4_noxref_g N_D_M20_noxref_g \
 N_D_M36_noxref_g N_D_M62_noxref_g N_D_M63_noxref_g N_D_M94_noxref_g \
 N_D_M95_noxref_g N_D_M126_noxref_g N_D_M127_noxref_g N_D_c_4502_n \
 N_D_c_4505_n N_D_c_4749_p N_D_c_4756_p N_D_c_4507_n N_D_c_4508_n N_D_c_4509_n \
 N_D_c_4510_n N_D_c_4482_n N_D_c_4567_n N_D_c_4570_n N_D_c_4770_p N_D_c_4777_p \
 N_D_c_4572_n N_D_c_4573_n N_D_c_4574_n N_D_c_4575_n N_D_c_4546_n N_D_c_4615_p \
 N_D_c_4617_p N_D_c_4790_p N_D_c_4797_p N_D_c_4621_p N_D_c_4623_p N_D_c_4624_p \
 N_D_c_4610_p N_D_c_4598_p N_D_c_4483_n N_D_c_4547_n N_D_c_4599_p )  \
 PM_TMRDFFRNQNX1\%D
x_PM_TMRDFFRNQNX1\%CLK ( N_CLK_c_4808_n N_CLK_c_4825_n N_CLK_c_4826_n \
 N_CLK_c_4843_n N_CLK_c_4844_n N_CLK_c_4861_n N_CLK_c_4862_n N_CLK_c_4879_n \
 N_CLK_c_4880_n N_CLK_c_4897_n CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK \
 CLK CLK CLK CLK N_CLK_c_4802_n N_CLK_c_4803_n N_CLK_c_4804_n N_CLK_c_4805_n \
 N_CLK_c_4806_n N_CLK_c_4807_n N_CLK_M1_noxref_g N_CLK_M9_noxref_g \
 N_CLK_M17_noxref_g N_CLK_M25_noxref_g N_CLK_M33_noxref_g N_CLK_M41_noxref_g \
 N_CLK_M56_noxref_g N_CLK_M57_noxref_g N_CLK_M72_noxref_g N_CLK_M73_noxref_g \
 N_CLK_M88_noxref_g N_CLK_M89_noxref_g N_CLK_M104_noxref_g N_CLK_M105_noxref_g \
 N_CLK_M120_noxref_g N_CLK_M121_noxref_g N_CLK_M136_noxref_g \
 N_CLK_M137_noxref_g N_CLK_c_5060_n N_CLK_c_5063_n N_CLK_c_5475_p \
 N_CLK_c_5482_p N_CLK_c_4952_n N_CLK_c_4953_n N_CLK_c_4954_n N_CLK_c_4955_n \
 N_CLK_c_4958_n N_CLK_c_4976_n N_CLK_c_4979_n N_CLK_c_5495_p N_CLK_c_5502_p \
 N_CLK_c_4981_n N_CLK_c_4982_n N_CLK_c_4983_n N_CLK_c_4984_n N_CLK_c_5070_n \
 N_CLK_c_5205_n N_CLK_c_5208_n N_CLK_c_5515_p N_CLK_c_5522_p N_CLK_c_5094_n \
 N_CLK_c_5095_n N_CLK_c_5096_n N_CLK_c_5097_n N_CLK_c_5100_n N_CLK_c_5118_n \
 N_CLK_c_5121_n N_CLK_c_5535_p N_CLK_c_5542_p N_CLK_c_5123_n N_CLK_c_5124_n \
 N_CLK_c_5125_n N_CLK_c_5126_n N_CLK_c_5215_n N_CLK_c_5363_p N_CLK_c_5365_p \
 N_CLK_c_5555_p N_CLK_c_5562_p N_CLK_c_5369_p N_CLK_c_5371_p N_CLK_c_5372_p \
 N_CLK_c_5265_p N_CLK_c_5250_p N_CLK_c_5426_p N_CLK_c_5428_p N_CLK_c_5575_p \
 N_CLK_c_5582_p N_CLK_c_5306_p N_CLK_c_5307_p N_CLK_c_5308_p N_CLK_c_5267_p \
 N_CLK_c_5332_p N_CLK_c_4959_n N_CLK_c_4986_n N_CLK_c_5101_n N_CLK_c_5128_n \
 N_CLK_c_5242_p N_CLK_c_5288_p )  PM_TMRDFFRNQNX1\%CLK
x_PM_TMRDFFRNQNX1\%noxref_14 ( N_noxref_14_c_5684_n N_noxref_14_c_5685_n \
 N_noxref_14_c_5659_n N_noxref_14_c_5660_n N_noxref_14_c_5611_n \
 N_noxref_14_c_5615_n N_noxref_14_c_5617_n N_noxref_14_c_5621_n \
 N_noxref_14_c_5587_n N_noxref_14_c_5704_p N_noxref_14_c_5625_n \
 N_noxref_14_c_5588_n N_noxref_14_c_5589_n N_noxref_14_c_5699_n \
 N_noxref_14_c_5779_p N_noxref_14_M35_noxref_g N_noxref_14_M43_noxref_g \
 N_noxref_14_M124_noxref_g N_noxref_14_M125_noxref_g N_noxref_14_M140_noxref_g \
 N_noxref_14_M141_noxref_g N_noxref_14_c_5590_n N_noxref_14_c_5592_n \
 N_noxref_14_c_5593_n N_noxref_14_c_5594_n N_noxref_14_c_5595_n \
 N_noxref_14_c_5596_n N_noxref_14_c_5597_n N_noxref_14_c_5599_n \
 N_noxref_14_c_5680_n N_noxref_14_c_5640_n N_noxref_14_c_5600_n \
 N_noxref_14_c_5602_n N_noxref_14_c_5603_n N_noxref_14_c_5604_n \
 N_noxref_14_c_5605_n N_noxref_14_c_5606_n N_noxref_14_c_5607_n \
 N_noxref_14_c_5609_n N_noxref_14_c_5717_p N_noxref_14_c_5642_n \
 N_noxref_14_M34_noxref_d N_noxref_14_M118_noxref_d N_noxref_14_M120_noxref_d \
 N_noxref_14_M122_noxref_d )  PM_TMRDFFRNQNX1\%noxref_14
x_PM_TMRDFFRNQNX1\%RN ( N_RN_c_5846_n N_RN_c_5854_n N_RN_c_5856_n \
 N_RN_c_5860_n N_RN_c_5861_n N_RN_c_5872_n N_RN_c_5873_n N_RN_c_5881_n \
 N_RN_c_5882_n N_RN_c_5886_n N_RN_c_5887_n N_RN_c_5898_n N_RN_c_5899_n \
 N_RN_c_5907_n N_RN_c_5908_n N_RN_c_5912_n RN RN RN RN RN RN RN RN RN RN \
 N_RN_c_5913_n N_RN_c_5914_n N_RN_c_5915_n N_RN_c_5916_n N_RN_c_5917_n \
 N_RN_c_5918_n N_RN_c_5919_n N_RN_c_5920_n N_RN_c_5921_n N_RN_M5_noxref_g \
 N_RN_M10_noxref_g N_RN_M12_noxref_g N_RN_M21_noxref_g N_RN_M26_noxref_g \
 N_RN_M28_noxref_g N_RN_M37_noxref_g N_RN_M42_noxref_g N_RN_M44_noxref_g \
 N_RN_M64_noxref_g N_RN_M65_noxref_g N_RN_M74_noxref_g N_RN_M75_noxref_g \
 N_RN_M78_noxref_g N_RN_M79_noxref_g N_RN_M96_noxref_g N_RN_M97_noxref_g \
 N_RN_M106_noxref_g N_RN_M107_noxref_g N_RN_M110_noxref_g N_RN_M111_noxref_g \
 N_RN_M128_noxref_g N_RN_M129_noxref_g N_RN_M138_noxref_g N_RN_M139_noxref_g \
 N_RN_M142_noxref_g N_RN_M143_noxref_g N_RN_c_5988_n N_RN_c_5989_n \
 N_RN_c_5990_n N_RN_c_5991_n N_RN_c_5992_n N_RN_c_5994_n N_RN_c_5995_n \
 N_RN_c_6075_n N_RN_c_6076_n N_RN_c_6077_n N_RN_c_6078_n N_RN_c_6079_n \
 N_RN_c_6081_n N_RN_c_6082_n N_RN_c_6029_n N_RN_c_6032_n N_RN_c_6631_p \
 N_RN_c_6639_p N_RN_c_6034_n N_RN_c_6035_n N_RN_c_6036_n N_RN_c_6037_n \
 N_RN_c_6084_n N_RN_c_6109_n N_RN_c_6110_n N_RN_c_6111_n N_RN_c_6112_n \
 N_RN_c_6113_n N_RN_c_6115_n N_RN_c_6116_n N_RN_c_6196_n N_RN_c_6197_n \
 N_RN_c_6198_n N_RN_c_6199_n N_RN_c_6200_n N_RN_c_6202_n N_RN_c_6203_n \
 N_RN_c_6149_n N_RN_c_6152_n N_RN_c_6712_p N_RN_c_6720_p N_RN_c_6154_n \
 N_RN_c_6155_n N_RN_c_6156_n N_RN_c_6157_n N_RN_c_6172_n N_RN_c_6268_n \
 N_RN_c_6269_n N_RN_c_6270_n N_RN_c_6513_p N_RN_c_6474_p N_RN_c_6515_p \
 N_RN_c_6475_p N_RN_c_6341_n N_RN_c_6342_n N_RN_c_6343_n N_RN_c_6436_p \
 N_RN_c_6412_p N_RN_c_6438_p N_RN_c_6413_p N_RN_c_6387_n N_RN_c_6390_n \
 N_RN_c_6789_p N_RN_c_6796_p N_RN_c_6392_n N_RN_c_6393_n N_RN_c_6394_n \
 N_RN_c_6395_n N_RN_c_6404_p N_RN_c_5997_n N_RN_c_5998_n N_RN_c_6000_n \
 N_RN_c_6085_n N_RN_c_6086_n N_RN_c_6088_n N_RN_c_6039_n N_RN_c_6118_n \
 N_RN_c_6119_n N_RN_c_6121_n N_RN_c_6205_n N_RN_c_6206_n N_RN_c_6208_n \
 N_RN_c_6159_n N_RN_c_6283_n N_RN_c_6285_n N_RN_c_6286_n N_RN_c_6363_n \
 N_RN_c_6365_n N_RN_c_6366_n N_RN_c_6397_n )  PM_TMRDFFRNQNX1\%RN
x_PM_TMRDFFRNQNX1\%noxref_16 ( N_noxref_16_c_6831_n N_noxref_16_c_6833_n \
 N_noxref_16_c_6834_n N_noxref_16_c_6962_n N_noxref_16_c_6836_n \
 N_noxref_16_c_6842_n N_noxref_16_c_6845_n N_noxref_16_c_6851_n \
 N_noxref_16_c_6854_n N_noxref_16_c_6855_n N_noxref_16_c_6801_n \
 N_noxref_16_c_6968_n N_noxref_16_c_6802_n N_noxref_16_c_6863_n \
 N_noxref_16_c_6867_n N_noxref_16_c_6869_n N_noxref_16_c_6873_n \
 N_noxref_16_c_6804_n N_noxref_16_c_7039_n N_noxref_16_c_6877_n \
 N_noxref_16_c_6878_n N_noxref_16_c_6882_n N_noxref_16_c_6884_n \
 N_noxref_16_c_6888_n N_noxref_16_c_6805_n N_noxref_16_c_7240_p \
 N_noxref_16_c_6892_n N_noxref_16_c_6806_n N_noxref_16_c_7181_p \
 N_noxref_16_c_6807_n N_noxref_16_c_6977_n N_noxref_16_c_7052_n \
 N_noxref_16_c_7054_n N_noxref_16_c_7179_p N_noxref_16_M32_noxref_g \
 N_noxref_16_M39_noxref_g N_noxref_16_M46_noxref_g N_noxref_16_M47_noxref_g \
 N_noxref_16_M118_noxref_g N_noxref_16_M119_noxref_g N_noxref_16_M132_noxref_g \
 N_noxref_16_M133_noxref_g N_noxref_16_M146_noxref_g N_noxref_16_M147_noxref_g \
 N_noxref_16_M148_noxref_g N_noxref_16_M149_noxref_g N_noxref_16_c_6809_n \
 N_noxref_16_c_6811_n N_noxref_16_c_6812_n N_noxref_16_c_6813_n \
 N_noxref_16_c_6814_n N_noxref_16_c_6815_n N_noxref_16_c_6816_n \
 N_noxref_16_c_6818_n N_noxref_16_c_6992_n N_noxref_16_c_6916_n \
 N_noxref_16_c_7136_p N_noxref_16_c_7138_p N_noxref_16_c_7139_p \
 N_noxref_16_c_6997_n N_noxref_16_c_7154_p N_noxref_16_c_7056_n \
 N_noxref_16_c_7144_p N_noxref_16_c_7116_p N_noxref_16_c_6819_n \
 N_noxref_16_c_6821_n N_noxref_16_c_6822_n N_noxref_16_c_6823_n \
 N_noxref_16_c_6824_n N_noxref_16_c_6825_n N_noxref_16_c_6826_n \
 N_noxref_16_c_6828_n N_noxref_16_c_7223_p N_noxref_16_c_7224_p \
 N_noxref_16_c_7225_p N_noxref_16_c_7169_p N_noxref_16_c_7226_p \
 N_noxref_16_c_7191_p N_noxref_16_c_7228_p N_noxref_16_c_7192_p \
 N_noxref_16_c_7057_n N_noxref_16_c_7124_p N_noxref_16_c_6998_n \
 N_noxref_16_c_6918_n N_noxref_16_c_7199_p N_noxref_16_c_7200_p \
 N_noxref_16_c_7170_p N_noxref_16_M42_noxref_d N_noxref_16_M45_noxref_d \
 N_noxref_16_M134_noxref_d N_noxref_16_M136_noxref_d N_noxref_16_M138_noxref_d \
 N_noxref_16_M140_noxref_d N_noxref_16_M142_noxref_d N_noxref_16_M144_noxref_d \
 )  PM_TMRDFFRNQNX1\%noxref_16
x_PM_TMRDFFRNQNX1\%noxref_17 ( N_noxref_17_c_7491_n N_noxref_17_c_7495_n \
 N_noxref_17_c_7362_n N_noxref_17_c_7529_n N_noxref_17_c_7559_n \
 N_noxref_17_c_7561_n N_noxref_17_c_7648_n N_noxref_17_c_7649_n \
 N_noxref_17_c_7650_n N_noxref_17_c_7651_n N_noxref_17_c_7652_n \
 N_noxref_17_c_7653_n N_noxref_17_c_7583_n N_noxref_17_c_7584_n \
 N_noxref_17_c_7363_n N_noxref_17_c_7368_n N_noxref_17_c_7301_n \
 N_noxref_17_c_7373_n N_noxref_17_c_7377_n N_noxref_17_c_7379_n \
 N_noxref_17_c_7302_n N_noxref_17_c_7713_n N_noxref_17_c_7303_n \
 N_noxref_17_c_7304_n N_noxref_17_c_7385_n N_noxref_17_c_7389_n \
 N_noxref_17_c_7391_n N_noxref_17_c_7395_n N_noxref_17_c_7305_n \
 N_noxref_17_c_7721_n N_noxref_17_c_7399_n N_noxref_17_c_7306_n \
 N_noxref_17_c_7403_n N_noxref_17_c_7407_n N_noxref_17_c_7409_n \
 N_noxref_17_c_7307_n N_noxref_17_c_7730_n N_noxref_17_c_7308_n \
 N_noxref_17_c_7309_n N_noxref_17_c_7310_n N_noxref_17_c_7313_n \
 N_noxref_17_c_7544_n N_noxref_17_c_7570_n N_noxref_17_c_7734_n \
 N_noxref_17_c_7824_n N_noxref_17_M29_noxref_g N_noxref_17_M34_noxref_g \
 N_noxref_17_M38_noxref_g N_noxref_17_M40_noxref_g N_noxref_17_M48_noxref_g \
 N_noxref_17_M50_noxref_g N_noxref_17_M112_noxref_g N_noxref_17_M113_noxref_g \
 N_noxref_17_M122_noxref_g N_noxref_17_M123_noxref_g N_noxref_17_M130_noxref_g \
 N_noxref_17_M131_noxref_g N_noxref_17_M134_noxref_g N_noxref_17_M135_noxref_g \
 N_noxref_17_M150_noxref_g N_noxref_17_M151_noxref_g N_noxref_17_M154_noxref_g \
 N_noxref_17_M155_noxref_g N_noxref_17_c_7510_n N_noxref_17_c_7511_n \
 N_noxref_17_c_7512_n N_noxref_17_c_7513_n N_noxref_17_c_7514_n \
 N_noxref_17_c_7516_n N_noxref_17_c_7517_n N_noxref_17_c_7614_n \
 N_noxref_17_c_7615_n N_noxref_17_c_7616_n N_noxref_17_c_7677_n \
 N_noxref_17_c_7678_n N_noxref_17_c_7680_n N_noxref_17_c_7681_n \
 N_noxref_17_c_7315_n N_noxref_17_c_7317_n N_noxref_17_c_7318_n \
 N_noxref_17_c_7319_n N_noxref_17_c_7320_n N_noxref_17_c_7321_n \
 N_noxref_17_c_7322_n N_noxref_17_c_7324_n N_noxref_17_c_7325_n \
 N_noxref_17_c_7327_n N_noxref_17_c_7328_n N_noxref_17_c_7329_n \
 N_noxref_17_c_7330_n N_noxref_17_c_7331_n N_noxref_17_c_7332_n \
 N_noxref_17_c_7334_n N_noxref_17_c_7627_n N_noxref_17_c_7447_n \
 N_noxref_17_c_7335_n N_noxref_17_c_7337_n N_noxref_17_c_7338_n \
 N_noxref_17_c_7339_n N_noxref_17_c_7340_n N_noxref_17_c_7341_n \
 N_noxref_17_c_7875_p N_noxref_17_c_7449_n N_noxref_17_c_7342_n \
 N_noxref_17_c_7344_n N_noxref_17_c_7345_n N_noxref_17_c_7347_n \
 N_noxref_17_c_7958_p N_noxref_17_c_7348_n N_noxref_17_c_7349_n \
 N_noxref_17_c_7350_n N_noxref_17_c_7351_n N_noxref_17_c_7353_n \
 N_noxref_17_c_7519_n N_noxref_17_c_7520_n N_noxref_17_c_7522_n \
 N_noxref_17_c_7633_n N_noxref_17_c_7635_n N_noxref_17_c_7636_n \
 N_noxref_17_c_7451_n N_noxref_17_c_7354_n N_noxref_17_c_7452_n \
 N_noxref_17_M31_noxref_d N_noxref_17_M37_noxref_d N_noxref_17_M39_noxref_d \
 N_noxref_17_M114_noxref_d N_noxref_17_M116_noxref_d N_noxref_17_M124_noxref_d \
 N_noxref_17_M126_noxref_d N_noxref_17_M128_noxref_d N_noxref_17_M130_noxref_d \
 N_noxref_17_M132_noxref_d )  PM_TMRDFFRNQNX1\%noxref_17
x_PM_TMRDFFRNQNX1\%noxref_18 ( N_noxref_18_c_8076_n N_noxref_18_c_8127_n \
 N_noxref_18_c_8077_n N_noxref_18_c_8079_n N_noxref_18_c_8064_n \
 N_noxref_18_c_8085_n N_noxref_18_c_8065_n N_noxref_18_c_8087_n \
 N_noxref_18_c_8091_n N_noxref_18_c_8093_n N_noxref_18_c_8066_n \
 N_noxref_18_c_8286_p N_noxref_18_c_8067_n N_noxref_18_c_8099_n \
 N_noxref_18_c_8068_n N_noxref_18_c_8070_n N_noxref_18_c_8188_n \
 N_noxref_18_c_8309_p N_noxref_18_M45_noxref_g N_noxref_18_M49_noxref_g \
 N_noxref_18_M53_noxref_g N_noxref_18_M144_noxref_g N_noxref_18_M145_noxref_g \
 N_noxref_18_M152_noxref_g N_noxref_18_M153_noxref_g N_noxref_18_M160_noxref_g \
 N_noxref_18_M161_noxref_g N_noxref_18_c_8137_n N_noxref_18_c_8138_n \
 N_noxref_18_c_8139_n N_noxref_18_c_8196_n N_noxref_18_c_8197_n \
 N_noxref_18_c_8199_n N_noxref_18_c_8200_n N_noxref_18_c_8250_n \
 N_noxref_18_c_8253_n N_noxref_18_c_8255_n N_noxref_18_c_8114_n \
 N_noxref_18_c_8340_p N_noxref_18_c_8341_p N_noxref_18_c_8259_n \
 N_noxref_18_c_8260_n N_noxref_18_c_8305_p N_noxref_18_c_8316_p \
 N_noxref_18_c_8307_p N_noxref_18_c_8357_p N_noxref_18_c_8348_p \
 N_noxref_18_c_8318_p N_noxref_18_c_8315_p N_noxref_18_c_8319_p \
 N_noxref_18_c_8140_n N_noxref_18_c_8143_n N_noxref_18_c_8144_n \
 N_noxref_18_c_8072_n N_noxref_18_c_8412_p N_noxref_18_c_8115_n \
 N_noxref_18_c_8293_p N_noxref_18_c_8359_p N_noxref_18_c_8299_p \
 N_noxref_18_M47_noxref_d N_noxref_18_M146_noxref_d N_noxref_18_M148_noxref_d ) \
 PM_TMRDFFRNQNX1\%noxref_18
x_PM_TMRDFFRNQNX1\%noxref_19 ( N_noxref_19_c_8424_n N_noxref_19_c_8430_n \
 N_noxref_19_c_8435_n N_noxref_19_c_8439_n N_noxref_19_c_8441_n \
 N_noxref_19_c_8444_n N_noxref_19_c_8470_n N_noxref_19_c_8446_n \
 N_noxref_19_c_8489_p N_noxref_19_M150_noxref_d N_noxref_19_M152_noxref_d \
 N_noxref_19_M154_noxref_s N_noxref_19_M155_noxref_d N_noxref_19_M157_noxref_d \
 )  PM_TMRDFFRNQNX1\%noxref_19
x_PM_TMRDFFRNQNX1\%noxref_20 ( N_noxref_20_c_8515_n N_noxref_20_c_8606_n \
 N_noxref_20_c_8516_n N_noxref_20_c_8608_n N_noxref_20_c_8536_n \
 N_noxref_20_c_8537_n N_noxref_20_c_8538_n N_noxref_20_c_8560_n \
 N_noxref_20_c_8564_n N_noxref_20_c_8566_n N_noxref_20_c_8539_n \
 N_noxref_20_c_8761_n N_noxref_20_c_8540_n N_noxref_20_c_8541_n \
 N_noxref_20_c_8543_n N_noxref_20_c_8633_n N_noxref_20_M13_noxref_g \
 N_noxref_20_M51_noxref_g N_noxref_20_M52_noxref_g N_noxref_20_M80_noxref_g \
 N_noxref_20_M81_noxref_g N_noxref_20_M156_noxref_g N_noxref_20_M157_noxref_g \
 N_noxref_20_M158_noxref_g N_noxref_20_M159_noxref_g N_noxref_20_c_8638_n \
 N_noxref_20_c_8639_n N_noxref_20_c_8640_n N_noxref_20_c_8641_n \
 N_noxref_20_c_8642_n N_noxref_20_c_8644_n N_noxref_20_c_8645_n \
 N_noxref_20_c_8825_n N_noxref_20_c_8828_n N_noxref_20_c_8901_p \
 N_noxref_20_c_8830_n N_noxref_20_c_8929_p N_noxref_20_c_8930_p \
 N_noxref_20_c_8584_n N_noxref_20_c_8834_n N_noxref_20_c_8835_n \
 N_noxref_20_c_8836_n N_noxref_20_c_8544_n N_noxref_20_c_8545_n \
 N_noxref_20_c_8547_n N_noxref_20_c_8866_n N_noxref_20_c_8548_n \
 N_noxref_20_c_8549_n N_noxref_20_c_8550_n N_noxref_20_c_8868_n \
 N_noxref_20_c_8585_n N_noxref_20_c_8551_n N_noxref_20_c_8553_n \
 N_noxref_20_c_8647_n N_noxref_20_c_8648_n N_noxref_20_c_8650_n \
 N_noxref_20_c_8554_n N_noxref_20_M15_noxref_d N_noxref_20_M82_noxref_d \
 N_noxref_20_M84_noxref_d )  PM_TMRDFFRNQNX1\%noxref_20
x_PM_TMRDFFRNQNX1\%noxref_21 ( N_noxref_21_c_9008_n N_noxref_21_c_9012_n \
 N_noxref_21_c_9023_n N_noxref_21_c_9014_n N_noxref_21_c_9015_n \
 N_noxref_21_c_9016_n N_noxref_21_c_9035_n N_noxref_21_c_9018_n \
 N_noxref_21_c_9036_n N_noxref_21_M154_noxref_d N_noxref_21_M156_noxref_d \
 N_noxref_21_M158_noxref_s N_noxref_21_M159_noxref_d N_noxref_21_M161_noxref_d \
 )  PM_TMRDFFRNQNX1\%noxref_21
x_PM_TMRDFFRNQNX1\%QN ( N_QN_c_9097_n N_QN_c_9104_n N_QN_c_9105_n \
 N_QN_c_9111_n QN QN QN QN QN QN QN QN N_QN_c_9164_n N_QN_c_9126_n \
 N_QN_c_9127_n N_QN_c_9113_n N_QN_c_9171_n N_QN_c_9172_n N_QN_M49_noxref_d \
 N_QN_M51_noxref_d N_QN_M53_noxref_d N_QN_M158_noxref_d N_QN_M160_noxref_d )  \
 PM_TMRDFFRNQNX1\%QN
x_PM_TMRDFFRNQNX1\%noxref_23 ( N_noxref_23_c_9282_n N_noxref_23_c_9266_n \
 N_noxref_23_c_9270_n N_noxref_23_c_9273_n N_noxref_23_c_9290_n \
 N_noxref_23_M0_noxref_s )  PM_TMRDFFRNQNX1\%noxref_23
x_PM_TMRDFFRNQNX1\%noxref_24 ( N_noxref_24_c_9312_n N_noxref_24_c_9314_n \
 N_noxref_24_c_9317_n N_noxref_24_c_9319_n N_noxref_24_c_9330_n \
 N_noxref_24_M1_noxref_d N_noxref_24_M2_noxref_s )  PM_TMRDFFRNQNX1\%noxref_24
x_PM_TMRDFFRNQNX1\%noxref_25 ( N_noxref_25_c_9379_n N_noxref_25_c_9364_n \
 N_noxref_25_c_9368_n N_noxref_25_c_9371_n N_noxref_25_c_9381_n \
 N_noxref_25_M3_noxref_s )  PM_TMRDFFRNQNX1\%noxref_25
x_PM_TMRDFFRNQNX1\%noxref_26 ( N_noxref_26_c_9416_n N_noxref_26_c_9418_n \
 N_noxref_26_c_9421_n N_noxref_26_c_9423_n N_noxref_26_c_9431_n \
 N_noxref_26_M4_noxref_d N_noxref_26_M5_noxref_s )  PM_TMRDFFRNQNX1\%noxref_26
x_PM_TMRDFFRNQNX1\%noxref_27 ( N_noxref_27_c_9487_n N_noxref_27_c_9469_n \
 N_noxref_27_c_9473_n N_noxref_27_c_9476_n N_noxref_27_c_9477_n \
 N_noxref_27_c_9479_n N_noxref_27_M6_noxref_s )  PM_TMRDFFRNQNX1\%noxref_27
x_PM_TMRDFFRNQNX1\%noxref_28 ( N_noxref_28_c_9535_n N_noxref_28_c_9520_n \
 N_noxref_28_c_9524_n N_noxref_28_c_9527_n N_noxref_28_c_9550_n \
 N_noxref_28_M8_noxref_s )  PM_TMRDFFRNQNX1\%noxref_28
x_PM_TMRDFFRNQNX1\%noxref_29 ( N_noxref_29_c_9569_n N_noxref_29_c_9571_n \
 N_noxref_29_c_9574_n N_noxref_29_c_9576_n N_noxref_29_c_9584_n \
 N_noxref_29_M9_noxref_d N_noxref_29_M10_noxref_s )  PM_TMRDFFRNQNX1\%noxref_29
x_PM_TMRDFFRNQNX1\%noxref_30 ( N_noxref_30_c_9637_n N_noxref_30_c_9622_n \
 N_noxref_30_c_9626_n N_noxref_30_c_9629_n N_noxref_30_c_9654_n \
 N_noxref_30_M11_noxref_s )  PM_TMRDFFRNQNX1\%noxref_30
x_PM_TMRDFFRNQNX1\%noxref_31 ( N_noxref_31_c_9674_n N_noxref_31_c_9676_n \
 N_noxref_31_c_9679_n N_noxref_31_c_9681_n N_noxref_31_c_9689_n \
 N_noxref_31_M12_noxref_d N_noxref_31_M13_noxref_s )  PM_TMRDFFRNQNX1\%noxref_31
x_PM_TMRDFFRNQNX1\%noxref_32 ( N_noxref_32_c_9744_n N_noxref_32_c_9726_n \
 N_noxref_32_c_9730_n N_noxref_32_c_9733_n N_noxref_32_c_9734_n \
 N_noxref_32_c_9736_n N_noxref_32_M14_noxref_s )  PM_TMRDFFRNQNX1\%noxref_32
x_PM_TMRDFFRNQNX1\%noxref_33 ( N_noxref_33_c_9793_n N_noxref_33_c_9777_n \
 N_noxref_33_c_9781_n N_noxref_33_c_9784_n N_noxref_33_c_9805_n \
 N_noxref_33_M16_noxref_s )  PM_TMRDFFRNQNX1\%noxref_33
x_PM_TMRDFFRNQNX1\%noxref_34 ( N_noxref_34_c_9826_n N_noxref_34_c_9828_n \
 N_noxref_34_c_9831_n N_noxref_34_c_9833_n N_noxref_34_c_9843_n \
 N_noxref_34_M17_noxref_d N_noxref_34_M18_noxref_s )  PM_TMRDFFRNQNX1\%noxref_34
x_PM_TMRDFFRNQNX1\%noxref_35 ( N_noxref_35_c_9894_n N_noxref_35_c_9878_n \
 N_noxref_35_c_9882_n N_noxref_35_c_9885_n N_noxref_35_c_9908_n \
 N_noxref_35_M19_noxref_s )  PM_TMRDFFRNQNX1\%noxref_35
x_PM_TMRDFFRNQNX1\%noxref_36 ( N_noxref_36_c_9927_n N_noxref_36_c_9929_n \
 N_noxref_36_c_9932_n N_noxref_36_c_9934_n N_noxref_36_c_9942_n \
 N_noxref_36_M20_noxref_d N_noxref_36_M21_noxref_s )  PM_TMRDFFRNQNX1\%noxref_36
x_PM_TMRDFFRNQNX1\%noxref_37 ( N_noxref_37_c_9998_n N_noxref_37_c_9980_n \
 N_noxref_37_c_9984_n N_noxref_37_c_9987_n N_noxref_37_c_9988_n \
 N_noxref_37_c_9990_n N_noxref_37_M22_noxref_s )  PM_TMRDFFRNQNX1\%noxref_37
x_PM_TMRDFFRNQNX1\%noxref_38 ( N_noxref_38_c_10046_n N_noxref_38_c_10031_n \
 N_noxref_38_c_10035_n N_noxref_38_c_10038_n N_noxref_38_c_10061_n \
 N_noxref_38_M24_noxref_s )  PM_TMRDFFRNQNX1\%noxref_38
x_PM_TMRDFFRNQNX1\%noxref_39 ( N_noxref_39_c_10080_n N_noxref_39_c_10082_n \
 N_noxref_39_c_10085_n N_noxref_39_c_10087_n N_noxref_39_c_10095_n \
 N_noxref_39_M25_noxref_d N_noxref_39_M26_noxref_s )  PM_TMRDFFRNQNX1\%noxref_39
x_PM_TMRDFFRNQNX1\%noxref_40 ( N_noxref_40_c_10148_n N_noxref_40_c_10133_n \
 N_noxref_40_c_10137_n N_noxref_40_c_10140_n N_noxref_40_c_10165_n \
 N_noxref_40_M27_noxref_s )  PM_TMRDFFRNQNX1\%noxref_40
x_PM_TMRDFFRNQNX1\%noxref_41 ( N_noxref_41_c_10185_n N_noxref_41_c_10187_n \
 N_noxref_41_c_10190_n N_noxref_41_c_10192_n N_noxref_41_c_10200_n \
 N_noxref_41_M28_noxref_d N_noxref_41_M29_noxref_s )  PM_TMRDFFRNQNX1\%noxref_41
x_PM_TMRDFFRNQNX1\%noxref_42 ( N_noxref_42_c_10255_n N_noxref_42_c_10237_n \
 N_noxref_42_c_10241_n N_noxref_42_c_10244_n N_noxref_42_c_10245_n \
 N_noxref_42_c_10247_n N_noxref_42_M30_noxref_s )  PM_TMRDFFRNQNX1\%noxref_42
x_PM_TMRDFFRNQNX1\%noxref_43 ( N_noxref_43_c_10312_n N_noxref_43_c_10288_n \
 N_noxref_43_c_10292_n N_noxref_43_c_10295_n N_noxref_43_c_10305_n \
 N_noxref_43_M32_noxref_s )  PM_TMRDFFRNQNX1\%noxref_43
x_PM_TMRDFFRNQNX1\%noxref_44 ( N_noxref_44_c_10337_n N_noxref_44_c_10339_n \
 N_noxref_44_c_10342_n N_noxref_44_c_10344_n N_noxref_44_c_10364_n \
 N_noxref_44_M33_noxref_d N_noxref_44_M34_noxref_s )  PM_TMRDFFRNQNX1\%noxref_44
x_PM_TMRDFFRNQNX1\%noxref_45 ( N_noxref_45_c_10412_n N_noxref_45_c_10389_n \
 N_noxref_45_c_10393_n N_noxref_45_c_10396_n N_noxref_45_c_10406_n \
 N_noxref_45_M35_noxref_s )  PM_TMRDFFRNQNX1\%noxref_45
x_PM_TMRDFFRNQNX1\%noxref_46 ( N_noxref_46_c_10438_n N_noxref_46_c_10440_n \
 N_noxref_46_c_10443_n N_noxref_46_c_10445_n N_noxref_46_c_10470_n \
 N_noxref_46_M36_noxref_d N_noxref_46_M37_noxref_s )  PM_TMRDFFRNQNX1\%noxref_46
x_PM_TMRDFFRNQNX1\%noxref_47 ( N_noxref_47_c_10509_n N_noxref_47_c_10491_n \
 N_noxref_47_c_10495_n N_noxref_47_c_10498_n N_noxref_47_c_10499_n \
 N_noxref_47_c_10501_n N_noxref_47_M38_noxref_s )  PM_TMRDFFRNQNX1\%noxref_47
x_PM_TMRDFFRNQNX1\%noxref_48 ( N_noxref_48_c_10565_n N_noxref_48_c_10542_n \
 N_noxref_48_c_10546_n N_noxref_48_c_10549_n N_noxref_48_c_10559_n \
 N_noxref_48_M40_noxref_s )  PM_TMRDFFRNQNX1\%noxref_48
x_PM_TMRDFFRNQNX1\%noxref_49 ( N_noxref_49_c_10591_n N_noxref_49_c_10593_n \
 N_noxref_49_c_10596_n N_noxref_49_c_10598_n N_noxref_49_c_10623_n \
 N_noxref_49_M41_noxref_d N_noxref_49_M42_noxref_s )  PM_TMRDFFRNQNX1\%noxref_49
x_PM_TMRDFFRNQNX1\%noxref_50 ( N_noxref_50_c_10659_n N_noxref_50_c_10644_n \
 N_noxref_50_c_10648_n N_noxref_50_c_10651_n N_noxref_50_c_10673_n \
 N_noxref_50_M43_noxref_s )  PM_TMRDFFRNQNX1\%noxref_50
x_PM_TMRDFFRNQNX1\%noxref_51 ( N_noxref_51_c_10695_n N_noxref_51_c_10697_n \
 N_noxref_51_c_10700_n N_noxref_51_c_10702_n N_noxref_51_c_10722_n \
 N_noxref_51_M44_noxref_d N_noxref_51_M45_noxref_s )  PM_TMRDFFRNQNX1\%noxref_51
x_PM_TMRDFFRNQNX1\%noxref_52 ( N_noxref_52_c_10765_n N_noxref_52_c_10747_n \
 N_noxref_52_c_10751_n N_noxref_52_c_10754_n N_noxref_52_c_10755_n \
 N_noxref_52_c_10757_n N_noxref_52_M46_noxref_s )  PM_TMRDFFRNQNX1\%noxref_52
x_PM_TMRDFFRNQNX1\%noxref_53 ( N_noxref_53_c_10816_n N_noxref_53_c_10798_n \
 N_noxref_53_c_10802_n N_noxref_53_c_10805_n N_noxref_53_c_10806_n \
 N_noxref_53_c_10808_n N_noxref_53_M48_noxref_s )  PM_TMRDFFRNQNX1\%noxref_53
x_PM_TMRDFFRNQNX1\%noxref_54 ( N_noxref_54_c_10872_n N_noxref_54_c_10855_n \
 N_noxref_54_c_10858_n N_noxref_54_c_10861_n N_noxref_54_c_10862_n \
 N_noxref_54_c_10864_n N_noxref_54_M50_noxref_s )  PM_TMRDFFRNQNX1\%noxref_54
x_PM_TMRDFFRNQNX1\%noxref_55 ( N_noxref_55_c_10937_n N_noxref_55_c_10910_n \
 N_noxref_55_c_10913_n N_noxref_55_c_10916_n N_noxref_55_c_10917_n \
 N_noxref_55_c_10919_n N_noxref_55_M52_noxref_s )  PM_TMRDFFRNQNX1\%noxref_55
cc_1 ( N_GND_c_1_p N_VDD_c_992_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_993_n ) capacitor c=0.00989031f //x=86.95 //y=0 \
 //x2=86.95 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_994_n ) capacitor c=0.00500587f //x=4.81 //y=0 \
 //x2=4.81 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_995_n ) capacitor c=0.0057235f //x=9.62 //y=0 \
 //x2=9.62 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_996_n ) capacitor c=0.0057235f //x=12.95 //y=0 \
 //x2=12.95 //y2=7.4
cc_6 ( N_GND_c_6_p N_VDD_c_997_n ) capacitor c=0.0057235f //x=17.76 //y=0 \
 //x2=17.76 //y2=7.4
cc_7 ( N_GND_c_7_p N_VDD_c_998_n ) capacitor c=0.00579636f //x=22.57 //y=0 \
 //x2=22.57 //y2=7.4
cc_8 ( N_GND_c_8_p N_VDD_c_999_n ) capacitor c=0.00989031f //x=25.9 //y=0 \
 //x2=25.9 //y2=7.4
cc_9 ( N_GND_c_9_p N_VDD_c_1000_n ) capacitor c=0.0057235f //x=30.71 //y=0 \
 //x2=30.71 //y2=7.4
cc_10 ( N_GND_c_10_p N_VDD_c_1001_n ) capacitor c=0.0057235f //x=35.52 //y=0 \
 //x2=35.52 //y2=7.4
cc_11 ( N_GND_c_11_p N_VDD_c_1002_n ) capacitor c=0.0057235f //x=38.85 //y=0 \
 //x2=38.85 //y2=7.4
cc_12 ( N_GND_c_12_p N_VDD_c_1003_n ) capacitor c=0.0057235f //x=43.66 //y=0 \
 //x2=43.66 //y2=7.4
cc_13 ( N_GND_c_13_p N_VDD_c_1004_n ) capacitor c=0.0057235f //x=48.47 //y=0 \
 //x2=48.47 //y2=7.4
cc_14 ( N_GND_c_14_p N_VDD_c_1005_n ) capacitor c=0.00989031f //x=51.8 //y=0 \
 //x2=51.8 //y2=7.4
cc_15 ( N_GND_c_15_p N_VDD_c_1006_n ) capacitor c=0.0057235f //x=56.61 //y=0 \
 //x2=56.61 //y2=7.4
cc_16 ( N_GND_c_16_p N_VDD_c_1007_n ) capacitor c=0.00474727f //x=61.42 //y=0 \
 //x2=61.42 //y2=7.4
cc_17 ( N_GND_c_17_p N_VDD_c_1008_n ) capacitor c=0.00474727f //x=64.75 //y=0 \
 //x2=64.75 //y2=7.4
cc_18 ( N_GND_c_18_p N_VDD_c_1009_n ) capacitor c=0.00474727f //x=69.56 //y=0 \
 //x2=69.56 //y2=7.4
cc_19 ( N_GND_c_19_p N_VDD_c_1010_n ) capacitor c=0.00474727f //x=74.37 //y=0 \
 //x2=74.37 //y2=7.4
cc_20 ( N_GND_c_20_p N_VDD_c_1011_n ) capacitor c=0.00802221f //x=77.7 //y=0 \
 //x2=77.7 //y2=7.4
cc_21 ( N_GND_c_21_p N_VDD_c_1012_n ) capacitor c=0.00482014f //x=81.03 //y=0 \
 //x2=81.03 //y2=7.4
cc_22 ( N_GND_c_22_p N_VDD_c_1013_n ) capacitor c=0.00553669f //x=84.36 //y=0 \
 //x2=84.36 //y2=7.4
cc_23 ( N_GND_c_23_p N_noxref_3_c_2093_n ) capacitor c=0.0265869f //x=86.95 \
 //y=0 //x2=8.765 //y2=3.33
cc_24 ( N_GND_c_24_p N_noxref_3_c_2093_n ) capacitor c=0.00174514f //x=4.64 \
 //y=0 //x2=8.765 //y2=3.33
cc_25 ( N_GND_c_25_p N_noxref_3_c_2093_n ) capacitor c=0.00152503f //x=5.8 \
 //y=0 //x2=8.765 //y2=3.33
cc_26 ( N_GND_c_3_p N_noxref_3_c_2093_n ) capacitor c=0.00820844f //x=4.81 \
 //y=0 //x2=8.765 //y2=3.33
cc_27 ( N_GND_c_23_p N_noxref_3_c_2097_n ) capacitor c=0.00172266f //x=86.95 \
 //y=0 //x2=3.445 //y2=3.33
cc_28 ( N_GND_c_4_p N_noxref_3_c_2098_n ) capacitor c=0.00505527f //x=9.62 \
 //y=0 //x2=10.615 //y2=3.33
cc_29 ( N_GND_c_3_p N_noxref_3_c_2099_n ) capacitor c=9.53263e-19 //x=4.81 \
 //y=0 //x2=3.33 //y2=2.08
cc_30 ( N_GND_c_4_p N_noxref_3_c_2100_n ) capacitor c=0.0405089f //x=9.62 \
 //y=0 //x2=8.795 //y2=1.665
cc_31 ( N_GND_c_4_p N_noxref_3_c_2101_n ) capacitor c=0.0130533f //x=9.62 \
 //y=0 //x2=10.73 //y2=2.08
cc_32 ( N_GND_c_32_p N_noxref_3_c_2102_n ) capacitor c=0.00135046f //x=10.715 \
 //y=0 //x2=10.535 //y2=0.865
cc_33 ( N_GND_M6_noxref_d N_noxref_3_c_2102_n ) capacitor c=0.00220047f \
 //x=10.61 //y=0.865 //x2=10.535 //y2=0.865
cc_34 ( N_GND_M6_noxref_d N_noxref_3_c_2104_n ) capacitor c=0.00255985f \
 //x=10.61 //y=0.865 //x2=10.535 //y2=1.21
cc_35 ( N_GND_c_4_p N_noxref_3_c_2105_n ) capacitor c=0.00189421f //x=9.62 \
 //y=0 //x2=10.535 //y2=1.52
cc_36 ( N_GND_c_4_p N_noxref_3_c_2106_n ) capacitor c=0.00992619f //x=9.62 \
 //y=0 //x2=10.535 //y2=1.915
cc_37 ( N_GND_M6_noxref_d N_noxref_3_c_2107_n ) capacitor c=0.0131326f \
 //x=10.61 //y=0.865 //x2=10.91 //y2=0.71
cc_38 ( N_GND_M6_noxref_d N_noxref_3_c_2108_n ) capacitor c=0.00193127f \
 //x=10.61 //y=0.865 //x2=10.91 //y2=1.365
cc_39 ( N_GND_c_39_p N_noxref_3_c_2109_n ) capacitor c=0.00130622f //x=12.78 \
 //y=0 //x2=11.065 //y2=0.865
cc_40 ( N_GND_M6_noxref_d N_noxref_3_c_2109_n ) capacitor c=0.00257848f \
 //x=10.61 //y=0.865 //x2=11.065 //y2=0.865
cc_41 ( N_GND_M6_noxref_d N_noxref_3_c_2111_n ) capacitor c=0.00255985f \
 //x=10.61 //y=0.865 //x2=11.065 //y2=1.21
cc_42 ( N_GND_c_4_p N_noxref_3_M5_noxref_d ) capacitor c=0.00591582f //x=9.62 \
 //y=0 //x2=8.205 //y2=0.915
cc_43 ( N_GND_c_5_p N_noxref_4_c_2343_n ) capacitor c=0.00505527f //x=12.95 \
 //y=0 //x2=13.945 //y2=3.33
cc_44 ( N_GND_c_5_p N_noxref_4_c_2344_n ) capacitor c=0.0410119f //x=12.95 \
 //y=0 //x2=12.125 //y2=1.655
cc_45 ( N_GND_c_4_p N_noxref_4_c_2345_n ) capacitor c=9.64732e-19 //x=9.62 \
 //y=0 //x2=12.21 //y2=3.33
cc_46 ( N_GND_c_5_p N_noxref_4_c_2346_n ) capacitor c=0.0130528f //x=12.95 \
 //y=0 //x2=14.06 //y2=2.08
cc_47 ( N_GND_c_47_p N_noxref_4_c_2347_n ) capacitor c=0.00132755f //x=13.94 \
 //y=0 //x2=13.76 //y2=0.875
cc_48 ( N_GND_M8_noxref_d N_noxref_4_c_2347_n ) capacitor c=0.00211996f \
 //x=13.835 //y=0.875 //x2=13.76 //y2=0.875
cc_49 ( N_GND_M8_noxref_d N_noxref_4_c_2349_n ) capacitor c=0.00255985f \
 //x=13.835 //y=0.875 //x2=13.76 //y2=1.22
cc_50 ( N_GND_c_5_p N_noxref_4_c_2350_n ) capacitor c=0.00195164f //x=12.95 \
 //y=0 //x2=13.76 //y2=1.53
cc_51 ( N_GND_c_5_p N_noxref_4_c_2351_n ) capacitor c=0.0110952f //x=12.95 \
 //y=0 //x2=13.76 //y2=1.915
cc_52 ( N_GND_M8_noxref_d N_noxref_4_c_2352_n ) capacitor c=0.0131341f \
 //x=13.835 //y=0.875 //x2=14.135 //y2=0.72
cc_53 ( N_GND_M8_noxref_d N_noxref_4_c_2353_n ) capacitor c=0.00193146f \
 //x=13.835 //y=0.875 //x2=14.135 //y2=1.375
cc_54 ( N_GND_c_54_p N_noxref_4_c_2354_n ) capacitor c=0.00129018f //x=17.59 \
 //y=0 //x2=14.29 //y2=0.875
cc_55 ( N_GND_M8_noxref_d N_noxref_4_c_2354_n ) capacitor c=0.00257848f \
 //x=13.835 //y=0.875 //x2=14.29 //y2=0.875
cc_56 ( N_GND_M8_noxref_d N_noxref_4_c_2356_n ) capacitor c=0.00255985f \
 //x=13.835 //y=0.875 //x2=14.29 //y2=1.22
cc_57 ( N_GND_c_4_p N_noxref_4_M7_noxref_d ) capacitor c=8.58106e-19 //x=9.62 \
 //y=0 //x2=11.58 //y2=0.905
cc_58 ( N_GND_c_5_p N_noxref_4_M7_noxref_d ) capacitor c=0.00616547f //x=12.95 \
 //y=0 //x2=11.58 //y2=0.905
cc_59 ( N_GND_M6_noxref_d N_noxref_4_M7_noxref_d ) capacitor c=0.00143464f \
 //x=10.61 //y=0.865 //x2=11.58 //y2=0.905
cc_60 ( N_GND_c_6_p N_noxref_5_c_2495_n ) capacitor c=0.0034979f //x=17.76 \
 //y=0 //x2=18.755 //y2=3.7
cc_61 ( N_GND_c_3_p N_noxref_5_c_2496_n ) capacitor c=0.0455868f //x=4.81 \
 //y=0 //x2=3.985 //y2=1.665
cc_62 ( N_GND_c_3_p N_noxref_5_c_2497_n ) capacitor c=0.0175021f //x=4.81 \
 //y=0 //x2=5.92 //y2=2.08
cc_63 ( N_GND_c_6_p N_noxref_5_c_2498_n ) capacitor c=0.0129883f //x=17.76 \
 //y=0 //x2=18.87 //y2=2.08
cc_64 ( N_GND_c_25_p N_noxref_5_c_2499_n ) capacitor c=0.00132755f //x=5.8 \
 //y=0 //x2=5.62 //y2=0.875
cc_65 ( N_GND_M3_noxref_d N_noxref_5_c_2499_n ) capacitor c=0.00211996f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=0.875
cc_66 ( N_GND_M3_noxref_d N_noxref_5_c_2501_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=1.22
cc_67 ( N_GND_c_3_p N_noxref_5_c_2502_n ) capacitor c=0.00204716f //x=4.81 \
 //y=0 //x2=5.62 //y2=1.53
cc_68 ( N_GND_c_3_p N_noxref_5_c_2503_n ) capacitor c=0.0118433f //x=4.81 \
 //y=0 //x2=5.62 //y2=1.915
cc_69 ( N_GND_M3_noxref_d N_noxref_5_c_2504_n ) capacitor c=0.0131341f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=0.72
cc_70 ( N_GND_M3_noxref_d N_noxref_5_c_2505_n ) capacitor c=0.00193146f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=1.375
cc_71 ( N_GND_c_71_p N_noxref_5_c_2506_n ) capacitor c=0.00129018f //x=9.45 \
 //y=0 //x2=6.15 //y2=0.875
cc_72 ( N_GND_M3_noxref_d N_noxref_5_c_2506_n ) capacitor c=0.00257848f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=0.875
cc_73 ( N_GND_M3_noxref_d N_noxref_5_c_2508_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=1.22
cc_74 ( N_GND_c_74_p N_noxref_5_c_2509_n ) capacitor c=0.00132755f //x=18.75 \
 //y=0 //x2=18.57 //y2=0.875
cc_75 ( N_GND_M11_noxref_d N_noxref_5_c_2509_n ) capacitor c=0.00211996f \
 //x=18.645 //y=0.875 //x2=18.57 //y2=0.875
cc_76 ( N_GND_M11_noxref_d N_noxref_5_c_2511_n ) capacitor c=0.00255985f \
 //x=18.645 //y=0.875 //x2=18.57 //y2=1.22
cc_77 ( N_GND_c_6_p N_noxref_5_c_2512_n ) capacitor c=0.00204716f //x=17.76 \
 //y=0 //x2=18.57 //y2=1.53
cc_78 ( N_GND_c_6_p N_noxref_5_c_2513_n ) capacitor c=0.0110952f //x=17.76 \
 //y=0 //x2=18.57 //y2=1.915
cc_79 ( N_GND_M11_noxref_d N_noxref_5_c_2514_n ) capacitor c=0.0131341f \
 //x=18.645 //y=0.875 //x2=18.945 //y2=0.72
cc_80 ( N_GND_M11_noxref_d N_noxref_5_c_2515_n ) capacitor c=0.00193146f \
 //x=18.645 //y=0.875 //x2=18.945 //y2=1.375
cc_81 ( N_GND_c_81_p N_noxref_5_c_2516_n ) capacitor c=0.00129018f //x=22.4 \
 //y=0 //x2=19.1 //y2=0.875
cc_82 ( N_GND_M11_noxref_d N_noxref_5_c_2516_n ) capacitor c=0.00257848f \
 //x=18.645 //y=0.875 //x2=19.1 //y2=0.875
cc_83 ( N_GND_M11_noxref_d N_noxref_5_c_2518_n ) capacitor c=0.00255985f \
 //x=18.645 //y=0.875 //x2=19.1 //y2=1.22
cc_84 ( N_GND_c_3_p N_noxref_5_M2_noxref_d ) capacitor c=0.00591582f //x=4.81 \
 //y=0 //x2=3.395 //y2=0.915
cc_85 ( N_GND_c_23_p N_noxref_6_c_2748_n ) capacitor c=0.0122686f //x=86.95 \
 //y=0 //x2=11.355 //y2=4.07
cc_86 ( N_GND_c_23_p N_noxref_6_c_2749_n ) capacitor c=0.0015877f //x=86.95 \
 //y=0 //x2=1.225 //y2=4.07
cc_87 ( N_GND_c_1_p N_noxref_6_c_2750_n ) capacitor c=0.0180363f //x=0.74 \
 //y=0 //x2=1.11 //y2=2.08
cc_88 ( N_GND_c_4_p N_noxref_6_c_2751_n ) capacitor c=5.78225e-19 //x=9.62 \
 //y=0 //x2=11.47 //y2=2.08
cc_89 ( N_GND_c_5_p N_noxref_6_c_2751_n ) capacitor c=5.32623e-19 //x=12.95 \
 //y=0 //x2=11.47 //y2=2.08
cc_90 ( N_GND_c_6_p N_noxref_6_c_2753_n ) capacitor c=0.0404734f //x=17.76 \
 //y=0 //x2=16.935 //y2=1.665
cc_91 ( N_GND_c_7_p N_noxref_6_c_2754_n ) capacitor c=0.0406661f //x=22.57 \
 //y=0 //x2=21.745 //y2=1.665
cc_92 ( N_GND_c_7_p N_noxref_6_c_2755_n ) capacitor c=0.0131041f //x=22.57 \
 //y=0 //x2=23.68 //y2=2.08
cc_93 ( N_GND_c_7_p N_noxref_6_c_2756_n ) capacitor c=5.41726e-19 //x=22.57 \
 //y=0 //x2=24.42 //y2=2.08
cc_94 ( N_GND_c_8_p N_noxref_6_c_2756_n ) capacitor c=5.32623e-19 //x=25.9 \
 //y=0 //x2=24.42 //y2=2.08
cc_95 ( N_GND_c_95_p N_noxref_6_c_2758_n ) capacitor c=0.00132755f //x=0.99 \
 //y=0 //x2=0.81 //y2=0.875
cc_96 ( N_GND_M0_noxref_d N_noxref_6_c_2758_n ) capacitor c=0.00211996f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=0.875
cc_97 ( N_GND_M0_noxref_d N_noxref_6_c_2760_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=1.22
cc_98 ( N_GND_c_1_p N_noxref_6_c_2761_n ) capacitor c=0.00295461f //x=0.74 \
 //y=0 //x2=0.81 //y2=1.53
cc_99 ( N_GND_c_1_p N_noxref_6_c_2762_n ) capacitor c=0.0134214f //x=0.74 \
 //y=0 //x2=0.81 //y2=1.915
cc_100 ( N_GND_M0_noxref_d N_noxref_6_c_2763_n ) capacitor c=0.0131341f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=0.72
cc_101 ( N_GND_M0_noxref_d N_noxref_6_c_2764_n ) capacitor c=0.00193146f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=1.375
cc_102 ( N_GND_c_24_p N_noxref_6_c_2765_n ) capacitor c=0.00129018f //x=4.64 \
 //y=0 //x2=1.34 //y2=0.875
cc_103 ( N_GND_M0_noxref_d N_noxref_6_c_2765_n ) capacitor c=0.00257848f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=0.875
cc_104 ( N_GND_M0_noxref_d N_noxref_6_c_2767_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=1.22
cc_105 ( N_GND_c_105_p N_noxref_6_c_2768_n ) capacitor c=0.00135046f \
 //x=23.665 //y=0 //x2=23.485 //y2=0.865
cc_106 ( N_GND_M14_noxref_d N_noxref_6_c_2768_n ) capacitor c=0.00220047f \
 //x=23.56 //y=0.865 //x2=23.485 //y2=0.865
cc_107 ( N_GND_M14_noxref_d N_noxref_6_c_2770_n ) capacitor c=0.00255985f \
 //x=23.56 //y=0.865 //x2=23.485 //y2=1.21
cc_108 ( N_GND_c_7_p N_noxref_6_c_2771_n ) capacitor c=0.00189421f //x=22.57 \
 //y=0 //x2=23.485 //y2=1.52
cc_109 ( N_GND_c_7_p N_noxref_6_c_2772_n ) capacitor c=0.00992619f //x=22.57 \
 //y=0 //x2=23.485 //y2=1.915
cc_110 ( N_GND_M14_noxref_d N_noxref_6_c_2773_n ) capacitor c=0.0131326f \
 //x=23.56 //y=0.865 //x2=23.86 //y2=0.71
cc_111 ( N_GND_M14_noxref_d N_noxref_6_c_2774_n ) capacitor c=0.00193127f \
 //x=23.56 //y=0.865 //x2=23.86 //y2=1.365
cc_112 ( N_GND_c_112_p N_noxref_6_c_2775_n ) capacitor c=0.00130622f //x=25.73 \
 //y=0 //x2=24.015 //y2=0.865
cc_113 ( N_GND_M14_noxref_d N_noxref_6_c_2775_n ) capacitor c=0.00257848f \
 //x=23.56 //y=0.865 //x2=24.015 //y2=0.865
cc_114 ( N_GND_M14_noxref_d N_noxref_6_c_2777_n ) capacitor c=0.00255985f \
 //x=23.56 //y=0.865 //x2=24.015 //y2=1.21
cc_115 ( N_GND_c_6_p N_noxref_6_M10_noxref_d ) capacitor c=0.00591582f \
 //x=17.76 //y=0 //x2=16.345 //y2=0.915
cc_116 ( N_GND_c_7_p N_noxref_6_M13_noxref_d ) capacitor c=0.00591582f \
 //x=22.57 //y=0 //x2=21.155 //y2=0.915
cc_117 ( N_GND_c_9_p N_noxref_7_c_3233_n ) capacitor c=5.32623e-19 //x=30.71 \
 //y=0 //x2=29.23 //y2=2.08
cc_118 ( N_GND_c_10_p N_noxref_7_c_3234_n ) capacitor c=0.0405089f //x=35.52 \
 //y=0 //x2=34.695 //y2=1.665
cc_119 ( N_GND_c_10_p N_noxref_7_c_3235_n ) capacitor c=0.0130533f //x=35.52 \
 //y=0 //x2=36.63 //y2=2.08
cc_120 ( N_GND_c_120_p N_noxref_7_c_3236_n ) capacitor c=0.00135046f \
 //x=36.615 //y=0 //x2=36.435 //y2=0.865
cc_121 ( N_GND_M22_noxref_d N_noxref_7_c_3236_n ) capacitor c=0.00220047f \
 //x=36.51 //y=0.865 //x2=36.435 //y2=0.865
cc_122 ( N_GND_M22_noxref_d N_noxref_7_c_3238_n ) capacitor c=0.00255985f \
 //x=36.51 //y=0.865 //x2=36.435 //y2=1.21
cc_123 ( N_GND_c_10_p N_noxref_7_c_3239_n ) capacitor c=0.00189421f //x=35.52 \
 //y=0 //x2=36.435 //y2=1.52
cc_124 ( N_GND_c_10_p N_noxref_7_c_3240_n ) capacitor c=0.00992619f //x=35.52 \
 //y=0 //x2=36.435 //y2=1.915
cc_125 ( N_GND_M22_noxref_d N_noxref_7_c_3241_n ) capacitor c=0.0131326f \
 //x=36.51 //y=0.865 //x2=36.81 //y2=0.71
cc_126 ( N_GND_M22_noxref_d N_noxref_7_c_3242_n ) capacitor c=0.00193127f \
 //x=36.51 //y=0.865 //x2=36.81 //y2=1.365
cc_127 ( N_GND_c_127_p N_noxref_7_c_3243_n ) capacitor c=0.00130622f //x=38.68 \
 //y=0 //x2=36.965 //y2=0.865
cc_128 ( N_GND_M22_noxref_d N_noxref_7_c_3243_n ) capacitor c=0.00257848f \
 //x=36.51 //y=0.865 //x2=36.965 //y2=0.865
cc_129 ( N_GND_M22_noxref_d N_noxref_7_c_3245_n ) capacitor c=0.00255985f \
 //x=36.51 //y=0.865 //x2=36.965 //y2=1.21
cc_130 ( N_GND_c_10_p N_noxref_7_M21_noxref_d ) capacitor c=0.00591582f \
 //x=35.52 //y=0 //x2=34.105 //y2=0.915
cc_131 ( N_GND_c_11_p N_noxref_8_c_3480_n ) capacitor c=0.0410119f //x=38.85 \
 //y=0 //x2=38.025 //y2=1.655
cc_132 ( N_GND_c_10_p N_noxref_8_c_3481_n ) capacitor c=9.64732e-19 //x=35.52 \
 //y=0 //x2=38.11 //y2=3.33
cc_133 ( N_GND_c_11_p N_noxref_8_c_3482_n ) capacitor c=0.0130528f //x=38.85 \
 //y=0 //x2=39.96 //y2=2.08
cc_134 ( N_GND_c_134_p N_noxref_8_c_3483_n ) capacitor c=0.00132755f //x=39.84 \
 //y=0 //x2=39.66 //y2=0.875
cc_135 ( N_GND_M24_noxref_d N_noxref_8_c_3483_n ) capacitor c=0.00211996f \
 //x=39.735 //y=0.875 //x2=39.66 //y2=0.875
cc_136 ( N_GND_M24_noxref_d N_noxref_8_c_3485_n ) capacitor c=0.00255985f \
 //x=39.735 //y=0.875 //x2=39.66 //y2=1.22
cc_137 ( N_GND_c_11_p N_noxref_8_c_3486_n ) capacitor c=0.00195164f //x=38.85 \
 //y=0 //x2=39.66 //y2=1.53
cc_138 ( N_GND_c_11_p N_noxref_8_c_3487_n ) capacitor c=0.0110952f //x=38.85 \
 //y=0 //x2=39.66 //y2=1.915
cc_139 ( N_GND_M24_noxref_d N_noxref_8_c_3488_n ) capacitor c=0.0131341f \
 //x=39.735 //y=0.875 //x2=40.035 //y2=0.72
cc_140 ( N_GND_M24_noxref_d N_noxref_8_c_3489_n ) capacitor c=0.00193146f \
 //x=39.735 //y=0.875 //x2=40.035 //y2=1.375
cc_141 ( N_GND_c_141_p N_noxref_8_c_3490_n ) capacitor c=0.00129018f //x=43.49 \
 //y=0 //x2=40.19 //y2=0.875
cc_142 ( N_GND_M24_noxref_d N_noxref_8_c_3490_n ) capacitor c=0.00257848f \
 //x=39.735 //y=0.875 //x2=40.19 //y2=0.875
cc_143 ( N_GND_M24_noxref_d N_noxref_8_c_3492_n ) capacitor c=0.00255985f \
 //x=39.735 //y=0.875 //x2=40.19 //y2=1.22
cc_144 ( N_GND_c_10_p N_noxref_8_M23_noxref_d ) capacitor c=8.58106e-19 \
 //x=35.52 //y=0 //x2=37.48 //y2=0.905
cc_145 ( N_GND_c_11_p N_noxref_8_M23_noxref_d ) capacitor c=0.00616547f \
 //x=38.85 //y=0 //x2=37.48 //y2=0.905
cc_146 ( N_GND_M22_noxref_d N_noxref_8_M23_noxref_d ) capacitor c=0.00143464f \
 //x=36.51 //y=0.865 //x2=37.48 //y2=0.905
cc_147 ( N_GND_c_9_p N_noxref_9_c_3633_n ) capacitor c=0.0406306f //x=30.71 \
 //y=0 //x2=29.885 //y2=1.665
cc_148 ( N_GND_c_9_p N_noxref_9_c_3634_n ) capacitor c=0.0129722f //x=30.71 \
 //y=0 //x2=31.82 //y2=2.08
cc_149 ( N_GND_c_12_p N_noxref_9_c_3635_n ) capacitor c=0.0129883f //x=43.66 \
 //y=0 //x2=44.77 //y2=2.08
cc_150 ( N_GND_c_150_p N_noxref_9_c_3636_n ) capacitor c=0.00132755f //x=31.7 \
 //y=0 //x2=31.52 //y2=0.875
cc_151 ( N_GND_M19_noxref_d N_noxref_9_c_3636_n ) capacitor c=0.00211996f \
 //x=31.595 //y=0.875 //x2=31.52 //y2=0.875
cc_152 ( N_GND_M19_noxref_d N_noxref_9_c_3638_n ) capacitor c=0.00255985f \
 //x=31.595 //y=0.875 //x2=31.52 //y2=1.22
cc_153 ( N_GND_c_9_p N_noxref_9_c_3639_n ) capacitor c=0.00204716f //x=30.71 \
 //y=0 //x2=31.52 //y2=1.53
cc_154 ( N_GND_c_9_p N_noxref_9_c_3640_n ) capacitor c=0.0110952f //x=30.71 \
 //y=0 //x2=31.52 //y2=1.915
cc_155 ( N_GND_M19_noxref_d N_noxref_9_c_3641_n ) capacitor c=0.0131341f \
 //x=31.595 //y=0.875 //x2=31.895 //y2=0.72
cc_156 ( N_GND_M19_noxref_d N_noxref_9_c_3642_n ) capacitor c=0.00193146f \
 //x=31.595 //y=0.875 //x2=31.895 //y2=1.375
cc_157 ( N_GND_c_157_p N_noxref_9_c_3643_n ) capacitor c=0.00129018f //x=35.35 \
 //y=0 //x2=32.05 //y2=0.875
cc_158 ( N_GND_M19_noxref_d N_noxref_9_c_3643_n ) capacitor c=0.00257848f \
 //x=31.595 //y=0.875 //x2=32.05 //y2=0.875
cc_159 ( N_GND_M19_noxref_d N_noxref_9_c_3645_n ) capacitor c=0.00255985f \
 //x=31.595 //y=0.875 //x2=32.05 //y2=1.22
cc_160 ( N_GND_c_160_p N_noxref_9_c_3646_n ) capacitor c=0.00132755f //x=44.65 \
 //y=0 //x2=44.47 //y2=0.875
cc_161 ( N_GND_M27_noxref_d N_noxref_9_c_3646_n ) capacitor c=0.00211996f \
 //x=44.545 //y=0.875 //x2=44.47 //y2=0.875
cc_162 ( N_GND_M27_noxref_d N_noxref_9_c_3648_n ) capacitor c=0.00255985f \
 //x=44.545 //y=0.875 //x2=44.47 //y2=1.22
cc_163 ( N_GND_c_12_p N_noxref_9_c_3649_n ) capacitor c=0.00204716f //x=43.66 \
 //y=0 //x2=44.47 //y2=1.53
cc_164 ( N_GND_c_12_p N_noxref_9_c_3650_n ) capacitor c=0.0110952f //x=43.66 \
 //y=0 //x2=44.47 //y2=1.915
cc_165 ( N_GND_M27_noxref_d N_noxref_9_c_3651_n ) capacitor c=0.0131341f \
 //x=44.545 //y=0.875 //x2=44.845 //y2=0.72
cc_166 ( N_GND_M27_noxref_d N_noxref_9_c_3652_n ) capacitor c=0.00193146f \
 //x=44.545 //y=0.875 //x2=44.845 //y2=1.375
cc_167 ( N_GND_c_167_p N_noxref_9_c_3653_n ) capacitor c=0.00129018f //x=48.3 \
 //y=0 //x2=45 //y2=0.875
cc_168 ( N_GND_M27_noxref_d N_noxref_9_c_3653_n ) capacitor c=0.00257848f \
 //x=44.545 //y=0.875 //x2=45 //y2=0.875
cc_169 ( N_GND_M27_noxref_d N_noxref_9_c_3655_n ) capacitor c=0.00255985f \
 //x=44.545 //y=0.875 //x2=45 //y2=1.22
cc_170 ( N_GND_c_9_p N_noxref_9_M18_noxref_d ) capacitor c=0.00591582f \
 //x=30.71 //y=0 //x2=29.295 //y2=0.915
cc_171 ( N_GND_c_13_p N_noxref_10_c_3895_n ) capacitor c=0.0406661f //x=48.47 \
 //y=0 //x2=47.645 //y2=1.665
cc_172 ( N_GND_c_13_p N_noxref_10_c_3896_n ) capacitor c=0.0131041f //x=48.47 \
 //y=0 //x2=49.58 //y2=2.08
cc_173 ( N_GND_c_173_p N_noxref_10_c_3897_n ) capacitor c=0.00135046f \
 //x=49.565 //y=0 //x2=49.385 //y2=0.865
cc_174 ( N_GND_M30_noxref_d N_noxref_10_c_3897_n ) capacitor c=0.00220047f \
 //x=49.46 //y=0.865 //x2=49.385 //y2=0.865
cc_175 ( N_GND_M30_noxref_d N_noxref_10_c_3899_n ) capacitor c=0.00255985f \
 //x=49.46 //y=0.865 //x2=49.385 //y2=1.21
cc_176 ( N_GND_c_13_p N_noxref_10_c_3900_n ) capacitor c=0.00189421f //x=48.47 \
 //y=0 //x2=49.385 //y2=1.52
cc_177 ( N_GND_c_13_p N_noxref_10_c_3901_n ) capacitor c=0.00992619f //x=48.47 \
 //y=0 //x2=49.385 //y2=1.915
cc_178 ( N_GND_M30_noxref_d N_noxref_10_c_3902_n ) capacitor c=0.0131326f \
 //x=49.46 //y=0.865 //x2=49.76 //y2=0.71
cc_179 ( N_GND_M30_noxref_d N_noxref_10_c_3903_n ) capacitor c=0.00193127f \
 //x=49.46 //y=0.865 //x2=49.76 //y2=1.365
cc_180 ( N_GND_c_180_p N_noxref_10_c_3904_n ) capacitor c=0.00130622f \
 //x=51.63 //y=0 //x2=49.915 //y2=0.865
cc_181 ( N_GND_M30_noxref_d N_noxref_10_c_3904_n ) capacitor c=0.00257848f \
 //x=49.46 //y=0.865 //x2=49.915 //y2=0.865
cc_182 ( N_GND_M30_noxref_d N_noxref_10_c_3906_n ) capacitor c=0.00255985f \
 //x=49.46 //y=0.865 //x2=49.915 //y2=1.21
cc_183 ( N_GND_c_13_p N_noxref_10_M29_noxref_d ) capacitor c=0.00591582f \
 //x=48.47 //y=0 //x2=47.055 //y2=0.915
cc_184 ( N_GND_c_8_p N_noxref_11_c_4058_n ) capacitor c=0.0130885f //x=25.9 \
 //y=0 //x2=27.01 //y2=2.08
cc_185 ( N_GND_c_10_p N_noxref_11_c_4059_n ) capacitor c=5.78225e-19 //x=35.52 \
 //y=0 //x2=37.37 //y2=2.08
cc_186 ( N_GND_c_11_p N_noxref_11_c_4059_n ) capacitor c=5.32623e-19 //x=38.85 \
 //y=0 //x2=37.37 //y2=2.08
cc_187 ( N_GND_c_12_p N_noxref_11_c_4061_n ) capacitor c=0.0404734f //x=43.66 \
 //y=0 //x2=42.835 //y2=1.665
cc_188 ( N_GND_c_13_p N_noxref_11_c_4062_n ) capacitor c=5.41726e-19 //x=48.47 \
 //y=0 //x2=50.32 //y2=2.08
cc_189 ( N_GND_c_14_p N_noxref_11_c_4062_n ) capacitor c=5.32623e-19 //x=51.8 \
 //y=0 //x2=50.32 //y2=2.08
cc_190 ( N_GND_c_190_p N_noxref_11_c_4064_n ) capacitor c=0.00132755f \
 //x=26.89 //y=0 //x2=26.71 //y2=0.875
cc_191 ( N_GND_M16_noxref_d N_noxref_11_c_4064_n ) capacitor c=0.00211996f \
 //x=26.785 //y=0.875 //x2=26.71 //y2=0.875
cc_192 ( N_GND_M16_noxref_d N_noxref_11_c_4066_n ) capacitor c=0.00255985f \
 //x=26.785 //y=0.875 //x2=26.71 //y2=1.22
cc_193 ( N_GND_c_8_p N_noxref_11_c_4067_n ) capacitor c=0.00195164f //x=25.9 \
 //y=0 //x2=26.71 //y2=1.53
cc_194 ( N_GND_c_8_p N_noxref_11_c_4068_n ) capacitor c=0.0112696f //x=25.9 \
 //y=0 //x2=26.71 //y2=1.915
cc_195 ( N_GND_M16_noxref_d N_noxref_11_c_4069_n ) capacitor c=0.0131341f \
 //x=26.785 //y=0.875 //x2=27.085 //y2=0.72
cc_196 ( N_GND_M16_noxref_d N_noxref_11_c_4070_n ) capacitor c=0.00193146f \
 //x=26.785 //y=0.875 //x2=27.085 //y2=1.375
cc_197 ( N_GND_c_197_p N_noxref_11_c_4071_n ) capacitor c=0.00129018f \
 //x=30.54 //y=0 //x2=27.24 //y2=0.875
cc_198 ( N_GND_M16_noxref_d N_noxref_11_c_4071_n ) capacitor c=0.00257848f \
 //x=26.785 //y=0.875 //x2=27.24 //y2=0.875
cc_199 ( N_GND_M16_noxref_d N_noxref_11_c_4073_n ) capacitor c=0.00255985f \
 //x=26.785 //y=0.875 //x2=27.24 //y2=1.22
cc_200 ( N_GND_c_12_p N_noxref_11_M26_noxref_d ) capacitor c=0.00591582f \
 //x=43.66 //y=0 //x2=42.245 //y2=0.915
cc_201 ( N_GND_c_23_p N_D_c_4434_n ) capacitor c=0.104609f //x=86.95 //y=0 \
 //x2=32.815 //y2=2.59
cc_202 ( N_GND_c_4_p N_D_c_4434_n ) capacitor c=0.0238274f //x=9.62 //y=0 \
 //x2=32.815 //y2=2.59
cc_203 ( N_GND_c_5_p N_D_c_4434_n ) capacitor c=0.0238274f //x=12.95 //y=0 \
 //x2=32.815 //y2=2.59
cc_204 ( N_GND_c_6_p N_D_c_4434_n ) capacitor c=0.0254584f //x=17.76 //y=0 \
 //x2=32.815 //y2=2.59
cc_205 ( N_GND_c_7_p N_D_c_4434_n ) capacitor c=0.0215583f //x=22.57 //y=0 \
 //x2=32.815 //y2=2.59
cc_206 ( N_GND_c_8_p N_D_c_4434_n ) capacitor c=0.0215583f //x=25.9 //y=0 \
 //x2=32.815 //y2=2.59
cc_207 ( N_GND_c_9_p N_D_c_4434_n ) capacitor c=0.0215583f //x=30.71 //y=0 \
 //x2=32.815 //y2=2.59
cc_208 ( N_GND_c_23_p N_D_c_4441_n ) capacitor c=0.00219703f //x=86.95 //y=0 \
 //x2=7.145 //y2=2.59
cc_209 ( N_GND_c_10_p N_D_c_4442_n ) capacitor c=0.0215583f //x=35.52 //y=0 \
 //x2=58.715 //y2=2.59
cc_210 ( N_GND_c_11_p N_D_c_4442_n ) capacitor c=0.0215583f //x=38.85 //y=0 \
 //x2=58.715 //y2=2.59
cc_211 ( N_GND_c_12_p N_D_c_4442_n ) capacitor c=0.0215583f //x=43.66 //y=0 \
 //x2=58.715 //y2=2.59
cc_212 ( N_GND_c_13_p N_D_c_4442_n ) capacitor c=0.0215583f //x=48.47 //y=0 \
 //x2=58.715 //y2=2.59
cc_213 ( N_GND_c_14_p N_D_c_4442_n ) capacitor c=0.0215583f //x=51.8 //y=0 \
 //x2=58.715 //y2=2.59
cc_214 ( N_GND_c_15_p N_D_c_4442_n ) capacitor c=0.0215583f //x=56.61 //y=0 \
 //x2=58.715 //y2=2.59
cc_215 ( N_GND_c_3_p N_D_c_4448_n ) capacitor c=0.00101246f //x=4.81 //y=0 \
 //x2=7.03 //y2=2.08
cc_216 ( N_GND_c_9_p N_D_c_4449_n ) capacitor c=5.31163e-19 //x=30.71 //y=0 \
 //x2=32.93 //y2=2.08
cc_217 ( N_GND_c_15_p N_D_c_4450_n ) capacitor c=5.31163e-19 //x=56.61 //y=0 \
 //x2=58.83 //y2=2.08
cc_218 ( N_GND_c_1_p N_CLK_c_4802_n ) capacitor c=7.64246e-19 //x=0.74 //y=0 \
 //x2=2.22 //y2=2.08
cc_219 ( N_GND_c_5_p N_CLK_c_4803_n ) capacitor c=4.89793e-19 //x=12.95 //y=0 \
 //x2=15.17 //y2=2.08
cc_220 ( N_GND_c_8_p N_CLK_c_4804_n ) capacitor c=4.59642e-19 //x=25.9 //y=0 \
 //x2=28.12 //y2=2.08
cc_221 ( N_GND_c_11_p N_CLK_c_4805_n ) capacitor c=4.89793e-19 //x=38.85 //y=0 \
 //x2=41.07 //y2=2.08
cc_222 ( N_GND_c_14_p N_CLK_c_4806_n ) capacitor c=4.59642e-19 //x=51.8 //y=0 \
 //x2=54.02 //y2=2.08
cc_223 ( N_GND_c_17_p N_CLK_c_4807_n ) capacitor c=6.04789e-19 //x=64.75 //y=0 \
 //x2=66.97 //y2=2.08
cc_224 ( N_GND_c_15_p N_noxref_14_c_5587_n ) capacitor c=0.0406306f //x=56.61 \
 //y=0 //x2=55.785 //y2=1.665
cc_225 ( N_GND_c_15_p N_noxref_14_c_5588_n ) capacitor c=0.0129722f //x=56.61 \
 //y=0 //x2=57.72 //y2=2.08
cc_226 ( N_GND_c_18_p N_noxref_14_c_5589_n ) capacitor c=0.0155796f //x=69.56 \
 //y=0 //x2=70.67 //y2=2.08
cc_227 ( N_GND_c_227_p N_noxref_14_c_5590_n ) capacitor c=0.00132755f //x=57.6 \
 //y=0 //x2=57.42 //y2=0.875
cc_228 ( N_GND_M35_noxref_d N_noxref_14_c_5590_n ) capacitor c=0.00211996f \
 //x=57.495 //y=0.875 //x2=57.42 //y2=0.875
cc_229 ( N_GND_M35_noxref_d N_noxref_14_c_5592_n ) capacitor c=0.00255985f \
 //x=57.495 //y=0.875 //x2=57.42 //y2=1.22
cc_230 ( N_GND_c_15_p N_noxref_14_c_5593_n ) capacitor c=0.00204716f //x=56.61 \
 //y=0 //x2=57.42 //y2=1.53
cc_231 ( N_GND_c_15_p N_noxref_14_c_5594_n ) capacitor c=0.0110952f //x=56.61 \
 //y=0 //x2=57.42 //y2=1.915
cc_232 ( N_GND_M35_noxref_d N_noxref_14_c_5595_n ) capacitor c=0.0131341f \
 //x=57.495 //y=0.875 //x2=57.795 //y2=0.72
cc_233 ( N_GND_M35_noxref_d N_noxref_14_c_5596_n ) capacitor c=0.00193146f \
 //x=57.495 //y=0.875 //x2=57.795 //y2=1.375
cc_234 ( N_GND_c_234_p N_noxref_14_c_5597_n ) capacitor c=0.00129018f \
 //x=61.25 //y=0 //x2=57.95 //y2=0.875
cc_235 ( N_GND_M35_noxref_d N_noxref_14_c_5597_n ) capacitor c=0.00257848f \
 //x=57.495 //y=0.875 //x2=57.95 //y2=0.875
cc_236 ( N_GND_M35_noxref_d N_noxref_14_c_5599_n ) capacitor c=0.00255985f \
 //x=57.495 //y=0.875 //x2=57.95 //y2=1.22
cc_237 ( N_GND_c_237_p N_noxref_14_c_5600_n ) capacitor c=0.00132755f \
 //x=70.55 //y=0 //x2=70.37 //y2=0.875
cc_238 ( N_GND_M43_noxref_d N_noxref_14_c_5600_n ) capacitor c=0.00211996f \
 //x=70.445 //y=0.875 //x2=70.37 //y2=0.875
cc_239 ( N_GND_M43_noxref_d N_noxref_14_c_5602_n ) capacitor c=0.00255985f \
 //x=70.445 //y=0.875 //x2=70.37 //y2=1.22
cc_240 ( N_GND_c_18_p N_noxref_14_c_5603_n ) capacitor c=0.00204716f //x=69.56 \
 //y=0 //x2=70.37 //y2=1.53
cc_241 ( N_GND_c_18_p N_noxref_14_c_5604_n ) capacitor c=0.0110952f //x=69.56 \
 //y=0 //x2=70.37 //y2=1.915
cc_242 ( N_GND_M43_noxref_d N_noxref_14_c_5605_n ) capacitor c=0.0131341f \
 //x=70.445 //y=0.875 //x2=70.745 //y2=0.72
cc_243 ( N_GND_M43_noxref_d N_noxref_14_c_5606_n ) capacitor c=0.00193146f \
 //x=70.445 //y=0.875 //x2=70.745 //y2=1.375
cc_244 ( N_GND_c_244_p N_noxref_14_c_5607_n ) capacitor c=0.00129018f //x=74.2 \
 //y=0 //x2=70.9 //y2=0.875
cc_245 ( N_GND_M43_noxref_d N_noxref_14_c_5607_n ) capacitor c=0.00257848f \
 //x=70.445 //y=0.875 //x2=70.9 //y2=0.875
cc_246 ( N_GND_M43_noxref_d N_noxref_14_c_5609_n ) capacitor c=0.00255985f \
 //x=70.445 //y=0.875 //x2=70.9 //y2=1.22
cc_247 ( N_GND_c_15_p N_noxref_14_M34_noxref_d ) capacitor c=0.00591582f \
 //x=56.61 //y=0 //x2=55.195 //y2=0.915
cc_248 ( N_GND_c_23_p N_RN_c_5846_n ) capacitor c=0.0754427f //x=86.95 //y=0 \
 //x2=16.165 //y2=2.22
cc_249 ( N_GND_c_71_p N_RN_c_5846_n ) capacitor c=0.00318526f //x=9.45 //y=0 \
 //x2=16.165 //y2=2.22
cc_250 ( N_GND_c_32_p N_RN_c_5846_n ) capacitor c=0.00347653f //x=10.715 //y=0 \
 //x2=16.165 //y2=2.22
cc_251 ( N_GND_c_39_p N_RN_c_5846_n ) capacitor c=0.00411932f //x=12.78 //y=0 \
 //x2=16.165 //y2=2.22
cc_252 ( N_GND_c_47_p N_RN_c_5846_n ) capacitor c=0.00274252f //x=13.94 //y=0 \
 //x2=16.165 //y2=2.22
cc_253 ( N_GND_c_54_p N_RN_c_5846_n ) capacitor c=0.00111309f //x=17.59 //y=0 \
 //x2=16.165 //y2=2.22
cc_254 ( N_GND_c_4_p N_RN_c_5846_n ) capacitor c=0.0379964f //x=9.62 //y=0 \
 //x2=16.165 //y2=2.22
cc_255 ( N_GND_c_5_p N_RN_c_5846_n ) capacitor c=0.0379964f //x=12.95 //y=0 \
 //x2=16.165 //y2=2.22
cc_256 ( N_GND_c_23_p N_RN_c_5854_n ) capacitor c=0.00221055f //x=86.95 //y=0 \
 //x2=8.255 //y2=2.22
cc_257 ( N_GND_c_71_p N_RN_c_5854_n ) capacitor c=4.19033e-19 //x=9.45 //y=0 \
 //x2=8.255 //y2=2.22
cc_258 ( N_GND_c_23_p N_RN_c_5856_n ) capacitor c=0.0336613f //x=86.95 //y=0 \
 //x2=19.865 //y2=2.22
cc_259 ( N_GND_c_54_p N_RN_c_5856_n ) capacitor c=0.00318526f //x=17.59 //y=0 \
 //x2=19.865 //y2=2.22
cc_260 ( N_GND_c_74_p N_RN_c_5856_n ) capacitor c=0.00274252f //x=18.75 //y=0 \
 //x2=19.865 //y2=2.22
cc_261 ( N_GND_c_6_p N_RN_c_5856_n ) capacitor c=0.0379964f //x=17.76 //y=0 \
 //x2=19.865 //y2=2.22
cc_262 ( N_GND_c_23_p N_RN_c_5860_n ) capacitor c=0.00195247f //x=86.95 //y=0 \
 //x2=16.395 //y2=2.22
cc_263 ( N_GND_c_23_p N_RN_c_5861_n ) capacitor c=0.131484f //x=86.95 //y=0 \
 //x2=33.925 //y2=2.22
cc_264 ( N_GND_c_81_p N_RN_c_5861_n ) capacitor c=0.00447829f //x=22.4 //y=0 \
 //x2=33.925 //y2=2.22
cc_265 ( N_GND_c_105_p N_RN_c_5861_n ) capacitor c=0.00347653f //x=23.665 \
 //y=0 //x2=33.925 //y2=2.22
cc_266 ( N_GND_c_112_p N_RN_c_5861_n ) capacitor c=0.00411932f //x=25.73 //y=0 \
 //x2=33.925 //y2=2.22
cc_267 ( N_GND_c_190_p N_RN_c_5861_n ) capacitor c=0.00274252f //x=26.89 //y=0 \
 //x2=33.925 //y2=2.22
cc_268 ( N_GND_c_197_p N_RN_c_5861_n ) capacitor c=0.00450506f //x=30.54 //y=0 \
 //x2=33.925 //y2=2.22
cc_269 ( N_GND_c_150_p N_RN_c_5861_n ) capacitor c=0.00274252f //x=31.7 //y=0 \
 //x2=33.925 //y2=2.22
cc_270 ( N_GND_c_157_p N_RN_c_5861_n ) capacitor c=0.00111309f //x=35.35 //y=0 \
 //x2=33.925 //y2=2.22
cc_271 ( N_GND_c_7_p N_RN_c_5861_n ) capacitor c=0.0379964f //x=22.57 //y=0 \
 //x2=33.925 //y2=2.22
cc_272 ( N_GND_c_8_p N_RN_c_5861_n ) capacitor c=0.0379964f //x=25.9 //y=0 \
 //x2=33.925 //y2=2.22
cc_273 ( N_GND_c_9_p N_RN_c_5861_n ) capacitor c=0.0379964f //x=30.71 //y=0 \
 //x2=33.925 //y2=2.22
cc_274 ( N_GND_c_23_p N_RN_c_5872_n ) capacitor c=0.00168059f //x=86.95 //y=0 \
 //x2=20.095 //y2=2.22
cc_275 ( N_GND_c_23_p N_RN_c_5873_n ) capacitor c=0.0754427f //x=86.95 //y=0 \
 //x2=42.065 //y2=2.22
cc_276 ( N_GND_c_157_p N_RN_c_5873_n ) capacitor c=0.00318526f //x=35.35 //y=0 \
 //x2=42.065 //y2=2.22
cc_277 ( N_GND_c_120_p N_RN_c_5873_n ) capacitor c=0.00347653f //x=36.615 \
 //y=0 //x2=42.065 //y2=2.22
cc_278 ( N_GND_c_127_p N_RN_c_5873_n ) capacitor c=0.00411932f //x=38.68 //y=0 \
 //x2=42.065 //y2=2.22
cc_279 ( N_GND_c_134_p N_RN_c_5873_n ) capacitor c=0.00274252f //x=39.84 //y=0 \
 //x2=42.065 //y2=2.22
cc_280 ( N_GND_c_141_p N_RN_c_5873_n ) capacitor c=0.00111309f //x=43.49 //y=0 \
 //x2=42.065 //y2=2.22
cc_281 ( N_GND_c_10_p N_RN_c_5873_n ) capacitor c=0.0379964f //x=35.52 //y=0 \
 //x2=42.065 //y2=2.22
cc_282 ( N_GND_c_11_p N_RN_c_5873_n ) capacitor c=0.0379964f //x=38.85 //y=0 \
 //x2=42.065 //y2=2.22
cc_283 ( N_GND_c_23_p N_RN_c_5881_n ) capacitor c=0.00195247f //x=86.95 //y=0 \
 //x2=34.155 //y2=2.22
cc_284 ( N_GND_c_23_p N_RN_c_5882_n ) capacitor c=0.0336613f //x=86.95 //y=0 \
 //x2=45.765 //y2=2.22
cc_285 ( N_GND_c_141_p N_RN_c_5882_n ) capacitor c=0.00318526f //x=43.49 //y=0 \
 //x2=45.765 //y2=2.22
cc_286 ( N_GND_c_160_p N_RN_c_5882_n ) capacitor c=0.00274252f //x=44.65 //y=0 \
 //x2=45.765 //y2=2.22
cc_287 ( N_GND_c_12_p N_RN_c_5882_n ) capacitor c=0.0379964f //x=43.66 //y=0 \
 //x2=45.765 //y2=2.22
cc_288 ( N_GND_c_23_p N_RN_c_5886_n ) capacitor c=0.00195247f //x=86.95 //y=0 \
 //x2=42.295 //y2=2.22
cc_289 ( N_GND_c_23_p N_RN_c_5887_n ) capacitor c=0.131484f //x=86.95 //y=0 \
 //x2=59.825 //y2=2.22
cc_290 ( N_GND_c_167_p N_RN_c_5887_n ) capacitor c=0.00447829f //x=48.3 //y=0 \
 //x2=59.825 //y2=2.22
cc_291 ( N_GND_c_173_p N_RN_c_5887_n ) capacitor c=0.00347653f //x=49.565 \
 //y=0 //x2=59.825 //y2=2.22
cc_292 ( N_GND_c_180_p N_RN_c_5887_n ) capacitor c=0.00411932f //x=51.63 //y=0 \
 //x2=59.825 //y2=2.22
cc_293 ( N_GND_c_293_p N_RN_c_5887_n ) capacitor c=0.00274252f //x=52.79 //y=0 \
 //x2=59.825 //y2=2.22
cc_294 ( N_GND_c_294_p N_RN_c_5887_n ) capacitor c=0.00450506f //x=56.44 //y=0 \
 //x2=59.825 //y2=2.22
cc_295 ( N_GND_c_227_p N_RN_c_5887_n ) capacitor c=0.00274252f //x=57.6 //y=0 \
 //x2=59.825 //y2=2.22
cc_296 ( N_GND_c_234_p N_RN_c_5887_n ) capacitor c=0.00111309f //x=61.25 //y=0 \
 //x2=59.825 //y2=2.22
cc_297 ( N_GND_c_13_p N_RN_c_5887_n ) capacitor c=0.0379964f //x=48.47 //y=0 \
 //x2=59.825 //y2=2.22
cc_298 ( N_GND_c_14_p N_RN_c_5887_n ) capacitor c=0.0379964f //x=51.8 //y=0 \
 //x2=59.825 //y2=2.22
cc_299 ( N_GND_c_15_p N_RN_c_5887_n ) capacitor c=0.0379964f //x=56.61 //y=0 \
 //x2=59.825 //y2=2.22
cc_300 ( N_GND_c_23_p N_RN_c_5898_n ) capacitor c=0.00168059f //x=86.95 //y=0 \
 //x2=45.995 //y2=2.22
cc_301 ( N_GND_c_23_p N_RN_c_5899_n ) capacitor c=0.0754427f //x=86.95 //y=0 \
 //x2=67.965 //y2=2.22
cc_302 ( N_GND_c_234_p N_RN_c_5899_n ) capacitor c=0.00318526f //x=61.25 //y=0 \
 //x2=67.965 //y2=2.22
cc_303 ( N_GND_c_303_p N_RN_c_5899_n ) capacitor c=0.00347653f //x=62.515 \
 //y=0 //x2=67.965 //y2=2.22
cc_304 ( N_GND_c_304_p N_RN_c_5899_n ) capacitor c=0.00411932f //x=64.58 //y=0 \
 //x2=67.965 //y2=2.22
cc_305 ( N_GND_c_305_p N_RN_c_5899_n ) capacitor c=0.00274252f //x=65.74 //y=0 \
 //x2=67.965 //y2=2.22
cc_306 ( N_GND_c_306_p N_RN_c_5899_n ) capacitor c=0.00111309f //x=69.39 //y=0 \
 //x2=67.965 //y2=2.22
cc_307 ( N_GND_c_16_p N_RN_c_5899_n ) capacitor c=0.0401775f //x=61.42 //y=0 \
 //x2=67.965 //y2=2.22
cc_308 ( N_GND_c_17_p N_RN_c_5899_n ) capacitor c=0.0401775f //x=64.75 //y=0 \
 //x2=67.965 //y2=2.22
cc_309 ( N_GND_c_23_p N_RN_c_5907_n ) capacitor c=0.00195247f //x=86.95 //y=0 \
 //x2=60.055 //y2=2.22
cc_310 ( N_GND_c_23_p N_RN_c_5908_n ) capacitor c=0.0355717f //x=86.95 //y=0 \
 //x2=71.665 //y2=2.22
cc_311 ( N_GND_c_306_p N_RN_c_5908_n ) capacitor c=0.00318526f //x=69.39 //y=0 \
 //x2=71.665 //y2=2.22
cc_312 ( N_GND_c_237_p N_RN_c_5908_n ) capacitor c=0.00274252f //x=70.55 //y=0 \
 //x2=71.665 //y2=2.22
cc_313 ( N_GND_c_18_p N_RN_c_5908_n ) capacitor c=0.0401775f //x=69.56 //y=0 \
 //x2=71.665 //y2=2.22
cc_314 ( N_GND_c_23_p N_RN_c_5912_n ) capacitor c=0.00195247f //x=86.95 //y=0 \
 //x2=68.195 //y2=2.22
cc_315 ( N_GND_c_4_p N_RN_c_5913_n ) capacitor c=6.79203e-19 //x=9.62 //y=0 \
 //x2=8.14 //y2=2.08
cc_316 ( N_GND_c_6_p N_RN_c_5914_n ) capacitor c=5.93203e-19 //x=17.76 //y=0 \
 //x2=16.28 //y2=2.08
cc_317 ( N_GND_c_6_p N_RN_c_5915_n ) capacitor c=4.79163e-19 //x=17.76 //y=0 \
 //x2=19.98 //y2=2.08
cc_318 ( N_GND_c_10_p N_RN_c_5916_n ) capacitor c=6.79203e-19 //x=35.52 //y=0 \
 //x2=34.04 //y2=2.08
cc_319 ( N_GND_c_12_p N_RN_c_5917_n ) capacitor c=5.93203e-19 //x=43.66 //y=0 \
 //x2=42.18 //y2=2.08
cc_320 ( N_GND_c_12_p N_RN_c_5918_n ) capacitor c=4.79163e-19 //x=43.66 //y=0 \
 //x2=45.88 //y2=2.08
cc_321 ( N_GND_c_16_p N_RN_c_5919_n ) capacitor c=0.0011655f //x=61.42 //y=0 \
 //x2=59.94 //y2=2.08
cc_322 ( N_GND_c_18_p N_RN_c_5920_n ) capacitor c=8.37259e-19 //x=69.56 //y=0 \
 //x2=68.08 //y2=2.08
cc_323 ( N_GND_c_18_p N_RN_c_5921_n ) capacitor c=5.94159e-19 //x=69.56 //y=0 \
 //x2=71.78 //y2=2.08
cc_324 ( N_GND_c_14_p N_noxref_16_c_6801_n ) capacitor c=0.0130885f //x=51.8 \
 //y=0 //x2=52.91 //y2=2.08
cc_325 ( N_GND_c_16_p N_noxref_16_c_6802_n ) capacitor c=7.4738e-19 //x=61.42 \
 //y=0 //x2=63.27 //y2=2.08
cc_326 ( N_GND_c_17_p N_noxref_16_c_6802_n ) capacitor c=7.76678e-19 //x=64.75 \
 //y=0 //x2=63.27 //y2=2.08
cc_327 ( N_GND_c_18_p N_noxref_16_c_6804_n ) capacitor c=0.0430857f //x=69.56 \
 //y=0 //x2=68.735 //y2=1.665
cc_328 ( N_GND_c_19_p N_noxref_16_c_6805_n ) capacitor c=0.0455978f //x=74.37 \
 //y=0 //x2=73.545 //y2=1.665
cc_329 ( N_GND_c_19_p N_noxref_16_c_6806_n ) capacitor c=0.0179404f //x=74.37 \
 //y=0 //x2=75.48 //y2=2.08
cc_330 ( N_GND_c_19_p N_noxref_16_c_6807_n ) capacitor c=9.2064e-19 //x=74.37 \
 //y=0 //x2=76.22 //y2=2.08
cc_331 ( N_GND_c_20_p N_noxref_16_c_6807_n ) capacitor c=9.53263e-19 //x=77.7 \
 //y=0 //x2=76.22 //y2=2.08
cc_332 ( N_GND_c_293_p N_noxref_16_c_6809_n ) capacitor c=0.00132755f \
 //x=52.79 //y=0 //x2=52.61 //y2=0.875
cc_333 ( N_GND_M32_noxref_d N_noxref_16_c_6809_n ) capacitor c=0.00211996f \
 //x=52.685 //y=0.875 //x2=52.61 //y2=0.875
cc_334 ( N_GND_M32_noxref_d N_noxref_16_c_6811_n ) capacitor c=0.00255985f \
 //x=52.685 //y=0.875 //x2=52.61 //y2=1.22
cc_335 ( N_GND_c_14_p N_noxref_16_c_6812_n ) capacitor c=0.00195164f //x=51.8 \
 //y=0 //x2=52.61 //y2=1.53
cc_336 ( N_GND_c_14_p N_noxref_16_c_6813_n ) capacitor c=0.0112696f //x=51.8 \
 //y=0 //x2=52.61 //y2=1.915
cc_337 ( N_GND_M32_noxref_d N_noxref_16_c_6814_n ) capacitor c=0.0131341f \
 //x=52.685 //y=0.875 //x2=52.985 //y2=0.72
cc_338 ( N_GND_M32_noxref_d N_noxref_16_c_6815_n ) capacitor c=0.00193146f \
 //x=52.685 //y=0.875 //x2=52.985 //y2=1.375
cc_339 ( N_GND_c_294_p N_noxref_16_c_6816_n ) capacitor c=0.00129018f \
 //x=56.44 //y=0 //x2=53.14 //y2=0.875
cc_340 ( N_GND_M32_noxref_d N_noxref_16_c_6816_n ) capacitor c=0.00257848f \
 //x=52.685 //y=0.875 //x2=53.14 //y2=0.875
cc_341 ( N_GND_M32_noxref_d N_noxref_16_c_6818_n ) capacitor c=0.00255985f \
 //x=52.685 //y=0.875 //x2=53.14 //y2=1.22
cc_342 ( N_GND_c_342_p N_noxref_16_c_6819_n ) capacitor c=0.00135046f \
 //x=75.465 //y=0 //x2=75.285 //y2=0.865
cc_343 ( N_GND_M46_noxref_d N_noxref_16_c_6819_n ) capacitor c=0.00220047f \
 //x=75.36 //y=0.865 //x2=75.285 //y2=0.865
cc_344 ( N_GND_M46_noxref_d N_noxref_16_c_6821_n ) capacitor c=0.00255985f \
 //x=75.36 //y=0.865 //x2=75.285 //y2=1.21
cc_345 ( N_GND_c_19_p N_noxref_16_c_6822_n ) capacitor c=0.00189421f //x=74.37 \
 //y=0 //x2=75.285 //y2=1.52
cc_346 ( N_GND_c_19_p N_noxref_16_c_6823_n ) capacitor c=0.0106743f //x=74.37 \
 //y=0 //x2=75.285 //y2=1.915
cc_347 ( N_GND_M46_noxref_d N_noxref_16_c_6824_n ) capacitor c=0.0131326f \
 //x=75.36 //y=0.865 //x2=75.66 //y2=0.71
cc_348 ( N_GND_M46_noxref_d N_noxref_16_c_6825_n ) capacitor c=0.00193127f \
 //x=75.36 //y=0.865 //x2=75.66 //y2=1.365
cc_349 ( N_GND_c_349_p N_noxref_16_c_6826_n ) capacitor c=0.00130622f \
 //x=77.53 //y=0 //x2=75.815 //y2=0.865
cc_350 ( N_GND_M46_noxref_d N_noxref_16_c_6826_n ) capacitor c=0.00257848f \
 //x=75.36 //y=0.865 //x2=75.815 //y2=0.865
cc_351 ( N_GND_M46_noxref_d N_noxref_16_c_6828_n ) capacitor c=0.00255985f \
 //x=75.36 //y=0.865 //x2=75.815 //y2=1.21
cc_352 ( N_GND_c_18_p N_noxref_16_M42_noxref_d ) capacitor c=0.00591582f \
 //x=69.56 //y=0 //x2=68.145 //y2=0.915
cc_353 ( N_GND_c_19_p N_noxref_16_M45_noxref_d ) capacitor c=0.00591582f \
 //x=74.37 //y=0 //x2=72.955 //y2=0.915
cc_354 ( N_GND_c_13_p N_noxref_17_c_7301_n ) capacitor c=6.18623e-19 //x=48.47 \
 //y=0 //x2=46.99 //y2=2.08
cc_355 ( N_GND_c_14_p N_noxref_17_c_7302_n ) capacitor c=0.0410119f //x=51.8 \
 //y=0 //x2=50.975 //y2=1.655
cc_356 ( N_GND_c_13_p N_noxref_17_c_7303_n ) capacitor c=9.64732e-19 //x=48.47 \
 //y=0 //x2=51.06 //y2=3.33
cc_357 ( N_GND_c_15_p N_noxref_17_c_7304_n ) capacitor c=5.32623e-19 //x=56.61 \
 //y=0 //x2=55.13 //y2=2.08
cc_358 ( N_GND_c_16_p N_noxref_17_c_7305_n ) capacitor c=0.0428194f //x=61.42 \
 //y=0 //x2=60.595 //y2=1.665
cc_359 ( N_GND_c_16_p N_noxref_17_c_7306_n ) capacitor c=0.0156446f //x=61.42 \
 //y=0 //x2=62.53 //y2=2.08
cc_360 ( N_GND_c_17_p N_noxref_17_c_7307_n ) capacitor c=0.0436242f //x=64.75 \
 //y=0 //x2=63.925 //y2=1.655
cc_361 ( N_GND_c_16_p N_noxref_17_c_7308_n ) capacitor c=9.64732e-19 //x=61.42 \
 //y=0 //x2=64.01 //y2=3.33
cc_362 ( N_GND_c_17_p N_noxref_17_c_7309_n ) capacitor c=0.0156442f //x=64.75 \
 //y=0 //x2=65.86 //y2=2.08
cc_363 ( N_GND_c_23_p N_noxref_17_c_7310_n ) capacitor c=2.98913e-19 //x=86.95 \
 //y=0 //x2=78.44 //y2=2.08
cc_364 ( N_GND_c_20_p N_noxref_17_c_7310_n ) capacitor c=0.0292135f //x=77.7 \
 //y=0 //x2=78.44 //y2=2.08
cc_365 ( N_GND_c_21_p N_noxref_17_c_7310_n ) capacitor c=3.10504e-19 //x=81.03 \
 //y=0 //x2=78.44 //y2=2.08
cc_366 ( N_GND_c_21_p N_noxref_17_c_7313_n ) capacitor c=0.0178945f //x=81.03 \
 //y=0 //x2=82.14 //y2=2.08
cc_367 ( N_GND_c_22_p N_noxref_17_c_7313_n ) capacitor c=7.87427e-19 //x=84.36 \
 //y=0 //x2=82.14 //y2=2.08
cc_368 ( N_GND_c_303_p N_noxref_17_c_7315_n ) capacitor c=0.00135046f \
 //x=62.515 //y=0 //x2=62.335 //y2=0.865
cc_369 ( N_GND_M38_noxref_d N_noxref_17_c_7315_n ) capacitor c=0.00220047f \
 //x=62.41 //y=0.865 //x2=62.335 //y2=0.865
cc_370 ( N_GND_M38_noxref_d N_noxref_17_c_7317_n ) capacitor c=0.00255985f \
 //x=62.41 //y=0.865 //x2=62.335 //y2=1.21
cc_371 ( N_GND_c_16_p N_noxref_17_c_7318_n ) capacitor c=0.00189421f //x=61.42 \
 //y=0 //x2=62.335 //y2=1.52
cc_372 ( N_GND_c_16_p N_noxref_17_c_7319_n ) capacitor c=0.00992619f //x=61.42 \
 //y=0 //x2=62.335 //y2=1.915
cc_373 ( N_GND_M38_noxref_d N_noxref_17_c_7320_n ) capacitor c=0.0131326f \
 //x=62.41 //y=0.865 //x2=62.71 //y2=0.71
cc_374 ( N_GND_M38_noxref_d N_noxref_17_c_7321_n ) capacitor c=0.00193127f \
 //x=62.41 //y=0.865 //x2=62.71 //y2=1.365
cc_375 ( N_GND_c_304_p N_noxref_17_c_7322_n ) capacitor c=0.00130622f \
 //x=64.58 //y=0 //x2=62.865 //y2=0.865
cc_376 ( N_GND_M38_noxref_d N_noxref_17_c_7322_n ) capacitor c=0.00257848f \
 //x=62.41 //y=0.865 //x2=62.865 //y2=0.865
cc_377 ( N_GND_M38_noxref_d N_noxref_17_c_7324_n ) capacitor c=0.00255985f \
 //x=62.41 //y=0.865 //x2=62.865 //y2=1.21
cc_378 ( N_GND_c_305_p N_noxref_17_c_7325_n ) capacitor c=0.00132755f \
 //x=65.74 //y=0 //x2=65.56 //y2=0.875
cc_379 ( N_GND_M40_noxref_d N_noxref_17_c_7325_n ) capacitor c=0.00211996f \
 //x=65.635 //y=0.875 //x2=65.56 //y2=0.875
cc_380 ( N_GND_M40_noxref_d N_noxref_17_c_7327_n ) capacitor c=0.00255985f \
 //x=65.635 //y=0.875 //x2=65.56 //y2=1.22
cc_381 ( N_GND_c_17_p N_noxref_17_c_7328_n ) capacitor c=0.00195164f //x=64.75 \
 //y=0 //x2=65.56 //y2=1.53
cc_382 ( N_GND_c_17_p N_noxref_17_c_7329_n ) capacitor c=0.0110952f //x=64.75 \
 //y=0 //x2=65.56 //y2=1.915
cc_383 ( N_GND_M40_noxref_d N_noxref_17_c_7330_n ) capacitor c=0.0131341f \
 //x=65.635 //y=0.875 //x2=65.935 //y2=0.72
cc_384 ( N_GND_M40_noxref_d N_noxref_17_c_7331_n ) capacitor c=0.00193146f \
 //x=65.635 //y=0.875 //x2=65.935 //y2=1.375
cc_385 ( N_GND_c_306_p N_noxref_17_c_7332_n ) capacitor c=0.00129018f \
 //x=69.39 //y=0 //x2=66.09 //y2=0.875
cc_386 ( N_GND_M40_noxref_d N_noxref_17_c_7332_n ) capacitor c=0.00257848f \
 //x=65.635 //y=0.875 //x2=66.09 //y2=0.875
cc_387 ( N_GND_M40_noxref_d N_noxref_17_c_7334_n ) capacitor c=0.00255985f \
 //x=65.635 //y=0.875 //x2=66.09 //y2=1.22
cc_388 ( N_GND_c_388_p N_noxref_17_c_7335_n ) capacitor c=0.0013864f \
 //x=78.795 //y=0 //x2=78.615 //y2=0.865
cc_389 ( N_GND_M48_noxref_d N_noxref_17_c_7335_n ) capacitor c=0.00220047f \
 //x=78.69 //y=0.865 //x2=78.615 //y2=0.865
cc_390 ( N_GND_M48_noxref_d N_noxref_17_c_7337_n ) capacitor c=0.00255985f \
 //x=78.69 //y=0.865 //x2=78.615 //y2=1.21
cc_391 ( N_GND_c_20_p N_noxref_17_c_7338_n ) capacitor c=0.0018059f //x=77.7 \
 //y=0 //x2=78.615 //y2=1.52
cc_392 ( N_GND_c_20_p N_noxref_17_c_7339_n ) capacitor c=0.00369987f //x=77.7 \
 //y=0 //x2=78.615 //y2=1.915
cc_393 ( N_GND_M48_noxref_d N_noxref_17_c_7340_n ) capacitor c=0.0131326f \
 //x=78.69 //y=0.865 //x2=78.99 //y2=0.71
cc_394 ( N_GND_M48_noxref_d N_noxref_17_c_7341_n ) capacitor c=0.00193127f \
 //x=78.69 //y=0.865 //x2=78.99 //y2=1.365
cc_395 ( N_GND_c_395_p N_noxref_17_c_7342_n ) capacitor c=0.00130622f \
 //x=80.86 //y=0 //x2=79.145 //y2=0.865
cc_396 ( N_GND_M48_noxref_d N_noxref_17_c_7342_n ) capacitor c=0.00257848f \
 //x=78.69 //y=0.865 //x2=79.145 //y2=0.865
cc_397 ( N_GND_M48_noxref_d N_noxref_17_c_7344_n ) capacitor c=0.00255985f \
 //x=78.69 //y=0.865 //x2=79.145 //y2=1.21
cc_398 ( N_GND_c_398_p N_noxref_17_c_7345_n ) capacitor c=0.00135046f \
 //x=82.125 //y=0 //x2=81.945 //y2=0.865
cc_399 ( N_GND_M50_noxref_d N_noxref_17_c_7345_n ) capacitor c=0.00220047f \
 //x=82.02 //y=0.865 //x2=81.945 //y2=0.865
cc_400 ( N_GND_M50_noxref_d N_noxref_17_c_7347_n ) capacitor c=0.00272336f \
 //x=82.02 //y=0.865 //x2=81.945 //y2=1.21
cc_401 ( N_GND_c_21_p N_noxref_17_c_7348_n ) capacitor c=0.0100605f //x=81.03 \
 //y=0 //x2=81.945 //y2=1.915
cc_402 ( N_GND_M50_noxref_d N_noxref_17_c_7349_n ) capacitor c=0.0131326f \
 //x=82.02 //y=0.865 //x2=82.32 //y2=0.71
cc_403 ( N_GND_M50_noxref_d N_noxref_17_c_7350_n ) capacitor c=0.00167494f \
 //x=82.02 //y=0.865 //x2=82.32 //y2=1.365
cc_404 ( N_GND_c_404_p N_noxref_17_c_7351_n ) capacitor c=0.00130622f \
 //x=84.19 //y=0 //x2=82.475 //y2=0.865
cc_405 ( N_GND_M50_noxref_d N_noxref_17_c_7351_n ) capacitor c=0.00257848f \
 //x=82.02 //y=0.865 //x2=82.475 //y2=0.865
cc_406 ( N_GND_M50_noxref_d N_noxref_17_c_7353_n ) capacitor c=0.00272336f \
 //x=82.02 //y=0.865 //x2=82.475 //y2=1.21
cc_407 ( N_GND_c_20_p N_noxref_17_c_7354_n ) capacitor c=0.01092f //x=77.7 \
 //y=0 //x2=78.44 //y2=2.08
cc_408 ( N_GND_c_13_p N_noxref_17_M31_noxref_d ) capacitor c=8.58106e-19 \
 //x=48.47 //y=0 //x2=50.43 //y2=0.905
cc_409 ( N_GND_c_14_p N_noxref_17_M31_noxref_d ) capacitor c=0.00616547f \
 //x=51.8 //y=0 //x2=50.43 //y2=0.905
cc_410 ( N_GND_M30_noxref_d N_noxref_17_M31_noxref_d ) capacitor c=0.00143464f \
 //x=49.46 //y=0.865 //x2=50.43 //y2=0.905
cc_411 ( N_GND_c_16_p N_noxref_17_M37_noxref_d ) capacitor c=0.00591582f \
 //x=61.42 //y=0 //x2=60.005 //y2=0.915
cc_412 ( N_GND_c_16_p N_noxref_17_M39_noxref_d ) capacitor c=8.58106e-19 \
 //x=61.42 //y=0 //x2=63.38 //y2=0.905
cc_413 ( N_GND_c_17_p N_noxref_17_M39_noxref_d ) capacitor c=0.00616547f \
 //x=64.75 //y=0 //x2=63.38 //y2=0.905
cc_414 ( N_GND_M38_noxref_d N_noxref_17_M39_noxref_d ) capacitor c=0.00143464f \
 //x=62.41 //y=0.865 //x2=63.38 //y2=0.905
cc_415 ( N_GND_c_22_p N_noxref_18_c_8064_n ) capacitor c=0.00281233f //x=84.36 \
 //y=0 //x2=86.095 //y2=4.07
cc_416 ( N_GND_c_19_p N_noxref_18_c_8065_n ) capacitor c=0.00128267f //x=74.37 \
 //y=0 //x2=72.89 //y2=2.08
cc_417 ( N_GND_c_20_p N_noxref_18_c_8066_n ) capacitor c=0.0462119f //x=77.7 \
 //y=0 //x2=76.875 //y2=1.655
cc_418 ( N_GND_c_19_p N_noxref_18_c_8067_n ) capacitor c=9.64732e-19 //x=74.37 \
 //y=0 //x2=76.96 //y2=3.7
cc_419 ( N_GND_c_20_p N_noxref_18_c_8068_n ) capacitor c=0.00123238f //x=77.7 \
 //y=0 //x2=79.55 //y2=2.08
cc_420 ( N_GND_c_21_p N_noxref_18_c_8068_n ) capacitor c=0.0125771f //x=81.03 \
 //y=0 //x2=79.55 //y2=2.08
cc_421 ( N_GND_c_2_p N_noxref_18_c_8070_n ) capacitor c=0.00128267f //x=86.95 \
 //y=0 //x2=86.21 //y2=2.08
cc_422 ( N_GND_c_22_p N_noxref_18_c_8070_n ) capacitor c=8.50308e-19 //x=84.36 \
 //y=0 //x2=86.21 //y2=2.08
cc_423 ( N_GND_c_21_p N_noxref_18_c_8072_n ) capacitor c=2.63786e-19 //x=81.03 \
 //y=0 //x2=79.55 //y2=2.08
cc_424 ( N_GND_c_19_p N_noxref_18_M47_noxref_d ) capacitor c=8.58106e-19 \
 //x=74.37 //y=0 //x2=76.33 //y2=0.905
cc_425 ( N_GND_c_20_p N_noxref_18_M47_noxref_d ) capacitor c=0.00616146f \
 //x=77.7 //y=0 //x2=76.33 //y2=0.905
cc_426 ( N_GND_M46_noxref_d N_noxref_18_M47_noxref_d ) capacitor c=0.00143464f \
 //x=75.36 //y=0.865 //x2=76.33 //y2=0.905
cc_427 ( N_GND_c_7_p N_noxref_20_c_8515_n ) capacitor c=0.00750857f //x=22.57 \
 //y=0 //x2=25.045 //y2=2.96
cc_428 ( N_GND_c_23_p N_noxref_20_c_8516_n ) capacitor c=0.0892844f //x=86.95 \
 //y=0 //x2=83.505 //y2=2.96
cc_429 ( N_GND_c_244_p N_noxref_20_c_8516_n ) capacitor c=0.00282695f //x=74.2 \
 //y=0 //x2=83.505 //y2=2.96
cc_430 ( N_GND_c_342_p N_noxref_20_c_8516_n ) capacitor c=0.00233429f \
 //x=75.465 //y=0 //x2=83.505 //y2=2.96
cc_431 ( N_GND_c_349_p N_noxref_20_c_8516_n ) capacitor c=0.00272473f \
 //x=77.53 //y=0 //x2=83.505 //y2=2.96
cc_432 ( N_GND_c_388_p N_noxref_20_c_8516_n ) capacitor c=0.0019279f \
 //x=78.795 //y=0 //x2=83.505 //y2=2.96
cc_433 ( N_GND_c_395_p N_noxref_20_c_8516_n ) capacitor c=6.3489e-19 //x=80.86 \
 //y=0 //x2=83.505 //y2=2.96
cc_434 ( N_GND_c_8_p N_noxref_20_c_8516_n ) capacitor c=0.00750857f //x=25.9 \
 //y=0 //x2=83.505 //y2=2.96
cc_435 ( N_GND_c_9_p N_noxref_20_c_8516_n ) capacitor c=0.00750857f //x=30.71 \
 //y=0 //x2=83.505 //y2=2.96
cc_436 ( N_GND_c_10_p N_noxref_20_c_8516_n ) capacitor c=0.00750857f //x=35.52 \
 //y=0 //x2=83.505 //y2=2.96
cc_437 ( N_GND_c_11_p N_noxref_20_c_8516_n ) capacitor c=0.00750857f //x=38.85 \
 //y=0 //x2=83.505 //y2=2.96
cc_438 ( N_GND_c_12_p N_noxref_20_c_8516_n ) capacitor c=0.00750857f //x=43.66 \
 //y=0 //x2=83.505 //y2=2.96
cc_439 ( N_GND_c_13_p N_noxref_20_c_8516_n ) capacitor c=0.00750857f //x=48.47 \
 //y=0 //x2=83.505 //y2=2.96
cc_440 ( N_GND_c_14_p N_noxref_20_c_8516_n ) capacitor c=0.00750857f //x=51.8 \
 //y=0 //x2=83.505 //y2=2.96
cc_441 ( N_GND_c_15_p N_noxref_20_c_8516_n ) capacitor c=0.00750857f //x=56.61 \
 //y=0 //x2=83.505 //y2=2.96
cc_442 ( N_GND_c_16_p N_noxref_20_c_8516_n ) capacitor c=0.00949826f //x=61.42 \
 //y=0 //x2=83.505 //y2=2.96
cc_443 ( N_GND_c_17_p N_noxref_20_c_8516_n ) capacitor c=0.00949826f //x=64.75 \
 //y=0 //x2=83.505 //y2=2.96
cc_444 ( N_GND_c_18_p N_noxref_20_c_8516_n ) capacitor c=0.00949826f //x=69.56 \
 //y=0 //x2=83.505 //y2=2.96
cc_445 ( N_GND_c_19_p N_noxref_20_c_8516_n ) capacitor c=0.0144849f //x=74.37 \
 //y=0 //x2=83.505 //y2=2.96
cc_446 ( N_GND_c_20_p N_noxref_20_c_8516_n ) capacitor c=0.0144849f //x=77.7 \
 //y=0 //x2=83.505 //y2=2.96
cc_447 ( N_GND_c_21_p N_noxref_20_c_8516_n ) capacitor c=0.0128764f //x=81.03 \
 //y=0 //x2=83.505 //y2=2.96
cc_448 ( N_GND_c_22_p N_noxref_20_c_8536_n ) capacitor c=0.0396043f //x=84.36 \
 //y=0 //x2=84.985 //y2=2.08
cc_449 ( N_GND_c_22_p N_noxref_20_c_8537_n ) capacitor c=0.00128384f //x=84.36 \
 //y=0 //x2=83.735 //y2=2.08
cc_450 ( N_GND_c_7_p N_noxref_20_c_8538_n ) capacitor c=6.18623e-19 //x=22.57 \
 //y=0 //x2=21.09 //y2=2.08
cc_451 ( N_GND_c_8_p N_noxref_20_c_8539_n ) capacitor c=0.0410119f //x=25.9 \
 //y=0 //x2=25.075 //y2=1.655
cc_452 ( N_GND_c_7_p N_noxref_20_c_8540_n ) capacitor c=9.64732e-19 //x=22.57 \
 //y=0 //x2=25.16 //y2=2.96
cc_453 ( N_GND_c_21_p N_noxref_20_c_8541_n ) capacitor c=6.95291e-19 //x=81.03 \
 //y=0 //x2=83.62 //y2=2.08
cc_454 ( N_GND_c_22_p N_noxref_20_c_8541_n ) capacitor c=0.0266762f //x=84.36 \
 //y=0 //x2=83.62 //y2=2.08
cc_455 ( N_GND_c_22_p N_noxref_20_c_8543_n ) capacitor c=0.0272331f //x=84.36 \
 //y=0 //x2=85.1 //y2=2.08
cc_456 ( N_GND_c_22_p N_noxref_20_c_8544_n ) capacitor c=0.0103285f //x=84.36 \
 //y=0 //x2=83.445 //y2=1.915
cc_457 ( N_GND_c_457_p N_noxref_20_c_8545_n ) capacitor c=0.0013864f \
 //x=85.455 //y=0 //x2=85.275 //y2=0.865
cc_458 ( N_GND_M52_noxref_d N_noxref_20_c_8545_n ) capacitor c=0.00220047f \
 //x=85.35 //y=0.865 //x2=85.275 //y2=0.865
cc_459 ( N_GND_M52_noxref_d N_noxref_20_c_8547_n ) capacitor c=0.00272336f \
 //x=85.35 //y=0.865 //x2=85.275 //y2=1.21
cc_460 ( N_GND_c_22_p N_noxref_20_c_8548_n ) capacitor c=0.00369763f //x=84.36 \
 //y=0 //x2=85.275 //y2=1.915
cc_461 ( N_GND_M52_noxref_d N_noxref_20_c_8549_n ) capacitor c=0.0131326f \
 //x=85.35 //y=0.865 //x2=85.65 //y2=0.71
cc_462 ( N_GND_M52_noxref_d N_noxref_20_c_8550_n ) capacitor c=0.00167494f \
 //x=85.35 //y=0.865 //x2=85.65 //y2=1.365
cc_463 ( N_GND_c_2_p N_noxref_20_c_8551_n ) capacitor c=0.00130622f //x=86.95 \
 //y=0 //x2=85.805 //y2=0.865
cc_464 ( N_GND_M52_noxref_d N_noxref_20_c_8551_n ) capacitor c=0.00257848f \
 //x=85.35 //y=0.865 //x2=85.805 //y2=0.865
cc_465 ( N_GND_M52_noxref_d N_noxref_20_c_8553_n ) capacitor c=0.00272336f \
 //x=85.35 //y=0.865 //x2=85.805 //y2=1.21
cc_466 ( N_GND_c_22_p N_noxref_20_c_8554_n ) capacitor c=0.00564759f //x=84.36 \
 //y=0 //x2=85.1 //y2=2.08
cc_467 ( N_GND_c_7_p N_noxref_20_M15_noxref_d ) capacitor c=8.58106e-19 \
 //x=22.57 //y=0 //x2=24.53 //y2=0.905
cc_468 ( N_GND_c_8_p N_noxref_20_M15_noxref_d ) capacitor c=0.00616547f \
 //x=25.9 //y=0 //x2=24.53 //y2=0.905
cc_469 ( N_GND_M14_noxref_d N_noxref_20_M15_noxref_d ) capacitor c=0.00143464f \
 //x=23.56 //y=0.865 //x2=24.53 //y2=0.905
cc_470 ( N_GND_c_23_p N_QN_c_9097_n ) capacitor c=0.0695894f //x=86.95 //y=0 \
 //x2=83.065 //y2=1.18
cc_471 ( N_GND_c_395_p N_QN_c_9097_n ) capacitor c=0.0081414f //x=80.86 //y=0 \
 //x2=83.065 //y2=1.18
cc_472 ( N_GND_c_398_p N_QN_c_9097_n ) capacitor c=0.0101988f //x=82.125 //y=0 \
 //x2=83.065 //y2=1.18
cc_473 ( N_GND_c_404_p N_QN_c_9097_n ) capacitor c=0.00469062f //x=84.19 //y=0 \
 //x2=83.065 //y2=1.18
cc_474 ( N_GND_c_2_p N_QN_c_9097_n ) capacitor c=0.00131455f //x=86.95 //y=0 \
 //x2=83.065 //y2=1.18
cc_475 ( N_GND_c_21_p N_QN_c_9097_n ) capacitor c=0.0412927f //x=81.03 //y=0 \
 //x2=83.065 //y2=1.18
cc_476 ( N_GND_M50_noxref_d N_QN_c_9097_n ) capacitor c=0.00960943f //x=82.02 \
 //y=0.865 //x2=83.065 //y2=1.18
cc_477 ( N_GND_c_23_p N_QN_c_9104_n ) capacitor c=0.00715563f //x=86.95 //y=0 \
 //x2=79.965 //y2=1.18
cc_478 ( N_GND_c_23_p N_QN_c_9105_n ) capacitor c=0.0769193f //x=86.95 //y=0 \
 //x2=86.395 //y2=1.18
cc_479 ( N_GND_c_404_p N_QN_c_9105_n ) capacitor c=0.00788597f //x=84.19 //y=0 \
 //x2=86.395 //y2=1.18
cc_480 ( N_GND_c_457_p N_QN_c_9105_n ) capacitor c=0.00974891f //x=85.455 \
 //y=0 //x2=86.395 //y2=1.18
cc_481 ( N_GND_c_2_p N_QN_c_9105_n ) capacitor c=0.00577463f //x=86.95 //y=0 \
 //x2=86.395 //y2=1.18
cc_482 ( N_GND_c_22_p N_QN_c_9105_n ) capacitor c=0.0384312f //x=84.36 //y=0 \
 //x2=86.395 //y2=1.18
cc_483 ( N_GND_M52_noxref_d N_QN_c_9105_n ) capacitor c=0.00960943f //x=85.35 \
 //y=0.865 //x2=86.395 //y2=1.18
cc_484 ( N_GND_c_23_p N_QN_c_9111_n ) capacitor c=0.00664346f //x=86.95 //y=0 \
 //x2=83.295 //y2=1.18
cc_485 ( N_GND_c_22_p QN ) capacitor c=0.00109945f //x=84.36 //y=0 //x2=86.95 \
 //y2=2.22
cc_486 ( N_GND_c_2_p N_QN_c_9113_n ) capacitor c=0.04686f //x=86.95 //y=0 \
 //x2=86.865 //y2=1.645
cc_487 ( N_GND_c_23_p N_QN_M49_noxref_d ) capacitor c=2.00936e-19 //x=86.95 \
 //y=0 //x2=79.66 //y2=0.905
cc_488 ( N_GND_c_21_p N_QN_M49_noxref_d ) capacitor c=0.00141366f //x=81.03 \
 //y=0 //x2=79.66 //y2=0.905
cc_489 ( N_GND_M48_noxref_d N_QN_M49_noxref_d ) capacitor c=0.00128667f \
 //x=78.69 //y=0.865 //x2=79.66 //y2=0.905
cc_490 ( N_GND_c_23_p N_QN_M51_noxref_d ) capacitor c=2.00936e-19 //x=86.95 \
 //y=0 //x2=82.99 //y2=0.905
cc_491 ( N_GND_c_22_p N_QN_M51_noxref_d ) capacitor c=0.0014176f //x=84.36 \
 //y=0 //x2=82.99 //y2=0.905
cc_492 ( N_GND_M50_noxref_d N_QN_M51_noxref_d ) capacitor c=0.0012247f \
 //x=82.02 //y=0.865 //x2=82.99 //y2=0.905
cc_493 ( N_GND_c_23_p N_QN_M53_noxref_d ) capacitor c=2.00936e-19 //x=86.95 \
 //y=0 //x2=86.32 //y2=0.905
cc_494 ( N_GND_c_2_p N_QN_M53_noxref_d ) capacitor c=0.00524992f //x=86.95 \
 //y=0 //x2=86.32 //y2=0.905
cc_495 ( N_GND_c_22_p N_QN_M53_noxref_d ) capacitor c=8.62423e-19 //x=84.36 \
 //y=0 //x2=86.32 //y2=0.905
cc_496 ( N_GND_M52_noxref_d N_QN_M53_noxref_d ) capacitor c=0.0012247f \
 //x=85.35 //y=0.865 //x2=86.32 //y2=0.905
cc_497 ( N_GND_c_23_p N_noxref_23_c_9266_n ) capacitor c=0.00618812f //x=86.95 \
 //y=0 //x2=1.475 //y2=1.59
cc_498 ( N_GND_c_95_p N_noxref_23_c_9266_n ) capacitor c=0.00110021f //x=0.99 \
 //y=0 //x2=1.475 //y2=1.59
cc_499 ( N_GND_c_24_p N_noxref_23_c_9266_n ) capacitor c=0.00179185f //x=4.64 \
 //y=0 //x2=1.475 //y2=1.59
cc_500 ( N_GND_M0_noxref_d N_noxref_23_c_9266_n ) capacitor c=0.00894788f \
 //x=0.885 //y=0.875 //x2=1.475 //y2=1.59
cc_501 ( N_GND_c_23_p N_noxref_23_c_9270_n ) capacitor c=0.00575184f //x=86.95 \
 //y=0 //x2=1.56 //y2=0.625
cc_502 ( N_GND_c_24_p N_noxref_23_c_9270_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=1.56 //y2=0.625
cc_503 ( N_GND_M0_noxref_d N_noxref_23_c_9270_n ) capacitor c=0.033954f \
 //x=0.885 //y=0.875 //x2=1.56 //y2=0.625
cc_504 ( N_GND_c_23_p N_noxref_23_c_9273_n ) capacitor c=0.0139021f //x=86.95 \
 //y=0 //x2=2.445 //y2=0.54
cc_505 ( N_GND_c_24_p N_noxref_23_c_9273_n ) capacitor c=0.0356078f //x=4.64 \
 //y=0 //x2=2.445 //y2=0.54
cc_506 ( N_GND_c_23_p N_noxref_23_M0_noxref_s ) capacitor c=0.0125336f \
 //x=86.95 //y=0 //x2=0.455 //y2=0.375
cc_507 ( N_GND_c_95_p N_noxref_23_M0_noxref_s ) capacitor c=0.0140218f \
 //x=0.99 //y=0 //x2=0.455 //y2=0.375
cc_508 ( N_GND_c_1_p N_noxref_23_M0_noxref_s ) capacitor c=0.0712607f //x=0.74 \
 //y=0 //x2=0.455 //y2=0.375
cc_509 ( N_GND_c_24_p N_noxref_23_M0_noxref_s ) capacitor c=0.0131422f \
 //x=4.64 //y=0 //x2=0.455 //y2=0.375
cc_510 ( N_GND_c_3_p N_noxref_23_M0_noxref_s ) capacitor c=3.31601e-19 \
 //x=4.81 //y=0 //x2=0.455 //y2=0.375
cc_511 ( N_GND_M0_noxref_d N_noxref_23_M0_noxref_s ) capacitor c=0.033718f \
 //x=0.885 //y=0.875 //x2=0.455 //y2=0.375
cc_512 ( N_GND_c_23_p N_noxref_24_c_9312_n ) capacitor c=0.00402784f //x=86.95 \
 //y=0 //x2=3.015 //y2=0.995
cc_513 ( N_GND_c_24_p N_noxref_24_c_9312_n ) capacitor c=0.00829979f //x=4.64 \
 //y=0 //x2=3.015 //y2=0.995
cc_514 ( N_GND_c_23_p N_noxref_24_c_9314_n ) capacitor c=0.00575184f //x=86.95 \
 //y=0 //x2=3.1 //y2=0.625
cc_515 ( N_GND_c_24_p N_noxref_24_c_9314_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=3.1 //y2=0.625
cc_516 ( N_GND_M0_noxref_d N_noxref_24_c_9314_n ) capacitor c=6.21394e-19 \
 //x=0.885 //y=0.875 //x2=3.1 //y2=0.625
cc_517 ( N_GND_c_23_p N_noxref_24_c_9317_n ) capacitor c=0.0118365f //x=86.95 \
 //y=0 //x2=3.985 //y2=0.54
cc_518 ( N_GND_c_24_p N_noxref_24_c_9317_n ) capacitor c=0.0365413f //x=4.64 \
 //y=0 //x2=3.985 //y2=0.54
cc_519 ( N_GND_c_23_p N_noxref_24_c_9319_n ) capacitor c=0.00287549f //x=86.95 \
 //y=0 //x2=4.07 //y2=0.625
cc_520 ( N_GND_c_24_p N_noxref_24_c_9319_n ) capacitor c=0.0142658f //x=4.64 \
 //y=0 //x2=4.07 //y2=0.625
cc_521 ( N_GND_c_3_p N_noxref_24_c_9319_n ) capacitor c=0.0404137f //x=4.81 \
 //y=0 //x2=4.07 //y2=0.625
cc_522 ( N_GND_M0_noxref_d N_noxref_24_M1_noxref_d ) capacitor c=0.00162435f \
 //x=0.885 //y=0.875 //x2=1.86 //y2=0.91
cc_523 ( N_GND_c_1_p N_noxref_24_M2_noxref_s ) capacitor c=8.16352e-19 \
 //x=0.74 //y=0 //x2=2.965 //y2=0.375
cc_524 ( N_GND_c_3_p N_noxref_24_M2_noxref_s ) capacitor c=0.00183204f \
 //x=4.81 //y=0 //x2=2.965 //y2=0.375
cc_525 ( N_GND_c_23_p N_noxref_25_c_9364_n ) capacitor c=0.00551063f //x=86.95 \
 //y=0 //x2=6.285 //y2=1.59
cc_526 ( N_GND_c_25_p N_noxref_25_c_9364_n ) capacitor c=0.00111576f //x=5.8 \
 //y=0 //x2=6.285 //y2=1.59
cc_527 ( N_GND_c_71_p N_noxref_25_c_9364_n ) capacitor c=0.0018074f //x=9.45 \
 //y=0 //x2=6.285 //y2=1.59
cc_528 ( N_GND_M3_noxref_d N_noxref_25_c_9364_n ) capacitor c=0.00887549f \
 //x=5.695 //y=0.875 //x2=6.285 //y2=1.59
cc_529 ( N_GND_c_23_p N_noxref_25_c_9368_n ) capacitor c=0.00287639f //x=86.95 \
 //y=0 //x2=6.37 //y2=0.625
cc_530 ( N_GND_c_71_p N_noxref_25_c_9368_n ) capacitor c=0.014327f //x=9.45 \
 //y=0 //x2=6.37 //y2=0.625
cc_531 ( N_GND_M3_noxref_d N_noxref_25_c_9368_n ) capacitor c=0.033954f \
 //x=5.695 //y=0.875 //x2=6.37 //y2=0.625
cc_532 ( N_GND_c_23_p N_noxref_25_c_9371_n ) capacitor c=0.0113713f //x=86.95 \
 //y=0 //x2=7.255 //y2=0.54
cc_533 ( N_GND_c_71_p N_noxref_25_c_9371_n ) capacitor c=0.0361671f //x=9.45 \
 //y=0 //x2=7.255 //y2=0.54
cc_534 ( N_GND_c_23_p N_noxref_25_M3_noxref_s ) capacitor c=0.00553362f \
 //x=86.95 //y=0 //x2=5.265 //y2=0.375
cc_535 ( N_GND_c_25_p N_noxref_25_M3_noxref_s ) capacitor c=0.014327f //x=5.8 \
 //y=0 //x2=5.265 //y2=0.375
cc_536 ( N_GND_c_71_p N_noxref_25_M3_noxref_s ) capacitor c=0.0137569f \
 //x=9.45 //y=0 //x2=5.265 //y2=0.375
cc_537 ( N_GND_c_3_p N_noxref_25_M3_noxref_s ) capacitor c=0.0696963f //x=4.81 \
 //y=0 //x2=5.265 //y2=0.375
cc_538 ( N_GND_c_4_p N_noxref_25_M3_noxref_s ) capacitor c=3.31601e-19 \
 //x=9.62 //y=0 //x2=5.265 //y2=0.375
cc_539 ( N_GND_M3_noxref_d N_noxref_25_M3_noxref_s ) capacitor c=0.033718f \
 //x=5.695 //y=0.875 //x2=5.265 //y2=0.375
cc_540 ( N_GND_c_23_p N_noxref_26_c_9416_n ) capacitor c=0.00364762f //x=86.95 \
 //y=0 //x2=7.825 //y2=0.995
cc_541 ( N_GND_c_71_p N_noxref_26_c_9416_n ) capacitor c=0.00940048f //x=9.45 \
 //y=0 //x2=7.825 //y2=0.995
cc_542 ( N_GND_c_23_p N_noxref_26_c_9418_n ) capacitor c=0.00266608f //x=86.95 \
 //y=0 //x2=7.91 //y2=0.625
cc_543 ( N_GND_c_71_p N_noxref_26_c_9418_n ) capacitor c=0.0141814f //x=9.45 \
 //y=0 //x2=7.91 //y2=0.625
cc_544 ( N_GND_M3_noxref_d N_noxref_26_c_9418_n ) capacitor c=6.21394e-19 \
 //x=5.695 //y=0.875 //x2=7.91 //y2=0.625
cc_545 ( N_GND_c_23_p N_noxref_26_c_9421_n ) capacitor c=0.0105197f //x=86.95 \
 //y=0 //x2=8.795 //y2=0.54
cc_546 ( N_GND_c_71_p N_noxref_26_c_9421_n ) capacitor c=0.036368f //x=9.45 \
 //y=0 //x2=8.795 //y2=0.54
cc_547 ( N_GND_c_23_p N_noxref_26_c_9423_n ) capacitor c=0.00254232f //x=86.95 \
 //y=0 //x2=8.88 //y2=0.625
cc_548 ( N_GND_c_71_p N_noxref_26_c_9423_n ) capacitor c=0.0140304f //x=9.45 \
 //y=0 //x2=8.88 //y2=0.625
cc_549 ( N_GND_c_4_p N_noxref_26_c_9423_n ) capacitor c=0.0404137f //x=9.62 \
 //y=0 //x2=8.88 //y2=0.625
cc_550 ( N_GND_M3_noxref_d N_noxref_26_M4_noxref_d ) capacitor c=0.00162435f \
 //x=5.695 //y=0.875 //x2=6.67 //y2=0.91
cc_551 ( N_GND_c_3_p N_noxref_26_M5_noxref_s ) capacitor c=8.16352e-19 \
 //x=4.81 //y=0 //x2=7.775 //y2=0.375
cc_552 ( N_GND_c_4_p N_noxref_26_M5_noxref_s ) capacitor c=0.00183576f \
 //x=9.62 //y=0 //x2=7.775 //y2=0.375
cc_553 ( N_GND_c_23_p N_noxref_27_c_9469_n ) capacitor c=0.00517234f //x=86.95 \
 //y=0 //x2=11.2 //y2=1.58
cc_554 ( N_GND_c_32_p N_noxref_27_c_9469_n ) capacitor c=0.00112872f \
 //x=10.715 //y=0 //x2=11.2 //y2=1.58
cc_555 ( N_GND_c_39_p N_noxref_27_c_9469_n ) capacitor c=0.0018229f //x=12.78 \
 //y=0 //x2=11.2 //y2=1.58
cc_556 ( N_GND_M6_noxref_d N_noxref_27_c_9469_n ) capacitor c=0.008625f \
 //x=10.61 //y=0.865 //x2=11.2 //y2=1.58
cc_557 ( N_GND_c_23_p N_noxref_27_c_9473_n ) capacitor c=0.00259029f //x=86.95 \
 //y=0 //x2=11.285 //y2=0.615
cc_558 ( N_GND_c_39_p N_noxref_27_c_9473_n ) capacitor c=0.0146901f //x=12.78 \
 //y=0 //x2=11.285 //y2=0.615
cc_559 ( N_GND_M6_noxref_d N_noxref_27_c_9473_n ) capacitor c=0.033812f \
 //x=10.61 //y=0.865 //x2=11.285 //y2=0.615
cc_560 ( N_GND_c_4_p N_noxref_27_c_9476_n ) capacitor c=2.91423e-19 //x=9.62 \
 //y=0 //x2=11.285 //y2=1.495
cc_561 ( N_GND_c_23_p N_noxref_27_c_9477_n ) capacitor c=0.0106919f //x=86.95 \
 //y=0 //x2=12.17 //y2=0.53
cc_562 ( N_GND_c_39_p N_noxref_27_c_9477_n ) capacitor c=0.0374253f //x=12.78 \
 //y=0 //x2=12.17 //y2=0.53
cc_563 ( N_GND_c_23_p N_noxref_27_c_9479_n ) capacitor c=0.00258845f //x=86.95 \
 //y=0 //x2=12.255 //y2=0.615
cc_564 ( N_GND_c_39_p N_noxref_27_c_9479_n ) capacitor c=0.0146256f //x=12.78 \
 //y=0 //x2=12.255 //y2=0.615
cc_565 ( N_GND_c_5_p N_noxref_27_c_9479_n ) capacitor c=0.0431718f //x=12.95 \
 //y=0 //x2=12.255 //y2=0.615
cc_566 ( N_GND_c_23_p N_noxref_27_M6_noxref_s ) capacitor c=0.00259029f \
 //x=86.95 //y=0 //x2=10.18 //y2=0.365
cc_567 ( N_GND_c_32_p N_noxref_27_M6_noxref_s ) capacitor c=0.0146901f \
 //x=10.715 //y=0 //x2=10.18 //y2=0.365
cc_568 ( N_GND_c_4_p N_noxref_27_M6_noxref_s ) capacitor c=0.0583534f //x=9.62 \
 //y=0 //x2=10.18 //y2=0.365
cc_569 ( N_GND_c_5_p N_noxref_27_M6_noxref_s ) capacitor c=0.00198098f \
 //x=12.95 //y=0 //x2=10.18 //y2=0.365
cc_570 ( N_GND_M6_noxref_d N_noxref_27_M6_noxref_s ) capacitor c=0.0334197f \
 //x=10.61 //y=0.865 //x2=10.18 //y2=0.365
cc_571 ( N_GND_c_23_p N_noxref_28_c_9520_n ) capacitor c=0.00517576f //x=86.95 \
 //y=0 //x2=14.425 //y2=1.59
cc_572 ( N_GND_c_47_p N_noxref_28_c_9520_n ) capacitor c=0.00111448f //x=13.94 \
 //y=0 //x2=14.425 //y2=1.59
cc_573 ( N_GND_c_54_p N_noxref_28_c_9520_n ) capacitor c=0.00180612f //x=17.59 \
 //y=0 //x2=14.425 //y2=1.59
cc_574 ( N_GND_M8_noxref_d N_noxref_28_c_9520_n ) capacitor c=0.00853078f \
 //x=13.835 //y=0.875 //x2=14.425 //y2=1.59
cc_575 ( N_GND_c_23_p N_noxref_28_c_9524_n ) capacitor c=0.00254475f //x=86.95 \
 //y=0 //x2=14.51 //y2=0.625
cc_576 ( N_GND_c_54_p N_noxref_28_c_9524_n ) capacitor c=0.0140928f //x=17.59 \
 //y=0 //x2=14.51 //y2=0.625
cc_577 ( N_GND_M8_noxref_d N_noxref_28_c_9524_n ) capacitor c=0.033954f \
 //x=13.835 //y=0.875 //x2=14.51 //y2=0.625
cc_578 ( N_GND_c_23_p N_noxref_28_c_9527_n ) capacitor c=0.0104506f //x=86.95 \
 //y=0 //x2=15.395 //y2=0.54
cc_579 ( N_GND_c_54_p N_noxref_28_c_9527_n ) capacitor c=0.0360726f //x=17.59 \
 //y=0 //x2=15.395 //y2=0.54
cc_580 ( N_GND_c_23_p N_noxref_28_M8_noxref_s ) capacitor c=0.00507657f \
 //x=86.95 //y=0 //x2=13.405 //y2=0.375
cc_581 ( N_GND_c_47_p N_noxref_28_M8_noxref_s ) capacitor c=0.0140928f \
 //x=13.94 //y=0 //x2=13.405 //y2=0.375
cc_582 ( N_GND_c_54_p N_noxref_28_M8_noxref_s ) capacitor c=0.0136651f \
 //x=17.59 //y=0 //x2=13.405 //y2=0.375
cc_583 ( N_GND_c_5_p N_noxref_28_M8_noxref_s ) capacitor c=0.0696963f \
 //x=12.95 //y=0 //x2=13.405 //y2=0.375
cc_584 ( N_GND_c_6_p N_noxref_28_M8_noxref_s ) capacitor c=3.31601e-19 \
 //x=17.76 //y=0 //x2=13.405 //y2=0.375
cc_585 ( N_GND_M8_noxref_d N_noxref_28_M8_noxref_s ) capacitor c=0.033718f \
 //x=13.835 //y=0.875 //x2=13.405 //y2=0.375
cc_586 ( N_GND_c_23_p N_noxref_29_c_9569_n ) capacitor c=0.00352952f //x=86.95 \
 //y=0 //x2=15.965 //y2=0.995
cc_587 ( N_GND_c_54_p N_noxref_29_c_9569_n ) capacitor c=0.00934524f //x=17.59 \
 //y=0 //x2=15.965 //y2=0.995
cc_588 ( N_GND_c_23_p N_noxref_29_c_9571_n ) capacitor c=0.00254475f //x=86.95 \
 //y=0 //x2=16.05 //y2=0.625
cc_589 ( N_GND_c_54_p N_noxref_29_c_9571_n ) capacitor c=0.0140928f //x=17.59 \
 //y=0 //x2=16.05 //y2=0.625
cc_590 ( N_GND_M8_noxref_d N_noxref_29_c_9571_n ) capacitor c=6.21394e-19 \
 //x=13.835 //y=0.875 //x2=16.05 //y2=0.625
cc_591 ( N_GND_c_23_p N_noxref_29_c_9574_n ) capacitor c=0.0105197f //x=86.95 \
 //y=0 //x2=16.935 //y2=0.54
cc_592 ( N_GND_c_54_p N_noxref_29_c_9574_n ) capacitor c=0.0364139f //x=17.59 \
 //y=0 //x2=16.935 //y2=0.54
cc_593 ( N_GND_c_23_p N_noxref_29_c_9576_n ) capacitor c=0.00254232f //x=86.95 \
 //y=0 //x2=17.02 //y2=0.625
cc_594 ( N_GND_c_54_p N_noxref_29_c_9576_n ) capacitor c=0.0140304f //x=17.59 \
 //y=0 //x2=17.02 //y2=0.625
cc_595 ( N_GND_c_6_p N_noxref_29_c_9576_n ) capacitor c=0.0404137f //x=17.76 \
 //y=0 //x2=17.02 //y2=0.625
cc_596 ( N_GND_M8_noxref_d N_noxref_29_M9_noxref_d ) capacitor c=0.00162435f \
 //x=13.835 //y=0.875 //x2=14.81 //y2=0.91
cc_597 ( N_GND_c_5_p N_noxref_29_M10_noxref_s ) capacitor c=8.16352e-19 \
 //x=12.95 //y=0 //x2=15.915 //y2=0.375
cc_598 ( N_GND_c_6_p N_noxref_29_M10_noxref_s ) capacitor c=0.00183204f \
 //x=17.76 //y=0 //x2=15.915 //y2=0.375
cc_599 ( N_GND_c_23_p N_noxref_30_c_9622_n ) capacitor c=0.00517576f //x=86.95 \
 //y=0 //x2=19.235 //y2=1.59
cc_600 ( N_GND_c_74_p N_noxref_30_c_9622_n ) capacitor c=0.00111448f //x=18.75 \
 //y=0 //x2=19.235 //y2=1.59
cc_601 ( N_GND_c_81_p N_noxref_30_c_9622_n ) capacitor c=0.00180612f //x=22.4 \
 //y=0 //x2=19.235 //y2=1.59
cc_602 ( N_GND_M11_noxref_d N_noxref_30_c_9622_n ) capacitor c=0.00853078f \
 //x=18.645 //y=0.875 //x2=19.235 //y2=1.59
cc_603 ( N_GND_c_23_p N_noxref_30_c_9626_n ) capacitor c=0.00254475f //x=86.95 \
 //y=0 //x2=19.32 //y2=0.625
cc_604 ( N_GND_c_81_p N_noxref_30_c_9626_n ) capacitor c=0.0140928f //x=22.4 \
 //y=0 //x2=19.32 //y2=0.625
cc_605 ( N_GND_M11_noxref_d N_noxref_30_c_9626_n ) capacitor c=0.033954f \
 //x=18.645 //y=0.875 //x2=19.32 //y2=0.625
cc_606 ( N_GND_c_23_p N_noxref_30_c_9629_n ) capacitor c=0.0104386f //x=86.95 \
 //y=0 //x2=20.205 //y2=0.54
cc_607 ( N_GND_c_81_p N_noxref_30_c_9629_n ) capacitor c=0.0360726f //x=22.4 \
 //y=0 //x2=20.205 //y2=0.54
cc_608 ( N_GND_c_23_p N_noxref_30_M11_noxref_s ) capacitor c=0.00507657f \
 //x=86.95 //y=0 //x2=18.215 //y2=0.375
cc_609 ( N_GND_c_74_p N_noxref_30_M11_noxref_s ) capacitor c=0.0140928f \
 //x=18.75 //y=0 //x2=18.215 //y2=0.375
cc_610 ( N_GND_c_81_p N_noxref_30_M11_noxref_s ) capacitor c=0.0131437f \
 //x=22.4 //y=0 //x2=18.215 //y2=0.375
cc_611 ( N_GND_c_6_p N_noxref_30_M11_noxref_s ) capacitor c=0.0696963f \
 //x=17.76 //y=0 //x2=18.215 //y2=0.375
cc_612 ( N_GND_c_7_p N_noxref_30_M11_noxref_s ) capacitor c=3.31601e-19 \
 //x=22.57 //y=0 //x2=18.215 //y2=0.375
cc_613 ( N_GND_M11_noxref_d N_noxref_30_M11_noxref_s ) capacitor c=0.033718f \
 //x=18.645 //y=0.875 //x2=18.215 //y2=0.375
cc_614 ( N_GND_c_23_p N_noxref_31_c_9674_n ) capacitor c=0.00352952f //x=86.95 \
 //y=0 //x2=20.775 //y2=0.995
cc_615 ( N_GND_c_81_p N_noxref_31_c_9674_n ) capacitor c=0.00934524f //x=22.4 \
 //y=0 //x2=20.775 //y2=0.995
cc_616 ( N_GND_c_23_p N_noxref_31_c_9676_n ) capacitor c=0.00254475f //x=86.95 \
 //y=0 //x2=20.86 //y2=0.625
cc_617 ( N_GND_c_81_p N_noxref_31_c_9676_n ) capacitor c=0.0140928f //x=22.4 \
 //y=0 //x2=20.86 //y2=0.625
cc_618 ( N_GND_M11_noxref_d N_noxref_31_c_9676_n ) capacitor c=6.21394e-19 \
 //x=18.645 //y=0.875 //x2=20.86 //y2=0.625
cc_619 ( N_GND_c_23_p N_noxref_31_c_9679_n ) capacitor c=0.0105317f //x=86.95 \
 //y=0 //x2=21.745 //y2=0.54
cc_620 ( N_GND_c_81_p N_noxref_31_c_9679_n ) capacitor c=0.036415f //x=22.4 \
 //y=0 //x2=21.745 //y2=0.54
cc_621 ( N_GND_c_23_p N_noxref_31_c_9681_n ) capacitor c=0.00254232f //x=86.95 \
 //y=0 //x2=21.83 //y2=0.625
cc_622 ( N_GND_c_81_p N_noxref_31_c_9681_n ) capacitor c=0.0140304f //x=22.4 \
 //y=0 //x2=21.83 //y2=0.625
cc_623 ( N_GND_c_7_p N_noxref_31_c_9681_n ) capacitor c=0.0404137f //x=22.57 \
 //y=0 //x2=21.83 //y2=0.625
cc_624 ( N_GND_M11_noxref_d N_noxref_31_M12_noxref_d ) capacitor c=0.00162435f \
 //x=18.645 //y=0.875 //x2=19.62 //y2=0.91
cc_625 ( N_GND_c_6_p N_noxref_31_M13_noxref_s ) capacitor c=8.16352e-19 \
 //x=17.76 //y=0 //x2=20.725 //y2=0.375
cc_626 ( N_GND_c_7_p N_noxref_31_M13_noxref_s ) capacitor c=0.00183576f \
 //x=22.57 //y=0 //x2=20.725 //y2=0.375
cc_627 ( N_GND_c_23_p N_noxref_32_c_9726_n ) capacitor c=0.00517234f //x=86.95 \
 //y=0 //x2=24.15 //y2=1.58
cc_628 ( N_GND_c_105_p N_noxref_32_c_9726_n ) capacitor c=0.00112872f \
 //x=23.665 //y=0 //x2=24.15 //y2=1.58
cc_629 ( N_GND_c_112_p N_noxref_32_c_9726_n ) capacitor c=0.0018229f //x=25.73 \
 //y=0 //x2=24.15 //y2=1.58
cc_630 ( N_GND_M14_noxref_d N_noxref_32_c_9726_n ) capacitor c=0.008625f \
 //x=23.56 //y=0.865 //x2=24.15 //y2=1.58
cc_631 ( N_GND_c_23_p N_noxref_32_c_9730_n ) capacitor c=0.00259029f //x=86.95 \
 //y=0 //x2=24.235 //y2=0.615
cc_632 ( N_GND_c_112_p N_noxref_32_c_9730_n ) capacitor c=0.0146901f //x=25.73 \
 //y=0 //x2=24.235 //y2=0.615
cc_633 ( N_GND_M14_noxref_d N_noxref_32_c_9730_n ) capacitor c=0.033812f \
 //x=23.56 //y=0.865 //x2=24.235 //y2=0.615
cc_634 ( N_GND_c_7_p N_noxref_32_c_9733_n ) capacitor c=2.91423e-19 //x=22.57 \
 //y=0 //x2=24.235 //y2=1.495
cc_635 ( N_GND_c_23_p N_noxref_32_c_9734_n ) capacitor c=0.0106919f //x=86.95 \
 //y=0 //x2=25.12 //y2=0.53
cc_636 ( N_GND_c_112_p N_noxref_32_c_9734_n ) capacitor c=0.0374253f //x=25.73 \
 //y=0 //x2=25.12 //y2=0.53
cc_637 ( N_GND_c_23_p N_noxref_32_c_9736_n ) capacitor c=0.00258845f //x=86.95 \
 //y=0 //x2=25.205 //y2=0.615
cc_638 ( N_GND_c_112_p N_noxref_32_c_9736_n ) capacitor c=0.0146256f //x=25.73 \
 //y=0 //x2=25.205 //y2=0.615
cc_639 ( N_GND_c_8_p N_noxref_32_c_9736_n ) capacitor c=0.0431718f //x=25.9 \
 //y=0 //x2=25.205 //y2=0.615
cc_640 ( N_GND_c_23_p N_noxref_32_M14_noxref_s ) capacitor c=0.00259029f \
 //x=86.95 //y=0 //x2=23.13 //y2=0.365
cc_641 ( N_GND_c_105_p N_noxref_32_M14_noxref_s ) capacitor c=0.0146901f \
 //x=23.665 //y=0 //x2=23.13 //y2=0.365
cc_642 ( N_GND_c_7_p N_noxref_32_M14_noxref_s ) capacitor c=0.0583534f \
 //x=22.57 //y=0 //x2=23.13 //y2=0.365
cc_643 ( N_GND_c_8_p N_noxref_32_M14_noxref_s ) capacitor c=0.00198098f \
 //x=25.9 //y=0 //x2=23.13 //y2=0.365
cc_644 ( N_GND_M14_noxref_d N_noxref_32_M14_noxref_s ) capacitor c=0.0334197f \
 //x=23.56 //y=0.865 //x2=23.13 //y2=0.365
cc_645 ( N_GND_c_23_p N_noxref_33_c_9777_n ) capacitor c=0.00517576f //x=86.95 \
 //y=0 //x2=27.375 //y2=1.59
cc_646 ( N_GND_c_190_p N_noxref_33_c_9777_n ) capacitor c=0.00111448f \
 //x=26.89 //y=0 //x2=27.375 //y2=1.59
cc_647 ( N_GND_c_197_p N_noxref_33_c_9777_n ) capacitor c=0.00180612f \
 //x=30.54 //y=0 //x2=27.375 //y2=1.59
cc_648 ( N_GND_M16_noxref_d N_noxref_33_c_9777_n ) capacitor c=0.00853078f \
 //x=26.785 //y=0.875 //x2=27.375 //y2=1.59
cc_649 ( N_GND_c_23_p N_noxref_33_c_9781_n ) capacitor c=0.00254475f //x=86.95 \
 //y=0 //x2=27.46 //y2=0.625
cc_650 ( N_GND_c_197_p N_noxref_33_c_9781_n ) capacitor c=0.0140928f //x=30.54 \
 //y=0 //x2=27.46 //y2=0.625
cc_651 ( N_GND_M16_noxref_d N_noxref_33_c_9781_n ) capacitor c=0.033954f \
 //x=26.785 //y=0.875 //x2=27.46 //y2=0.625
cc_652 ( N_GND_c_23_p N_noxref_33_c_9784_n ) capacitor c=0.0104506f //x=86.95 \
 //y=0 //x2=28.345 //y2=0.54
cc_653 ( N_GND_c_197_p N_noxref_33_c_9784_n ) capacitor c=0.0360726f //x=30.54 \
 //y=0 //x2=28.345 //y2=0.54
cc_654 ( N_GND_c_23_p N_noxref_33_M16_noxref_s ) capacitor c=0.00507657f \
 //x=86.95 //y=0 //x2=26.355 //y2=0.375
cc_655 ( N_GND_c_190_p N_noxref_33_M16_noxref_s ) capacitor c=0.0140928f \
 //x=26.89 //y=0 //x2=26.355 //y2=0.375
cc_656 ( N_GND_c_197_p N_noxref_33_M16_noxref_s ) capacitor c=0.0136651f \
 //x=30.54 //y=0 //x2=26.355 //y2=0.375
cc_657 ( N_GND_c_8_p N_noxref_33_M16_noxref_s ) capacitor c=0.0696963f \
 //x=25.9 //y=0 //x2=26.355 //y2=0.375
cc_658 ( N_GND_c_9_p N_noxref_33_M16_noxref_s ) capacitor c=3.31601e-19 \
 //x=30.71 //y=0 //x2=26.355 //y2=0.375
cc_659 ( N_GND_M16_noxref_d N_noxref_33_M16_noxref_s ) capacitor c=0.033718f \
 //x=26.785 //y=0.875 //x2=26.355 //y2=0.375
cc_660 ( N_GND_c_23_p N_noxref_34_c_9826_n ) capacitor c=0.00352952f //x=86.95 \
 //y=0 //x2=28.915 //y2=0.995
cc_661 ( N_GND_c_197_p N_noxref_34_c_9826_n ) capacitor c=0.00934524f \
 //x=30.54 //y=0 //x2=28.915 //y2=0.995
cc_662 ( N_GND_c_23_p N_noxref_34_c_9828_n ) capacitor c=0.00254475f //x=86.95 \
 //y=0 //x2=29 //y2=0.625
cc_663 ( N_GND_c_197_p N_noxref_34_c_9828_n ) capacitor c=0.0140928f //x=30.54 \
 //y=0 //x2=29 //y2=0.625
cc_664 ( N_GND_M16_noxref_d N_noxref_34_c_9828_n ) capacitor c=6.21394e-19 \
 //x=26.785 //y=0.875 //x2=29 //y2=0.625
cc_665 ( N_GND_c_23_p N_noxref_34_c_9831_n ) capacitor c=0.0105317f //x=86.95 \
 //y=0 //x2=29.885 //y2=0.54
cc_666 ( N_GND_c_197_p N_noxref_34_c_9831_n ) capacitor c=0.036415f //x=30.54 \
 //y=0 //x2=29.885 //y2=0.54
cc_667 ( N_GND_c_23_p N_noxref_34_c_9833_n ) capacitor c=0.00254232f //x=86.95 \
 //y=0 //x2=29.97 //y2=0.625
cc_668 ( N_GND_c_197_p N_noxref_34_c_9833_n ) capacitor c=0.0140304f //x=30.54 \
 //y=0 //x2=29.97 //y2=0.625
cc_669 ( N_GND_c_9_p N_noxref_34_c_9833_n ) capacitor c=0.0404137f //x=30.71 \
 //y=0 //x2=29.97 //y2=0.625
cc_670 ( N_GND_M16_noxref_d N_noxref_34_M17_noxref_d ) capacitor c=0.00162435f \
 //x=26.785 //y=0.875 //x2=27.76 //y2=0.91
cc_671 ( N_GND_c_8_p N_noxref_34_M18_noxref_s ) capacitor c=8.16352e-19 \
 //x=25.9 //y=0 //x2=28.865 //y2=0.375
cc_672 ( N_GND_c_9_p N_noxref_34_M18_noxref_s ) capacitor c=0.00183204f \
 //x=30.71 //y=0 //x2=28.865 //y2=0.375
cc_673 ( N_GND_c_23_p N_noxref_35_c_9878_n ) capacitor c=0.00517576f //x=86.95 \
 //y=0 //x2=32.185 //y2=1.59
cc_674 ( N_GND_c_150_p N_noxref_35_c_9878_n ) capacitor c=0.00111448f //x=31.7 \
 //y=0 //x2=32.185 //y2=1.59
cc_675 ( N_GND_c_157_p N_noxref_35_c_9878_n ) capacitor c=0.00180612f \
 //x=35.35 //y=0 //x2=32.185 //y2=1.59
cc_676 ( N_GND_M19_noxref_d N_noxref_35_c_9878_n ) capacitor c=0.00853078f \
 //x=31.595 //y=0.875 //x2=32.185 //y2=1.59
cc_677 ( N_GND_c_23_p N_noxref_35_c_9882_n ) capacitor c=0.00254475f //x=86.95 \
 //y=0 //x2=32.27 //y2=0.625
cc_678 ( N_GND_c_157_p N_noxref_35_c_9882_n ) capacitor c=0.0140928f //x=35.35 \
 //y=0 //x2=32.27 //y2=0.625
cc_679 ( N_GND_M19_noxref_d N_noxref_35_c_9882_n ) capacitor c=0.033954f \
 //x=31.595 //y=0.875 //x2=32.27 //y2=0.625
cc_680 ( N_GND_c_23_p N_noxref_35_c_9885_n ) capacitor c=0.0104506f //x=86.95 \
 //y=0 //x2=33.155 //y2=0.54
cc_681 ( N_GND_c_157_p N_noxref_35_c_9885_n ) capacitor c=0.0360726f //x=35.35 \
 //y=0 //x2=33.155 //y2=0.54
cc_682 ( N_GND_c_23_p N_noxref_35_M19_noxref_s ) capacitor c=0.00507657f \
 //x=86.95 //y=0 //x2=31.165 //y2=0.375
cc_683 ( N_GND_c_150_p N_noxref_35_M19_noxref_s ) capacitor c=0.0140928f \
 //x=31.7 //y=0 //x2=31.165 //y2=0.375
cc_684 ( N_GND_c_157_p N_noxref_35_M19_noxref_s ) capacitor c=0.0136651f \
 //x=35.35 //y=0 //x2=31.165 //y2=0.375
cc_685 ( N_GND_c_9_p N_noxref_35_M19_noxref_s ) capacitor c=0.0696963f \
 //x=30.71 //y=0 //x2=31.165 //y2=0.375
cc_686 ( N_GND_c_10_p N_noxref_35_M19_noxref_s ) capacitor c=3.31601e-19 \
 //x=35.52 //y=0 //x2=31.165 //y2=0.375
cc_687 ( N_GND_M19_noxref_d N_noxref_35_M19_noxref_s ) capacitor c=0.033718f \
 //x=31.595 //y=0.875 //x2=31.165 //y2=0.375
cc_688 ( N_GND_c_23_p N_noxref_36_c_9927_n ) capacitor c=0.00352952f //x=86.95 \
 //y=0 //x2=33.725 //y2=0.995
cc_689 ( N_GND_c_157_p N_noxref_36_c_9927_n ) capacitor c=0.00934524f \
 //x=35.35 //y=0 //x2=33.725 //y2=0.995
cc_690 ( N_GND_c_23_p N_noxref_36_c_9929_n ) capacitor c=0.00254475f //x=86.95 \
 //y=0 //x2=33.81 //y2=0.625
cc_691 ( N_GND_c_157_p N_noxref_36_c_9929_n ) capacitor c=0.0140928f //x=35.35 \
 //y=0 //x2=33.81 //y2=0.625
cc_692 ( N_GND_M19_noxref_d N_noxref_36_c_9929_n ) capacitor c=6.21394e-19 \
 //x=31.595 //y=0.875 //x2=33.81 //y2=0.625
cc_693 ( N_GND_c_23_p N_noxref_36_c_9932_n ) capacitor c=0.0105197f //x=86.95 \
 //y=0 //x2=34.695 //y2=0.54
cc_694 ( N_GND_c_157_p N_noxref_36_c_9932_n ) capacitor c=0.036368f //x=35.35 \
 //y=0 //x2=34.695 //y2=0.54
cc_695 ( N_GND_c_23_p N_noxref_36_c_9934_n ) capacitor c=0.00254232f //x=86.95 \
 //y=0 //x2=34.78 //y2=0.625
cc_696 ( N_GND_c_157_p N_noxref_36_c_9934_n ) capacitor c=0.0140304f //x=35.35 \
 //y=0 //x2=34.78 //y2=0.625
cc_697 ( N_GND_c_10_p N_noxref_36_c_9934_n ) capacitor c=0.0404137f //x=35.52 \
 //y=0 //x2=34.78 //y2=0.625
cc_698 ( N_GND_M19_noxref_d N_noxref_36_M20_noxref_d ) capacitor c=0.00162435f \
 //x=31.595 //y=0.875 //x2=32.57 //y2=0.91
cc_699 ( N_GND_c_9_p N_noxref_36_M21_noxref_s ) capacitor c=8.16352e-19 \
 //x=30.71 //y=0 //x2=33.675 //y2=0.375
cc_700 ( N_GND_c_10_p N_noxref_36_M21_noxref_s ) capacitor c=0.00183576f \
 //x=35.52 //y=0 //x2=33.675 //y2=0.375
cc_701 ( N_GND_c_23_p N_noxref_37_c_9980_n ) capacitor c=0.00517234f //x=86.95 \
 //y=0 //x2=37.1 //y2=1.58
cc_702 ( N_GND_c_120_p N_noxref_37_c_9980_n ) capacitor c=0.00112872f \
 //x=36.615 //y=0 //x2=37.1 //y2=1.58
cc_703 ( N_GND_c_127_p N_noxref_37_c_9980_n ) capacitor c=0.0018229f //x=38.68 \
 //y=0 //x2=37.1 //y2=1.58
cc_704 ( N_GND_M22_noxref_d N_noxref_37_c_9980_n ) capacitor c=0.008625f \
 //x=36.51 //y=0.865 //x2=37.1 //y2=1.58
cc_705 ( N_GND_c_23_p N_noxref_37_c_9984_n ) capacitor c=0.00259029f //x=86.95 \
 //y=0 //x2=37.185 //y2=0.615
cc_706 ( N_GND_c_127_p N_noxref_37_c_9984_n ) capacitor c=0.0146901f //x=38.68 \
 //y=0 //x2=37.185 //y2=0.615
cc_707 ( N_GND_M22_noxref_d N_noxref_37_c_9984_n ) capacitor c=0.033812f \
 //x=36.51 //y=0.865 //x2=37.185 //y2=0.615
cc_708 ( N_GND_c_10_p N_noxref_37_c_9987_n ) capacitor c=2.91423e-19 //x=35.52 \
 //y=0 //x2=37.185 //y2=1.495
cc_709 ( N_GND_c_23_p N_noxref_37_c_9988_n ) capacitor c=0.0106919f //x=86.95 \
 //y=0 //x2=38.07 //y2=0.53
cc_710 ( N_GND_c_127_p N_noxref_37_c_9988_n ) capacitor c=0.0374253f //x=38.68 \
 //y=0 //x2=38.07 //y2=0.53
cc_711 ( N_GND_c_23_p N_noxref_37_c_9990_n ) capacitor c=0.00258845f //x=86.95 \
 //y=0 //x2=38.155 //y2=0.615
cc_712 ( N_GND_c_127_p N_noxref_37_c_9990_n ) capacitor c=0.0146256f //x=38.68 \
 //y=0 //x2=38.155 //y2=0.615
cc_713 ( N_GND_c_11_p N_noxref_37_c_9990_n ) capacitor c=0.0431718f //x=38.85 \
 //y=0 //x2=38.155 //y2=0.615
cc_714 ( N_GND_c_23_p N_noxref_37_M22_noxref_s ) capacitor c=0.00259029f \
 //x=86.95 //y=0 //x2=36.08 //y2=0.365
cc_715 ( N_GND_c_120_p N_noxref_37_M22_noxref_s ) capacitor c=0.0146901f \
 //x=36.615 //y=0 //x2=36.08 //y2=0.365
cc_716 ( N_GND_c_10_p N_noxref_37_M22_noxref_s ) capacitor c=0.0583534f \
 //x=35.52 //y=0 //x2=36.08 //y2=0.365
cc_717 ( N_GND_c_11_p N_noxref_37_M22_noxref_s ) capacitor c=0.00198098f \
 //x=38.85 //y=0 //x2=36.08 //y2=0.365
cc_718 ( N_GND_M22_noxref_d N_noxref_37_M22_noxref_s ) capacitor c=0.0334197f \
 //x=36.51 //y=0.865 //x2=36.08 //y2=0.365
cc_719 ( N_GND_c_23_p N_noxref_38_c_10031_n ) capacitor c=0.00517576f \
 //x=86.95 //y=0 //x2=40.325 //y2=1.59
cc_720 ( N_GND_c_134_p N_noxref_38_c_10031_n ) capacitor c=0.00111448f \
 //x=39.84 //y=0 //x2=40.325 //y2=1.59
cc_721 ( N_GND_c_141_p N_noxref_38_c_10031_n ) capacitor c=0.00180612f \
 //x=43.49 //y=0 //x2=40.325 //y2=1.59
cc_722 ( N_GND_M24_noxref_d N_noxref_38_c_10031_n ) capacitor c=0.00853078f \
 //x=39.735 //y=0.875 //x2=40.325 //y2=1.59
cc_723 ( N_GND_c_23_p N_noxref_38_c_10035_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=40.41 //y2=0.625
cc_724 ( N_GND_c_141_p N_noxref_38_c_10035_n ) capacitor c=0.0140928f \
 //x=43.49 //y=0 //x2=40.41 //y2=0.625
cc_725 ( N_GND_M24_noxref_d N_noxref_38_c_10035_n ) capacitor c=0.033954f \
 //x=39.735 //y=0.875 //x2=40.41 //y2=0.625
cc_726 ( N_GND_c_23_p N_noxref_38_c_10038_n ) capacitor c=0.0104506f //x=86.95 \
 //y=0 //x2=41.295 //y2=0.54
cc_727 ( N_GND_c_141_p N_noxref_38_c_10038_n ) capacitor c=0.0360726f \
 //x=43.49 //y=0 //x2=41.295 //y2=0.54
cc_728 ( N_GND_c_23_p N_noxref_38_M24_noxref_s ) capacitor c=0.00507657f \
 //x=86.95 //y=0 //x2=39.305 //y2=0.375
cc_729 ( N_GND_c_134_p N_noxref_38_M24_noxref_s ) capacitor c=0.0140928f \
 //x=39.84 //y=0 //x2=39.305 //y2=0.375
cc_730 ( N_GND_c_141_p N_noxref_38_M24_noxref_s ) capacitor c=0.0131437f \
 //x=43.49 //y=0 //x2=39.305 //y2=0.375
cc_731 ( N_GND_c_11_p N_noxref_38_M24_noxref_s ) capacitor c=0.0696963f \
 //x=38.85 //y=0 //x2=39.305 //y2=0.375
cc_732 ( N_GND_c_12_p N_noxref_38_M24_noxref_s ) capacitor c=3.31601e-19 \
 //x=43.66 //y=0 //x2=39.305 //y2=0.375
cc_733 ( N_GND_M24_noxref_d N_noxref_38_M24_noxref_s ) capacitor c=0.033718f \
 //x=39.735 //y=0.875 //x2=39.305 //y2=0.375
cc_734 ( N_GND_c_23_p N_noxref_39_c_10080_n ) capacitor c=0.00352952f \
 //x=86.95 //y=0 //x2=41.865 //y2=0.995
cc_735 ( N_GND_c_141_p N_noxref_39_c_10080_n ) capacitor c=0.00934524f \
 //x=43.49 //y=0 //x2=41.865 //y2=0.995
cc_736 ( N_GND_c_23_p N_noxref_39_c_10082_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=41.95 //y2=0.625
cc_737 ( N_GND_c_141_p N_noxref_39_c_10082_n ) capacitor c=0.0140928f \
 //x=43.49 //y=0 //x2=41.95 //y2=0.625
cc_738 ( N_GND_M24_noxref_d N_noxref_39_c_10082_n ) capacitor c=6.21394e-19 \
 //x=39.735 //y=0.875 //x2=41.95 //y2=0.625
cc_739 ( N_GND_c_23_p N_noxref_39_c_10085_n ) capacitor c=0.0105197f //x=86.95 \
 //y=0 //x2=42.835 //y2=0.54
cc_740 ( N_GND_c_141_p N_noxref_39_c_10085_n ) capacitor c=0.0364139f \
 //x=43.49 //y=0 //x2=42.835 //y2=0.54
cc_741 ( N_GND_c_23_p N_noxref_39_c_10087_n ) capacitor c=0.00254232f \
 //x=86.95 //y=0 //x2=42.92 //y2=0.625
cc_742 ( N_GND_c_141_p N_noxref_39_c_10087_n ) capacitor c=0.0140304f \
 //x=43.49 //y=0 //x2=42.92 //y2=0.625
cc_743 ( N_GND_c_12_p N_noxref_39_c_10087_n ) capacitor c=0.0404137f //x=43.66 \
 //y=0 //x2=42.92 //y2=0.625
cc_744 ( N_GND_M24_noxref_d N_noxref_39_M25_noxref_d ) capacitor c=0.00162435f \
 //x=39.735 //y=0.875 //x2=40.71 //y2=0.91
cc_745 ( N_GND_c_11_p N_noxref_39_M26_noxref_s ) capacitor c=8.16352e-19 \
 //x=38.85 //y=0 //x2=41.815 //y2=0.375
cc_746 ( N_GND_c_12_p N_noxref_39_M26_noxref_s ) capacitor c=0.00183204f \
 //x=43.66 //y=0 //x2=41.815 //y2=0.375
cc_747 ( N_GND_c_23_p N_noxref_40_c_10133_n ) capacitor c=0.00517576f \
 //x=86.95 //y=0 //x2=45.135 //y2=1.59
cc_748 ( N_GND_c_160_p N_noxref_40_c_10133_n ) capacitor c=0.00111448f \
 //x=44.65 //y=0 //x2=45.135 //y2=1.59
cc_749 ( N_GND_c_167_p N_noxref_40_c_10133_n ) capacitor c=0.00180612f \
 //x=48.3 //y=0 //x2=45.135 //y2=1.59
cc_750 ( N_GND_M27_noxref_d N_noxref_40_c_10133_n ) capacitor c=0.00853078f \
 //x=44.545 //y=0.875 //x2=45.135 //y2=1.59
cc_751 ( N_GND_c_23_p N_noxref_40_c_10137_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=45.22 //y2=0.625
cc_752 ( N_GND_c_167_p N_noxref_40_c_10137_n ) capacitor c=0.0140928f //x=48.3 \
 //y=0 //x2=45.22 //y2=0.625
cc_753 ( N_GND_M27_noxref_d N_noxref_40_c_10137_n ) capacitor c=0.033954f \
 //x=44.545 //y=0.875 //x2=45.22 //y2=0.625
cc_754 ( N_GND_c_23_p N_noxref_40_c_10140_n ) capacitor c=0.0104386f //x=86.95 \
 //y=0 //x2=46.105 //y2=0.54
cc_755 ( N_GND_c_167_p N_noxref_40_c_10140_n ) capacitor c=0.0360726f //x=48.3 \
 //y=0 //x2=46.105 //y2=0.54
cc_756 ( N_GND_c_23_p N_noxref_40_M27_noxref_s ) capacitor c=0.00507657f \
 //x=86.95 //y=0 //x2=44.115 //y2=0.375
cc_757 ( N_GND_c_160_p N_noxref_40_M27_noxref_s ) capacitor c=0.0140928f \
 //x=44.65 //y=0 //x2=44.115 //y2=0.375
cc_758 ( N_GND_c_167_p N_noxref_40_M27_noxref_s ) capacitor c=0.0136651f \
 //x=48.3 //y=0 //x2=44.115 //y2=0.375
cc_759 ( N_GND_c_12_p N_noxref_40_M27_noxref_s ) capacitor c=0.0696963f \
 //x=43.66 //y=0 //x2=44.115 //y2=0.375
cc_760 ( N_GND_c_13_p N_noxref_40_M27_noxref_s ) capacitor c=3.31601e-19 \
 //x=48.47 //y=0 //x2=44.115 //y2=0.375
cc_761 ( N_GND_M27_noxref_d N_noxref_40_M27_noxref_s ) capacitor c=0.033718f \
 //x=44.545 //y=0.875 //x2=44.115 //y2=0.375
cc_762 ( N_GND_c_23_p N_noxref_41_c_10185_n ) capacitor c=0.00352952f \
 //x=86.95 //y=0 //x2=46.675 //y2=0.995
cc_763 ( N_GND_c_167_p N_noxref_41_c_10185_n ) capacitor c=0.00934524f \
 //x=48.3 //y=0 //x2=46.675 //y2=0.995
cc_764 ( N_GND_c_23_p N_noxref_41_c_10187_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=46.76 //y2=0.625
cc_765 ( N_GND_c_167_p N_noxref_41_c_10187_n ) capacitor c=0.0140928f //x=48.3 \
 //y=0 //x2=46.76 //y2=0.625
cc_766 ( N_GND_M27_noxref_d N_noxref_41_c_10187_n ) capacitor c=6.21394e-19 \
 //x=44.545 //y=0.875 //x2=46.76 //y2=0.625
cc_767 ( N_GND_c_23_p N_noxref_41_c_10190_n ) capacitor c=0.0105317f //x=86.95 \
 //y=0 //x2=47.645 //y2=0.54
cc_768 ( N_GND_c_167_p N_noxref_41_c_10190_n ) capacitor c=0.036415f //x=48.3 \
 //y=0 //x2=47.645 //y2=0.54
cc_769 ( N_GND_c_23_p N_noxref_41_c_10192_n ) capacitor c=0.00254232f \
 //x=86.95 //y=0 //x2=47.73 //y2=0.625
cc_770 ( N_GND_c_167_p N_noxref_41_c_10192_n ) capacitor c=0.0140304f //x=48.3 \
 //y=0 //x2=47.73 //y2=0.625
cc_771 ( N_GND_c_13_p N_noxref_41_c_10192_n ) capacitor c=0.0404137f //x=48.47 \
 //y=0 //x2=47.73 //y2=0.625
cc_772 ( N_GND_M27_noxref_d N_noxref_41_M28_noxref_d ) capacitor c=0.00162435f \
 //x=44.545 //y=0.875 //x2=45.52 //y2=0.91
cc_773 ( N_GND_c_12_p N_noxref_41_M29_noxref_s ) capacitor c=8.16352e-19 \
 //x=43.66 //y=0 //x2=46.625 //y2=0.375
cc_774 ( N_GND_c_13_p N_noxref_41_M29_noxref_s ) capacitor c=0.00183576f \
 //x=48.47 //y=0 //x2=46.625 //y2=0.375
cc_775 ( N_GND_c_23_p N_noxref_42_c_10237_n ) capacitor c=0.00517234f \
 //x=86.95 //y=0 //x2=50.05 //y2=1.58
cc_776 ( N_GND_c_173_p N_noxref_42_c_10237_n ) capacitor c=0.00112872f \
 //x=49.565 //y=0 //x2=50.05 //y2=1.58
cc_777 ( N_GND_c_180_p N_noxref_42_c_10237_n ) capacitor c=0.0018229f \
 //x=51.63 //y=0 //x2=50.05 //y2=1.58
cc_778 ( N_GND_M30_noxref_d N_noxref_42_c_10237_n ) capacitor c=0.008625f \
 //x=49.46 //y=0.865 //x2=50.05 //y2=1.58
cc_779 ( N_GND_c_23_p N_noxref_42_c_10241_n ) capacitor c=0.00259029f \
 //x=86.95 //y=0 //x2=50.135 //y2=0.615
cc_780 ( N_GND_c_180_p N_noxref_42_c_10241_n ) capacitor c=0.0146901f \
 //x=51.63 //y=0 //x2=50.135 //y2=0.615
cc_781 ( N_GND_M30_noxref_d N_noxref_42_c_10241_n ) capacitor c=0.033812f \
 //x=49.46 //y=0.865 //x2=50.135 //y2=0.615
cc_782 ( N_GND_c_13_p N_noxref_42_c_10244_n ) capacitor c=2.91423e-19 \
 //x=48.47 //y=0 //x2=50.135 //y2=1.495
cc_783 ( N_GND_c_23_p N_noxref_42_c_10245_n ) capacitor c=0.0106919f //x=86.95 \
 //y=0 //x2=51.02 //y2=0.53
cc_784 ( N_GND_c_180_p N_noxref_42_c_10245_n ) capacitor c=0.0374253f \
 //x=51.63 //y=0 //x2=51.02 //y2=0.53
cc_785 ( N_GND_c_23_p N_noxref_42_c_10247_n ) capacitor c=0.00258845f \
 //x=86.95 //y=0 //x2=51.105 //y2=0.615
cc_786 ( N_GND_c_180_p N_noxref_42_c_10247_n ) capacitor c=0.0146256f \
 //x=51.63 //y=0 //x2=51.105 //y2=0.615
cc_787 ( N_GND_c_14_p N_noxref_42_c_10247_n ) capacitor c=0.0431718f //x=51.8 \
 //y=0 //x2=51.105 //y2=0.615
cc_788 ( N_GND_c_23_p N_noxref_42_M30_noxref_s ) capacitor c=0.00259029f \
 //x=86.95 //y=0 //x2=49.03 //y2=0.365
cc_789 ( N_GND_c_173_p N_noxref_42_M30_noxref_s ) capacitor c=0.0146901f \
 //x=49.565 //y=0 //x2=49.03 //y2=0.365
cc_790 ( N_GND_c_13_p N_noxref_42_M30_noxref_s ) capacitor c=0.0583534f \
 //x=48.47 //y=0 //x2=49.03 //y2=0.365
cc_791 ( N_GND_c_14_p N_noxref_42_M30_noxref_s ) capacitor c=0.00198098f \
 //x=51.8 //y=0 //x2=49.03 //y2=0.365
cc_792 ( N_GND_M30_noxref_d N_noxref_42_M30_noxref_s ) capacitor c=0.0334197f \
 //x=49.46 //y=0.865 //x2=49.03 //y2=0.365
cc_793 ( N_GND_c_23_p N_noxref_43_c_10288_n ) capacitor c=0.00517576f \
 //x=86.95 //y=0 //x2=53.275 //y2=1.59
cc_794 ( N_GND_c_293_p N_noxref_43_c_10288_n ) capacitor c=0.00111448f \
 //x=52.79 //y=0 //x2=53.275 //y2=1.59
cc_795 ( N_GND_c_294_p N_noxref_43_c_10288_n ) capacitor c=0.00180612f \
 //x=56.44 //y=0 //x2=53.275 //y2=1.59
cc_796 ( N_GND_M32_noxref_d N_noxref_43_c_10288_n ) capacitor c=0.00853078f \
 //x=52.685 //y=0.875 //x2=53.275 //y2=1.59
cc_797 ( N_GND_c_23_p N_noxref_43_c_10292_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=53.36 //y2=0.625
cc_798 ( N_GND_c_294_p N_noxref_43_c_10292_n ) capacitor c=0.0140928f \
 //x=56.44 //y=0 //x2=53.36 //y2=0.625
cc_799 ( N_GND_M32_noxref_d N_noxref_43_c_10292_n ) capacitor c=0.033954f \
 //x=52.685 //y=0.875 //x2=53.36 //y2=0.625
cc_800 ( N_GND_c_23_p N_noxref_43_c_10295_n ) capacitor c=0.0104506f //x=86.95 \
 //y=0 //x2=54.245 //y2=0.54
cc_801 ( N_GND_c_294_p N_noxref_43_c_10295_n ) capacitor c=0.0360726f \
 //x=56.44 //y=0 //x2=54.245 //y2=0.54
cc_802 ( N_GND_c_23_p N_noxref_43_M32_noxref_s ) capacitor c=0.00507657f \
 //x=86.95 //y=0 //x2=52.255 //y2=0.375
cc_803 ( N_GND_c_293_p N_noxref_43_M32_noxref_s ) capacitor c=0.0140928f \
 //x=52.79 //y=0 //x2=52.255 //y2=0.375
cc_804 ( N_GND_c_294_p N_noxref_43_M32_noxref_s ) capacitor c=0.0131437f \
 //x=56.44 //y=0 //x2=52.255 //y2=0.375
cc_805 ( N_GND_c_14_p N_noxref_43_M32_noxref_s ) capacitor c=0.0696963f \
 //x=51.8 //y=0 //x2=52.255 //y2=0.375
cc_806 ( N_GND_c_15_p N_noxref_43_M32_noxref_s ) capacitor c=3.31601e-19 \
 //x=56.61 //y=0 //x2=52.255 //y2=0.375
cc_807 ( N_GND_M32_noxref_d N_noxref_43_M32_noxref_s ) capacitor c=0.033718f \
 //x=52.685 //y=0.875 //x2=52.255 //y2=0.375
cc_808 ( N_GND_c_23_p N_noxref_44_c_10337_n ) capacitor c=0.00352952f \
 //x=86.95 //y=0 //x2=54.815 //y2=0.995
cc_809 ( N_GND_c_294_p N_noxref_44_c_10337_n ) capacitor c=0.00934524f \
 //x=56.44 //y=0 //x2=54.815 //y2=0.995
cc_810 ( N_GND_c_23_p N_noxref_44_c_10339_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=54.9 //y2=0.625
cc_811 ( N_GND_c_294_p N_noxref_44_c_10339_n ) capacitor c=0.0140928f \
 //x=56.44 //y=0 //x2=54.9 //y2=0.625
cc_812 ( N_GND_M32_noxref_d N_noxref_44_c_10339_n ) capacitor c=6.21394e-19 \
 //x=52.685 //y=0.875 //x2=54.9 //y2=0.625
cc_813 ( N_GND_c_23_p N_noxref_44_c_10342_n ) capacitor c=0.0105317f //x=86.95 \
 //y=0 //x2=55.785 //y2=0.54
cc_814 ( N_GND_c_294_p N_noxref_44_c_10342_n ) capacitor c=0.036415f //x=56.44 \
 //y=0 //x2=55.785 //y2=0.54
cc_815 ( N_GND_c_23_p N_noxref_44_c_10344_n ) capacitor c=0.00254232f \
 //x=86.95 //y=0 //x2=55.87 //y2=0.625
cc_816 ( N_GND_c_294_p N_noxref_44_c_10344_n ) capacitor c=0.0140304f \
 //x=56.44 //y=0 //x2=55.87 //y2=0.625
cc_817 ( N_GND_c_15_p N_noxref_44_c_10344_n ) capacitor c=0.0404137f //x=56.61 \
 //y=0 //x2=55.87 //y2=0.625
cc_818 ( N_GND_M32_noxref_d N_noxref_44_M33_noxref_d ) capacitor c=0.00162435f \
 //x=52.685 //y=0.875 //x2=53.66 //y2=0.91
cc_819 ( N_GND_c_14_p N_noxref_44_M34_noxref_s ) capacitor c=8.16352e-19 \
 //x=51.8 //y=0 //x2=54.765 //y2=0.375
cc_820 ( N_GND_c_15_p N_noxref_44_M34_noxref_s ) capacitor c=0.00183204f \
 //x=56.61 //y=0 //x2=54.765 //y2=0.375
cc_821 ( N_GND_c_23_p N_noxref_45_c_10389_n ) capacitor c=0.00517576f \
 //x=86.95 //y=0 //x2=58.085 //y2=1.59
cc_822 ( N_GND_c_227_p N_noxref_45_c_10389_n ) capacitor c=0.00111448f \
 //x=57.6 //y=0 //x2=58.085 //y2=1.59
cc_823 ( N_GND_c_234_p N_noxref_45_c_10389_n ) capacitor c=0.00180612f \
 //x=61.25 //y=0 //x2=58.085 //y2=1.59
cc_824 ( N_GND_M35_noxref_d N_noxref_45_c_10389_n ) capacitor c=0.00853078f \
 //x=57.495 //y=0.875 //x2=58.085 //y2=1.59
cc_825 ( N_GND_c_23_p N_noxref_45_c_10393_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=58.17 //y2=0.625
cc_826 ( N_GND_c_234_p N_noxref_45_c_10393_n ) capacitor c=0.0140928f \
 //x=61.25 //y=0 //x2=58.17 //y2=0.625
cc_827 ( N_GND_M35_noxref_d N_noxref_45_c_10393_n ) capacitor c=0.033954f \
 //x=57.495 //y=0.875 //x2=58.17 //y2=0.625
cc_828 ( N_GND_c_23_p N_noxref_45_c_10396_n ) capacitor c=0.0104506f //x=86.95 \
 //y=0 //x2=59.055 //y2=0.54
cc_829 ( N_GND_c_234_p N_noxref_45_c_10396_n ) capacitor c=0.0360726f \
 //x=61.25 //y=0 //x2=59.055 //y2=0.54
cc_830 ( N_GND_c_23_p N_noxref_45_M35_noxref_s ) capacitor c=0.00507657f \
 //x=86.95 //y=0 //x2=57.065 //y2=0.375
cc_831 ( N_GND_c_227_p N_noxref_45_M35_noxref_s ) capacitor c=0.0140928f \
 //x=57.6 //y=0 //x2=57.065 //y2=0.375
cc_832 ( N_GND_c_234_p N_noxref_45_M35_noxref_s ) capacitor c=0.0131437f \
 //x=61.25 //y=0 //x2=57.065 //y2=0.375
cc_833 ( N_GND_c_15_p N_noxref_45_M35_noxref_s ) capacitor c=0.0696963f \
 //x=56.61 //y=0 //x2=57.065 //y2=0.375
cc_834 ( N_GND_c_16_p N_noxref_45_M35_noxref_s ) capacitor c=3.31601e-19 \
 //x=61.42 //y=0 //x2=57.065 //y2=0.375
cc_835 ( N_GND_M35_noxref_d N_noxref_45_M35_noxref_s ) capacitor c=0.033718f \
 //x=57.495 //y=0.875 //x2=57.065 //y2=0.375
cc_836 ( N_GND_c_23_p N_noxref_46_c_10438_n ) capacitor c=0.00352952f \
 //x=86.95 //y=0 //x2=59.625 //y2=0.995
cc_837 ( N_GND_c_234_p N_noxref_46_c_10438_n ) capacitor c=0.00934524f \
 //x=61.25 //y=0 //x2=59.625 //y2=0.995
cc_838 ( N_GND_c_23_p N_noxref_46_c_10440_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=59.71 //y2=0.625
cc_839 ( N_GND_c_234_p N_noxref_46_c_10440_n ) capacitor c=0.0140928f \
 //x=61.25 //y=0 //x2=59.71 //y2=0.625
cc_840 ( N_GND_M35_noxref_d N_noxref_46_c_10440_n ) capacitor c=6.21394e-19 \
 //x=57.495 //y=0.875 //x2=59.71 //y2=0.625
cc_841 ( N_GND_c_23_p N_noxref_46_c_10443_n ) capacitor c=0.0105197f //x=86.95 \
 //y=0 //x2=60.595 //y2=0.54
cc_842 ( N_GND_c_234_p N_noxref_46_c_10443_n ) capacitor c=0.036368f //x=61.25 \
 //y=0 //x2=60.595 //y2=0.54
cc_843 ( N_GND_c_23_p N_noxref_46_c_10445_n ) capacitor c=0.00254232f \
 //x=86.95 //y=0 //x2=60.68 //y2=0.625
cc_844 ( N_GND_c_234_p N_noxref_46_c_10445_n ) capacitor c=0.0140304f \
 //x=61.25 //y=0 //x2=60.68 //y2=0.625
cc_845 ( N_GND_c_16_p N_noxref_46_c_10445_n ) capacitor c=0.0404137f //x=61.42 \
 //y=0 //x2=60.68 //y2=0.625
cc_846 ( N_GND_M35_noxref_d N_noxref_46_M36_noxref_d ) capacitor c=0.00162435f \
 //x=57.495 //y=0.875 //x2=58.47 //y2=0.91
cc_847 ( N_GND_c_15_p N_noxref_46_M37_noxref_s ) capacitor c=8.16352e-19 \
 //x=56.61 //y=0 //x2=59.575 //y2=0.375
cc_848 ( N_GND_c_16_p N_noxref_46_M37_noxref_s ) capacitor c=0.00183576f \
 //x=61.42 //y=0 //x2=59.575 //y2=0.375
cc_849 ( N_GND_c_23_p N_noxref_47_c_10491_n ) capacitor c=0.00517234f \
 //x=86.95 //y=0 //x2=63 //y2=1.58
cc_850 ( N_GND_c_303_p N_noxref_47_c_10491_n ) capacitor c=0.00112872f \
 //x=62.515 //y=0 //x2=63 //y2=1.58
cc_851 ( N_GND_c_304_p N_noxref_47_c_10491_n ) capacitor c=0.0018229f \
 //x=64.58 //y=0 //x2=63 //y2=1.58
cc_852 ( N_GND_M38_noxref_d N_noxref_47_c_10491_n ) capacitor c=0.008625f \
 //x=62.41 //y=0.865 //x2=63 //y2=1.58
cc_853 ( N_GND_c_23_p N_noxref_47_c_10495_n ) capacitor c=0.00259029f \
 //x=86.95 //y=0 //x2=63.085 //y2=0.615
cc_854 ( N_GND_c_304_p N_noxref_47_c_10495_n ) capacitor c=0.0146901f \
 //x=64.58 //y=0 //x2=63.085 //y2=0.615
cc_855 ( N_GND_M38_noxref_d N_noxref_47_c_10495_n ) capacitor c=0.033812f \
 //x=62.41 //y=0.865 //x2=63.085 //y2=0.615
cc_856 ( N_GND_c_16_p N_noxref_47_c_10498_n ) capacitor c=2.91423e-19 \
 //x=61.42 //y=0 //x2=63.085 //y2=1.495
cc_857 ( N_GND_c_23_p N_noxref_47_c_10499_n ) capacitor c=0.0106919f //x=86.95 \
 //y=0 //x2=63.97 //y2=0.53
cc_858 ( N_GND_c_304_p N_noxref_47_c_10499_n ) capacitor c=0.0374253f \
 //x=64.58 //y=0 //x2=63.97 //y2=0.53
cc_859 ( N_GND_c_23_p N_noxref_47_c_10501_n ) capacitor c=0.00258845f \
 //x=86.95 //y=0 //x2=64.055 //y2=0.615
cc_860 ( N_GND_c_304_p N_noxref_47_c_10501_n ) capacitor c=0.0146256f \
 //x=64.58 //y=0 //x2=64.055 //y2=0.615
cc_861 ( N_GND_c_17_p N_noxref_47_c_10501_n ) capacitor c=0.0431718f //x=64.75 \
 //y=0 //x2=64.055 //y2=0.615
cc_862 ( N_GND_c_23_p N_noxref_47_M38_noxref_s ) capacitor c=0.00259029f \
 //x=86.95 //y=0 //x2=61.98 //y2=0.365
cc_863 ( N_GND_c_303_p N_noxref_47_M38_noxref_s ) capacitor c=0.0146901f \
 //x=62.515 //y=0 //x2=61.98 //y2=0.365
cc_864 ( N_GND_c_16_p N_noxref_47_M38_noxref_s ) capacitor c=0.0583534f \
 //x=61.42 //y=0 //x2=61.98 //y2=0.365
cc_865 ( N_GND_c_17_p N_noxref_47_M38_noxref_s ) capacitor c=0.00198098f \
 //x=64.75 //y=0 //x2=61.98 //y2=0.365
cc_866 ( N_GND_M38_noxref_d N_noxref_47_M38_noxref_s ) capacitor c=0.0334197f \
 //x=62.41 //y=0.865 //x2=61.98 //y2=0.365
cc_867 ( N_GND_c_23_p N_noxref_48_c_10542_n ) capacitor c=0.00517576f \
 //x=86.95 //y=0 //x2=66.225 //y2=1.59
cc_868 ( N_GND_c_305_p N_noxref_48_c_10542_n ) capacitor c=0.00111448f \
 //x=65.74 //y=0 //x2=66.225 //y2=1.59
cc_869 ( N_GND_c_306_p N_noxref_48_c_10542_n ) capacitor c=0.00180612f \
 //x=69.39 //y=0 //x2=66.225 //y2=1.59
cc_870 ( N_GND_M40_noxref_d N_noxref_48_c_10542_n ) capacitor c=0.00853078f \
 //x=65.635 //y=0.875 //x2=66.225 //y2=1.59
cc_871 ( N_GND_c_23_p N_noxref_48_c_10546_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=66.31 //y2=0.625
cc_872 ( N_GND_c_306_p N_noxref_48_c_10546_n ) capacitor c=0.0140928f \
 //x=69.39 //y=0 //x2=66.31 //y2=0.625
cc_873 ( N_GND_M40_noxref_d N_noxref_48_c_10546_n ) capacitor c=0.033954f \
 //x=65.635 //y=0.875 //x2=66.31 //y2=0.625
cc_874 ( N_GND_c_23_p N_noxref_48_c_10549_n ) capacitor c=0.0104506f //x=86.95 \
 //y=0 //x2=67.195 //y2=0.54
cc_875 ( N_GND_c_306_p N_noxref_48_c_10549_n ) capacitor c=0.0360726f \
 //x=69.39 //y=0 //x2=67.195 //y2=0.54
cc_876 ( N_GND_c_23_p N_noxref_48_M40_noxref_s ) capacitor c=0.00507657f \
 //x=86.95 //y=0 //x2=65.205 //y2=0.375
cc_877 ( N_GND_c_305_p N_noxref_48_M40_noxref_s ) capacitor c=0.0140928f \
 //x=65.74 //y=0 //x2=65.205 //y2=0.375
cc_878 ( N_GND_c_306_p N_noxref_48_M40_noxref_s ) capacitor c=0.0131437f \
 //x=69.39 //y=0 //x2=65.205 //y2=0.375
cc_879 ( N_GND_c_17_p N_noxref_48_M40_noxref_s ) capacitor c=0.0696963f \
 //x=64.75 //y=0 //x2=65.205 //y2=0.375
cc_880 ( N_GND_c_18_p N_noxref_48_M40_noxref_s ) capacitor c=3.31601e-19 \
 //x=69.56 //y=0 //x2=65.205 //y2=0.375
cc_881 ( N_GND_M40_noxref_d N_noxref_48_M40_noxref_s ) capacitor c=0.033718f \
 //x=65.635 //y=0.875 //x2=65.205 //y2=0.375
cc_882 ( N_GND_c_23_p N_noxref_49_c_10591_n ) capacitor c=0.00352952f \
 //x=86.95 //y=0 //x2=67.765 //y2=0.995
cc_883 ( N_GND_c_306_p N_noxref_49_c_10591_n ) capacitor c=0.00934524f \
 //x=69.39 //y=0 //x2=67.765 //y2=0.995
cc_884 ( N_GND_c_23_p N_noxref_49_c_10593_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=67.85 //y2=0.625
cc_885 ( N_GND_c_306_p N_noxref_49_c_10593_n ) capacitor c=0.0140928f \
 //x=69.39 //y=0 //x2=67.85 //y2=0.625
cc_886 ( N_GND_M40_noxref_d N_noxref_49_c_10593_n ) capacitor c=6.21394e-19 \
 //x=65.635 //y=0.875 //x2=67.85 //y2=0.625
cc_887 ( N_GND_c_23_p N_noxref_49_c_10596_n ) capacitor c=0.0105197f //x=86.95 \
 //y=0 //x2=68.735 //y2=0.54
cc_888 ( N_GND_c_306_p N_noxref_49_c_10596_n ) capacitor c=0.0364139f \
 //x=69.39 //y=0 //x2=68.735 //y2=0.54
cc_889 ( N_GND_c_23_p N_noxref_49_c_10598_n ) capacitor c=0.00254232f \
 //x=86.95 //y=0 //x2=68.82 //y2=0.625
cc_890 ( N_GND_c_306_p N_noxref_49_c_10598_n ) capacitor c=0.0140304f \
 //x=69.39 //y=0 //x2=68.82 //y2=0.625
cc_891 ( N_GND_c_18_p N_noxref_49_c_10598_n ) capacitor c=0.0404137f //x=69.56 \
 //y=0 //x2=68.82 //y2=0.625
cc_892 ( N_GND_M40_noxref_d N_noxref_49_M41_noxref_d ) capacitor c=0.00162435f \
 //x=65.635 //y=0.875 //x2=66.61 //y2=0.91
cc_893 ( N_GND_c_17_p N_noxref_49_M42_noxref_s ) capacitor c=8.16352e-19 \
 //x=64.75 //y=0 //x2=67.715 //y2=0.375
cc_894 ( N_GND_c_18_p N_noxref_49_M42_noxref_s ) capacitor c=0.00183204f \
 //x=69.56 //y=0 //x2=67.715 //y2=0.375
cc_895 ( N_GND_c_23_p N_noxref_50_c_10644_n ) capacitor c=0.00517576f \
 //x=86.95 //y=0 //x2=71.035 //y2=1.59
cc_896 ( N_GND_c_237_p N_noxref_50_c_10644_n ) capacitor c=0.00111448f \
 //x=70.55 //y=0 //x2=71.035 //y2=1.59
cc_897 ( N_GND_c_244_p N_noxref_50_c_10644_n ) capacitor c=0.00180612f \
 //x=74.2 //y=0 //x2=71.035 //y2=1.59
cc_898 ( N_GND_M43_noxref_d N_noxref_50_c_10644_n ) capacitor c=0.00853078f \
 //x=70.445 //y=0.875 //x2=71.035 //y2=1.59
cc_899 ( N_GND_c_23_p N_noxref_50_c_10648_n ) capacitor c=0.00254475f \
 //x=86.95 //y=0 //x2=71.12 //y2=0.625
cc_900 ( N_GND_c_244_p N_noxref_50_c_10648_n ) capacitor c=0.0140928f //x=74.2 \
 //y=0 //x2=71.12 //y2=0.625
cc_901 ( N_GND_M43_noxref_d N_noxref_50_c_10648_n ) capacitor c=0.033954f \
 //x=70.445 //y=0.875 //x2=71.12 //y2=0.625
cc_902 ( N_GND_c_23_p N_noxref_50_c_10651_n ) capacitor c=0.0105304f //x=86.95 \
 //y=0 //x2=72.005 //y2=0.54
cc_903 ( N_GND_c_244_p N_noxref_50_c_10651_n ) capacitor c=0.0361183f //x=74.2 \
 //y=0 //x2=72.005 //y2=0.54
cc_904 ( N_GND_c_23_p N_noxref_50_M43_noxref_s ) capacitor c=0.00531539f \
 //x=86.95 //y=0 //x2=70.015 //y2=0.375
cc_905 ( N_GND_c_237_p N_noxref_50_M43_noxref_s ) capacitor c=0.0140928f \
 //x=70.55 //y=0 //x2=70.015 //y2=0.375
cc_906 ( N_GND_c_244_p N_noxref_50_M43_noxref_s ) capacitor c=0.0133155f \
 //x=74.2 //y=0 //x2=70.015 //y2=0.375
cc_907 ( N_GND_c_18_p N_noxref_50_M43_noxref_s ) capacitor c=0.0696963f \
 //x=69.56 //y=0 //x2=70.015 //y2=0.375
cc_908 ( N_GND_c_19_p N_noxref_50_M43_noxref_s ) capacitor c=3.31601e-19 \
 //x=74.37 //y=0 //x2=70.015 //y2=0.375
cc_909 ( N_GND_M43_noxref_d N_noxref_50_M43_noxref_s ) capacitor c=0.033718f \
 //x=70.445 //y=0.875 //x2=70.015 //y2=0.375
cc_910 ( N_GND_c_23_p N_noxref_51_c_10695_n ) capacitor c=0.00375441f \
 //x=86.95 //y=0 //x2=72.575 //y2=0.995
cc_911 ( N_GND_c_244_p N_noxref_51_c_10695_n ) capacitor c=0.00944862f \
 //x=74.2 //y=0 //x2=72.575 //y2=0.995
cc_912 ( N_GND_c_23_p N_noxref_51_c_10697_n ) capacitor c=0.00277579f \
 //x=86.95 //y=0 //x2=72.66 //y2=0.625
cc_913 ( N_GND_c_244_p N_noxref_51_c_10697_n ) capacitor c=0.0142586f //x=74.2 \
 //y=0 //x2=72.66 //y2=0.625
cc_914 ( N_GND_M43_noxref_d N_noxref_51_c_10697_n ) capacitor c=6.21394e-19 \
 //x=70.445 //y=0.875 //x2=72.66 //y2=0.625
cc_915 ( N_GND_c_23_p N_noxref_51_c_10700_n ) capacitor c=0.0114469f //x=86.95 \
 //y=0 //x2=73.545 //y2=0.54
cc_916 ( N_GND_c_244_p N_noxref_51_c_10700_n ) capacitor c=0.0365589f //x=74.2 \
 //y=0 //x2=73.545 //y2=0.54
cc_917 ( N_GND_c_23_p N_noxref_51_c_10702_n ) capacitor c=0.00277442f \
 //x=86.95 //y=0 //x2=73.63 //y2=0.625
cc_918 ( N_GND_c_244_p N_noxref_51_c_10702_n ) capacitor c=0.014197f //x=74.2 \
 //y=0 //x2=73.63 //y2=0.625
cc_919 ( N_GND_c_19_p N_noxref_51_c_10702_n ) capacitor c=0.0404137f //x=74.37 \
 //y=0 //x2=73.63 //y2=0.625
cc_920 ( N_GND_M43_noxref_d N_noxref_51_M44_noxref_d ) capacitor c=0.00162435f \
 //x=70.445 //y=0.875 //x2=71.42 //y2=0.91
cc_921 ( N_GND_c_18_p N_noxref_51_M45_noxref_s ) capacitor c=8.16352e-19 \
 //x=69.56 //y=0 //x2=72.525 //y2=0.375
cc_922 ( N_GND_c_19_p N_noxref_51_M45_noxref_s ) capacitor c=0.00183576f \
 //x=74.37 //y=0 //x2=72.525 //y2=0.375
cc_923 ( N_GND_c_23_p N_noxref_52_c_10747_n ) capacitor c=0.00542069f \
 //x=86.95 //y=0 //x2=75.95 //y2=1.58
cc_924 ( N_GND_c_342_p N_noxref_52_c_10747_n ) capacitor c=0.00112963f \
 //x=75.465 //y=0 //x2=75.95 //y2=1.58
cc_925 ( N_GND_c_349_p N_noxref_52_c_10747_n ) capacitor c=0.00182382f \
 //x=77.53 //y=0 //x2=75.95 //y2=1.58
cc_926 ( N_GND_M46_noxref_d N_noxref_52_c_10747_n ) capacitor c=0.00890129f \
 //x=75.36 //y=0.865 //x2=75.95 //y2=1.58
cc_927 ( N_GND_c_23_p N_noxref_52_c_10751_n ) capacitor c=0.00282937f \
 //x=86.95 //y=0 //x2=76.035 //y2=0.615
cc_928 ( N_GND_c_349_p N_noxref_52_c_10751_n ) capacitor c=0.0148639f \
 //x=77.53 //y=0 //x2=76.035 //y2=0.615
cc_929 ( N_GND_M46_noxref_d N_noxref_52_c_10751_n ) capacitor c=0.033812f \
 //x=75.36 //y=0.865 //x2=76.035 //y2=0.615
cc_930 ( N_GND_c_19_p N_noxref_52_c_10754_n ) capacitor c=2.91423e-19 \
 //x=74.37 //y=0 //x2=76.035 //y2=1.495
cc_931 ( N_GND_c_23_p N_noxref_52_c_10755_n ) capacitor c=0.0116329f //x=86.95 \
 //y=0 //x2=76.92 //y2=0.53
cc_932 ( N_GND_c_349_p N_noxref_52_c_10755_n ) capacitor c=0.0375167f \
 //x=77.53 //y=0 //x2=76.92 //y2=0.53
cc_933 ( N_GND_c_23_p N_noxref_52_c_10757_n ) capacitor c=0.00282863f \
 //x=86.95 //y=0 //x2=77.005 //y2=0.615
cc_934 ( N_GND_c_349_p N_noxref_52_c_10757_n ) capacitor c=0.0148003f \
 //x=77.53 //y=0 //x2=77.005 //y2=0.615
cc_935 ( N_GND_c_20_p N_noxref_52_c_10757_n ) capacitor c=0.0427915f //x=77.7 \
 //y=0 //x2=77.005 //y2=0.615
cc_936 ( N_GND_c_23_p N_noxref_52_M46_noxref_s ) capacitor c=0.00282937f \
 //x=86.95 //y=0 //x2=74.93 //y2=0.365
cc_937 ( N_GND_c_342_p N_noxref_52_M46_noxref_s ) capacitor c=0.0148639f \
 //x=75.465 //y=0 //x2=74.93 //y2=0.365
cc_938 ( N_GND_c_19_p N_noxref_52_M46_noxref_s ) capacitor c=0.0583534f \
 //x=74.37 //y=0 //x2=74.93 //y2=0.365
cc_939 ( N_GND_c_20_p N_noxref_52_M46_noxref_s ) capacitor c=0.00198098f \
 //x=77.7 //y=0 //x2=74.93 //y2=0.365
cc_940 ( N_GND_M46_noxref_d N_noxref_52_M46_noxref_s ) capacitor c=0.0334197f \
 //x=75.36 //y=0.865 //x2=74.93 //y2=0.365
cc_941 ( N_GND_c_23_p N_noxref_53_c_10798_n ) capacitor c=0.00547799f \
 //x=86.95 //y=0 //x2=79.28 //y2=1.58
cc_942 ( N_GND_c_388_p N_noxref_53_c_10798_n ) capacitor c=0.00112964f \
 //x=78.795 //y=0 //x2=79.28 //y2=1.58
cc_943 ( N_GND_c_395_p N_noxref_53_c_10798_n ) capacitor c=0.00182382f \
 //x=80.86 //y=0 //x2=79.28 //y2=1.58
cc_944 ( N_GND_M48_noxref_d N_noxref_53_c_10798_n ) capacitor c=0.0092166f \
 //x=78.69 //y=0.865 //x2=79.28 //y2=1.58
cc_945 ( N_GND_c_23_p N_noxref_53_c_10802_n ) capacitor c=0.00282937f \
 //x=86.95 //y=0 //x2=79.365 //y2=0.615
cc_946 ( N_GND_c_395_p N_noxref_53_c_10802_n ) capacitor c=0.0148639f \
 //x=80.86 //y=0 //x2=79.365 //y2=0.615
cc_947 ( N_GND_M48_noxref_d N_noxref_53_c_10802_n ) capacitor c=0.0336822f \
 //x=78.69 //y=0.865 //x2=79.365 //y2=0.615
cc_948 ( N_GND_c_20_p N_noxref_53_c_10805_n ) capacitor c=2.91423e-19 //x=77.7 \
 //y=0 //x2=79.365 //y2=1.495
cc_949 ( N_GND_c_23_p N_noxref_53_c_10806_n ) capacitor c=0.00972782f \
 //x=86.95 //y=0 //x2=80.25 //y2=0.53
cc_950 ( N_GND_c_395_p N_noxref_53_c_10806_n ) capacitor c=0.0375243f \
 //x=80.86 //y=0 //x2=80.25 //y2=0.53
cc_951 ( N_GND_c_23_p N_noxref_53_c_10808_n ) capacitor c=0.00212661f \
 //x=86.95 //y=0 //x2=80.335 //y2=0.615
cc_952 ( N_GND_c_395_p N_noxref_53_c_10808_n ) capacitor c=0.0143168f \
 //x=80.86 //y=0 //x2=80.335 //y2=0.615
cc_953 ( N_GND_c_21_p N_noxref_53_c_10808_n ) capacitor c=0.0554337f //x=81.03 \
 //y=0 //x2=80.335 //y2=0.615
cc_954 ( N_GND_c_23_p N_noxref_53_M48_noxref_s ) capacitor c=0.00282937f \
 //x=86.95 //y=0 //x2=78.26 //y2=0.365
cc_955 ( N_GND_c_388_p N_noxref_53_M48_noxref_s ) capacitor c=0.0148639f \
 //x=78.795 //y=0 //x2=78.26 //y2=0.365
cc_956 ( N_GND_c_20_p N_noxref_53_M48_noxref_s ) capacitor c=0.0587986f \
 //x=77.7 //y=0 //x2=78.26 //y2=0.365
cc_957 ( N_GND_c_21_p N_noxref_53_M48_noxref_s ) capacitor c=0.00181744f \
 //x=81.03 //y=0 //x2=78.26 //y2=0.365
cc_958 ( N_GND_M48_noxref_d N_noxref_53_M48_noxref_s ) capacitor c=0.0333456f \
 //x=78.69 //y=0.865 //x2=78.26 //y2=0.365
cc_959 ( N_GND_c_398_p N_noxref_54_c_10855_n ) capacitor c=8.01905e-19 \
 //x=82.125 //y=0 //x2=82.61 //y2=1.58
cc_960 ( N_GND_c_404_p N_noxref_54_c_10855_n ) capacitor c=0.00161527f \
 //x=84.19 //y=0 //x2=82.61 //y2=1.58
cc_961 ( N_GND_M50_noxref_d N_noxref_54_c_10855_n ) capacitor c=0.0073276f \
 //x=82.02 //y=0.865 //x2=82.61 //y2=1.58
cc_962 ( N_GND_c_23_p N_noxref_54_c_10858_n ) capacitor c=0.00212661f \
 //x=86.95 //y=0 //x2=82.695 //y2=0.615
cc_963 ( N_GND_c_404_p N_noxref_54_c_10858_n ) capacitor c=0.0143168f \
 //x=84.19 //y=0 //x2=82.695 //y2=0.615
cc_964 ( N_GND_M50_noxref_d N_noxref_54_c_10858_n ) capacitor c=0.0336587f \
 //x=82.02 //y=0.865 //x2=82.695 //y2=0.615
cc_965 ( N_GND_c_21_p N_noxref_54_c_10861_n ) capacitor c=2.91423e-19 \
 //x=81.03 //y=0 //x2=82.695 //y2=1.495
cc_966 ( N_GND_c_23_p N_noxref_54_c_10862_n ) capacitor c=0.00884129f \
 //x=86.95 //y=0 //x2=83.58 //y2=0.53
cc_967 ( N_GND_c_404_p N_noxref_54_c_10862_n ) capacitor c=0.0373651f \
 //x=84.19 //y=0 //x2=83.58 //y2=0.53
cc_968 ( N_GND_c_23_p N_noxref_54_c_10864_n ) capacitor c=0.00212661f \
 //x=86.95 //y=0 //x2=83.665 //y2=0.615
cc_969 ( N_GND_c_404_p N_noxref_54_c_10864_n ) capacitor c=0.0143168f \
 //x=84.19 //y=0 //x2=83.665 //y2=0.615
cc_970 ( N_GND_c_22_p N_noxref_54_c_10864_n ) capacitor c=0.0548042f //x=84.36 \
 //y=0 //x2=83.665 //y2=0.615
cc_971 ( N_GND_c_23_p N_noxref_54_M50_noxref_s ) capacitor c=0.00212661f \
 //x=86.95 //y=0 //x2=81.59 //y2=0.365
cc_972 ( N_GND_c_398_p N_noxref_54_M50_noxref_s ) capacitor c=0.0143168f \
 //x=82.125 //y=0 //x2=81.59 //y2=0.365
cc_973 ( N_GND_c_21_p N_noxref_54_M50_noxref_s ) capacitor c=0.0561194f \
 //x=81.03 //y=0 //x2=81.59 //y2=0.365
cc_974 ( N_GND_c_22_p N_noxref_54_M50_noxref_s ) capacitor c=0.0022128f \
 //x=84.36 //y=0 //x2=81.59 //y2=0.365
cc_975 ( N_GND_M50_noxref_d N_noxref_54_M50_noxref_s ) capacitor c=0.0332904f \
 //x=82.02 //y=0.865 //x2=81.59 //y2=0.365
cc_976 ( N_GND_c_457_p N_noxref_55_c_10910_n ) capacitor c=8.01912e-19 \
 //x=85.455 //y=0 //x2=85.94 //y2=1.58
cc_977 ( N_GND_c_2_p N_noxref_55_c_10910_n ) capacitor c=0.00161527f //x=86.95 \
 //y=0 //x2=85.94 //y2=1.58
cc_978 ( N_GND_M52_noxref_d N_noxref_55_c_10910_n ) capacitor c=0.0073482f \
 //x=85.35 //y=0.865 //x2=85.94 //y2=1.58
cc_979 ( N_GND_c_23_p N_noxref_55_c_10913_n ) capacitor c=0.00212661f \
 //x=86.95 //y=0 //x2=86.025 //y2=0.615
cc_980 ( N_GND_c_2_p N_noxref_55_c_10913_n ) capacitor c=0.0143168f //x=86.95 \
 //y=0 //x2=86.025 //y2=0.615
cc_981 ( N_GND_M52_noxref_d N_noxref_55_c_10913_n ) capacitor c=0.0336587f \
 //x=85.35 //y=0.865 //x2=86.025 //y2=0.615
cc_982 ( N_GND_c_22_p N_noxref_55_c_10916_n ) capacitor c=2.91423e-19 \
 //x=84.36 //y=0 //x2=86.025 //y2=1.495
cc_983 ( N_GND_c_23_p N_noxref_55_c_10917_n ) capacitor c=0.0127012f //x=86.95 \
 //y=0 //x2=86.91 //y2=0.53
cc_984 ( N_GND_c_2_p N_noxref_55_c_10917_n ) capacitor c=0.0371788f //x=86.95 \
 //y=0 //x2=86.91 //y2=0.53
cc_985 ( N_GND_c_23_p N_noxref_55_c_10919_n ) capacitor c=0.00719686f \
 //x=86.95 //y=0 //x2=86.995 //y2=0.615
cc_986 ( N_GND_c_2_p N_noxref_55_c_10919_n ) capacitor c=0.0581858f //x=86.95 \
 //y=0 //x2=86.995 //y2=0.615
cc_987 ( N_GND_c_23_p N_noxref_55_M52_noxref_s ) capacitor c=0.00212661f \
 //x=86.95 //y=0 //x2=84.92 //y2=0.365
cc_988 ( N_GND_c_457_p N_noxref_55_M52_noxref_s ) capacitor c=0.0143168f \
 //x=85.455 //y=0 //x2=84.92 //y2=0.365
cc_989 ( N_GND_c_2_p N_noxref_55_M52_noxref_s ) capacitor c=0.00202267f \
 //x=86.95 //y=0 //x2=84.92 //y2=0.365
cc_990 ( N_GND_c_22_p N_noxref_55_M52_noxref_s ) capacitor c=0.0555228f \
 //x=84.36 //y=0 //x2=84.92 //y2=0.365
cc_991 ( N_GND_M52_noxref_d N_noxref_55_M52_noxref_s ) capacitor c=0.0332904f \
 //x=85.35 //y=0.865 //x2=84.92 //y2=0.365
cc_992 ( N_VDD_c_994_n N_noxref_3_c_2099_n ) capacitor c=6.58823e-19 //x=4.81 \
 //y=7.4 //x2=3.33 //y2=2.08
cc_993 ( N_VDD_c_1015_p N_noxref_3_c_2114_n ) capacitor c=0.00444892f \
 //x=86.95 //y=7.4 //x2=7.135 //y2=5.155
cc_994 ( N_VDD_c_1016_p N_noxref_3_c_2114_n ) capacitor c=4.31931e-19 \
 //x=6.695 //y=7.4 //x2=7.135 //y2=5.155
cc_995 ( N_VDD_c_1017_p N_noxref_3_c_2114_n ) capacitor c=4.31931e-19 \
 //x=7.575 //y=7.4 //x2=7.135 //y2=5.155
cc_996 ( N_VDD_M61_noxref_d N_noxref_3_c_2114_n ) capacitor c=0.0112985f \
 //x=6.635 //y=5.02 //x2=7.135 //y2=5.155
cc_997 ( N_VDD_c_994_n N_noxref_3_c_2118_n ) capacitor c=0.00863585f //x=4.81 \
 //y=7.4 //x2=6.425 //y2=5.155
cc_998 ( N_VDD_M60_noxref_s N_noxref_3_c_2118_n ) capacitor c=0.0831083f \
 //x=5.765 //y=5.02 //x2=6.425 //y2=5.155
cc_999 ( N_VDD_c_1015_p N_noxref_3_c_2120_n ) capacitor c=0.0044221f //x=86.95 \
 //y=7.4 //x2=8.015 //y2=5.155
cc_1000 ( N_VDD_c_1017_p N_noxref_3_c_2120_n ) capacitor c=4.31931e-19 \
 //x=7.575 //y=7.4 //x2=8.015 //y2=5.155
cc_1001 ( N_VDD_c_1023_p N_noxref_3_c_2120_n ) capacitor c=4.31931e-19 \
 //x=8.455 //y=7.4 //x2=8.015 //y2=5.155
cc_1002 ( N_VDD_M63_noxref_d N_noxref_3_c_2120_n ) capacitor c=0.0112985f \
 //x=7.515 //y=5.02 //x2=8.015 //y2=5.155
cc_1003 ( N_VDD_c_1015_p N_noxref_3_c_2124_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=8.795 //y2=5.155
cc_1004 ( N_VDD_c_1023_p N_noxref_3_c_2124_n ) capacitor c=7.46626e-19 \
 //x=8.455 //y=7.4 //x2=8.795 //y2=5.155
cc_1005 ( N_VDD_c_1027_p N_noxref_3_c_2124_n ) capacitor c=0.00198565f \
 //x=9.45 //y=7.4 //x2=8.795 //y2=5.155
cc_1006 ( N_VDD_M65_noxref_d N_noxref_3_c_2124_n ) capacitor c=0.0112985f \
 //x=8.395 //y=5.02 //x2=8.795 //y2=5.155
cc_1007 ( N_VDD_c_995_n N_noxref_3_c_2128_n ) capacitor c=0.0426864f //x=9.62 \
 //y=7.4 //x2=8.88 //y2=3.33
cc_1008 ( N_VDD_c_1015_p N_noxref_3_c_2101_n ) capacitor c=0.00125279f \
 //x=86.95 //y=7.4 //x2=10.73 //y2=2.08
cc_1009 ( N_VDD_c_1031_p N_noxref_3_c_2101_n ) capacitor c=2.87256e-19 \
 //x=11.205 //y=7.4 //x2=10.73 //y2=2.08
cc_1010 ( N_VDD_c_995_n N_noxref_3_c_2101_n ) capacitor c=0.0134208f //x=9.62 \
 //y=7.4 //x2=10.73 //y2=2.08
cc_1011 ( N_VDD_c_1033_p N_noxref_3_M58_noxref_g ) capacitor c=0.00675175f \
 //x=3.645 //y=7.4 //x2=3.07 //y2=6.02
cc_1012 ( N_VDD_M57_noxref_d N_noxref_3_M58_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=3.07 //y2=6.02
cc_1013 ( N_VDD_c_1033_p N_noxref_3_M59_noxref_g ) capacitor c=0.00675379f \
 //x=3.645 //y=7.4 //x2=3.51 //y2=6.02
cc_1014 ( N_VDD_M59_noxref_d N_noxref_3_M59_noxref_g ) capacitor c=0.0394719f \
 //x=3.585 //y=5.02 //x2=3.51 //y2=6.02
cc_1015 ( N_VDD_c_1031_p N_noxref_3_M66_noxref_g ) capacitor c=0.00726866f \
 //x=11.205 //y=7.4 //x2=10.63 //y2=6.02
cc_1016 ( N_VDD_M66_noxref_s N_noxref_3_M66_noxref_g ) capacitor c=0.054195f \
 //x=10.275 //y=5.02 //x2=10.63 //y2=6.02
cc_1017 ( N_VDD_c_1031_p N_noxref_3_M67_noxref_g ) capacitor c=0.00672952f \
 //x=11.205 //y=7.4 //x2=11.07 //y2=6.02
cc_1018 ( N_VDD_M67_noxref_d N_noxref_3_M67_noxref_g ) capacitor c=0.015318f \
 //x=11.145 //y=5.02 //x2=11.07 //y2=6.02
cc_1019 ( N_VDD_c_995_n N_noxref_3_c_2140_n ) capacitor c=0.0154093f //x=9.62 \
 //y=7.4 //x2=10.73 //y2=4.7
cc_1020 ( N_VDD_c_1015_p N_noxref_3_M60_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=6.195 //y2=5.02
cc_1021 ( N_VDD_c_1016_p N_noxref_3_M60_noxref_d ) capacitor c=0.014035f \
 //x=6.695 //y=7.4 //x2=6.195 //y2=5.02
cc_1022 ( N_VDD_M61_noxref_d N_noxref_3_M60_noxref_d ) capacitor c=0.0664752f \
 //x=6.635 //y=5.02 //x2=6.195 //y2=5.02
cc_1023 ( N_VDD_c_1015_p N_noxref_3_M62_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=7.075 //y2=5.02
cc_1024 ( N_VDD_c_1017_p N_noxref_3_M62_noxref_d ) capacitor c=0.014035f \
 //x=7.575 //y=7.4 //x2=7.075 //y2=5.02
cc_1025 ( N_VDD_c_995_n N_noxref_3_M62_noxref_d ) capacitor c=4.9285e-19 \
 //x=9.62 //y=7.4 //x2=7.075 //y2=5.02
cc_1026 ( N_VDD_M60_noxref_s N_noxref_3_M62_noxref_d ) capacitor c=0.00130656f \
 //x=5.765 //y=5.02 //x2=7.075 //y2=5.02
cc_1027 ( N_VDD_M61_noxref_d N_noxref_3_M62_noxref_d ) capacitor c=0.0664752f \
 //x=6.635 //y=5.02 //x2=7.075 //y2=5.02
cc_1028 ( N_VDD_M63_noxref_d N_noxref_3_M62_noxref_d ) capacitor c=0.0664752f \
 //x=7.515 //y=5.02 //x2=7.075 //y2=5.02
cc_1029 ( N_VDD_c_1015_p N_noxref_3_M64_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=7.955 //y2=5.02
cc_1030 ( N_VDD_c_1023_p N_noxref_3_M64_noxref_d ) capacitor c=0.014035f \
 //x=8.455 //y=7.4 //x2=7.955 //y2=5.02
cc_1031 ( N_VDD_c_995_n N_noxref_3_M64_noxref_d ) capacitor c=0.00939849f \
 //x=9.62 //y=7.4 //x2=7.955 //y2=5.02
cc_1032 ( N_VDD_M63_noxref_d N_noxref_3_M64_noxref_d ) capacitor c=0.0664752f \
 //x=7.515 //y=5.02 //x2=7.955 //y2=5.02
cc_1033 ( N_VDD_M65_noxref_d N_noxref_3_M64_noxref_d ) capacitor c=0.0664752f \
 //x=8.395 //y=5.02 //x2=7.955 //y2=5.02
cc_1034 ( N_VDD_M66_noxref_s N_noxref_3_M64_noxref_d ) capacitor c=4.52683e-19 \
 //x=10.275 //y=5.02 //x2=7.955 //y2=5.02
cc_1035 ( N_VDD_c_1015_p N_noxref_4_c_2360_n ) capacitor c=0.00453663f \
 //x=86.95 //y=7.4 //x2=11.645 //y2=5.2
cc_1036 ( N_VDD_c_1031_p N_noxref_4_c_2360_n ) capacitor c=4.48391e-19 \
 //x=11.205 //y=7.4 //x2=11.645 //y2=5.2
cc_1037 ( N_VDD_c_1059_p N_noxref_4_c_2360_n ) capacitor c=4.48391e-19 \
 //x=12.085 //y=7.4 //x2=11.645 //y2=5.2
cc_1038 ( N_VDD_M67_noxref_d N_noxref_4_c_2360_n ) capacitor c=0.0124542f \
 //x=11.145 //y=5.02 //x2=11.645 //y2=5.2
cc_1039 ( N_VDD_c_995_n N_noxref_4_c_2364_n ) capacitor c=0.00985474f //x=9.62 \
 //y=7.4 //x2=10.935 //y2=5.2
cc_1040 ( N_VDD_M66_noxref_s N_noxref_4_c_2364_n ) capacitor c=0.087833f \
 //x=10.275 //y=5.02 //x2=10.935 //y2=5.2
cc_1041 ( N_VDD_c_1015_p N_noxref_4_c_2366_n ) capacitor c=0.00301575f \
 //x=86.95 //y=7.4 //x2=12.125 //y2=5.2
cc_1042 ( N_VDD_c_1059_p N_noxref_4_c_2366_n ) capacitor c=7.72068e-19 \
 //x=12.085 //y=7.4 //x2=12.125 //y2=5.2
cc_1043 ( N_VDD_M69_noxref_d N_noxref_4_c_2366_n ) capacitor c=0.0158515f \
 //x=12.025 //y=5.02 //x2=12.125 //y2=5.2
cc_1044 ( N_VDD_c_995_n N_noxref_4_c_2345_n ) capacitor c=0.00151618f //x=9.62 \
 //y=7.4 //x2=12.21 //y2=3.33
cc_1045 ( N_VDD_c_996_n N_noxref_4_c_2345_n ) capacitor c=0.0428942f //x=12.95 \
 //y=7.4 //x2=12.21 //y2=3.33
cc_1046 ( N_VDD_c_1015_p N_noxref_4_c_2346_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=14.06 //y2=2.08
cc_1047 ( N_VDD_c_996_n N_noxref_4_c_2346_n ) capacitor c=0.0133749f //x=12.95 \
 //y=7.4 //x2=14.06 //y2=2.08
cc_1048 ( N_VDD_M70_noxref_s N_noxref_4_c_2346_n ) capacitor c=0.0125322f \
 //x=13.905 //y=5.02 //x2=14.06 //y2=2.08
cc_1049 ( N_VDD_c_1071_p N_noxref_4_M70_noxref_g ) capacitor c=0.00749687f \
 //x=14.835 //y=7.4 //x2=14.26 //y2=6.02
cc_1050 ( N_VDD_M70_noxref_s N_noxref_4_M70_noxref_g ) capacitor c=0.0477201f \
 //x=13.905 //y=5.02 //x2=14.26 //y2=6.02
cc_1051 ( N_VDD_c_1071_p N_noxref_4_M71_noxref_g ) capacitor c=0.00675175f \
 //x=14.835 //y=7.4 //x2=14.7 //y2=6.02
cc_1052 ( N_VDD_M71_noxref_d N_noxref_4_M71_noxref_g ) capacitor c=0.015318f \
 //x=14.775 //y=5.02 //x2=14.7 //y2=6.02
cc_1053 ( N_VDD_c_996_n N_noxref_4_c_2378_n ) capacitor c=0.00757682f \
 //x=12.95 //y=7.4 //x2=14.335 //y2=4.79
cc_1054 ( N_VDD_M70_noxref_s N_noxref_4_c_2378_n ) capacitor c=0.00444914f \
 //x=13.905 //y=5.02 //x2=14.335 //y2=4.79
cc_1055 ( N_VDD_c_1015_p N_noxref_4_M66_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=10.705 //y2=5.02
cc_1056 ( N_VDD_c_1031_p N_noxref_4_M66_noxref_d ) capacitor c=0.0140317f \
 //x=11.205 //y=7.4 //x2=10.705 //y2=5.02
cc_1057 ( N_VDD_c_996_n N_noxref_4_M66_noxref_d ) capacitor c=6.94454e-19 \
 //x=12.95 //y=7.4 //x2=10.705 //y2=5.02
cc_1058 ( N_VDD_M67_noxref_d N_noxref_4_M66_noxref_d ) capacitor c=0.0664752f \
 //x=11.145 //y=5.02 //x2=10.705 //y2=5.02
cc_1059 ( N_VDD_c_1015_p N_noxref_4_M68_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=11.585 //y2=5.02
cc_1060 ( N_VDD_c_1059_p N_noxref_4_M68_noxref_d ) capacitor c=0.0140317f \
 //x=12.085 //y=7.4 //x2=11.585 //y2=5.02
cc_1061 ( N_VDD_c_996_n N_noxref_4_M68_noxref_d ) capacitor c=0.0120541f \
 //x=12.95 //y=7.4 //x2=11.585 //y2=5.02
cc_1062 ( N_VDD_M66_noxref_s N_noxref_4_M68_noxref_d ) capacitor c=0.00111971f \
 //x=10.275 //y=5.02 //x2=11.585 //y2=5.02
cc_1063 ( N_VDD_M67_noxref_d N_noxref_4_M68_noxref_d ) capacitor c=0.0664752f \
 //x=11.145 //y=5.02 //x2=11.585 //y2=5.02
cc_1064 ( N_VDD_M69_noxref_d N_noxref_4_M68_noxref_d ) capacitor c=0.0664752f \
 //x=12.025 //y=5.02 //x2=11.585 //y2=5.02
cc_1065 ( N_VDD_M70_noxref_s N_noxref_4_M68_noxref_d ) capacitor c=3.73257e-19 \
 //x=13.905 //y=5.02 //x2=11.585 //y2=5.02
cc_1066 ( N_VDD_c_1015_p N_noxref_5_c_2520_n ) capacitor c=0.00449316f \
 //x=86.95 //y=7.4 //x2=2.325 //y2=5.155
cc_1067 ( N_VDD_c_1089_p N_noxref_5_c_2520_n ) capacitor c=4.32228e-19 \
 //x=1.885 //y=7.4 //x2=2.325 //y2=5.155
cc_1068 ( N_VDD_c_1090_p N_noxref_5_c_2520_n ) capacitor c=4.31906e-19 \
 //x=2.765 //y=7.4 //x2=2.325 //y2=5.155
cc_1069 ( N_VDD_M55_noxref_d N_noxref_5_c_2520_n ) capacitor c=0.0115147f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_1070 ( N_VDD_c_992_n N_noxref_5_c_2524_n ) capacitor c=0.00880189f //x=0.74 \
 //y=7.4 //x2=1.615 //y2=5.155
cc_1071 ( N_VDD_M54_noxref_s N_noxref_5_c_2524_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_1072 ( N_VDD_c_1015_p N_noxref_5_c_2526_n ) capacitor c=0.0044221f \
 //x=86.95 //y=7.4 //x2=3.205 //y2=5.155
cc_1073 ( N_VDD_c_1090_p N_noxref_5_c_2526_n ) capacitor c=4.31931e-19 \
 //x=2.765 //y=7.4 //x2=3.205 //y2=5.155
cc_1074 ( N_VDD_c_1033_p N_noxref_5_c_2526_n ) capacitor c=4.31931e-19 \
 //x=3.645 //y=7.4 //x2=3.205 //y2=5.155
cc_1075 ( N_VDD_M57_noxref_d N_noxref_5_c_2526_n ) capacitor c=0.0112985f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_1076 ( N_VDD_c_1015_p N_noxref_5_c_2530_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=3.985 //y2=5.155
cc_1077 ( N_VDD_c_1033_p N_noxref_5_c_2530_n ) capacitor c=7.46626e-19 \
 //x=3.645 //y=7.4 //x2=3.985 //y2=5.155
cc_1078 ( N_VDD_c_1100_p N_noxref_5_c_2530_n ) capacitor c=0.00198565f \
 //x=4.64 //y=7.4 //x2=3.985 //y2=5.155
cc_1079 ( N_VDD_M59_noxref_d N_noxref_5_c_2530_n ) capacitor c=0.0112985f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_1080 ( N_VDD_c_994_n N_noxref_5_c_2534_n ) capacitor c=0.0427116f //x=4.81 \
 //y=7.4 //x2=4.07 //y2=3.7
cc_1081 ( N_VDD_c_1015_p N_noxref_5_c_2497_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=5.92 //y2=2.08
cc_1082 ( N_VDD_c_994_n N_noxref_5_c_2497_n ) capacitor c=0.0134711f //x=4.81 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_1083 ( N_VDD_M60_noxref_s N_noxref_5_c_2497_n ) capacitor c=0.0120327f \
 //x=5.765 //y=5.02 //x2=5.92 //y2=2.08
cc_1084 ( N_VDD_c_1015_p N_noxref_5_c_2498_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=18.87 //y2=2.08
cc_1085 ( N_VDD_c_997_n N_noxref_5_c_2498_n ) capacitor c=0.0134269f //x=17.76 \
 //y=7.4 //x2=18.87 //y2=2.08
cc_1086 ( N_VDD_M76_noxref_s N_noxref_5_c_2498_n ) capacitor c=0.0125322f \
 //x=18.715 //y=5.02 //x2=18.87 //y2=2.08
cc_1087 ( N_VDD_c_1016_p N_noxref_5_M60_noxref_g ) capacitor c=0.00749687f \
 //x=6.695 //y=7.4 //x2=6.12 //y2=6.02
cc_1088 ( N_VDD_M60_noxref_s N_noxref_5_M60_noxref_g ) capacitor c=0.0477201f \
 //x=5.765 //y=5.02 //x2=6.12 //y2=6.02
cc_1089 ( N_VDD_c_1016_p N_noxref_5_M61_noxref_g ) capacitor c=0.00675175f \
 //x=6.695 //y=7.4 //x2=6.56 //y2=6.02
cc_1090 ( N_VDD_M61_noxref_d N_noxref_5_M61_noxref_g ) capacitor c=0.015318f \
 //x=6.635 //y=5.02 //x2=6.56 //y2=6.02
cc_1091 ( N_VDD_c_1113_p N_noxref_5_M76_noxref_g ) capacitor c=0.00749687f \
 //x=19.645 //y=7.4 //x2=19.07 //y2=6.02
cc_1092 ( N_VDD_M76_noxref_s N_noxref_5_M76_noxref_g ) capacitor c=0.0477201f \
 //x=18.715 //y=5.02 //x2=19.07 //y2=6.02
cc_1093 ( N_VDD_c_1113_p N_noxref_5_M77_noxref_g ) capacitor c=0.00675175f \
 //x=19.645 //y=7.4 //x2=19.51 //y2=6.02
cc_1094 ( N_VDD_M77_noxref_d N_noxref_5_M77_noxref_g ) capacitor c=0.015318f \
 //x=19.585 //y=5.02 //x2=19.51 //y2=6.02
cc_1095 ( N_VDD_c_994_n N_noxref_5_c_2549_n ) capacitor c=0.00757682f //x=4.81 \
 //y=7.4 //x2=6.195 //y2=4.79
cc_1096 ( N_VDD_M60_noxref_s N_noxref_5_c_2549_n ) capacitor c=0.00444914f \
 //x=5.765 //y=5.02 //x2=6.195 //y2=4.79
cc_1097 ( N_VDD_c_997_n N_noxref_5_c_2551_n ) capacitor c=0.00757682f \
 //x=17.76 //y=7.4 //x2=19.145 //y2=4.79
cc_1098 ( N_VDD_M76_noxref_s N_noxref_5_c_2551_n ) capacitor c=0.00444914f \
 //x=18.715 //y=5.02 //x2=19.145 //y2=4.79
cc_1099 ( N_VDD_c_1015_p N_noxref_5_M54_noxref_d ) capacitor c=0.00285091f \
 //x=86.95 //y=7.4 //x2=1.385 //y2=5.02
cc_1100 ( N_VDD_c_1089_p N_noxref_5_M54_noxref_d ) capacitor c=0.0141016f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_1101 ( N_VDD_M55_noxref_d N_noxref_5_M54_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_1102 ( N_VDD_c_1015_p N_noxref_5_M56_noxref_d ) capacitor c=0.00275186f \
 //x=86.95 //y=7.4 //x2=2.265 //y2=5.02
cc_1103 ( N_VDD_c_1090_p N_noxref_5_M56_noxref_d ) capacitor c=0.0140346f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_1104 ( N_VDD_c_994_n N_noxref_5_M56_noxref_d ) capacitor c=4.9285e-19 \
 //x=4.81 //y=7.4 //x2=2.265 //y2=5.02
cc_1105 ( N_VDD_M54_noxref_s N_noxref_5_M56_noxref_d ) capacitor c=0.00130656f \
 //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_1106 ( N_VDD_M55_noxref_d N_noxref_5_M56_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_1107 ( N_VDD_M57_noxref_d N_noxref_5_M56_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_1108 ( N_VDD_c_1015_p N_noxref_5_M58_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=3.145 //y2=5.02
cc_1109 ( N_VDD_c_1033_p N_noxref_5_M58_noxref_d ) capacitor c=0.0137384f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_1110 ( N_VDD_c_994_n N_noxref_5_M58_noxref_d ) capacitor c=0.00939849f \
 //x=4.81 //y=7.4 //x2=3.145 //y2=5.02
cc_1111 ( N_VDD_M57_noxref_d N_noxref_5_M58_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_1112 ( N_VDD_M59_noxref_d N_noxref_5_M58_noxref_d ) capacitor c=0.0664752f \
 //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_1113 ( N_VDD_M60_noxref_s N_noxref_5_M58_noxref_d ) capacitor c=3.57641e-19 \
 //x=5.765 //y=5.02 //x2=3.145 //y2=5.02
cc_1114 ( N_VDD_c_1015_p N_noxref_6_c_2748_n ) capacitor c=0.0425735f \
 //x=86.95 //y=7.4 //x2=11.355 //y2=4.07
cc_1115 ( N_VDD_c_1089_p N_noxref_6_c_2748_n ) capacitor c=0.00113322f \
 //x=1.885 //y=7.4 //x2=11.355 //y2=4.07
cc_1116 ( N_VDD_c_994_n N_noxref_6_c_2748_n ) capacitor c=0.0140578f //x=4.81 \
 //y=7.4 //x2=11.355 //y2=4.07
cc_1117 ( N_VDD_c_995_n N_noxref_6_c_2748_n ) capacitor c=0.0140578f //x=9.62 \
 //y=7.4 //x2=11.355 //y2=4.07
cc_1118 ( N_VDD_c_1015_p N_noxref_6_c_2749_n ) capacitor c=0.00189266f \
 //x=86.95 //y=7.4 //x2=1.225 //y2=4.07
cc_1119 ( N_VDD_c_992_n N_noxref_6_c_2749_n ) capacitor c=0.0017219f //x=0.74 \
 //y=7.4 //x2=1.225 //y2=4.07
cc_1120 ( N_VDD_M54_noxref_s N_noxref_6_c_2749_n ) capacitor c=0.00128242f \
 //x=0.955 //y=5.02 //x2=1.225 //y2=4.07
cc_1121 ( N_VDD_c_996_n N_noxref_6_c_2787_n ) capacitor c=0.0140578f //x=12.95 \
 //y=7.4 //x2=16.905 //y2=4.07
cc_1122 ( N_VDD_c_997_n N_noxref_6_c_2788_n ) capacitor c=0.0140578f //x=17.76 \
 //y=7.4 //x2=21.715 //y2=4.07
cc_1123 ( N_VDD_c_997_n N_noxref_6_c_2789_n ) capacitor c=0.00104972f \
 //x=17.76 //y=7.4 //x2=17.135 //y2=4.07
cc_1124 ( N_VDD_c_998_n N_noxref_6_c_2790_n ) capacitor c=0.0145592f //x=22.57 \
 //y=7.4 //x2=23.565 //y2=4.07
cc_1125 ( N_VDD_c_998_n N_noxref_6_c_2791_n ) capacitor c=5.12647e-19 \
 //x=22.57 //y=7.4 //x2=21.945 //y2=4.07
cc_1126 ( N_VDD_c_998_n N_noxref_6_c_2792_n ) capacitor c=3.58282e-19 \
 //x=22.57 //y=7.4 //x2=23.795 //y2=4.07
cc_1127 ( N_VDD_c_1015_p N_noxref_6_c_2750_n ) capacitor c=9.2251e-19 \
 //x=86.95 //y=7.4 //x2=1.11 //y2=2.08
cc_1128 ( N_VDD_c_992_n N_noxref_6_c_2750_n ) capacitor c=0.0159723f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_1129 ( N_VDD_M54_noxref_s N_noxref_6_c_2750_n ) capacitor c=0.0122951f \
 //x=0.955 //y=5.02 //x2=1.11 //y2=2.08
cc_1130 ( N_VDD_c_995_n N_noxref_6_c_2751_n ) capacitor c=4.57806e-19 //x=9.62 \
 //y=7.4 //x2=11.47 //y2=2.08
cc_1131 ( N_VDD_c_996_n N_noxref_6_c_2751_n ) capacitor c=3.21957e-19 \
 //x=12.95 //y=7.4 //x2=11.47 //y2=2.08
cc_1132 ( N_VDD_c_1015_p N_noxref_6_c_2798_n ) capacitor c=0.00444751f \
 //x=86.95 //y=7.4 //x2=15.275 //y2=5.155
cc_1133 ( N_VDD_c_1071_p N_noxref_6_c_2798_n ) capacitor c=4.31931e-19 \
 //x=14.835 //y=7.4 //x2=15.275 //y2=5.155
cc_1134 ( N_VDD_c_1156_p N_noxref_6_c_2798_n ) capacitor c=4.31906e-19 \
 //x=15.715 //y=7.4 //x2=15.275 //y2=5.155
cc_1135 ( N_VDD_M71_noxref_d N_noxref_6_c_2798_n ) capacitor c=0.0112985f \
 //x=14.775 //y=5.02 //x2=15.275 //y2=5.155
cc_1136 ( N_VDD_c_996_n N_noxref_6_c_2802_n ) capacitor c=0.00863585f \
 //x=12.95 //y=7.4 //x2=14.565 //y2=5.155
cc_1137 ( N_VDD_M70_noxref_s N_noxref_6_c_2802_n ) capacitor c=0.0831083f \
 //x=13.905 //y=5.02 //x2=14.565 //y2=5.155
cc_1138 ( N_VDD_c_1015_p N_noxref_6_c_2804_n ) capacitor c=0.0044221f \
 //x=86.95 //y=7.4 //x2=16.155 //y2=5.155
cc_1139 ( N_VDD_c_1156_p N_noxref_6_c_2804_n ) capacitor c=4.31931e-19 \
 //x=15.715 //y=7.4 //x2=16.155 //y2=5.155
cc_1140 ( N_VDD_c_1162_p N_noxref_6_c_2804_n ) capacitor c=4.31931e-19 \
 //x=16.595 //y=7.4 //x2=16.155 //y2=5.155
cc_1141 ( N_VDD_M73_noxref_d N_noxref_6_c_2804_n ) capacitor c=0.0112985f \
 //x=15.655 //y=5.02 //x2=16.155 //y2=5.155
cc_1142 ( N_VDD_c_1015_p N_noxref_6_c_2808_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=16.935 //y2=5.155
cc_1143 ( N_VDD_c_1162_p N_noxref_6_c_2808_n ) capacitor c=7.46626e-19 \
 //x=16.595 //y=7.4 //x2=16.935 //y2=5.155
cc_1144 ( N_VDD_c_1166_p N_noxref_6_c_2808_n ) capacitor c=0.00198565f \
 //x=17.59 //y=7.4 //x2=16.935 //y2=5.155
cc_1145 ( N_VDD_M75_noxref_d N_noxref_6_c_2808_n ) capacitor c=0.0112985f \
 //x=16.535 //y=5.02 //x2=16.935 //y2=5.155
cc_1146 ( N_VDD_c_997_n N_noxref_6_c_2812_n ) capacitor c=0.0429118f //x=17.76 \
 //y=7.4 //x2=17.02 //y2=4.07
cc_1147 ( N_VDD_c_1015_p N_noxref_6_c_2813_n ) capacitor c=0.00444892f \
 //x=86.95 //y=7.4 //x2=20.085 //y2=5.155
cc_1148 ( N_VDD_c_1113_p N_noxref_6_c_2813_n ) capacitor c=4.31931e-19 \
 //x=19.645 //y=7.4 //x2=20.085 //y2=5.155
cc_1149 ( N_VDD_c_1171_p N_noxref_6_c_2813_n ) capacitor c=4.31931e-19 \
 //x=20.525 //y=7.4 //x2=20.085 //y2=5.155
cc_1150 ( N_VDD_M77_noxref_d N_noxref_6_c_2813_n ) capacitor c=0.0112985f \
 //x=19.585 //y=5.02 //x2=20.085 //y2=5.155
cc_1151 ( N_VDD_c_997_n N_noxref_6_c_2817_n ) capacitor c=0.00863585f \
 //x=17.76 //y=7.4 //x2=19.375 //y2=5.155
cc_1152 ( N_VDD_M76_noxref_s N_noxref_6_c_2817_n ) capacitor c=0.0831083f \
 //x=18.715 //y=5.02 //x2=19.375 //y2=5.155
cc_1153 ( N_VDD_c_1015_p N_noxref_6_c_2819_n ) capacitor c=0.0044221f \
 //x=86.95 //y=7.4 //x2=20.965 //y2=5.155
cc_1154 ( N_VDD_c_1171_p N_noxref_6_c_2819_n ) capacitor c=4.31931e-19 \
 //x=20.525 //y=7.4 //x2=20.965 //y2=5.155
cc_1155 ( N_VDD_c_1177_p N_noxref_6_c_2819_n ) capacitor c=4.31931e-19 \
 //x=21.405 //y=7.4 //x2=20.965 //y2=5.155
cc_1156 ( N_VDD_M79_noxref_d N_noxref_6_c_2819_n ) capacitor c=0.0112985f \
 //x=20.465 //y=5.02 //x2=20.965 //y2=5.155
cc_1157 ( N_VDD_c_1015_p N_noxref_6_c_2823_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=21.745 //y2=5.155
cc_1158 ( N_VDD_c_1177_p N_noxref_6_c_2823_n ) capacitor c=7.46626e-19 \
 //x=21.405 //y=7.4 //x2=21.745 //y2=5.155
cc_1159 ( N_VDD_c_1181_p N_noxref_6_c_2823_n ) capacitor c=0.00198565f \
 //x=22.4 //y=7.4 //x2=21.745 //y2=5.155
cc_1160 ( N_VDD_M81_noxref_d N_noxref_6_c_2823_n ) capacitor c=0.0112985f \
 //x=21.345 //y=5.02 //x2=21.745 //y2=5.155
cc_1161 ( N_VDD_c_998_n N_noxref_6_c_2827_n ) capacitor c=0.0430224f //x=22.57 \
 //y=7.4 //x2=21.83 //y2=4.07
cc_1162 ( N_VDD_c_1015_p N_noxref_6_c_2755_n ) capacitor c=0.00125279f \
 //x=86.95 //y=7.4 //x2=23.68 //y2=2.08
cc_1163 ( N_VDD_c_1185_p N_noxref_6_c_2755_n ) capacitor c=2.87256e-19 \
 //x=24.155 //y=7.4 //x2=23.68 //y2=2.08
cc_1164 ( N_VDD_c_998_n N_noxref_6_c_2755_n ) capacitor c=0.0134064f //x=22.57 \
 //y=7.4 //x2=23.68 //y2=2.08
cc_1165 ( N_VDD_c_998_n N_noxref_6_c_2756_n ) capacitor c=4.5519e-19 //x=22.57 \
 //y=7.4 //x2=24.42 //y2=2.08
cc_1166 ( N_VDD_c_999_n N_noxref_6_c_2756_n ) capacitor c=4.17938e-19 //x=25.9 \
 //y=7.4 //x2=24.42 //y2=2.08
cc_1167 ( N_VDD_c_1089_p N_noxref_6_M54_noxref_g ) capacitor c=0.00749687f \
 //x=1.885 //y=7.4 //x2=1.31 //y2=6.02
cc_1168 ( N_VDD_M54_noxref_s N_noxref_6_M54_noxref_g ) capacitor c=0.0477201f \
 //x=0.955 //y=5.02 //x2=1.31 //y2=6.02
cc_1169 ( N_VDD_c_1089_p N_noxref_6_M55_noxref_g ) capacitor c=0.00675175f \
 //x=1.885 //y=7.4 //x2=1.75 //y2=6.02
cc_1170 ( N_VDD_M55_noxref_d N_noxref_6_M55_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=1.75 //y2=6.02
cc_1171 ( N_VDD_c_1059_p N_noxref_6_M68_noxref_g ) capacitor c=0.00673971f \
 //x=12.085 //y=7.4 //x2=11.51 //y2=6.02
cc_1172 ( N_VDD_M67_noxref_d N_noxref_6_M68_noxref_g ) capacitor c=0.015318f \
 //x=11.145 //y=5.02 //x2=11.51 //y2=6.02
cc_1173 ( N_VDD_c_1059_p N_noxref_6_M69_noxref_g ) capacitor c=0.00672952f \
 //x=12.085 //y=7.4 //x2=11.95 //y2=6.02
cc_1174 ( N_VDD_c_996_n N_noxref_6_M69_noxref_g ) capacitor c=0.00928743f \
 //x=12.95 //y=7.4 //x2=11.95 //y2=6.02
cc_1175 ( N_VDD_M69_noxref_d N_noxref_6_M69_noxref_g ) capacitor c=0.0430452f \
 //x=12.025 //y=5.02 //x2=11.95 //y2=6.02
cc_1176 ( N_VDD_c_1185_p N_noxref_6_M82_noxref_g ) capacitor c=0.00726866f \
 //x=24.155 //y=7.4 //x2=23.58 //y2=6.02
cc_1177 ( N_VDD_M82_noxref_s N_noxref_6_M82_noxref_g ) capacitor c=0.054195f \
 //x=23.225 //y=5.02 //x2=23.58 //y2=6.02
cc_1178 ( N_VDD_c_1185_p N_noxref_6_M83_noxref_g ) capacitor c=0.00672952f \
 //x=24.155 //y=7.4 //x2=24.02 //y2=6.02
cc_1179 ( N_VDD_M83_noxref_d N_noxref_6_M83_noxref_g ) capacitor c=0.015318f \
 //x=24.095 //y=5.02 //x2=24.02 //y2=6.02
cc_1180 ( N_VDD_c_1202_p N_noxref_6_M84_noxref_g ) capacitor c=0.00673971f \
 //x=25.035 //y=7.4 //x2=24.46 //y2=6.02
cc_1181 ( N_VDD_M83_noxref_d N_noxref_6_M84_noxref_g ) capacitor c=0.015318f \
 //x=24.095 //y=5.02 //x2=24.46 //y2=6.02
cc_1182 ( N_VDD_c_1202_p N_noxref_6_M85_noxref_g ) capacitor c=0.00672952f \
 //x=25.035 //y=7.4 //x2=24.9 //y2=6.02
cc_1183 ( N_VDD_c_999_n N_noxref_6_M85_noxref_g ) capacitor c=0.00928743f \
 //x=25.9 //y=7.4 //x2=24.9 //y2=6.02
cc_1184 ( N_VDD_M85_noxref_d N_noxref_6_M85_noxref_g ) capacitor c=0.0430452f \
 //x=24.975 //y=5.02 //x2=24.9 //y2=6.02
cc_1185 ( N_VDD_c_992_n N_noxref_6_c_2851_n ) capacitor c=0.00757682f //x=0.74 \
 //y=7.4 //x2=1.385 //y2=4.79
cc_1186 ( N_VDD_M54_noxref_s N_noxref_6_c_2851_n ) capacitor c=0.00445117f \
 //x=0.955 //y=5.02 //x2=1.385 //y2=4.79
cc_1187 ( N_VDD_c_998_n N_noxref_6_c_2853_n ) capacitor c=0.0154093f //x=22.57 \
 //y=7.4 //x2=23.68 //y2=4.7
cc_1188 ( N_VDD_c_1015_p N_noxref_6_M70_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=14.335 //y2=5.02
cc_1189 ( N_VDD_c_1071_p N_noxref_6_M70_noxref_d ) capacitor c=0.014035f \
 //x=14.835 //y=7.4 //x2=14.335 //y2=5.02
cc_1190 ( N_VDD_M71_noxref_d N_noxref_6_M70_noxref_d ) capacitor c=0.0664752f \
 //x=14.775 //y=5.02 //x2=14.335 //y2=5.02
cc_1191 ( N_VDD_c_1015_p N_noxref_6_M72_noxref_d ) capacitor c=0.00275186f \
 //x=86.95 //y=7.4 //x2=15.215 //y2=5.02
cc_1192 ( N_VDD_c_1156_p N_noxref_6_M72_noxref_d ) capacitor c=0.0140346f \
 //x=15.715 //y=7.4 //x2=15.215 //y2=5.02
cc_1193 ( N_VDD_c_997_n N_noxref_6_M72_noxref_d ) capacitor c=4.9285e-19 \
 //x=17.76 //y=7.4 //x2=15.215 //y2=5.02
cc_1194 ( N_VDD_M70_noxref_s N_noxref_6_M72_noxref_d ) capacitor c=0.00130656f \
 //x=13.905 //y=5.02 //x2=15.215 //y2=5.02
cc_1195 ( N_VDD_M71_noxref_d N_noxref_6_M72_noxref_d ) capacitor c=0.0664752f \
 //x=14.775 //y=5.02 //x2=15.215 //y2=5.02
cc_1196 ( N_VDD_M73_noxref_d N_noxref_6_M72_noxref_d ) capacitor c=0.0664752f \
 //x=15.655 //y=5.02 //x2=15.215 //y2=5.02
cc_1197 ( N_VDD_c_1015_p N_noxref_6_M74_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=16.095 //y2=5.02
cc_1198 ( N_VDD_c_1162_p N_noxref_6_M74_noxref_d ) capacitor c=0.014035f \
 //x=16.595 //y=7.4 //x2=16.095 //y2=5.02
cc_1199 ( N_VDD_c_997_n N_noxref_6_M74_noxref_d ) capacitor c=0.00939849f \
 //x=17.76 //y=7.4 //x2=16.095 //y2=5.02
cc_1200 ( N_VDD_M73_noxref_d N_noxref_6_M74_noxref_d ) capacitor c=0.0664752f \
 //x=15.655 //y=5.02 //x2=16.095 //y2=5.02
cc_1201 ( N_VDD_M75_noxref_d N_noxref_6_M74_noxref_d ) capacitor c=0.0664752f \
 //x=16.535 //y=5.02 //x2=16.095 //y2=5.02
cc_1202 ( N_VDD_M76_noxref_s N_noxref_6_M74_noxref_d ) capacitor c=3.57641e-19 \
 //x=18.715 //y=5.02 //x2=16.095 //y2=5.02
cc_1203 ( N_VDD_c_1015_p N_noxref_6_M76_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=19.145 //y2=5.02
cc_1204 ( N_VDD_c_1113_p N_noxref_6_M76_noxref_d ) capacitor c=0.014035f \
 //x=19.645 //y=7.4 //x2=19.145 //y2=5.02
cc_1205 ( N_VDD_M77_noxref_d N_noxref_6_M76_noxref_d ) capacitor c=0.0664752f \
 //x=19.585 //y=5.02 //x2=19.145 //y2=5.02
cc_1206 ( N_VDD_c_1015_p N_noxref_6_M78_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=20.025 //y2=5.02
cc_1207 ( N_VDD_c_1171_p N_noxref_6_M78_noxref_d ) capacitor c=0.014035f \
 //x=20.525 //y=7.4 //x2=20.025 //y2=5.02
cc_1208 ( N_VDD_c_998_n N_noxref_6_M78_noxref_d ) capacitor c=4.9285e-19 \
 //x=22.57 //y=7.4 //x2=20.025 //y2=5.02
cc_1209 ( N_VDD_M76_noxref_s N_noxref_6_M78_noxref_d ) capacitor c=0.00130656f \
 //x=18.715 //y=5.02 //x2=20.025 //y2=5.02
cc_1210 ( N_VDD_M77_noxref_d N_noxref_6_M78_noxref_d ) capacitor c=0.0664752f \
 //x=19.585 //y=5.02 //x2=20.025 //y2=5.02
cc_1211 ( N_VDD_M79_noxref_d N_noxref_6_M78_noxref_d ) capacitor c=0.0664752f \
 //x=20.465 //y=5.02 //x2=20.025 //y2=5.02
cc_1212 ( N_VDD_c_1015_p N_noxref_6_M80_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=20.905 //y2=5.02
cc_1213 ( N_VDD_c_1177_p N_noxref_6_M80_noxref_d ) capacitor c=0.0137384f \
 //x=21.405 //y=7.4 //x2=20.905 //y2=5.02
cc_1214 ( N_VDD_c_998_n N_noxref_6_M80_noxref_d ) capacitor c=0.00939849f \
 //x=22.57 //y=7.4 //x2=20.905 //y2=5.02
cc_1215 ( N_VDD_M79_noxref_d N_noxref_6_M80_noxref_d ) capacitor c=0.0664752f \
 //x=20.465 //y=5.02 //x2=20.905 //y2=5.02
cc_1216 ( N_VDD_M81_noxref_d N_noxref_6_M80_noxref_d ) capacitor c=0.0664752f \
 //x=21.345 //y=5.02 //x2=20.905 //y2=5.02
cc_1217 ( N_VDD_M82_noxref_s N_noxref_6_M80_noxref_d ) capacitor c=4.52683e-19 \
 //x=23.225 //y=5.02 //x2=20.905 //y2=5.02
cc_1218 ( N_VDD_c_1000_n N_noxref_7_c_3233_n ) capacitor c=6.58823e-19 \
 //x=30.71 //y=7.4 //x2=29.23 //y2=2.08
cc_1219 ( N_VDD_c_1015_p N_noxref_7_c_3248_n ) capacitor c=0.00444892f \
 //x=86.95 //y=7.4 //x2=33.035 //y2=5.155
cc_1220 ( N_VDD_c_1242_p N_noxref_7_c_3248_n ) capacitor c=4.31931e-19 \
 //x=32.595 //y=7.4 //x2=33.035 //y2=5.155
cc_1221 ( N_VDD_c_1243_p N_noxref_7_c_3248_n ) capacitor c=4.31931e-19 \
 //x=33.475 //y=7.4 //x2=33.035 //y2=5.155
cc_1222 ( N_VDD_M93_noxref_d N_noxref_7_c_3248_n ) capacitor c=0.0112985f \
 //x=32.535 //y=5.02 //x2=33.035 //y2=5.155
cc_1223 ( N_VDD_c_1000_n N_noxref_7_c_3252_n ) capacitor c=0.00863585f \
 //x=30.71 //y=7.4 //x2=32.325 //y2=5.155
cc_1224 ( N_VDD_M92_noxref_s N_noxref_7_c_3252_n ) capacitor c=0.0831083f \
 //x=31.665 //y=5.02 //x2=32.325 //y2=5.155
cc_1225 ( N_VDD_c_1015_p N_noxref_7_c_3254_n ) capacitor c=0.0044221f \
 //x=86.95 //y=7.4 //x2=33.915 //y2=5.155
cc_1226 ( N_VDD_c_1243_p N_noxref_7_c_3254_n ) capacitor c=4.31931e-19 \
 //x=33.475 //y=7.4 //x2=33.915 //y2=5.155
cc_1227 ( N_VDD_c_1249_p N_noxref_7_c_3254_n ) capacitor c=4.31931e-19 \
 //x=34.355 //y=7.4 //x2=33.915 //y2=5.155
cc_1228 ( N_VDD_M95_noxref_d N_noxref_7_c_3254_n ) capacitor c=0.0112985f \
 //x=33.415 //y=5.02 //x2=33.915 //y2=5.155
cc_1229 ( N_VDD_c_1015_p N_noxref_7_c_3258_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=34.695 //y2=5.155
cc_1230 ( N_VDD_c_1249_p N_noxref_7_c_3258_n ) capacitor c=7.46626e-19 \
 //x=34.355 //y=7.4 //x2=34.695 //y2=5.155
cc_1231 ( N_VDD_c_1253_p N_noxref_7_c_3258_n ) capacitor c=0.00198565f \
 //x=35.35 //y=7.4 //x2=34.695 //y2=5.155
cc_1232 ( N_VDD_M97_noxref_d N_noxref_7_c_3258_n ) capacitor c=0.0112985f \
 //x=34.295 //y=5.02 //x2=34.695 //y2=5.155
cc_1233 ( N_VDD_c_1001_n N_noxref_7_c_3262_n ) capacitor c=0.0426864f \
 //x=35.52 //y=7.4 //x2=34.78 //y2=3.33
cc_1234 ( N_VDD_c_1015_p N_noxref_7_c_3235_n ) capacitor c=0.00125279f \
 //x=86.95 //y=7.4 //x2=36.63 //y2=2.08
cc_1235 ( N_VDD_c_1257_p N_noxref_7_c_3235_n ) capacitor c=2.87256e-19 \
 //x=37.105 //y=7.4 //x2=36.63 //y2=2.08
cc_1236 ( N_VDD_c_1001_n N_noxref_7_c_3235_n ) capacitor c=0.0134208f \
 //x=35.52 //y=7.4 //x2=36.63 //y2=2.08
cc_1237 ( N_VDD_c_1259_p N_noxref_7_M90_noxref_g ) capacitor c=0.00675175f \
 //x=29.545 //y=7.4 //x2=28.97 //y2=6.02
cc_1238 ( N_VDD_M89_noxref_d N_noxref_7_M90_noxref_g ) capacitor c=0.015318f \
 //x=28.605 //y=5.02 //x2=28.97 //y2=6.02
cc_1239 ( N_VDD_c_1259_p N_noxref_7_M91_noxref_g ) capacitor c=0.00675379f \
 //x=29.545 //y=7.4 //x2=29.41 //y2=6.02
cc_1240 ( N_VDD_M91_noxref_d N_noxref_7_M91_noxref_g ) capacitor c=0.0394719f \
 //x=29.485 //y=5.02 //x2=29.41 //y2=6.02
cc_1241 ( N_VDD_c_1257_p N_noxref_7_M98_noxref_g ) capacitor c=0.00726866f \
 //x=37.105 //y=7.4 //x2=36.53 //y2=6.02
cc_1242 ( N_VDD_M98_noxref_s N_noxref_7_M98_noxref_g ) capacitor c=0.054195f \
 //x=36.175 //y=5.02 //x2=36.53 //y2=6.02
cc_1243 ( N_VDD_c_1257_p N_noxref_7_M99_noxref_g ) capacitor c=0.00672952f \
 //x=37.105 //y=7.4 //x2=36.97 //y2=6.02
cc_1244 ( N_VDD_M99_noxref_d N_noxref_7_M99_noxref_g ) capacitor c=0.015318f \
 //x=37.045 //y=5.02 //x2=36.97 //y2=6.02
cc_1245 ( N_VDD_c_1001_n N_noxref_7_c_3274_n ) capacitor c=0.0154093f \
 //x=35.52 //y=7.4 //x2=36.63 //y2=4.7
cc_1246 ( N_VDD_c_1015_p N_noxref_7_M92_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=32.095 //y2=5.02
cc_1247 ( N_VDD_c_1242_p N_noxref_7_M92_noxref_d ) capacitor c=0.014035f \
 //x=32.595 //y=7.4 //x2=32.095 //y2=5.02
cc_1248 ( N_VDD_M93_noxref_d N_noxref_7_M92_noxref_d ) capacitor c=0.0664752f \
 //x=32.535 //y=5.02 //x2=32.095 //y2=5.02
cc_1249 ( N_VDD_c_1015_p N_noxref_7_M94_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=32.975 //y2=5.02
cc_1250 ( N_VDD_c_1243_p N_noxref_7_M94_noxref_d ) capacitor c=0.014035f \
 //x=33.475 //y=7.4 //x2=32.975 //y2=5.02
cc_1251 ( N_VDD_c_1001_n N_noxref_7_M94_noxref_d ) capacitor c=4.9285e-19 \
 //x=35.52 //y=7.4 //x2=32.975 //y2=5.02
cc_1252 ( N_VDD_M92_noxref_s N_noxref_7_M94_noxref_d ) capacitor c=0.00130656f \
 //x=31.665 //y=5.02 //x2=32.975 //y2=5.02
cc_1253 ( N_VDD_M93_noxref_d N_noxref_7_M94_noxref_d ) capacitor c=0.0664752f \
 //x=32.535 //y=5.02 //x2=32.975 //y2=5.02
cc_1254 ( N_VDD_M95_noxref_d N_noxref_7_M94_noxref_d ) capacitor c=0.0664752f \
 //x=33.415 //y=5.02 //x2=32.975 //y2=5.02
cc_1255 ( N_VDD_c_1015_p N_noxref_7_M96_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=33.855 //y2=5.02
cc_1256 ( N_VDD_c_1249_p N_noxref_7_M96_noxref_d ) capacitor c=0.014035f \
 //x=34.355 //y=7.4 //x2=33.855 //y2=5.02
cc_1257 ( N_VDD_c_1001_n N_noxref_7_M96_noxref_d ) capacitor c=0.00939849f \
 //x=35.52 //y=7.4 //x2=33.855 //y2=5.02
cc_1258 ( N_VDD_M95_noxref_d N_noxref_7_M96_noxref_d ) capacitor c=0.0664752f \
 //x=33.415 //y=5.02 //x2=33.855 //y2=5.02
cc_1259 ( N_VDD_M97_noxref_d N_noxref_7_M96_noxref_d ) capacitor c=0.0664752f \
 //x=34.295 //y=5.02 //x2=33.855 //y2=5.02
cc_1260 ( N_VDD_M98_noxref_s N_noxref_7_M96_noxref_d ) capacitor c=4.52683e-19 \
 //x=36.175 //y=5.02 //x2=33.855 //y2=5.02
cc_1261 ( N_VDD_c_1015_p N_noxref_8_c_3496_n ) capacitor c=0.00453663f \
 //x=86.95 //y=7.4 //x2=37.545 //y2=5.2
cc_1262 ( N_VDD_c_1257_p N_noxref_8_c_3496_n ) capacitor c=4.48391e-19 \
 //x=37.105 //y=7.4 //x2=37.545 //y2=5.2
cc_1263 ( N_VDD_c_1285_p N_noxref_8_c_3496_n ) capacitor c=4.48391e-19 \
 //x=37.985 //y=7.4 //x2=37.545 //y2=5.2
cc_1264 ( N_VDD_M99_noxref_d N_noxref_8_c_3496_n ) capacitor c=0.0124542f \
 //x=37.045 //y=5.02 //x2=37.545 //y2=5.2
cc_1265 ( N_VDD_c_1001_n N_noxref_8_c_3500_n ) capacitor c=0.00985474f \
 //x=35.52 //y=7.4 //x2=36.835 //y2=5.2
cc_1266 ( N_VDD_M98_noxref_s N_noxref_8_c_3500_n ) capacitor c=0.087833f \
 //x=36.175 //y=5.02 //x2=36.835 //y2=5.2
cc_1267 ( N_VDD_c_1015_p N_noxref_8_c_3502_n ) capacitor c=0.00301575f \
 //x=86.95 //y=7.4 //x2=38.025 //y2=5.2
cc_1268 ( N_VDD_c_1285_p N_noxref_8_c_3502_n ) capacitor c=7.72068e-19 \
 //x=37.985 //y=7.4 //x2=38.025 //y2=5.2
cc_1269 ( N_VDD_M101_noxref_d N_noxref_8_c_3502_n ) capacitor c=0.0158515f \
 //x=37.925 //y=5.02 //x2=38.025 //y2=5.2
cc_1270 ( N_VDD_c_1001_n N_noxref_8_c_3481_n ) capacitor c=0.00151618f \
 //x=35.52 //y=7.4 //x2=38.11 //y2=3.33
cc_1271 ( N_VDD_c_1002_n N_noxref_8_c_3481_n ) capacitor c=0.0428942f \
 //x=38.85 //y=7.4 //x2=38.11 //y2=3.33
cc_1272 ( N_VDD_c_1015_p N_noxref_8_c_3482_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=39.96 //y2=2.08
cc_1273 ( N_VDD_c_1002_n N_noxref_8_c_3482_n ) capacitor c=0.0133749f \
 //x=38.85 //y=7.4 //x2=39.96 //y2=2.08
cc_1274 ( N_VDD_M102_noxref_s N_noxref_8_c_3482_n ) capacitor c=0.0126798f \
 //x=39.805 //y=5.02 //x2=39.96 //y2=2.08
cc_1275 ( N_VDD_c_1297_p N_noxref_8_M102_noxref_g ) capacitor c=0.00749687f \
 //x=40.735 //y=7.4 //x2=40.16 //y2=6.02
cc_1276 ( N_VDD_M102_noxref_s N_noxref_8_M102_noxref_g ) capacitor \
 c=0.0477201f //x=39.805 //y=5.02 //x2=40.16 //y2=6.02
cc_1277 ( N_VDD_c_1297_p N_noxref_8_M103_noxref_g ) capacitor c=0.00675175f \
 //x=40.735 //y=7.4 //x2=40.6 //y2=6.02
cc_1278 ( N_VDD_M103_noxref_d N_noxref_8_M103_noxref_g ) capacitor c=0.015318f \
 //x=40.675 //y=5.02 //x2=40.6 //y2=6.02
cc_1279 ( N_VDD_c_1002_n N_noxref_8_c_3514_n ) capacitor c=0.00757682f \
 //x=38.85 //y=7.4 //x2=40.235 //y2=4.79
cc_1280 ( N_VDD_M102_noxref_s N_noxref_8_c_3514_n ) capacitor c=0.00444914f \
 //x=39.805 //y=5.02 //x2=40.235 //y2=4.79
cc_1281 ( N_VDD_c_1015_p N_noxref_8_M98_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=36.605 //y2=5.02
cc_1282 ( N_VDD_c_1257_p N_noxref_8_M98_noxref_d ) capacitor c=0.0140317f \
 //x=37.105 //y=7.4 //x2=36.605 //y2=5.02
cc_1283 ( N_VDD_c_1002_n N_noxref_8_M98_noxref_d ) capacitor c=6.94454e-19 \
 //x=38.85 //y=7.4 //x2=36.605 //y2=5.02
cc_1284 ( N_VDD_M99_noxref_d N_noxref_8_M98_noxref_d ) capacitor c=0.0664752f \
 //x=37.045 //y=5.02 //x2=36.605 //y2=5.02
cc_1285 ( N_VDD_c_1015_p N_noxref_8_M100_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=37.485 //y2=5.02
cc_1286 ( N_VDD_c_1285_p N_noxref_8_M100_noxref_d ) capacitor c=0.0140317f \
 //x=37.985 //y=7.4 //x2=37.485 //y2=5.02
cc_1287 ( N_VDD_c_1002_n N_noxref_8_M100_noxref_d ) capacitor c=0.0120541f \
 //x=38.85 //y=7.4 //x2=37.485 //y2=5.02
cc_1288 ( N_VDD_M98_noxref_s N_noxref_8_M100_noxref_d ) capacitor \
 c=0.00111971f //x=36.175 //y=5.02 //x2=37.485 //y2=5.02
cc_1289 ( N_VDD_M99_noxref_d N_noxref_8_M100_noxref_d ) capacitor c=0.0664752f \
 //x=37.045 //y=5.02 //x2=37.485 //y2=5.02
cc_1290 ( N_VDD_M101_noxref_d N_noxref_8_M100_noxref_d ) capacitor \
 c=0.0664752f //x=37.925 //y=5.02 //x2=37.485 //y2=5.02
cc_1291 ( N_VDD_M102_noxref_s N_noxref_8_M100_noxref_d ) capacitor \
 c=3.73257e-19 //x=39.805 //y=5.02 //x2=37.485 //y2=5.02
cc_1292 ( N_VDD_c_1015_p N_noxref_9_c_3657_n ) capacitor c=0.00444751f \
 //x=86.95 //y=7.4 //x2=28.225 //y2=5.155
cc_1293 ( N_VDD_c_1315_p N_noxref_9_c_3657_n ) capacitor c=4.31931e-19 \
 //x=27.785 //y=7.4 //x2=28.225 //y2=5.155
cc_1294 ( N_VDD_c_1316_p N_noxref_9_c_3657_n ) capacitor c=4.31906e-19 \
 //x=28.665 //y=7.4 //x2=28.225 //y2=5.155
cc_1295 ( N_VDD_M87_noxref_d N_noxref_9_c_3657_n ) capacitor c=0.0112985f \
 //x=27.725 //y=5.02 //x2=28.225 //y2=5.155
cc_1296 ( N_VDD_c_999_n N_noxref_9_c_3661_n ) capacitor c=0.00863585f //x=25.9 \
 //y=7.4 //x2=27.515 //y2=5.155
cc_1297 ( N_VDD_M86_noxref_s N_noxref_9_c_3661_n ) capacitor c=0.0831083f \
 //x=26.855 //y=5.02 //x2=27.515 //y2=5.155
cc_1298 ( N_VDD_c_1015_p N_noxref_9_c_3663_n ) capacitor c=0.0044221f \
 //x=86.95 //y=7.4 //x2=29.105 //y2=5.155
cc_1299 ( N_VDD_c_1316_p N_noxref_9_c_3663_n ) capacitor c=4.31931e-19 \
 //x=28.665 //y=7.4 //x2=29.105 //y2=5.155
cc_1300 ( N_VDD_c_1259_p N_noxref_9_c_3663_n ) capacitor c=4.31931e-19 \
 //x=29.545 //y=7.4 //x2=29.105 //y2=5.155
cc_1301 ( N_VDD_M89_noxref_d N_noxref_9_c_3663_n ) capacitor c=0.0112985f \
 //x=28.605 //y=5.02 //x2=29.105 //y2=5.155
cc_1302 ( N_VDD_c_1015_p N_noxref_9_c_3667_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=29.885 //y2=5.155
cc_1303 ( N_VDD_c_1259_p N_noxref_9_c_3667_n ) capacitor c=7.46626e-19 \
 //x=29.545 //y=7.4 //x2=29.885 //y2=5.155
cc_1304 ( N_VDD_c_1326_p N_noxref_9_c_3667_n ) capacitor c=0.00198565f \
 //x=30.54 //y=7.4 //x2=29.885 //y2=5.155
cc_1305 ( N_VDD_M91_noxref_d N_noxref_9_c_3667_n ) capacitor c=0.0112985f \
 //x=29.485 //y=5.02 //x2=29.885 //y2=5.155
cc_1306 ( N_VDD_c_1000_n N_noxref_9_c_3671_n ) capacitor c=0.0427116f \
 //x=30.71 //y=7.4 //x2=29.97 //y2=3.7
cc_1307 ( N_VDD_c_1015_p N_noxref_9_c_3634_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=31.82 //y2=2.08
cc_1308 ( N_VDD_c_1000_n N_noxref_9_c_3634_n ) capacitor c=0.0134711f \
 //x=30.71 //y=7.4 //x2=31.82 //y2=2.08
cc_1309 ( N_VDD_M92_noxref_s N_noxref_9_c_3634_n ) capacitor c=0.0126798f \
 //x=31.665 //y=5.02 //x2=31.82 //y2=2.08
cc_1310 ( N_VDD_c_1015_p N_noxref_9_c_3635_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=44.77 //y2=2.08
cc_1311 ( N_VDD_c_1003_n N_noxref_9_c_3635_n ) capacitor c=0.0134269f \
 //x=43.66 //y=7.4 //x2=44.77 //y2=2.08
cc_1312 ( N_VDD_M108_noxref_s N_noxref_9_c_3635_n ) capacitor c=0.0125322f \
 //x=44.615 //y=5.02 //x2=44.77 //y2=2.08
cc_1313 ( N_VDD_c_1242_p N_noxref_9_M92_noxref_g ) capacitor c=0.00749687f \
 //x=32.595 //y=7.4 //x2=32.02 //y2=6.02
cc_1314 ( N_VDD_M92_noxref_s N_noxref_9_M92_noxref_g ) capacitor c=0.0477201f \
 //x=31.665 //y=5.02 //x2=32.02 //y2=6.02
cc_1315 ( N_VDD_c_1242_p N_noxref_9_M93_noxref_g ) capacitor c=0.00675175f \
 //x=32.595 //y=7.4 //x2=32.46 //y2=6.02
cc_1316 ( N_VDD_M93_noxref_d N_noxref_9_M93_noxref_g ) capacitor c=0.015318f \
 //x=32.535 //y=5.02 //x2=32.46 //y2=6.02
cc_1317 ( N_VDD_c_1339_p N_noxref_9_M108_noxref_g ) capacitor c=0.00749687f \
 //x=45.545 //y=7.4 //x2=44.97 //y2=6.02
cc_1318 ( N_VDD_M108_noxref_s N_noxref_9_M108_noxref_g ) capacitor \
 c=0.0477201f //x=44.615 //y=5.02 //x2=44.97 //y2=6.02
cc_1319 ( N_VDD_c_1339_p N_noxref_9_M109_noxref_g ) capacitor c=0.00675175f \
 //x=45.545 //y=7.4 //x2=45.41 //y2=6.02
cc_1320 ( N_VDD_M109_noxref_d N_noxref_9_M109_noxref_g ) capacitor c=0.015318f \
 //x=45.485 //y=5.02 //x2=45.41 //y2=6.02
cc_1321 ( N_VDD_c_1000_n N_noxref_9_c_3686_n ) capacitor c=0.00757682f \
 //x=30.71 //y=7.4 //x2=32.095 //y2=4.79
cc_1322 ( N_VDD_M92_noxref_s N_noxref_9_c_3686_n ) capacitor c=0.00444914f \
 //x=31.665 //y=5.02 //x2=32.095 //y2=4.79
cc_1323 ( N_VDD_c_1003_n N_noxref_9_c_3688_n ) capacitor c=0.00757682f \
 //x=43.66 //y=7.4 //x2=45.045 //y2=4.79
cc_1324 ( N_VDD_M108_noxref_s N_noxref_9_c_3688_n ) capacitor c=0.00444914f \
 //x=44.615 //y=5.02 //x2=45.045 //y2=4.79
cc_1325 ( N_VDD_c_1015_p N_noxref_9_M86_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=27.285 //y2=5.02
cc_1326 ( N_VDD_c_1315_p N_noxref_9_M86_noxref_d ) capacitor c=0.014035f \
 //x=27.785 //y=7.4 //x2=27.285 //y2=5.02
cc_1327 ( N_VDD_M87_noxref_d N_noxref_9_M86_noxref_d ) capacitor c=0.0664752f \
 //x=27.725 //y=5.02 //x2=27.285 //y2=5.02
cc_1328 ( N_VDD_c_1015_p N_noxref_9_M88_noxref_d ) capacitor c=0.00275186f \
 //x=86.95 //y=7.4 //x2=28.165 //y2=5.02
cc_1329 ( N_VDD_c_1316_p N_noxref_9_M88_noxref_d ) capacitor c=0.0140346f \
 //x=28.665 //y=7.4 //x2=28.165 //y2=5.02
cc_1330 ( N_VDD_c_1000_n N_noxref_9_M88_noxref_d ) capacitor c=4.9285e-19 \
 //x=30.71 //y=7.4 //x2=28.165 //y2=5.02
cc_1331 ( N_VDD_M86_noxref_s N_noxref_9_M88_noxref_d ) capacitor c=0.00130656f \
 //x=26.855 //y=5.02 //x2=28.165 //y2=5.02
cc_1332 ( N_VDD_M87_noxref_d N_noxref_9_M88_noxref_d ) capacitor c=0.0664752f \
 //x=27.725 //y=5.02 //x2=28.165 //y2=5.02
cc_1333 ( N_VDD_M89_noxref_d N_noxref_9_M88_noxref_d ) capacitor c=0.0664752f \
 //x=28.605 //y=5.02 //x2=28.165 //y2=5.02
cc_1334 ( N_VDD_c_1015_p N_noxref_9_M90_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=29.045 //y2=5.02
cc_1335 ( N_VDD_c_1259_p N_noxref_9_M90_noxref_d ) capacitor c=0.0137384f \
 //x=29.545 //y=7.4 //x2=29.045 //y2=5.02
cc_1336 ( N_VDD_c_1000_n N_noxref_9_M90_noxref_d ) capacitor c=0.00939849f \
 //x=30.71 //y=7.4 //x2=29.045 //y2=5.02
cc_1337 ( N_VDD_M89_noxref_d N_noxref_9_M90_noxref_d ) capacitor c=0.0664752f \
 //x=28.605 //y=5.02 //x2=29.045 //y2=5.02
cc_1338 ( N_VDD_M91_noxref_d N_noxref_9_M90_noxref_d ) capacitor c=0.0664752f \
 //x=29.485 //y=5.02 //x2=29.045 //y2=5.02
cc_1339 ( N_VDD_M92_noxref_s N_noxref_9_M90_noxref_d ) capacitor c=3.57641e-19 \
 //x=31.665 //y=5.02 //x2=29.045 //y2=5.02
cc_1340 ( N_VDD_c_1015_p N_noxref_10_c_3908_n ) capacitor c=0.00444892f \
 //x=86.95 //y=7.4 //x2=45.985 //y2=5.155
cc_1341 ( N_VDD_c_1339_p N_noxref_10_c_3908_n ) capacitor c=4.31931e-19 \
 //x=45.545 //y=7.4 //x2=45.985 //y2=5.155
cc_1342 ( N_VDD_c_1364_p N_noxref_10_c_3908_n ) capacitor c=4.31931e-19 \
 //x=46.425 //y=7.4 //x2=45.985 //y2=5.155
cc_1343 ( N_VDD_M109_noxref_d N_noxref_10_c_3908_n ) capacitor c=0.0112985f \
 //x=45.485 //y=5.02 //x2=45.985 //y2=5.155
cc_1344 ( N_VDD_c_1003_n N_noxref_10_c_3912_n ) capacitor c=0.00863585f \
 //x=43.66 //y=7.4 //x2=45.275 //y2=5.155
cc_1345 ( N_VDD_M108_noxref_s N_noxref_10_c_3912_n ) capacitor c=0.0831083f \
 //x=44.615 //y=5.02 //x2=45.275 //y2=5.155
cc_1346 ( N_VDD_c_1015_p N_noxref_10_c_3914_n ) capacitor c=0.0044221f \
 //x=86.95 //y=7.4 //x2=46.865 //y2=5.155
cc_1347 ( N_VDD_c_1364_p N_noxref_10_c_3914_n ) capacitor c=4.31931e-19 \
 //x=46.425 //y=7.4 //x2=46.865 //y2=5.155
cc_1348 ( N_VDD_c_1370_p N_noxref_10_c_3914_n ) capacitor c=4.31931e-19 \
 //x=47.305 //y=7.4 //x2=46.865 //y2=5.155
cc_1349 ( N_VDD_M111_noxref_d N_noxref_10_c_3914_n ) capacitor c=0.0112985f \
 //x=46.365 //y=5.02 //x2=46.865 //y2=5.155
cc_1350 ( N_VDD_c_1015_p N_noxref_10_c_3918_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=47.645 //y2=5.155
cc_1351 ( N_VDD_c_1370_p N_noxref_10_c_3918_n ) capacitor c=7.46626e-19 \
 //x=47.305 //y=7.4 //x2=47.645 //y2=5.155
cc_1352 ( N_VDD_c_1374_p N_noxref_10_c_3918_n ) capacitor c=0.00198565f \
 //x=48.3 //y=7.4 //x2=47.645 //y2=5.155
cc_1353 ( N_VDD_M113_noxref_d N_noxref_10_c_3918_n ) capacitor c=0.0112985f \
 //x=47.245 //y=5.02 //x2=47.645 //y2=5.155
cc_1354 ( N_VDD_c_1004_n N_noxref_10_c_3922_n ) capacitor c=0.0426864f \
 //x=48.47 //y=7.4 //x2=47.73 //y2=3.7
cc_1355 ( N_VDD_c_1015_p N_noxref_10_c_3896_n ) capacitor c=0.00125279f \
 //x=86.95 //y=7.4 //x2=49.58 //y2=2.08
cc_1356 ( N_VDD_c_1378_p N_noxref_10_c_3896_n ) capacitor c=2.87256e-19 \
 //x=50.055 //y=7.4 //x2=49.58 //y2=2.08
cc_1357 ( N_VDD_c_1004_n N_noxref_10_c_3896_n ) capacitor c=0.0134208f \
 //x=48.47 //y=7.4 //x2=49.58 //y2=2.08
cc_1358 ( N_VDD_c_1378_p N_noxref_10_M114_noxref_g ) capacitor c=0.00726866f \
 //x=50.055 //y=7.4 //x2=49.48 //y2=6.02
cc_1359 ( N_VDD_M114_noxref_s N_noxref_10_M114_noxref_g ) capacitor \
 c=0.054195f //x=49.125 //y=5.02 //x2=49.48 //y2=6.02
cc_1360 ( N_VDD_c_1378_p N_noxref_10_M115_noxref_g ) capacitor c=0.00672952f \
 //x=50.055 //y=7.4 //x2=49.92 //y2=6.02
cc_1361 ( N_VDD_M115_noxref_d N_noxref_10_M115_noxref_g ) capacitor \
 c=0.015318f //x=49.995 //y=5.02 //x2=49.92 //y2=6.02
cc_1362 ( N_VDD_c_1004_n N_noxref_10_c_3930_n ) capacitor c=0.0154093f \
 //x=48.47 //y=7.4 //x2=49.58 //y2=4.7
cc_1363 ( N_VDD_c_1015_p N_noxref_10_M108_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=45.045 //y2=5.02
cc_1364 ( N_VDD_c_1339_p N_noxref_10_M108_noxref_d ) capacitor c=0.014035f \
 //x=45.545 //y=7.4 //x2=45.045 //y2=5.02
cc_1365 ( N_VDD_M109_noxref_d N_noxref_10_M108_noxref_d ) capacitor \
 c=0.0664752f //x=45.485 //y=5.02 //x2=45.045 //y2=5.02
cc_1366 ( N_VDD_c_1015_p N_noxref_10_M110_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=45.925 //y2=5.02
cc_1367 ( N_VDD_c_1364_p N_noxref_10_M110_noxref_d ) capacitor c=0.014035f \
 //x=46.425 //y=7.4 //x2=45.925 //y2=5.02
cc_1368 ( N_VDD_c_1004_n N_noxref_10_M110_noxref_d ) capacitor c=4.9285e-19 \
 //x=48.47 //y=7.4 //x2=45.925 //y2=5.02
cc_1369 ( N_VDD_M108_noxref_s N_noxref_10_M110_noxref_d ) capacitor \
 c=0.00130656f //x=44.615 //y=5.02 //x2=45.925 //y2=5.02
cc_1370 ( N_VDD_M109_noxref_d N_noxref_10_M110_noxref_d ) capacitor \
 c=0.0664752f //x=45.485 //y=5.02 //x2=45.925 //y2=5.02
cc_1371 ( N_VDD_M111_noxref_d N_noxref_10_M110_noxref_d ) capacitor \
 c=0.0664752f //x=46.365 //y=5.02 //x2=45.925 //y2=5.02
cc_1372 ( N_VDD_c_1015_p N_noxref_10_M112_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=46.805 //y2=5.02
cc_1373 ( N_VDD_c_1370_p N_noxref_10_M112_noxref_d ) capacitor c=0.0137384f \
 //x=47.305 //y=7.4 //x2=46.805 //y2=5.02
cc_1374 ( N_VDD_c_1004_n N_noxref_10_M112_noxref_d ) capacitor c=0.00939849f \
 //x=48.47 //y=7.4 //x2=46.805 //y2=5.02
cc_1375 ( N_VDD_M111_noxref_d N_noxref_10_M112_noxref_d ) capacitor \
 c=0.0664752f //x=46.365 //y=5.02 //x2=46.805 //y2=5.02
cc_1376 ( N_VDD_M113_noxref_d N_noxref_10_M112_noxref_d ) capacitor \
 c=0.0664752f //x=47.245 //y=5.02 //x2=46.805 //y2=5.02
cc_1377 ( N_VDD_M114_noxref_s N_noxref_10_M112_noxref_d ) capacitor \
 c=4.52683e-19 //x=49.125 //y=5.02 //x2=46.805 //y2=5.02
cc_1378 ( N_VDD_c_1000_n N_noxref_11_c_4075_n ) capacitor c=0.0140578f \
 //x=30.71 //y=7.4 //x2=37.255 //y2=4.07
cc_1379 ( N_VDD_c_1001_n N_noxref_11_c_4075_n ) capacitor c=0.0140578f \
 //x=35.52 //y=7.4 //x2=37.255 //y2=4.07
cc_1380 ( N_VDD_c_999_n N_noxref_11_c_4077_n ) capacitor c=0.00116746f \
 //x=25.9 //y=7.4 //x2=27.125 //y2=4.07
cc_1381 ( N_VDD_c_1002_n N_noxref_11_c_4078_n ) capacitor c=0.0140578f \
 //x=38.85 //y=7.4 //x2=42.805 //y2=4.07
cc_1382 ( N_VDD_c_1003_n N_noxref_11_c_4079_n ) capacitor c=0.0140578f \
 //x=43.66 //y=7.4 //x2=50.205 //y2=4.07
cc_1383 ( N_VDD_c_1004_n N_noxref_11_c_4079_n ) capacitor c=0.0140578f \
 //x=48.47 //y=7.4 //x2=50.205 //y2=4.07
cc_1384 ( N_VDD_c_1003_n N_noxref_11_c_4081_n ) capacitor c=0.00104972f \
 //x=43.66 //y=7.4 //x2=43.035 //y2=4.07
cc_1385 ( N_VDD_c_1015_p N_noxref_11_c_4058_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=27.01 //y2=2.08
cc_1386 ( N_VDD_c_999_n N_noxref_11_c_4058_n ) capacitor c=0.0137129f //x=25.9 \
 //y=7.4 //x2=27.01 //y2=2.08
cc_1387 ( N_VDD_M86_noxref_s N_noxref_11_c_4058_n ) capacitor c=0.0120327f \
 //x=26.855 //y=5.02 //x2=27.01 //y2=2.08
cc_1388 ( N_VDD_c_1001_n N_noxref_11_c_4059_n ) capacitor c=4.57806e-19 \
 //x=35.52 //y=7.4 //x2=37.37 //y2=2.08
cc_1389 ( N_VDD_c_1002_n N_noxref_11_c_4059_n ) capacitor c=3.21957e-19 \
 //x=38.85 //y=7.4 //x2=37.37 //y2=2.08
cc_1390 ( N_VDD_c_1015_p N_noxref_11_c_4087_n ) capacitor c=0.00444751f \
 //x=86.95 //y=7.4 //x2=41.175 //y2=5.155
cc_1391 ( N_VDD_c_1297_p N_noxref_11_c_4087_n ) capacitor c=4.31931e-19 \
 //x=40.735 //y=7.4 //x2=41.175 //y2=5.155
cc_1392 ( N_VDD_c_1414_p N_noxref_11_c_4087_n ) capacitor c=4.31906e-19 \
 //x=41.615 //y=7.4 //x2=41.175 //y2=5.155
cc_1393 ( N_VDD_M103_noxref_d N_noxref_11_c_4087_n ) capacitor c=0.0112985f \
 //x=40.675 //y=5.02 //x2=41.175 //y2=5.155
cc_1394 ( N_VDD_c_1002_n N_noxref_11_c_4091_n ) capacitor c=0.00863585f \
 //x=38.85 //y=7.4 //x2=40.465 //y2=5.155
cc_1395 ( N_VDD_M102_noxref_s N_noxref_11_c_4091_n ) capacitor c=0.0831083f \
 //x=39.805 //y=5.02 //x2=40.465 //y2=5.155
cc_1396 ( N_VDD_c_1015_p N_noxref_11_c_4093_n ) capacitor c=0.0044221f \
 //x=86.95 //y=7.4 //x2=42.055 //y2=5.155
cc_1397 ( N_VDD_c_1414_p N_noxref_11_c_4093_n ) capacitor c=4.31931e-19 \
 //x=41.615 //y=7.4 //x2=42.055 //y2=5.155
cc_1398 ( N_VDD_c_1420_p N_noxref_11_c_4093_n ) capacitor c=4.31931e-19 \
 //x=42.495 //y=7.4 //x2=42.055 //y2=5.155
cc_1399 ( N_VDD_M105_noxref_d N_noxref_11_c_4093_n ) capacitor c=0.0112985f \
 //x=41.555 //y=5.02 //x2=42.055 //y2=5.155
cc_1400 ( N_VDD_c_1015_p N_noxref_11_c_4097_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=42.835 //y2=5.155
cc_1401 ( N_VDD_c_1420_p N_noxref_11_c_4097_n ) capacitor c=7.46626e-19 \
 //x=42.495 //y=7.4 //x2=42.835 //y2=5.155
cc_1402 ( N_VDD_c_1424_p N_noxref_11_c_4097_n ) capacitor c=0.00198565f \
 //x=43.49 //y=7.4 //x2=42.835 //y2=5.155
cc_1403 ( N_VDD_M107_noxref_d N_noxref_11_c_4097_n ) capacitor c=0.0112985f \
 //x=42.435 //y=5.02 //x2=42.835 //y2=5.155
cc_1404 ( N_VDD_c_1003_n N_noxref_11_c_4101_n ) capacitor c=0.0429118f \
 //x=43.66 //y=7.4 //x2=42.92 //y2=4.07
cc_1405 ( N_VDD_c_1004_n N_noxref_11_c_4062_n ) capacitor c=4.57806e-19 \
 //x=48.47 //y=7.4 //x2=50.32 //y2=2.08
cc_1406 ( N_VDD_c_1005_n N_noxref_11_c_4062_n ) capacitor c=4.17938e-19 \
 //x=51.8 //y=7.4 //x2=50.32 //y2=2.08
cc_1407 ( N_VDD_c_1315_p N_noxref_11_M86_noxref_g ) capacitor c=0.00749687f \
 //x=27.785 //y=7.4 //x2=27.21 //y2=6.02
cc_1408 ( N_VDD_M86_noxref_s N_noxref_11_M86_noxref_g ) capacitor c=0.0477201f \
 //x=26.855 //y=5.02 //x2=27.21 //y2=6.02
cc_1409 ( N_VDD_c_1315_p N_noxref_11_M87_noxref_g ) capacitor c=0.00675175f \
 //x=27.785 //y=7.4 //x2=27.65 //y2=6.02
cc_1410 ( N_VDD_M87_noxref_d N_noxref_11_M87_noxref_g ) capacitor c=0.015318f \
 //x=27.725 //y=5.02 //x2=27.65 //y2=6.02
cc_1411 ( N_VDD_c_1285_p N_noxref_11_M100_noxref_g ) capacitor c=0.00673971f \
 //x=37.985 //y=7.4 //x2=37.41 //y2=6.02
cc_1412 ( N_VDD_M99_noxref_d N_noxref_11_M100_noxref_g ) capacitor c=0.015318f \
 //x=37.045 //y=5.02 //x2=37.41 //y2=6.02
cc_1413 ( N_VDD_c_1285_p N_noxref_11_M101_noxref_g ) capacitor c=0.00672952f \
 //x=37.985 //y=7.4 //x2=37.85 //y2=6.02
cc_1414 ( N_VDD_c_1002_n N_noxref_11_M101_noxref_g ) capacitor c=0.00928743f \
 //x=38.85 //y=7.4 //x2=37.85 //y2=6.02
cc_1415 ( N_VDD_M101_noxref_d N_noxref_11_M101_noxref_g ) capacitor \
 c=0.0430452f //x=37.925 //y=5.02 //x2=37.85 //y2=6.02
cc_1416 ( N_VDD_c_1438_p N_noxref_11_M116_noxref_g ) capacitor c=0.00673971f \
 //x=50.935 //y=7.4 //x2=50.36 //y2=6.02
cc_1417 ( N_VDD_M115_noxref_d N_noxref_11_M116_noxref_g ) capacitor \
 c=0.015318f //x=49.995 //y=5.02 //x2=50.36 //y2=6.02
cc_1418 ( N_VDD_c_1438_p N_noxref_11_M117_noxref_g ) capacitor c=0.00672952f \
 //x=50.935 //y=7.4 //x2=50.8 //y2=6.02
cc_1419 ( N_VDD_c_1005_n N_noxref_11_M117_noxref_g ) capacitor c=0.00928743f \
 //x=51.8 //y=7.4 //x2=50.8 //y2=6.02
cc_1420 ( N_VDD_M117_noxref_d N_noxref_11_M117_noxref_g ) capacitor \
 c=0.0430452f //x=50.875 //y=5.02 //x2=50.8 //y2=6.02
cc_1421 ( N_VDD_c_999_n N_noxref_11_c_4118_n ) capacitor c=0.00757682f \
 //x=25.9 //y=7.4 //x2=27.285 //y2=4.79
cc_1422 ( N_VDD_M86_noxref_s N_noxref_11_c_4118_n ) capacitor c=0.00444914f \
 //x=26.855 //y=5.02 //x2=27.285 //y2=4.79
cc_1423 ( N_VDD_c_1015_p N_noxref_11_M102_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=40.235 //y2=5.02
cc_1424 ( N_VDD_c_1297_p N_noxref_11_M102_noxref_d ) capacitor c=0.014035f \
 //x=40.735 //y=7.4 //x2=40.235 //y2=5.02
cc_1425 ( N_VDD_M103_noxref_d N_noxref_11_M102_noxref_d ) capacitor \
 c=0.0664752f //x=40.675 //y=5.02 //x2=40.235 //y2=5.02
cc_1426 ( N_VDD_c_1015_p N_noxref_11_M104_noxref_d ) capacitor c=0.00275186f \
 //x=86.95 //y=7.4 //x2=41.115 //y2=5.02
cc_1427 ( N_VDD_c_1414_p N_noxref_11_M104_noxref_d ) capacitor c=0.0140346f \
 //x=41.615 //y=7.4 //x2=41.115 //y2=5.02
cc_1428 ( N_VDD_c_1003_n N_noxref_11_M104_noxref_d ) capacitor c=4.9285e-19 \
 //x=43.66 //y=7.4 //x2=41.115 //y2=5.02
cc_1429 ( N_VDD_M102_noxref_s N_noxref_11_M104_noxref_d ) capacitor \
 c=0.00130656f //x=39.805 //y=5.02 //x2=41.115 //y2=5.02
cc_1430 ( N_VDD_M103_noxref_d N_noxref_11_M104_noxref_d ) capacitor \
 c=0.0664752f //x=40.675 //y=5.02 //x2=41.115 //y2=5.02
cc_1431 ( N_VDD_M105_noxref_d N_noxref_11_M104_noxref_d ) capacitor \
 c=0.0664752f //x=41.555 //y=5.02 //x2=41.115 //y2=5.02
cc_1432 ( N_VDD_c_1015_p N_noxref_11_M106_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=41.995 //y2=5.02
cc_1433 ( N_VDD_c_1420_p N_noxref_11_M106_noxref_d ) capacitor c=0.014035f \
 //x=42.495 //y=7.4 //x2=41.995 //y2=5.02
cc_1434 ( N_VDD_c_1003_n N_noxref_11_M106_noxref_d ) capacitor c=0.00939849f \
 //x=43.66 //y=7.4 //x2=41.995 //y2=5.02
cc_1435 ( N_VDD_M105_noxref_d N_noxref_11_M106_noxref_d ) capacitor \
 c=0.0664752f //x=41.555 //y=5.02 //x2=41.995 //y2=5.02
cc_1436 ( N_VDD_M107_noxref_d N_noxref_11_M106_noxref_d ) capacitor \
 c=0.0664752f //x=42.435 //y=5.02 //x2=41.995 //y2=5.02
cc_1437 ( N_VDD_M108_noxref_s N_noxref_11_M106_noxref_d ) capacitor \
 c=3.57641e-19 //x=44.615 //y=5.02 //x2=41.995 //y2=5.02
cc_1438 ( N_VDD_c_1015_p N_D_c_4448_n ) capacitor c=2.03486e-19 //x=86.95 \
 //y=7.4 //x2=7.03 //y2=2.08
cc_1439 ( N_VDD_c_994_n N_D_c_4448_n ) capacitor c=5.89117e-19 //x=4.81 \
 //y=7.4 //x2=7.03 //y2=2.08
cc_1440 ( N_VDD_c_1015_p N_D_c_4449_n ) capacitor c=2.03486e-19 //x=86.95 \
 //y=7.4 //x2=32.93 //y2=2.08
cc_1441 ( N_VDD_c_1000_n N_D_c_4449_n ) capacitor c=5.89117e-19 //x=30.71 \
 //y=7.4 //x2=32.93 //y2=2.08
cc_1442 ( N_VDD_c_1015_p N_D_c_4450_n ) capacitor c=2.03486e-19 //x=86.95 \
 //y=7.4 //x2=58.83 //y2=2.08
cc_1443 ( N_VDD_c_1006_n N_D_c_4450_n ) capacitor c=5.89117e-19 //x=56.61 \
 //y=7.4 //x2=58.83 //y2=2.08
cc_1444 ( N_VDD_c_1017_p N_D_M62_noxref_g ) capacitor c=0.00676195f //x=7.575 \
 //y=7.4 //x2=7 //y2=6.02
cc_1445 ( N_VDD_M61_noxref_d N_D_M62_noxref_g ) capacitor c=0.015318f \
 //x=6.635 //y=5.02 //x2=7 //y2=6.02
cc_1446 ( N_VDD_c_1017_p N_D_M63_noxref_g ) capacitor c=0.00675175f //x=7.575 \
 //y=7.4 //x2=7.44 //y2=6.02
cc_1447 ( N_VDD_M63_noxref_d N_D_M63_noxref_g ) capacitor c=0.015318f \
 //x=7.515 //y=5.02 //x2=7.44 //y2=6.02
cc_1448 ( N_VDD_c_1243_p N_D_M94_noxref_g ) capacitor c=0.00676195f //x=33.475 \
 //y=7.4 //x2=32.9 //y2=6.02
cc_1449 ( N_VDD_M93_noxref_d N_D_M94_noxref_g ) capacitor c=0.015318f \
 //x=32.535 //y=5.02 //x2=32.9 //y2=6.02
cc_1450 ( N_VDD_c_1243_p N_D_M95_noxref_g ) capacitor c=0.00675175f //x=33.475 \
 //y=7.4 //x2=33.34 //y2=6.02
cc_1451 ( N_VDD_M95_noxref_d N_D_M95_noxref_g ) capacitor c=0.015318f \
 //x=33.415 //y=5.02 //x2=33.34 //y2=6.02
cc_1452 ( N_VDD_c_1474_p N_D_M126_noxref_g ) capacitor c=0.00676195f \
 //x=59.375 //y=7.4 //x2=58.8 //y2=6.02
cc_1453 ( N_VDD_M125_noxref_d N_D_M126_noxref_g ) capacitor c=0.015318f \
 //x=58.435 //y=5.02 //x2=58.8 //y2=6.02
cc_1454 ( N_VDD_c_1474_p N_D_M127_noxref_g ) capacitor c=0.00675175f \
 //x=59.375 //y=7.4 //x2=59.24 //y2=6.02
cc_1455 ( N_VDD_M127_noxref_d N_D_M127_noxref_g ) capacitor c=0.015318f \
 //x=59.315 //y=5.02 //x2=59.24 //y2=6.02
cc_1456 ( N_VDD_c_1015_p N_CLK_c_4808_n ) capacitor c=0.0956945f //x=86.95 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1457 ( N_VDD_c_1100_p N_CLK_c_4808_n ) capacitor c=0.00258496f //x=4.64 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1458 ( N_VDD_c_1480_p N_CLK_c_4808_n ) capacitor c=0.00328994f //x=5.815 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1459 ( N_VDD_c_1016_p N_CLK_c_4808_n ) capacitor c=0.00135925f //x=6.695 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1460 ( N_VDD_c_1027_p N_CLK_c_4808_n ) capacitor c=0.00258496f //x=9.45 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1461 ( N_VDD_c_1483_p N_CLK_c_4808_n ) capacitor c=0.00209689f //x=10.325 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1462 ( N_VDD_c_1031_p N_CLK_c_4808_n ) capacitor c=7.81728e-19 //x=11.205 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1463 ( N_VDD_c_1485_p N_CLK_c_4808_n ) capacitor c=0.00205475f //x=12.78 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1464 ( N_VDD_c_1486_p N_CLK_c_4808_n ) capacitor c=0.00328994f //x=13.955 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1465 ( N_VDD_c_1071_p N_CLK_c_4808_n ) capacitor c=0.00135925f //x=14.835 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1466 ( N_VDD_c_994_n N_CLK_c_4808_n ) capacitor c=0.0389825f //x=4.81 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1467 ( N_VDD_c_995_n N_CLK_c_4808_n ) capacitor c=0.0389825f //x=9.62 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1468 ( N_VDD_c_996_n N_CLK_c_4808_n ) capacitor c=0.0389825f //x=12.95 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_1469 ( N_VDD_M60_noxref_s N_CLK_c_4808_n ) capacitor c=0.00179496f \
 //x=5.765 //y=5.02 //x2=15.055 //y2=4.44
cc_1470 ( N_VDD_M66_noxref_s N_CLK_c_4808_n ) capacitor c=0.00541054f \
 //x=10.275 //y=5.02 //x2=15.055 //y2=4.44
cc_1471 ( N_VDD_M69_noxref_d N_CLK_c_4808_n ) capacitor c=6.7165e-19 \
 //x=12.025 //y=5.02 //x2=15.055 //y2=4.44
cc_1472 ( N_VDD_M70_noxref_s N_CLK_c_4808_n ) capacitor c=0.00179496f \
 //x=13.905 //y=5.02 //x2=15.055 //y2=4.44
cc_1473 ( N_VDD_c_1015_p N_CLK_c_4825_n ) capacitor c=0.00146064f //x=86.95 \
 //y=7.4 //x2=2.335 //y2=4.44
cc_1474 ( N_VDD_c_1015_p N_CLK_c_4826_n ) capacitor c=0.0956945f //x=86.95 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1475 ( N_VDD_c_1166_p N_CLK_c_4826_n ) capacitor c=0.00258496f //x=17.59 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1476 ( N_VDD_c_1498_p N_CLK_c_4826_n ) capacitor c=0.00328994f //x=18.765 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1477 ( N_VDD_c_1113_p N_CLK_c_4826_n ) capacitor c=0.00135925f //x=19.645 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1478 ( N_VDD_c_1181_p N_CLK_c_4826_n ) capacitor c=0.00258496f //x=22.4 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1479 ( N_VDD_c_1501_p N_CLK_c_4826_n ) capacitor c=0.00209689f //x=23.275 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1480 ( N_VDD_c_1185_p N_CLK_c_4826_n ) capacitor c=7.81728e-19 //x=24.155 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1481 ( N_VDD_c_1503_p N_CLK_c_4826_n ) capacitor c=0.00205475f //x=25.73 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1482 ( N_VDD_c_1504_p N_CLK_c_4826_n ) capacitor c=0.00328994f //x=26.905 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1483 ( N_VDD_c_1315_p N_CLK_c_4826_n ) capacitor c=0.00135925f //x=27.785 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1484 ( N_VDD_c_997_n N_CLK_c_4826_n ) capacitor c=0.0389825f //x=17.76 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1485 ( N_VDD_c_998_n N_CLK_c_4826_n ) capacitor c=0.0389825f //x=22.57 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1486 ( N_VDD_c_999_n N_CLK_c_4826_n ) capacitor c=0.0404757f //x=25.9 \
 //y=7.4 //x2=28.005 //y2=4.44
cc_1487 ( N_VDD_M76_noxref_s N_CLK_c_4826_n ) capacitor c=0.00179496f \
 //x=18.715 //y=5.02 //x2=28.005 //y2=4.44
cc_1488 ( N_VDD_M82_noxref_s N_CLK_c_4826_n ) capacitor c=0.00541054f \
 //x=23.225 //y=5.02 //x2=28.005 //y2=4.44
cc_1489 ( N_VDD_M85_noxref_d N_CLK_c_4826_n ) capacitor c=6.7165e-19 \
 //x=24.975 //y=5.02 //x2=28.005 //y2=4.44
cc_1490 ( N_VDD_M86_noxref_s N_CLK_c_4826_n ) capacitor c=0.00179496f \
 //x=26.855 //y=5.02 //x2=28.005 //y2=4.44
cc_1491 ( N_VDD_c_1015_p N_CLK_c_4843_n ) capacitor c=0.00120845f //x=86.95 \
 //y=7.4 //x2=15.285 //y2=4.44
cc_1492 ( N_VDD_c_1015_p N_CLK_c_4844_n ) capacitor c=0.0956945f //x=86.95 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1493 ( N_VDD_c_1326_p N_CLK_c_4844_n ) capacitor c=0.00258496f //x=30.54 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1494 ( N_VDD_c_1516_p N_CLK_c_4844_n ) capacitor c=0.00328994f //x=31.715 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1495 ( N_VDD_c_1242_p N_CLK_c_4844_n ) capacitor c=0.00135925f //x=32.595 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1496 ( N_VDD_c_1253_p N_CLK_c_4844_n ) capacitor c=0.00258496f //x=35.35 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1497 ( N_VDD_c_1519_p N_CLK_c_4844_n ) capacitor c=0.00209689f //x=36.225 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1498 ( N_VDD_c_1257_p N_CLK_c_4844_n ) capacitor c=7.81728e-19 //x=37.105 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1499 ( N_VDD_c_1521_p N_CLK_c_4844_n ) capacitor c=0.00205475f //x=38.68 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1500 ( N_VDD_c_1522_p N_CLK_c_4844_n ) capacitor c=0.00328994f //x=39.855 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1501 ( N_VDD_c_1297_p N_CLK_c_4844_n ) capacitor c=0.00135925f //x=40.735 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1502 ( N_VDD_c_1000_n N_CLK_c_4844_n ) capacitor c=0.0389825f //x=30.71 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1503 ( N_VDD_c_1001_n N_CLK_c_4844_n ) capacitor c=0.0389825f //x=35.52 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1504 ( N_VDD_c_1002_n N_CLK_c_4844_n ) capacitor c=0.0389825f //x=38.85 \
 //y=7.4 //x2=40.955 //y2=4.44
cc_1505 ( N_VDD_M92_noxref_s N_CLK_c_4844_n ) capacitor c=0.00179496f \
 //x=31.665 //y=5.02 //x2=40.955 //y2=4.44
cc_1506 ( N_VDD_M98_noxref_s N_CLK_c_4844_n ) capacitor c=0.00541054f \
 //x=36.175 //y=5.02 //x2=40.955 //y2=4.44
cc_1507 ( N_VDD_M101_noxref_d N_CLK_c_4844_n ) capacitor c=6.7165e-19 \
 //x=37.925 //y=5.02 //x2=40.955 //y2=4.44
cc_1508 ( N_VDD_M102_noxref_s N_CLK_c_4844_n ) capacitor c=0.00179496f \
 //x=39.805 //y=5.02 //x2=40.955 //y2=4.44
cc_1509 ( N_VDD_c_1015_p N_CLK_c_4861_n ) capacitor c=0.00120845f //x=86.95 \
 //y=7.4 //x2=28.235 //y2=4.44
cc_1510 ( N_VDD_c_1015_p N_CLK_c_4862_n ) capacitor c=0.0956945f //x=86.95 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1511 ( N_VDD_c_1424_p N_CLK_c_4862_n ) capacitor c=0.00258496f //x=43.49 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1512 ( N_VDD_c_1534_p N_CLK_c_4862_n ) capacitor c=0.00328994f //x=44.665 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1513 ( N_VDD_c_1339_p N_CLK_c_4862_n ) capacitor c=0.00135925f //x=45.545 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1514 ( N_VDD_c_1374_p N_CLK_c_4862_n ) capacitor c=0.00258496f //x=48.3 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1515 ( N_VDD_c_1537_p N_CLK_c_4862_n ) capacitor c=0.00209689f //x=49.175 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1516 ( N_VDD_c_1378_p N_CLK_c_4862_n ) capacitor c=7.81728e-19 //x=50.055 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1517 ( N_VDD_c_1539_p N_CLK_c_4862_n ) capacitor c=0.00205475f //x=51.63 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1518 ( N_VDD_c_1540_p N_CLK_c_4862_n ) capacitor c=0.00328994f //x=52.805 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1519 ( N_VDD_c_1541_p N_CLK_c_4862_n ) capacitor c=0.00135925f //x=53.685 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1520 ( N_VDD_c_1003_n N_CLK_c_4862_n ) capacitor c=0.0389825f //x=43.66 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1521 ( N_VDD_c_1004_n N_CLK_c_4862_n ) capacitor c=0.0389825f //x=48.47 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1522 ( N_VDD_c_1005_n N_CLK_c_4862_n ) capacitor c=0.0392569f //x=51.8 \
 //y=7.4 //x2=53.905 //y2=4.44
cc_1523 ( N_VDD_M108_noxref_s N_CLK_c_4862_n ) capacitor c=0.00179496f \
 //x=44.615 //y=5.02 //x2=53.905 //y2=4.44
cc_1524 ( N_VDD_M114_noxref_s N_CLK_c_4862_n ) capacitor c=0.00541054f \
 //x=49.125 //y=5.02 //x2=53.905 //y2=4.44
cc_1525 ( N_VDD_M117_noxref_d N_CLK_c_4862_n ) capacitor c=6.7165e-19 \
 //x=50.875 //y=5.02 //x2=53.905 //y2=4.44
cc_1526 ( N_VDD_M118_noxref_s N_CLK_c_4862_n ) capacitor c=0.00179496f \
 //x=52.755 //y=5.02 //x2=53.905 //y2=4.44
cc_1527 ( N_VDD_c_1015_p N_CLK_c_4879_n ) capacitor c=0.00120845f //x=86.95 \
 //y=7.4 //x2=41.185 //y2=4.44
cc_1528 ( N_VDD_c_1015_p N_CLK_c_4880_n ) capacitor c=0.0971263f //x=86.95 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1529 ( N_VDD_c_1551_p N_CLK_c_4880_n ) capacitor c=0.00258496f //x=56.44 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1530 ( N_VDD_c_1552_p N_CLK_c_4880_n ) capacitor c=0.00328994f //x=57.615 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1531 ( N_VDD_c_1553_p N_CLK_c_4880_n ) capacitor c=0.00135925f //x=58.495 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1532 ( N_VDD_c_1554_p N_CLK_c_4880_n ) capacitor c=0.00258496f //x=61.25 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1533 ( N_VDD_c_1555_p N_CLK_c_4880_n ) capacitor c=0.00209689f //x=62.125 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1534 ( N_VDD_c_1556_p N_CLK_c_4880_n ) capacitor c=7.81728e-19 //x=63.005 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1535 ( N_VDD_c_1557_p N_CLK_c_4880_n ) capacitor c=0.00205475f //x=64.58 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1536 ( N_VDD_c_1558_p N_CLK_c_4880_n ) capacitor c=0.00328994f //x=65.755 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1537 ( N_VDD_c_1559_p N_CLK_c_4880_n ) capacitor c=0.00135925f //x=66.635 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1538 ( N_VDD_c_1006_n N_CLK_c_4880_n ) capacitor c=0.0389825f //x=56.61 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1539 ( N_VDD_c_1007_n N_CLK_c_4880_n ) capacitor c=0.0389825f //x=61.42 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1540 ( N_VDD_c_1008_n N_CLK_c_4880_n ) capacitor c=0.0389825f //x=64.75 \
 //y=7.4 //x2=66.855 //y2=4.44
cc_1541 ( N_VDD_M124_noxref_s N_CLK_c_4880_n ) capacitor c=0.00179496f \
 //x=57.565 //y=5.02 //x2=66.855 //y2=4.44
cc_1542 ( N_VDD_M130_noxref_s N_CLK_c_4880_n ) capacitor c=0.00541054f \
 //x=62.075 //y=5.02 //x2=66.855 //y2=4.44
cc_1543 ( N_VDD_M133_noxref_d N_CLK_c_4880_n ) capacitor c=6.7165e-19 \
 //x=63.825 //y=5.02 //x2=66.855 //y2=4.44
cc_1544 ( N_VDD_M134_noxref_s N_CLK_c_4880_n ) capacitor c=0.00179496f \
 //x=65.705 //y=5.02 //x2=66.855 //y2=4.44
cc_1545 ( N_VDD_c_1015_p N_CLK_c_4897_n ) capacitor c=0.00120845f //x=86.95 \
 //y=7.4 //x2=54.135 //y2=4.44
cc_1546 ( N_VDD_c_1015_p N_CLK_c_4802_n ) capacitor c=2.03287e-19 //x=86.95 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_1547 ( N_VDD_c_992_n N_CLK_c_4802_n ) capacitor c=9.53425e-19 //x=0.74 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_1548 ( N_VDD_c_1015_p N_CLK_c_4803_n ) capacitor c=2.03287e-19 //x=86.95 \
 //y=7.4 //x2=15.17 //y2=2.08
cc_1549 ( N_VDD_c_996_n N_CLK_c_4803_n ) capacitor c=6.15921e-19 //x=12.95 \
 //y=7.4 //x2=15.17 //y2=2.08
cc_1550 ( N_VDD_c_1015_p N_CLK_c_4804_n ) capacitor c=2.03287e-19 //x=86.95 \
 //y=7.4 //x2=28.12 //y2=2.08
cc_1551 ( N_VDD_c_999_n N_CLK_c_4804_n ) capacitor c=7.21466e-19 //x=25.9 \
 //y=7.4 //x2=28.12 //y2=2.08
cc_1552 ( N_VDD_c_1015_p N_CLK_c_4805_n ) capacitor c=2.03287e-19 //x=86.95 \
 //y=7.4 //x2=41.07 //y2=2.08
cc_1553 ( N_VDD_c_1002_n N_CLK_c_4805_n ) capacitor c=6.15921e-19 //x=38.85 \
 //y=7.4 //x2=41.07 //y2=2.08
cc_1554 ( N_VDD_c_1015_p N_CLK_c_4806_n ) capacitor c=2.03287e-19 //x=86.95 \
 //y=7.4 //x2=54.02 //y2=2.08
cc_1555 ( N_VDD_c_1005_n N_CLK_c_4806_n ) capacitor c=7.21466e-19 //x=51.8 \
 //y=7.4 //x2=54.02 //y2=2.08
cc_1556 ( N_VDD_c_1015_p N_CLK_c_4807_n ) capacitor c=2.03287e-19 //x=86.95 \
 //y=7.4 //x2=66.97 //y2=2.08
cc_1557 ( N_VDD_c_1008_n N_CLK_c_4807_n ) capacitor c=6.15921e-19 //x=64.75 \
 //y=7.4 //x2=66.97 //y2=2.08
cc_1558 ( N_VDD_c_1090_p N_CLK_M56_noxref_g ) capacitor c=0.00676195f \
 //x=2.765 //y=7.4 //x2=2.19 //y2=6.02
cc_1559 ( N_VDD_M55_noxref_d N_CLK_M56_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=2.19 //y2=6.02
cc_1560 ( N_VDD_c_1090_p N_CLK_M57_noxref_g ) capacitor c=0.00675175f \
 //x=2.765 //y=7.4 //x2=2.63 //y2=6.02
cc_1561 ( N_VDD_M57_noxref_d N_CLK_M57_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=2.63 //y2=6.02
cc_1562 ( N_VDD_c_1156_p N_CLK_M72_noxref_g ) capacitor c=0.00676195f \
 //x=15.715 //y=7.4 //x2=15.14 //y2=6.02
cc_1563 ( N_VDD_M71_noxref_d N_CLK_M72_noxref_g ) capacitor c=0.015318f \
 //x=14.775 //y=5.02 //x2=15.14 //y2=6.02
cc_1564 ( N_VDD_c_1156_p N_CLK_M73_noxref_g ) capacitor c=0.00675175f \
 //x=15.715 //y=7.4 //x2=15.58 //y2=6.02
cc_1565 ( N_VDD_M73_noxref_d N_CLK_M73_noxref_g ) capacitor c=0.015318f \
 //x=15.655 //y=5.02 //x2=15.58 //y2=6.02
cc_1566 ( N_VDD_c_1316_p N_CLK_M88_noxref_g ) capacitor c=0.00676195f \
 //x=28.665 //y=7.4 //x2=28.09 //y2=6.02
cc_1567 ( N_VDD_M87_noxref_d N_CLK_M88_noxref_g ) capacitor c=0.015318f \
 //x=27.725 //y=5.02 //x2=28.09 //y2=6.02
cc_1568 ( N_VDD_c_1316_p N_CLK_M89_noxref_g ) capacitor c=0.00675175f \
 //x=28.665 //y=7.4 //x2=28.53 //y2=6.02
cc_1569 ( N_VDD_M89_noxref_d N_CLK_M89_noxref_g ) capacitor c=0.015318f \
 //x=28.605 //y=5.02 //x2=28.53 //y2=6.02
cc_1570 ( N_VDD_c_1414_p N_CLK_M104_noxref_g ) capacitor c=0.00676195f \
 //x=41.615 //y=7.4 //x2=41.04 //y2=6.02
cc_1571 ( N_VDD_M103_noxref_d N_CLK_M104_noxref_g ) capacitor c=0.015318f \
 //x=40.675 //y=5.02 //x2=41.04 //y2=6.02
cc_1572 ( N_VDD_c_1414_p N_CLK_M105_noxref_g ) capacitor c=0.00675175f \
 //x=41.615 //y=7.4 //x2=41.48 //y2=6.02
cc_1573 ( N_VDD_M105_noxref_d N_CLK_M105_noxref_g ) capacitor c=0.015318f \
 //x=41.555 //y=5.02 //x2=41.48 //y2=6.02
cc_1574 ( N_VDD_c_1596_p N_CLK_M120_noxref_g ) capacitor c=0.00676195f \
 //x=54.565 //y=7.4 //x2=53.99 //y2=6.02
cc_1575 ( N_VDD_M119_noxref_d N_CLK_M120_noxref_g ) capacitor c=0.015318f \
 //x=53.625 //y=5.02 //x2=53.99 //y2=6.02
cc_1576 ( N_VDD_c_1596_p N_CLK_M121_noxref_g ) capacitor c=0.00675175f \
 //x=54.565 //y=7.4 //x2=54.43 //y2=6.02
cc_1577 ( N_VDD_M121_noxref_d N_CLK_M121_noxref_g ) capacitor c=0.015318f \
 //x=54.505 //y=5.02 //x2=54.43 //y2=6.02
cc_1578 ( N_VDD_c_1600_p N_CLK_M136_noxref_g ) capacitor c=0.00676195f \
 //x=67.515 //y=7.4 //x2=66.94 //y2=6.02
cc_1579 ( N_VDD_M135_noxref_d N_CLK_M136_noxref_g ) capacitor c=0.015318f \
 //x=66.575 //y=5.02 //x2=66.94 //y2=6.02
cc_1580 ( N_VDD_c_1600_p N_CLK_M137_noxref_g ) capacitor c=0.00675175f \
 //x=67.515 //y=7.4 //x2=67.38 //y2=6.02
cc_1581 ( N_VDD_M137_noxref_d N_CLK_M137_noxref_g ) capacitor c=0.015318f \
 //x=67.455 //y=5.02 //x2=67.38 //y2=6.02
cc_1582 ( N_VDD_c_1015_p N_noxref_14_c_5611_n ) capacitor c=0.00444751f \
 //x=86.95 //y=7.4 //x2=54.125 //y2=5.155
cc_1583 ( N_VDD_c_1541_p N_noxref_14_c_5611_n ) capacitor c=4.31931e-19 \
 //x=53.685 //y=7.4 //x2=54.125 //y2=5.155
cc_1584 ( N_VDD_c_1596_p N_noxref_14_c_5611_n ) capacitor c=4.31906e-19 \
 //x=54.565 //y=7.4 //x2=54.125 //y2=5.155
cc_1585 ( N_VDD_M119_noxref_d N_noxref_14_c_5611_n ) capacitor c=0.0112985f \
 //x=53.625 //y=5.02 //x2=54.125 //y2=5.155
cc_1586 ( N_VDD_c_1005_n N_noxref_14_c_5615_n ) capacitor c=0.00863585f \
 //x=51.8 //y=7.4 //x2=53.415 //y2=5.155
cc_1587 ( N_VDD_M118_noxref_s N_noxref_14_c_5615_n ) capacitor c=0.0831083f \
 //x=52.755 //y=5.02 //x2=53.415 //y2=5.155
cc_1588 ( N_VDD_c_1015_p N_noxref_14_c_5617_n ) capacitor c=0.0044221f \
 //x=86.95 //y=7.4 //x2=55.005 //y2=5.155
cc_1589 ( N_VDD_c_1596_p N_noxref_14_c_5617_n ) capacitor c=4.31931e-19 \
 //x=54.565 //y=7.4 //x2=55.005 //y2=5.155
cc_1590 ( N_VDD_c_1612_p N_noxref_14_c_5617_n ) capacitor c=4.31931e-19 \
 //x=55.445 //y=7.4 //x2=55.005 //y2=5.155
cc_1591 ( N_VDD_M121_noxref_d N_noxref_14_c_5617_n ) capacitor c=0.0112985f \
 //x=54.505 //y=5.02 //x2=55.005 //y2=5.155
cc_1592 ( N_VDD_c_1015_p N_noxref_14_c_5621_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=55.785 //y2=5.155
cc_1593 ( N_VDD_c_1612_p N_noxref_14_c_5621_n ) capacitor c=7.46626e-19 \
 //x=55.445 //y=7.4 //x2=55.785 //y2=5.155
cc_1594 ( N_VDD_c_1551_p N_noxref_14_c_5621_n ) capacitor c=0.00198565f \
 //x=56.44 //y=7.4 //x2=55.785 //y2=5.155
cc_1595 ( N_VDD_M123_noxref_d N_noxref_14_c_5621_n ) capacitor c=0.0112985f \
 //x=55.385 //y=5.02 //x2=55.785 //y2=5.155
cc_1596 ( N_VDD_c_1006_n N_noxref_14_c_5625_n ) capacitor c=0.0427116f \
 //x=56.61 //y=7.4 //x2=55.87 //y2=3.7
cc_1597 ( N_VDD_c_1015_p N_noxref_14_c_5588_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=57.72 //y2=2.08
cc_1598 ( N_VDD_c_1006_n N_noxref_14_c_5588_n ) capacitor c=0.0134711f \
 //x=56.61 //y=7.4 //x2=57.72 //y2=2.08
cc_1599 ( N_VDD_M124_noxref_s N_noxref_14_c_5588_n ) capacitor c=0.0126798f \
 //x=57.565 //y=5.02 //x2=57.72 //y2=2.08
cc_1600 ( N_VDD_c_1015_p N_noxref_14_c_5589_n ) capacitor c=9.23542e-19 \
 //x=86.95 //y=7.4 //x2=70.67 //y2=2.08
cc_1601 ( N_VDD_c_1009_n N_noxref_14_c_5589_n ) capacitor c=0.0160182f \
 //x=69.56 //y=7.4 //x2=70.67 //y2=2.08
cc_1602 ( N_VDD_M140_noxref_s N_noxref_14_c_5589_n ) capacitor c=0.0128378f \
 //x=70.515 //y=5.02 //x2=70.67 //y2=2.08
cc_1603 ( N_VDD_c_1553_p N_noxref_14_M124_noxref_g ) capacitor c=0.00749687f \
 //x=58.495 //y=7.4 //x2=57.92 //y2=6.02
cc_1604 ( N_VDD_M124_noxref_s N_noxref_14_M124_noxref_g ) capacitor \
 c=0.0477201f //x=57.565 //y=5.02 //x2=57.92 //y2=6.02
cc_1605 ( N_VDD_c_1553_p N_noxref_14_M125_noxref_g ) capacitor c=0.00675175f \
 //x=58.495 //y=7.4 //x2=58.36 //y2=6.02
cc_1606 ( N_VDD_M125_noxref_d N_noxref_14_M125_noxref_g ) capacitor \
 c=0.015318f //x=58.435 //y=5.02 //x2=58.36 //y2=6.02
cc_1607 ( N_VDD_c_1629_p N_noxref_14_M140_noxref_g ) capacitor c=0.00749687f \
 //x=71.445 //y=7.4 //x2=70.87 //y2=6.02
cc_1608 ( N_VDD_M140_noxref_s N_noxref_14_M140_noxref_g ) capacitor \
 c=0.0477201f //x=70.515 //y=5.02 //x2=70.87 //y2=6.02
cc_1609 ( N_VDD_c_1629_p N_noxref_14_M141_noxref_g ) capacitor c=0.00675175f \
 //x=71.445 //y=7.4 //x2=71.31 //y2=6.02
cc_1610 ( N_VDD_M141_noxref_d N_noxref_14_M141_noxref_g ) capacitor \
 c=0.015318f //x=71.385 //y=5.02 //x2=71.31 //y2=6.02
cc_1611 ( N_VDD_c_1006_n N_noxref_14_c_5640_n ) capacitor c=0.00757682f \
 //x=56.61 //y=7.4 //x2=57.995 //y2=4.79
cc_1612 ( N_VDD_M124_noxref_s N_noxref_14_c_5640_n ) capacitor c=0.00444914f \
 //x=57.565 //y=5.02 //x2=57.995 //y2=4.79
cc_1613 ( N_VDD_c_1009_n N_noxref_14_c_5642_n ) capacitor c=0.00757682f \
 //x=69.56 //y=7.4 //x2=70.945 //y2=4.79
cc_1614 ( N_VDD_M140_noxref_s N_noxref_14_c_5642_n ) capacitor c=0.00445134f \
 //x=70.515 //y=5.02 //x2=70.945 //y2=4.79
cc_1615 ( N_VDD_c_1015_p N_noxref_14_M118_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=53.185 //y2=5.02
cc_1616 ( N_VDD_c_1541_p N_noxref_14_M118_noxref_d ) capacitor c=0.014035f \
 //x=53.685 //y=7.4 //x2=53.185 //y2=5.02
cc_1617 ( N_VDD_M119_noxref_d N_noxref_14_M118_noxref_d ) capacitor \
 c=0.0664752f //x=53.625 //y=5.02 //x2=53.185 //y2=5.02
cc_1618 ( N_VDD_c_1015_p N_noxref_14_M120_noxref_d ) capacitor c=0.00275186f \
 //x=86.95 //y=7.4 //x2=54.065 //y2=5.02
cc_1619 ( N_VDD_c_1596_p N_noxref_14_M120_noxref_d ) capacitor c=0.0140346f \
 //x=54.565 //y=7.4 //x2=54.065 //y2=5.02
cc_1620 ( N_VDD_c_1006_n N_noxref_14_M120_noxref_d ) capacitor c=4.9285e-19 \
 //x=56.61 //y=7.4 //x2=54.065 //y2=5.02
cc_1621 ( N_VDD_M118_noxref_s N_noxref_14_M120_noxref_d ) capacitor \
 c=0.00130656f //x=52.755 //y=5.02 //x2=54.065 //y2=5.02
cc_1622 ( N_VDD_M119_noxref_d N_noxref_14_M120_noxref_d ) capacitor \
 c=0.0664752f //x=53.625 //y=5.02 //x2=54.065 //y2=5.02
cc_1623 ( N_VDD_M121_noxref_d N_noxref_14_M120_noxref_d ) capacitor \
 c=0.0664752f //x=54.505 //y=5.02 //x2=54.065 //y2=5.02
cc_1624 ( N_VDD_c_1015_p N_noxref_14_M122_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=54.945 //y2=5.02
cc_1625 ( N_VDD_c_1612_p N_noxref_14_M122_noxref_d ) capacitor c=0.0137384f \
 //x=55.445 //y=7.4 //x2=54.945 //y2=5.02
cc_1626 ( N_VDD_c_1006_n N_noxref_14_M122_noxref_d ) capacitor c=0.00939849f \
 //x=56.61 //y=7.4 //x2=54.945 //y2=5.02
cc_1627 ( N_VDD_M121_noxref_d N_noxref_14_M122_noxref_d ) capacitor \
 c=0.0664752f //x=54.505 //y=5.02 //x2=54.945 //y2=5.02
cc_1628 ( N_VDD_M123_noxref_d N_noxref_14_M122_noxref_d ) capacitor \
 c=0.0664752f //x=55.385 //y=5.02 //x2=54.945 //y2=5.02
cc_1629 ( N_VDD_M124_noxref_s N_noxref_14_M122_noxref_d ) capacitor \
 c=3.57641e-19 //x=57.565 //y=5.02 //x2=54.945 //y2=5.02
cc_1630 ( N_VDD_c_995_n N_RN_c_5913_n ) capacitor c=6.09414e-19 //x=9.62 \
 //y=7.4 //x2=8.14 //y2=2.08
cc_1631 ( N_VDD_c_997_n N_RN_c_5914_n ) capacitor c=7.21146e-19 //x=17.76 \
 //y=7.4 //x2=16.28 //y2=2.08
cc_1632 ( N_VDD_c_1015_p N_RN_c_5915_n ) capacitor c=2.03486e-19 //x=86.95 \
 //y=7.4 //x2=19.98 //y2=2.08
cc_1633 ( N_VDD_c_997_n N_RN_c_5915_n ) capacitor c=6.15067e-19 //x=17.76 \
 //y=7.4 //x2=19.98 //y2=2.08
cc_1634 ( N_VDD_c_1001_n N_RN_c_5916_n ) capacitor c=6.09414e-19 //x=35.52 \
 //y=7.4 //x2=34.04 //y2=2.08
cc_1635 ( N_VDD_c_1003_n N_RN_c_5917_n ) capacitor c=7.21146e-19 //x=43.66 \
 //y=7.4 //x2=42.18 //y2=2.08
cc_1636 ( N_VDD_c_1015_p N_RN_c_5918_n ) capacitor c=2.03486e-19 //x=86.95 \
 //y=7.4 //x2=45.88 //y2=2.08
cc_1637 ( N_VDD_c_1003_n N_RN_c_5918_n ) capacitor c=6.15067e-19 //x=43.66 \
 //y=7.4 //x2=45.88 //y2=2.08
cc_1638 ( N_VDD_c_1007_n N_RN_c_5919_n ) capacitor c=6.09414e-19 //x=61.42 \
 //y=7.4 //x2=59.94 //y2=2.08
cc_1639 ( N_VDD_c_1009_n N_RN_c_5920_n ) capacitor c=0.00120861f //x=69.56 \
 //y=7.4 //x2=68.08 //y2=2.08
cc_1640 ( N_VDD_c_1015_p N_RN_c_5921_n ) capacitor c=2.05828e-19 //x=86.95 \
 //y=7.4 //x2=71.78 //y2=2.08
cc_1641 ( N_VDD_c_1009_n N_RN_c_5921_n ) capacitor c=7.30063e-19 //x=69.56 \
 //y=7.4 //x2=71.78 //y2=2.08
cc_1642 ( N_VDD_c_1023_p N_RN_M64_noxref_g ) capacitor c=0.00675175f //x=8.455 \
 //y=7.4 //x2=7.88 //y2=6.02
cc_1643 ( N_VDD_M63_noxref_d N_RN_M64_noxref_g ) capacitor c=0.015318f \
 //x=7.515 //y=5.02 //x2=7.88 //y2=6.02
cc_1644 ( N_VDD_c_1023_p N_RN_M65_noxref_g ) capacitor c=0.00675379f //x=8.455 \
 //y=7.4 //x2=8.32 //y2=6.02
cc_1645 ( N_VDD_M65_noxref_d N_RN_M65_noxref_g ) capacitor c=0.0394719f \
 //x=8.395 //y=5.02 //x2=8.32 //y2=6.02
cc_1646 ( N_VDD_c_1162_p N_RN_M74_noxref_g ) capacitor c=0.00675175f \
 //x=16.595 //y=7.4 //x2=16.02 //y2=6.02
cc_1647 ( N_VDD_M73_noxref_d N_RN_M74_noxref_g ) capacitor c=0.015318f \
 //x=15.655 //y=5.02 //x2=16.02 //y2=6.02
cc_1648 ( N_VDD_c_1162_p N_RN_M75_noxref_g ) capacitor c=0.00675379f \
 //x=16.595 //y=7.4 //x2=16.46 //y2=6.02
cc_1649 ( N_VDD_M75_noxref_d N_RN_M75_noxref_g ) capacitor c=0.0394719f \
 //x=16.535 //y=5.02 //x2=16.46 //y2=6.02
cc_1650 ( N_VDD_c_1171_p N_RN_M78_noxref_g ) capacitor c=0.00676195f \
 //x=20.525 //y=7.4 //x2=19.95 //y2=6.02
cc_1651 ( N_VDD_M77_noxref_d N_RN_M78_noxref_g ) capacitor c=0.015318f \
 //x=19.585 //y=5.02 //x2=19.95 //y2=6.02
cc_1652 ( N_VDD_c_1171_p N_RN_M79_noxref_g ) capacitor c=0.00675175f \
 //x=20.525 //y=7.4 //x2=20.39 //y2=6.02
cc_1653 ( N_VDD_M79_noxref_d N_RN_M79_noxref_g ) capacitor c=0.015318f \
 //x=20.465 //y=5.02 //x2=20.39 //y2=6.02
cc_1654 ( N_VDD_c_1249_p N_RN_M96_noxref_g ) capacitor c=0.00675175f \
 //x=34.355 //y=7.4 //x2=33.78 //y2=6.02
cc_1655 ( N_VDD_M95_noxref_d N_RN_M96_noxref_g ) capacitor c=0.015318f \
 //x=33.415 //y=5.02 //x2=33.78 //y2=6.02
cc_1656 ( N_VDD_c_1249_p N_RN_M97_noxref_g ) capacitor c=0.00675379f \
 //x=34.355 //y=7.4 //x2=34.22 //y2=6.02
cc_1657 ( N_VDD_M97_noxref_d N_RN_M97_noxref_g ) capacitor c=0.0394719f \
 //x=34.295 //y=5.02 //x2=34.22 //y2=6.02
cc_1658 ( N_VDD_c_1420_p N_RN_M106_noxref_g ) capacitor c=0.00675175f \
 //x=42.495 //y=7.4 //x2=41.92 //y2=6.02
cc_1659 ( N_VDD_M105_noxref_d N_RN_M106_noxref_g ) capacitor c=0.015318f \
 //x=41.555 //y=5.02 //x2=41.92 //y2=6.02
cc_1660 ( N_VDD_c_1420_p N_RN_M107_noxref_g ) capacitor c=0.00675379f \
 //x=42.495 //y=7.4 //x2=42.36 //y2=6.02
cc_1661 ( N_VDD_M107_noxref_d N_RN_M107_noxref_g ) capacitor c=0.0394719f \
 //x=42.435 //y=5.02 //x2=42.36 //y2=6.02
cc_1662 ( N_VDD_c_1364_p N_RN_M110_noxref_g ) capacitor c=0.00676195f \
 //x=46.425 //y=7.4 //x2=45.85 //y2=6.02
cc_1663 ( N_VDD_M109_noxref_d N_RN_M110_noxref_g ) capacitor c=0.015318f \
 //x=45.485 //y=5.02 //x2=45.85 //y2=6.02
cc_1664 ( N_VDD_c_1364_p N_RN_M111_noxref_g ) capacitor c=0.00675175f \
 //x=46.425 //y=7.4 //x2=46.29 //y2=6.02
cc_1665 ( N_VDD_M111_noxref_d N_RN_M111_noxref_g ) capacitor c=0.015318f \
 //x=46.365 //y=5.02 //x2=46.29 //y2=6.02
cc_1666 ( N_VDD_c_1688_p N_RN_M128_noxref_g ) capacitor c=0.00675175f \
 //x=60.255 //y=7.4 //x2=59.68 //y2=6.02
cc_1667 ( N_VDD_M127_noxref_d N_RN_M128_noxref_g ) capacitor c=0.015318f \
 //x=59.315 //y=5.02 //x2=59.68 //y2=6.02
cc_1668 ( N_VDD_c_1688_p N_RN_M129_noxref_g ) capacitor c=0.00675379f \
 //x=60.255 //y=7.4 //x2=60.12 //y2=6.02
cc_1669 ( N_VDD_M129_noxref_d N_RN_M129_noxref_g ) capacitor c=0.0394719f \
 //x=60.195 //y=5.02 //x2=60.12 //y2=6.02
cc_1670 ( N_VDD_c_1692_p N_RN_M138_noxref_g ) capacitor c=0.00675175f \
 //x=68.395 //y=7.4 //x2=67.82 //y2=6.02
cc_1671 ( N_VDD_M137_noxref_d N_RN_M138_noxref_g ) capacitor c=0.015318f \
 //x=67.455 //y=5.02 //x2=67.82 //y2=6.02
cc_1672 ( N_VDD_c_1692_p N_RN_M139_noxref_g ) capacitor c=0.00675379f \
 //x=68.395 //y=7.4 //x2=68.26 //y2=6.02
cc_1673 ( N_VDD_M139_noxref_d N_RN_M139_noxref_g ) capacitor c=0.0394719f \
 //x=68.335 //y=5.02 //x2=68.26 //y2=6.02
cc_1674 ( N_VDD_c_1696_p N_RN_M142_noxref_g ) capacitor c=0.00676195f \
 //x=72.325 //y=7.4 //x2=71.75 //y2=6.02
cc_1675 ( N_VDD_M141_noxref_d N_RN_M142_noxref_g ) capacitor c=0.015318f \
 //x=71.385 //y=5.02 //x2=71.75 //y2=6.02
cc_1676 ( N_VDD_c_1696_p N_RN_M143_noxref_g ) capacitor c=0.00675175f \
 //x=72.325 //y=7.4 //x2=72.19 //y2=6.02
cc_1677 ( N_VDD_M143_noxref_d N_RN_M143_noxref_g ) capacitor c=0.015318f \
 //x=72.265 //y=5.02 //x2=72.19 //y2=6.02
cc_1678 ( N_VDD_c_1006_n N_noxref_16_c_6831_n ) capacitor c=0.0140578f \
 //x=56.61 //y=7.4 //x2=63.155 //y2=4.07
cc_1679 ( N_VDD_c_1007_n N_noxref_16_c_6831_n ) capacitor c=0.0140578f \
 //x=61.42 //y=7.4 //x2=63.155 //y2=4.07
cc_1680 ( N_VDD_c_1005_n N_noxref_16_c_6833_n ) capacitor c=0.00116746f \
 //x=51.8 //y=7.4 //x2=53.025 //y2=4.07
cc_1681 ( N_VDD_c_1015_p N_noxref_16_c_6834_n ) capacitor c=0.0256485f \
 //x=86.95 //y=7.4 //x2=68.705 //y2=4.07
cc_1682 ( N_VDD_c_1008_n N_noxref_16_c_6834_n ) capacitor c=0.0140578f \
 //x=64.75 //y=7.4 //x2=68.705 //y2=4.07
cc_1683 ( N_VDD_c_1015_p N_noxref_16_c_6836_n ) capacitor c=0.0316106f \
 //x=86.95 //y=7.4 //x2=73.515 //y2=4.07
cc_1684 ( N_VDD_c_1706_p N_noxref_16_c_6836_n ) capacitor c=0.0016229f \
 //x=69.39 //y=7.4 //x2=73.515 //y2=4.07
cc_1685 ( N_VDD_c_1707_p N_noxref_16_c_6836_n ) capacitor c=0.0027159f \
 //x=70.565 //y=7.4 //x2=73.515 //y2=4.07
cc_1686 ( N_VDD_c_1629_p N_noxref_16_c_6836_n ) capacitor c=0.00113459f \
 //x=71.445 //y=7.4 //x2=73.515 //y2=4.07
cc_1687 ( N_VDD_c_1009_n N_noxref_16_c_6836_n ) capacitor c=0.0269494f \
 //x=69.56 //y=7.4 //x2=73.515 //y2=4.07
cc_1688 ( N_VDD_M140_noxref_s N_noxref_16_c_6836_n ) capacitor c=0.00122826f \
 //x=70.515 //y=5.02 //x2=73.515 //y2=4.07
cc_1689 ( N_VDD_c_1015_p N_noxref_16_c_6842_n ) capacitor c=0.00175338f \
 //x=86.95 //y=7.4 //x2=68.935 //y2=4.07
cc_1690 ( N_VDD_c_1706_p N_noxref_16_c_6842_n ) capacitor c=5.20513e-19 \
 //x=69.39 //y=7.4 //x2=68.935 //y2=4.07
cc_1691 ( N_VDD_c_1009_n N_noxref_16_c_6842_n ) capacitor c=0.00104972f \
 //x=69.56 //y=7.4 //x2=68.935 //y2=4.07
cc_1692 ( N_VDD_c_1015_p N_noxref_16_c_6845_n ) capacitor c=0.0114971f \
 //x=86.95 //y=7.4 //x2=75.365 //y2=4.07
cc_1693 ( N_VDD_c_1715_p N_noxref_16_c_6845_n ) capacitor c=0.0016229f \
 //x=74.2 //y=7.4 //x2=75.365 //y2=4.07
cc_1694 ( N_VDD_c_1716_p N_noxref_16_c_6845_n ) capacitor c=0.00172186f \
 //x=75.075 //y=7.4 //x2=75.365 //y2=4.07
cc_1695 ( N_VDD_c_1717_p N_noxref_16_c_6845_n ) capacitor c=2.43243e-19 \
 //x=75.955 //y=7.4 //x2=75.365 //y2=4.07
cc_1696 ( N_VDD_c_1010_n N_noxref_16_c_6845_n ) capacitor c=0.0269494f \
 //x=74.37 //y=7.4 //x2=75.365 //y2=4.07
cc_1697 ( N_VDD_M146_noxref_s N_noxref_16_c_6845_n ) capacitor c=0.00363031f \
 //x=75.025 //y=5.02 //x2=75.365 //y2=4.07
cc_1698 ( N_VDD_c_1015_p N_noxref_16_c_6851_n ) capacitor c=0.00175338f \
 //x=86.95 //y=7.4 //x2=73.745 //y2=4.07
cc_1699 ( N_VDD_c_1715_p N_noxref_16_c_6851_n ) capacitor c=5.20513e-19 \
 //x=74.2 //y=7.4 //x2=73.745 //y2=4.07
cc_1700 ( N_VDD_c_1010_n N_noxref_16_c_6851_n ) capacitor c=5.12647e-19 \
 //x=74.37 //y=7.4 //x2=73.745 //y2=4.07
cc_1701 ( N_VDD_c_1015_p N_noxref_16_c_6854_n ) capacitor c=0.00560422f \
 //x=86.95 //y=7.4 //x2=76.105 //y2=4.07
cc_1702 ( N_VDD_c_1015_p N_noxref_16_c_6855_n ) capacitor c=0.0015497f \
 //x=86.95 //y=7.4 //x2=75.595 //y2=4.07
cc_1703 ( N_VDD_c_1717_p N_noxref_16_c_6855_n ) capacitor c=4.18761e-19 \
 //x=75.955 //y=7.4 //x2=75.595 //y2=4.07
cc_1704 ( N_VDD_c_1010_n N_noxref_16_c_6855_n ) capacitor c=3.58282e-19 \
 //x=74.37 //y=7.4 //x2=75.595 //y2=4.07
cc_1705 ( N_VDD_c_1015_p N_noxref_16_c_6801_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=52.91 //y2=2.08
cc_1706 ( N_VDD_c_1005_n N_noxref_16_c_6801_n ) capacitor c=0.0137129f \
 //x=51.8 //y=7.4 //x2=52.91 //y2=2.08
cc_1707 ( N_VDD_M118_noxref_s N_noxref_16_c_6801_n ) capacitor c=0.0120327f \
 //x=52.755 //y=5.02 //x2=52.91 //y2=2.08
cc_1708 ( N_VDD_c_1007_n N_noxref_16_c_6802_n ) capacitor c=4.57806e-19 \
 //x=61.42 //y=7.4 //x2=63.27 //y2=2.08
cc_1709 ( N_VDD_c_1008_n N_noxref_16_c_6802_n ) capacitor c=3.21957e-19 \
 //x=64.75 //y=7.4 //x2=63.27 //y2=2.08
cc_1710 ( N_VDD_c_1015_p N_noxref_16_c_6863_n ) capacitor c=0.00444751f \
 //x=86.95 //y=7.4 //x2=67.075 //y2=5.155
cc_1711 ( N_VDD_c_1559_p N_noxref_16_c_6863_n ) capacitor c=4.31931e-19 \
 //x=66.635 //y=7.4 //x2=67.075 //y2=5.155
cc_1712 ( N_VDD_c_1600_p N_noxref_16_c_6863_n ) capacitor c=4.31906e-19 \
 //x=67.515 //y=7.4 //x2=67.075 //y2=5.155
cc_1713 ( N_VDD_M135_noxref_d N_noxref_16_c_6863_n ) capacitor c=0.0112985f \
 //x=66.575 //y=5.02 //x2=67.075 //y2=5.155
cc_1714 ( N_VDD_c_1008_n N_noxref_16_c_6867_n ) capacitor c=0.00863585f \
 //x=64.75 //y=7.4 //x2=66.365 //y2=5.155
cc_1715 ( N_VDD_M134_noxref_s N_noxref_16_c_6867_n ) capacitor c=0.0831083f \
 //x=65.705 //y=5.02 //x2=66.365 //y2=5.155
cc_1716 ( N_VDD_c_1015_p N_noxref_16_c_6869_n ) capacitor c=0.00448996f \
 //x=86.95 //y=7.4 //x2=67.955 //y2=5.155
cc_1717 ( N_VDD_c_1600_p N_noxref_16_c_6869_n ) capacitor c=4.32228e-19 \
 //x=67.515 //y=7.4 //x2=67.955 //y2=5.155
cc_1718 ( N_VDD_c_1692_p N_noxref_16_c_6869_n ) capacitor c=4.32228e-19 \
 //x=68.395 //y=7.4 //x2=67.955 //y2=5.155
cc_1719 ( N_VDD_M137_noxref_d N_noxref_16_c_6869_n ) capacitor c=0.0115147f \
 //x=67.455 //y=5.02 //x2=67.955 //y2=5.155
cc_1720 ( N_VDD_c_1015_p N_noxref_16_c_6873_n ) capacitor c=0.00442469f \
 //x=86.95 //y=7.4 //x2=68.735 //y2=5.155
cc_1721 ( N_VDD_c_1692_p N_noxref_16_c_6873_n ) capacitor c=7.47666e-19 \
 //x=68.395 //y=7.4 //x2=68.735 //y2=5.155
cc_1722 ( N_VDD_c_1706_p N_noxref_16_c_6873_n ) capacitor c=0.00198959f \
 //x=69.39 //y=7.4 //x2=68.735 //y2=5.155
cc_1723 ( N_VDD_M139_noxref_d N_noxref_16_c_6873_n ) capacitor c=0.0115147f \
 //x=68.335 //y=5.02 //x2=68.735 //y2=5.155
cc_1724 ( N_VDD_c_1009_n N_noxref_16_c_6877_n ) capacitor c=0.0452313f \
 //x=69.56 //y=7.4 //x2=68.82 //y2=4.07
cc_1725 ( N_VDD_c_1015_p N_noxref_16_c_6878_n ) capacitor c=0.004515f \
 //x=86.95 //y=7.4 //x2=71.885 //y2=5.155
cc_1726 ( N_VDD_c_1629_p N_noxref_16_c_6878_n ) capacitor c=4.32228e-19 \
 //x=71.445 //y=7.4 //x2=71.885 //y2=5.155
cc_1727 ( N_VDD_c_1696_p N_noxref_16_c_6878_n ) capacitor c=4.32228e-19 \
 //x=72.325 //y=7.4 //x2=71.885 //y2=5.155
cc_1728 ( N_VDD_M141_noxref_d N_noxref_16_c_6878_n ) capacitor c=0.0115147f \
 //x=71.385 //y=5.02 //x2=71.885 //y2=5.155
cc_1729 ( N_VDD_c_1009_n N_noxref_16_c_6882_n ) capacitor c=0.00863585f \
 //x=69.56 //y=7.4 //x2=71.175 //y2=5.155
cc_1730 ( N_VDD_M140_noxref_s N_noxref_16_c_6882_n ) capacitor c=0.0831083f \
 //x=70.515 //y=5.02 //x2=71.175 //y2=5.155
cc_1731 ( N_VDD_c_1015_p N_noxref_16_c_6884_n ) capacitor c=0.00448996f \
 //x=86.95 //y=7.4 //x2=72.765 //y2=5.155
cc_1732 ( N_VDD_c_1696_p N_noxref_16_c_6884_n ) capacitor c=4.32228e-19 \
 //x=72.325 //y=7.4 //x2=72.765 //y2=5.155
cc_1733 ( N_VDD_c_1755_p N_noxref_16_c_6884_n ) capacitor c=4.32228e-19 \
 //x=73.205 //y=7.4 //x2=72.765 //y2=5.155
cc_1734 ( N_VDD_M143_noxref_d N_noxref_16_c_6884_n ) capacitor c=0.0115147f \
 //x=72.265 //y=5.02 //x2=72.765 //y2=5.155
cc_1735 ( N_VDD_c_1015_p N_noxref_16_c_6888_n ) capacitor c=0.00442469f \
 //x=86.95 //y=7.4 //x2=73.545 //y2=5.155
cc_1736 ( N_VDD_c_1755_p N_noxref_16_c_6888_n ) capacitor c=7.47666e-19 \
 //x=73.205 //y=7.4 //x2=73.545 //y2=5.155
cc_1737 ( N_VDD_c_1715_p N_noxref_16_c_6888_n ) capacitor c=0.00198959f \
 //x=74.2 //y=7.4 //x2=73.545 //y2=5.155
cc_1738 ( N_VDD_M145_noxref_d N_noxref_16_c_6888_n ) capacitor c=0.0115147f \
 //x=73.145 //y=5.02 //x2=73.545 //y2=5.155
cc_1739 ( N_VDD_c_1010_n N_noxref_16_c_6892_n ) capacitor c=0.0456347f \
 //x=74.37 //y=7.4 //x2=73.63 //y2=4.07
cc_1740 ( N_VDD_c_1015_p N_noxref_16_c_6806_n ) capacitor c=0.00126142f \
 //x=86.95 //y=7.4 //x2=75.48 //y2=2.08
cc_1741 ( N_VDD_c_1717_p N_noxref_16_c_6806_n ) capacitor c=2.8777e-19 \
 //x=75.955 //y=7.4 //x2=75.48 //y2=2.08
cc_1742 ( N_VDD_c_1010_n N_noxref_16_c_6806_n ) capacitor c=0.0159978f \
 //x=74.37 //y=7.4 //x2=75.48 //y2=2.08
cc_1743 ( N_VDD_c_1010_n N_noxref_16_c_6807_n ) capacitor c=6.24345e-19 \
 //x=74.37 //y=7.4 //x2=76.22 //y2=2.08
cc_1744 ( N_VDD_c_1011_n N_noxref_16_c_6807_n ) capacitor c=9.09239e-19 \
 //x=77.7 //y=7.4 //x2=76.22 //y2=2.08
cc_1745 ( N_VDD_c_1541_p N_noxref_16_M118_noxref_g ) capacitor c=0.00749687f \
 //x=53.685 //y=7.4 //x2=53.11 //y2=6.02
cc_1746 ( N_VDD_M118_noxref_s N_noxref_16_M118_noxref_g ) capacitor \
 c=0.0477201f //x=52.755 //y=5.02 //x2=53.11 //y2=6.02
cc_1747 ( N_VDD_c_1541_p N_noxref_16_M119_noxref_g ) capacitor c=0.00675175f \
 //x=53.685 //y=7.4 //x2=53.55 //y2=6.02
cc_1748 ( N_VDD_M119_noxref_d N_noxref_16_M119_noxref_g ) capacitor \
 c=0.015318f //x=53.625 //y=5.02 //x2=53.55 //y2=6.02
cc_1749 ( N_VDD_c_1771_p N_noxref_16_M132_noxref_g ) capacitor c=0.00673971f \
 //x=63.885 //y=7.4 //x2=63.31 //y2=6.02
cc_1750 ( N_VDD_M131_noxref_d N_noxref_16_M132_noxref_g ) capacitor \
 c=0.015318f //x=62.945 //y=5.02 //x2=63.31 //y2=6.02
cc_1751 ( N_VDD_c_1771_p N_noxref_16_M133_noxref_g ) capacitor c=0.00672952f \
 //x=63.885 //y=7.4 //x2=63.75 //y2=6.02
cc_1752 ( N_VDD_c_1008_n N_noxref_16_M133_noxref_g ) capacitor c=0.00928743f \
 //x=64.75 //y=7.4 //x2=63.75 //y2=6.02
cc_1753 ( N_VDD_M133_noxref_d N_noxref_16_M133_noxref_g ) capacitor \
 c=0.0430452f //x=63.825 //y=5.02 //x2=63.75 //y2=6.02
cc_1754 ( N_VDD_c_1717_p N_noxref_16_M146_noxref_g ) capacitor c=0.00726866f \
 //x=75.955 //y=7.4 //x2=75.38 //y2=6.02
cc_1755 ( N_VDD_M146_noxref_s N_noxref_16_M146_noxref_g ) capacitor \
 c=0.054195f //x=75.025 //y=5.02 //x2=75.38 //y2=6.02
cc_1756 ( N_VDD_c_1717_p N_noxref_16_M147_noxref_g ) capacitor c=0.00672952f \
 //x=75.955 //y=7.4 //x2=75.82 //y2=6.02
cc_1757 ( N_VDD_M147_noxref_d N_noxref_16_M147_noxref_g ) capacitor \
 c=0.015318f //x=75.895 //y=5.02 //x2=75.82 //y2=6.02
cc_1758 ( N_VDD_c_1780_p N_noxref_16_M148_noxref_g ) capacitor c=0.00673971f \
 //x=76.835 //y=7.4 //x2=76.26 //y2=6.02
cc_1759 ( N_VDD_M147_noxref_d N_noxref_16_M148_noxref_g ) capacitor \
 c=0.015318f //x=75.895 //y=5.02 //x2=76.26 //y2=6.02
cc_1760 ( N_VDD_c_1780_p N_noxref_16_M149_noxref_g ) capacitor c=0.00672952f \
 //x=76.835 //y=7.4 //x2=76.7 //y2=6.02
cc_1761 ( N_VDD_c_1011_n N_noxref_16_M149_noxref_g ) capacitor c=0.00814158f \
 //x=77.7 //y=7.4 //x2=76.7 //y2=6.02
cc_1762 ( N_VDD_M149_noxref_d N_noxref_16_M149_noxref_g ) capacitor \
 c=0.0430452f //x=76.775 //y=5.02 //x2=76.7 //y2=6.02
cc_1763 ( N_VDD_c_1005_n N_noxref_16_c_6916_n ) capacitor c=0.00757682f \
 //x=51.8 //y=7.4 //x2=53.185 //y2=4.79
cc_1764 ( N_VDD_M118_noxref_s N_noxref_16_c_6916_n ) capacitor c=0.00444914f \
 //x=52.755 //y=5.02 //x2=53.185 //y2=4.79
cc_1765 ( N_VDD_c_1010_n N_noxref_16_c_6918_n ) capacitor c=0.0154093f \
 //x=74.37 //y=7.4 //x2=75.48 //y2=4.7
cc_1766 ( N_VDD_c_1015_p N_noxref_16_M134_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=66.135 //y2=5.02
cc_1767 ( N_VDD_c_1559_p N_noxref_16_M134_noxref_d ) capacitor c=0.014035f \
 //x=66.635 //y=7.4 //x2=66.135 //y2=5.02
cc_1768 ( N_VDD_M135_noxref_d N_noxref_16_M134_noxref_d ) capacitor \
 c=0.0664752f //x=66.575 //y=5.02 //x2=66.135 //y2=5.02
cc_1769 ( N_VDD_c_1015_p N_noxref_16_M136_noxref_d ) capacitor c=0.00282723f \
 //x=86.95 //y=7.4 //x2=67.015 //y2=5.02
cc_1770 ( N_VDD_c_1600_p N_noxref_16_M136_noxref_d ) capacitor c=0.0140856f \
 //x=67.515 //y=7.4 //x2=67.015 //y2=5.02
cc_1771 ( N_VDD_c_1009_n N_noxref_16_M136_noxref_d ) capacitor c=4.9285e-19 \
 //x=69.56 //y=7.4 //x2=67.015 //y2=5.02
cc_1772 ( N_VDD_M134_noxref_s N_noxref_16_M136_noxref_d ) capacitor \
 c=0.00130656f //x=65.705 //y=5.02 //x2=67.015 //y2=5.02
cc_1773 ( N_VDD_M135_noxref_d N_noxref_16_M136_noxref_d ) capacitor \
 c=0.0664752f //x=66.575 //y=5.02 //x2=67.015 //y2=5.02
cc_1774 ( N_VDD_M137_noxref_d N_noxref_16_M136_noxref_d ) capacitor \
 c=0.0664752f //x=67.455 //y=5.02 //x2=67.015 //y2=5.02
cc_1775 ( N_VDD_c_1015_p N_noxref_16_M138_noxref_d ) capacitor c=0.00285091f \
 //x=86.95 //y=7.4 //x2=67.895 //y2=5.02
cc_1776 ( N_VDD_c_1692_p N_noxref_16_M138_noxref_d ) capacitor c=0.0138051f \
 //x=68.395 //y=7.4 //x2=67.895 //y2=5.02
cc_1777 ( N_VDD_c_1009_n N_noxref_16_M138_noxref_d ) capacitor c=0.00939849f \
 //x=69.56 //y=7.4 //x2=67.895 //y2=5.02
cc_1778 ( N_VDD_M137_noxref_d N_noxref_16_M138_noxref_d ) capacitor \
 c=0.0664752f //x=67.455 //y=5.02 //x2=67.895 //y2=5.02
cc_1779 ( N_VDD_M139_noxref_d N_noxref_16_M138_noxref_d ) capacitor \
 c=0.0664752f //x=68.335 //y=5.02 //x2=67.895 //y2=5.02
cc_1780 ( N_VDD_M140_noxref_s N_noxref_16_M138_noxref_d ) capacitor \
 c=3.57641e-19 //x=70.515 //y=5.02 //x2=67.895 //y2=5.02
cc_1781 ( N_VDD_c_1015_p N_noxref_16_M140_noxref_d ) capacitor c=0.00285091f \
 //x=86.95 //y=7.4 //x2=70.945 //y2=5.02
cc_1782 ( N_VDD_c_1629_p N_noxref_16_M140_noxref_d ) capacitor c=0.0141016f \
 //x=71.445 //y=7.4 //x2=70.945 //y2=5.02
cc_1783 ( N_VDD_M141_noxref_d N_noxref_16_M140_noxref_d ) capacitor \
 c=0.0664752f //x=71.385 //y=5.02 //x2=70.945 //y2=5.02
cc_1784 ( N_VDD_c_1015_p N_noxref_16_M142_noxref_d ) capacitor c=0.00285091f \
 //x=86.95 //y=7.4 //x2=71.825 //y2=5.02
cc_1785 ( N_VDD_c_1696_p N_noxref_16_M142_noxref_d ) capacitor c=0.0141016f \
 //x=72.325 //y=7.4 //x2=71.825 //y2=5.02
cc_1786 ( N_VDD_c_1010_n N_noxref_16_M142_noxref_d ) capacitor c=4.9285e-19 \
 //x=74.37 //y=7.4 //x2=71.825 //y2=5.02
cc_1787 ( N_VDD_M140_noxref_s N_noxref_16_M142_noxref_d ) capacitor \
 c=0.00130656f //x=70.515 //y=5.02 //x2=71.825 //y2=5.02
cc_1788 ( N_VDD_M141_noxref_d N_noxref_16_M142_noxref_d ) capacitor \
 c=0.0664752f //x=71.385 //y=5.02 //x2=71.825 //y2=5.02
cc_1789 ( N_VDD_M143_noxref_d N_noxref_16_M142_noxref_d ) capacitor \
 c=0.0664752f //x=72.265 //y=5.02 //x2=71.825 //y2=5.02
cc_1790 ( N_VDD_c_1015_p N_noxref_16_M144_noxref_d ) capacitor c=0.00285091f \
 //x=86.95 //y=7.4 //x2=72.705 //y2=5.02
cc_1791 ( N_VDD_c_1755_p N_noxref_16_M144_noxref_d ) capacitor c=0.0138051f \
 //x=73.205 //y=7.4 //x2=72.705 //y2=5.02
cc_1792 ( N_VDD_c_1010_n N_noxref_16_M144_noxref_d ) capacitor c=0.00939849f \
 //x=74.37 //y=7.4 //x2=72.705 //y2=5.02
cc_1793 ( N_VDD_M143_noxref_d N_noxref_16_M144_noxref_d ) capacitor \
 c=0.0664752f //x=72.265 //y=5.02 //x2=72.705 //y2=5.02
cc_1794 ( N_VDD_M145_noxref_d N_noxref_16_M144_noxref_d ) capacitor \
 c=0.0664752f //x=73.145 //y=5.02 //x2=72.705 //y2=5.02
cc_1795 ( N_VDD_M146_noxref_s N_noxref_16_M144_noxref_d ) capacitor \
 c=4.52683e-19 //x=75.025 //y=5.02 //x2=72.705 //y2=5.02
cc_1796 ( N_VDD_c_1005_n N_noxref_17_c_7362_n ) capacitor c=0.0045786f \
 //x=51.8 //y=7.4 //x2=55.015 //y2=3.33
cc_1797 ( N_VDD_c_1015_p N_noxref_17_c_7363_n ) capacitor c=0.014626f \
 //x=86.95 //y=7.4 //x2=82.025 //y2=4.44
cc_1798 ( N_VDD_c_1820_p N_noxref_17_c_7363_n ) capacitor c=0.00134165f \
 //x=79.285 //y=7.4 //x2=82.025 //y2=4.44
cc_1799 ( N_VDD_c_1012_n N_noxref_17_c_7363_n ) capacitor c=0.03415f //x=81.03 \
 //y=7.4 //x2=82.025 //y2=4.44
cc_1800 ( N_VDD_M150_noxref_s N_noxref_17_c_7363_n ) capacitor c=6.29527e-19 \
 //x=78.355 //y=5.025 //x2=82.025 //y2=4.44
cc_1801 ( N_VDD_M153_noxref_d N_noxref_17_c_7363_n ) capacitor c=0.0033086f \
 //x=80.105 //y=5.025 //x2=82.025 //y2=4.44
cc_1802 ( N_VDD_c_1015_p N_noxref_17_c_7368_n ) capacitor c=0.00166343f \
 //x=86.95 //y=7.4 //x2=78.555 //y2=4.44
cc_1803 ( N_VDD_c_1825_p N_noxref_17_c_7368_n ) capacitor c=4.53049e-19 \
 //x=78.405 //y=7.4 //x2=78.555 //y2=4.44
cc_1804 ( N_VDD_c_1011_n N_noxref_17_c_7368_n ) capacitor c=0.00910381f \
 //x=77.7 //y=7.4 //x2=78.555 //y2=4.44
cc_1805 ( N_VDD_M150_noxref_s N_noxref_17_c_7368_n ) capacitor c=0.00225389f \
 //x=78.355 //y=5.025 //x2=78.555 //y2=4.44
cc_1806 ( N_VDD_c_1004_n N_noxref_17_c_7301_n ) capacitor c=6.09414e-19 \
 //x=48.47 //y=7.4 //x2=46.99 //y2=2.08
cc_1807 ( N_VDD_c_1015_p N_noxref_17_c_7373_n ) capacitor c=0.00453663f \
 //x=86.95 //y=7.4 //x2=50.495 //y2=5.2
cc_1808 ( N_VDD_c_1378_p N_noxref_17_c_7373_n ) capacitor c=4.48391e-19 \
 //x=50.055 //y=7.4 //x2=50.495 //y2=5.2
cc_1809 ( N_VDD_c_1438_p N_noxref_17_c_7373_n ) capacitor c=4.48391e-19 \
 //x=50.935 //y=7.4 //x2=50.495 //y2=5.2
cc_1810 ( N_VDD_M115_noxref_d N_noxref_17_c_7373_n ) capacitor c=0.0124542f \
 //x=49.995 //y=5.02 //x2=50.495 //y2=5.2
cc_1811 ( N_VDD_c_1004_n N_noxref_17_c_7377_n ) capacitor c=0.00985474f \
 //x=48.47 //y=7.4 //x2=49.785 //y2=5.2
cc_1812 ( N_VDD_M114_noxref_s N_noxref_17_c_7377_n ) capacitor c=0.087833f \
 //x=49.125 //y=5.02 //x2=49.785 //y2=5.2
cc_1813 ( N_VDD_c_1015_p N_noxref_17_c_7379_n ) capacitor c=0.00301575f \
 //x=86.95 //y=7.4 //x2=50.975 //y2=5.2
cc_1814 ( N_VDD_c_1438_p N_noxref_17_c_7379_n ) capacitor c=7.72068e-19 \
 //x=50.935 //y=7.4 //x2=50.975 //y2=5.2
cc_1815 ( N_VDD_M117_noxref_d N_noxref_17_c_7379_n ) capacitor c=0.0158515f \
 //x=50.875 //y=5.02 //x2=50.975 //y2=5.2
cc_1816 ( N_VDD_c_1004_n N_noxref_17_c_7303_n ) capacitor c=0.00151618f \
 //x=48.47 //y=7.4 //x2=51.06 //y2=3.33
cc_1817 ( N_VDD_c_1005_n N_noxref_17_c_7303_n ) capacitor c=0.0433069f \
 //x=51.8 //y=7.4 //x2=51.06 //y2=3.33
cc_1818 ( N_VDD_c_1006_n N_noxref_17_c_7304_n ) capacitor c=6.58823e-19 \
 //x=56.61 //y=7.4 //x2=55.13 //y2=2.08
cc_1819 ( N_VDD_c_1015_p N_noxref_17_c_7385_n ) capacitor c=0.00444892f \
 //x=86.95 //y=7.4 //x2=58.935 //y2=5.155
cc_1820 ( N_VDD_c_1553_p N_noxref_17_c_7385_n ) capacitor c=4.31931e-19 \
 //x=58.495 //y=7.4 //x2=58.935 //y2=5.155
cc_1821 ( N_VDD_c_1474_p N_noxref_17_c_7385_n ) capacitor c=4.31931e-19 \
 //x=59.375 //y=7.4 //x2=58.935 //y2=5.155
cc_1822 ( N_VDD_M125_noxref_d N_noxref_17_c_7385_n ) capacitor c=0.0112985f \
 //x=58.435 //y=5.02 //x2=58.935 //y2=5.155
cc_1823 ( N_VDD_c_1006_n N_noxref_17_c_7389_n ) capacitor c=0.00863585f \
 //x=56.61 //y=7.4 //x2=58.225 //y2=5.155
cc_1824 ( N_VDD_M124_noxref_s N_noxref_17_c_7389_n ) capacitor c=0.0831083f \
 //x=57.565 //y=5.02 //x2=58.225 //y2=5.155
cc_1825 ( N_VDD_c_1015_p N_noxref_17_c_7391_n ) capacitor c=0.0044221f \
 //x=86.95 //y=7.4 //x2=59.815 //y2=5.155
cc_1826 ( N_VDD_c_1474_p N_noxref_17_c_7391_n ) capacitor c=4.31931e-19 \
 //x=59.375 //y=7.4 //x2=59.815 //y2=5.155
cc_1827 ( N_VDD_c_1688_p N_noxref_17_c_7391_n ) capacitor c=4.31931e-19 \
 //x=60.255 //y=7.4 //x2=59.815 //y2=5.155
cc_1828 ( N_VDD_M127_noxref_d N_noxref_17_c_7391_n ) capacitor c=0.0112985f \
 //x=59.315 //y=5.02 //x2=59.815 //y2=5.155
cc_1829 ( N_VDD_c_1015_p N_noxref_17_c_7395_n ) capacitor c=0.00434174f \
 //x=86.95 //y=7.4 //x2=60.595 //y2=5.155
cc_1830 ( N_VDD_c_1688_p N_noxref_17_c_7395_n ) capacitor c=7.46626e-19 \
 //x=60.255 //y=7.4 //x2=60.595 //y2=5.155
cc_1831 ( N_VDD_c_1554_p N_noxref_17_c_7395_n ) capacitor c=0.00198565f \
 //x=61.25 //y=7.4 //x2=60.595 //y2=5.155
cc_1832 ( N_VDD_M129_noxref_d N_noxref_17_c_7395_n ) capacitor c=0.0112985f \
 //x=60.195 //y=5.02 //x2=60.595 //y2=5.155
cc_1833 ( N_VDD_c_1007_n N_noxref_17_c_7399_n ) capacitor c=0.0426864f \
 //x=61.42 //y=7.4 //x2=60.68 //y2=3.33
cc_1834 ( N_VDD_c_1015_p N_noxref_17_c_7306_n ) capacitor c=0.00125279f \
 //x=86.95 //y=7.4 //x2=62.53 //y2=2.08
cc_1835 ( N_VDD_c_1556_p N_noxref_17_c_7306_n ) capacitor c=2.87256e-19 \
 //x=63.005 //y=7.4 //x2=62.53 //y2=2.08
cc_1836 ( N_VDD_c_1007_n N_noxref_17_c_7306_n ) capacitor c=0.0134208f \
 //x=61.42 //y=7.4 //x2=62.53 //y2=2.08
cc_1837 ( N_VDD_c_1015_p N_noxref_17_c_7403_n ) capacitor c=0.00453663f \
 //x=86.95 //y=7.4 //x2=63.445 //y2=5.2
cc_1838 ( N_VDD_c_1556_p N_noxref_17_c_7403_n ) capacitor c=4.48391e-19 \
 //x=63.005 //y=7.4 //x2=63.445 //y2=5.2
cc_1839 ( N_VDD_c_1771_p N_noxref_17_c_7403_n ) capacitor c=4.48391e-19 \
 //x=63.885 //y=7.4 //x2=63.445 //y2=5.2
cc_1840 ( N_VDD_M131_noxref_d N_noxref_17_c_7403_n ) capacitor c=0.0124542f \
 //x=62.945 //y=5.02 //x2=63.445 //y2=5.2
cc_1841 ( N_VDD_c_1007_n N_noxref_17_c_7407_n ) capacitor c=0.00985474f \
 //x=61.42 //y=7.4 //x2=62.735 //y2=5.2
cc_1842 ( N_VDD_M130_noxref_s N_noxref_17_c_7407_n ) capacitor c=0.087833f \
 //x=62.075 //y=5.02 //x2=62.735 //y2=5.2
cc_1843 ( N_VDD_c_1015_p N_noxref_17_c_7409_n ) capacitor c=0.00301575f \
 //x=86.95 //y=7.4 //x2=63.925 //y2=5.2
cc_1844 ( N_VDD_c_1771_p N_noxref_17_c_7409_n ) capacitor c=7.72068e-19 \
 //x=63.885 //y=7.4 //x2=63.925 //y2=5.2
cc_1845 ( N_VDD_M133_noxref_d N_noxref_17_c_7409_n ) capacitor c=0.0158515f \
 //x=63.825 //y=5.02 //x2=63.925 //y2=5.2
cc_1846 ( N_VDD_c_1007_n N_noxref_17_c_7308_n ) capacitor c=0.00151618f \
 //x=61.42 //y=7.4 //x2=64.01 //y2=3.33
cc_1847 ( N_VDD_c_1008_n N_noxref_17_c_7308_n ) capacitor c=0.0428942f \
 //x=64.75 //y=7.4 //x2=64.01 //y2=3.33
cc_1848 ( N_VDD_c_1015_p N_noxref_17_c_7309_n ) capacitor c=9.10347e-19 \
 //x=86.95 //y=7.4 //x2=65.86 //y2=2.08
cc_1849 ( N_VDD_c_1008_n N_noxref_17_c_7309_n ) capacitor c=0.0133749f \
 //x=64.75 //y=7.4 //x2=65.86 //y2=2.08
cc_1850 ( N_VDD_M134_noxref_s N_noxref_17_c_7309_n ) capacitor c=0.0125322f \
 //x=65.705 //y=5.02 //x2=65.86 //y2=2.08
cc_1851 ( N_VDD_c_1015_p N_noxref_17_c_7310_n ) capacitor c=0.00142825f \
 //x=86.95 //y=7.4 //x2=78.44 //y2=2.08
cc_1852 ( N_VDD_c_1011_n N_noxref_17_c_7310_n ) capacitor c=0.0250258f \
 //x=77.7 //y=7.4 //x2=78.44 //y2=2.08
cc_1853 ( N_VDD_c_1012_n N_noxref_17_c_7310_n ) capacitor c=4.17679e-19 \
 //x=81.03 //y=7.4 //x2=78.44 //y2=2.08
cc_1854 ( N_VDD_M150_noxref_s N_noxref_17_c_7310_n ) capacitor c=0.0117177f \
 //x=78.355 //y=5.025 //x2=78.44 //y2=2.08
cc_1855 ( N_VDD_c_1012_n N_noxref_17_c_7313_n ) capacitor c=0.0131686f \
 //x=81.03 //y=7.4 //x2=82.14 //y2=2.08
cc_1856 ( N_VDD_c_1013_n N_noxref_17_c_7313_n ) capacitor c=0.00133861f \
 //x=84.36 //y=7.4 //x2=82.14 //y2=2.08
cc_1857 ( N_VDD_c_1370_p N_noxref_17_M112_noxref_g ) capacitor c=0.00675175f \
 //x=47.305 //y=7.4 //x2=46.73 //y2=6.02
cc_1858 ( N_VDD_M111_noxref_d N_noxref_17_M112_noxref_g ) capacitor \
 c=0.015318f //x=46.365 //y=5.02 //x2=46.73 //y2=6.02
cc_1859 ( N_VDD_c_1370_p N_noxref_17_M113_noxref_g ) capacitor c=0.00675379f \
 //x=47.305 //y=7.4 //x2=47.17 //y2=6.02
cc_1860 ( N_VDD_M113_noxref_d N_noxref_17_M113_noxref_g ) capacitor \
 c=0.0394719f //x=47.245 //y=5.02 //x2=47.17 //y2=6.02
cc_1861 ( N_VDD_c_1612_p N_noxref_17_M122_noxref_g ) capacitor c=0.00675175f \
 //x=55.445 //y=7.4 //x2=54.87 //y2=6.02
cc_1862 ( N_VDD_M121_noxref_d N_noxref_17_M122_noxref_g ) capacitor \
 c=0.015318f //x=54.505 //y=5.02 //x2=54.87 //y2=6.02
cc_1863 ( N_VDD_c_1612_p N_noxref_17_M123_noxref_g ) capacitor c=0.00675379f \
 //x=55.445 //y=7.4 //x2=55.31 //y2=6.02
cc_1864 ( N_VDD_M123_noxref_d N_noxref_17_M123_noxref_g ) capacitor \
 c=0.0394719f //x=55.385 //y=5.02 //x2=55.31 //y2=6.02
cc_1865 ( N_VDD_c_1556_p N_noxref_17_M130_noxref_g ) capacitor c=0.00726866f \
 //x=63.005 //y=7.4 //x2=62.43 //y2=6.02
cc_1866 ( N_VDD_M130_noxref_s N_noxref_17_M130_noxref_g ) capacitor \
 c=0.054195f //x=62.075 //y=5.02 //x2=62.43 //y2=6.02
cc_1867 ( N_VDD_c_1556_p N_noxref_17_M131_noxref_g ) capacitor c=0.00672952f \
 //x=63.005 //y=7.4 //x2=62.87 //y2=6.02
cc_1868 ( N_VDD_M131_noxref_d N_noxref_17_M131_noxref_g ) capacitor \
 c=0.015318f //x=62.945 //y=5.02 //x2=62.87 //y2=6.02
cc_1869 ( N_VDD_c_1559_p N_noxref_17_M134_noxref_g ) capacitor c=0.00749687f \
 //x=66.635 //y=7.4 //x2=66.06 //y2=6.02
cc_1870 ( N_VDD_M134_noxref_s N_noxref_17_M134_noxref_g ) capacitor \
 c=0.0477201f //x=65.705 //y=5.02 //x2=66.06 //y2=6.02
cc_1871 ( N_VDD_c_1559_p N_noxref_17_M135_noxref_g ) capacitor c=0.00675175f \
 //x=66.635 //y=7.4 //x2=66.5 //y2=6.02
cc_1872 ( N_VDD_M135_noxref_d N_noxref_17_M135_noxref_g ) capacitor \
 c=0.015318f //x=66.575 //y=5.02 //x2=66.5 //y2=6.02
cc_1873 ( N_VDD_c_1820_p N_noxref_17_M150_noxref_g ) capacitor c=0.00754867f \
 //x=79.285 //y=7.4 //x2=78.71 //y2=6.025
cc_1874 ( N_VDD_c_1011_n N_noxref_17_M150_noxref_g ) capacitor c=0.00684066f \
 //x=77.7 //y=7.4 //x2=78.71 //y2=6.025
cc_1875 ( N_VDD_M150_noxref_s N_noxref_17_M150_noxref_g ) capacitor \
 c=0.0547553f //x=78.355 //y=5.025 //x2=78.71 //y2=6.025
cc_1876 ( N_VDD_c_1820_p N_noxref_17_M151_noxref_g ) capacitor c=0.00678153f \
 //x=79.285 //y=7.4 //x2=79.15 //y2=6.025
cc_1877 ( N_VDD_M151_noxref_d N_noxref_17_M151_noxref_g ) capacitor \
 c=0.015501f //x=79.225 //y=5.025 //x2=79.15 //y2=6.025
cc_1878 ( N_VDD_c_1900_p N_noxref_17_M154_noxref_g ) capacitor c=0.00513227f \
 //x=84.19 //y=7.4 //x2=82.03 //y2=6.025
cc_1879 ( N_VDD_c_1012_n N_noxref_17_M154_noxref_g ) capacitor c=0.00316281f \
 //x=81.03 //y=7.4 //x2=82.03 //y2=6.025
cc_1880 ( N_VDD_c_1900_p N_noxref_17_M155_noxref_g ) capacitor c=0.00512552f \
 //x=84.19 //y=7.4 //x2=82.47 //y2=6.025
cc_1881 ( N_VDD_c_1008_n N_noxref_17_c_7447_n ) capacitor c=0.00757682f \
 //x=64.75 //y=7.4 //x2=66.135 //y2=4.79
cc_1882 ( N_VDD_M134_noxref_s N_noxref_17_c_7447_n ) capacitor c=0.00444914f \
 //x=65.705 //y=5.02 //x2=66.135 //y2=4.79
cc_1883 ( N_VDD_c_1011_n N_noxref_17_c_7449_n ) capacitor c=0.0110236f \
 //x=77.7 //y=7.4 //x2=78.785 //y2=4.795
cc_1884 ( N_VDD_M150_noxref_s N_noxref_17_c_7449_n ) capacitor c=0.00628155f \
 //x=78.355 //y=5.025 //x2=78.785 //y2=4.795
cc_1885 ( N_VDD_c_1007_n N_noxref_17_c_7451_n ) capacitor c=0.0154093f \
 //x=61.42 //y=7.4 //x2=62.53 //y2=4.7
cc_1886 ( N_VDD_c_1012_n N_noxref_17_c_7452_n ) capacitor c=0.0115029f \
 //x=81.03 //y=7.4 //x2=82.14 //y2=4.705
cc_1887 ( N_VDD_c_1015_p N_noxref_17_M114_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=49.555 //y2=5.02
cc_1888 ( N_VDD_c_1378_p N_noxref_17_M114_noxref_d ) capacitor c=0.0140317f \
 //x=50.055 //y=7.4 //x2=49.555 //y2=5.02
cc_1889 ( N_VDD_c_1005_n N_noxref_17_M114_noxref_d ) capacitor c=6.94454e-19 \
 //x=51.8 //y=7.4 //x2=49.555 //y2=5.02
cc_1890 ( N_VDD_M115_noxref_d N_noxref_17_M114_noxref_d ) capacitor \
 c=0.0664752f //x=49.995 //y=5.02 //x2=49.555 //y2=5.02
cc_1891 ( N_VDD_c_1015_p N_noxref_17_M116_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=50.435 //y2=5.02
cc_1892 ( N_VDD_c_1438_p N_noxref_17_M116_noxref_d ) capacitor c=0.0140317f \
 //x=50.935 //y=7.4 //x2=50.435 //y2=5.02
cc_1893 ( N_VDD_c_1005_n N_noxref_17_M116_noxref_d ) capacitor c=0.0120541f \
 //x=51.8 //y=7.4 //x2=50.435 //y2=5.02
cc_1894 ( N_VDD_M114_noxref_s N_noxref_17_M116_noxref_d ) capacitor \
 c=0.00111971f //x=49.125 //y=5.02 //x2=50.435 //y2=5.02
cc_1895 ( N_VDD_M115_noxref_d N_noxref_17_M116_noxref_d ) capacitor \
 c=0.0664752f //x=49.995 //y=5.02 //x2=50.435 //y2=5.02
cc_1896 ( N_VDD_M117_noxref_d N_noxref_17_M116_noxref_d ) capacitor \
 c=0.0664752f //x=50.875 //y=5.02 //x2=50.435 //y2=5.02
cc_1897 ( N_VDD_M118_noxref_s N_noxref_17_M116_noxref_d ) capacitor \
 c=3.73257e-19 //x=52.755 //y=5.02 //x2=50.435 //y2=5.02
cc_1898 ( N_VDD_c_1015_p N_noxref_17_M124_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=57.995 //y2=5.02
cc_1899 ( N_VDD_c_1553_p N_noxref_17_M124_noxref_d ) capacitor c=0.014035f \
 //x=58.495 //y=7.4 //x2=57.995 //y2=5.02
cc_1900 ( N_VDD_M125_noxref_d N_noxref_17_M124_noxref_d ) capacitor \
 c=0.0664752f //x=58.435 //y=5.02 //x2=57.995 //y2=5.02
cc_1901 ( N_VDD_c_1015_p N_noxref_17_M126_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=58.875 //y2=5.02
cc_1902 ( N_VDD_c_1474_p N_noxref_17_M126_noxref_d ) capacitor c=0.014035f \
 //x=59.375 //y=7.4 //x2=58.875 //y2=5.02
cc_1903 ( N_VDD_c_1007_n N_noxref_17_M126_noxref_d ) capacitor c=4.9285e-19 \
 //x=61.42 //y=7.4 //x2=58.875 //y2=5.02
cc_1904 ( N_VDD_M124_noxref_s N_noxref_17_M126_noxref_d ) capacitor \
 c=0.00130656f //x=57.565 //y=5.02 //x2=58.875 //y2=5.02
cc_1905 ( N_VDD_M125_noxref_d N_noxref_17_M126_noxref_d ) capacitor \
 c=0.0664752f //x=58.435 //y=5.02 //x2=58.875 //y2=5.02
cc_1906 ( N_VDD_M127_noxref_d N_noxref_17_M126_noxref_d ) capacitor \
 c=0.0664752f //x=59.315 //y=5.02 //x2=58.875 //y2=5.02
cc_1907 ( N_VDD_c_1015_p N_noxref_17_M128_noxref_d ) capacitor c=0.00275235f \
 //x=86.95 //y=7.4 //x2=59.755 //y2=5.02
cc_1908 ( N_VDD_c_1688_p N_noxref_17_M128_noxref_d ) capacitor c=0.014035f \
 //x=60.255 //y=7.4 //x2=59.755 //y2=5.02
cc_1909 ( N_VDD_c_1007_n N_noxref_17_M128_noxref_d ) capacitor c=0.00939849f \
 //x=61.42 //y=7.4 //x2=59.755 //y2=5.02
cc_1910 ( N_VDD_M127_noxref_d N_noxref_17_M128_noxref_d ) capacitor \
 c=0.0664752f //x=59.315 //y=5.02 //x2=59.755 //y2=5.02
cc_1911 ( N_VDD_M129_noxref_d N_noxref_17_M128_noxref_d ) capacitor \
 c=0.0664752f //x=60.195 //y=5.02 //x2=59.755 //y2=5.02
cc_1912 ( N_VDD_M130_noxref_s N_noxref_17_M128_noxref_d ) capacitor \
 c=4.52683e-19 //x=62.075 //y=5.02 //x2=59.755 //y2=5.02
cc_1913 ( N_VDD_c_1015_p N_noxref_17_M130_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=62.505 //y2=5.02
cc_1914 ( N_VDD_c_1556_p N_noxref_17_M130_noxref_d ) capacitor c=0.0140317f \
 //x=63.005 //y=7.4 //x2=62.505 //y2=5.02
cc_1915 ( N_VDD_c_1008_n N_noxref_17_M130_noxref_d ) capacitor c=6.94454e-19 \
 //x=64.75 //y=7.4 //x2=62.505 //y2=5.02
cc_1916 ( N_VDD_M131_noxref_d N_noxref_17_M130_noxref_d ) capacitor \
 c=0.0664752f //x=62.945 //y=5.02 //x2=62.505 //y2=5.02
cc_1917 ( N_VDD_c_1015_p N_noxref_17_M132_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=63.385 //y2=5.02
cc_1918 ( N_VDD_c_1771_p N_noxref_17_M132_noxref_d ) capacitor c=0.0140317f \
 //x=63.885 //y=7.4 //x2=63.385 //y2=5.02
cc_1919 ( N_VDD_c_1008_n N_noxref_17_M132_noxref_d ) capacitor c=0.0120541f \
 //x=64.75 //y=7.4 //x2=63.385 //y2=5.02
cc_1920 ( N_VDD_M130_noxref_s N_noxref_17_M132_noxref_d ) capacitor \
 c=0.00111971f //x=62.075 //y=5.02 //x2=63.385 //y2=5.02
cc_1921 ( N_VDD_M131_noxref_d N_noxref_17_M132_noxref_d ) capacitor \
 c=0.0664752f //x=62.945 //y=5.02 //x2=63.385 //y2=5.02
cc_1922 ( N_VDD_M133_noxref_d N_noxref_17_M132_noxref_d ) capacitor \
 c=0.0664752f //x=63.825 //y=5.02 //x2=63.385 //y2=5.02
cc_1923 ( N_VDD_M134_noxref_s N_noxref_17_M132_noxref_d ) capacitor \
 c=3.73257e-19 //x=65.705 //y=5.02 //x2=63.385 //y2=5.02
cc_1924 ( N_VDD_c_1015_p N_noxref_18_c_8076_n ) capacitor c=0.0146576f \
 //x=86.95 //y=7.4 //x2=76.845 //y2=3.7
cc_1925 ( N_VDD_c_1015_p N_noxref_18_c_8077_n ) capacitor c=0.010327f \
 //x=86.95 //y=7.4 //x2=79.435 //y2=3.7
cc_1926 ( N_VDD_c_1011_n N_noxref_18_c_8077_n ) capacitor c=0.0109524f \
 //x=77.7 //y=7.4 //x2=79.435 //y2=3.7
cc_1927 ( N_VDD_c_1015_p N_noxref_18_c_8079_n ) capacitor c=0.00154061f \
 //x=86.95 //y=7.4 //x2=77.075 //y2=3.7
cc_1928 ( N_VDD_M149_noxref_d N_noxref_18_c_8079_n ) capacitor c=4.05358e-19 \
 //x=76.775 //y=5.02 //x2=77.075 //y2=3.7
cc_1929 ( N_VDD_c_1015_p N_noxref_18_c_8064_n ) capacitor c=0.0151699f \
 //x=86.95 //y=7.4 //x2=86.095 //y2=4.07
cc_1930 ( N_VDD_c_993_n N_noxref_18_c_8064_n ) capacitor c=4.075e-19 //x=86.95 \
 //y=7.4 //x2=86.095 //y2=4.07
cc_1931 ( N_VDD_c_1012_n N_noxref_18_c_8064_n ) capacitor c=0.0150456f \
 //x=81.03 //y=7.4 //x2=86.095 //y2=4.07
cc_1932 ( N_VDD_c_1013_n N_noxref_18_c_8064_n ) capacitor c=0.0225025f \
 //x=84.36 //y=7.4 //x2=86.095 //y2=4.07
cc_1933 ( N_VDD_c_1012_n N_noxref_18_c_8085_n ) capacitor c=5.4458e-19 \
 //x=81.03 //y=7.4 //x2=79.665 //y2=4.07
cc_1934 ( N_VDD_c_1010_n N_noxref_18_c_8065_n ) capacitor c=8.79202e-19 \
 //x=74.37 //y=7.4 //x2=72.89 //y2=2.08
cc_1935 ( N_VDD_c_1015_p N_noxref_18_c_8087_n ) capacitor c=0.00459955f \
 //x=86.95 //y=7.4 //x2=76.395 //y2=5.2
cc_1936 ( N_VDD_c_1717_p N_noxref_18_c_8087_n ) capacitor c=4.48705e-19 \
 //x=75.955 //y=7.4 //x2=76.395 //y2=5.2
cc_1937 ( N_VDD_c_1780_p N_noxref_18_c_8087_n ) capacitor c=4.48693e-19 \
 //x=76.835 //y=7.4 //x2=76.395 //y2=5.2
cc_1938 ( N_VDD_M147_noxref_d N_noxref_18_c_8087_n ) capacitor c=0.01269f \
 //x=75.895 //y=5.02 //x2=76.395 //y2=5.2
cc_1939 ( N_VDD_c_1010_n N_noxref_18_c_8091_n ) capacitor c=0.00985474f \
 //x=74.37 //y=7.4 //x2=75.685 //y2=5.2
cc_1940 ( N_VDD_M146_noxref_s N_noxref_18_c_8091_n ) capacitor c=0.087833f \
 //x=75.025 //y=5.02 //x2=75.685 //y2=5.2
cc_1941 ( N_VDD_c_1015_p N_noxref_18_c_8093_n ) capacitor c=0.00311875f \
 //x=86.95 //y=7.4 //x2=76.875 //y2=5.2
cc_1942 ( N_VDD_c_1780_p N_noxref_18_c_8093_n ) capacitor c=7.21492e-19 \
 //x=76.835 //y=7.4 //x2=76.875 //y2=5.2
cc_1943 ( N_VDD_M149_noxref_d N_noxref_18_c_8093_n ) capacitor c=0.0163364f \
 //x=76.775 //y=5.02 //x2=76.875 //y2=5.2
cc_1944 ( N_VDD_M150_noxref_s N_noxref_18_c_8093_n ) capacitor c=5.34061e-19 \
 //x=78.355 //y=5.025 //x2=76.875 //y2=5.2
cc_1945 ( N_VDD_c_1010_n N_noxref_18_c_8067_n ) capacitor c=0.00151618f \
 //x=74.37 //y=7.4 //x2=76.96 //y2=3.7
cc_1946 ( N_VDD_c_1011_n N_noxref_18_c_8067_n ) capacitor c=0.0449408f \
 //x=77.7 //y=7.4 //x2=76.96 //y2=3.7
cc_1947 ( N_VDD_c_1012_n N_noxref_18_c_8099_n ) capacitor c=0.00491684f \
 //x=81.03 //y=7.4 //x2=79.55 //y2=4.54
cc_1948 ( N_VDD_c_1011_n N_noxref_18_c_8068_n ) capacitor c=0.00113585f \
 //x=77.7 //y=7.4 //x2=79.55 //y2=2.08
cc_1949 ( N_VDD_c_1012_n N_noxref_18_c_8068_n ) capacitor c=0.0042566f \
 //x=81.03 //y=7.4 //x2=79.55 //y2=2.08
cc_1950 ( N_VDD_c_993_n N_noxref_18_c_8070_n ) capacitor c=6.69172e-19 \
 //x=86.95 //y=7.4 //x2=86.21 //y2=2.08
cc_1951 ( N_VDD_c_1013_n N_noxref_18_c_8070_n ) capacitor c=0.00116377f \
 //x=84.36 //y=7.4 //x2=86.21 //y2=2.08
cc_1952 ( N_VDD_c_1755_p N_noxref_18_M144_noxref_g ) capacitor c=0.00675175f \
 //x=73.205 //y=7.4 //x2=72.63 //y2=6.02
cc_1953 ( N_VDD_M143_noxref_d N_noxref_18_M144_noxref_g ) capacitor \
 c=0.015318f //x=72.265 //y=5.02 //x2=72.63 //y2=6.02
cc_1954 ( N_VDD_c_1755_p N_noxref_18_M145_noxref_g ) capacitor c=0.00675379f \
 //x=73.205 //y=7.4 //x2=73.07 //y2=6.02
cc_1955 ( N_VDD_M145_noxref_d N_noxref_18_M145_noxref_g ) capacitor \
 c=0.0394719f //x=73.145 //y=5.02 //x2=73.07 //y2=6.02
cc_1956 ( N_VDD_c_1978_p N_noxref_18_M152_noxref_g ) capacitor c=0.0067918f \
 //x=80.165 //y=7.4 //x2=79.59 //y2=6.025
cc_1957 ( N_VDD_M151_noxref_d N_noxref_18_M152_noxref_g ) capacitor \
 c=0.015526f //x=79.225 //y=5.025 //x2=79.59 //y2=6.025
cc_1958 ( N_VDD_c_1978_p N_noxref_18_M153_noxref_g ) capacitor c=0.00754867f \
 //x=80.165 //y=7.4 //x2=80.03 //y2=6.025
cc_1959 ( N_VDD_M153_noxref_d N_noxref_18_M153_noxref_g ) capacitor \
 c=0.0537676f //x=80.105 //y=5.025 //x2=80.03 //y2=6.025
cc_1960 ( N_VDD_c_993_n N_noxref_18_M160_noxref_g ) capacitor c=0.00513565f \
 //x=86.95 //y=7.4 //x2=86.25 //y2=6.025
cc_1961 ( N_VDD_c_993_n N_noxref_18_M161_noxref_g ) capacitor c=0.0309137f \
 //x=86.95 //y=7.4 //x2=86.69 //y2=6.025
cc_1962 ( N_VDD_c_1012_n N_noxref_18_c_8114_n ) capacitor c=0.00985898f \
 //x=81.03 //y=7.4 //x2=79.955 //y2=4.795
cc_1963 ( N_VDD_c_1012_n N_noxref_18_c_8115_n ) capacitor c=2.76772e-19 \
 //x=81.03 //y=7.4 //x2=79.59 //y2=4.705
cc_1964 ( N_VDD_c_1015_p N_noxref_18_M146_noxref_d ) capacitor c=0.0028472f \
 //x=86.95 //y=7.4 //x2=75.455 //y2=5.02
cc_1965 ( N_VDD_c_1717_p N_noxref_18_M146_noxref_d ) capacitor c=0.014096f \
 //x=75.955 //y=7.4 //x2=75.455 //y2=5.02
cc_1966 ( N_VDD_c_1011_n N_noxref_18_M146_noxref_d ) capacitor c=6.94454e-19 \
 //x=77.7 //y=7.4 //x2=75.455 //y2=5.02
cc_1967 ( N_VDD_M147_noxref_d N_noxref_18_M146_noxref_d ) capacitor \
 c=0.0664752f //x=75.895 //y=5.02 //x2=75.455 //y2=5.02
cc_1968 ( N_VDD_c_1015_p N_noxref_18_M148_noxref_d ) capacitor c=0.00294217f \
 //x=86.95 //y=7.4 //x2=76.335 //y2=5.02
cc_1969 ( N_VDD_c_1780_p N_noxref_18_M148_noxref_d ) capacitor c=0.0138379f \
 //x=76.835 //y=7.4 //x2=76.335 //y2=5.02
cc_1970 ( N_VDD_c_1011_n N_noxref_18_M148_noxref_d ) capacitor c=0.0120518f \
 //x=77.7 //y=7.4 //x2=76.335 //y2=5.02
cc_1971 ( N_VDD_M146_noxref_s N_noxref_18_M148_noxref_d ) capacitor \
 c=0.00111971f //x=75.025 //y=5.02 //x2=76.335 //y2=5.02
cc_1972 ( N_VDD_M147_noxref_d N_noxref_18_M148_noxref_d ) capacitor \
 c=0.0664752f //x=75.895 //y=5.02 //x2=76.335 //y2=5.02
cc_1973 ( N_VDD_M149_noxref_d N_noxref_18_M148_noxref_d ) capacitor \
 c=0.0664752f //x=76.775 //y=5.02 //x2=76.335 //y2=5.02
cc_1974 ( N_VDD_M150_noxref_s N_noxref_18_M148_noxref_d ) capacitor \
 c=4.54243e-19 //x=78.355 //y=5.025 //x2=76.335 //y2=5.02
cc_1975 ( N_VDD_c_1015_p N_noxref_19_c_8424_n ) capacitor c=0.0206457f \
 //x=86.95 //y=7.4 //x2=81.695 //y2=5.21
cc_1976 ( N_VDD_c_1978_p N_noxref_19_c_8424_n ) capacitor c=0.00213763f \
 //x=80.165 //y=7.4 //x2=81.695 //y2=5.21
cc_1977 ( N_VDD_c_1999_p N_noxref_19_c_8424_n ) capacitor c=0.003172f \
 //x=80.86 //y=7.4 //x2=81.695 //y2=5.21
cc_1978 ( N_VDD_c_1900_p N_noxref_19_c_8424_n ) capacitor c=0.00424633f \
 //x=84.19 //y=7.4 //x2=81.695 //y2=5.21
cc_1979 ( N_VDD_c_1012_n N_noxref_19_c_8424_n ) capacitor c=0.0430305f \
 //x=81.03 //y=7.4 //x2=81.695 //y2=5.21
cc_1980 ( N_VDD_M153_noxref_d N_noxref_19_c_8424_n ) capacitor c=0.0197937f \
 //x=80.105 //y=5.025 //x2=81.695 //y2=5.21
cc_1981 ( N_VDD_c_1015_p N_noxref_19_c_8430_n ) capacitor c=0.00274812f \
 //x=86.95 //y=7.4 //x2=79.925 //y2=5.21
cc_1982 ( N_VDD_c_1978_p N_noxref_19_c_8430_n ) capacitor c=0.00107267f \
 //x=80.165 //y=7.4 //x2=79.925 //y2=5.21
cc_1983 ( N_VDD_c_1011_n N_noxref_19_c_8430_n ) capacitor c=2.89592e-19 \
 //x=77.7 //y=7.4 //x2=79.925 //y2=5.21
cc_1984 ( N_VDD_c_1012_n N_noxref_19_c_8430_n ) capacitor c=3.35418e-19 \
 //x=81.03 //y=7.4 //x2=79.925 //y2=5.21
cc_1985 ( N_VDD_M153_noxref_d N_noxref_19_c_8430_n ) capacitor c=6.02701e-19 \
 //x=80.105 //y=5.025 //x2=79.925 //y2=5.21
cc_1986 ( N_VDD_c_1015_p N_noxref_19_c_8435_n ) capacitor c=0.00453889f \
 //x=86.95 //y=7.4 //x2=79.725 //y2=5.21
cc_1987 ( N_VDD_c_1820_p N_noxref_19_c_8435_n ) capacitor c=4.52207e-19 \
 //x=79.285 //y=7.4 //x2=79.725 //y2=5.21
cc_1988 ( N_VDD_c_1978_p N_noxref_19_c_8435_n ) capacitor c=4.11408e-19 \
 //x=80.165 //y=7.4 //x2=79.725 //y2=5.21
cc_1989 ( N_VDD_M151_noxref_d N_noxref_19_c_8435_n ) capacitor c=0.0127968f \
 //x=79.225 //y=5.025 //x2=79.725 //y2=5.21
cc_1990 ( N_VDD_c_1011_n N_noxref_19_c_8439_n ) capacitor c=0.00914165f \
 //x=77.7 //y=7.4 //x2=79.015 //y2=5.21
cc_1991 ( N_VDD_M150_noxref_s N_noxref_19_c_8439_n ) capacitor c=0.0872987f \
 //x=78.355 //y=5.025 //x2=79.015 //y2=5.21
cc_1992 ( N_VDD_c_1011_n N_noxref_19_c_8441_n ) capacitor c=6.3991e-19 \
 //x=77.7 //y=7.4 //x2=79.81 //y2=5.295
cc_1993 ( N_VDD_c_1012_n N_noxref_19_c_8441_n ) capacitor c=0.00985441f \
 //x=81.03 //y=7.4 //x2=79.81 //y2=5.295
cc_1994 ( N_VDD_M153_noxref_d N_noxref_19_c_8441_n ) capacitor c=0.0873334f \
 //x=80.105 //y=5.025 //x2=79.81 //y2=5.295
cc_1995 ( N_VDD_c_1012_n N_noxref_19_c_8444_n ) capacitor c=0.0674112f \
 //x=81.03 //y=7.4 //x2=81.81 //y2=5.21
cc_1996 ( N_VDD_M153_noxref_d N_noxref_19_c_8444_n ) capacitor c=0.00235009f \
 //x=80.105 //y=5.025 //x2=81.81 //y2=5.21
cc_1997 ( N_VDD_c_1015_p N_noxref_19_c_8446_n ) capacitor c=0.0296174f \
 //x=86.95 //y=7.4 //x2=81.895 //y2=6.91
cc_1998 ( N_VDD_c_1900_p N_noxref_19_c_8446_n ) capacitor c=0.109938f \
 //x=84.19 //y=7.4 //x2=81.895 //y2=6.91
cc_1999 ( N_VDD_c_1015_p N_noxref_19_M150_noxref_d ) capacitor c=0.00291898f \
 //x=86.95 //y=7.4 //x2=78.785 //y2=5.025
cc_2000 ( N_VDD_c_1820_p N_noxref_19_M150_noxref_d ) capacitor c=0.0137097f \
 //x=79.285 //y=7.4 //x2=78.785 //y2=5.025
cc_2001 ( N_VDD_M151_noxref_d N_noxref_19_M150_noxref_d ) capacitor \
 c=0.067695f //x=79.225 //y=5.025 //x2=78.785 //y2=5.025
cc_2002 ( N_VDD_M153_noxref_d N_noxref_19_M150_noxref_d ) capacitor \
 c=0.00105738f //x=80.105 //y=5.025 //x2=78.785 //y2=5.025
cc_2003 ( N_VDD_c_1015_p N_noxref_19_M152_noxref_d ) capacitor c=0.00241371f \
 //x=86.95 //y=7.4 //x2=79.665 //y2=5.025
cc_2004 ( N_VDD_c_1978_p N_noxref_19_M152_noxref_d ) capacitor c=0.01268f \
 //x=80.165 //y=7.4 //x2=79.665 //y2=5.025
cc_2005 ( N_VDD_M150_noxref_s N_noxref_19_M152_noxref_d ) capacitor \
 c=0.00103189f //x=78.355 //y=5.025 //x2=79.665 //y2=5.025
cc_2006 ( N_VDD_M151_noxref_d N_noxref_19_M152_noxref_d ) capacitor \
 c=0.0653408f //x=79.225 //y=5.025 //x2=79.665 //y2=5.025
cc_2007 ( N_VDD_c_1012_n N_noxref_19_M155_noxref_d ) capacitor c=8.96067e-19 \
 //x=81.03 //y=7.4 //x2=82.545 //y2=5.025
cc_2008 ( N_VDD_c_1013_n N_noxref_19_M155_noxref_d ) capacitor c=8.88629e-19 \
 //x=84.36 //y=7.4 //x2=82.545 //y2=5.025
cc_2009 ( N_VDD_c_1013_n N_noxref_19_M157_noxref_d ) capacitor c=0.0575594f \
 //x=84.36 //y=7.4 //x2=83.425 //y2=5.025
cc_2010 ( N_VDD_c_999_n N_noxref_20_c_8516_n ) capacitor c=0.00315988f \
 //x=25.9 //y=7.4 //x2=83.505 //y2=2.96
cc_2011 ( N_VDD_c_998_n N_noxref_20_c_8538_n ) capacitor c=6.35146e-19 \
 //x=22.57 //y=7.4 //x2=21.09 //y2=2.08
cc_2012 ( N_VDD_c_1015_p N_noxref_20_c_8560_n ) capacitor c=0.00453663f \
 //x=86.95 //y=7.4 //x2=24.595 //y2=5.2
cc_2013 ( N_VDD_c_1185_p N_noxref_20_c_8560_n ) capacitor c=4.48391e-19 \
 //x=24.155 //y=7.4 //x2=24.595 //y2=5.2
cc_2014 ( N_VDD_c_1202_p N_noxref_20_c_8560_n ) capacitor c=4.48391e-19 \
 //x=25.035 //y=7.4 //x2=24.595 //y2=5.2
cc_2015 ( N_VDD_M83_noxref_d N_noxref_20_c_8560_n ) capacitor c=0.0124542f \
 //x=24.095 //y=5.02 //x2=24.595 //y2=5.2
cc_2016 ( N_VDD_c_998_n N_noxref_20_c_8564_n ) capacitor c=0.00985474f \
 //x=22.57 //y=7.4 //x2=23.885 //y2=5.2
cc_2017 ( N_VDD_M82_noxref_s N_noxref_20_c_8564_n ) capacitor c=0.087833f \
 //x=23.225 //y=5.02 //x2=23.885 //y2=5.2
cc_2018 ( N_VDD_c_1015_p N_noxref_20_c_8566_n ) capacitor c=0.00301575f \
 //x=86.95 //y=7.4 //x2=25.075 //y2=5.2
cc_2019 ( N_VDD_c_1202_p N_noxref_20_c_8566_n ) capacitor c=7.72068e-19 \
 //x=25.035 //y=7.4 //x2=25.075 //y2=5.2
cc_2020 ( N_VDD_M85_noxref_d N_noxref_20_c_8566_n ) capacitor c=0.0158515f \
 //x=24.975 //y=5.02 //x2=25.075 //y2=5.2
cc_2021 ( N_VDD_c_998_n N_noxref_20_c_8540_n ) capacitor c=0.00151618f \
 //x=22.57 //y=7.4 //x2=25.16 //y2=2.96
cc_2022 ( N_VDD_c_999_n N_noxref_20_c_8540_n ) capacitor c=0.0433069f //x=25.9 \
 //y=7.4 //x2=25.16 //y2=2.96
cc_2023 ( N_VDD_c_1012_n N_noxref_20_c_8541_n ) capacitor c=7.57423e-19 \
 //x=81.03 //y=7.4 //x2=83.62 //y2=2.08
cc_2024 ( N_VDD_c_1013_n N_noxref_20_c_8541_n ) capacitor c=0.0263215f \
 //x=84.36 //y=7.4 //x2=83.62 //y2=2.08
cc_2025 ( N_VDD_c_1013_n N_noxref_20_c_8543_n ) capacitor c=0.0263871f \
 //x=84.36 //y=7.4 //x2=85.1 //y2=2.08
cc_2026 ( N_VDD_c_1177_p N_noxref_20_M80_noxref_g ) capacitor c=0.00675175f \
 //x=21.405 //y=7.4 //x2=20.83 //y2=6.02
cc_2027 ( N_VDD_M79_noxref_d N_noxref_20_M80_noxref_g ) capacitor c=0.015318f \
 //x=20.465 //y=5.02 //x2=20.83 //y2=6.02
cc_2028 ( N_VDD_c_1177_p N_noxref_20_M81_noxref_g ) capacitor c=0.00675379f \
 //x=21.405 //y=7.4 //x2=21.27 //y2=6.02
cc_2029 ( N_VDD_M81_noxref_d N_noxref_20_M81_noxref_g ) capacitor c=0.0394719f \
 //x=21.345 //y=5.02 //x2=21.27 //y2=6.02
cc_2030 ( N_VDD_c_1900_p N_noxref_20_M156_noxref_g ) capacitor c=0.00512552f \
 //x=84.19 //y=7.4 //x2=82.91 //y2=6.025
cc_2031 ( N_VDD_c_1900_p N_noxref_20_M157_noxref_g ) capacitor c=0.00512552f \
 //x=84.19 //y=7.4 //x2=83.35 //y2=6.025
cc_2032 ( N_VDD_c_1013_n N_noxref_20_M157_noxref_g ) capacitor c=0.010355f \
 //x=84.36 //y=7.4 //x2=83.35 //y2=6.025
cc_2033 ( N_VDD_c_993_n N_noxref_20_M158_noxref_g ) capacitor c=0.00512552f \
 //x=86.95 //y=7.4 //x2=85.37 //y2=6.025
cc_2034 ( N_VDD_c_1013_n N_noxref_20_M158_noxref_g ) capacitor c=0.00767856f \
 //x=84.36 //y=7.4 //x2=85.37 //y2=6.025
cc_2035 ( N_VDD_c_993_n N_noxref_20_M159_noxref_g ) capacitor c=0.00512552f \
 //x=86.95 //y=7.4 //x2=85.81 //y2=6.025
cc_2036 ( N_VDD_c_1013_n N_noxref_20_c_8584_n ) capacitor c=0.00803198f \
 //x=84.36 //y=7.4 //x2=83.35 //y2=4.87
cc_2037 ( N_VDD_c_1013_n N_noxref_20_c_8585_n ) capacitor c=0.00803198f \
 //x=84.36 //y=7.4 //x2=85.445 //y2=4.795
cc_2038 ( N_VDD_c_1015_p N_noxref_20_M82_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=23.655 //y2=5.02
cc_2039 ( N_VDD_c_1185_p N_noxref_20_M82_noxref_d ) capacitor c=0.0140317f \
 //x=24.155 //y=7.4 //x2=23.655 //y2=5.02
cc_2040 ( N_VDD_c_999_n N_noxref_20_M82_noxref_d ) capacitor c=6.94454e-19 \
 //x=25.9 //y=7.4 //x2=23.655 //y2=5.02
cc_2041 ( N_VDD_M83_noxref_d N_noxref_20_M82_noxref_d ) capacitor c=0.0664752f \
 //x=24.095 //y=5.02 //x2=23.655 //y2=5.02
cc_2042 ( N_VDD_c_1015_p N_noxref_20_M84_noxref_d ) capacitor c=0.00275225f \
 //x=86.95 //y=7.4 //x2=24.535 //y2=5.02
cc_2043 ( N_VDD_c_1202_p N_noxref_20_M84_noxref_d ) capacitor c=0.0140317f \
 //x=25.035 //y=7.4 //x2=24.535 //y2=5.02
cc_2044 ( N_VDD_c_999_n N_noxref_20_M84_noxref_d ) capacitor c=0.0120541f \
 //x=25.9 //y=7.4 //x2=24.535 //y2=5.02
cc_2045 ( N_VDD_M82_noxref_s N_noxref_20_M84_noxref_d ) capacitor \
 c=0.00111971f //x=23.225 //y=5.02 //x2=24.535 //y2=5.02
cc_2046 ( N_VDD_M83_noxref_d N_noxref_20_M84_noxref_d ) capacitor c=0.0664752f \
 //x=24.095 //y=5.02 //x2=24.535 //y2=5.02
cc_2047 ( N_VDD_M85_noxref_d N_noxref_20_M84_noxref_d ) capacitor c=0.0664752f \
 //x=24.975 //y=5.02 //x2=24.535 //y2=5.02
cc_2048 ( N_VDD_M86_noxref_s N_noxref_20_M84_noxref_d ) capacitor \
 c=3.73257e-19 //x=26.855 //y=5.02 //x2=24.535 //y2=5.02
cc_2049 ( N_VDD_c_1015_p N_noxref_21_c_9008_n ) capacitor c=0.0212729f \
 //x=86.95 //y=7.4 //x2=85.035 //y2=5.21
cc_2050 ( N_VDD_c_1900_p N_noxref_21_c_9008_n ) capacitor c=0.00386143f \
 //x=84.19 //y=7.4 //x2=85.035 //y2=5.21
cc_2051 ( N_VDD_c_993_n N_noxref_21_c_9008_n ) capacitor c=0.00403412f \
 //x=86.95 //y=7.4 //x2=85.035 //y2=5.21
cc_2052 ( N_VDD_c_1013_n N_noxref_21_c_9008_n ) capacitor c=0.0473381f \
 //x=84.36 //y=7.4 //x2=85.035 //y2=5.21
cc_2053 ( N_VDD_c_1015_p N_noxref_21_c_9012_n ) capacitor c=0.00264311f \
 //x=86.95 //y=7.4 //x2=83.245 //y2=5.21
cc_2054 ( N_VDD_c_1013_n N_noxref_21_c_9012_n ) capacitor c=6.67754e-19 \
 //x=84.36 //y=7.4 //x2=83.245 //y2=5.21
cc_2055 ( N_VDD_c_1012_n N_noxref_21_c_9014_n ) capacitor c=0.00662411f \
 //x=81.03 //y=7.4 //x2=82.335 //y2=5.21
cc_2056 ( N_VDD_c_1013_n N_noxref_21_c_9015_n ) capacitor c=0.00999961f \
 //x=84.36 //y=7.4 //x2=83.13 //y2=5.295
cc_2057 ( N_VDD_c_993_n N_noxref_21_c_9016_n ) capacitor c=6.48751e-19 \
 //x=86.95 //y=7.4 //x2=85.15 //y2=5.21
cc_2058 ( N_VDD_c_1013_n N_noxref_21_c_9016_n ) capacitor c=0.0664301f \
 //x=84.36 //y=7.4 //x2=85.15 //y2=5.21
cc_2059 ( N_VDD_c_1015_p N_noxref_21_c_9018_n ) capacitor c=0.043423f \
 //x=86.95 //y=7.4 //x2=85.235 //y2=6.91
cc_2060 ( N_VDD_c_993_n N_noxref_21_c_9018_n ) capacitor c=0.108124f //x=86.95 \
 //y=7.4 //x2=85.235 //y2=6.91
cc_2061 ( N_VDD_c_993_n N_noxref_21_M159_noxref_d ) capacitor c=8.96067e-19 \
 //x=86.95 //y=7.4 //x2=85.885 //y2=5.025
cc_2062 ( N_VDD_c_1013_n N_noxref_21_M159_noxref_d ) capacitor c=8.88629e-19 \
 //x=84.36 //y=7.4 //x2=85.885 //y2=5.025
cc_2063 ( N_VDD_c_993_n N_noxref_21_M161_noxref_d ) capacitor c=0.0529764f \
 //x=86.95 //y=7.4 //x2=86.765 //y2=5.025
cc_2064 ( N_VDD_c_993_n QN ) capacitor c=0.0470629f //x=86.95 //y=7.4 \
 //x2=86.95 //y2=2.22
cc_2065 ( N_VDD_c_1013_n QN ) capacitor c=0.00147633f //x=84.36 //y=7.4 \
 //x2=86.95 //y2=2.22
cc_2066 ( N_VDD_c_1013_n N_QN_c_9126_n ) capacitor c=0.00660621f //x=84.36 \
 //y=7.4 //x2=85.675 //y2=5.21
cc_2067 ( N_VDD_c_1015_p N_QN_c_9127_n ) capacitor c=0.00240012f //x=86.95 \
 //y=7.4 //x2=86.865 //y2=5.21
cc_2068 ( N_VDD_c_993_n N_QN_c_9127_n ) capacitor c=0.00136974f //x=86.95 \
 //y=7.4 //x2=86.865 //y2=5.21
cc_2069 ( N_VDD_c_993_n N_QN_M158_noxref_d ) capacitor c=6.67979e-19 //x=86.95 \
 //y=7.4 //x2=85.445 //y2=5.025
cc_2070 ( N_VDD_c_993_n N_QN_M160_noxref_d ) capacitor c=0.0099096f //x=86.95 \
 //y=7.4 //x2=86.325 //y2=5.025
cc_2071 ( N_noxref_3_c_2098_n N_noxref_4_c_2391_n ) capacitor c=0.011463f \
 //x=10.615 //y=3.33 //x2=12.325 //y2=3.33
cc_2072 ( N_noxref_3_M67_noxref_g N_noxref_4_c_2360_n ) capacitor c=0.0169521f \
 //x=11.07 //y=6.02 //x2=11.645 //y2=5.2
cc_2073 ( N_noxref_3_c_2101_n N_noxref_4_c_2364_n ) capacitor c=0.00539951f \
 //x=10.73 //y=2.08 //x2=10.935 //y2=5.2
cc_2074 ( N_noxref_3_M66_noxref_g N_noxref_4_c_2364_n ) capacitor c=0.0177326f \
 //x=10.63 //y=6.02 //x2=10.935 //y2=5.2
cc_2075 ( N_noxref_3_c_2140_n N_noxref_4_c_2364_n ) capacitor c=0.00581252f \
 //x=10.73 //y=4.7 //x2=10.935 //y2=5.2
cc_2076 ( N_noxref_3_c_2128_n N_noxref_4_c_2345_n ) capacitor c=3.52729e-19 \
 //x=8.88 //y=3.33 //x2=12.21 //y2=3.33
cc_2077 ( N_noxref_3_c_2101_n N_noxref_4_c_2345_n ) capacitor c=0.0027152f \
 //x=10.73 //y=2.08 //x2=12.21 //y2=3.33
cc_2078 ( N_noxref_3_M67_noxref_g N_noxref_4_M66_noxref_d ) capacitor \
 c=0.0173476f //x=11.07 //y=6.02 //x2=10.705 //y2=5.02
cc_2079 ( N_noxref_3_c_2093_n N_noxref_5_c_2568_n ) capacitor c=0.146539f \
 //x=8.765 //y=3.33 //x2=5.805 //y2=3.7
cc_2080 ( N_noxref_3_c_2093_n N_noxref_5_c_2569_n ) capacitor c=0.0294746f \
 //x=8.765 //y=3.33 //x2=4.185 //y2=3.7
cc_2081 ( N_noxref_3_c_2099_n N_noxref_5_c_2569_n ) capacitor c=0.00687545f \
 //x=3.33 //y=2.08 //x2=4.185 //y2=3.7
cc_2082 ( N_noxref_3_c_2093_n N_noxref_5_c_2495_n ) capacitor c=0.238435f \
 //x=8.765 //y=3.33 //x2=18.755 //y2=3.7
cc_2083 ( N_noxref_3_c_2098_n N_noxref_5_c_2495_n ) capacitor c=0.175734f \
 //x=10.615 //y=3.33 //x2=18.755 //y2=3.7
cc_2084 ( N_noxref_3_c_2169_p N_noxref_5_c_2495_n ) capacitor c=0.0268386f \
 //x=8.995 //y=3.33 //x2=18.755 //y2=3.7
cc_2085 ( N_noxref_3_c_2128_n N_noxref_5_c_2495_n ) capacitor c=0.0206044f \
 //x=8.88 //y=3.33 //x2=18.755 //y2=3.7
cc_2086 ( N_noxref_3_c_2101_n N_noxref_5_c_2495_n ) capacitor c=0.0205831f \
 //x=10.73 //y=2.08 //x2=18.755 //y2=3.7
cc_2087 ( N_noxref_3_c_2093_n N_noxref_5_c_2576_n ) capacitor c=0.0266966f \
 //x=8.765 //y=3.33 //x2=6.035 //y2=3.7
cc_2088 ( N_noxref_3_M58_noxref_g N_noxref_5_c_2526_n ) capacitor c=0.01736f \
 //x=3.07 //y=6.02 //x2=3.205 //y2=5.155
cc_2089 ( N_noxref_3_c_2118_n N_noxref_5_c_2530_n ) capacitor c=3.10026e-19 \
 //x=6.425 //y=5.155 //x2=3.985 //y2=5.155
cc_2090 ( N_noxref_3_M59_noxref_g N_noxref_5_c_2530_n ) capacitor c=0.0194981f \
 //x=3.51 //y=6.02 //x2=3.985 //y2=5.155
cc_2091 ( N_noxref_3_c_2176_p N_noxref_5_c_2530_n ) capacitor c=0.00201851f \
 //x=3.33 //y=4.7 //x2=3.985 //y2=5.155
cc_2092 ( N_noxref_3_c_2177_p N_noxref_5_c_2496_n ) capacitor c=0.00359704f \
 //x=3.695 //y=1.415 //x2=3.985 //y2=1.665
cc_2093 ( N_noxref_3_c_2178_p N_noxref_5_c_2496_n ) capacitor c=0.00457401f \
 //x=3.85 //y=1.26 //x2=3.985 //y2=1.665
cc_2094 ( N_noxref_3_c_2093_n N_noxref_5_c_2583_n ) capacitor c=0.00628992f \
 //x=8.765 //y=3.33 //x2=3.67 //y2=1.665
cc_2095 ( N_noxref_3_c_2093_n N_noxref_5_c_2534_n ) capacitor c=0.0260398f \
 //x=8.765 //y=3.33 //x2=4.07 //y2=3.7
cc_2096 ( N_noxref_3_c_2097_n N_noxref_5_c_2534_n ) capacitor c=0.00179385f \
 //x=3.445 //y=3.33 //x2=4.07 //y2=3.7
cc_2097 ( N_noxref_3_c_2099_n N_noxref_5_c_2534_n ) capacitor c=0.0831612f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_2098 ( N_noxref_3_c_2183_p N_noxref_5_c_2534_n ) capacitor c=0.00877984f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_2099 ( N_noxref_3_c_2184_p N_noxref_5_c_2534_n ) capacitor c=0.00283672f \
 //x=3.33 //y=1.915 //x2=4.07 //y2=3.7
cc_2100 ( N_noxref_3_c_2176_p N_noxref_5_c_2534_n ) capacitor c=0.013693f \
 //x=3.33 //y=4.7 //x2=4.07 //y2=3.7
cc_2101 ( N_noxref_3_c_2093_n N_noxref_5_c_2497_n ) capacitor c=0.0268062f \
 //x=8.765 //y=3.33 //x2=5.92 //y2=2.08
cc_2102 ( N_noxref_3_c_2099_n N_noxref_5_c_2497_n ) capacitor c=9.66956e-19 \
 //x=3.33 //y=2.08 //x2=5.92 //y2=2.08
cc_2103 ( N_noxref_3_c_2099_n N_noxref_5_c_2592_n ) capacitor c=0.0171303f \
 //x=3.33 //y=2.08 //x2=3.29 //y2=5.155
cc_2104 ( N_noxref_3_c_2176_p N_noxref_5_c_2592_n ) capacitor c=0.00475601f \
 //x=3.33 //y=4.7 //x2=3.29 //y2=5.155
cc_2105 ( N_noxref_3_c_2118_n N_noxref_5_M60_noxref_g ) capacitor c=0.0213876f \
 //x=6.425 //y=5.155 //x2=6.12 //y2=6.02
cc_2106 ( N_noxref_3_c_2114_n N_noxref_5_M61_noxref_g ) capacitor c=0.0168349f \
 //x=7.135 //y=5.155 //x2=6.56 //y2=6.02
cc_2107 ( N_noxref_3_M60_noxref_d N_noxref_5_M61_noxref_g ) capacitor \
 c=0.0180032f //x=6.195 //y=5.02 //x2=6.56 //y2=6.02
cc_2108 ( N_noxref_3_c_2118_n N_noxref_5_c_2597_n ) capacitor c=0.00428486f \
 //x=6.425 //y=5.155 //x2=6.485 //y2=4.79
cc_2109 ( N_noxref_3_c_2194_p N_noxref_5_M2_noxref_d ) capacitor c=0.00217566f \
 //x=3.32 //y=0.915 //x2=3.395 //y2=0.915
cc_2110 ( N_noxref_3_c_2195_p N_noxref_5_M2_noxref_d ) capacitor c=0.0034598f \
 //x=3.32 //y=1.26 //x2=3.395 //y2=0.915
cc_2111 ( N_noxref_3_c_2196_p N_noxref_5_M2_noxref_d ) capacitor c=0.00544291f \
 //x=3.32 //y=1.57 //x2=3.395 //y2=0.915
cc_2112 ( N_noxref_3_c_2197_p N_noxref_5_M2_noxref_d ) capacitor c=0.00241102f \
 //x=3.695 //y=0.76 //x2=3.395 //y2=0.915
cc_2113 ( N_noxref_3_c_2177_p N_noxref_5_M2_noxref_d ) capacitor c=0.0140297f \
 //x=3.695 //y=1.415 //x2=3.395 //y2=0.915
cc_2114 ( N_noxref_3_c_2199_p N_noxref_5_M2_noxref_d ) capacitor c=0.00219619f \
 //x=3.85 //y=0.915 //x2=3.395 //y2=0.915
cc_2115 ( N_noxref_3_c_2178_p N_noxref_5_M2_noxref_d ) capacitor c=0.00603828f \
 //x=3.85 //y=1.26 //x2=3.395 //y2=0.915
cc_2116 ( N_noxref_3_c_2184_p N_noxref_5_M2_noxref_d ) capacitor c=0.00661782f \
 //x=3.33 //y=1.915 //x2=3.395 //y2=0.915
cc_2117 ( N_noxref_3_M58_noxref_g N_noxref_5_M58_noxref_d ) capacitor \
 c=0.0180032f //x=3.07 //y=6.02 //x2=3.145 //y2=5.02
cc_2118 ( N_noxref_3_M59_noxref_g N_noxref_5_M58_noxref_d ) capacitor \
 c=0.0194246f //x=3.51 //y=6.02 //x2=3.145 //y2=5.02
cc_2119 ( N_noxref_3_c_2093_n N_noxref_6_c_2748_n ) capacitor c=0.0558554f \
 //x=8.765 //y=3.33 //x2=11.355 //y2=4.07
cc_2120 ( N_noxref_3_c_2097_n N_noxref_6_c_2748_n ) capacitor c=0.0135672f \
 //x=3.445 //y=3.33 //x2=11.355 //y2=4.07
cc_2121 ( N_noxref_3_c_2098_n N_noxref_6_c_2748_n ) capacitor c=0.010979f \
 //x=10.615 //y=3.33 //x2=11.355 //y2=4.07
cc_2122 ( N_noxref_3_c_2169_p N_noxref_6_c_2748_n ) capacitor c=4.80262e-19 \
 //x=8.995 //y=3.33 //x2=11.355 //y2=4.07
cc_2123 ( N_noxref_3_c_2099_n N_noxref_6_c_2748_n ) capacitor c=0.0206302f \
 //x=3.33 //y=2.08 //x2=11.355 //y2=4.07
cc_2124 ( N_noxref_3_c_2128_n N_noxref_6_c_2748_n ) capacitor c=0.0181982f \
 //x=8.88 //y=3.33 //x2=11.355 //y2=4.07
cc_2125 ( N_noxref_3_c_2101_n N_noxref_6_c_2748_n ) capacitor c=0.0184765f \
 //x=10.73 //y=2.08 //x2=11.355 //y2=4.07
cc_2126 ( N_noxref_3_c_2101_n N_noxref_6_c_2891_n ) capacitor c=0.00179385f \
 //x=10.73 //y=2.08 //x2=11.585 //y2=4.07
cc_2127 ( N_noxref_3_c_2099_n N_noxref_6_c_2750_n ) capacitor c=0.00175117f \
 //x=3.33 //y=2.08 //x2=1.11 //y2=2.08
cc_2128 ( N_noxref_3_c_2101_n N_noxref_6_c_2893_n ) capacitor c=0.00400249f \
 //x=10.73 //y=2.08 //x2=11.47 //y2=4.535
cc_2129 ( N_noxref_3_c_2140_n N_noxref_6_c_2893_n ) capacitor c=0.00417994f \
 //x=10.73 //y=4.7 //x2=11.47 //y2=4.535
cc_2130 ( N_noxref_3_c_2098_n N_noxref_6_c_2751_n ) capacitor c=0.00318578f \
 //x=10.615 //y=3.33 //x2=11.47 //y2=2.08
cc_2131 ( N_noxref_3_c_2128_n N_noxref_6_c_2751_n ) capacitor c=9.69022e-19 \
 //x=8.88 //y=3.33 //x2=11.47 //y2=2.08
cc_2132 ( N_noxref_3_c_2101_n N_noxref_6_c_2751_n ) capacitor c=0.0746656f \
 //x=10.73 //y=2.08 //x2=11.47 //y2=2.08
cc_2133 ( N_noxref_3_c_2106_n N_noxref_6_c_2751_n ) capacitor c=0.00284029f \
 //x=10.535 //y=1.915 //x2=11.47 //y2=2.08
cc_2134 ( N_noxref_3_M66_noxref_g N_noxref_6_M68_noxref_g ) capacitor \
 c=0.0104611f //x=10.63 //y=6.02 //x2=11.51 //y2=6.02
cc_2135 ( N_noxref_3_M67_noxref_g N_noxref_6_M68_noxref_g ) capacitor \
 c=0.106811f //x=11.07 //y=6.02 //x2=11.51 //y2=6.02
cc_2136 ( N_noxref_3_M67_noxref_g N_noxref_6_M69_noxref_g ) capacitor \
 c=0.0100341f //x=11.07 //y=6.02 //x2=11.95 //y2=6.02
cc_2137 ( N_noxref_3_c_2102_n N_noxref_6_c_2902_n ) capacitor c=4.86506e-19 \
 //x=10.535 //y=0.865 //x2=11.505 //y2=0.905
cc_2138 ( N_noxref_3_c_2104_n N_noxref_6_c_2902_n ) capacitor c=0.00152104f \
 //x=10.535 //y=1.21 //x2=11.505 //y2=0.905
cc_2139 ( N_noxref_3_c_2109_n N_noxref_6_c_2902_n ) capacitor c=0.0151475f \
 //x=11.065 //y=0.865 //x2=11.505 //y2=0.905
cc_2140 ( N_noxref_3_c_2105_n N_noxref_6_c_2905_n ) capacitor c=0.00109982f \
 //x=10.535 //y=1.52 //x2=11.505 //y2=1.25
cc_2141 ( N_noxref_3_c_2111_n N_noxref_6_c_2905_n ) capacitor c=0.0111064f \
 //x=11.065 //y=1.21 //x2=11.505 //y2=1.25
cc_2142 ( N_noxref_3_c_2105_n N_noxref_6_c_2907_n ) capacitor c=9.57794e-19 \
 //x=10.535 //y=1.52 //x2=11.505 //y2=1.56
cc_2143 ( N_noxref_3_c_2106_n N_noxref_6_c_2907_n ) capacitor c=0.00662747f \
 //x=10.535 //y=1.915 //x2=11.505 //y2=1.56
cc_2144 ( N_noxref_3_c_2111_n N_noxref_6_c_2907_n ) capacitor c=0.00862358f \
 //x=11.065 //y=1.21 //x2=11.505 //y2=1.56
cc_2145 ( N_noxref_3_c_2109_n N_noxref_6_c_2910_n ) capacitor c=0.00124821f \
 //x=11.065 //y=0.865 //x2=12.035 //y2=0.905
cc_2146 ( N_noxref_3_c_2111_n N_noxref_6_c_2911_n ) capacitor c=0.00200715f \
 //x=11.065 //y=1.21 //x2=12.035 //y2=1.25
cc_2147 ( N_noxref_3_c_2101_n N_noxref_6_c_2912_n ) capacitor c=0.00282278f \
 //x=10.73 //y=2.08 //x2=11.47 //y2=2.08
cc_2148 ( N_noxref_3_c_2106_n N_noxref_6_c_2912_n ) capacitor c=0.0172771f \
 //x=10.535 //y=1.915 //x2=11.47 //y2=2.08
cc_2149 ( N_noxref_3_c_2101_n N_noxref_6_c_2914_n ) capacitor c=0.00344981f \
 //x=10.73 //y=2.08 //x2=11.5 //y2=4.7
cc_2150 ( N_noxref_3_c_2140_n N_noxref_6_c_2914_n ) capacitor c=0.0293367f \
 //x=10.73 //y=4.7 //x2=11.5 //y2=4.7
cc_2151 ( N_noxref_3_c_2093_n N_D_c_4434_n ) capacitor c=0.0674719f //x=8.765 \
 //y=3.33 //x2=32.815 //y2=2.59
cc_2152 ( N_noxref_3_c_2098_n N_D_c_4434_n ) capacitor c=0.0838995f //x=10.615 \
 //y=3.33 //x2=32.815 //y2=2.59
cc_2153 ( N_noxref_3_c_2169_p N_D_c_4434_n ) capacitor c=0.0120889f //x=8.995 \
 //y=3.33 //x2=32.815 //y2=2.59
cc_2154 ( N_noxref_3_c_2128_n N_D_c_4434_n ) capacitor c=0.0192483f //x=8.88 \
 //y=3.33 //x2=32.815 //y2=2.59
cc_2155 ( N_noxref_3_c_2101_n N_D_c_4434_n ) capacitor c=0.0204451f //x=10.73 \
 //y=2.08 //x2=32.815 //y2=2.59
cc_2156 ( N_noxref_3_c_2093_n N_D_c_4441_n ) capacitor c=0.0133087f //x=8.765 \
 //y=3.33 //x2=7.145 //y2=2.59
cc_2157 ( N_noxref_3_c_2093_n N_D_c_4448_n ) capacitor c=0.0217085f //x=8.765 \
 //y=3.33 //x2=7.03 //y2=2.08
cc_2158 ( N_noxref_3_c_2114_n N_D_c_4448_n ) capacitor c=0.0144268f //x=7.135 \
 //y=5.155 //x2=7.03 //y2=2.08
cc_2159 ( N_noxref_3_c_2128_n N_D_c_4448_n ) capacitor c=0.00244556f //x=8.88 \
 //y=3.33 //x2=7.03 //y2=2.08
cc_2160 ( N_noxref_3_c_2114_n N_D_M62_noxref_g ) capacitor c=0.0165266f \
 //x=7.135 //y=5.155 //x2=7 //y2=6.02
cc_2161 ( N_noxref_3_M62_noxref_d N_D_M62_noxref_g ) capacitor c=0.0180032f \
 //x=7.075 //y=5.02 //x2=7 //y2=6.02
cc_2162 ( N_noxref_3_c_2120_n N_D_M63_noxref_g ) capacitor c=0.01736f \
 //x=8.015 //y=5.155 //x2=7.44 //y2=6.02
cc_2163 ( N_noxref_3_M62_noxref_d N_D_M63_noxref_g ) capacitor c=0.0180032f \
 //x=7.075 //y=5.02 //x2=7.44 //y2=6.02
cc_2164 ( N_noxref_3_c_2249_p N_D_c_4482_n ) capacitor c=0.00426767f //x=7.22 \
 //y=5.155 //x2=7.365 //y2=4.79
cc_2165 ( N_noxref_3_c_2114_n N_D_c_4483_n ) capacitor c=0.00322054f //x=7.135 \
 //y=5.155 //x2=7.03 //y2=4.7
cc_2166 ( N_noxref_3_c_2093_n N_CLK_c_4808_n ) capacitor c=0.00360213f \
 //x=8.765 //y=3.33 //x2=15.055 //y2=4.44
cc_2167 ( N_noxref_3_c_2097_n N_CLK_c_4808_n ) capacitor c=4.49102e-19 \
 //x=3.445 //y=3.33 //x2=15.055 //y2=4.44
cc_2168 ( N_noxref_3_c_2099_n N_CLK_c_4808_n ) capacitor c=0.0200057f //x=3.33 \
 //y=2.08 //x2=15.055 //y2=4.44
cc_2169 ( N_noxref_3_c_2114_n N_CLK_c_4808_n ) capacitor c=0.032141f //x=7.135 \
 //y=5.155 //x2=15.055 //y2=4.44
cc_2170 ( N_noxref_3_c_2118_n N_CLK_c_4808_n ) capacitor c=0.0230136f \
 //x=6.425 //y=5.155 //x2=15.055 //y2=4.44
cc_2171 ( N_noxref_3_c_2124_n N_CLK_c_4808_n ) capacitor c=0.0183122f \
 //x=8.795 //y=5.155 //x2=15.055 //y2=4.44
cc_2172 ( N_noxref_3_c_2128_n N_CLK_c_4808_n ) capacitor c=0.0210274f //x=8.88 \
 //y=3.33 //x2=15.055 //y2=4.44
cc_2173 ( N_noxref_3_c_2101_n N_CLK_c_4808_n ) capacitor c=0.0198304f \
 //x=10.73 //y=2.08 //x2=15.055 //y2=4.44
cc_2174 ( N_noxref_3_c_2176_p N_CLK_c_4808_n ) capacitor c=0.0111881f //x=3.33 \
 //y=4.7 //x2=15.055 //y2=4.44
cc_2175 ( N_noxref_3_c_2140_n N_CLK_c_4808_n ) capacitor c=0.0107057f \
 //x=10.73 //y=4.7 //x2=15.055 //y2=4.44
cc_2176 ( N_noxref_3_c_2099_n N_CLK_c_4825_n ) capacitor c=0.00153281f \
 //x=3.33 //y=2.08 //x2=2.335 //y2=4.44
cc_2177 ( N_noxref_3_c_2097_n N_CLK_c_4802_n ) capacitor c=0.00526349f \
 //x=3.445 //y=3.33 //x2=2.22 //y2=2.08
cc_2178 ( N_noxref_3_c_2099_n N_CLK_c_4802_n ) capacitor c=0.0511464f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_2179 ( N_noxref_3_c_2183_p N_CLK_c_4802_n ) capacitor c=0.00228632f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=2.08
cc_2180 ( N_noxref_3_c_2176_p N_CLK_c_4802_n ) capacitor c=0.00218014f \
 //x=3.33 //y=4.7 //x2=2.22 //y2=2.08
cc_2181 ( N_noxref_3_M58_noxref_g N_CLK_M56_noxref_g ) capacitor c=0.0101598f \
 //x=3.07 //y=6.02 //x2=2.19 //y2=6.02
cc_2182 ( N_noxref_3_M58_noxref_g N_CLK_M57_noxref_g ) capacitor c=0.0602553f \
 //x=3.07 //y=6.02 //x2=2.63 //y2=6.02
cc_2183 ( N_noxref_3_M59_noxref_g N_CLK_M57_noxref_g ) capacitor c=0.0101598f \
 //x=3.51 //y=6.02 //x2=2.63 //y2=6.02
cc_2184 ( N_noxref_3_c_2194_p N_CLK_c_4952_n ) capacitor c=0.00456962f \
 //x=3.32 //y=0.915 //x2=2.31 //y2=0.91
cc_2185 ( N_noxref_3_c_2195_p N_CLK_c_4953_n ) capacitor c=0.00438372f \
 //x=3.32 //y=1.26 //x2=2.31 //y2=1.22
cc_2186 ( N_noxref_3_c_2196_p N_CLK_c_4954_n ) capacitor c=0.00438372f \
 //x=3.32 //y=1.57 //x2=2.31 //y2=1.45
cc_2187 ( N_noxref_3_c_2099_n N_CLK_c_4955_n ) capacitor c=0.0023343f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_2188 ( N_noxref_3_c_2183_p N_CLK_c_4955_n ) capacitor c=0.00933826f \
 //x=3.33 //y=2.08 //x2=2.31 //y2=1.915
cc_2189 ( N_noxref_3_c_2184_p N_CLK_c_4955_n ) capacitor c=0.00438372f \
 //x=3.33 //y=1.915 //x2=2.31 //y2=1.915
cc_2190 ( N_noxref_3_c_2176_p N_CLK_c_4958_n ) capacitor c=0.0611812f //x=3.33 \
 //y=4.7 //x2=2.555 //y2=4.79
cc_2191 ( N_noxref_3_c_2099_n N_CLK_c_4959_n ) capacitor c=0.00142741f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=4.7
cc_2192 ( N_noxref_3_c_2176_p N_CLK_c_4959_n ) capacitor c=0.00487508f \
 //x=3.33 //y=4.7 //x2=2.22 //y2=4.7
cc_2193 ( N_noxref_3_c_2093_n N_RN_c_5846_n ) capacitor c=0.00399667f \
 //x=8.765 //y=3.33 //x2=16.165 //y2=2.22
cc_2194 ( N_noxref_3_c_2098_n N_RN_c_5846_n ) capacitor c=0.00800271f \
 //x=10.615 //y=3.33 //x2=16.165 //y2=2.22
cc_2195 ( N_noxref_3_c_2169_p N_RN_c_5846_n ) capacitor c=3.9466e-19 //x=8.995 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_2196 ( N_noxref_3_c_2281_p N_RN_c_5846_n ) capacitor c=0.016327f //x=8.48 \
 //y=1.665 //x2=16.165 //y2=2.22
cc_2197 ( N_noxref_3_c_2128_n N_RN_c_5846_n ) capacitor c=0.0197307f //x=8.88 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_2198 ( N_noxref_3_c_2101_n N_RN_c_5846_n ) capacitor c=0.0185012f //x=10.73 \
 //y=2.08 //x2=16.165 //y2=2.22
cc_2199 ( N_noxref_3_c_2106_n N_RN_c_5846_n ) capacitor c=0.00894156f \
 //x=10.535 //y=1.915 //x2=16.165 //y2=2.22
cc_2200 ( N_noxref_3_c_2093_n N_RN_c_5854_n ) capacitor c=7.40016e-19 \
 //x=8.765 //y=3.33 //x2=8.255 //y2=2.22
cc_2201 ( N_noxref_3_c_2128_n N_RN_c_5854_n ) capacitor c=0.00184436f //x=8.88 \
 //y=3.33 //x2=8.255 //y2=2.22
cc_2202 ( N_noxref_3_c_2093_n N_RN_c_5913_n ) capacitor c=0.0203592f //x=8.765 \
 //y=3.33 //x2=8.14 //y2=2.08
cc_2203 ( N_noxref_3_c_2169_p N_RN_c_5913_n ) capacitor c=0.00131333f \
 //x=8.995 //y=3.33 //x2=8.14 //y2=2.08
cc_2204 ( N_noxref_3_c_2128_n N_RN_c_5913_n ) capacitor c=0.077845f //x=8.88 \
 //y=3.33 //x2=8.14 //y2=2.08
cc_2205 ( N_noxref_3_c_2101_n N_RN_c_5913_n ) capacitor c=7.44267e-19 \
 //x=10.73 //y=2.08 //x2=8.14 //y2=2.08
cc_2206 ( N_noxref_3_c_2291_p N_RN_c_5913_n ) capacitor c=0.0166016f //x=8.1 \
 //y=5.155 //x2=8.14 //y2=2.08
cc_2207 ( N_noxref_3_c_2120_n N_RN_M64_noxref_g ) capacitor c=0.01736f \
 //x=8.015 //y=5.155 //x2=7.88 //y2=6.02
cc_2208 ( N_noxref_3_M64_noxref_d N_RN_M64_noxref_g ) capacitor c=0.0180032f \
 //x=7.955 //y=5.02 //x2=7.88 //y2=6.02
cc_2209 ( N_noxref_3_c_2124_n N_RN_M65_noxref_g ) capacitor c=0.0194981f \
 //x=8.795 //y=5.155 //x2=8.32 //y2=6.02
cc_2210 ( N_noxref_3_M64_noxref_d N_RN_M65_noxref_g ) capacitor c=0.0194246f \
 //x=7.955 //y=5.02 //x2=8.32 //y2=6.02
cc_2211 ( N_noxref_3_M5_noxref_d N_RN_c_5988_n ) capacitor c=0.00217566f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=0.915
cc_2212 ( N_noxref_3_M5_noxref_d N_RN_c_5989_n ) capacitor c=0.0034598f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=1.26
cc_2213 ( N_noxref_3_M5_noxref_d N_RN_c_5990_n ) capacitor c=0.00546784f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=1.57
cc_2214 ( N_noxref_3_M5_noxref_d N_RN_c_5991_n ) capacitor c=0.00241102f \
 //x=8.205 //y=0.915 //x2=8.505 //y2=0.76
cc_2215 ( N_noxref_3_c_2100_n N_RN_c_5992_n ) capacitor c=0.00371277f \
 //x=8.795 //y=1.665 //x2=8.505 //y2=1.415
cc_2216 ( N_noxref_3_M5_noxref_d N_RN_c_5992_n ) capacitor c=0.0138621f \
 //x=8.205 //y=0.915 //x2=8.505 //y2=1.415
cc_2217 ( N_noxref_3_M5_noxref_d N_RN_c_5994_n ) capacitor c=0.00219619f \
 //x=8.205 //y=0.915 //x2=8.66 //y2=0.915
cc_2218 ( N_noxref_3_c_2100_n N_RN_c_5995_n ) capacitor c=0.00457401f \
 //x=8.795 //y=1.665 //x2=8.66 //y2=1.26
cc_2219 ( N_noxref_3_M5_noxref_d N_RN_c_5995_n ) capacitor c=0.00603828f \
 //x=8.205 //y=0.915 //x2=8.66 //y2=1.26
cc_2220 ( N_noxref_3_c_2128_n N_RN_c_5997_n ) capacitor c=0.00709342f //x=8.88 \
 //y=3.33 //x2=8.14 //y2=2.08
cc_2221 ( N_noxref_3_c_2128_n N_RN_c_5998_n ) capacitor c=0.00283672f //x=8.88 \
 //y=3.33 //x2=8.14 //y2=1.915
cc_2222 ( N_noxref_3_M5_noxref_d N_RN_c_5998_n ) capacitor c=0.00661782f \
 //x=8.205 //y=0.915 //x2=8.14 //y2=1.915
cc_2223 ( N_noxref_3_c_2124_n N_RN_c_6000_n ) capacitor c=0.00201851f \
 //x=8.795 //y=5.155 //x2=8.14 //y2=4.7
cc_2224 ( N_noxref_3_c_2128_n N_RN_c_6000_n ) capacitor c=0.013844f //x=8.88 \
 //y=3.33 //x2=8.14 //y2=4.7
cc_2225 ( N_noxref_3_c_2291_p N_RN_c_6000_n ) capacitor c=0.00475601f //x=8.1 \
 //y=5.155 //x2=8.14 //y2=4.7
cc_2226 ( N_noxref_3_c_2093_n N_noxref_24_c_9317_n ) capacitor c=2.45218e-19 \
 //x=8.765 //y=3.33 //x2=3.985 //y2=0.54
cc_2227 ( N_noxref_3_c_2099_n N_noxref_24_c_9317_n ) capacitor c=0.00208521f \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_2228 ( N_noxref_3_c_2194_p N_noxref_24_c_9317_n ) capacitor c=0.0194423f \
 //x=3.32 //y=0.915 //x2=3.985 //y2=0.54
cc_2229 ( N_noxref_3_c_2199_p N_noxref_24_c_9317_n ) capacitor c=0.00656458f \
 //x=3.85 //y=0.915 //x2=3.985 //y2=0.54
cc_2230 ( N_noxref_3_c_2183_p N_noxref_24_c_9317_n ) capacitor c=2.20712e-19 \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_2231 ( N_noxref_3_c_2195_p N_noxref_24_c_9330_n ) capacitor c=0.00538829f \
 //x=3.32 //y=1.26 //x2=3.1 //y2=0.995
cc_2232 ( N_noxref_3_c_2194_p N_noxref_24_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=0.915 //x2=2.965 //y2=0.375
cc_2233 ( N_noxref_3_c_2196_p N_noxref_24_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=1.57 //x2=2.965 //y2=0.375
cc_2234 ( N_noxref_3_c_2199_p N_noxref_24_M2_noxref_s ) capacitor c=0.0143002f \
 //x=3.85 //y=0.915 //x2=2.965 //y2=0.375
cc_2235 ( N_noxref_3_c_2178_p N_noxref_24_M2_noxref_s ) capacitor \
 c=0.00290153f //x=3.85 //y=1.26 //x2=2.965 //y2=0.375
cc_2236 ( N_noxref_3_c_2093_n N_noxref_25_c_9379_n ) capacitor c=0.00243521f \
 //x=8.765 //y=3.33 //x2=5.4 //y2=1.505
cc_2237 ( N_noxref_3_c_2093_n N_noxref_25_c_9364_n ) capacitor c=0.0103731f \
 //x=8.765 //y=3.33 //x2=6.285 //y2=1.59
cc_2238 ( N_noxref_3_c_2093_n N_noxref_25_c_9381_n ) capacitor c=0.00504206f \
 //x=8.765 //y=3.33 //x2=7.255 //y2=1.59
cc_2239 ( N_noxref_3_c_2093_n N_noxref_25_M3_noxref_s ) capacitor \
 c=0.00243521f //x=8.765 //y=3.33 //x2=5.265 //y2=0.375
cc_2240 ( N_noxref_3_M5_noxref_d N_noxref_25_M3_noxref_s ) capacitor \
 c=0.00309936f //x=8.205 //y=0.915 //x2=5.265 //y2=0.375
cc_2241 ( N_noxref_3_c_2100_n N_noxref_26_c_9421_n ) capacitor c=0.00457167f \
 //x=8.795 //y=1.665 //x2=8.795 //y2=0.54
cc_2242 ( N_noxref_3_M5_noxref_d N_noxref_26_c_9421_n ) capacitor c=0.0115903f \
 //x=8.205 //y=0.915 //x2=8.795 //y2=0.54
cc_2243 ( N_noxref_3_c_2281_p N_noxref_26_c_9431_n ) capacitor c=0.020048f \
 //x=8.48 //y=1.665 //x2=7.91 //y2=0.995
cc_2244 ( N_noxref_3_M5_noxref_d N_noxref_26_M4_noxref_d ) capacitor \
 c=5.27807e-19 //x=8.205 //y=0.915 //x2=6.67 //y2=0.91
cc_2245 ( N_noxref_3_c_2100_n N_noxref_26_M5_noxref_s ) capacitor c=0.0196084f \
 //x=8.795 //y=1.665 //x2=7.775 //y2=0.375
cc_2246 ( N_noxref_3_M5_noxref_d N_noxref_26_M5_noxref_s ) capacitor \
 c=0.0426444f //x=8.205 //y=0.915 //x2=7.775 //y2=0.375
cc_2247 ( N_noxref_3_c_2100_n N_noxref_27_c_9487_n ) capacitor c=3.04182e-19 \
 //x=8.795 //y=1.665 //x2=10.315 //y2=1.495
cc_2248 ( N_noxref_3_c_2106_n N_noxref_27_c_9487_n ) capacitor c=0.0034165f \
 //x=10.535 //y=1.915 //x2=10.315 //y2=1.495
cc_2249 ( N_noxref_3_c_2101_n N_noxref_27_c_9469_n ) capacitor c=0.011618f \
 //x=10.73 //y=2.08 //x2=11.2 //y2=1.58
cc_2250 ( N_noxref_3_c_2105_n N_noxref_27_c_9469_n ) capacitor c=0.00696403f \
 //x=10.535 //y=1.52 //x2=11.2 //y2=1.58
cc_2251 ( N_noxref_3_c_2106_n N_noxref_27_c_9469_n ) capacitor c=0.0174694f \
 //x=10.535 //y=1.915 //x2=11.2 //y2=1.58
cc_2252 ( N_noxref_3_c_2108_n N_noxref_27_c_9469_n ) capacitor c=0.00776811f \
 //x=10.91 //y=1.365 //x2=11.2 //y2=1.58
cc_2253 ( N_noxref_3_c_2111_n N_noxref_27_c_9469_n ) capacitor c=0.00339872f \
 //x=11.065 //y=1.21 //x2=11.2 //y2=1.58
cc_2254 ( N_noxref_3_c_2106_n N_noxref_27_c_9476_n ) capacitor c=6.71402e-19 \
 //x=10.535 //y=1.915 //x2=11.285 //y2=1.495
cc_2255 ( N_noxref_3_c_2102_n N_noxref_27_M6_noxref_s ) capacitor c=0.0327502f \
 //x=10.535 //y=0.865 //x2=10.18 //y2=0.365
cc_2256 ( N_noxref_3_c_2105_n N_noxref_27_M6_noxref_s ) capacitor \
 c=3.48408e-19 //x=10.535 //y=1.52 //x2=10.18 //y2=0.365
cc_2257 ( N_noxref_3_c_2109_n N_noxref_27_M6_noxref_s ) capacitor c=0.0120759f \
 //x=11.065 //y=0.865 //x2=10.18 //y2=0.365
cc_2258 ( N_noxref_4_c_2343_n N_noxref_5_c_2495_n ) capacitor c=0.176049f \
 //x=13.945 //y=3.33 //x2=18.755 //y2=3.7
cc_2259 ( N_noxref_4_c_2391_n N_noxref_5_c_2495_n ) capacitor c=0.0293967f \
 //x=12.325 //y=3.33 //x2=18.755 //y2=3.7
cc_2260 ( N_noxref_4_c_2345_n N_noxref_5_c_2495_n ) capacitor c=0.0206034f \
 //x=12.21 //y=3.33 //x2=18.755 //y2=3.7
cc_2261 ( N_noxref_4_c_2346_n N_noxref_5_c_2495_n ) capacitor c=0.0216236f \
 //x=14.06 //y=2.08 //x2=18.755 //y2=3.7
cc_2262 ( N_noxref_4_c_2343_n N_noxref_6_c_2787_n ) capacitor c=0.0107156f \
 //x=13.945 //y=3.33 //x2=16.905 //y2=4.07
cc_2263 ( N_noxref_4_c_2391_n N_noxref_6_c_2787_n ) capacitor c=8.88358e-19 \
 //x=12.325 //y=3.33 //x2=16.905 //y2=4.07
cc_2264 ( N_noxref_4_c_2345_n N_noxref_6_c_2787_n ) capacitor c=0.0181936f \
 //x=12.21 //y=3.33 //x2=16.905 //y2=4.07
cc_2265 ( N_noxref_4_c_2346_n N_noxref_6_c_2787_n ) capacitor c=0.019517f \
 //x=14.06 //y=2.08 //x2=16.905 //y2=4.07
cc_2266 ( N_noxref_4_c_2345_n N_noxref_6_c_2891_n ) capacitor c=0.00179385f \
 //x=12.21 //y=3.33 //x2=11.585 //y2=4.07
cc_2267 ( N_noxref_4_c_2360_n N_noxref_6_c_2893_n ) capacitor c=0.0126603f \
 //x=11.645 //y=5.2 //x2=11.47 //y2=4.535
cc_2268 ( N_noxref_4_c_2345_n N_noxref_6_c_2893_n ) capacitor c=0.0101115f \
 //x=12.21 //y=3.33 //x2=11.47 //y2=4.535
cc_2269 ( N_noxref_4_c_2391_n N_noxref_6_c_2751_n ) capacitor c=0.00329059f \
 //x=12.325 //y=3.33 //x2=11.47 //y2=2.08
cc_2270 ( N_noxref_4_c_2345_n N_noxref_6_c_2751_n ) capacitor c=0.0696877f \
 //x=12.21 //y=3.33 //x2=11.47 //y2=2.08
cc_2271 ( N_noxref_4_c_2346_n N_noxref_6_c_2751_n ) capacitor c=9.69022e-19 \
 //x=14.06 //y=2.08 //x2=11.47 //y2=2.08
cc_2272 ( N_noxref_4_M71_noxref_g N_noxref_6_c_2798_n ) capacitor c=0.0168349f \
 //x=14.7 //y=6.02 //x2=15.275 //y2=5.155
cc_2273 ( N_noxref_4_c_2345_n N_noxref_6_c_2802_n ) capacitor c=2.97874e-19 \
 //x=12.21 //y=3.33 //x2=14.565 //y2=5.155
cc_2274 ( N_noxref_4_M70_noxref_g N_noxref_6_c_2802_n ) capacitor c=0.0213876f \
 //x=14.26 //y=6.02 //x2=14.565 //y2=5.155
cc_2275 ( N_noxref_4_c_2416_p N_noxref_6_c_2802_n ) capacitor c=0.00428486f \
 //x=14.625 //y=4.79 //x2=14.565 //y2=5.155
cc_2276 ( N_noxref_4_c_2360_n N_noxref_6_M68_noxref_g ) capacitor c=0.0166421f \
 //x=11.645 //y=5.2 //x2=11.51 //y2=6.02
cc_2277 ( N_noxref_4_M68_noxref_d N_noxref_6_M68_noxref_g ) capacitor \
 c=0.0173476f //x=11.585 //y=5.02 //x2=11.51 //y2=6.02
cc_2278 ( N_noxref_4_c_2366_n N_noxref_6_M69_noxref_g ) capacitor c=0.018922f \
 //x=12.125 //y=5.2 //x2=11.95 //y2=6.02
cc_2279 ( N_noxref_4_M68_noxref_d N_noxref_6_M69_noxref_g ) capacitor \
 c=0.0179769f //x=11.585 //y=5.02 //x2=11.95 //y2=6.02
cc_2280 ( N_noxref_4_M7_noxref_d N_noxref_6_c_2902_n ) capacitor c=0.00217566f \
 //x=11.58 //y=0.905 //x2=11.505 //y2=0.905
cc_2281 ( N_noxref_4_M7_noxref_d N_noxref_6_c_2905_n ) capacitor c=0.0034598f \
 //x=11.58 //y=0.905 //x2=11.505 //y2=1.25
cc_2282 ( N_noxref_4_M7_noxref_d N_noxref_6_c_2907_n ) capacitor c=0.0066953f \
 //x=11.58 //y=0.905 //x2=11.505 //y2=1.56
cc_2283 ( N_noxref_4_c_2345_n N_noxref_6_c_2937_n ) capacitor c=0.0142673f \
 //x=12.21 //y=3.33 //x2=11.875 //y2=4.79
cc_2284 ( N_noxref_4_c_2425_p N_noxref_6_c_2937_n ) capacitor c=0.00407665f \
 //x=11.73 //y=5.2 //x2=11.875 //y2=4.79
cc_2285 ( N_noxref_4_M7_noxref_d N_noxref_6_c_2939_n ) capacitor c=0.00241102f \
 //x=11.58 //y=0.905 //x2=11.88 //y2=0.75
cc_2286 ( N_noxref_4_c_2344_n N_noxref_6_c_2940_n ) capacitor c=0.00371277f \
 //x=12.125 //y=1.655 //x2=11.88 //y2=1.405
cc_2287 ( N_noxref_4_M7_noxref_d N_noxref_6_c_2940_n ) capacitor c=0.0137169f \
 //x=11.58 //y=0.905 //x2=11.88 //y2=1.405
cc_2288 ( N_noxref_4_M7_noxref_d N_noxref_6_c_2910_n ) capacitor c=0.00132245f \
 //x=11.58 //y=0.905 //x2=12.035 //y2=0.905
cc_2289 ( N_noxref_4_c_2344_n N_noxref_6_c_2911_n ) capacitor c=0.00457401f \
 //x=12.125 //y=1.655 //x2=12.035 //y2=1.25
cc_2290 ( N_noxref_4_M7_noxref_d N_noxref_6_c_2911_n ) capacitor c=0.00566463f \
 //x=11.58 //y=0.905 //x2=12.035 //y2=1.25
cc_2291 ( N_noxref_4_c_2345_n N_noxref_6_c_2912_n ) capacitor c=0.00731987f \
 //x=12.21 //y=3.33 //x2=11.47 //y2=2.08
cc_2292 ( N_noxref_4_c_2345_n N_noxref_6_c_2946_n ) capacitor c=0.00306024f \
 //x=12.21 //y=3.33 //x2=11.47 //y2=1.915
cc_2293 ( N_noxref_4_M7_noxref_d N_noxref_6_c_2946_n ) capacitor c=0.00660593f \
 //x=11.58 //y=0.905 //x2=11.47 //y2=1.915
cc_2294 ( N_noxref_4_c_2360_n N_noxref_6_c_2914_n ) capacitor c=0.00346527f \
 //x=11.645 //y=5.2 //x2=11.5 //y2=4.7
cc_2295 ( N_noxref_4_c_2345_n N_noxref_6_c_2914_n ) capacitor c=0.00517969f \
 //x=12.21 //y=3.33 //x2=11.5 //y2=4.7
cc_2296 ( N_noxref_4_M71_noxref_g N_noxref_6_M70_noxref_d ) capacitor \
 c=0.0180032f //x=14.7 //y=6.02 //x2=14.335 //y2=5.02
cc_2297 ( N_noxref_4_c_2343_n N_D_c_4434_n ) capacitor c=0.0844336f //x=13.945 \
 //y=3.33 //x2=32.815 //y2=2.59
cc_2298 ( N_noxref_4_c_2391_n N_D_c_4434_n ) capacitor c=0.0133398f //x=12.325 \
 //y=3.33 //x2=32.815 //y2=2.59
cc_2299 ( N_noxref_4_c_2345_n N_D_c_4434_n ) capacitor c=0.019254f //x=12.21 \
 //y=3.33 //x2=32.815 //y2=2.59
cc_2300 ( N_noxref_4_c_2346_n N_D_c_4434_n ) capacitor c=0.0214832f //x=14.06 \
 //y=2.08 //x2=32.815 //y2=2.59
cc_2301 ( N_noxref_4_c_2360_n N_CLK_c_4808_n ) capacitor c=0.0185297f \
 //x=11.645 //y=5.2 //x2=15.055 //y2=4.44
cc_2302 ( N_noxref_4_c_2364_n N_CLK_c_4808_n ) capacitor c=0.018142f \
 //x=10.935 //y=5.2 //x2=15.055 //y2=4.44
cc_2303 ( N_noxref_4_c_2345_n N_CLK_c_4808_n ) capacitor c=0.0208321f \
 //x=12.21 //y=3.33 //x2=15.055 //y2=4.44
cc_2304 ( N_noxref_4_c_2346_n N_CLK_c_4808_n ) capacitor c=0.0208709f \
 //x=14.06 //y=2.08 //x2=15.055 //y2=4.44
cc_2305 ( N_noxref_4_c_2378_n N_CLK_c_4808_n ) capacitor c=0.0166984f \
 //x=14.335 //y=4.79 //x2=15.055 //y2=4.44
cc_2306 ( N_noxref_4_c_2346_n N_CLK_c_4843_n ) capacitor c=0.00153281f \
 //x=14.06 //y=2.08 //x2=15.285 //y2=4.44
cc_2307 ( N_noxref_4_c_2343_n N_CLK_c_4803_n ) capacitor c=0.00520283f \
 //x=13.945 //y=3.33 //x2=15.17 //y2=2.08
cc_2308 ( N_noxref_4_c_2345_n N_CLK_c_4803_n ) capacitor c=5.77178e-19 \
 //x=12.21 //y=3.33 //x2=15.17 //y2=2.08
cc_2309 ( N_noxref_4_c_2346_n N_CLK_c_4803_n ) capacitor c=0.0446069f \
 //x=14.06 //y=2.08 //x2=15.17 //y2=2.08
cc_2310 ( N_noxref_4_c_2351_n N_CLK_c_4803_n ) capacitor c=0.00210802f \
 //x=13.76 //y=1.915 //x2=15.17 //y2=2.08
cc_2311 ( N_noxref_4_c_2416_p N_CLK_c_4803_n ) capacitor c=0.00147352f \
 //x=14.625 //y=4.79 //x2=15.17 //y2=2.08
cc_2312 ( N_noxref_4_c_2378_n N_CLK_c_4803_n ) capacitor c=0.00141297f \
 //x=14.335 //y=4.79 //x2=15.17 //y2=2.08
cc_2313 ( N_noxref_4_M70_noxref_g N_CLK_M72_noxref_g ) capacitor c=0.0105869f \
 //x=14.26 //y=6.02 //x2=15.14 //y2=6.02
cc_2314 ( N_noxref_4_M71_noxref_g N_CLK_M72_noxref_g ) capacitor c=0.10632f \
 //x=14.7 //y=6.02 //x2=15.14 //y2=6.02
cc_2315 ( N_noxref_4_M71_noxref_g N_CLK_M73_noxref_g ) capacitor c=0.0101598f \
 //x=14.7 //y=6.02 //x2=15.58 //y2=6.02
cc_2316 ( N_noxref_4_c_2347_n N_CLK_c_4976_n ) capacitor c=5.72482e-19 \
 //x=13.76 //y=0.875 //x2=14.735 //y2=0.91
cc_2317 ( N_noxref_4_c_2349_n N_CLK_c_4976_n ) capacitor c=0.00149976f \
 //x=13.76 //y=1.22 //x2=14.735 //y2=0.91
cc_2318 ( N_noxref_4_c_2354_n N_CLK_c_4976_n ) capacitor c=0.0160123f \
 //x=14.29 //y=0.875 //x2=14.735 //y2=0.91
cc_2319 ( N_noxref_4_c_2350_n N_CLK_c_4979_n ) capacitor c=0.00111227f \
 //x=13.76 //y=1.53 //x2=14.735 //y2=1.22
cc_2320 ( N_noxref_4_c_2356_n N_CLK_c_4979_n ) capacitor c=0.0124075f \
 //x=14.29 //y=1.22 //x2=14.735 //y2=1.22
cc_2321 ( N_noxref_4_c_2354_n N_CLK_c_4981_n ) capacitor c=0.00103227f \
 //x=14.29 //y=0.875 //x2=15.26 //y2=0.91
cc_2322 ( N_noxref_4_c_2356_n N_CLK_c_4982_n ) capacitor c=0.0010154f \
 //x=14.29 //y=1.22 //x2=15.26 //y2=1.22
cc_2323 ( N_noxref_4_c_2356_n N_CLK_c_4983_n ) capacitor c=9.23422e-19 \
 //x=14.29 //y=1.22 //x2=15.26 //y2=1.45
cc_2324 ( N_noxref_4_c_2346_n N_CLK_c_4984_n ) capacitor c=0.00203769f \
 //x=14.06 //y=2.08 //x2=15.26 //y2=1.915
cc_2325 ( N_noxref_4_c_2351_n N_CLK_c_4984_n ) capacitor c=0.00834532f \
 //x=13.76 //y=1.915 //x2=15.26 //y2=1.915
cc_2326 ( N_noxref_4_c_2346_n N_CLK_c_4986_n ) capacitor c=0.00183762f \
 //x=14.06 //y=2.08 //x2=15.17 //y2=4.7
cc_2327 ( N_noxref_4_c_2416_p N_CLK_c_4986_n ) capacitor c=0.0168581f \
 //x=14.625 //y=4.79 //x2=15.17 //y2=4.7
cc_2328 ( N_noxref_4_c_2378_n N_CLK_c_4986_n ) capacitor c=0.00484466f \
 //x=14.335 //y=4.79 //x2=15.17 //y2=4.7
cc_2329 ( N_noxref_4_c_2343_n N_RN_c_5846_n ) capacitor c=0.00736619f \
 //x=13.945 //y=3.33 //x2=16.165 //y2=2.22
cc_2330 ( N_noxref_4_c_2391_n N_RN_c_5846_n ) capacitor c=6.29463e-19 \
 //x=12.325 //y=3.33 //x2=16.165 //y2=2.22
cc_2331 ( N_noxref_4_c_2472_p N_RN_c_5846_n ) capacitor c=0.0146822f \
 //x=11.855 //y=1.655 //x2=16.165 //y2=2.22
cc_2332 ( N_noxref_4_c_2345_n N_RN_c_5846_n ) capacitor c=0.0199049f //x=12.21 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_2333 ( N_noxref_4_c_2346_n N_RN_c_5846_n ) capacitor c=0.0192695f //x=14.06 \
 //y=2.08 //x2=16.165 //y2=2.22
cc_2334 ( N_noxref_4_c_2351_n N_RN_c_5846_n ) capacitor c=0.011987f //x=13.76 \
 //y=1.915 //x2=16.165 //y2=2.22
cc_2335 ( N_noxref_4_c_2346_n N_RN_c_5914_n ) capacitor c=0.00117207f \
 //x=14.06 //y=2.08 //x2=16.28 //y2=2.08
cc_2336 ( N_noxref_4_c_2472_p N_noxref_27_c_9487_n ) capacitor c=3.15806e-19 \
 //x=11.855 //y=1.655 //x2=10.315 //y2=1.495
cc_2337 ( N_noxref_4_c_2472_p N_noxref_27_c_9476_n ) capacitor c=0.020324f \
 //x=11.855 //y=1.655 //x2=11.285 //y2=1.495
cc_2338 ( N_noxref_4_c_2344_n N_noxref_27_c_9477_n ) capacitor c=0.00457164f \
 //x=12.125 //y=1.655 //x2=12.17 //y2=0.53
cc_2339 ( N_noxref_4_M7_noxref_d N_noxref_27_c_9477_n ) capacitor c=0.0115831f \
 //x=11.58 //y=0.905 //x2=12.17 //y2=0.53
cc_2340 ( N_noxref_4_c_2344_n N_noxref_27_M6_noxref_s ) capacitor c=0.013435f \
 //x=12.125 //y=1.655 //x2=10.18 //y2=0.365
cc_2341 ( N_noxref_4_M7_noxref_d N_noxref_27_M6_noxref_s ) capacitor \
 c=0.0439476f //x=11.58 //y=0.905 //x2=10.18 //y2=0.365
cc_2342 ( N_noxref_4_c_2344_n N_noxref_28_c_9535_n ) capacitor c=4.08644e-19 \
 //x=12.125 //y=1.655 //x2=13.54 //y2=1.505
cc_2343 ( N_noxref_4_c_2351_n N_noxref_28_c_9535_n ) capacitor c=0.0034165f \
 //x=13.76 //y=1.915 //x2=13.54 //y2=1.505
cc_2344 ( N_noxref_4_c_2346_n N_noxref_28_c_9520_n ) capacitor c=0.0115578f \
 //x=14.06 //y=2.08 //x2=14.425 //y2=1.59
cc_2345 ( N_noxref_4_c_2350_n N_noxref_28_c_9520_n ) capacitor c=0.00697148f \
 //x=13.76 //y=1.53 //x2=14.425 //y2=1.59
cc_2346 ( N_noxref_4_c_2351_n N_noxref_28_c_9520_n ) capacitor c=0.0204849f \
 //x=13.76 //y=1.915 //x2=14.425 //y2=1.59
cc_2347 ( N_noxref_4_c_2353_n N_noxref_28_c_9520_n ) capacitor c=0.00610316f \
 //x=14.135 //y=1.375 //x2=14.425 //y2=1.59
cc_2348 ( N_noxref_4_c_2356_n N_noxref_28_c_9520_n ) capacitor c=0.00698822f \
 //x=14.29 //y=1.22 //x2=14.425 //y2=1.59
cc_2349 ( N_noxref_4_c_2347_n N_noxref_28_M8_noxref_s ) capacitor c=0.0327271f \
 //x=13.76 //y=0.875 //x2=13.405 //y2=0.375
cc_2350 ( N_noxref_4_c_2350_n N_noxref_28_M8_noxref_s ) capacitor \
 c=7.99997e-19 //x=13.76 //y=1.53 //x2=13.405 //y2=0.375
cc_2351 ( N_noxref_4_c_2351_n N_noxref_28_M8_noxref_s ) capacitor \
 c=0.00122123f //x=13.76 //y=1.915 //x2=13.405 //y2=0.375
cc_2352 ( N_noxref_4_c_2354_n N_noxref_28_M8_noxref_s ) capacitor c=0.0121427f \
 //x=14.29 //y=0.875 //x2=13.405 //y2=0.375
cc_2353 ( N_noxref_4_M7_noxref_d N_noxref_28_M8_noxref_s ) capacitor \
 c=2.53688e-19 //x=11.58 //y=0.905 //x2=13.405 //y2=0.375
cc_2354 ( N_noxref_5_c_2568_n N_noxref_6_c_2748_n ) capacitor c=0.147447f \
 //x=5.805 //y=3.7 //x2=11.355 //y2=4.07
cc_2355 ( N_noxref_5_c_2569_n N_noxref_6_c_2748_n ) capacitor c=0.0294294f \
 //x=4.185 //y=3.7 //x2=11.355 //y2=4.07
cc_2356 ( N_noxref_5_c_2495_n N_noxref_6_c_2748_n ) capacitor c=0.467539f \
 //x=18.755 //y=3.7 //x2=11.355 //y2=4.07
cc_2357 ( N_noxref_5_c_2576_n N_noxref_6_c_2748_n ) capacitor c=0.0264476f \
 //x=6.035 //y=3.7 //x2=11.355 //y2=4.07
cc_2358 ( N_noxref_5_c_2524_n N_noxref_6_c_2748_n ) capacitor c=0.0154449f \
 //x=1.615 //y=5.155 //x2=11.355 //y2=4.07
cc_2359 ( N_noxref_5_c_2534_n N_noxref_6_c_2748_n ) capacitor c=0.0200328f \
 //x=4.07 //y=3.7 //x2=11.355 //y2=4.07
cc_2360 ( N_noxref_5_c_2497_n N_noxref_6_c_2748_n ) capacitor c=0.0213516f \
 //x=5.92 //y=2.08 //x2=11.355 //y2=4.07
cc_2361 ( N_noxref_5_c_2495_n N_noxref_6_c_2787_n ) capacitor c=0.468066f \
 //x=18.755 //y=3.7 //x2=16.905 //y2=4.07
cc_2362 ( N_noxref_5_c_2495_n N_noxref_6_c_2891_n ) capacitor c=0.0267832f \
 //x=18.755 //y=3.7 //x2=11.585 //y2=4.07
cc_2363 ( N_noxref_5_c_2495_n N_noxref_6_c_2788_n ) capacitor c=0.176507f \
 //x=18.755 //y=3.7 //x2=21.715 //y2=4.07
cc_2364 ( N_noxref_5_c_2498_n N_noxref_6_c_2788_n ) capacitor c=0.0213324f \
 //x=18.87 //y=2.08 //x2=21.715 //y2=4.07
cc_2365 ( N_noxref_5_c_2495_n N_noxref_6_c_2789_n ) capacitor c=0.0268461f \
 //x=18.755 //y=3.7 //x2=17.135 //y2=4.07
cc_2366 ( N_noxref_5_c_2498_n N_noxref_6_c_2789_n ) capacitor c=2.98083e-19 \
 //x=18.87 //y=2.08 //x2=17.135 //y2=4.07
cc_2367 ( N_noxref_5_c_2495_n N_noxref_6_c_2751_n ) capacitor c=0.0226566f \
 //x=18.755 //y=3.7 //x2=11.47 //y2=2.08
cc_2368 ( N_noxref_5_c_2495_n N_noxref_6_c_2812_n ) capacitor c=0.0251381f \
 //x=18.755 //y=3.7 //x2=17.02 //y2=4.07
cc_2369 ( N_noxref_5_c_2498_n N_noxref_6_c_2812_n ) capacitor c=0.0141021f \
 //x=18.87 //y=2.08 //x2=17.02 //y2=4.07
cc_2370 ( N_noxref_5_M77_noxref_g N_noxref_6_c_2813_n ) capacitor c=0.0168349f \
 //x=19.51 //y=6.02 //x2=20.085 //y2=5.155
cc_2371 ( N_noxref_5_M76_noxref_g N_noxref_6_c_2817_n ) capacitor c=0.0213876f \
 //x=19.07 //y=6.02 //x2=19.375 //y2=5.155
cc_2372 ( N_noxref_5_c_2630_p N_noxref_6_c_2817_n ) capacitor c=0.00428486f \
 //x=19.435 //y=4.79 //x2=19.375 //y2=5.155
cc_2373 ( N_noxref_5_c_2524_n N_noxref_6_M54_noxref_g ) capacitor c=0.0213876f \
 //x=1.615 //y=5.155 //x2=1.31 //y2=6.02
cc_2374 ( N_noxref_5_c_2520_n N_noxref_6_M55_noxref_g ) capacitor c=0.0178794f \
 //x=2.325 //y=5.155 //x2=1.75 //y2=6.02
cc_2375 ( N_noxref_5_M54_noxref_d N_noxref_6_M55_noxref_g ) capacitor \
 c=0.0180032f //x=1.385 //y=5.02 //x2=1.75 //y2=6.02
cc_2376 ( N_noxref_5_c_2524_n N_noxref_6_c_2973_n ) capacitor c=0.00429591f \
 //x=1.615 //y=5.155 //x2=1.675 //y2=4.79
cc_2377 ( N_noxref_5_M77_noxref_g N_noxref_6_M76_noxref_d ) capacitor \
 c=0.0180032f //x=19.51 //y=6.02 //x2=19.145 //y2=5.02
cc_2378 ( N_noxref_5_c_2495_n N_D_c_4434_n ) capacitor c=0.194153f //x=18.755 \
 //y=3.7 //x2=32.815 //y2=2.59
cc_2379 ( N_noxref_5_c_2498_n N_D_c_4434_n ) capacitor c=0.0227777f //x=18.87 \
 //y=2.08 //x2=32.815 //y2=2.59
cc_2380 ( N_noxref_5_c_2495_n N_D_c_4441_n ) capacitor c=7.19251e-19 \
 //x=18.755 //y=3.7 //x2=7.145 //y2=2.59
cc_2381 ( N_noxref_5_c_2497_n N_D_c_4441_n ) capacitor c=0.00526349f //x=5.92 \
 //y=2.08 //x2=7.145 //y2=2.59
cc_2382 ( N_noxref_5_c_2495_n N_D_c_4448_n ) capacitor c=0.0190398f //x=18.755 \
 //y=3.7 //x2=7.03 //y2=2.08
cc_2383 ( N_noxref_5_c_2576_n N_D_c_4448_n ) capacitor c=9.95819e-19 //x=6.035 \
 //y=3.7 //x2=7.03 //y2=2.08
cc_2384 ( N_noxref_5_c_2534_n N_D_c_4448_n ) capacitor c=4.0219e-19 //x=4.07 \
 //y=3.7 //x2=7.03 //y2=2.08
cc_2385 ( N_noxref_5_c_2497_n N_D_c_4448_n ) capacitor c=0.0464235f //x=5.92 \
 //y=2.08 //x2=7.03 //y2=2.08
cc_2386 ( N_noxref_5_c_2503_n N_D_c_4448_n ) capacitor c=0.00238338f //x=5.62 \
 //y=1.915 //x2=7.03 //y2=2.08
cc_2387 ( N_noxref_5_c_2597_n N_D_c_4448_n ) capacitor c=0.00147352f //x=6.485 \
 //y=4.79 //x2=7.03 //y2=2.08
cc_2388 ( N_noxref_5_c_2549_n N_D_c_4448_n ) capacitor c=0.00142741f //x=6.195 \
 //y=4.79 //x2=7.03 //y2=2.08
cc_2389 ( N_noxref_5_M60_noxref_g N_D_M62_noxref_g ) capacitor c=0.0105869f \
 //x=6.12 //y=6.02 //x2=7 //y2=6.02
cc_2390 ( N_noxref_5_M61_noxref_g N_D_M62_noxref_g ) capacitor c=0.10632f \
 //x=6.56 //y=6.02 //x2=7 //y2=6.02
cc_2391 ( N_noxref_5_M61_noxref_g N_D_M63_noxref_g ) capacitor c=0.0101598f \
 //x=6.56 //y=6.02 //x2=7.44 //y2=6.02
cc_2392 ( N_noxref_5_c_2499_n N_D_c_4502_n ) capacitor c=5.72482e-19 //x=5.62 \
 //y=0.875 //x2=6.595 //y2=0.91
cc_2393 ( N_noxref_5_c_2501_n N_D_c_4502_n ) capacitor c=0.00149976f //x=5.62 \
 //y=1.22 //x2=6.595 //y2=0.91
cc_2394 ( N_noxref_5_c_2506_n N_D_c_4502_n ) capacitor c=0.0160123f //x=6.15 \
 //y=0.875 //x2=6.595 //y2=0.91
cc_2395 ( N_noxref_5_c_2502_n N_D_c_4505_n ) capacitor c=0.00111227f //x=5.62 \
 //y=1.53 //x2=6.595 //y2=1.22
cc_2396 ( N_noxref_5_c_2508_n N_D_c_4505_n ) capacitor c=0.0124075f //x=6.15 \
 //y=1.22 //x2=6.595 //y2=1.22
cc_2397 ( N_noxref_5_c_2506_n N_D_c_4507_n ) capacitor c=0.00103227f //x=6.15 \
 //y=0.875 //x2=7.12 //y2=0.91
cc_2398 ( N_noxref_5_c_2508_n N_D_c_4508_n ) capacitor c=0.0010154f //x=6.15 \
 //y=1.22 //x2=7.12 //y2=1.22
cc_2399 ( N_noxref_5_c_2508_n N_D_c_4509_n ) capacitor c=9.23422e-19 //x=6.15 \
 //y=1.22 //x2=7.12 //y2=1.45
cc_2400 ( N_noxref_5_c_2497_n N_D_c_4510_n ) capacitor c=0.00231304f //x=5.92 \
 //y=2.08 //x2=7.12 //y2=1.915
cc_2401 ( N_noxref_5_c_2503_n N_D_c_4510_n ) capacitor c=0.00964411f //x=5.62 \
 //y=1.915 //x2=7.12 //y2=1.915
cc_2402 ( N_noxref_5_c_2497_n N_D_c_4483_n ) capacitor c=0.00183762f //x=5.92 \
 //y=2.08 //x2=7.03 //y2=4.7
cc_2403 ( N_noxref_5_c_2597_n N_D_c_4483_n ) capacitor c=0.0168581f //x=6.485 \
 //y=4.79 //x2=7.03 //y2=4.7
cc_2404 ( N_noxref_5_c_2549_n N_D_c_4483_n ) capacitor c=0.00484466f //x=6.195 \
 //y=4.79 //x2=7.03 //y2=4.7
cc_2405 ( N_noxref_5_c_2568_n N_CLK_c_4808_n ) capacitor c=0.00910993f \
 //x=5.805 //y=3.7 //x2=15.055 //y2=4.44
cc_2406 ( N_noxref_5_c_2569_n N_CLK_c_4808_n ) capacitor c=7.95009e-19 \
 //x=4.185 //y=3.7 //x2=15.055 //y2=4.44
cc_2407 ( N_noxref_5_c_2495_n N_CLK_c_4808_n ) capacitor c=0.0658043f \
 //x=18.755 //y=3.7 //x2=15.055 //y2=4.44
cc_2408 ( N_noxref_5_c_2576_n N_CLK_c_4808_n ) capacitor c=6.59178e-19 \
 //x=6.035 //y=3.7 //x2=15.055 //y2=4.44
cc_2409 ( N_noxref_5_c_2530_n N_CLK_c_4808_n ) capacitor c=0.0183122f \
 //x=3.985 //y=5.155 //x2=15.055 //y2=4.44
cc_2410 ( N_noxref_5_c_2534_n N_CLK_c_4808_n ) capacitor c=0.0210274f //x=4.07 \
 //y=3.7 //x2=15.055 //y2=4.44
cc_2411 ( N_noxref_5_c_2497_n N_CLK_c_4808_n ) capacitor c=0.0208709f //x=5.92 \
 //y=2.08 //x2=15.055 //y2=4.44
cc_2412 ( N_noxref_5_c_2670_p N_CLK_c_4808_n ) capacitor c=0.0311227f //x=2.41 \
 //y=5.155 //x2=15.055 //y2=4.44
cc_2413 ( N_noxref_5_c_2549_n N_CLK_c_4808_n ) capacitor c=0.0166984f \
 //x=6.195 //y=4.79 //x2=15.055 //y2=4.44
cc_2414 ( N_noxref_5_c_2520_n N_CLK_c_4825_n ) capacitor c=0.00330099f \
 //x=2.325 //y=5.155 //x2=2.335 //y2=4.44
cc_2415 ( N_noxref_5_c_2495_n N_CLK_c_4826_n ) capacitor c=0.0254092f \
 //x=18.755 //y=3.7 //x2=28.005 //y2=4.44
cc_2416 ( N_noxref_5_c_2498_n N_CLK_c_4826_n ) capacitor c=0.0208709f \
 //x=18.87 //y=2.08 //x2=28.005 //y2=4.44
cc_2417 ( N_noxref_5_c_2551_n N_CLK_c_4826_n ) capacitor c=0.0166984f \
 //x=19.145 //y=4.79 //x2=28.005 //y2=4.44
cc_2418 ( N_noxref_5_c_2495_n N_CLK_c_4843_n ) capacitor c=6.6036e-19 \
 //x=18.755 //y=3.7 //x2=15.285 //y2=4.44
cc_2419 ( N_noxref_5_c_2520_n N_CLK_c_4802_n ) capacitor c=0.014564f //x=2.325 \
 //y=5.155 //x2=2.22 //y2=2.08
cc_2420 ( N_noxref_5_c_2534_n N_CLK_c_4802_n ) capacitor c=0.00319363f \
 //x=4.07 //y=3.7 //x2=2.22 //y2=2.08
cc_2421 ( N_noxref_5_c_2495_n N_CLK_c_4803_n ) capacitor c=0.0228956f \
 //x=18.755 //y=3.7 //x2=15.17 //y2=2.08
cc_2422 ( N_noxref_5_c_2520_n N_CLK_M56_noxref_g ) capacitor c=0.016514f \
 //x=2.325 //y=5.155 //x2=2.19 //y2=6.02
cc_2423 ( N_noxref_5_M56_noxref_d N_CLK_M56_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.19 //y2=6.02
cc_2424 ( N_noxref_5_c_2526_n N_CLK_M57_noxref_g ) capacitor c=0.01736f \
 //x=3.205 //y=5.155 //x2=2.63 //y2=6.02
cc_2425 ( N_noxref_5_M56_noxref_d N_CLK_M57_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.63 //y2=6.02
cc_2426 ( N_noxref_5_c_2670_p N_CLK_c_4958_n ) capacitor c=0.00426767f \
 //x=2.41 //y=5.155 //x2=2.555 //y2=4.79
cc_2427 ( N_noxref_5_c_2520_n N_CLK_c_4959_n ) capacitor c=0.00322046f \
 //x=2.325 //y=5.155 //x2=2.22 //y2=4.7
cc_2428 ( N_noxref_5_c_2495_n N_RN_c_5846_n ) capacitor c=0.0190175f \
 //x=18.755 //y=3.7 //x2=16.165 //y2=2.22
cc_2429 ( N_noxref_5_c_2495_n N_RN_c_5856_n ) capacitor c=0.00896425f \
 //x=18.755 //y=3.7 //x2=19.865 //y2=2.22
cc_2430 ( N_noxref_5_c_2498_n N_RN_c_5856_n ) capacitor c=0.0192695f //x=18.87 \
 //y=2.08 //x2=19.865 //y2=2.22
cc_2431 ( N_noxref_5_c_2513_n N_RN_c_5856_n ) capacitor c=0.011987f //x=18.57 \
 //y=1.915 //x2=19.865 //y2=2.22
cc_2432 ( N_noxref_5_c_2495_n N_RN_c_5860_n ) capacitor c=4.25768e-19 \
 //x=18.755 //y=3.7 //x2=16.395 //y2=2.22
cc_2433 ( N_noxref_5_c_2498_n N_RN_c_5872_n ) capacitor c=0.00100368f \
 //x=18.87 //y=2.08 //x2=20.095 //y2=2.22
cc_2434 ( N_noxref_5_c_2513_n N_RN_c_5872_n ) capacitor c=2.11894e-19 \
 //x=18.57 //y=1.915 //x2=20.095 //y2=2.22
cc_2435 ( N_noxref_5_c_2495_n N_RN_c_5913_n ) capacitor c=0.0179999f \
 //x=18.755 //y=3.7 //x2=8.14 //y2=2.08
cc_2436 ( N_noxref_5_c_2497_n N_RN_c_5913_n ) capacitor c=0.00125649f //x=5.92 \
 //y=2.08 //x2=8.14 //y2=2.08
cc_2437 ( N_noxref_5_c_2495_n N_RN_c_5914_n ) capacitor c=0.0218601f \
 //x=18.755 //y=3.7 //x2=16.28 //y2=2.08
cc_2438 ( N_noxref_5_c_2498_n N_RN_c_5914_n ) capacitor c=8.87185e-19 \
 //x=18.87 //y=2.08 //x2=16.28 //y2=2.08
cc_2439 ( N_noxref_5_c_2495_n N_RN_c_5915_n ) capacitor c=0.00526349f \
 //x=18.755 //y=3.7 //x2=19.98 //y2=2.08
cc_2440 ( N_noxref_5_c_2498_n N_RN_c_5915_n ) capacitor c=0.0467233f //x=18.87 \
 //y=2.08 //x2=19.98 //y2=2.08
cc_2441 ( N_noxref_5_c_2513_n N_RN_c_5915_n ) capacitor c=0.00208635f \
 //x=18.57 //y=1.915 //x2=19.98 //y2=2.08
cc_2442 ( N_noxref_5_c_2630_p N_RN_c_5915_n ) capacitor c=0.00147352f \
 //x=19.435 //y=4.79 //x2=19.98 //y2=2.08
cc_2443 ( N_noxref_5_c_2551_n N_RN_c_5915_n ) capacitor c=0.00142741f \
 //x=19.145 //y=4.79 //x2=19.98 //y2=2.08
cc_2444 ( N_noxref_5_M76_noxref_g N_RN_M78_noxref_g ) capacitor c=0.0105869f \
 //x=19.07 //y=6.02 //x2=19.95 //y2=6.02
cc_2445 ( N_noxref_5_M77_noxref_g N_RN_M78_noxref_g ) capacitor c=0.10632f \
 //x=19.51 //y=6.02 //x2=19.95 //y2=6.02
cc_2446 ( N_noxref_5_M77_noxref_g N_RN_M79_noxref_g ) capacitor c=0.0101598f \
 //x=19.51 //y=6.02 //x2=20.39 //y2=6.02
cc_2447 ( N_noxref_5_c_2509_n N_RN_c_6029_n ) capacitor c=5.72482e-19 \
 //x=18.57 //y=0.875 //x2=19.545 //y2=0.91
cc_2448 ( N_noxref_5_c_2511_n N_RN_c_6029_n ) capacitor c=0.00149976f \
 //x=18.57 //y=1.22 //x2=19.545 //y2=0.91
cc_2449 ( N_noxref_5_c_2516_n N_RN_c_6029_n ) capacitor c=0.0160123f //x=19.1 \
 //y=0.875 //x2=19.545 //y2=0.91
cc_2450 ( N_noxref_5_c_2512_n N_RN_c_6032_n ) capacitor c=0.00111227f \
 //x=18.57 //y=1.53 //x2=19.545 //y2=1.22
cc_2451 ( N_noxref_5_c_2518_n N_RN_c_6032_n ) capacitor c=0.0124075f //x=19.1 \
 //y=1.22 //x2=19.545 //y2=1.22
cc_2452 ( N_noxref_5_c_2516_n N_RN_c_6034_n ) capacitor c=0.00103227f //x=19.1 \
 //y=0.875 //x2=20.07 //y2=0.91
cc_2453 ( N_noxref_5_c_2518_n N_RN_c_6035_n ) capacitor c=0.0010154f //x=19.1 \
 //y=1.22 //x2=20.07 //y2=1.22
cc_2454 ( N_noxref_5_c_2518_n N_RN_c_6036_n ) capacitor c=9.23422e-19 //x=19.1 \
 //y=1.22 //x2=20.07 //y2=1.45
cc_2455 ( N_noxref_5_c_2498_n N_RN_c_6037_n ) capacitor c=0.00203769f \
 //x=18.87 //y=2.08 //x2=20.07 //y2=1.915
cc_2456 ( N_noxref_5_c_2513_n N_RN_c_6037_n ) capacitor c=0.00834532f \
 //x=18.57 //y=1.915 //x2=20.07 //y2=1.915
cc_2457 ( N_noxref_5_c_2498_n N_RN_c_6039_n ) capacitor c=0.00183762f \
 //x=18.87 //y=2.08 //x2=19.98 //y2=4.7
cc_2458 ( N_noxref_5_c_2630_p N_RN_c_6039_n ) capacitor c=0.0168581f \
 //x=19.435 //y=4.79 //x2=19.98 //y2=4.7
cc_2459 ( N_noxref_5_c_2551_n N_RN_c_6039_n ) capacitor c=0.00484466f \
 //x=19.145 //y=4.79 //x2=19.98 //y2=4.7
cc_2460 ( N_noxref_5_c_2498_n N_noxref_20_c_8538_n ) capacitor c=0.0013672f \
 //x=18.87 //y=2.08 //x2=21.09 //y2=2.08
cc_2461 ( N_noxref_5_M2_noxref_d N_noxref_23_M0_noxref_s ) capacitor \
 c=0.00309936f //x=3.395 //y=0.915 //x2=0.455 //y2=0.375
cc_2462 ( N_noxref_5_c_2496_n N_noxref_24_c_9317_n ) capacitor c=0.00466084f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_2463 ( N_noxref_5_M2_noxref_d N_noxref_24_c_9317_n ) capacitor c=0.0117786f \
 //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_2464 ( N_noxref_5_c_2583_n N_noxref_24_c_9330_n ) capacitor c=0.0200405f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_2465 ( N_noxref_5_M2_noxref_d N_noxref_24_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_2466 ( N_noxref_5_c_2496_n N_noxref_24_M2_noxref_s ) capacitor c=0.0207678f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_2467 ( N_noxref_5_M2_noxref_d N_noxref_24_M2_noxref_s ) capacitor \
 c=0.0426368f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
cc_2468 ( N_noxref_5_c_2496_n N_noxref_25_c_9379_n ) capacitor c=3.84569e-19 \
 //x=3.985 //y=1.665 //x2=5.4 //y2=1.505
cc_2469 ( N_noxref_5_c_2503_n N_noxref_25_c_9379_n ) capacitor c=0.0034165f \
 //x=5.62 //y=1.915 //x2=5.4 //y2=1.505
cc_2470 ( N_noxref_5_c_2497_n N_noxref_25_c_9364_n ) capacitor c=0.0125801f \
 //x=5.92 //y=2.08 //x2=6.285 //y2=1.59
cc_2471 ( N_noxref_5_c_2502_n N_noxref_25_c_9364_n ) capacitor c=0.00703864f \
 //x=5.62 //y=1.53 //x2=6.285 //y2=1.59
cc_2472 ( N_noxref_5_c_2503_n N_noxref_25_c_9364_n ) capacitor c=0.0245895f \
 //x=5.62 //y=1.915 //x2=6.285 //y2=1.59
cc_2473 ( N_noxref_5_c_2505_n N_noxref_25_c_9364_n ) capacitor c=0.00708583f \
 //x=5.995 //y=1.375 //x2=6.285 //y2=1.59
cc_2474 ( N_noxref_5_c_2508_n N_noxref_25_c_9364_n ) capacitor c=0.00698822f \
 //x=6.15 //y=1.22 //x2=6.285 //y2=1.59
cc_2475 ( N_noxref_5_c_2499_n N_noxref_25_M3_noxref_s ) capacitor c=0.0327271f \
 //x=5.62 //y=0.875 //x2=5.265 //y2=0.375
cc_2476 ( N_noxref_5_c_2502_n N_noxref_25_M3_noxref_s ) capacitor \
 c=7.99997e-19 //x=5.62 //y=1.53 //x2=5.265 //y2=0.375
cc_2477 ( N_noxref_5_c_2503_n N_noxref_25_M3_noxref_s ) capacitor \
 c=0.00122123f //x=5.62 //y=1.915 //x2=5.265 //y2=0.375
cc_2478 ( N_noxref_5_c_2506_n N_noxref_25_M3_noxref_s ) capacitor c=0.0121427f \
 //x=6.15 //y=0.875 //x2=5.265 //y2=0.375
cc_2479 ( N_noxref_5_M2_noxref_d N_noxref_25_M3_noxref_s ) capacitor \
 c=2.55333e-19 //x=3.395 //y=0.915 //x2=5.265 //y2=0.375
cc_2480 ( N_noxref_5_c_2513_n N_noxref_30_c_9637_n ) capacitor c=0.0034165f \
 //x=18.57 //y=1.915 //x2=18.35 //y2=1.505
cc_2481 ( N_noxref_5_c_2498_n N_noxref_30_c_9622_n ) capacitor c=0.0115578f \
 //x=18.87 //y=2.08 //x2=19.235 //y2=1.59
cc_2482 ( N_noxref_5_c_2512_n N_noxref_30_c_9622_n ) capacitor c=0.00697148f \
 //x=18.57 //y=1.53 //x2=19.235 //y2=1.59
cc_2483 ( N_noxref_5_c_2513_n N_noxref_30_c_9622_n ) capacitor c=0.0204849f \
 //x=18.57 //y=1.915 //x2=19.235 //y2=1.59
cc_2484 ( N_noxref_5_c_2515_n N_noxref_30_c_9622_n ) capacitor c=0.00610316f \
 //x=18.945 //y=1.375 //x2=19.235 //y2=1.59
cc_2485 ( N_noxref_5_c_2518_n N_noxref_30_c_9622_n ) capacitor c=0.00698822f \
 //x=19.1 //y=1.22 //x2=19.235 //y2=1.59
cc_2486 ( N_noxref_5_c_2509_n N_noxref_30_M11_noxref_s ) capacitor \
 c=0.0327271f //x=18.57 //y=0.875 //x2=18.215 //y2=0.375
cc_2487 ( N_noxref_5_c_2512_n N_noxref_30_M11_noxref_s ) capacitor \
 c=7.99997e-19 //x=18.57 //y=1.53 //x2=18.215 //y2=0.375
cc_2488 ( N_noxref_5_c_2513_n N_noxref_30_M11_noxref_s ) capacitor \
 c=0.00122123f //x=18.57 //y=1.915 //x2=18.215 //y2=0.375
cc_2489 ( N_noxref_5_c_2516_n N_noxref_30_M11_noxref_s ) capacitor \
 c=0.0121427f //x=19.1 //y=0.875 //x2=18.215 //y2=0.375
cc_2490 ( N_noxref_6_c_2975_p N_noxref_11_c_4077_n ) capacitor c=0.00648968f \
 //x=24.305 //y=4.07 //x2=27.125 //y2=4.07
cc_2491 ( N_noxref_6_c_2756_n N_noxref_11_c_4058_n ) capacitor c=8.45344e-19 \
 //x=24.42 //y=2.08 //x2=27.01 //y2=2.08
cc_2492 ( N_noxref_6_c_2748_n N_D_c_4434_n ) capacitor c=0.00334753f \
 //x=11.355 //y=4.07 //x2=32.815 //y2=2.59
cc_2493 ( N_noxref_6_c_2787_n N_D_c_4434_n ) capacitor c=0.0188674f //x=16.905 \
 //y=4.07 //x2=32.815 //y2=2.59
cc_2494 ( N_noxref_6_c_2891_n N_D_c_4434_n ) capacitor c=3.04562e-19 \
 //x=11.585 //y=4.07 //x2=32.815 //y2=2.59
cc_2495 ( N_noxref_6_c_2788_n N_D_c_4434_n ) capacitor c=0.0497112f //x=21.715 \
 //y=4.07 //x2=32.815 //y2=2.59
cc_2496 ( N_noxref_6_c_2789_n N_D_c_4434_n ) capacitor c=3.16222e-19 \
 //x=17.135 //y=4.07 //x2=32.815 //y2=2.59
cc_2497 ( N_noxref_6_c_2790_n N_D_c_4434_n ) capacitor c=0.00467819f \
 //x=23.565 //y=4.07 //x2=32.815 //y2=2.59
cc_2498 ( N_noxref_6_c_2791_n N_D_c_4434_n ) capacitor c=2.97275e-19 \
 //x=21.945 //y=4.07 //x2=32.815 //y2=2.59
cc_2499 ( N_noxref_6_c_2975_p N_D_c_4434_n ) capacitor c=0.00410116f \
 //x=24.305 //y=4.07 //x2=32.815 //y2=2.59
cc_2500 ( N_noxref_6_c_2792_n N_D_c_4434_n ) capacitor c=3.35912e-19 \
 //x=23.795 //y=4.07 //x2=32.815 //y2=2.59
cc_2501 ( N_noxref_6_c_2751_n N_D_c_4434_n ) capacitor c=0.0207818f //x=11.47 \
 //y=2.08 //x2=32.815 //y2=2.59
cc_2502 ( N_noxref_6_c_2812_n N_D_c_4434_n ) capacitor c=0.0204505f //x=17.02 \
 //y=4.07 //x2=32.815 //y2=2.59
cc_2503 ( N_noxref_6_c_2827_n N_D_c_4434_n ) capacitor c=0.0165903f //x=21.83 \
 //y=4.07 //x2=32.815 //y2=2.59
cc_2504 ( N_noxref_6_c_2755_n N_D_c_4434_n ) capacitor c=0.0177889f //x=23.68 \
 //y=2.08 //x2=32.815 //y2=2.59
cc_2505 ( N_noxref_6_c_2756_n N_D_c_4434_n ) capacitor c=0.0169241f //x=24.42 \
 //y=2.08 //x2=32.815 //y2=2.59
cc_2506 ( N_noxref_6_c_2748_n N_D_c_4448_n ) capacitor c=0.0190126f //x=11.355 \
 //y=4.07 //x2=7.03 //y2=2.08
cc_2507 ( N_noxref_6_c_2748_n N_CLK_c_4808_n ) capacitor c=0.784553f \
 //x=11.355 //y=4.07 //x2=15.055 //y2=4.44
cc_2508 ( N_noxref_6_c_2787_n N_CLK_c_4808_n ) capacitor c=0.302855f \
 //x=16.905 //y=4.07 //x2=15.055 //y2=4.44
cc_2509 ( N_noxref_6_c_2891_n N_CLK_c_4808_n ) capacitor c=0.0263375f \
 //x=11.585 //y=4.07 //x2=15.055 //y2=4.44
cc_2510 ( N_noxref_6_c_2893_n N_CLK_c_4808_n ) capacitor c=0.0016972f \
 //x=11.47 //y=4.535 //x2=15.055 //y2=4.44
cc_2511 ( N_noxref_6_c_2751_n N_CLK_c_4808_n ) capacitor c=0.0207534f \
 //x=11.47 //y=2.08 //x2=15.055 //y2=4.44
cc_2512 ( N_noxref_6_c_2802_n N_CLK_c_4808_n ) capacitor c=0.0219114f \
 //x=14.565 //y=5.155 //x2=15.055 //y2=4.44
cc_2513 ( N_noxref_6_c_2937_n N_CLK_c_4808_n ) capacitor c=0.00960248f \
 //x=11.875 //y=4.79 //x2=15.055 //y2=4.44
cc_2514 ( N_noxref_6_c_2914_n N_CLK_c_4808_n ) capacitor c=0.00203982f \
 //x=11.5 //y=4.7 //x2=15.055 //y2=4.44
cc_2515 ( N_noxref_6_c_2748_n N_CLK_c_4825_n ) capacitor c=0.0291328f \
 //x=11.355 //y=4.07 //x2=2.335 //y2=4.44
cc_2516 ( N_noxref_6_c_2750_n N_CLK_c_4825_n ) capacitor c=0.00551083f \
 //x=1.11 //y=2.08 //x2=2.335 //y2=4.44
cc_2517 ( N_noxref_6_c_2787_n N_CLK_c_4826_n ) capacitor c=0.140035f \
 //x=16.905 //y=4.07 //x2=28.005 //y2=4.44
cc_2518 ( N_noxref_6_c_2788_n N_CLK_c_4826_n ) capacitor c=0.398434f \
 //x=21.715 //y=4.07 //x2=28.005 //y2=4.44
cc_2519 ( N_noxref_6_c_2789_n N_CLK_c_4826_n ) capacitor c=0.0265915f \
 //x=17.135 //y=4.07 //x2=28.005 //y2=4.44
cc_2520 ( N_noxref_6_c_2790_n N_CLK_c_4826_n ) capacitor c=0.143555f \
 //x=23.565 //y=4.07 //x2=28.005 //y2=4.44
cc_2521 ( N_noxref_6_c_2791_n N_CLK_c_4826_n ) capacitor c=0.0265915f \
 //x=21.945 //y=4.07 //x2=28.005 //y2=4.44
cc_2522 ( N_noxref_6_c_2975_p N_CLK_c_4826_n ) capacitor c=0.073184f \
 //x=24.305 //y=4.07 //x2=28.005 //y2=4.44
cc_2523 ( N_noxref_6_c_2792_n N_CLK_c_4826_n ) capacitor c=0.0263778f \
 //x=23.795 //y=4.07 //x2=28.005 //y2=4.44
cc_2524 ( N_noxref_6_c_2808_n N_CLK_c_4826_n ) capacitor c=0.0183122f \
 //x=16.935 //y=5.155 //x2=28.005 //y2=4.44
cc_2525 ( N_noxref_6_c_2812_n N_CLK_c_4826_n ) capacitor c=0.022862f //x=17.02 \
 //y=4.07 //x2=28.005 //y2=4.44
cc_2526 ( N_noxref_6_c_2813_n N_CLK_c_4826_n ) capacitor c=0.032141f \
 //x=20.085 //y=5.155 //x2=28.005 //y2=4.44
cc_2527 ( N_noxref_6_c_2817_n N_CLK_c_4826_n ) capacitor c=0.0230136f \
 //x=19.375 //y=5.155 //x2=28.005 //y2=4.44
cc_2528 ( N_noxref_6_c_2823_n N_CLK_c_4826_n ) capacitor c=0.0183122f \
 //x=21.745 //y=5.155 //x2=28.005 //y2=4.44
cc_2529 ( N_noxref_6_c_2827_n N_CLK_c_4826_n ) capacitor c=0.022862f //x=21.83 \
 //y=4.07 //x2=28.005 //y2=4.44
cc_2530 ( N_noxref_6_c_2755_n N_CLK_c_4826_n ) capacitor c=0.0216667f \
 //x=23.68 //y=2.08 //x2=28.005 //y2=4.44
cc_2531 ( N_noxref_6_c_3016_p N_CLK_c_4826_n ) capacitor c=0.0016972f \
 //x=24.42 //y=4.535 //x2=28.005 //y2=4.44
cc_2532 ( N_noxref_6_c_2756_n N_CLK_c_4826_n ) capacitor c=0.0207552f \
 //x=24.42 //y=2.08 //x2=28.005 //y2=4.44
cc_2533 ( N_noxref_6_c_3018_p N_CLK_c_4826_n ) capacitor c=0.0311227f \
 //x=15.36 //y=5.155 //x2=28.005 //y2=4.44
cc_2534 ( N_noxref_6_c_3019_p N_CLK_c_4826_n ) capacitor c=0.00720343f \
 //x=24.825 //y=4.79 //x2=28.005 //y2=4.44
cc_2535 ( N_noxref_6_c_2853_n N_CLK_c_4826_n ) capacitor c=0.0107036f \
 //x=23.68 //y=4.7 //x2=28.005 //y2=4.44
cc_2536 ( N_noxref_6_c_3021_p N_CLK_c_4826_n ) capacitor c=0.0019199f \
 //x=24.45 //y=4.7 //x2=28.005 //y2=4.44
cc_2537 ( N_noxref_6_c_2787_n N_CLK_c_4843_n ) capacitor c=0.026534f \
 //x=16.905 //y=4.07 //x2=15.285 //y2=4.44
cc_2538 ( N_noxref_6_c_2798_n N_CLK_c_4843_n ) capacitor c=0.00241768f \
 //x=15.275 //y=5.155 //x2=15.285 //y2=4.44
cc_2539 ( N_noxref_6_c_2748_n N_CLK_c_4802_n ) capacitor c=0.0265867f \
 //x=11.355 //y=4.07 //x2=2.22 //y2=2.08
cc_2540 ( N_noxref_6_c_2749_n N_CLK_c_4802_n ) capacitor c=0.00128547f \
 //x=1.225 //y=4.07 //x2=2.22 //y2=2.08
cc_2541 ( N_noxref_6_c_2750_n N_CLK_c_4802_n ) capacitor c=0.0535714f //x=1.11 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_2542 ( N_noxref_6_c_2762_n N_CLK_c_4802_n ) capacitor c=0.00238338f \
 //x=0.81 //y=1.915 //x2=2.22 //y2=2.08
cc_2543 ( N_noxref_6_c_2973_n N_CLK_c_4802_n ) capacitor c=0.00147352f \
 //x=1.675 //y=4.79 //x2=2.22 //y2=2.08
cc_2544 ( N_noxref_6_c_2851_n N_CLK_c_4802_n ) capacitor c=0.00141297f \
 //x=1.385 //y=4.79 //x2=2.22 //y2=2.08
cc_2545 ( N_noxref_6_c_2787_n N_CLK_c_4803_n ) capacitor c=0.0208526f \
 //x=16.905 //y=4.07 //x2=15.17 //y2=2.08
cc_2546 ( N_noxref_6_c_2798_n N_CLK_c_4803_n ) capacitor c=0.0143918f \
 //x=15.275 //y=5.155 //x2=15.17 //y2=2.08
cc_2547 ( N_noxref_6_c_2812_n N_CLK_c_4803_n ) capacitor c=0.00272321f \
 //x=17.02 //y=4.07 //x2=15.17 //y2=2.08
cc_2548 ( N_noxref_6_M54_noxref_g N_CLK_M56_noxref_g ) capacitor c=0.0105869f \
 //x=1.31 //y=6.02 //x2=2.19 //y2=6.02
cc_2549 ( N_noxref_6_M55_noxref_g N_CLK_M56_noxref_g ) capacitor c=0.10632f \
 //x=1.75 //y=6.02 //x2=2.19 //y2=6.02
cc_2550 ( N_noxref_6_M55_noxref_g N_CLK_M57_noxref_g ) capacitor c=0.0101598f \
 //x=1.75 //y=6.02 //x2=2.63 //y2=6.02
cc_2551 ( N_noxref_6_c_2798_n N_CLK_M72_noxref_g ) capacitor c=0.016514f \
 //x=15.275 //y=5.155 //x2=15.14 //y2=6.02
cc_2552 ( N_noxref_6_M72_noxref_d N_CLK_M72_noxref_g ) capacitor c=0.0180032f \
 //x=15.215 //y=5.02 //x2=15.14 //y2=6.02
cc_2553 ( N_noxref_6_c_2804_n N_CLK_M73_noxref_g ) capacitor c=0.01736f \
 //x=16.155 //y=5.155 //x2=15.58 //y2=6.02
cc_2554 ( N_noxref_6_M72_noxref_d N_CLK_M73_noxref_g ) capacitor c=0.0180032f \
 //x=15.215 //y=5.02 //x2=15.58 //y2=6.02
cc_2555 ( N_noxref_6_c_2758_n N_CLK_c_5060_n ) capacitor c=5.72482e-19 \
 //x=0.81 //y=0.875 //x2=1.785 //y2=0.91
cc_2556 ( N_noxref_6_c_2760_n N_CLK_c_5060_n ) capacitor c=0.00149976f \
 //x=0.81 //y=1.22 //x2=1.785 //y2=0.91
cc_2557 ( N_noxref_6_c_2765_n N_CLK_c_5060_n ) capacitor c=0.0160123f //x=1.34 \
 //y=0.875 //x2=1.785 //y2=0.91
cc_2558 ( N_noxref_6_c_2761_n N_CLK_c_5063_n ) capacitor c=0.00111227f \
 //x=0.81 //y=1.53 //x2=1.785 //y2=1.22
cc_2559 ( N_noxref_6_c_2767_n N_CLK_c_5063_n ) capacitor c=0.0124075f //x=1.34 \
 //y=1.22 //x2=1.785 //y2=1.22
cc_2560 ( N_noxref_6_c_2765_n N_CLK_c_4952_n ) capacitor c=0.00103227f \
 //x=1.34 //y=0.875 //x2=2.31 //y2=0.91
cc_2561 ( N_noxref_6_c_2767_n N_CLK_c_4953_n ) capacitor c=0.0010154f //x=1.34 \
 //y=1.22 //x2=2.31 //y2=1.22
cc_2562 ( N_noxref_6_c_2767_n N_CLK_c_4954_n ) capacitor c=9.23422e-19 \
 //x=1.34 //y=1.22 //x2=2.31 //y2=1.45
cc_2563 ( N_noxref_6_c_2750_n N_CLK_c_4955_n ) capacitor c=0.00231304f \
 //x=1.11 //y=2.08 //x2=2.31 //y2=1.915
cc_2564 ( N_noxref_6_c_2762_n N_CLK_c_4955_n ) capacitor c=0.00964411f \
 //x=0.81 //y=1.915 //x2=2.31 //y2=1.915
cc_2565 ( N_noxref_6_c_3018_p N_CLK_c_5070_n ) capacitor c=0.00426767f \
 //x=15.36 //y=5.155 //x2=15.505 //y2=4.79
cc_2566 ( N_noxref_6_c_2748_n N_CLK_c_4959_n ) capacitor c=6.38735e-19 \
 //x=11.355 //y=4.07 //x2=2.22 //y2=4.7
cc_2567 ( N_noxref_6_c_2750_n N_CLK_c_4959_n ) capacitor c=0.00183762f \
 //x=1.11 //y=2.08 //x2=2.22 //y2=4.7
cc_2568 ( N_noxref_6_c_2973_n N_CLK_c_4959_n ) capacitor c=0.0168581f \
 //x=1.675 //y=4.79 //x2=2.22 //y2=4.7
cc_2569 ( N_noxref_6_c_2851_n N_CLK_c_4959_n ) capacitor c=0.00484466f \
 //x=1.385 //y=4.79 //x2=2.22 //y2=4.7
cc_2570 ( N_noxref_6_c_2798_n N_CLK_c_4986_n ) capacitor c=0.00322046f \
 //x=15.275 //y=5.155 //x2=15.17 //y2=4.7
cc_2571 ( N_noxref_6_c_2751_n N_RN_c_5846_n ) capacitor c=0.0178519f //x=11.47 \
 //y=2.08 //x2=16.165 //y2=2.22
cc_2572 ( N_noxref_6_c_2940_n N_RN_c_5846_n ) capacitor c=3.11115e-19 \
 //x=11.88 //y=1.405 //x2=16.165 //y2=2.22
cc_2573 ( N_noxref_6_c_2912_n N_RN_c_5846_n ) capacitor c=0.00570799f \
 //x=11.47 //y=2.08 //x2=16.165 //y2=2.22
cc_2574 ( N_noxref_6_c_2788_n N_RN_c_5856_n ) capacitor c=0.00501936f \
 //x=21.715 //y=4.07 //x2=19.865 //y2=2.22
cc_2575 ( N_noxref_6_c_3060_p N_RN_c_5856_n ) capacitor c=0.016327f //x=16.62 \
 //y=1.665 //x2=19.865 //y2=2.22
cc_2576 ( N_noxref_6_c_2812_n N_RN_c_5856_n ) capacitor c=0.0197307f //x=17.02 \
 //y=4.07 //x2=19.865 //y2=2.22
cc_2577 ( N_noxref_6_c_2812_n N_RN_c_5860_n ) capacitor c=0.0012045f //x=17.02 \
 //y=4.07 //x2=16.395 //y2=2.22
cc_2578 ( N_noxref_6_c_2788_n N_RN_c_5861_n ) capacitor c=0.00559167f \
 //x=21.715 //y=4.07 //x2=33.925 //y2=2.22
cc_2579 ( N_noxref_6_c_3064_p N_RN_c_5861_n ) capacitor c=0.016327f //x=21.43 \
 //y=1.665 //x2=33.925 //y2=2.22
cc_2580 ( N_noxref_6_c_2827_n N_RN_c_5861_n ) capacitor c=0.0197307f //x=21.83 \
 //y=4.07 //x2=33.925 //y2=2.22
cc_2581 ( N_noxref_6_c_2755_n N_RN_c_5861_n ) capacitor c=0.0185072f //x=23.68 \
 //y=2.08 //x2=33.925 //y2=2.22
cc_2582 ( N_noxref_6_c_2756_n N_RN_c_5861_n ) capacitor c=0.0178578f //x=24.42 \
 //y=2.08 //x2=33.925 //y2=2.22
cc_2583 ( N_noxref_6_c_2772_n N_RN_c_5861_n ) capacitor c=0.00892609f \
 //x=23.485 //y=1.915 //x2=33.925 //y2=2.22
cc_2584 ( N_noxref_6_c_3069_p N_RN_c_5861_n ) capacitor c=3.11115e-19 \
 //x=24.83 //y=1.405 //x2=33.925 //y2=2.22
cc_2585 ( N_noxref_6_c_3070_p N_RN_c_5861_n ) capacitor c=0.00569252f \
 //x=24.42 //y=2.08 //x2=33.925 //y2=2.22
cc_2586 ( N_noxref_6_c_2788_n N_RN_c_5872_n ) capacitor c=4.24963e-19 \
 //x=21.715 //y=4.07 //x2=20.095 //y2=2.22
cc_2587 ( N_noxref_6_c_2748_n N_RN_c_5913_n ) capacitor c=0.0179722f \
 //x=11.355 //y=4.07 //x2=8.14 //y2=2.08
cc_2588 ( N_noxref_6_c_2787_n N_RN_c_5914_n ) capacitor c=0.0179722f \
 //x=16.905 //y=4.07 //x2=16.28 //y2=2.08
cc_2589 ( N_noxref_6_c_2789_n N_RN_c_5914_n ) capacitor c=0.00179385f \
 //x=17.135 //y=4.07 //x2=16.28 //y2=2.08
cc_2590 ( N_noxref_6_c_2812_n N_RN_c_5914_n ) capacitor c=0.0801183f //x=17.02 \
 //y=4.07 //x2=16.28 //y2=2.08
cc_2591 ( N_noxref_6_c_3076_p N_RN_c_5914_n ) capacitor c=0.0171303f //x=16.24 \
 //y=5.155 //x2=16.28 //y2=2.08
cc_2592 ( N_noxref_6_c_2788_n N_RN_c_5915_n ) capacitor c=0.023857f //x=21.715 \
 //y=4.07 //x2=19.98 //y2=2.08
cc_2593 ( N_noxref_6_c_2812_n N_RN_c_5915_n ) capacitor c=7.03136e-19 \
 //x=17.02 //y=4.07 //x2=19.98 //y2=2.08
cc_2594 ( N_noxref_6_c_2813_n N_RN_c_5915_n ) capacitor c=0.0144268f \
 //x=20.085 //y=5.155 //x2=19.98 //y2=2.08
cc_2595 ( N_noxref_6_c_2827_n N_RN_c_5915_n ) capacitor c=0.00295341f \
 //x=21.83 //y=4.07 //x2=19.98 //y2=2.08
cc_2596 ( N_noxref_6_c_2804_n N_RN_M74_noxref_g ) capacitor c=0.01736f \
 //x=16.155 //y=5.155 //x2=16.02 //y2=6.02
cc_2597 ( N_noxref_6_M74_noxref_d N_RN_M74_noxref_g ) capacitor c=0.0180032f \
 //x=16.095 //y=5.02 //x2=16.02 //y2=6.02
cc_2598 ( N_noxref_6_c_2808_n N_RN_M75_noxref_g ) capacitor c=0.0194981f \
 //x=16.935 //y=5.155 //x2=16.46 //y2=6.02
cc_2599 ( N_noxref_6_M74_noxref_d N_RN_M75_noxref_g ) capacitor c=0.0194246f \
 //x=16.095 //y=5.02 //x2=16.46 //y2=6.02
cc_2600 ( N_noxref_6_c_2813_n N_RN_M78_noxref_g ) capacitor c=0.0165266f \
 //x=20.085 //y=5.155 //x2=19.95 //y2=6.02
cc_2601 ( N_noxref_6_M78_noxref_d N_RN_M78_noxref_g ) capacitor c=0.0180032f \
 //x=20.025 //y=5.02 //x2=19.95 //y2=6.02
cc_2602 ( N_noxref_6_c_2819_n N_RN_M79_noxref_g ) capacitor c=0.01736f \
 //x=20.965 //y=5.155 //x2=20.39 //y2=6.02
cc_2603 ( N_noxref_6_M78_noxref_d N_RN_M79_noxref_g ) capacitor c=0.0180032f \
 //x=20.025 //y=5.02 //x2=20.39 //y2=6.02
cc_2604 ( N_noxref_6_M10_noxref_d N_RN_c_6075_n ) capacitor c=0.00217566f \
 //x=16.345 //y=0.915 //x2=16.27 //y2=0.915
cc_2605 ( N_noxref_6_M10_noxref_d N_RN_c_6076_n ) capacitor c=0.0034598f \
 //x=16.345 //y=0.915 //x2=16.27 //y2=1.26
cc_2606 ( N_noxref_6_M10_noxref_d N_RN_c_6077_n ) capacitor c=0.00546784f \
 //x=16.345 //y=0.915 //x2=16.27 //y2=1.57
cc_2607 ( N_noxref_6_M10_noxref_d N_RN_c_6078_n ) capacitor c=0.00241102f \
 //x=16.345 //y=0.915 //x2=16.645 //y2=0.76
cc_2608 ( N_noxref_6_c_2753_n N_RN_c_6079_n ) capacitor c=0.00371277f \
 //x=16.935 //y=1.665 //x2=16.645 //y2=1.415
cc_2609 ( N_noxref_6_M10_noxref_d N_RN_c_6079_n ) capacitor c=0.0138621f \
 //x=16.345 //y=0.915 //x2=16.645 //y2=1.415
cc_2610 ( N_noxref_6_M10_noxref_d N_RN_c_6081_n ) capacitor c=0.00219619f \
 //x=16.345 //y=0.915 //x2=16.8 //y2=0.915
cc_2611 ( N_noxref_6_c_2753_n N_RN_c_6082_n ) capacitor c=0.00457401f \
 //x=16.935 //y=1.665 //x2=16.8 //y2=1.26
cc_2612 ( N_noxref_6_M10_noxref_d N_RN_c_6082_n ) capacitor c=0.00603828f \
 //x=16.345 //y=0.915 //x2=16.8 //y2=1.26
cc_2613 ( N_noxref_6_c_3098_p N_RN_c_6084_n ) capacitor c=0.00426767f \
 //x=20.17 //y=5.155 //x2=20.315 //y2=4.79
cc_2614 ( N_noxref_6_c_2812_n N_RN_c_6085_n ) capacitor c=0.00709342f \
 //x=17.02 //y=4.07 //x2=16.28 //y2=2.08
cc_2615 ( N_noxref_6_c_2812_n N_RN_c_6086_n ) capacitor c=0.00283672f \
 //x=17.02 //y=4.07 //x2=16.28 //y2=1.915
cc_2616 ( N_noxref_6_M10_noxref_d N_RN_c_6086_n ) capacitor c=0.00661782f \
 //x=16.345 //y=0.915 //x2=16.28 //y2=1.915
cc_2617 ( N_noxref_6_c_2808_n N_RN_c_6088_n ) capacitor c=0.00201851f \
 //x=16.935 //y=5.155 //x2=16.28 //y2=4.7
cc_2618 ( N_noxref_6_c_2812_n N_RN_c_6088_n ) capacitor c=0.013693f //x=17.02 \
 //y=4.07 //x2=16.28 //y2=4.7
cc_2619 ( N_noxref_6_c_3076_p N_RN_c_6088_n ) capacitor c=0.00475601f \
 //x=16.24 //y=5.155 //x2=16.28 //y2=4.7
cc_2620 ( N_noxref_6_c_2813_n N_RN_c_6039_n ) capacitor c=0.00322054f \
 //x=20.085 //y=5.155 //x2=19.98 //y2=4.7
cc_2621 ( N_noxref_6_c_2788_n N_noxref_20_c_8515_n ) capacitor c=0.0142808f \
 //x=21.715 //y=4.07 //x2=25.045 //y2=2.96
cc_2622 ( N_noxref_6_c_2790_n N_noxref_20_c_8515_n ) capacitor c=0.0512827f \
 //x=23.565 //y=4.07 //x2=25.045 //y2=2.96
cc_2623 ( N_noxref_6_c_2791_n N_noxref_20_c_8515_n ) capacitor c=0.00700854f \
 //x=21.945 //y=4.07 //x2=25.045 //y2=2.96
cc_2624 ( N_noxref_6_c_2975_p N_noxref_20_c_8515_n ) capacitor c=0.022067f \
 //x=24.305 //y=4.07 //x2=25.045 //y2=2.96
cc_2625 ( N_noxref_6_c_2792_n N_noxref_20_c_8515_n ) capacitor c=0.0068108f \
 //x=23.795 //y=4.07 //x2=25.045 //y2=2.96
cc_2626 ( N_noxref_6_c_2827_n N_noxref_20_c_8515_n ) capacitor c=0.0227185f \
 //x=21.83 //y=4.07 //x2=25.045 //y2=2.96
cc_2627 ( N_noxref_6_c_2755_n N_noxref_20_c_8515_n ) capacitor c=0.0226688f \
 //x=23.68 //y=2.08 //x2=25.045 //y2=2.96
cc_2628 ( N_noxref_6_c_2756_n N_noxref_20_c_8515_n ) capacitor c=0.0209033f \
 //x=24.42 //y=2.08 //x2=25.045 //y2=2.96
cc_2629 ( N_noxref_6_c_2788_n N_noxref_20_c_8606_n ) capacitor c=0.00780534f \
 //x=21.715 //y=4.07 //x2=21.205 //y2=2.96
cc_2630 ( N_noxref_6_c_2827_n N_noxref_20_c_8606_n ) capacitor c=0.00117715f \
 //x=21.83 //y=4.07 //x2=21.205 //y2=2.96
cc_2631 ( N_noxref_6_c_2756_n N_noxref_20_c_8608_n ) capacitor c=0.00117715f \
 //x=24.42 //y=2.08 //x2=25.275 //y2=2.96
cc_2632 ( N_noxref_6_c_2788_n N_noxref_20_c_8538_n ) capacitor c=0.0219251f \
 //x=21.715 //y=4.07 //x2=21.09 //y2=2.08
cc_2633 ( N_noxref_6_c_2791_n N_noxref_20_c_8538_n ) capacitor c=0.00131333f \
 //x=21.945 //y=4.07 //x2=21.09 //y2=2.08
cc_2634 ( N_noxref_6_c_2827_n N_noxref_20_c_8538_n ) capacitor c=0.0801459f \
 //x=21.83 //y=4.07 //x2=21.09 //y2=2.08
cc_2635 ( N_noxref_6_c_2755_n N_noxref_20_c_8538_n ) capacitor c=7.99641e-19 \
 //x=23.68 //y=2.08 //x2=21.09 //y2=2.08
cc_2636 ( N_noxref_6_c_3121_p N_noxref_20_c_8538_n ) capacitor c=0.0171303f \
 //x=21.05 //y=5.155 //x2=21.09 //y2=2.08
cc_2637 ( N_noxref_6_c_3016_p N_noxref_20_c_8560_n ) capacitor c=0.0126603f \
 //x=24.42 //y=4.535 //x2=24.595 //y2=5.2
cc_2638 ( N_noxref_6_M83_noxref_g N_noxref_20_c_8560_n ) capacitor \
 c=0.0169686f //x=24.02 //y=6.02 //x2=24.595 //y2=5.2
cc_2639 ( N_noxref_6_M84_noxref_g N_noxref_20_c_8560_n ) capacitor \
 c=0.0166421f //x=24.46 //y=6.02 //x2=24.595 //y2=5.2
cc_2640 ( N_noxref_6_c_3021_p N_noxref_20_c_8560_n ) capacitor c=0.00346527f \
 //x=24.45 //y=4.7 //x2=24.595 //y2=5.2
cc_2641 ( N_noxref_6_c_2755_n N_noxref_20_c_8564_n ) capacitor c=0.00521572f \
 //x=23.68 //y=2.08 //x2=23.885 //y2=5.2
cc_2642 ( N_noxref_6_M82_noxref_g N_noxref_20_c_8564_n ) capacitor \
 c=0.0177326f //x=23.58 //y=6.02 //x2=23.885 //y2=5.2
cc_2643 ( N_noxref_6_c_2853_n N_noxref_20_c_8564_n ) capacitor c=0.00581252f \
 //x=23.68 //y=4.7 //x2=23.885 //y2=5.2
cc_2644 ( N_noxref_6_M85_noxref_g N_noxref_20_c_8566_n ) capacitor c=0.018922f \
 //x=24.9 //y=6.02 //x2=25.075 //y2=5.2
cc_2645 ( N_noxref_6_c_3069_p N_noxref_20_c_8539_n ) capacitor c=0.00371277f \
 //x=24.83 //y=1.405 //x2=25.075 //y2=1.655
cc_2646 ( N_noxref_6_c_3131_p N_noxref_20_c_8539_n ) capacitor c=0.00457401f \
 //x=24.985 //y=1.25 //x2=25.075 //y2=1.655
cc_2647 ( N_noxref_6_c_2975_p N_noxref_20_c_8540_n ) capacitor c=0.00423741f \
 //x=24.305 //y=4.07 //x2=25.16 //y2=2.96
cc_2648 ( N_noxref_6_c_2827_n N_noxref_20_c_8540_n ) capacitor c=3.52729e-19 \
 //x=21.83 //y=4.07 //x2=25.16 //y2=2.96
cc_2649 ( N_noxref_6_c_2755_n N_noxref_20_c_8540_n ) capacitor c=0.00318426f \
 //x=23.68 //y=2.08 //x2=25.16 //y2=2.96
cc_2650 ( N_noxref_6_c_3016_p N_noxref_20_c_8540_n ) capacitor c=0.0101115f \
 //x=24.42 //y=4.535 //x2=25.16 //y2=2.96
cc_2651 ( N_noxref_6_c_2756_n N_noxref_20_c_8540_n ) capacitor c=0.0723476f \
 //x=24.42 //y=2.08 //x2=25.16 //y2=2.96
cc_2652 ( N_noxref_6_c_3019_p N_noxref_20_c_8540_n ) capacitor c=0.0142673f \
 //x=24.825 //y=4.79 //x2=25.16 //y2=2.96
cc_2653 ( N_noxref_6_c_3070_p N_noxref_20_c_8540_n ) capacitor c=0.00731987f \
 //x=24.42 //y=2.08 //x2=25.16 //y2=2.96
cc_2654 ( N_noxref_6_c_3139_p N_noxref_20_c_8540_n ) capacitor c=0.00306024f \
 //x=24.42 //y=1.915 //x2=25.16 //y2=2.96
cc_2655 ( N_noxref_6_c_3021_p N_noxref_20_c_8540_n ) capacitor c=0.00517969f \
 //x=24.45 //y=4.7 //x2=25.16 //y2=2.96
cc_2656 ( N_noxref_6_c_3019_p N_noxref_20_c_8633_n ) capacitor c=0.00407665f \
 //x=24.825 //y=4.79 //x2=24.68 //y2=5.2
cc_2657 ( N_noxref_6_c_2819_n N_noxref_20_M80_noxref_g ) capacitor c=0.01736f \
 //x=20.965 //y=5.155 //x2=20.83 //y2=6.02
cc_2658 ( N_noxref_6_M80_noxref_d N_noxref_20_M80_noxref_g ) capacitor \
 c=0.0180032f //x=20.905 //y=5.02 //x2=20.83 //y2=6.02
cc_2659 ( N_noxref_6_c_2823_n N_noxref_20_M81_noxref_g ) capacitor \
 c=0.0194981f //x=21.745 //y=5.155 //x2=21.27 //y2=6.02
cc_2660 ( N_noxref_6_M80_noxref_d N_noxref_20_M81_noxref_g ) capacitor \
 c=0.0194246f //x=20.905 //y=5.02 //x2=21.27 //y2=6.02
cc_2661 ( N_noxref_6_M13_noxref_d N_noxref_20_c_8638_n ) capacitor \
 c=0.00217566f //x=21.155 //y=0.915 //x2=21.08 //y2=0.915
cc_2662 ( N_noxref_6_M13_noxref_d N_noxref_20_c_8639_n ) capacitor \
 c=0.0034598f //x=21.155 //y=0.915 //x2=21.08 //y2=1.26
cc_2663 ( N_noxref_6_M13_noxref_d N_noxref_20_c_8640_n ) capacitor \
 c=0.00546784f //x=21.155 //y=0.915 //x2=21.08 //y2=1.57
cc_2664 ( N_noxref_6_M13_noxref_d N_noxref_20_c_8641_n ) capacitor \
 c=0.00241102f //x=21.155 //y=0.915 //x2=21.455 //y2=0.76
cc_2665 ( N_noxref_6_c_2754_n N_noxref_20_c_8642_n ) capacitor c=0.00371277f \
 //x=21.745 //y=1.665 //x2=21.455 //y2=1.415
cc_2666 ( N_noxref_6_M13_noxref_d N_noxref_20_c_8642_n ) capacitor \
 c=0.0138621f //x=21.155 //y=0.915 //x2=21.455 //y2=1.415
cc_2667 ( N_noxref_6_M13_noxref_d N_noxref_20_c_8644_n ) capacitor \
 c=0.00219619f //x=21.155 //y=0.915 //x2=21.61 //y2=0.915
cc_2668 ( N_noxref_6_c_2754_n N_noxref_20_c_8645_n ) capacitor c=0.00457401f \
 //x=21.745 //y=1.665 //x2=21.61 //y2=1.26
cc_2669 ( N_noxref_6_M13_noxref_d N_noxref_20_c_8645_n ) capacitor \
 c=0.00603828f //x=21.155 //y=0.915 //x2=21.61 //y2=1.26
cc_2670 ( N_noxref_6_c_2827_n N_noxref_20_c_8647_n ) capacitor c=0.00709342f \
 //x=21.83 //y=4.07 //x2=21.09 //y2=2.08
cc_2671 ( N_noxref_6_c_2827_n N_noxref_20_c_8648_n ) capacitor c=0.00283672f \
 //x=21.83 //y=4.07 //x2=21.09 //y2=1.915
cc_2672 ( N_noxref_6_M13_noxref_d N_noxref_20_c_8648_n ) capacitor \
 c=0.00661782f //x=21.155 //y=0.915 //x2=21.09 //y2=1.915
cc_2673 ( N_noxref_6_c_2823_n N_noxref_20_c_8650_n ) capacitor c=0.00201851f \
 //x=21.745 //y=5.155 //x2=21.09 //y2=4.7
cc_2674 ( N_noxref_6_c_2827_n N_noxref_20_c_8650_n ) capacitor c=0.013844f \
 //x=21.83 //y=4.07 //x2=21.09 //y2=4.7
cc_2675 ( N_noxref_6_c_3121_p N_noxref_20_c_8650_n ) capacitor c=0.00475601f \
 //x=21.05 //y=5.155 //x2=21.09 //y2=4.7
cc_2676 ( N_noxref_6_c_3161_p N_noxref_20_M15_noxref_d ) capacitor \
 c=0.00217566f //x=24.455 //y=0.905 //x2=24.53 //y2=0.905
cc_2677 ( N_noxref_6_c_3162_p N_noxref_20_M15_noxref_d ) capacitor \
 c=0.0034598f //x=24.455 //y=1.25 //x2=24.53 //y2=0.905
cc_2678 ( N_noxref_6_c_3163_p N_noxref_20_M15_noxref_d ) capacitor \
 c=0.0066953f //x=24.455 //y=1.56 //x2=24.53 //y2=0.905
cc_2679 ( N_noxref_6_c_3164_p N_noxref_20_M15_noxref_d ) capacitor \
 c=0.00241102f //x=24.83 //y=0.75 //x2=24.53 //y2=0.905
cc_2680 ( N_noxref_6_c_3069_p N_noxref_20_M15_noxref_d ) capacitor \
 c=0.0137169f //x=24.83 //y=1.405 //x2=24.53 //y2=0.905
cc_2681 ( N_noxref_6_c_3166_p N_noxref_20_M15_noxref_d ) capacitor \
 c=0.00132245f //x=24.985 //y=0.905 //x2=24.53 //y2=0.905
cc_2682 ( N_noxref_6_c_3131_p N_noxref_20_M15_noxref_d ) capacitor \
 c=0.00566463f //x=24.985 //y=1.25 //x2=24.53 //y2=0.905
cc_2683 ( N_noxref_6_c_3139_p N_noxref_20_M15_noxref_d ) capacitor \
 c=0.00660593f //x=24.42 //y=1.915 //x2=24.53 //y2=0.905
cc_2684 ( N_noxref_6_M83_noxref_g N_noxref_20_M82_noxref_d ) capacitor \
 c=0.0173476f //x=24.02 //y=6.02 //x2=23.655 //y2=5.02
cc_2685 ( N_noxref_6_M84_noxref_g N_noxref_20_M84_noxref_d ) capacitor \
 c=0.0173476f //x=24.46 //y=6.02 //x2=24.535 //y2=5.02
cc_2686 ( N_noxref_6_M85_noxref_g N_noxref_20_M84_noxref_d ) capacitor \
 c=0.0179769f //x=24.9 //y=6.02 //x2=24.535 //y2=5.02
cc_2687 ( N_noxref_6_c_2762_n N_noxref_23_c_9282_n ) capacitor c=0.0034165f \
 //x=0.81 //y=1.915 //x2=0.59 //y2=1.505
cc_2688 ( N_noxref_6_c_2748_n N_noxref_23_c_9266_n ) capacitor c=0.00179505f \
 //x=11.355 //y=4.07 //x2=1.475 //y2=1.59
cc_2689 ( N_noxref_6_c_2749_n N_noxref_23_c_9266_n ) capacitor c=0.00102628f \
 //x=1.225 //y=4.07 //x2=1.475 //y2=1.59
cc_2690 ( N_noxref_6_c_2750_n N_noxref_23_c_9266_n ) capacitor c=0.0122033f \
 //x=1.11 //y=2.08 //x2=1.475 //y2=1.59
cc_2691 ( N_noxref_6_c_2761_n N_noxref_23_c_9266_n ) capacitor c=0.00703864f \
 //x=0.81 //y=1.53 //x2=1.475 //y2=1.59
cc_2692 ( N_noxref_6_c_2762_n N_noxref_23_c_9266_n ) capacitor c=0.0259045f \
 //x=0.81 //y=1.915 //x2=1.475 //y2=1.59
cc_2693 ( N_noxref_6_c_2764_n N_noxref_23_c_9266_n ) capacitor c=0.00708583f \
 //x=1.185 //y=1.375 //x2=1.475 //y2=1.59
cc_2694 ( N_noxref_6_c_2767_n N_noxref_23_c_9266_n ) capacitor c=0.00698822f \
 //x=1.34 //y=1.22 //x2=1.475 //y2=1.59
cc_2695 ( N_noxref_6_c_2748_n N_noxref_23_c_9290_n ) capacitor c=0.0058169f \
 //x=11.355 //y=4.07 //x2=2.445 //y2=1.59
cc_2696 ( N_noxref_6_c_2748_n N_noxref_23_M0_noxref_s ) capacitor \
 c=0.00262629f //x=11.355 //y=4.07 //x2=0.455 //y2=0.375
cc_2697 ( N_noxref_6_c_2758_n N_noxref_23_M0_noxref_s ) capacitor c=0.0327271f \
 //x=0.81 //y=0.875 //x2=0.455 //y2=0.375
cc_2698 ( N_noxref_6_c_2761_n N_noxref_23_M0_noxref_s ) capacitor \
 c=7.99997e-19 //x=0.81 //y=1.53 //x2=0.455 //y2=0.375
cc_2699 ( N_noxref_6_c_2762_n N_noxref_23_M0_noxref_s ) capacitor \
 c=0.00122123f //x=0.81 //y=1.915 //x2=0.455 //y2=0.375
cc_2700 ( N_noxref_6_c_2765_n N_noxref_23_M0_noxref_s ) capacitor c=0.0121427f \
 //x=1.34 //y=0.875 //x2=0.455 //y2=0.375
cc_2701 ( N_noxref_6_c_2748_n N_noxref_24_c_9312_n ) capacitor c=0.0020922f \
 //x=11.355 //y=4.07 //x2=3.015 //y2=0.995
cc_2702 ( N_noxref_6_c_2748_n N_noxref_24_M2_noxref_s ) capacitor \
 c=0.00143334f //x=11.355 //y=4.07 //x2=2.965 //y2=0.375
cc_2703 ( N_noxref_6_c_2907_n N_noxref_27_c_9476_n ) capacitor c=0.00623646f \
 //x=11.505 //y=1.56 //x2=11.285 //y2=1.495
cc_2704 ( N_noxref_6_c_2912_n N_noxref_27_c_9476_n ) capacitor c=0.00173579f \
 //x=11.47 //y=2.08 //x2=11.285 //y2=1.495
cc_2705 ( N_noxref_6_c_2751_n N_noxref_27_c_9477_n ) capacitor c=0.00156605f \
 //x=11.47 //y=2.08 //x2=12.17 //y2=0.53
cc_2706 ( N_noxref_6_c_2902_n N_noxref_27_c_9477_n ) capacitor c=0.0188655f \
 //x=11.505 //y=0.905 //x2=12.17 //y2=0.53
cc_2707 ( N_noxref_6_c_2910_n N_noxref_27_c_9477_n ) capacitor c=0.00656458f \
 //x=12.035 //y=0.905 //x2=12.17 //y2=0.53
cc_2708 ( N_noxref_6_c_2912_n N_noxref_27_c_9477_n ) capacitor c=2.1838e-19 \
 //x=11.47 //y=2.08 //x2=12.17 //y2=0.53
cc_2709 ( N_noxref_6_c_2902_n N_noxref_27_M6_noxref_s ) capacitor \
 c=0.00623646f //x=11.505 //y=0.905 //x2=10.18 //y2=0.365
cc_2710 ( N_noxref_6_c_2910_n N_noxref_27_M6_noxref_s ) capacitor c=0.0143002f \
 //x=12.035 //y=0.905 //x2=10.18 //y2=0.365
cc_2711 ( N_noxref_6_c_2911_n N_noxref_27_M6_noxref_s ) capacitor \
 c=0.00290153f //x=12.035 //y=1.25 //x2=10.18 //y2=0.365
cc_2712 ( N_noxref_6_M10_noxref_d N_noxref_28_M8_noxref_s ) capacitor \
 c=0.00309936f //x=16.345 //y=0.915 //x2=13.405 //y2=0.375
cc_2713 ( N_noxref_6_c_2753_n N_noxref_29_c_9574_n ) capacitor c=0.00457167f \
 //x=16.935 //y=1.665 //x2=16.935 //y2=0.54
cc_2714 ( N_noxref_6_M10_noxref_d N_noxref_29_c_9574_n ) capacitor \
 c=0.0115903f //x=16.345 //y=0.915 //x2=16.935 //y2=0.54
cc_2715 ( N_noxref_6_c_3060_p N_noxref_29_c_9584_n ) capacitor c=0.0200405f \
 //x=16.62 //y=1.665 //x2=16.05 //y2=0.995
cc_2716 ( N_noxref_6_M10_noxref_d N_noxref_29_M9_noxref_d ) capacitor \
 c=5.27807e-19 //x=16.345 //y=0.915 //x2=14.81 //y2=0.91
cc_2717 ( N_noxref_6_c_2753_n N_noxref_29_M10_noxref_s ) capacitor \
 c=0.0196084f //x=16.935 //y=1.665 //x2=15.915 //y2=0.375
cc_2718 ( N_noxref_6_M10_noxref_d N_noxref_29_M10_noxref_s ) capacitor \
 c=0.0426368f //x=16.345 //y=0.915 //x2=15.915 //y2=0.375
cc_2719 ( N_noxref_6_c_2753_n N_noxref_30_c_9637_n ) capacitor c=3.84569e-19 \
 //x=16.935 //y=1.665 //x2=18.35 //y2=1.505
cc_2720 ( N_noxref_6_M10_noxref_d N_noxref_30_M11_noxref_s ) capacitor \
 c=2.55333e-19 //x=16.345 //y=0.915 //x2=18.215 //y2=0.375
cc_2721 ( N_noxref_6_M13_noxref_d N_noxref_30_M11_noxref_s ) capacitor \
 c=0.00309936f //x=21.155 //y=0.915 //x2=18.215 //y2=0.375
cc_2722 ( N_noxref_6_c_2754_n N_noxref_31_c_9679_n ) capacitor c=0.00457167f \
 //x=21.745 //y=1.665 //x2=21.745 //y2=0.54
cc_2723 ( N_noxref_6_M13_noxref_d N_noxref_31_c_9679_n ) capacitor \
 c=0.0115903f //x=21.155 //y=0.915 //x2=21.745 //y2=0.54
cc_2724 ( N_noxref_6_c_3064_p N_noxref_31_c_9689_n ) capacitor c=0.020048f \
 //x=21.43 //y=1.665 //x2=20.86 //y2=0.995
cc_2725 ( N_noxref_6_M13_noxref_d N_noxref_31_M12_noxref_d ) capacitor \
 c=5.27807e-19 //x=21.155 //y=0.915 //x2=19.62 //y2=0.91
cc_2726 ( N_noxref_6_c_2754_n N_noxref_31_M13_noxref_s ) capacitor \
 c=0.0196084f //x=21.745 //y=1.665 //x2=20.725 //y2=0.375
cc_2727 ( N_noxref_6_M13_noxref_d N_noxref_31_M13_noxref_s ) capacitor \
 c=0.0426444f //x=21.155 //y=0.915 //x2=20.725 //y2=0.375
cc_2728 ( N_noxref_6_c_2754_n N_noxref_32_c_9744_n ) capacitor c=3.04182e-19 \
 //x=21.745 //y=1.665 //x2=23.265 //y2=1.495
cc_2729 ( N_noxref_6_c_2772_n N_noxref_32_c_9744_n ) capacitor c=0.0034165f \
 //x=23.485 //y=1.915 //x2=23.265 //y2=1.495
cc_2730 ( N_noxref_6_c_2755_n N_noxref_32_c_9726_n ) capacitor c=0.011618f \
 //x=23.68 //y=2.08 //x2=24.15 //y2=1.58
cc_2731 ( N_noxref_6_c_2771_n N_noxref_32_c_9726_n ) capacitor c=0.00696403f \
 //x=23.485 //y=1.52 //x2=24.15 //y2=1.58
cc_2732 ( N_noxref_6_c_2772_n N_noxref_32_c_9726_n ) capacitor c=0.0174694f \
 //x=23.485 //y=1.915 //x2=24.15 //y2=1.58
cc_2733 ( N_noxref_6_c_2774_n N_noxref_32_c_9726_n ) capacitor c=0.00776811f \
 //x=23.86 //y=1.365 //x2=24.15 //y2=1.58
cc_2734 ( N_noxref_6_c_2777_n N_noxref_32_c_9726_n ) capacitor c=0.00339872f \
 //x=24.015 //y=1.21 //x2=24.15 //y2=1.58
cc_2735 ( N_noxref_6_c_2772_n N_noxref_32_c_9733_n ) capacitor c=6.71402e-19 \
 //x=23.485 //y=1.915 //x2=24.235 //y2=1.495
cc_2736 ( N_noxref_6_c_3163_p N_noxref_32_c_9733_n ) capacitor c=0.00623646f \
 //x=24.455 //y=1.56 //x2=24.235 //y2=1.495
cc_2737 ( N_noxref_6_c_3070_p N_noxref_32_c_9733_n ) capacitor c=0.00173579f \
 //x=24.42 //y=2.08 //x2=24.235 //y2=1.495
cc_2738 ( N_noxref_6_c_2756_n N_noxref_32_c_9734_n ) capacitor c=0.00156605f \
 //x=24.42 //y=2.08 //x2=25.12 //y2=0.53
cc_2739 ( N_noxref_6_c_3161_p N_noxref_32_c_9734_n ) capacitor c=0.0188655f \
 //x=24.455 //y=0.905 //x2=25.12 //y2=0.53
cc_2740 ( N_noxref_6_c_3166_p N_noxref_32_c_9734_n ) capacitor c=0.00656458f \
 //x=24.985 //y=0.905 //x2=25.12 //y2=0.53
cc_2741 ( N_noxref_6_c_3070_p N_noxref_32_c_9734_n ) capacitor c=2.1838e-19 \
 //x=24.42 //y=2.08 //x2=25.12 //y2=0.53
cc_2742 ( N_noxref_6_c_2768_n N_noxref_32_M14_noxref_s ) capacitor \
 c=0.0327502f //x=23.485 //y=0.865 //x2=23.13 //y2=0.365
cc_2743 ( N_noxref_6_c_2771_n N_noxref_32_M14_noxref_s ) capacitor \
 c=3.48408e-19 //x=23.485 //y=1.52 //x2=23.13 //y2=0.365
cc_2744 ( N_noxref_6_c_2775_n N_noxref_32_M14_noxref_s ) capacitor \
 c=0.0120759f //x=24.015 //y=0.865 //x2=23.13 //y2=0.365
cc_2745 ( N_noxref_6_c_3161_p N_noxref_32_M14_noxref_s ) capacitor \
 c=0.00623646f //x=24.455 //y=0.905 //x2=23.13 //y2=0.365
cc_2746 ( N_noxref_6_c_3166_p N_noxref_32_M14_noxref_s ) capacitor \
 c=0.0143002f //x=24.985 //y=0.905 //x2=23.13 //y2=0.365
cc_2747 ( N_noxref_6_c_3131_p N_noxref_32_M14_noxref_s ) capacitor \
 c=0.00290153f //x=24.985 //y=1.25 //x2=23.13 //y2=0.365
cc_2748 ( N_noxref_7_c_3290_p N_noxref_8_c_3527_n ) capacitor c=0.011463f \
 //x=36.515 //y=3.33 //x2=38.225 //y2=3.33
cc_2749 ( N_noxref_7_M99_noxref_g N_noxref_8_c_3496_n ) capacitor c=0.0169521f \
 //x=36.97 //y=6.02 //x2=37.545 //y2=5.2
cc_2750 ( N_noxref_7_c_3235_n N_noxref_8_c_3500_n ) capacitor c=0.00539951f \
 //x=36.63 //y=2.08 //x2=36.835 //y2=5.2
cc_2751 ( N_noxref_7_M98_noxref_g N_noxref_8_c_3500_n ) capacitor c=0.0177326f \
 //x=36.53 //y=6.02 //x2=36.835 //y2=5.2
cc_2752 ( N_noxref_7_c_3274_n N_noxref_8_c_3500_n ) capacitor c=0.00581252f \
 //x=36.63 //y=4.7 //x2=36.835 //y2=5.2
cc_2753 ( N_noxref_7_c_3262_n N_noxref_8_c_3481_n ) capacitor c=3.52729e-19 \
 //x=34.78 //y=3.33 //x2=38.11 //y2=3.33
cc_2754 ( N_noxref_7_c_3235_n N_noxref_8_c_3481_n ) capacitor c=0.00250675f \
 //x=36.63 //y=2.08 //x2=38.11 //y2=3.33
cc_2755 ( N_noxref_7_M99_noxref_g N_noxref_8_M98_noxref_d ) capacitor \
 c=0.0173476f //x=36.97 //y=6.02 //x2=36.605 //y2=5.02
cc_2756 ( N_noxref_7_c_3298_p N_noxref_9_c_3705_n ) capacitor c=0.146539f \
 //x=34.665 //y=3.33 //x2=31.705 //y2=3.7
cc_2757 ( N_noxref_7_c_3298_p N_noxref_9_c_3706_n ) capacitor c=0.0294746f \
 //x=34.665 //y=3.33 //x2=30.085 //y2=3.7
cc_2758 ( N_noxref_7_c_3233_n N_noxref_9_c_3706_n ) capacitor c=0.00687545f \
 //x=29.23 //y=2.08 //x2=30.085 //y2=3.7
cc_2759 ( N_noxref_7_c_3298_p N_noxref_9_c_3708_n ) capacitor c=0.238435f \
 //x=34.665 //y=3.33 //x2=44.655 //y2=3.7
cc_2760 ( N_noxref_7_c_3290_p N_noxref_9_c_3708_n ) capacitor c=0.175734f \
 //x=36.515 //y=3.33 //x2=44.655 //y2=3.7
cc_2761 ( N_noxref_7_c_3303_p N_noxref_9_c_3708_n ) capacitor c=0.0268386f \
 //x=34.895 //y=3.33 //x2=44.655 //y2=3.7
cc_2762 ( N_noxref_7_c_3262_n N_noxref_9_c_3708_n ) capacitor c=0.0206044f \
 //x=34.78 //y=3.33 //x2=44.655 //y2=3.7
cc_2763 ( N_noxref_7_c_3235_n N_noxref_9_c_3708_n ) capacitor c=0.0205831f \
 //x=36.63 //y=2.08 //x2=44.655 //y2=3.7
cc_2764 ( N_noxref_7_c_3298_p N_noxref_9_c_3713_n ) capacitor c=0.0266966f \
 //x=34.665 //y=3.33 //x2=31.935 //y2=3.7
cc_2765 ( N_noxref_7_M90_noxref_g N_noxref_9_c_3663_n ) capacitor c=0.01736f \
 //x=28.97 //y=6.02 //x2=29.105 //y2=5.155
cc_2766 ( N_noxref_7_c_3252_n N_noxref_9_c_3667_n ) capacitor c=3.10026e-19 \
 //x=32.325 //y=5.155 //x2=29.885 //y2=5.155
cc_2767 ( N_noxref_7_M91_noxref_g N_noxref_9_c_3667_n ) capacitor c=0.0194981f \
 //x=29.41 //y=6.02 //x2=29.885 //y2=5.155
cc_2768 ( N_noxref_7_c_3310_p N_noxref_9_c_3667_n ) capacitor c=0.00201851f \
 //x=29.23 //y=4.7 //x2=29.885 //y2=5.155
cc_2769 ( N_noxref_7_c_3311_p N_noxref_9_c_3633_n ) capacitor c=0.00371277f \
 //x=29.595 //y=1.415 //x2=29.885 //y2=1.665
cc_2770 ( N_noxref_7_c_3312_p N_noxref_9_c_3633_n ) capacitor c=0.00457401f \
 //x=29.75 //y=1.26 //x2=29.885 //y2=1.665
cc_2771 ( N_noxref_7_c_3298_p N_noxref_9_c_3671_n ) capacitor c=0.0206036f \
 //x=34.665 //y=3.33 //x2=29.97 //y2=3.7
cc_2772 ( N_noxref_7_c_3314_p N_noxref_9_c_3671_n ) capacitor c=0.00179385f \
 //x=29.345 //y=3.33 //x2=29.97 //y2=3.7
cc_2773 ( N_noxref_7_c_3233_n N_noxref_9_c_3671_n ) capacitor c=0.0760319f \
 //x=29.23 //y=2.08 //x2=29.97 //y2=3.7
cc_2774 ( N_noxref_7_c_3316_p N_noxref_9_c_3671_n ) capacitor c=0.00731987f \
 //x=29.23 //y=2.08 //x2=29.97 //y2=3.7
cc_2775 ( N_noxref_7_c_3317_p N_noxref_9_c_3671_n ) capacitor c=0.00283672f \
 //x=29.23 //y=1.915 //x2=29.97 //y2=3.7
cc_2776 ( N_noxref_7_c_3310_p N_noxref_9_c_3671_n ) capacitor c=0.013693f \
 //x=29.23 //y=4.7 //x2=29.97 //y2=3.7
cc_2777 ( N_noxref_7_c_3298_p N_noxref_9_c_3634_n ) capacitor c=0.021615f \
 //x=34.665 //y=3.33 //x2=31.82 //y2=2.08
cc_2778 ( N_noxref_7_c_3233_n N_noxref_9_c_3634_n ) capacitor c=8.46099e-19 \
 //x=29.23 //y=2.08 //x2=31.82 //y2=2.08
cc_2779 ( N_noxref_7_c_3233_n N_noxref_9_c_3728_n ) capacitor c=0.0166016f \
 //x=29.23 //y=2.08 //x2=29.19 //y2=5.155
cc_2780 ( N_noxref_7_c_3310_p N_noxref_9_c_3728_n ) capacitor c=0.00475601f \
 //x=29.23 //y=4.7 //x2=29.19 //y2=5.155
cc_2781 ( N_noxref_7_c_3252_n N_noxref_9_M92_noxref_g ) capacitor c=0.0213876f \
 //x=32.325 //y=5.155 //x2=32.02 //y2=6.02
cc_2782 ( N_noxref_7_c_3248_n N_noxref_9_M93_noxref_g ) capacitor c=0.0168349f \
 //x=33.035 //y=5.155 //x2=32.46 //y2=6.02
cc_2783 ( N_noxref_7_M92_noxref_d N_noxref_9_M93_noxref_g ) capacitor \
 c=0.0180032f //x=32.095 //y=5.02 //x2=32.46 //y2=6.02
cc_2784 ( N_noxref_7_c_3252_n N_noxref_9_c_3733_n ) capacitor c=0.00428486f \
 //x=32.325 //y=5.155 //x2=32.385 //y2=4.79
cc_2785 ( N_noxref_7_c_3327_p N_noxref_9_M18_noxref_d ) capacitor \
 c=0.00217566f //x=29.22 //y=0.915 //x2=29.295 //y2=0.915
cc_2786 ( N_noxref_7_c_3328_p N_noxref_9_M18_noxref_d ) capacitor c=0.0034598f \
 //x=29.22 //y=1.26 //x2=29.295 //y2=0.915
cc_2787 ( N_noxref_7_c_3329_p N_noxref_9_M18_noxref_d ) capacitor \
 c=0.00546784f //x=29.22 //y=1.57 //x2=29.295 //y2=0.915
cc_2788 ( N_noxref_7_c_3330_p N_noxref_9_M18_noxref_d ) capacitor \
 c=0.00241102f //x=29.595 //y=0.76 //x2=29.295 //y2=0.915
cc_2789 ( N_noxref_7_c_3311_p N_noxref_9_M18_noxref_d ) capacitor c=0.0138621f \
 //x=29.595 //y=1.415 //x2=29.295 //y2=0.915
cc_2790 ( N_noxref_7_c_3332_p N_noxref_9_M18_noxref_d ) capacitor \
 c=0.00219619f //x=29.75 //y=0.915 //x2=29.295 //y2=0.915
cc_2791 ( N_noxref_7_c_3312_p N_noxref_9_M18_noxref_d ) capacitor \
 c=0.00603828f //x=29.75 //y=1.26 //x2=29.295 //y2=0.915
cc_2792 ( N_noxref_7_c_3317_p N_noxref_9_M18_noxref_d ) capacitor \
 c=0.00661782f //x=29.23 //y=1.915 //x2=29.295 //y2=0.915
cc_2793 ( N_noxref_7_M90_noxref_g N_noxref_9_M90_noxref_d ) capacitor \
 c=0.0180032f //x=28.97 //y=6.02 //x2=29.045 //y2=5.02
cc_2794 ( N_noxref_7_M91_noxref_g N_noxref_9_M90_noxref_d ) capacitor \
 c=0.0194246f //x=29.41 //y=6.02 //x2=29.045 //y2=5.02
cc_2795 ( N_noxref_7_c_3298_p N_noxref_11_c_4075_n ) capacitor c=0.0558554f \
 //x=34.665 //y=3.33 //x2=37.255 //y2=4.07
cc_2796 ( N_noxref_7_c_3314_p N_noxref_11_c_4075_n ) capacitor c=0.0135672f \
 //x=29.345 //y=3.33 //x2=37.255 //y2=4.07
cc_2797 ( N_noxref_7_c_3290_p N_noxref_11_c_4075_n ) capacitor c=0.010979f \
 //x=36.515 //y=3.33 //x2=37.255 //y2=4.07
cc_2798 ( N_noxref_7_c_3303_p N_noxref_11_c_4075_n ) capacitor c=4.80262e-19 \
 //x=34.895 //y=3.33 //x2=37.255 //y2=4.07
cc_2799 ( N_noxref_7_c_3233_n N_noxref_11_c_4075_n ) capacitor c=0.0206302f \
 //x=29.23 //y=2.08 //x2=37.255 //y2=4.07
cc_2800 ( N_noxref_7_c_3262_n N_noxref_11_c_4075_n ) capacitor c=0.0181982f \
 //x=34.78 //y=3.33 //x2=37.255 //y2=4.07
cc_2801 ( N_noxref_7_c_3235_n N_noxref_11_c_4075_n ) capacitor c=0.0184765f \
 //x=36.63 //y=2.08 //x2=37.255 //y2=4.07
cc_2802 ( N_noxref_7_c_3235_n N_noxref_11_c_4144_n ) capacitor c=0.00179385f \
 //x=36.63 //y=2.08 //x2=37.485 //y2=4.07
cc_2803 ( N_noxref_7_c_3233_n N_noxref_11_c_4058_n ) capacitor c=0.00133538f \
 //x=29.23 //y=2.08 //x2=27.01 //y2=2.08
cc_2804 ( N_noxref_7_c_3235_n N_noxref_11_c_4146_n ) capacitor c=0.00400249f \
 //x=36.63 //y=2.08 //x2=37.37 //y2=4.535
cc_2805 ( N_noxref_7_c_3274_n N_noxref_11_c_4146_n ) capacitor c=0.00417994f \
 //x=36.63 //y=4.7 //x2=37.37 //y2=4.535
cc_2806 ( N_noxref_7_c_3290_p N_noxref_11_c_4059_n ) capacitor c=0.00318578f \
 //x=36.515 //y=3.33 //x2=37.37 //y2=2.08
cc_2807 ( N_noxref_7_c_3262_n N_noxref_11_c_4059_n ) capacitor c=8.48165e-19 \
 //x=34.78 //y=3.33 //x2=37.37 //y2=2.08
cc_2808 ( N_noxref_7_c_3235_n N_noxref_11_c_4059_n ) capacitor c=0.0721686f \
 //x=36.63 //y=2.08 //x2=37.37 //y2=2.08
cc_2809 ( N_noxref_7_c_3240_n N_noxref_11_c_4059_n ) capacitor c=0.00284029f \
 //x=36.435 //y=1.915 //x2=37.37 //y2=2.08
cc_2810 ( N_noxref_7_M98_noxref_g N_noxref_11_M100_noxref_g ) capacitor \
 c=0.0104611f //x=36.53 //y=6.02 //x2=37.41 //y2=6.02
cc_2811 ( N_noxref_7_M99_noxref_g N_noxref_11_M100_noxref_g ) capacitor \
 c=0.106811f //x=36.97 //y=6.02 //x2=37.41 //y2=6.02
cc_2812 ( N_noxref_7_M99_noxref_g N_noxref_11_M101_noxref_g ) capacitor \
 c=0.0100341f //x=36.97 //y=6.02 //x2=37.85 //y2=6.02
cc_2813 ( N_noxref_7_c_3236_n N_noxref_11_c_4155_n ) capacitor c=4.86506e-19 \
 //x=36.435 //y=0.865 //x2=37.405 //y2=0.905
cc_2814 ( N_noxref_7_c_3238_n N_noxref_11_c_4155_n ) capacitor c=0.00152104f \
 //x=36.435 //y=1.21 //x2=37.405 //y2=0.905
cc_2815 ( N_noxref_7_c_3243_n N_noxref_11_c_4155_n ) capacitor c=0.0151475f \
 //x=36.965 //y=0.865 //x2=37.405 //y2=0.905
cc_2816 ( N_noxref_7_c_3239_n N_noxref_11_c_4158_n ) capacitor c=0.00109982f \
 //x=36.435 //y=1.52 //x2=37.405 //y2=1.25
cc_2817 ( N_noxref_7_c_3245_n N_noxref_11_c_4158_n ) capacitor c=0.0111064f \
 //x=36.965 //y=1.21 //x2=37.405 //y2=1.25
cc_2818 ( N_noxref_7_c_3239_n N_noxref_11_c_4160_n ) capacitor c=9.57794e-19 \
 //x=36.435 //y=1.52 //x2=37.405 //y2=1.56
cc_2819 ( N_noxref_7_c_3240_n N_noxref_11_c_4160_n ) capacitor c=0.00662747f \
 //x=36.435 //y=1.915 //x2=37.405 //y2=1.56
cc_2820 ( N_noxref_7_c_3245_n N_noxref_11_c_4160_n ) capacitor c=0.00862358f \
 //x=36.965 //y=1.21 //x2=37.405 //y2=1.56
cc_2821 ( N_noxref_7_c_3243_n N_noxref_11_c_4163_n ) capacitor c=0.00124821f \
 //x=36.965 //y=0.865 //x2=37.935 //y2=0.905
cc_2822 ( N_noxref_7_c_3245_n N_noxref_11_c_4164_n ) capacitor c=0.00200715f \
 //x=36.965 //y=1.21 //x2=37.935 //y2=1.25
cc_2823 ( N_noxref_7_c_3235_n N_noxref_11_c_4165_n ) capacitor c=0.00282278f \
 //x=36.63 //y=2.08 //x2=37.37 //y2=2.08
cc_2824 ( N_noxref_7_c_3240_n N_noxref_11_c_4165_n ) capacitor c=0.0172771f \
 //x=36.435 //y=1.915 //x2=37.37 //y2=2.08
cc_2825 ( N_noxref_7_c_3235_n N_noxref_11_c_4167_n ) capacitor c=0.00344981f \
 //x=36.63 //y=2.08 //x2=37.4 //y2=4.7
cc_2826 ( N_noxref_7_c_3274_n N_noxref_11_c_4167_n ) capacitor c=0.0293367f \
 //x=36.63 //y=4.7 //x2=37.4 //y2=4.7
cc_2827 ( N_noxref_7_c_3298_p N_D_c_4434_n ) capacitor c=0.0262386f //x=34.665 \
 //y=3.33 //x2=32.815 //y2=2.59
cc_2828 ( N_noxref_7_c_3314_p N_D_c_4434_n ) capacitor c=9.8111e-19 //x=29.345 \
 //y=3.33 //x2=32.815 //y2=2.59
cc_2829 ( N_noxref_7_c_3233_n N_D_c_4434_n ) capacitor c=0.0179628f //x=29.23 \
 //y=2.08 //x2=32.815 //y2=2.59
cc_2830 ( N_noxref_7_c_3298_p N_D_c_4442_n ) capacitor c=0.0153535f //x=34.665 \
 //y=3.33 //x2=58.715 //y2=2.59
cc_2831 ( N_noxref_7_c_3290_p N_D_c_4442_n ) capacitor c=0.0125403f //x=36.515 \
 //y=3.33 //x2=58.715 //y2=2.59
cc_2832 ( N_noxref_7_c_3303_p N_D_c_4442_n ) capacitor c=5.76706e-19 \
 //x=34.895 //y=3.33 //x2=58.715 //y2=2.59
cc_2833 ( N_noxref_7_c_3262_n N_D_c_4442_n ) capacitor c=0.0165903f //x=34.78 \
 //y=3.33 //x2=58.715 //y2=2.59
cc_2834 ( N_noxref_7_c_3235_n N_D_c_4442_n ) capacitor c=0.0177872f //x=36.63 \
 //y=2.08 //x2=58.715 //y2=2.59
cc_2835 ( N_noxref_7_c_3298_p N_D_c_4538_n ) capacitor c=6.65036e-19 \
 //x=34.665 //y=3.33 //x2=33.045 //y2=2.59
cc_2836 ( N_noxref_7_c_3298_p N_D_c_4449_n ) capacitor c=0.0190562f //x=34.665 \
 //y=3.33 //x2=32.93 //y2=2.08
cc_2837 ( N_noxref_7_c_3248_n N_D_c_4449_n ) capacitor c=0.0146f //x=33.035 \
 //y=5.155 //x2=32.93 //y2=2.08
cc_2838 ( N_noxref_7_c_3262_n N_D_c_4449_n ) capacitor c=0.0022276f //x=34.78 \
 //y=3.33 //x2=32.93 //y2=2.08
cc_2839 ( N_noxref_7_c_3248_n N_D_M94_noxref_g ) capacitor c=0.0165266f \
 //x=33.035 //y=5.155 //x2=32.9 //y2=6.02
cc_2840 ( N_noxref_7_M94_noxref_d N_D_M94_noxref_g ) capacitor c=0.0180032f \
 //x=32.975 //y=5.02 //x2=32.9 //y2=6.02
cc_2841 ( N_noxref_7_c_3254_n N_D_M95_noxref_g ) capacitor c=0.01736f \
 //x=33.915 //y=5.155 //x2=33.34 //y2=6.02
cc_2842 ( N_noxref_7_M94_noxref_d N_D_M95_noxref_g ) capacitor c=0.0180032f \
 //x=32.975 //y=5.02 //x2=33.34 //y2=6.02
cc_2843 ( N_noxref_7_c_3385_p N_D_c_4546_n ) capacitor c=0.00426767f //x=33.12 \
 //y=5.155 //x2=33.265 //y2=4.79
cc_2844 ( N_noxref_7_c_3248_n N_D_c_4547_n ) capacitor c=0.00322054f \
 //x=33.035 //y=5.155 //x2=32.93 //y2=4.7
cc_2845 ( N_noxref_7_c_3298_p N_CLK_c_4844_n ) capacitor c=0.00360213f \
 //x=34.665 //y=3.33 //x2=40.955 //y2=4.44
cc_2846 ( N_noxref_7_c_3314_p N_CLK_c_4844_n ) capacitor c=4.49102e-19 \
 //x=29.345 //y=3.33 //x2=40.955 //y2=4.44
cc_2847 ( N_noxref_7_c_3233_n N_CLK_c_4844_n ) capacitor c=0.0200057f \
 //x=29.23 //y=2.08 //x2=40.955 //y2=4.44
cc_2848 ( N_noxref_7_c_3248_n N_CLK_c_4844_n ) capacitor c=0.032141f \
 //x=33.035 //y=5.155 //x2=40.955 //y2=4.44
cc_2849 ( N_noxref_7_c_3252_n N_CLK_c_4844_n ) capacitor c=0.0230136f \
 //x=32.325 //y=5.155 //x2=40.955 //y2=4.44
cc_2850 ( N_noxref_7_c_3258_n N_CLK_c_4844_n ) capacitor c=0.0183122f \
 //x=34.695 //y=5.155 //x2=40.955 //y2=4.44
cc_2851 ( N_noxref_7_c_3262_n N_CLK_c_4844_n ) capacitor c=0.0210274f \
 //x=34.78 //y=3.33 //x2=40.955 //y2=4.44
cc_2852 ( N_noxref_7_c_3235_n N_CLK_c_4844_n ) capacitor c=0.0198304f \
 //x=36.63 //y=2.08 //x2=40.955 //y2=4.44
cc_2853 ( N_noxref_7_c_3310_p N_CLK_c_4844_n ) capacitor c=0.0111881f \
 //x=29.23 //y=4.7 //x2=40.955 //y2=4.44
cc_2854 ( N_noxref_7_c_3274_n N_CLK_c_4844_n ) capacitor c=0.0107057f \
 //x=36.63 //y=4.7 //x2=40.955 //y2=4.44
cc_2855 ( N_noxref_7_c_3233_n N_CLK_c_4861_n ) capacitor c=0.00153281f \
 //x=29.23 //y=2.08 //x2=28.235 //y2=4.44
cc_2856 ( N_noxref_7_c_3314_p N_CLK_c_4804_n ) capacitor c=0.00526349f \
 //x=29.345 //y=3.33 //x2=28.12 //y2=2.08
cc_2857 ( N_noxref_7_c_3233_n N_CLK_c_4804_n ) capacitor c=0.0443839f \
 //x=29.23 //y=2.08 //x2=28.12 //y2=2.08
cc_2858 ( N_noxref_7_c_3316_p N_CLK_c_4804_n ) capacitor c=0.00201097f \
 //x=29.23 //y=2.08 //x2=28.12 //y2=2.08
cc_2859 ( N_noxref_7_c_3310_p N_CLK_c_4804_n ) capacitor c=0.00218014f \
 //x=29.23 //y=4.7 //x2=28.12 //y2=2.08
cc_2860 ( N_noxref_7_M90_noxref_g N_CLK_M88_noxref_g ) capacitor c=0.0101598f \
 //x=28.97 //y=6.02 //x2=28.09 //y2=6.02
cc_2861 ( N_noxref_7_M90_noxref_g N_CLK_M89_noxref_g ) capacitor c=0.0602553f \
 //x=28.97 //y=6.02 //x2=28.53 //y2=6.02
cc_2862 ( N_noxref_7_M91_noxref_g N_CLK_M89_noxref_g ) capacitor c=0.0101598f \
 //x=29.41 //y=6.02 //x2=28.53 //y2=6.02
cc_2863 ( N_noxref_7_c_3327_p N_CLK_c_5094_n ) capacitor c=0.00456962f \
 //x=29.22 //y=0.915 //x2=28.21 //y2=0.91
cc_2864 ( N_noxref_7_c_3328_p N_CLK_c_5095_n ) capacitor c=0.00438372f \
 //x=29.22 //y=1.26 //x2=28.21 //y2=1.22
cc_2865 ( N_noxref_7_c_3329_p N_CLK_c_5096_n ) capacitor c=0.00438372f \
 //x=29.22 //y=1.57 //x2=28.21 //y2=1.45
cc_2866 ( N_noxref_7_c_3233_n N_CLK_c_5097_n ) capacitor c=0.00205895f \
 //x=29.23 //y=2.08 //x2=28.21 //y2=1.915
cc_2867 ( N_noxref_7_c_3316_p N_CLK_c_5097_n ) capacitor c=0.00828003f \
 //x=29.23 //y=2.08 //x2=28.21 //y2=1.915
cc_2868 ( N_noxref_7_c_3317_p N_CLK_c_5097_n ) capacitor c=0.00438372f \
 //x=29.23 //y=1.915 //x2=28.21 //y2=1.915
cc_2869 ( N_noxref_7_c_3310_p N_CLK_c_5100_n ) capacitor c=0.0611812f \
 //x=29.23 //y=4.7 //x2=28.455 //y2=4.79
cc_2870 ( N_noxref_7_c_3233_n N_CLK_c_5101_n ) capacitor c=0.00142741f \
 //x=29.23 //y=2.08 //x2=28.12 //y2=4.7
cc_2871 ( N_noxref_7_c_3310_p N_CLK_c_5101_n ) capacitor c=0.00487508f \
 //x=29.23 //y=4.7 //x2=28.12 //y2=4.7
cc_2872 ( N_noxref_7_c_3233_n N_RN_c_5861_n ) capacitor c=0.0186201f //x=29.23 \
 //y=2.08 //x2=33.925 //y2=2.22
cc_2873 ( N_noxref_7_c_3311_p N_RN_c_5861_n ) capacitor c=3.13485e-19 \
 //x=29.595 //y=1.415 //x2=33.925 //y2=2.22
cc_2874 ( N_noxref_7_c_3316_p N_RN_c_5861_n ) capacitor c=0.00584491f \
 //x=29.23 //y=2.08 //x2=33.925 //y2=2.22
cc_2875 ( N_noxref_7_c_3417_p N_RN_c_5873_n ) capacitor c=0.016327f //x=34.38 \
 //y=1.665 //x2=42.065 //y2=2.22
cc_2876 ( N_noxref_7_c_3262_n N_RN_c_5873_n ) capacitor c=0.0197307f //x=34.78 \
 //y=3.33 //x2=42.065 //y2=2.22
cc_2877 ( N_noxref_7_c_3235_n N_RN_c_5873_n ) capacitor c=0.0185012f //x=36.63 \
 //y=2.08 //x2=42.065 //y2=2.22
cc_2878 ( N_noxref_7_c_3240_n N_RN_c_5873_n ) capacitor c=0.00894156f \
 //x=36.435 //y=1.915 //x2=42.065 //y2=2.22
cc_2879 ( N_noxref_7_c_3262_n N_RN_c_5881_n ) capacitor c=0.00184436f \
 //x=34.78 //y=3.33 //x2=34.155 //y2=2.22
cc_2880 ( N_noxref_7_c_3298_p N_RN_c_5916_n ) capacitor c=0.0180187f \
 //x=34.665 //y=3.33 //x2=34.04 //y2=2.08
cc_2881 ( N_noxref_7_c_3303_p N_RN_c_5916_n ) capacitor c=0.00131333f \
 //x=34.895 //y=3.33 //x2=34.04 //y2=2.08
cc_2882 ( N_noxref_7_c_3262_n N_RN_c_5916_n ) capacitor c=0.075348f //x=34.78 \
 //y=3.33 //x2=34.04 //y2=2.08
cc_2883 ( N_noxref_7_c_3235_n N_RN_c_5916_n ) capacitor c=6.23409e-19 \
 //x=36.63 //y=2.08 //x2=34.04 //y2=2.08
cc_2884 ( N_noxref_7_c_3426_p N_RN_c_5916_n ) capacitor c=0.0171303f //x=34 \
 //y=5.155 //x2=34.04 //y2=2.08
cc_2885 ( N_noxref_7_c_3254_n N_RN_M96_noxref_g ) capacitor c=0.01736f \
 //x=33.915 //y=5.155 //x2=33.78 //y2=6.02
cc_2886 ( N_noxref_7_M96_noxref_d N_RN_M96_noxref_g ) capacitor c=0.0180032f \
 //x=33.855 //y=5.02 //x2=33.78 //y2=6.02
cc_2887 ( N_noxref_7_c_3258_n N_RN_M97_noxref_g ) capacitor c=0.0194981f \
 //x=34.695 //y=5.155 //x2=34.22 //y2=6.02
cc_2888 ( N_noxref_7_M96_noxref_d N_RN_M97_noxref_g ) capacitor c=0.0194246f \
 //x=33.855 //y=5.02 //x2=34.22 //y2=6.02
cc_2889 ( N_noxref_7_M21_noxref_d N_RN_c_6109_n ) capacitor c=0.00217566f \
 //x=34.105 //y=0.915 //x2=34.03 //y2=0.915
cc_2890 ( N_noxref_7_M21_noxref_d N_RN_c_6110_n ) capacitor c=0.0034598f \
 //x=34.105 //y=0.915 //x2=34.03 //y2=1.26
cc_2891 ( N_noxref_7_M21_noxref_d N_RN_c_6111_n ) capacitor c=0.00546784f \
 //x=34.105 //y=0.915 //x2=34.03 //y2=1.57
cc_2892 ( N_noxref_7_M21_noxref_d N_RN_c_6112_n ) capacitor c=0.00241102f \
 //x=34.105 //y=0.915 //x2=34.405 //y2=0.76
cc_2893 ( N_noxref_7_c_3234_n N_RN_c_6113_n ) capacitor c=0.00371277f \
 //x=34.695 //y=1.665 //x2=34.405 //y2=1.415
cc_2894 ( N_noxref_7_M21_noxref_d N_RN_c_6113_n ) capacitor c=0.0138621f \
 //x=34.105 //y=0.915 //x2=34.405 //y2=1.415
cc_2895 ( N_noxref_7_M21_noxref_d N_RN_c_6115_n ) capacitor c=0.00219619f \
 //x=34.105 //y=0.915 //x2=34.56 //y2=0.915
cc_2896 ( N_noxref_7_c_3234_n N_RN_c_6116_n ) capacitor c=0.00457401f \
 //x=34.695 //y=1.665 //x2=34.56 //y2=1.26
cc_2897 ( N_noxref_7_M21_noxref_d N_RN_c_6116_n ) capacitor c=0.00603828f \
 //x=34.105 //y=0.915 //x2=34.56 //y2=1.26
cc_2898 ( N_noxref_7_c_3262_n N_RN_c_6118_n ) capacitor c=0.00709342f \
 //x=34.78 //y=3.33 //x2=34.04 //y2=2.08
cc_2899 ( N_noxref_7_c_3262_n N_RN_c_6119_n ) capacitor c=0.00283672f \
 //x=34.78 //y=3.33 //x2=34.04 //y2=1.915
cc_2900 ( N_noxref_7_M21_noxref_d N_RN_c_6119_n ) capacitor c=0.00661782f \
 //x=34.105 //y=0.915 //x2=34.04 //y2=1.915
cc_2901 ( N_noxref_7_c_3258_n N_RN_c_6121_n ) capacitor c=0.00201851f \
 //x=34.695 //y=5.155 //x2=34.04 //y2=4.7
cc_2902 ( N_noxref_7_c_3262_n N_RN_c_6121_n ) capacitor c=0.013844f //x=34.78 \
 //y=3.33 //x2=34.04 //y2=4.7
cc_2903 ( N_noxref_7_c_3426_p N_RN_c_6121_n ) capacitor c=0.00475601f //x=34 \
 //y=5.155 //x2=34.04 //y2=4.7
cc_2904 ( N_noxref_7_c_3298_p N_noxref_20_c_8516_n ) capacitor c=0.466581f \
 //x=34.665 //y=3.33 //x2=83.505 //y2=2.96
cc_2905 ( N_noxref_7_c_3314_p N_noxref_20_c_8516_n ) capacitor c=0.0291389f \
 //x=29.345 //y=3.33 //x2=83.505 //y2=2.96
cc_2906 ( N_noxref_7_c_3290_p N_noxref_20_c_8516_n ) capacitor c=0.173514f \
 //x=36.515 //y=3.33 //x2=83.505 //y2=2.96
cc_2907 ( N_noxref_7_c_3303_p N_noxref_20_c_8516_n ) capacitor c=0.0266688f \
 //x=34.895 //y=3.33 //x2=83.505 //y2=2.96
cc_2908 ( N_noxref_7_c_3233_n N_noxref_20_c_8516_n ) capacitor c=0.0198264f \
 //x=29.23 //y=2.08 //x2=83.505 //y2=2.96
cc_2909 ( N_noxref_7_c_3262_n N_noxref_20_c_8516_n ) capacitor c=0.0206002f \
 //x=34.78 //y=3.33 //x2=83.505 //y2=2.96
cc_2910 ( N_noxref_7_c_3235_n N_noxref_20_c_8516_n ) capacitor c=0.0205758f \
 //x=36.63 //y=2.08 //x2=83.505 //y2=2.96
cc_2911 ( N_noxref_7_c_3233_n N_noxref_34_c_9831_n ) capacitor c=0.00204385f \
 //x=29.23 //y=2.08 //x2=29.885 //y2=0.54
cc_2912 ( N_noxref_7_c_3327_p N_noxref_34_c_9831_n ) capacitor c=0.0194423f \
 //x=29.22 //y=0.915 //x2=29.885 //y2=0.54
cc_2913 ( N_noxref_7_c_3332_p N_noxref_34_c_9831_n ) capacitor c=0.00656458f \
 //x=29.75 //y=0.915 //x2=29.885 //y2=0.54
cc_2914 ( N_noxref_7_c_3316_p N_noxref_34_c_9831_n ) capacitor c=2.20712e-19 \
 //x=29.23 //y=2.08 //x2=29.885 //y2=0.54
cc_2915 ( N_noxref_7_c_3328_p N_noxref_34_c_9843_n ) capacitor c=0.00538829f \
 //x=29.22 //y=1.26 //x2=29 //y2=0.995
cc_2916 ( N_noxref_7_c_3327_p N_noxref_34_M18_noxref_s ) capacitor \
 c=0.00538829f //x=29.22 //y=0.915 //x2=28.865 //y2=0.375
cc_2917 ( N_noxref_7_c_3329_p N_noxref_34_M18_noxref_s ) capacitor \
 c=0.00538829f //x=29.22 //y=1.57 //x2=28.865 //y2=0.375
cc_2918 ( N_noxref_7_c_3332_p N_noxref_34_M18_noxref_s ) capacitor \
 c=0.0143002f //x=29.75 //y=0.915 //x2=28.865 //y2=0.375
cc_2919 ( N_noxref_7_c_3312_p N_noxref_34_M18_noxref_s ) capacitor \
 c=0.00290153f //x=29.75 //y=1.26 //x2=28.865 //y2=0.375
cc_2920 ( N_noxref_7_M21_noxref_d N_noxref_35_M19_noxref_s ) capacitor \
 c=0.00309936f //x=34.105 //y=0.915 //x2=31.165 //y2=0.375
cc_2921 ( N_noxref_7_c_3234_n N_noxref_36_c_9932_n ) capacitor c=0.00457167f \
 //x=34.695 //y=1.665 //x2=34.695 //y2=0.54
cc_2922 ( N_noxref_7_M21_noxref_d N_noxref_36_c_9932_n ) capacitor \
 c=0.0115903f //x=34.105 //y=0.915 //x2=34.695 //y2=0.54
cc_2923 ( N_noxref_7_c_3417_p N_noxref_36_c_9942_n ) capacitor c=0.020048f \
 //x=34.38 //y=1.665 //x2=33.81 //y2=0.995
cc_2924 ( N_noxref_7_M21_noxref_d N_noxref_36_M20_noxref_d ) capacitor \
 c=5.27807e-19 //x=34.105 //y=0.915 //x2=32.57 //y2=0.91
cc_2925 ( N_noxref_7_c_3234_n N_noxref_36_M21_noxref_s ) capacitor \
 c=0.0196084f //x=34.695 //y=1.665 //x2=33.675 //y2=0.375
cc_2926 ( N_noxref_7_M21_noxref_d N_noxref_36_M21_noxref_s ) capacitor \
 c=0.0426444f //x=34.105 //y=0.915 //x2=33.675 //y2=0.375
cc_2927 ( N_noxref_7_c_3234_n N_noxref_37_c_9998_n ) capacitor c=3.04182e-19 \
 //x=34.695 //y=1.665 //x2=36.215 //y2=1.495
cc_2928 ( N_noxref_7_c_3240_n N_noxref_37_c_9998_n ) capacitor c=0.0034165f \
 //x=36.435 //y=1.915 //x2=36.215 //y2=1.495
cc_2929 ( N_noxref_7_c_3235_n N_noxref_37_c_9980_n ) capacitor c=0.0111916f \
 //x=36.63 //y=2.08 //x2=37.1 //y2=1.58
cc_2930 ( N_noxref_7_c_3239_n N_noxref_37_c_9980_n ) capacitor c=0.00696403f \
 //x=36.435 //y=1.52 //x2=37.1 //y2=1.58
cc_2931 ( N_noxref_7_c_3240_n N_noxref_37_c_9980_n ) capacitor c=0.0174694f \
 //x=36.435 //y=1.915 //x2=37.1 //y2=1.58
cc_2932 ( N_noxref_7_c_3242_n N_noxref_37_c_9980_n ) capacitor c=0.00776811f \
 //x=36.81 //y=1.365 //x2=37.1 //y2=1.58
cc_2933 ( N_noxref_7_c_3245_n N_noxref_37_c_9980_n ) capacitor c=0.00339872f \
 //x=36.965 //y=1.21 //x2=37.1 //y2=1.58
cc_2934 ( N_noxref_7_c_3240_n N_noxref_37_c_9987_n ) capacitor c=6.71402e-19 \
 //x=36.435 //y=1.915 //x2=37.185 //y2=1.495
cc_2935 ( N_noxref_7_c_3236_n N_noxref_37_M22_noxref_s ) capacitor \
 c=0.0327502f //x=36.435 //y=0.865 //x2=36.08 //y2=0.365
cc_2936 ( N_noxref_7_c_3239_n N_noxref_37_M22_noxref_s ) capacitor \
 c=3.48408e-19 //x=36.435 //y=1.52 //x2=36.08 //y2=0.365
cc_2937 ( N_noxref_7_c_3243_n N_noxref_37_M22_noxref_s ) capacitor \
 c=0.0120759f //x=36.965 //y=0.865 //x2=36.08 //y2=0.365
cc_2938 ( N_noxref_8_c_3535_p N_noxref_9_c_3708_n ) capacitor c=0.176049f \
 //x=39.845 //y=3.33 //x2=44.655 //y2=3.7
cc_2939 ( N_noxref_8_c_3527_n N_noxref_9_c_3708_n ) capacitor c=0.0293967f \
 //x=38.225 //y=3.33 //x2=44.655 //y2=3.7
cc_2940 ( N_noxref_8_c_3481_n N_noxref_9_c_3708_n ) capacitor c=0.0206034f \
 //x=38.11 //y=3.33 //x2=44.655 //y2=3.7
cc_2941 ( N_noxref_8_c_3482_n N_noxref_9_c_3708_n ) capacitor c=0.0216236f \
 //x=39.96 //y=2.08 //x2=44.655 //y2=3.7
cc_2942 ( N_noxref_8_c_3535_p N_noxref_11_c_4078_n ) capacitor c=0.0107156f \
 //x=39.845 //y=3.33 //x2=42.805 //y2=4.07
cc_2943 ( N_noxref_8_c_3527_n N_noxref_11_c_4078_n ) capacitor c=8.88358e-19 \
 //x=38.225 //y=3.33 //x2=42.805 //y2=4.07
cc_2944 ( N_noxref_8_c_3481_n N_noxref_11_c_4078_n ) capacitor c=0.0181936f \
 //x=38.11 //y=3.33 //x2=42.805 //y2=4.07
cc_2945 ( N_noxref_8_c_3482_n N_noxref_11_c_4078_n ) capacitor c=0.019517f \
 //x=39.96 //y=2.08 //x2=42.805 //y2=4.07
cc_2946 ( N_noxref_8_c_3481_n N_noxref_11_c_4144_n ) capacitor c=0.00179385f \
 //x=38.11 //y=3.33 //x2=37.485 //y2=4.07
cc_2947 ( N_noxref_8_c_3496_n N_noxref_11_c_4146_n ) capacitor c=0.0127164f \
 //x=37.545 //y=5.2 //x2=37.37 //y2=4.535
cc_2948 ( N_noxref_8_c_3481_n N_noxref_11_c_4146_n ) capacitor c=0.0101115f \
 //x=38.11 //y=3.33 //x2=37.37 //y2=4.535
cc_2949 ( N_noxref_8_c_3527_n N_noxref_11_c_4059_n ) capacitor c=0.00329059f \
 //x=38.225 //y=3.33 //x2=37.37 //y2=2.08
cc_2950 ( N_noxref_8_c_3481_n N_noxref_11_c_4059_n ) capacitor c=0.0671907f \
 //x=38.11 //y=3.33 //x2=37.37 //y2=2.08
cc_2951 ( N_noxref_8_c_3482_n N_noxref_11_c_4059_n ) capacitor c=8.48165e-19 \
 //x=39.96 //y=2.08 //x2=37.37 //y2=2.08
cc_2952 ( N_noxref_8_M103_noxref_g N_noxref_11_c_4087_n ) capacitor \
 c=0.0168349f //x=40.6 //y=6.02 //x2=41.175 //y2=5.155
cc_2953 ( N_noxref_8_c_3481_n N_noxref_11_c_4091_n ) capacitor c=2.97874e-19 \
 //x=38.11 //y=3.33 //x2=40.465 //y2=5.155
cc_2954 ( N_noxref_8_M102_noxref_g N_noxref_11_c_4091_n ) capacitor \
 c=0.0213876f //x=40.16 //y=6.02 //x2=40.465 //y2=5.155
cc_2955 ( N_noxref_8_c_3552_p N_noxref_11_c_4091_n ) capacitor c=0.00428486f \
 //x=40.525 //y=4.79 //x2=40.465 //y2=5.155
cc_2956 ( N_noxref_8_c_3496_n N_noxref_11_M100_noxref_g ) capacitor \
 c=0.0166421f //x=37.545 //y=5.2 //x2=37.41 //y2=6.02
cc_2957 ( N_noxref_8_M100_noxref_d N_noxref_11_M100_noxref_g ) capacitor \
 c=0.0173476f //x=37.485 //y=5.02 //x2=37.41 //y2=6.02
cc_2958 ( N_noxref_8_c_3502_n N_noxref_11_M101_noxref_g ) capacitor \
 c=0.018922f //x=38.025 //y=5.2 //x2=37.85 //y2=6.02
cc_2959 ( N_noxref_8_M100_noxref_d N_noxref_11_M101_noxref_g ) capacitor \
 c=0.0179769f //x=37.485 //y=5.02 //x2=37.85 //y2=6.02
cc_2960 ( N_noxref_8_M23_noxref_d N_noxref_11_c_4155_n ) capacitor \
 c=0.00217566f //x=37.48 //y=0.905 //x2=37.405 //y2=0.905
cc_2961 ( N_noxref_8_M23_noxref_d N_noxref_11_c_4158_n ) capacitor \
 c=0.0034598f //x=37.48 //y=0.905 //x2=37.405 //y2=1.25
cc_2962 ( N_noxref_8_M23_noxref_d N_noxref_11_c_4160_n ) capacitor \
 c=0.0066953f //x=37.48 //y=0.905 //x2=37.405 //y2=1.56
cc_2963 ( N_noxref_8_c_3481_n N_noxref_11_c_4190_n ) capacitor c=0.0142673f \
 //x=38.11 //y=3.33 //x2=37.775 //y2=4.79
cc_2964 ( N_noxref_8_c_3561_p N_noxref_11_c_4190_n ) capacitor c=0.00407665f \
 //x=37.63 //y=5.2 //x2=37.775 //y2=4.79
cc_2965 ( N_noxref_8_M23_noxref_d N_noxref_11_c_4192_n ) capacitor \
 c=0.00241102f //x=37.48 //y=0.905 //x2=37.78 //y2=0.75
cc_2966 ( N_noxref_8_c_3480_n N_noxref_11_c_4193_n ) capacitor c=0.00371277f \
 //x=38.025 //y=1.655 //x2=37.78 //y2=1.405
cc_2967 ( N_noxref_8_M23_noxref_d N_noxref_11_c_4193_n ) capacitor \
 c=0.0137169f //x=37.48 //y=0.905 //x2=37.78 //y2=1.405
cc_2968 ( N_noxref_8_M23_noxref_d N_noxref_11_c_4163_n ) capacitor \
 c=0.00132245f //x=37.48 //y=0.905 //x2=37.935 //y2=0.905
cc_2969 ( N_noxref_8_c_3480_n N_noxref_11_c_4164_n ) capacitor c=0.00457401f \
 //x=38.025 //y=1.655 //x2=37.935 //y2=1.25
cc_2970 ( N_noxref_8_M23_noxref_d N_noxref_11_c_4164_n ) capacitor \
 c=0.00566463f //x=37.48 //y=0.905 //x2=37.935 //y2=1.25
cc_2971 ( N_noxref_8_c_3481_n N_noxref_11_c_4165_n ) capacitor c=0.00731987f \
 //x=38.11 //y=3.33 //x2=37.37 //y2=2.08
cc_2972 ( N_noxref_8_c_3481_n N_noxref_11_c_4199_n ) capacitor c=0.00306024f \
 //x=38.11 //y=3.33 //x2=37.37 //y2=1.915
cc_2973 ( N_noxref_8_M23_noxref_d N_noxref_11_c_4199_n ) capacitor \
 c=0.00660593f //x=37.48 //y=0.905 //x2=37.37 //y2=1.915
cc_2974 ( N_noxref_8_c_3496_n N_noxref_11_c_4167_n ) capacitor c=0.00346527f \
 //x=37.545 //y=5.2 //x2=37.4 //y2=4.7
cc_2975 ( N_noxref_8_c_3481_n N_noxref_11_c_4167_n ) capacitor c=0.00517969f \
 //x=38.11 //y=3.33 //x2=37.4 //y2=4.7
cc_2976 ( N_noxref_8_M103_noxref_g N_noxref_11_M102_noxref_d ) capacitor \
 c=0.0180032f //x=40.6 //y=6.02 //x2=40.235 //y2=5.02
cc_2977 ( N_noxref_8_c_3535_p N_D_c_4442_n ) capacitor c=0.0119007f //x=39.845 \
 //y=3.33 //x2=58.715 //y2=2.59
cc_2978 ( N_noxref_8_c_3527_n N_D_c_4442_n ) capacitor c=8.92472e-19 \
 //x=38.225 //y=3.33 //x2=58.715 //y2=2.59
cc_2979 ( N_noxref_8_c_3481_n N_D_c_4442_n ) capacitor c=0.0165961f //x=38.11 \
 //y=3.33 //x2=58.715 //y2=2.59
cc_2980 ( N_noxref_8_c_3482_n N_D_c_4442_n ) capacitor c=0.0188253f //x=39.96 \
 //y=2.08 //x2=58.715 //y2=2.59
cc_2981 ( N_noxref_8_c_3496_n N_CLK_c_4844_n ) capacitor c=0.0185297f \
 //x=37.545 //y=5.2 //x2=40.955 //y2=4.44
cc_2982 ( N_noxref_8_c_3500_n N_CLK_c_4844_n ) capacitor c=0.018142f \
 //x=36.835 //y=5.2 //x2=40.955 //y2=4.44
cc_2983 ( N_noxref_8_c_3481_n N_CLK_c_4844_n ) capacitor c=0.0208321f \
 //x=38.11 //y=3.33 //x2=40.955 //y2=4.44
cc_2984 ( N_noxref_8_c_3482_n N_CLK_c_4844_n ) capacitor c=0.0208709f \
 //x=39.96 //y=2.08 //x2=40.955 //y2=4.44
cc_2985 ( N_noxref_8_c_3514_n N_CLK_c_4844_n ) capacitor c=0.0166984f \
 //x=40.235 //y=4.79 //x2=40.955 //y2=4.44
cc_2986 ( N_noxref_8_c_3482_n N_CLK_c_4879_n ) capacitor c=0.00153281f \
 //x=39.96 //y=2.08 //x2=41.185 //y2=4.44
cc_2987 ( N_noxref_8_c_3535_p N_CLK_c_4805_n ) capacitor c=0.00520283f \
 //x=39.845 //y=3.33 //x2=41.07 //y2=2.08
cc_2988 ( N_noxref_8_c_3481_n N_CLK_c_4805_n ) capacitor c=5.10318e-19 \
 //x=38.11 //y=3.33 //x2=41.07 //y2=2.08
cc_2989 ( N_noxref_8_c_3482_n N_CLK_c_4805_n ) capacitor c=0.0422272f \
 //x=39.96 //y=2.08 //x2=41.07 //y2=2.08
cc_2990 ( N_noxref_8_c_3487_n N_CLK_c_4805_n ) capacitor c=0.00210802f \
 //x=39.66 //y=1.915 //x2=41.07 //y2=2.08
cc_2991 ( N_noxref_8_c_3552_p N_CLK_c_4805_n ) capacitor c=0.00147352f \
 //x=40.525 //y=4.79 //x2=41.07 //y2=2.08
cc_2992 ( N_noxref_8_c_3514_n N_CLK_c_4805_n ) capacitor c=0.00141297f \
 //x=40.235 //y=4.79 //x2=41.07 //y2=2.08
cc_2993 ( N_noxref_8_M102_noxref_g N_CLK_M104_noxref_g ) capacitor \
 c=0.0105869f //x=40.16 //y=6.02 //x2=41.04 //y2=6.02
cc_2994 ( N_noxref_8_M103_noxref_g N_CLK_M104_noxref_g ) capacitor c=0.10632f \
 //x=40.6 //y=6.02 //x2=41.04 //y2=6.02
cc_2995 ( N_noxref_8_M103_noxref_g N_CLK_M105_noxref_g ) capacitor \
 c=0.0101598f //x=40.6 //y=6.02 //x2=41.48 //y2=6.02
cc_2996 ( N_noxref_8_c_3483_n N_CLK_c_5118_n ) capacitor c=5.72482e-19 \
 //x=39.66 //y=0.875 //x2=40.635 //y2=0.91
cc_2997 ( N_noxref_8_c_3485_n N_CLK_c_5118_n ) capacitor c=0.00149976f \
 //x=39.66 //y=1.22 //x2=40.635 //y2=0.91
cc_2998 ( N_noxref_8_c_3490_n N_CLK_c_5118_n ) capacitor c=0.0160123f \
 //x=40.19 //y=0.875 //x2=40.635 //y2=0.91
cc_2999 ( N_noxref_8_c_3486_n N_CLK_c_5121_n ) capacitor c=0.00111227f \
 //x=39.66 //y=1.53 //x2=40.635 //y2=1.22
cc_3000 ( N_noxref_8_c_3492_n N_CLK_c_5121_n ) capacitor c=0.0124075f \
 //x=40.19 //y=1.22 //x2=40.635 //y2=1.22
cc_3001 ( N_noxref_8_c_3490_n N_CLK_c_5123_n ) capacitor c=0.00103227f \
 //x=40.19 //y=0.875 //x2=41.16 //y2=0.91
cc_3002 ( N_noxref_8_c_3492_n N_CLK_c_5124_n ) capacitor c=0.0010154f \
 //x=40.19 //y=1.22 //x2=41.16 //y2=1.22
cc_3003 ( N_noxref_8_c_3492_n N_CLK_c_5125_n ) capacitor c=9.23422e-19 \
 //x=40.19 //y=1.22 //x2=41.16 //y2=1.45
cc_3004 ( N_noxref_8_c_3482_n N_CLK_c_5126_n ) capacitor c=0.00203769f \
 //x=39.96 //y=2.08 //x2=41.16 //y2=1.915
cc_3005 ( N_noxref_8_c_3487_n N_CLK_c_5126_n ) capacitor c=0.00834532f \
 //x=39.66 //y=1.915 //x2=41.16 //y2=1.915
cc_3006 ( N_noxref_8_c_3482_n N_CLK_c_5128_n ) capacitor c=0.00183762f \
 //x=39.96 //y=2.08 //x2=41.07 //y2=4.7
cc_3007 ( N_noxref_8_c_3552_p N_CLK_c_5128_n ) capacitor c=0.0168581f \
 //x=40.525 //y=4.79 //x2=41.07 //y2=4.7
cc_3008 ( N_noxref_8_c_3514_n N_CLK_c_5128_n ) capacitor c=0.00484466f \
 //x=40.235 //y=4.79 //x2=41.07 //y2=4.7
cc_3009 ( N_noxref_8_c_3606_p N_RN_c_5873_n ) capacitor c=0.0146822f \
 //x=37.755 //y=1.655 //x2=42.065 //y2=2.22
cc_3010 ( N_noxref_8_c_3481_n N_RN_c_5873_n ) capacitor c=0.0199049f //x=38.11 \
 //y=3.33 //x2=42.065 //y2=2.22
cc_3011 ( N_noxref_8_c_3482_n N_RN_c_5873_n ) capacitor c=0.0192695f //x=39.96 \
 //y=2.08 //x2=42.065 //y2=2.22
cc_3012 ( N_noxref_8_c_3487_n N_RN_c_5873_n ) capacitor c=0.011987f //x=39.66 \
 //y=1.915 //x2=42.065 //y2=2.22
cc_3013 ( N_noxref_8_c_3482_n N_RN_c_5917_n ) capacitor c=0.00107158f \
 //x=39.96 //y=2.08 //x2=42.18 //y2=2.08
cc_3014 ( N_noxref_8_c_3535_p N_noxref_20_c_8516_n ) capacitor c=0.173984f \
 //x=39.845 //y=3.33 //x2=83.505 //y2=2.96
cc_3015 ( N_noxref_8_c_3527_n N_noxref_20_c_8516_n ) capacitor c=0.0292689f \
 //x=38.225 //y=3.33 //x2=83.505 //y2=2.96
cc_3016 ( N_noxref_8_c_3481_n N_noxref_20_c_8516_n ) capacitor c=0.0206014f \
 //x=38.11 //y=3.33 //x2=83.505 //y2=2.96
cc_3017 ( N_noxref_8_c_3482_n N_noxref_20_c_8516_n ) capacitor c=0.0216162f \
 //x=39.96 //y=2.08 //x2=83.505 //y2=2.96
cc_3018 ( N_noxref_8_c_3606_p N_noxref_37_c_9998_n ) capacitor c=3.15806e-19 \
 //x=37.755 //y=1.655 //x2=36.215 //y2=1.495
cc_3019 ( N_noxref_8_c_3606_p N_noxref_37_c_9987_n ) capacitor c=0.020324f \
 //x=37.755 //y=1.655 //x2=37.185 //y2=1.495
cc_3020 ( N_noxref_8_c_3480_n N_noxref_37_c_9988_n ) capacitor c=0.00457164f \
 //x=38.025 //y=1.655 //x2=38.07 //y2=0.53
cc_3021 ( N_noxref_8_M23_noxref_d N_noxref_37_c_9988_n ) capacitor \
 c=0.0115831f //x=37.48 //y=0.905 //x2=38.07 //y2=0.53
cc_3022 ( N_noxref_8_c_3480_n N_noxref_37_M22_noxref_s ) capacitor c=0.013435f \
 //x=38.025 //y=1.655 //x2=36.08 //y2=0.365
cc_3023 ( N_noxref_8_M23_noxref_d N_noxref_37_M22_noxref_s ) capacitor \
 c=0.0439476f //x=37.48 //y=0.905 //x2=36.08 //y2=0.365
cc_3024 ( N_noxref_8_c_3480_n N_noxref_38_c_10046_n ) capacitor c=4.08644e-19 \
 //x=38.025 //y=1.655 //x2=39.44 //y2=1.505
cc_3025 ( N_noxref_8_c_3487_n N_noxref_38_c_10046_n ) capacitor c=0.0034165f \
 //x=39.66 //y=1.915 //x2=39.44 //y2=1.505
cc_3026 ( N_noxref_8_c_3482_n N_noxref_38_c_10031_n ) capacitor c=0.0115578f \
 //x=39.96 //y=2.08 //x2=40.325 //y2=1.59
cc_3027 ( N_noxref_8_c_3486_n N_noxref_38_c_10031_n ) capacitor c=0.00697148f \
 //x=39.66 //y=1.53 //x2=40.325 //y2=1.59
cc_3028 ( N_noxref_8_c_3487_n N_noxref_38_c_10031_n ) capacitor c=0.0204849f \
 //x=39.66 //y=1.915 //x2=40.325 //y2=1.59
cc_3029 ( N_noxref_8_c_3489_n N_noxref_38_c_10031_n ) capacitor c=0.00610316f \
 //x=40.035 //y=1.375 //x2=40.325 //y2=1.59
cc_3030 ( N_noxref_8_c_3492_n N_noxref_38_c_10031_n ) capacitor c=0.00698822f \
 //x=40.19 //y=1.22 //x2=40.325 //y2=1.59
cc_3031 ( N_noxref_8_c_3483_n N_noxref_38_M24_noxref_s ) capacitor \
 c=0.0327271f //x=39.66 //y=0.875 //x2=39.305 //y2=0.375
cc_3032 ( N_noxref_8_c_3486_n N_noxref_38_M24_noxref_s ) capacitor \
 c=7.99997e-19 //x=39.66 //y=1.53 //x2=39.305 //y2=0.375
cc_3033 ( N_noxref_8_c_3487_n N_noxref_38_M24_noxref_s ) capacitor \
 c=0.00122123f //x=39.66 //y=1.915 //x2=39.305 //y2=0.375
cc_3034 ( N_noxref_8_c_3490_n N_noxref_38_M24_noxref_s ) capacitor \
 c=0.0121427f //x=40.19 //y=0.875 //x2=39.305 //y2=0.375
cc_3035 ( N_noxref_8_M23_noxref_d N_noxref_38_M24_noxref_s ) capacitor \
 c=2.53688e-19 //x=37.48 //y=0.905 //x2=39.305 //y2=0.375
cc_3036 ( N_noxref_9_c_3708_n N_noxref_10_c_3946_n ) capacitor c=0.00564994f \
 //x=44.655 //y=3.7 //x2=47.845 //y2=3.7
cc_3037 ( N_noxref_9_M109_noxref_g N_noxref_10_c_3908_n ) capacitor \
 c=0.0168349f //x=45.41 //y=6.02 //x2=45.985 //y2=5.155
cc_3038 ( N_noxref_9_M108_noxref_g N_noxref_10_c_3912_n ) capacitor \
 c=0.0213876f //x=44.97 //y=6.02 //x2=45.275 //y2=5.155
cc_3039 ( N_noxref_9_c_3751_p N_noxref_10_c_3912_n ) capacitor c=0.00428486f \
 //x=45.335 //y=4.79 //x2=45.275 //y2=5.155
cc_3040 ( N_noxref_9_M109_noxref_g N_noxref_10_M108_noxref_d ) capacitor \
 c=0.0180032f //x=45.41 //y=6.02 //x2=45.045 //y2=5.02
cc_3041 ( N_noxref_9_c_3705_n N_noxref_11_c_4075_n ) capacitor c=0.147447f \
 //x=31.705 //y=3.7 //x2=37.255 //y2=4.07
cc_3042 ( N_noxref_9_c_3706_n N_noxref_11_c_4075_n ) capacitor c=0.0294294f \
 //x=30.085 //y=3.7 //x2=37.255 //y2=4.07
cc_3043 ( N_noxref_9_c_3708_n N_noxref_11_c_4075_n ) capacitor c=0.467539f \
 //x=44.655 //y=3.7 //x2=37.255 //y2=4.07
cc_3044 ( N_noxref_9_c_3713_n N_noxref_11_c_4075_n ) capacitor c=0.0264476f \
 //x=31.935 //y=3.7 //x2=37.255 //y2=4.07
cc_3045 ( N_noxref_9_c_3671_n N_noxref_11_c_4075_n ) capacitor c=0.0200328f \
 //x=29.97 //y=3.7 //x2=37.255 //y2=4.07
cc_3046 ( N_noxref_9_c_3634_n N_noxref_11_c_4075_n ) capacitor c=0.0213516f \
 //x=31.82 //y=2.08 //x2=37.255 //y2=4.07
cc_3047 ( N_noxref_9_c_3708_n N_noxref_11_c_4078_n ) capacitor c=0.468066f \
 //x=44.655 //y=3.7 //x2=42.805 //y2=4.07
cc_3048 ( N_noxref_9_c_3708_n N_noxref_11_c_4144_n ) capacitor c=0.0267832f \
 //x=44.655 //y=3.7 //x2=37.485 //y2=4.07
cc_3049 ( N_noxref_9_c_3708_n N_noxref_11_c_4079_n ) capacitor c=0.176507f \
 //x=44.655 //y=3.7 //x2=50.205 //y2=4.07
cc_3050 ( N_noxref_9_c_3635_n N_noxref_11_c_4079_n ) capacitor c=0.0213324f \
 //x=44.77 //y=2.08 //x2=50.205 //y2=4.07
cc_3051 ( N_noxref_9_c_3708_n N_noxref_11_c_4081_n ) capacitor c=0.0268461f \
 //x=44.655 //y=3.7 //x2=43.035 //y2=4.07
cc_3052 ( N_noxref_9_c_3635_n N_noxref_11_c_4081_n ) capacitor c=3.50683e-19 \
 //x=44.77 //y=2.08 //x2=43.035 //y2=4.07
cc_3053 ( N_noxref_9_c_3708_n N_noxref_11_c_4059_n ) capacitor c=0.0211371f \
 //x=44.655 //y=3.7 //x2=37.37 //y2=2.08
cc_3054 ( N_noxref_9_c_3708_n N_noxref_11_c_4101_n ) capacitor c=0.0236196f \
 //x=44.655 //y=3.7 //x2=42.92 //y2=4.07
cc_3055 ( N_noxref_9_c_3635_n N_noxref_11_c_4101_n ) capacitor c=0.0123451f \
 //x=44.77 //y=2.08 //x2=42.92 //y2=4.07
cc_3056 ( N_noxref_9_c_3661_n N_noxref_11_M86_noxref_g ) capacitor \
 c=0.0213876f //x=27.515 //y=5.155 //x2=27.21 //y2=6.02
cc_3057 ( N_noxref_9_c_3657_n N_noxref_11_M87_noxref_g ) capacitor \
 c=0.0168349f //x=28.225 //y=5.155 //x2=27.65 //y2=6.02
cc_3058 ( N_noxref_9_M86_noxref_d N_noxref_11_M87_noxref_g ) capacitor \
 c=0.0180032f //x=27.285 //y=5.02 //x2=27.65 //y2=6.02
cc_3059 ( N_noxref_9_c_3661_n N_noxref_11_c_4222_n ) capacitor c=0.00428486f \
 //x=27.515 //y=5.155 //x2=27.575 //y2=4.79
cc_3060 ( N_noxref_9_c_3671_n N_D_c_4434_n ) capacitor c=0.0165903f //x=29.97 \
 //y=3.7 //x2=32.815 //y2=2.59
cc_3061 ( N_noxref_9_c_3634_n N_D_c_4434_n ) capacitor c=0.0188253f //x=31.82 \
 //y=2.08 //x2=32.815 //y2=2.59
cc_3062 ( N_noxref_9_c_3708_n N_D_c_4442_n ) capacitor c=0.0324441f //x=44.655 \
 //y=3.7 //x2=58.715 //y2=2.59
cc_3063 ( N_noxref_9_c_3635_n N_D_c_4442_n ) capacitor c=0.0188253f //x=44.77 \
 //y=2.08 //x2=58.715 //y2=2.59
cc_3064 ( N_noxref_9_c_3634_n N_D_c_4538_n ) capacitor c=0.00128547f //x=31.82 \
 //y=2.08 //x2=33.045 //y2=2.59
cc_3065 ( N_noxref_9_c_3708_n N_D_c_4449_n ) capacitor c=0.0190398f //x=44.655 \
 //y=3.7 //x2=32.93 //y2=2.08
cc_3066 ( N_noxref_9_c_3713_n N_D_c_4449_n ) capacitor c=9.95819e-19 \
 //x=31.935 //y=3.7 //x2=32.93 //y2=2.08
cc_3067 ( N_noxref_9_c_3671_n N_D_c_4449_n ) capacitor c=3.3533e-19 //x=29.97 \
 //y=3.7 //x2=32.93 //y2=2.08
cc_3068 ( N_noxref_9_c_3634_n N_D_c_4449_n ) capacitor c=0.0413373f //x=31.82 \
 //y=2.08 //x2=32.93 //y2=2.08
cc_3069 ( N_noxref_9_c_3640_n N_D_c_4449_n ) capacitor c=0.00210802f //x=31.52 \
 //y=1.915 //x2=32.93 //y2=2.08
cc_3070 ( N_noxref_9_c_3733_n N_D_c_4449_n ) capacitor c=0.00147352f \
 //x=32.385 //y=4.79 //x2=32.93 //y2=2.08
cc_3071 ( N_noxref_9_c_3686_n N_D_c_4449_n ) capacitor c=0.00142741f \
 //x=32.095 //y=4.79 //x2=32.93 //y2=2.08
cc_3072 ( N_noxref_9_M92_noxref_g N_D_M94_noxref_g ) capacitor c=0.0105869f \
 //x=32.02 //y=6.02 //x2=32.9 //y2=6.02
cc_3073 ( N_noxref_9_M93_noxref_g N_D_M94_noxref_g ) capacitor c=0.10632f \
 //x=32.46 //y=6.02 //x2=32.9 //y2=6.02
cc_3074 ( N_noxref_9_M93_noxref_g N_D_M95_noxref_g ) capacitor c=0.0101598f \
 //x=32.46 //y=6.02 //x2=33.34 //y2=6.02
cc_3075 ( N_noxref_9_c_3636_n N_D_c_4567_n ) capacitor c=5.72482e-19 //x=31.52 \
 //y=0.875 //x2=32.495 //y2=0.91
cc_3076 ( N_noxref_9_c_3638_n N_D_c_4567_n ) capacitor c=0.00149976f //x=31.52 \
 //y=1.22 //x2=32.495 //y2=0.91
cc_3077 ( N_noxref_9_c_3643_n N_D_c_4567_n ) capacitor c=0.0160123f //x=32.05 \
 //y=0.875 //x2=32.495 //y2=0.91
cc_3078 ( N_noxref_9_c_3639_n N_D_c_4570_n ) capacitor c=0.00111227f //x=31.52 \
 //y=1.53 //x2=32.495 //y2=1.22
cc_3079 ( N_noxref_9_c_3645_n N_D_c_4570_n ) capacitor c=0.0124075f //x=32.05 \
 //y=1.22 //x2=32.495 //y2=1.22
cc_3080 ( N_noxref_9_c_3643_n N_D_c_4572_n ) capacitor c=0.00103227f //x=32.05 \
 //y=0.875 //x2=33.02 //y2=0.91
cc_3081 ( N_noxref_9_c_3645_n N_D_c_4573_n ) capacitor c=0.0010154f //x=32.05 \
 //y=1.22 //x2=33.02 //y2=1.22
cc_3082 ( N_noxref_9_c_3645_n N_D_c_4574_n ) capacitor c=9.23422e-19 //x=32.05 \
 //y=1.22 //x2=33.02 //y2=1.45
cc_3083 ( N_noxref_9_c_3634_n N_D_c_4575_n ) capacitor c=0.00203769f //x=31.82 \
 //y=2.08 //x2=33.02 //y2=1.915
cc_3084 ( N_noxref_9_c_3640_n N_D_c_4575_n ) capacitor c=0.00834532f //x=31.52 \
 //y=1.915 //x2=33.02 //y2=1.915
cc_3085 ( N_noxref_9_c_3634_n N_D_c_4547_n ) capacitor c=0.00183762f //x=31.82 \
 //y=2.08 //x2=32.93 //y2=4.7
cc_3086 ( N_noxref_9_c_3733_n N_D_c_4547_n ) capacitor c=0.0168581f //x=32.385 \
 //y=4.79 //x2=32.93 //y2=4.7
cc_3087 ( N_noxref_9_c_3686_n N_D_c_4547_n ) capacitor c=0.00484466f \
 //x=32.095 //y=4.79 //x2=32.93 //y2=4.7
cc_3088 ( N_noxref_9_c_3661_n N_CLK_c_4826_n ) capacitor c=0.0219114f \
 //x=27.515 //y=5.155 //x2=28.005 //y2=4.44
cc_3089 ( N_noxref_9_c_3705_n N_CLK_c_4844_n ) capacitor c=0.00910993f \
 //x=31.705 //y=3.7 //x2=40.955 //y2=4.44
cc_3090 ( N_noxref_9_c_3706_n N_CLK_c_4844_n ) capacitor c=7.95009e-19 \
 //x=30.085 //y=3.7 //x2=40.955 //y2=4.44
cc_3091 ( N_noxref_9_c_3708_n N_CLK_c_4844_n ) capacitor c=0.0658043f \
 //x=44.655 //y=3.7 //x2=40.955 //y2=4.44
cc_3092 ( N_noxref_9_c_3713_n N_CLK_c_4844_n ) capacitor c=6.59178e-19 \
 //x=31.935 //y=3.7 //x2=40.955 //y2=4.44
cc_3093 ( N_noxref_9_c_3667_n N_CLK_c_4844_n ) capacitor c=0.0183122f \
 //x=29.885 //y=5.155 //x2=40.955 //y2=4.44
cc_3094 ( N_noxref_9_c_3671_n N_CLK_c_4844_n ) capacitor c=0.0210274f \
 //x=29.97 //y=3.7 //x2=40.955 //y2=4.44
cc_3095 ( N_noxref_9_c_3634_n N_CLK_c_4844_n ) capacitor c=0.0208709f \
 //x=31.82 //y=2.08 //x2=40.955 //y2=4.44
cc_3096 ( N_noxref_9_c_3808_p N_CLK_c_4844_n ) capacitor c=0.0311227f \
 //x=28.31 //y=5.155 //x2=40.955 //y2=4.44
cc_3097 ( N_noxref_9_c_3686_n N_CLK_c_4844_n ) capacitor c=0.0166984f \
 //x=32.095 //y=4.79 //x2=40.955 //y2=4.44
cc_3098 ( N_noxref_9_c_3657_n N_CLK_c_4861_n ) capacitor c=0.00241768f \
 //x=28.225 //y=5.155 //x2=28.235 //y2=4.44
cc_3099 ( N_noxref_9_c_3708_n N_CLK_c_4862_n ) capacitor c=0.0254092f \
 //x=44.655 //y=3.7 //x2=53.905 //y2=4.44
cc_3100 ( N_noxref_9_c_3635_n N_CLK_c_4862_n ) capacitor c=0.0208709f \
 //x=44.77 //y=2.08 //x2=53.905 //y2=4.44
cc_3101 ( N_noxref_9_c_3688_n N_CLK_c_4862_n ) capacitor c=0.0166984f \
 //x=45.045 //y=4.79 //x2=53.905 //y2=4.44
cc_3102 ( N_noxref_9_c_3708_n N_CLK_c_4879_n ) capacitor c=6.6036e-19 \
 //x=44.655 //y=3.7 //x2=41.185 //y2=4.44
cc_3103 ( N_noxref_9_c_3657_n N_CLK_c_4804_n ) capacitor c=0.0143918f \
 //x=28.225 //y=5.155 //x2=28.12 //y2=2.08
cc_3104 ( N_noxref_9_c_3671_n N_CLK_c_4804_n ) capacitor c=0.00264025f \
 //x=29.97 //y=3.7 //x2=28.12 //y2=2.08
cc_3105 ( N_noxref_9_c_3708_n N_CLK_c_4805_n ) capacitor c=0.0213788f \
 //x=44.655 //y=3.7 //x2=41.07 //y2=2.08
cc_3106 ( N_noxref_9_c_3657_n N_CLK_M88_noxref_g ) capacitor c=0.016514f \
 //x=28.225 //y=5.155 //x2=28.09 //y2=6.02
cc_3107 ( N_noxref_9_M88_noxref_d N_CLK_M88_noxref_g ) capacitor c=0.0180032f \
 //x=28.165 //y=5.02 //x2=28.09 //y2=6.02
cc_3108 ( N_noxref_9_c_3663_n N_CLK_M89_noxref_g ) capacitor c=0.01736f \
 //x=29.105 //y=5.155 //x2=28.53 //y2=6.02
cc_3109 ( N_noxref_9_M88_noxref_d N_CLK_M89_noxref_g ) capacitor c=0.0180032f \
 //x=28.165 //y=5.02 //x2=28.53 //y2=6.02
cc_3110 ( N_noxref_9_c_3808_p N_CLK_c_5100_n ) capacitor c=0.00426767f \
 //x=28.31 //y=5.155 //x2=28.455 //y2=4.79
cc_3111 ( N_noxref_9_c_3657_n N_CLK_c_5101_n ) capacitor c=0.00322046f \
 //x=28.225 //y=5.155 //x2=28.12 //y2=4.7
cc_3112 ( N_noxref_9_c_3824_p N_RN_c_5861_n ) capacitor c=0.016327f //x=29.57 \
 //y=1.665 //x2=33.925 //y2=2.22
cc_3113 ( N_noxref_9_c_3671_n N_RN_c_5861_n ) capacitor c=0.0197307f //x=29.97 \
 //y=3.7 //x2=33.925 //y2=2.22
cc_3114 ( N_noxref_9_c_3634_n N_RN_c_5861_n ) capacitor c=0.0192695f //x=31.82 \
 //y=2.08 //x2=33.925 //y2=2.22
cc_3115 ( N_noxref_9_c_3640_n N_RN_c_5861_n ) capacitor c=0.011987f //x=31.52 \
 //y=1.915 //x2=33.925 //y2=2.22
cc_3116 ( N_noxref_9_c_3635_n N_RN_c_5882_n ) capacitor c=0.0192695f //x=44.77 \
 //y=2.08 //x2=45.765 //y2=2.22
cc_3117 ( N_noxref_9_c_3650_n N_RN_c_5882_n ) capacitor c=0.011987f //x=44.47 \
 //y=1.915 //x2=45.765 //y2=2.22
cc_3118 ( N_noxref_9_c_3635_n N_RN_c_5898_n ) capacitor c=0.00100368f \
 //x=44.77 //y=2.08 //x2=45.995 //y2=2.22
cc_3119 ( N_noxref_9_c_3650_n N_RN_c_5898_n ) capacitor c=2.11894e-19 \
 //x=44.47 //y=1.915 //x2=45.995 //y2=2.22
cc_3120 ( N_noxref_9_c_3708_n N_RN_c_5916_n ) capacitor c=0.0179999f \
 //x=44.655 //y=3.7 //x2=34.04 //y2=2.08
cc_3121 ( N_noxref_9_c_3634_n N_RN_c_5916_n ) capacitor c=9.0823e-19 //x=31.82 \
 //y=2.08 //x2=34.04 //y2=2.08
cc_3122 ( N_noxref_9_c_3708_n N_RN_c_5917_n ) capacitor c=0.0203405f \
 //x=44.655 //y=3.7 //x2=42.18 //y2=2.08
cc_3123 ( N_noxref_9_c_3635_n N_RN_c_5917_n ) capacitor c=7.66327e-19 \
 //x=44.77 //y=2.08 //x2=42.18 //y2=2.08
cc_3124 ( N_noxref_9_c_3708_n N_RN_c_5918_n ) capacitor c=0.00311593f \
 //x=44.655 //y=3.7 //x2=45.88 //y2=2.08
cc_3125 ( N_noxref_9_c_3635_n N_RN_c_5918_n ) capacitor c=0.0449982f //x=44.77 \
 //y=2.08 //x2=45.88 //y2=2.08
cc_3126 ( N_noxref_9_c_3650_n N_RN_c_5918_n ) capacitor c=0.00208635f \
 //x=44.47 //y=1.915 //x2=45.88 //y2=2.08
cc_3127 ( N_noxref_9_c_3751_p N_RN_c_5918_n ) capacitor c=0.00147352f \
 //x=45.335 //y=4.79 //x2=45.88 //y2=2.08
cc_3128 ( N_noxref_9_c_3688_n N_RN_c_5918_n ) capacitor c=0.00142741f \
 //x=45.045 //y=4.79 //x2=45.88 //y2=2.08
cc_3129 ( N_noxref_9_M108_noxref_g N_RN_M110_noxref_g ) capacitor c=0.0105869f \
 //x=44.97 //y=6.02 //x2=45.85 //y2=6.02
cc_3130 ( N_noxref_9_M109_noxref_g N_RN_M110_noxref_g ) capacitor c=0.10632f \
 //x=45.41 //y=6.02 //x2=45.85 //y2=6.02
cc_3131 ( N_noxref_9_M109_noxref_g N_RN_M111_noxref_g ) capacitor c=0.0101598f \
 //x=45.41 //y=6.02 //x2=46.29 //y2=6.02
cc_3132 ( N_noxref_9_c_3646_n N_RN_c_6149_n ) capacitor c=5.72482e-19 \
 //x=44.47 //y=0.875 //x2=45.445 //y2=0.91
cc_3133 ( N_noxref_9_c_3648_n N_RN_c_6149_n ) capacitor c=0.00149976f \
 //x=44.47 //y=1.22 //x2=45.445 //y2=0.91
cc_3134 ( N_noxref_9_c_3653_n N_RN_c_6149_n ) capacitor c=0.0160123f //x=45 \
 //y=0.875 //x2=45.445 //y2=0.91
cc_3135 ( N_noxref_9_c_3649_n N_RN_c_6152_n ) capacitor c=0.00111227f \
 //x=44.47 //y=1.53 //x2=45.445 //y2=1.22
cc_3136 ( N_noxref_9_c_3655_n N_RN_c_6152_n ) capacitor c=0.0124075f //x=45 \
 //y=1.22 //x2=45.445 //y2=1.22
cc_3137 ( N_noxref_9_c_3653_n N_RN_c_6154_n ) capacitor c=0.00103227f //x=45 \
 //y=0.875 //x2=45.97 //y2=0.91
cc_3138 ( N_noxref_9_c_3655_n N_RN_c_6155_n ) capacitor c=0.0010154f //x=45 \
 //y=1.22 //x2=45.97 //y2=1.22
cc_3139 ( N_noxref_9_c_3655_n N_RN_c_6156_n ) capacitor c=9.23422e-19 //x=45 \
 //y=1.22 //x2=45.97 //y2=1.45
cc_3140 ( N_noxref_9_c_3635_n N_RN_c_6157_n ) capacitor c=0.00203769f \
 //x=44.77 //y=2.08 //x2=45.97 //y2=1.915
cc_3141 ( N_noxref_9_c_3650_n N_RN_c_6157_n ) capacitor c=0.00834532f \
 //x=44.47 //y=1.915 //x2=45.97 //y2=1.915
cc_3142 ( N_noxref_9_c_3635_n N_RN_c_6159_n ) capacitor c=0.00183762f \
 //x=44.77 //y=2.08 //x2=45.88 //y2=4.7
cc_3143 ( N_noxref_9_c_3751_p N_RN_c_6159_n ) capacitor c=0.0168581f \
 //x=45.335 //y=4.79 //x2=45.88 //y2=4.7
cc_3144 ( N_noxref_9_c_3688_n N_RN_c_6159_n ) capacitor c=0.00484466f \
 //x=45.045 //y=4.79 //x2=45.88 //y2=4.7
cc_3145 ( N_noxref_9_c_3635_n N_noxref_17_c_7301_n ) capacitor c=0.00121487f \
 //x=44.77 //y=2.08 //x2=46.99 //y2=2.08
cc_3146 ( N_noxref_9_c_3705_n N_noxref_20_c_8516_n ) capacitor c=0.0108826f \
 //x=31.705 //y=3.7 //x2=83.505 //y2=2.96
cc_3147 ( N_noxref_9_c_3706_n N_noxref_20_c_8516_n ) capacitor c=7.98411e-19 \
 //x=30.085 //y=3.7 //x2=83.505 //y2=2.96
cc_3148 ( N_noxref_9_c_3708_n N_noxref_20_c_8516_n ) capacitor c=0.308195f \
 //x=44.655 //y=3.7 //x2=83.505 //y2=2.96
cc_3149 ( N_noxref_9_c_3713_n N_noxref_20_c_8516_n ) capacitor c=5.46757e-19 \
 //x=31.935 //y=3.7 //x2=83.505 //y2=2.96
cc_3150 ( N_noxref_9_c_3671_n N_noxref_20_c_8516_n ) capacitor c=0.0187656f \
 //x=29.97 //y=3.7 //x2=83.505 //y2=2.96
cc_3151 ( N_noxref_9_c_3634_n N_noxref_20_c_8516_n ) capacitor c=0.0197816f \
 //x=31.82 //y=2.08 //x2=83.505 //y2=2.96
cc_3152 ( N_noxref_9_c_3635_n N_noxref_20_c_8516_n ) capacitor c=0.0224129f \
 //x=44.77 //y=2.08 //x2=83.505 //y2=2.96
cc_3153 ( N_noxref_9_c_3661_n N_noxref_20_c_8540_n ) capacitor c=2.97874e-19 \
 //x=27.515 //y=5.155 //x2=25.16 //y2=2.96
cc_3154 ( N_noxref_9_M18_noxref_d N_noxref_33_M16_noxref_s ) capacitor \
 c=0.00309936f //x=29.295 //y=0.915 //x2=26.355 //y2=0.375
cc_3155 ( N_noxref_9_c_3633_n N_noxref_34_c_9831_n ) capacitor c=0.00457167f \
 //x=29.885 //y=1.665 //x2=29.885 //y2=0.54
cc_3156 ( N_noxref_9_M18_noxref_d N_noxref_34_c_9831_n ) capacitor \
 c=0.0115903f //x=29.295 //y=0.915 //x2=29.885 //y2=0.54
cc_3157 ( N_noxref_9_c_3824_p N_noxref_34_c_9843_n ) capacitor c=0.0200405f \
 //x=29.57 //y=1.665 //x2=29 //y2=0.995
cc_3158 ( N_noxref_9_M18_noxref_d N_noxref_34_M17_noxref_d ) capacitor \
 c=5.27807e-19 //x=29.295 //y=0.915 //x2=27.76 //y2=0.91
cc_3159 ( N_noxref_9_c_3633_n N_noxref_34_M18_noxref_s ) capacitor \
 c=0.0196084f //x=29.885 //y=1.665 //x2=28.865 //y2=0.375
cc_3160 ( N_noxref_9_M18_noxref_d N_noxref_34_M18_noxref_s ) capacitor \
 c=0.0426368f //x=29.295 //y=0.915 //x2=28.865 //y2=0.375
cc_3161 ( N_noxref_9_c_3633_n N_noxref_35_c_9894_n ) capacitor c=3.84569e-19 \
 //x=29.885 //y=1.665 //x2=31.3 //y2=1.505
cc_3162 ( N_noxref_9_c_3640_n N_noxref_35_c_9894_n ) capacitor c=0.0034165f \
 //x=31.52 //y=1.915 //x2=31.3 //y2=1.505
cc_3163 ( N_noxref_9_c_3634_n N_noxref_35_c_9878_n ) capacitor c=0.0115578f \
 //x=31.82 //y=2.08 //x2=32.185 //y2=1.59
cc_3164 ( N_noxref_9_c_3639_n N_noxref_35_c_9878_n ) capacitor c=0.00697148f \
 //x=31.52 //y=1.53 //x2=32.185 //y2=1.59
cc_3165 ( N_noxref_9_c_3640_n N_noxref_35_c_9878_n ) capacitor c=0.0204849f \
 //x=31.52 //y=1.915 //x2=32.185 //y2=1.59
cc_3166 ( N_noxref_9_c_3642_n N_noxref_35_c_9878_n ) capacitor c=0.00610316f \
 //x=31.895 //y=1.375 //x2=32.185 //y2=1.59
cc_3167 ( N_noxref_9_c_3645_n N_noxref_35_c_9878_n ) capacitor c=0.00698822f \
 //x=32.05 //y=1.22 //x2=32.185 //y2=1.59
cc_3168 ( N_noxref_9_c_3636_n N_noxref_35_M19_noxref_s ) capacitor \
 c=0.0327271f //x=31.52 //y=0.875 //x2=31.165 //y2=0.375
cc_3169 ( N_noxref_9_c_3639_n N_noxref_35_M19_noxref_s ) capacitor \
 c=7.99997e-19 //x=31.52 //y=1.53 //x2=31.165 //y2=0.375
cc_3170 ( N_noxref_9_c_3640_n N_noxref_35_M19_noxref_s ) capacitor \
 c=0.00122123f //x=31.52 //y=1.915 //x2=31.165 //y2=0.375
cc_3171 ( N_noxref_9_c_3643_n N_noxref_35_M19_noxref_s ) capacitor \
 c=0.0121427f //x=32.05 //y=0.875 //x2=31.165 //y2=0.375
cc_3172 ( N_noxref_9_M18_noxref_d N_noxref_35_M19_noxref_s ) capacitor \
 c=2.55333e-19 //x=29.295 //y=0.915 //x2=31.165 //y2=0.375
cc_3173 ( N_noxref_9_c_3650_n N_noxref_40_c_10148_n ) capacitor c=0.0034165f \
 //x=44.47 //y=1.915 //x2=44.25 //y2=1.505
cc_3174 ( N_noxref_9_c_3635_n N_noxref_40_c_10133_n ) capacitor c=0.0115578f \
 //x=44.77 //y=2.08 //x2=45.135 //y2=1.59
cc_3175 ( N_noxref_9_c_3649_n N_noxref_40_c_10133_n ) capacitor c=0.00697148f \
 //x=44.47 //y=1.53 //x2=45.135 //y2=1.59
cc_3176 ( N_noxref_9_c_3650_n N_noxref_40_c_10133_n ) capacitor c=0.0204849f \
 //x=44.47 //y=1.915 //x2=45.135 //y2=1.59
cc_3177 ( N_noxref_9_c_3652_n N_noxref_40_c_10133_n ) capacitor c=0.00610316f \
 //x=44.845 //y=1.375 //x2=45.135 //y2=1.59
cc_3178 ( N_noxref_9_c_3655_n N_noxref_40_c_10133_n ) capacitor c=0.00698822f \
 //x=45 //y=1.22 //x2=45.135 //y2=1.59
cc_3179 ( N_noxref_9_c_3646_n N_noxref_40_M27_noxref_s ) capacitor \
 c=0.0327271f //x=44.47 //y=0.875 //x2=44.115 //y2=0.375
cc_3180 ( N_noxref_9_c_3649_n N_noxref_40_M27_noxref_s ) capacitor \
 c=7.99997e-19 //x=44.47 //y=1.53 //x2=44.115 //y2=0.375
cc_3181 ( N_noxref_9_c_3650_n N_noxref_40_M27_noxref_s ) capacitor \
 c=0.00122123f //x=44.47 //y=1.915 //x2=44.115 //y2=0.375
cc_3182 ( N_noxref_9_c_3653_n N_noxref_40_M27_noxref_s ) capacitor \
 c=0.0121427f //x=45 //y=0.875 //x2=44.115 //y2=0.375
cc_3183 ( N_noxref_10_c_3951_p N_noxref_11_c_4079_n ) capacitor c=0.176083f \
 //x=49.465 //y=3.7 //x2=50.205 //y2=4.07
cc_3184 ( N_noxref_10_c_3946_n N_noxref_11_c_4079_n ) capacitor c=0.0294294f \
 //x=47.845 //y=3.7 //x2=50.205 //y2=4.07
cc_3185 ( N_noxref_10_c_3922_n N_noxref_11_c_4079_n ) capacitor c=0.0200135f \
 //x=47.73 //y=3.7 //x2=50.205 //y2=4.07
cc_3186 ( N_noxref_10_c_3896_n N_noxref_11_c_4079_n ) capacitor c=0.0216244f \
 //x=49.58 //y=2.08 //x2=50.205 //y2=4.07
cc_3187 ( N_noxref_10_c_3912_n N_noxref_11_c_4097_n ) capacitor c=3.10026e-19 \
 //x=45.275 //y=5.155 //x2=42.835 //y2=5.155
cc_3188 ( N_noxref_10_c_3896_n N_noxref_11_c_4228_n ) capacitor c=0.00400249f \
 //x=49.58 //y=2.08 //x2=50.32 //y2=4.535
cc_3189 ( N_noxref_10_c_3930_n N_noxref_11_c_4228_n ) capacitor c=0.00417994f \
 //x=49.58 //y=4.7 //x2=50.32 //y2=4.535
cc_3190 ( N_noxref_10_c_3951_p N_noxref_11_c_4062_n ) capacitor c=0.00720056f \
 //x=49.465 //y=3.7 //x2=50.32 //y2=2.08
cc_3191 ( N_noxref_10_c_3922_n N_noxref_11_c_4062_n ) capacitor c=9.52757e-19 \
 //x=47.73 //y=3.7 //x2=50.32 //y2=2.08
cc_3192 ( N_noxref_10_c_3896_n N_noxref_11_c_4062_n ) capacitor c=0.07134f \
 //x=49.58 //y=2.08 //x2=50.32 //y2=2.08
cc_3193 ( N_noxref_10_c_3901_n N_noxref_11_c_4062_n ) capacitor c=0.00284029f \
 //x=49.385 //y=1.915 //x2=50.32 //y2=2.08
cc_3194 ( N_noxref_10_M114_noxref_g N_noxref_11_M116_noxref_g ) capacitor \
 c=0.0104611f //x=49.48 //y=6.02 //x2=50.36 //y2=6.02
cc_3195 ( N_noxref_10_M115_noxref_g N_noxref_11_M116_noxref_g ) capacitor \
 c=0.106811f //x=49.92 //y=6.02 //x2=50.36 //y2=6.02
cc_3196 ( N_noxref_10_M115_noxref_g N_noxref_11_M117_noxref_g ) capacitor \
 c=0.0100341f //x=49.92 //y=6.02 //x2=50.8 //y2=6.02
cc_3197 ( N_noxref_10_c_3897_n N_noxref_11_c_4237_n ) capacitor c=4.86506e-19 \
 //x=49.385 //y=0.865 //x2=50.355 //y2=0.905
cc_3198 ( N_noxref_10_c_3899_n N_noxref_11_c_4237_n ) capacitor c=0.00152104f \
 //x=49.385 //y=1.21 //x2=50.355 //y2=0.905
cc_3199 ( N_noxref_10_c_3904_n N_noxref_11_c_4237_n ) capacitor c=0.0151475f \
 //x=49.915 //y=0.865 //x2=50.355 //y2=0.905
cc_3200 ( N_noxref_10_c_3900_n N_noxref_11_c_4240_n ) capacitor c=0.00109982f \
 //x=49.385 //y=1.52 //x2=50.355 //y2=1.25
cc_3201 ( N_noxref_10_c_3906_n N_noxref_11_c_4240_n ) capacitor c=0.0111064f \
 //x=49.915 //y=1.21 //x2=50.355 //y2=1.25
cc_3202 ( N_noxref_10_c_3900_n N_noxref_11_c_4242_n ) capacitor c=9.57794e-19 \
 //x=49.385 //y=1.52 //x2=50.355 //y2=1.56
cc_3203 ( N_noxref_10_c_3901_n N_noxref_11_c_4242_n ) capacitor c=0.00662747f \
 //x=49.385 //y=1.915 //x2=50.355 //y2=1.56
cc_3204 ( N_noxref_10_c_3906_n N_noxref_11_c_4242_n ) capacitor c=0.00862358f \
 //x=49.915 //y=1.21 //x2=50.355 //y2=1.56
cc_3205 ( N_noxref_10_c_3904_n N_noxref_11_c_4245_n ) capacitor c=0.00124821f \
 //x=49.915 //y=0.865 //x2=50.885 //y2=0.905
cc_3206 ( N_noxref_10_c_3906_n N_noxref_11_c_4246_n ) capacitor c=0.00200715f \
 //x=49.915 //y=1.21 //x2=50.885 //y2=1.25
cc_3207 ( N_noxref_10_c_3896_n N_noxref_11_c_4247_n ) capacitor c=0.00282278f \
 //x=49.58 //y=2.08 //x2=50.32 //y2=2.08
cc_3208 ( N_noxref_10_c_3901_n N_noxref_11_c_4247_n ) capacitor c=0.0172771f \
 //x=49.385 //y=1.915 //x2=50.32 //y2=2.08
cc_3209 ( N_noxref_10_c_3896_n N_noxref_11_c_4249_n ) capacitor c=0.00344981f \
 //x=49.58 //y=2.08 //x2=50.35 //y2=4.7
cc_3210 ( N_noxref_10_c_3930_n N_noxref_11_c_4249_n ) capacitor c=0.0293367f \
 //x=49.58 //y=4.7 //x2=50.35 //y2=4.7
cc_3211 ( N_noxref_10_c_3922_n N_D_c_4442_n ) capacitor c=0.0165903f //x=47.73 \
 //y=3.7 //x2=58.715 //y2=2.59
cc_3212 ( N_noxref_10_c_3896_n N_D_c_4442_n ) capacitor c=0.0177872f //x=49.58 \
 //y=2.08 //x2=58.715 //y2=2.59
cc_3213 ( N_noxref_10_c_3951_p N_CLK_c_4862_n ) capacitor c=0.0103783f \
 //x=49.465 //y=3.7 //x2=53.905 //y2=4.44
cc_3214 ( N_noxref_10_c_3946_n N_CLK_c_4862_n ) capacitor c=7.95009e-19 \
 //x=47.845 //y=3.7 //x2=53.905 //y2=4.44
cc_3215 ( N_noxref_10_c_3908_n N_CLK_c_4862_n ) capacitor c=0.032141f \
 //x=45.985 //y=5.155 //x2=53.905 //y2=4.44
cc_3216 ( N_noxref_10_c_3912_n N_CLK_c_4862_n ) capacitor c=0.0230136f \
 //x=45.275 //y=5.155 //x2=53.905 //y2=4.44
cc_3217 ( N_noxref_10_c_3918_n N_CLK_c_4862_n ) capacitor c=0.0183122f \
 //x=47.645 //y=5.155 //x2=53.905 //y2=4.44
cc_3218 ( N_noxref_10_c_3922_n N_CLK_c_4862_n ) capacitor c=0.0210274f \
 //x=47.73 //y=3.7 //x2=53.905 //y2=4.44
cc_3219 ( N_noxref_10_c_3896_n N_CLK_c_4862_n ) capacitor c=0.0198304f \
 //x=49.58 //y=2.08 //x2=53.905 //y2=4.44
cc_3220 ( N_noxref_10_c_3930_n N_CLK_c_4862_n ) capacitor c=0.0107057f \
 //x=49.58 //y=4.7 //x2=53.905 //y2=4.44
cc_3221 ( N_noxref_10_c_3989_p N_RN_c_5887_n ) capacitor c=0.016327f //x=47.33 \
 //y=1.665 //x2=59.825 //y2=2.22
cc_3222 ( N_noxref_10_c_3922_n N_RN_c_5887_n ) capacitor c=0.0197307f \
 //x=47.73 //y=3.7 //x2=59.825 //y2=2.22
cc_3223 ( N_noxref_10_c_3896_n N_RN_c_5887_n ) capacitor c=0.0185012f \
 //x=49.58 //y=2.08 //x2=59.825 //y2=2.22
cc_3224 ( N_noxref_10_c_3901_n N_RN_c_5887_n ) capacitor c=0.00894156f \
 //x=49.385 //y=1.915 //x2=59.825 //y2=2.22
cc_3225 ( N_noxref_10_c_3908_n N_RN_c_5918_n ) capacitor c=0.0144268f \
 //x=45.985 //y=5.155 //x2=45.88 //y2=2.08
cc_3226 ( N_noxref_10_c_3922_n N_RN_c_5918_n ) capacitor c=0.00255845f \
 //x=47.73 //y=3.7 //x2=45.88 //y2=2.08
cc_3227 ( N_noxref_10_c_3908_n N_RN_M110_noxref_g ) capacitor c=0.0165266f \
 //x=45.985 //y=5.155 //x2=45.85 //y2=6.02
cc_3228 ( N_noxref_10_M110_noxref_d N_RN_M110_noxref_g ) capacitor \
 c=0.0180032f //x=45.925 //y=5.02 //x2=45.85 //y2=6.02
cc_3229 ( N_noxref_10_c_3914_n N_RN_M111_noxref_g ) capacitor c=0.01736f \
 //x=46.865 //y=5.155 //x2=46.29 //y2=6.02
cc_3230 ( N_noxref_10_M110_noxref_d N_RN_M111_noxref_g ) capacitor \
 c=0.0180032f //x=45.925 //y=5.02 //x2=46.29 //y2=6.02
cc_3231 ( N_noxref_10_c_3999_p N_RN_c_6172_n ) capacitor c=0.00426767f \
 //x=46.07 //y=5.155 //x2=46.215 //y2=4.79
cc_3232 ( N_noxref_10_c_3908_n N_RN_c_6159_n ) capacitor c=0.00322054f \
 //x=45.985 //y=5.155 //x2=45.88 //y2=4.7
cc_3233 ( N_noxref_10_c_3951_p N_noxref_17_c_7491_n ) capacitor c=0.17564f \
 //x=49.465 //y=3.7 //x2=50.945 //y2=3.33
cc_3234 ( N_noxref_10_c_3946_n N_noxref_17_c_7491_n ) capacitor c=0.0294746f \
 //x=47.845 //y=3.7 //x2=50.945 //y2=3.33
cc_3235 ( N_noxref_10_c_3922_n N_noxref_17_c_7491_n ) capacitor c=0.0206036f \
 //x=47.73 //y=3.7 //x2=50.945 //y2=3.33
cc_3236 ( N_noxref_10_c_3896_n N_noxref_17_c_7491_n ) capacitor c=0.020575f \
 //x=49.58 //y=2.08 //x2=50.945 //y2=3.33
cc_3237 ( N_noxref_10_c_3922_n N_noxref_17_c_7495_n ) capacitor c=0.00117715f \
 //x=47.73 //y=3.7 //x2=47.105 //y2=3.33
cc_3238 ( N_noxref_10_c_3946_n N_noxref_17_c_7301_n ) capacitor c=0.00456439f \
 //x=47.845 //y=3.7 //x2=46.99 //y2=2.08
cc_3239 ( N_noxref_10_c_3922_n N_noxref_17_c_7301_n ) capacitor c=0.0769087f \
 //x=47.73 //y=3.7 //x2=46.99 //y2=2.08
cc_3240 ( N_noxref_10_c_3896_n N_noxref_17_c_7301_n ) capacitor c=8.82143e-19 \
 //x=49.58 //y=2.08 //x2=46.99 //y2=2.08
cc_3241 ( N_noxref_10_c_4009_p N_noxref_17_c_7301_n ) capacitor c=0.0166016f \
 //x=46.95 //y=5.155 //x2=46.99 //y2=2.08
cc_3242 ( N_noxref_10_M115_noxref_g N_noxref_17_c_7373_n ) capacitor \
 c=0.0169521f //x=49.92 //y=6.02 //x2=50.495 //y2=5.2
cc_3243 ( N_noxref_10_c_3896_n N_noxref_17_c_7377_n ) capacitor c=0.00521572f \
 //x=49.58 //y=2.08 //x2=49.785 //y2=5.2
cc_3244 ( N_noxref_10_M114_noxref_g N_noxref_17_c_7377_n ) capacitor \
 c=0.0177326f //x=49.48 //y=6.02 //x2=49.785 //y2=5.2
cc_3245 ( N_noxref_10_c_3930_n N_noxref_17_c_7377_n ) capacitor c=0.00581252f \
 //x=49.58 //y=4.7 //x2=49.785 //y2=5.2
cc_3246 ( N_noxref_10_c_3922_n N_noxref_17_c_7303_n ) capacitor c=3.52729e-19 \
 //x=47.73 //y=3.7 //x2=51.06 //y2=3.33
cc_3247 ( N_noxref_10_c_3896_n N_noxref_17_c_7303_n ) capacitor c=0.00318542f \
 //x=49.58 //y=2.08 //x2=51.06 //y2=3.33
cc_3248 ( N_noxref_10_c_3914_n N_noxref_17_M112_noxref_g ) capacitor \
 c=0.01736f //x=46.865 //y=5.155 //x2=46.73 //y2=6.02
cc_3249 ( N_noxref_10_M112_noxref_d N_noxref_17_M112_noxref_g ) capacitor \
 c=0.0180032f //x=46.805 //y=5.02 //x2=46.73 //y2=6.02
cc_3250 ( N_noxref_10_c_3918_n N_noxref_17_M113_noxref_g ) capacitor \
 c=0.0194981f //x=47.645 //y=5.155 //x2=47.17 //y2=6.02
cc_3251 ( N_noxref_10_M112_noxref_d N_noxref_17_M113_noxref_g ) capacitor \
 c=0.0194246f //x=46.805 //y=5.02 //x2=47.17 //y2=6.02
cc_3252 ( N_noxref_10_M29_noxref_d N_noxref_17_c_7510_n ) capacitor \
 c=0.00217566f //x=47.055 //y=0.915 //x2=46.98 //y2=0.915
cc_3253 ( N_noxref_10_M29_noxref_d N_noxref_17_c_7511_n ) capacitor \
 c=0.0034598f //x=47.055 //y=0.915 //x2=46.98 //y2=1.26
cc_3254 ( N_noxref_10_M29_noxref_d N_noxref_17_c_7512_n ) capacitor \
 c=0.00546784f //x=47.055 //y=0.915 //x2=46.98 //y2=1.57
cc_3255 ( N_noxref_10_M29_noxref_d N_noxref_17_c_7513_n ) capacitor \
 c=0.00241102f //x=47.055 //y=0.915 //x2=47.355 //y2=0.76
cc_3256 ( N_noxref_10_c_3895_n N_noxref_17_c_7514_n ) capacitor c=0.00371277f \
 //x=47.645 //y=1.665 //x2=47.355 //y2=1.415
cc_3257 ( N_noxref_10_M29_noxref_d N_noxref_17_c_7514_n ) capacitor \
 c=0.0138621f //x=47.055 //y=0.915 //x2=47.355 //y2=1.415
cc_3258 ( N_noxref_10_M29_noxref_d N_noxref_17_c_7516_n ) capacitor \
 c=0.00219619f //x=47.055 //y=0.915 //x2=47.51 //y2=0.915
cc_3259 ( N_noxref_10_c_3895_n N_noxref_17_c_7517_n ) capacitor c=0.00457401f \
 //x=47.645 //y=1.665 //x2=47.51 //y2=1.26
cc_3260 ( N_noxref_10_M29_noxref_d N_noxref_17_c_7517_n ) capacitor \
 c=0.00603828f //x=47.055 //y=0.915 //x2=47.51 //y2=1.26
cc_3261 ( N_noxref_10_c_3922_n N_noxref_17_c_7519_n ) capacitor c=0.00709342f \
 //x=47.73 //y=3.7 //x2=46.99 //y2=2.08
cc_3262 ( N_noxref_10_c_3922_n N_noxref_17_c_7520_n ) capacitor c=0.00283672f \
 //x=47.73 //y=3.7 //x2=46.99 //y2=1.915
cc_3263 ( N_noxref_10_M29_noxref_d N_noxref_17_c_7520_n ) capacitor \
 c=0.00661782f //x=47.055 //y=0.915 //x2=46.99 //y2=1.915
cc_3264 ( N_noxref_10_c_3918_n N_noxref_17_c_7522_n ) capacitor c=0.00201851f \
 //x=47.645 //y=5.155 //x2=46.99 //y2=4.7
cc_3265 ( N_noxref_10_c_3922_n N_noxref_17_c_7522_n ) capacitor c=0.013844f \
 //x=47.73 //y=3.7 //x2=46.99 //y2=4.7
cc_3266 ( N_noxref_10_c_4009_p N_noxref_17_c_7522_n ) capacitor c=0.00475601f \
 //x=46.95 //y=5.155 //x2=46.99 //y2=4.7
cc_3267 ( N_noxref_10_M115_noxref_g N_noxref_17_M114_noxref_d ) capacitor \
 c=0.0173476f //x=49.92 //y=6.02 //x2=49.555 //y2=5.02
cc_3268 ( N_noxref_10_c_3951_p N_noxref_20_c_8516_n ) capacitor c=0.0119727f \
 //x=49.465 //y=3.7 //x2=83.505 //y2=2.96
cc_3269 ( N_noxref_10_c_3946_n N_noxref_20_c_8516_n ) capacitor c=7.98411e-19 \
 //x=47.845 //y=3.7 //x2=83.505 //y2=2.96
cc_3270 ( N_noxref_10_c_3922_n N_noxref_20_c_8516_n ) capacitor c=0.0187656f \
 //x=47.73 //y=3.7 //x2=83.505 //y2=2.96
cc_3271 ( N_noxref_10_c_3896_n N_noxref_20_c_8516_n ) capacitor c=0.0187412f \
 //x=49.58 //y=2.08 //x2=83.505 //y2=2.96
cc_3272 ( N_noxref_10_M29_noxref_d N_noxref_40_M27_noxref_s ) capacitor \
 c=0.00309936f //x=47.055 //y=0.915 //x2=44.115 //y2=0.375
cc_3273 ( N_noxref_10_c_3895_n N_noxref_41_c_10190_n ) capacitor c=0.00457167f \
 //x=47.645 //y=1.665 //x2=47.645 //y2=0.54
cc_3274 ( N_noxref_10_M29_noxref_d N_noxref_41_c_10190_n ) capacitor \
 c=0.0115903f //x=47.055 //y=0.915 //x2=47.645 //y2=0.54
cc_3275 ( N_noxref_10_c_3989_p N_noxref_41_c_10200_n ) capacitor c=0.020048f \
 //x=47.33 //y=1.665 //x2=46.76 //y2=0.995
cc_3276 ( N_noxref_10_M29_noxref_d N_noxref_41_M28_noxref_d ) capacitor \
 c=5.27807e-19 //x=47.055 //y=0.915 //x2=45.52 //y2=0.91
cc_3277 ( N_noxref_10_c_3895_n N_noxref_41_M29_noxref_s ) capacitor \
 c=0.0196084f //x=47.645 //y=1.665 //x2=46.625 //y2=0.375
cc_3278 ( N_noxref_10_M29_noxref_d N_noxref_41_M29_noxref_s ) capacitor \
 c=0.0426444f //x=47.055 //y=0.915 //x2=46.625 //y2=0.375
cc_3279 ( N_noxref_10_c_3895_n N_noxref_42_c_10255_n ) capacitor c=3.04182e-19 \
 //x=47.645 //y=1.665 //x2=49.165 //y2=1.495
cc_3280 ( N_noxref_10_c_3901_n N_noxref_42_c_10255_n ) capacitor c=0.0034165f \
 //x=49.385 //y=1.915 //x2=49.165 //y2=1.495
cc_3281 ( N_noxref_10_c_3896_n N_noxref_42_c_10237_n ) capacitor c=0.0111916f \
 //x=49.58 //y=2.08 //x2=50.05 //y2=1.58
cc_3282 ( N_noxref_10_c_3900_n N_noxref_42_c_10237_n ) capacitor c=0.00696403f \
 //x=49.385 //y=1.52 //x2=50.05 //y2=1.58
cc_3283 ( N_noxref_10_c_3901_n N_noxref_42_c_10237_n ) capacitor c=0.0174694f \
 //x=49.385 //y=1.915 //x2=50.05 //y2=1.58
cc_3284 ( N_noxref_10_c_3903_n N_noxref_42_c_10237_n ) capacitor c=0.00776811f \
 //x=49.76 //y=1.365 //x2=50.05 //y2=1.58
cc_3285 ( N_noxref_10_c_3906_n N_noxref_42_c_10237_n ) capacitor c=0.00339872f \
 //x=49.915 //y=1.21 //x2=50.05 //y2=1.58
cc_3286 ( N_noxref_10_c_3901_n N_noxref_42_c_10244_n ) capacitor c=6.71402e-19 \
 //x=49.385 //y=1.915 //x2=50.135 //y2=1.495
cc_3287 ( N_noxref_10_c_3897_n N_noxref_42_M30_noxref_s ) capacitor \
 c=0.0327502f //x=49.385 //y=0.865 //x2=49.03 //y2=0.365
cc_3288 ( N_noxref_10_c_3900_n N_noxref_42_M30_noxref_s ) capacitor \
 c=3.48408e-19 //x=49.385 //y=1.52 //x2=49.03 //y2=0.365
cc_3289 ( N_noxref_10_c_3904_n N_noxref_42_M30_noxref_s ) capacitor \
 c=0.0120759f //x=49.915 //y=0.865 //x2=49.03 //y2=0.365
cc_3290 ( N_noxref_11_c_4075_n N_D_c_4434_n ) capacitor c=0.011848f //x=37.255 \
 //y=4.07 //x2=32.815 //y2=2.59
cc_3291 ( N_noxref_11_c_4077_n N_D_c_4434_n ) capacitor c=4.25679e-19 \
 //x=27.125 //y=4.07 //x2=32.815 //y2=2.59
cc_3292 ( N_noxref_11_c_4058_n N_D_c_4434_n ) capacitor c=0.0188253f //x=27.01 \
 //y=2.08 //x2=32.815 //y2=2.59
cc_3293 ( N_noxref_11_c_4079_n N_D_c_4442_n ) capacitor c=0.01173f //x=50.205 \
 //y=4.07 //x2=58.715 //y2=2.59
cc_3294 ( N_noxref_11_c_4059_n N_D_c_4442_n ) capacitor c=0.0169223f //x=37.37 \
 //y=2.08 //x2=58.715 //y2=2.59
cc_3295 ( N_noxref_11_c_4101_n N_D_c_4442_n ) capacitor c=0.0165903f //x=42.92 \
 //y=4.07 //x2=58.715 //y2=2.59
cc_3296 ( N_noxref_11_c_4062_n N_D_c_4442_n ) capacitor c=0.0169223f //x=50.32 \
 //y=2.08 //x2=58.715 //y2=2.59
cc_3297 ( N_noxref_11_c_4075_n N_D_c_4449_n ) capacitor c=0.0190126f \
 //x=37.255 //y=4.07 //x2=32.93 //y2=2.08
cc_3298 ( N_noxref_11_c_4075_n N_CLK_c_4826_n ) capacitor c=0.076217f \
 //x=37.255 //y=4.07 //x2=28.005 //y2=4.44
cc_3299 ( N_noxref_11_c_4077_n N_CLK_c_4826_n ) capacitor c=0.0290178f \
 //x=27.125 //y=4.07 //x2=28.005 //y2=4.44
cc_3300 ( N_noxref_11_c_4058_n N_CLK_c_4826_n ) capacitor c=0.0227055f \
 //x=27.01 //y=2.08 //x2=28.005 //y2=4.44
cc_3301 ( N_noxref_11_c_4118_n N_CLK_c_4826_n ) capacitor c=0.0166959f \
 //x=27.285 //y=4.79 //x2=28.005 //y2=4.44
cc_3302 ( N_noxref_11_c_4075_n N_CLK_c_4844_n ) capacitor c=0.784553f \
 //x=37.255 //y=4.07 //x2=40.955 //y2=4.44
cc_3303 ( N_noxref_11_c_4078_n N_CLK_c_4844_n ) capacitor c=0.302855f \
 //x=42.805 //y=4.07 //x2=40.955 //y2=4.44
cc_3304 ( N_noxref_11_c_4144_n N_CLK_c_4844_n ) capacitor c=0.0263375f \
 //x=37.485 //y=4.07 //x2=40.955 //y2=4.44
cc_3305 ( N_noxref_11_c_4146_n N_CLK_c_4844_n ) capacitor c=0.0016972f \
 //x=37.37 //y=4.535 //x2=40.955 //y2=4.44
cc_3306 ( N_noxref_11_c_4059_n N_CLK_c_4844_n ) capacitor c=0.0207534f \
 //x=37.37 //y=2.08 //x2=40.955 //y2=4.44
cc_3307 ( N_noxref_11_c_4091_n N_CLK_c_4844_n ) capacitor c=0.0219114f \
 //x=40.465 //y=5.155 //x2=40.955 //y2=4.44
cc_3308 ( N_noxref_11_c_4190_n N_CLK_c_4844_n ) capacitor c=0.00960248f \
 //x=37.775 //y=4.79 //x2=40.955 //y2=4.44
cc_3309 ( N_noxref_11_c_4167_n N_CLK_c_4844_n ) capacitor c=0.00203982f \
 //x=37.4 //y=4.7 //x2=40.955 //y2=4.44
cc_3310 ( N_noxref_11_c_4075_n N_CLK_c_4861_n ) capacitor c=0.026534f \
 //x=37.255 //y=4.07 //x2=28.235 //y2=4.44
cc_3311 ( N_noxref_11_c_4058_n N_CLK_c_4861_n ) capacitor c=0.00153281f \
 //x=27.01 //y=2.08 //x2=28.235 //y2=4.44
cc_3312 ( N_noxref_11_c_4078_n N_CLK_c_4862_n ) capacitor c=0.140035f \
 //x=42.805 //y=4.07 //x2=53.905 //y2=4.44
cc_3313 ( N_noxref_11_c_4079_n N_CLK_c_4862_n ) capacitor c=0.654031f \
 //x=50.205 //y=4.07 //x2=53.905 //y2=4.44
cc_3314 ( N_noxref_11_c_4081_n N_CLK_c_4862_n ) capacitor c=0.0265915f \
 //x=43.035 //y=4.07 //x2=53.905 //y2=4.44
cc_3315 ( N_noxref_11_c_4097_n N_CLK_c_4862_n ) capacitor c=0.0183122f \
 //x=42.835 //y=5.155 //x2=53.905 //y2=4.44
cc_3316 ( N_noxref_11_c_4101_n N_CLK_c_4862_n ) capacitor c=0.022862f \
 //x=42.92 //y=4.07 //x2=53.905 //y2=4.44
cc_3317 ( N_noxref_11_c_4228_n N_CLK_c_4862_n ) capacitor c=0.0016972f \
 //x=50.32 //y=4.535 //x2=53.905 //y2=4.44
cc_3318 ( N_noxref_11_c_4062_n N_CLK_c_4862_n ) capacitor c=0.0207534f \
 //x=50.32 //y=2.08 //x2=53.905 //y2=4.44
cc_3319 ( N_noxref_11_c_4280_p N_CLK_c_4862_n ) capacitor c=0.0311227f \
 //x=41.26 //y=5.155 //x2=53.905 //y2=4.44
cc_3320 ( N_noxref_11_c_4281_p N_CLK_c_4862_n ) capacitor c=0.00720343f \
 //x=50.725 //y=4.79 //x2=53.905 //y2=4.44
cc_3321 ( N_noxref_11_c_4249_n N_CLK_c_4862_n ) capacitor c=0.0019199f \
 //x=50.35 //y=4.7 //x2=53.905 //y2=4.44
cc_3322 ( N_noxref_11_c_4078_n N_CLK_c_4879_n ) capacitor c=0.026534f \
 //x=42.805 //y=4.07 //x2=41.185 //y2=4.44
cc_3323 ( N_noxref_11_c_4087_n N_CLK_c_4879_n ) capacitor c=0.00241768f \
 //x=41.175 //y=5.155 //x2=41.185 //y2=4.44
cc_3324 ( N_noxref_11_c_4075_n N_CLK_c_4804_n ) capacitor c=0.0247116f \
 //x=37.255 //y=4.07 //x2=28.12 //y2=2.08
cc_3325 ( N_noxref_11_c_4077_n N_CLK_c_4804_n ) capacitor c=0.00128547f \
 //x=27.125 //y=4.07 //x2=28.12 //y2=2.08
cc_3326 ( N_noxref_11_c_4058_n N_CLK_c_4804_n ) capacitor c=0.0456686f \
 //x=27.01 //y=2.08 //x2=28.12 //y2=2.08
cc_3327 ( N_noxref_11_c_4068_n N_CLK_c_4804_n ) capacitor c=0.00210802f \
 //x=26.71 //y=1.915 //x2=28.12 //y2=2.08
cc_3328 ( N_noxref_11_c_4222_n N_CLK_c_4804_n ) capacitor c=0.00147352f \
 //x=27.575 //y=4.79 //x2=28.12 //y2=2.08
cc_3329 ( N_noxref_11_c_4118_n N_CLK_c_4804_n ) capacitor c=0.00141297f \
 //x=27.285 //y=4.79 //x2=28.12 //y2=2.08
cc_3330 ( N_noxref_11_c_4078_n N_CLK_c_4805_n ) capacitor c=0.0208526f \
 //x=42.805 //y=4.07 //x2=41.07 //y2=2.08
cc_3331 ( N_noxref_11_c_4087_n N_CLK_c_4805_n ) capacitor c=0.014564f \
 //x=41.175 //y=5.155 //x2=41.07 //y2=2.08
cc_3332 ( N_noxref_11_c_4101_n N_CLK_c_4805_n ) capacitor c=0.00256882f \
 //x=42.92 //y=4.07 //x2=41.07 //y2=2.08
cc_3333 ( N_noxref_11_M86_noxref_g N_CLK_M88_noxref_g ) capacitor c=0.0105869f \
 //x=27.21 //y=6.02 //x2=28.09 //y2=6.02
cc_3334 ( N_noxref_11_M87_noxref_g N_CLK_M88_noxref_g ) capacitor c=0.10632f \
 //x=27.65 //y=6.02 //x2=28.09 //y2=6.02
cc_3335 ( N_noxref_11_M87_noxref_g N_CLK_M89_noxref_g ) capacitor c=0.0101598f \
 //x=27.65 //y=6.02 //x2=28.53 //y2=6.02
cc_3336 ( N_noxref_11_c_4087_n N_CLK_M104_noxref_g ) capacitor c=0.016514f \
 //x=41.175 //y=5.155 //x2=41.04 //y2=6.02
cc_3337 ( N_noxref_11_M104_noxref_d N_CLK_M104_noxref_g ) capacitor \
 c=0.0180032f //x=41.115 //y=5.02 //x2=41.04 //y2=6.02
cc_3338 ( N_noxref_11_c_4093_n N_CLK_M105_noxref_g ) capacitor c=0.01736f \
 //x=42.055 //y=5.155 //x2=41.48 //y2=6.02
cc_3339 ( N_noxref_11_M104_noxref_d N_CLK_M105_noxref_g ) capacitor \
 c=0.0180032f //x=41.115 //y=5.02 //x2=41.48 //y2=6.02
cc_3340 ( N_noxref_11_c_4064_n N_CLK_c_5205_n ) capacitor c=5.72482e-19 \
 //x=26.71 //y=0.875 //x2=27.685 //y2=0.91
cc_3341 ( N_noxref_11_c_4066_n N_CLK_c_5205_n ) capacitor c=0.00149976f \
 //x=26.71 //y=1.22 //x2=27.685 //y2=0.91
cc_3342 ( N_noxref_11_c_4071_n N_CLK_c_5205_n ) capacitor c=0.0160123f \
 //x=27.24 //y=0.875 //x2=27.685 //y2=0.91
cc_3343 ( N_noxref_11_c_4067_n N_CLK_c_5208_n ) capacitor c=0.00111227f \
 //x=26.71 //y=1.53 //x2=27.685 //y2=1.22
cc_3344 ( N_noxref_11_c_4073_n N_CLK_c_5208_n ) capacitor c=0.0124075f \
 //x=27.24 //y=1.22 //x2=27.685 //y2=1.22
cc_3345 ( N_noxref_11_c_4071_n N_CLK_c_5094_n ) capacitor c=0.00103227f \
 //x=27.24 //y=0.875 //x2=28.21 //y2=0.91
cc_3346 ( N_noxref_11_c_4073_n N_CLK_c_5095_n ) capacitor c=0.0010154f \
 //x=27.24 //y=1.22 //x2=28.21 //y2=1.22
cc_3347 ( N_noxref_11_c_4073_n N_CLK_c_5096_n ) capacitor c=9.23422e-19 \
 //x=27.24 //y=1.22 //x2=28.21 //y2=1.45
cc_3348 ( N_noxref_11_c_4058_n N_CLK_c_5097_n ) capacitor c=0.00203769f \
 //x=27.01 //y=2.08 //x2=28.21 //y2=1.915
cc_3349 ( N_noxref_11_c_4068_n N_CLK_c_5097_n ) capacitor c=0.00834532f \
 //x=26.71 //y=1.915 //x2=28.21 //y2=1.915
cc_3350 ( N_noxref_11_c_4280_p N_CLK_c_5215_n ) capacitor c=0.00426767f \
 //x=41.26 //y=5.155 //x2=41.405 //y2=4.79
cc_3351 ( N_noxref_11_c_4058_n N_CLK_c_5101_n ) capacitor c=0.00183762f \
 //x=27.01 //y=2.08 //x2=28.12 //y2=4.7
cc_3352 ( N_noxref_11_c_4222_n N_CLK_c_5101_n ) capacitor c=0.0168581f \
 //x=27.575 //y=4.79 //x2=28.12 //y2=4.7
cc_3353 ( N_noxref_11_c_4118_n N_CLK_c_5101_n ) capacitor c=0.00484466f \
 //x=27.285 //y=4.79 //x2=28.12 //y2=4.7
cc_3354 ( N_noxref_11_c_4087_n N_CLK_c_5128_n ) capacitor c=0.00322046f \
 //x=41.175 //y=5.155 //x2=41.07 //y2=4.7
cc_3355 ( N_noxref_11_c_4058_n N_RN_c_5861_n ) capacitor c=0.0192695f \
 //x=27.01 //y=2.08 //x2=33.925 //y2=2.22
cc_3356 ( N_noxref_11_c_4068_n N_RN_c_5861_n ) capacitor c=0.011987f //x=26.71 \
 //y=1.915 //x2=33.925 //y2=2.22
cc_3357 ( N_noxref_11_c_4059_n N_RN_c_5873_n ) capacitor c=0.0178519f \
 //x=37.37 //y=2.08 //x2=42.065 //y2=2.22
cc_3358 ( N_noxref_11_c_4193_n N_RN_c_5873_n ) capacitor c=3.11115e-19 \
 //x=37.78 //y=1.405 //x2=42.065 //y2=2.22
cc_3359 ( N_noxref_11_c_4165_n N_RN_c_5873_n ) capacitor c=0.00570799f \
 //x=37.37 //y=2.08 //x2=42.065 //y2=2.22
cc_3360 ( N_noxref_11_c_4321_p N_RN_c_5882_n ) capacitor c=0.016327f //x=42.52 \
 //y=1.665 //x2=45.765 //y2=2.22
cc_3361 ( N_noxref_11_c_4101_n N_RN_c_5882_n ) capacitor c=0.0197307f \
 //x=42.92 //y=4.07 //x2=45.765 //y2=2.22
cc_3362 ( N_noxref_11_c_4101_n N_RN_c_5886_n ) capacitor c=0.0012045f \
 //x=42.92 //y=4.07 //x2=42.295 //y2=2.22
cc_3363 ( N_noxref_11_c_4062_n N_RN_c_5887_n ) capacitor c=0.0178519f \
 //x=50.32 //y=2.08 //x2=59.825 //y2=2.22
cc_3364 ( N_noxref_11_c_4325_p N_RN_c_5887_n ) capacitor c=3.11115e-19 \
 //x=50.73 //y=1.405 //x2=59.825 //y2=2.22
cc_3365 ( N_noxref_11_c_4247_n N_RN_c_5887_n ) capacitor c=0.00570799f \
 //x=50.32 //y=2.08 //x2=59.825 //y2=2.22
cc_3366 ( N_noxref_11_c_4075_n N_RN_c_5916_n ) capacitor c=0.0179722f \
 //x=37.255 //y=4.07 //x2=34.04 //y2=2.08
cc_3367 ( N_noxref_11_c_4078_n N_RN_c_5917_n ) capacitor c=0.0179722f \
 //x=42.805 //y=4.07 //x2=42.18 //y2=2.08
cc_3368 ( N_noxref_11_c_4081_n N_RN_c_5917_n ) capacitor c=0.00179385f \
 //x=43.035 //y=4.07 //x2=42.18 //y2=2.08
cc_3369 ( N_noxref_11_c_4101_n N_RN_c_5917_n ) capacitor c=0.0776213f \
 //x=42.92 //y=4.07 //x2=42.18 //y2=2.08
cc_3370 ( N_noxref_11_c_4331_p N_RN_c_5917_n ) capacitor c=0.0171303f \
 //x=42.14 //y=5.155 //x2=42.18 //y2=2.08
cc_3371 ( N_noxref_11_c_4079_n N_RN_c_5918_n ) capacitor c=0.0228716f \
 //x=50.205 //y=4.07 //x2=45.88 //y2=2.08
cc_3372 ( N_noxref_11_c_4101_n N_RN_c_5918_n ) capacitor c=6.36276e-19 \
 //x=42.92 //y=4.07 //x2=45.88 //y2=2.08
cc_3373 ( N_noxref_11_c_4093_n N_RN_M106_noxref_g ) capacitor c=0.01736f \
 //x=42.055 //y=5.155 //x2=41.92 //y2=6.02
cc_3374 ( N_noxref_11_M106_noxref_d N_RN_M106_noxref_g ) capacitor \
 c=0.0180032f //x=41.995 //y=5.02 //x2=41.92 //y2=6.02
cc_3375 ( N_noxref_11_c_4097_n N_RN_M107_noxref_g ) capacitor c=0.0194981f \
 //x=42.835 //y=5.155 //x2=42.36 //y2=6.02
cc_3376 ( N_noxref_11_M106_noxref_d N_RN_M107_noxref_g ) capacitor \
 c=0.0194246f //x=41.995 //y=5.02 //x2=42.36 //y2=6.02
cc_3377 ( N_noxref_11_M26_noxref_d N_RN_c_6196_n ) capacitor c=0.00217566f \
 //x=42.245 //y=0.915 //x2=42.17 //y2=0.915
cc_3378 ( N_noxref_11_M26_noxref_d N_RN_c_6197_n ) capacitor c=0.0034598f \
 //x=42.245 //y=0.915 //x2=42.17 //y2=1.26
cc_3379 ( N_noxref_11_M26_noxref_d N_RN_c_6198_n ) capacitor c=0.00546784f \
 //x=42.245 //y=0.915 //x2=42.17 //y2=1.57
cc_3380 ( N_noxref_11_M26_noxref_d N_RN_c_6199_n ) capacitor c=0.00241102f \
 //x=42.245 //y=0.915 //x2=42.545 //y2=0.76
cc_3381 ( N_noxref_11_c_4061_n N_RN_c_6200_n ) capacitor c=0.00371277f \
 //x=42.835 //y=1.665 //x2=42.545 //y2=1.415
cc_3382 ( N_noxref_11_M26_noxref_d N_RN_c_6200_n ) capacitor c=0.0138621f \
 //x=42.245 //y=0.915 //x2=42.545 //y2=1.415
cc_3383 ( N_noxref_11_M26_noxref_d N_RN_c_6202_n ) capacitor c=0.00219619f \
 //x=42.245 //y=0.915 //x2=42.7 //y2=0.915
cc_3384 ( N_noxref_11_c_4061_n N_RN_c_6203_n ) capacitor c=0.00457401f \
 //x=42.835 //y=1.665 //x2=42.7 //y2=1.26
cc_3385 ( N_noxref_11_M26_noxref_d N_RN_c_6203_n ) capacitor c=0.00603828f \
 //x=42.245 //y=0.915 //x2=42.7 //y2=1.26
cc_3386 ( N_noxref_11_c_4101_n N_RN_c_6205_n ) capacitor c=0.00709342f \
 //x=42.92 //y=4.07 //x2=42.18 //y2=2.08
cc_3387 ( N_noxref_11_c_4101_n N_RN_c_6206_n ) capacitor c=0.00283672f \
 //x=42.92 //y=4.07 //x2=42.18 //y2=1.915
cc_3388 ( N_noxref_11_M26_noxref_d N_RN_c_6206_n ) capacitor c=0.00661782f \
 //x=42.245 //y=0.915 //x2=42.18 //y2=1.915
cc_3389 ( N_noxref_11_c_4097_n N_RN_c_6208_n ) capacitor c=0.00201851f \
 //x=42.835 //y=5.155 //x2=42.18 //y2=4.7
cc_3390 ( N_noxref_11_c_4101_n N_RN_c_6208_n ) capacitor c=0.013693f //x=42.92 \
 //y=4.07 //x2=42.18 //y2=4.7
cc_3391 ( N_noxref_11_c_4331_p N_RN_c_6208_n ) capacitor c=0.00475601f \
 //x=42.14 //y=5.155 //x2=42.18 //y2=4.7
cc_3392 ( N_noxref_11_c_4079_n N_noxref_16_c_6833_n ) capacitor c=0.00649178f \
 //x=50.205 //y=4.07 //x2=53.025 //y2=4.07
cc_3393 ( N_noxref_11_c_4062_n N_noxref_16_c_6801_n ) capacitor c=8.49059e-19 \
 //x=50.32 //y=2.08 //x2=52.91 //y2=2.08
cc_3394 ( N_noxref_11_c_4079_n N_noxref_17_c_7491_n ) capacitor c=0.0661065f \
 //x=50.205 //y=4.07 //x2=50.945 //y2=3.33
cc_3395 ( N_noxref_11_c_4062_n N_noxref_17_c_7491_n ) capacitor c=0.019633f \
 //x=50.32 //y=2.08 //x2=50.945 //y2=3.33
cc_3396 ( N_noxref_11_c_4079_n N_noxref_17_c_7495_n ) capacitor c=0.0135672f \
 //x=50.205 //y=4.07 //x2=47.105 //y2=3.33
cc_3397 ( N_noxref_11_c_4062_n N_noxref_17_c_7529_n ) capacitor c=0.00117715f \
 //x=50.32 //y=2.08 //x2=51.175 //y2=3.33
cc_3398 ( N_noxref_11_c_4079_n N_noxref_17_c_7301_n ) capacitor c=0.0206302f \
 //x=50.205 //y=4.07 //x2=46.99 //y2=2.08
cc_3399 ( N_noxref_11_c_4228_n N_noxref_17_c_7373_n ) capacitor c=0.0127164f \
 //x=50.32 //y=4.535 //x2=50.495 //y2=5.2
cc_3400 ( N_noxref_11_M116_noxref_g N_noxref_17_c_7373_n ) capacitor \
 c=0.0166421f //x=50.36 //y=6.02 //x2=50.495 //y2=5.2
cc_3401 ( N_noxref_11_c_4249_n N_noxref_17_c_7373_n ) capacitor c=0.00346527f \
 //x=50.35 //y=4.7 //x2=50.495 //y2=5.2
cc_3402 ( N_noxref_11_M117_noxref_g N_noxref_17_c_7379_n ) capacitor \
 c=0.018922f //x=50.8 //y=6.02 //x2=50.975 //y2=5.2
cc_3403 ( N_noxref_11_c_4325_p N_noxref_17_c_7302_n ) capacitor c=0.00371277f \
 //x=50.73 //y=1.405 //x2=50.975 //y2=1.655
cc_3404 ( N_noxref_11_c_4246_n N_noxref_17_c_7302_n ) capacitor c=0.00457401f \
 //x=50.885 //y=1.25 //x2=50.975 //y2=1.655
cc_3405 ( N_noxref_11_c_4079_n N_noxref_17_c_7303_n ) capacitor c=0.00423741f \
 //x=50.205 //y=4.07 //x2=51.06 //y2=3.33
cc_3406 ( N_noxref_11_c_4228_n N_noxref_17_c_7303_n ) capacitor c=0.0101115f \
 //x=50.32 //y=4.535 //x2=51.06 //y2=3.33
cc_3407 ( N_noxref_11_c_4062_n N_noxref_17_c_7303_n ) capacitor c=0.0693397f \
 //x=50.32 //y=2.08 //x2=51.06 //y2=3.33
cc_3408 ( N_noxref_11_c_4281_p N_noxref_17_c_7303_n ) capacitor c=0.0142673f \
 //x=50.725 //y=4.79 //x2=51.06 //y2=3.33
cc_3409 ( N_noxref_11_c_4247_n N_noxref_17_c_7303_n ) capacitor c=0.00731987f \
 //x=50.32 //y=2.08 //x2=51.06 //y2=3.33
cc_3410 ( N_noxref_11_c_4371_p N_noxref_17_c_7303_n ) capacitor c=0.00306024f \
 //x=50.32 //y=1.915 //x2=51.06 //y2=3.33
cc_3411 ( N_noxref_11_c_4249_n N_noxref_17_c_7303_n ) capacitor c=0.00517969f \
 //x=50.35 //y=4.7 //x2=51.06 //y2=3.33
cc_3412 ( N_noxref_11_c_4281_p N_noxref_17_c_7544_n ) capacitor c=0.00407665f \
 //x=50.725 //y=4.79 //x2=50.58 //y2=5.2
cc_3413 ( N_noxref_11_c_4237_n N_noxref_17_M31_noxref_d ) capacitor \
 c=0.00217566f //x=50.355 //y=0.905 //x2=50.43 //y2=0.905
cc_3414 ( N_noxref_11_c_4240_n N_noxref_17_M31_noxref_d ) capacitor \
 c=0.0034598f //x=50.355 //y=1.25 //x2=50.43 //y2=0.905
cc_3415 ( N_noxref_11_c_4242_n N_noxref_17_M31_noxref_d ) capacitor \
 c=0.0066953f //x=50.355 //y=1.56 //x2=50.43 //y2=0.905
cc_3416 ( N_noxref_11_c_4377_p N_noxref_17_M31_noxref_d ) capacitor \
 c=0.00241102f //x=50.73 //y=0.75 //x2=50.43 //y2=0.905
cc_3417 ( N_noxref_11_c_4325_p N_noxref_17_M31_noxref_d ) capacitor \
 c=0.0137169f //x=50.73 //y=1.405 //x2=50.43 //y2=0.905
cc_3418 ( N_noxref_11_c_4245_n N_noxref_17_M31_noxref_d ) capacitor \
 c=0.00132245f //x=50.885 //y=0.905 //x2=50.43 //y2=0.905
cc_3419 ( N_noxref_11_c_4246_n N_noxref_17_M31_noxref_d ) capacitor \
 c=0.00566463f //x=50.885 //y=1.25 //x2=50.43 //y2=0.905
cc_3420 ( N_noxref_11_c_4371_p N_noxref_17_M31_noxref_d ) capacitor \
 c=0.00660593f //x=50.32 //y=1.915 //x2=50.43 //y2=0.905
cc_3421 ( N_noxref_11_M116_noxref_g N_noxref_17_M116_noxref_d ) capacitor \
 c=0.0173476f //x=50.36 //y=6.02 //x2=50.435 //y2=5.02
cc_3422 ( N_noxref_11_M117_noxref_g N_noxref_17_M116_noxref_d ) capacitor \
 c=0.0179769f //x=50.8 //y=6.02 //x2=50.435 //y2=5.02
cc_3423 ( N_noxref_11_c_4075_n N_noxref_20_c_8516_n ) capacitor c=0.0615741f \
 //x=37.255 //y=4.07 //x2=83.505 //y2=2.96
cc_3424 ( N_noxref_11_c_4077_n N_noxref_20_c_8516_n ) capacitor c=0.00776275f \
 //x=27.125 //y=4.07 //x2=83.505 //y2=2.96
cc_3425 ( N_noxref_11_c_4078_n N_noxref_20_c_8516_n ) capacitor c=0.0212588f \
 //x=42.805 //y=4.07 //x2=83.505 //y2=2.96
cc_3426 ( N_noxref_11_c_4144_n N_noxref_20_c_8516_n ) capacitor c=3.56521e-19 \
 //x=37.485 //y=4.07 //x2=83.505 //y2=2.96
cc_3427 ( N_noxref_11_c_4079_n N_noxref_20_c_8516_n ) capacitor c=0.0690095f \
 //x=50.205 //y=4.07 //x2=83.505 //y2=2.96
cc_3428 ( N_noxref_11_c_4081_n N_noxref_20_c_8516_n ) capacitor c=3.54204e-19 \
 //x=43.035 //y=4.07 //x2=83.505 //y2=2.96
cc_3429 ( N_noxref_11_c_4058_n N_noxref_20_c_8516_n ) capacitor c=0.0237066f \
 //x=27.01 //y=2.08 //x2=83.505 //y2=2.96
cc_3430 ( N_noxref_11_c_4059_n N_noxref_20_c_8516_n ) capacitor c=0.019291f \
 //x=37.37 //y=2.08 //x2=83.505 //y2=2.96
cc_3431 ( N_noxref_11_c_4101_n N_noxref_20_c_8516_n ) capacitor c=0.0210801f \
 //x=42.92 //y=4.07 //x2=83.505 //y2=2.96
cc_3432 ( N_noxref_11_c_4062_n N_noxref_20_c_8516_n ) capacitor c=0.0169513f \
 //x=50.32 //y=2.08 //x2=83.505 //y2=2.96
cc_3433 ( N_noxref_11_c_4058_n N_noxref_20_c_8608_n ) capacitor c=7.01366e-19 \
 //x=27.01 //y=2.08 //x2=25.275 //y2=2.96
cc_3434 ( N_noxref_11_c_4077_n N_noxref_20_c_8540_n ) capacitor c=0.00103915f \
 //x=27.125 //y=4.07 //x2=25.16 //y2=2.96
cc_3435 ( N_noxref_11_c_4058_n N_noxref_20_c_8540_n ) capacitor c=0.0148922f \
 //x=27.01 //y=2.08 //x2=25.16 //y2=2.96
cc_3436 ( N_noxref_11_c_4068_n N_noxref_33_c_9793_n ) capacitor c=0.0034165f \
 //x=26.71 //y=1.915 //x2=26.49 //y2=1.505
cc_3437 ( N_noxref_11_c_4058_n N_noxref_33_c_9777_n ) capacitor c=0.0115578f \
 //x=27.01 //y=2.08 //x2=27.375 //y2=1.59
cc_3438 ( N_noxref_11_c_4067_n N_noxref_33_c_9777_n ) capacitor c=0.00697148f \
 //x=26.71 //y=1.53 //x2=27.375 //y2=1.59
cc_3439 ( N_noxref_11_c_4068_n N_noxref_33_c_9777_n ) capacitor c=0.0204849f \
 //x=26.71 //y=1.915 //x2=27.375 //y2=1.59
cc_3440 ( N_noxref_11_c_4070_n N_noxref_33_c_9777_n ) capacitor c=0.00610316f \
 //x=27.085 //y=1.375 //x2=27.375 //y2=1.59
cc_3441 ( N_noxref_11_c_4073_n N_noxref_33_c_9777_n ) capacitor c=0.00698822f \
 //x=27.24 //y=1.22 //x2=27.375 //y2=1.59
cc_3442 ( N_noxref_11_c_4064_n N_noxref_33_M16_noxref_s ) capacitor \
 c=0.0327271f //x=26.71 //y=0.875 //x2=26.355 //y2=0.375
cc_3443 ( N_noxref_11_c_4067_n N_noxref_33_M16_noxref_s ) capacitor \
 c=7.99997e-19 //x=26.71 //y=1.53 //x2=26.355 //y2=0.375
cc_3444 ( N_noxref_11_c_4068_n N_noxref_33_M16_noxref_s ) capacitor \
 c=0.00122123f //x=26.71 //y=1.915 //x2=26.355 //y2=0.375
cc_3445 ( N_noxref_11_c_4071_n N_noxref_33_M16_noxref_s ) capacitor \
 c=0.0121427f //x=27.24 //y=0.875 //x2=26.355 //y2=0.375
cc_3446 ( N_noxref_11_c_4160_n N_noxref_37_c_9987_n ) capacitor c=0.00623646f \
 //x=37.405 //y=1.56 //x2=37.185 //y2=1.495
cc_3447 ( N_noxref_11_c_4165_n N_noxref_37_c_9987_n ) capacitor c=0.00173579f \
 //x=37.37 //y=2.08 //x2=37.185 //y2=1.495
cc_3448 ( N_noxref_11_c_4059_n N_noxref_37_c_9988_n ) capacitor c=0.00156605f \
 //x=37.37 //y=2.08 //x2=38.07 //y2=0.53
cc_3449 ( N_noxref_11_c_4155_n N_noxref_37_c_9988_n ) capacitor c=0.0188655f \
 //x=37.405 //y=0.905 //x2=38.07 //y2=0.53
cc_3450 ( N_noxref_11_c_4163_n N_noxref_37_c_9988_n ) capacitor c=0.00656458f \
 //x=37.935 //y=0.905 //x2=38.07 //y2=0.53
cc_3451 ( N_noxref_11_c_4165_n N_noxref_37_c_9988_n ) capacitor c=2.1838e-19 \
 //x=37.37 //y=2.08 //x2=38.07 //y2=0.53
cc_3452 ( N_noxref_11_c_4155_n N_noxref_37_M22_noxref_s ) capacitor \
 c=0.00623646f //x=37.405 //y=0.905 //x2=36.08 //y2=0.365
cc_3453 ( N_noxref_11_c_4163_n N_noxref_37_M22_noxref_s ) capacitor \
 c=0.0143002f //x=37.935 //y=0.905 //x2=36.08 //y2=0.365
cc_3454 ( N_noxref_11_c_4164_n N_noxref_37_M22_noxref_s ) capacitor \
 c=0.00290153f //x=37.935 //y=1.25 //x2=36.08 //y2=0.365
cc_3455 ( N_noxref_11_M26_noxref_d N_noxref_38_M24_noxref_s ) capacitor \
 c=0.00309936f //x=42.245 //y=0.915 //x2=39.305 //y2=0.375
cc_3456 ( N_noxref_11_c_4061_n N_noxref_39_c_10085_n ) capacitor c=0.00457167f \
 //x=42.835 //y=1.665 //x2=42.835 //y2=0.54
cc_3457 ( N_noxref_11_M26_noxref_d N_noxref_39_c_10085_n ) capacitor \
 c=0.0115903f //x=42.245 //y=0.915 //x2=42.835 //y2=0.54
cc_3458 ( N_noxref_11_c_4321_p N_noxref_39_c_10095_n ) capacitor c=0.0200405f \
 //x=42.52 //y=1.665 //x2=41.95 //y2=0.995
cc_3459 ( N_noxref_11_M26_noxref_d N_noxref_39_M25_noxref_d ) capacitor \
 c=5.27807e-19 //x=42.245 //y=0.915 //x2=40.71 //y2=0.91
cc_3460 ( N_noxref_11_c_4061_n N_noxref_39_M26_noxref_s ) capacitor \
 c=0.0196084f //x=42.835 //y=1.665 //x2=41.815 //y2=0.375
cc_3461 ( N_noxref_11_M26_noxref_d N_noxref_39_M26_noxref_s ) capacitor \
 c=0.0426368f //x=42.245 //y=0.915 //x2=41.815 //y2=0.375
cc_3462 ( N_noxref_11_c_4061_n N_noxref_40_c_10148_n ) capacitor c=3.84569e-19 \
 //x=42.835 //y=1.665 //x2=44.25 //y2=1.505
cc_3463 ( N_noxref_11_M26_noxref_d N_noxref_40_M27_noxref_s ) capacitor \
 c=2.55333e-19 //x=42.245 //y=0.915 //x2=44.115 //y2=0.375
cc_3464 ( N_noxref_11_c_4242_n N_noxref_42_c_10244_n ) capacitor c=0.00623646f \
 //x=50.355 //y=1.56 //x2=50.135 //y2=1.495
cc_3465 ( N_noxref_11_c_4247_n N_noxref_42_c_10244_n ) capacitor c=0.00173579f \
 //x=50.32 //y=2.08 //x2=50.135 //y2=1.495
cc_3466 ( N_noxref_11_c_4062_n N_noxref_42_c_10245_n ) capacitor c=0.00156605f \
 //x=50.32 //y=2.08 //x2=51.02 //y2=0.53
cc_3467 ( N_noxref_11_c_4237_n N_noxref_42_c_10245_n ) capacitor c=0.0188655f \
 //x=50.355 //y=0.905 //x2=51.02 //y2=0.53
cc_3468 ( N_noxref_11_c_4245_n N_noxref_42_c_10245_n ) capacitor c=0.00656458f \
 //x=50.885 //y=0.905 //x2=51.02 //y2=0.53
cc_3469 ( N_noxref_11_c_4247_n N_noxref_42_c_10245_n ) capacitor c=2.1838e-19 \
 //x=50.32 //y=2.08 //x2=51.02 //y2=0.53
cc_3470 ( N_noxref_11_c_4237_n N_noxref_42_M30_noxref_s ) capacitor \
 c=0.00623646f //x=50.355 //y=0.905 //x2=49.03 //y2=0.365
cc_3471 ( N_noxref_11_c_4245_n N_noxref_42_M30_noxref_s ) capacitor \
 c=0.0143002f //x=50.885 //y=0.905 //x2=49.03 //y2=0.365
cc_3472 ( N_noxref_11_c_4246_n N_noxref_42_M30_noxref_s ) capacitor \
 c=0.00290153f //x=50.885 //y=1.25 //x2=49.03 //y2=0.365
cc_3473 ( N_D_c_4448_n N_CLK_c_4808_n ) capacitor c=0.0210462f //x=7.03 \
 //y=2.08 //x2=15.055 //y2=4.44
cc_3474 ( N_D_c_4482_n N_CLK_c_4808_n ) capacitor c=0.0085986f //x=7.365 \
 //y=4.79 //x2=15.055 //y2=4.44
cc_3475 ( N_D_c_4483_n N_CLK_c_4808_n ) capacitor c=0.00293313f //x=7.03 \
 //y=4.7 //x2=15.055 //y2=4.44
cc_3476 ( N_D_c_4434_n N_CLK_c_4826_n ) capacitor c=0.0185184f //x=32.815 \
 //y=2.59 //x2=28.005 //y2=4.44
cc_3477 ( N_D_c_4449_n N_CLK_c_4844_n ) capacitor c=0.0210462f //x=32.93 \
 //y=2.08 //x2=40.955 //y2=4.44
cc_3478 ( N_D_c_4546_n N_CLK_c_4844_n ) capacitor c=0.0085986f //x=33.265 \
 //y=4.79 //x2=40.955 //y2=4.44
cc_3479 ( N_D_c_4547_n N_CLK_c_4844_n ) capacitor c=0.00293313f //x=32.93 \
 //y=4.7 //x2=40.955 //y2=4.44
cc_3480 ( N_D_c_4450_n N_CLK_c_4880_n ) capacitor c=0.0210462f //x=58.83 \
 //y=2.08 //x2=66.855 //y2=4.44
cc_3481 ( N_D_c_4598_p N_CLK_c_4880_n ) capacitor c=0.00862724f //x=59.165 \
 //y=4.79 //x2=66.855 //y2=4.44
cc_3482 ( N_D_c_4599_p N_CLK_c_4880_n ) capacitor c=0.00293313f //x=58.83 \
 //y=4.7 //x2=66.855 //y2=4.44
cc_3483 ( N_D_c_4434_n N_CLK_c_4803_n ) capacitor c=0.0228599f //x=32.815 \
 //y=2.59 //x2=15.17 //y2=2.08
cc_3484 ( N_D_c_4434_n N_CLK_c_4804_n ) capacitor c=0.0190006f //x=32.815 \
 //y=2.59 //x2=28.12 //y2=2.08
cc_3485 ( N_D_c_4442_n N_CLK_c_4805_n ) capacitor c=0.0190006f //x=58.715 \
 //y=2.59 //x2=41.07 //y2=2.08
cc_3486 ( N_D_c_4442_n N_CLK_c_4806_n ) capacitor c=0.0190006f //x=58.715 \
 //y=2.59 //x2=54.02 //y2=2.08
cc_3487 ( N_D_c_4450_n N_noxref_14_c_5659_n ) capacitor c=0.0190398f //x=58.83 \
 //y=2.08 //x2=70.555 //y2=3.7
cc_3488 ( N_D_c_4450_n N_noxref_14_c_5660_n ) capacitor c=9.95819e-19 \
 //x=58.83 //y=2.08 //x2=57.835 //y2=3.7
cc_3489 ( N_D_c_4442_n N_noxref_14_c_5625_n ) capacitor c=0.0165903f \
 //x=58.715 //y=2.59 //x2=55.87 //y2=3.7
cc_3490 ( N_D_c_4450_n N_noxref_14_c_5625_n ) capacitor c=3.3533e-19 //x=58.83 \
 //y=2.08 //x2=55.87 //y2=3.7
cc_3491 ( N_D_c_4442_n N_noxref_14_c_5588_n ) capacitor c=0.0201108f \
 //x=58.715 //y=2.59 //x2=57.72 //y2=2.08
cc_3492 ( N_D_c_4450_n N_noxref_14_c_5588_n ) capacitor c=0.0413373f //x=58.83 \
 //y=2.08 //x2=57.72 //y2=2.08
cc_3493 ( N_D_c_4610_p N_noxref_14_c_5588_n ) capacitor c=0.00203769f \
 //x=58.92 //y=1.915 //x2=57.72 //y2=2.08
cc_3494 ( N_D_c_4599_p N_noxref_14_c_5588_n ) capacitor c=0.00183762f \
 //x=58.83 //y=4.7 //x2=57.72 //y2=2.08
cc_3495 ( N_D_M126_noxref_g N_noxref_14_M124_noxref_g ) capacitor c=0.0105869f \
 //x=58.8 //y=6.02 //x2=57.92 //y2=6.02
cc_3496 ( N_D_M126_noxref_g N_noxref_14_M125_noxref_g ) capacitor c=0.10632f \
 //x=58.8 //y=6.02 //x2=58.36 //y2=6.02
cc_3497 ( N_D_M127_noxref_g N_noxref_14_M125_noxref_g ) capacitor c=0.0101598f \
 //x=59.24 //y=6.02 //x2=58.36 //y2=6.02
cc_3498 ( N_D_c_4615_p N_noxref_14_c_5590_n ) capacitor c=5.72482e-19 \
 //x=58.395 //y=0.91 //x2=57.42 //y2=0.875
cc_3499 ( N_D_c_4615_p N_noxref_14_c_5592_n ) capacitor c=0.00149976f \
 //x=58.395 //y=0.91 //x2=57.42 //y2=1.22
cc_3500 ( N_D_c_4617_p N_noxref_14_c_5593_n ) capacitor c=0.00111227f \
 //x=58.395 //y=1.22 //x2=57.42 //y2=1.53
cc_3501 ( N_D_c_4450_n N_noxref_14_c_5594_n ) capacitor c=0.00210802f \
 //x=58.83 //y=2.08 //x2=57.42 //y2=1.915
cc_3502 ( N_D_c_4610_p N_noxref_14_c_5594_n ) capacitor c=0.00834532f \
 //x=58.92 //y=1.915 //x2=57.42 //y2=1.915
cc_3503 ( N_D_c_4615_p N_noxref_14_c_5597_n ) capacitor c=0.0160123f \
 //x=58.395 //y=0.91 //x2=57.95 //y2=0.875
cc_3504 ( N_D_c_4621_p N_noxref_14_c_5597_n ) capacitor c=0.00103227f \
 //x=58.92 //y=0.91 //x2=57.95 //y2=0.875
cc_3505 ( N_D_c_4617_p N_noxref_14_c_5599_n ) capacitor c=0.0124075f \
 //x=58.395 //y=1.22 //x2=57.95 //y2=1.22
cc_3506 ( N_D_c_4623_p N_noxref_14_c_5599_n ) capacitor c=0.0010154f //x=58.92 \
 //y=1.22 //x2=57.95 //y2=1.22
cc_3507 ( N_D_c_4624_p N_noxref_14_c_5599_n ) capacitor c=9.23422e-19 \
 //x=58.92 //y=1.45 //x2=57.95 //y2=1.22
cc_3508 ( N_D_c_4450_n N_noxref_14_c_5680_n ) capacitor c=0.00147352f \
 //x=58.83 //y=2.08 //x2=58.285 //y2=4.79
cc_3509 ( N_D_c_4599_p N_noxref_14_c_5680_n ) capacitor c=0.0168581f //x=58.83 \
 //y=4.7 //x2=58.285 //y2=4.79
cc_3510 ( N_D_c_4450_n N_noxref_14_c_5640_n ) capacitor c=0.00142741f \
 //x=58.83 //y=2.08 //x2=57.995 //y2=4.79
cc_3511 ( N_D_c_4599_p N_noxref_14_c_5640_n ) capacitor c=0.00484466f \
 //x=58.83 //y=4.7 //x2=57.995 //y2=4.79
cc_3512 ( N_D_c_4434_n N_RN_c_5846_n ) capacitor c=0.688138f //x=32.815 \
 //y=2.59 //x2=16.165 //y2=2.22
cc_3513 ( N_D_c_4434_n N_RN_c_5854_n ) capacitor c=0.029141f //x=32.815 \
 //y=2.59 //x2=8.255 //y2=2.22
cc_3514 ( N_D_c_4448_n N_RN_c_5854_n ) capacitor c=0.00558344f //x=7.03 \
 //y=2.08 //x2=8.255 //y2=2.22
cc_3515 ( N_D_c_4510_n N_RN_c_5854_n ) capacitor c=0.00341397f //x=7.12 \
 //y=1.915 //x2=8.255 //y2=2.22
cc_3516 ( N_D_c_4434_n N_RN_c_5856_n ) capacitor c=0.302834f //x=32.815 \
 //y=2.59 //x2=19.865 //y2=2.22
cc_3517 ( N_D_c_4434_n N_RN_c_5860_n ) capacitor c=0.026528f //x=32.815 \
 //y=2.59 //x2=16.395 //y2=2.22
cc_3518 ( N_D_c_4434_n N_RN_c_5861_n ) capacitor c=1.10611f //x=32.815 \
 //y=2.59 //x2=33.925 //y2=2.22
cc_3519 ( N_D_c_4442_n N_RN_c_5861_n ) capacitor c=0.0764156f //x=58.715 \
 //y=2.59 //x2=33.925 //y2=2.22
cc_3520 ( N_D_c_4538_n N_RN_c_5861_n ) capacitor c=0.0263455f //x=33.045 \
 //y=2.59 //x2=33.925 //y2=2.22
cc_3521 ( N_D_c_4449_n N_RN_c_5861_n ) capacitor c=0.021223f //x=32.93 \
 //y=2.08 //x2=33.925 //y2=2.22
cc_3522 ( N_D_c_4575_n N_RN_c_5861_n ) capacitor c=0.00583058f //x=33.02 \
 //y=1.915 //x2=33.925 //y2=2.22
cc_3523 ( N_D_c_4434_n N_RN_c_5872_n ) capacitor c=0.0265257f //x=32.815 \
 //y=2.59 //x2=20.095 //y2=2.22
cc_3524 ( N_D_c_4442_n N_RN_c_5873_n ) capacitor c=0.688138f //x=58.715 \
 //y=2.59 //x2=42.065 //y2=2.22
cc_3525 ( N_D_c_4442_n N_RN_c_5881_n ) capacitor c=0.026528f //x=58.715 \
 //y=2.59 //x2=34.155 //y2=2.22
cc_3526 ( N_D_c_4449_n N_RN_c_5881_n ) capacitor c=0.00165648f //x=32.93 \
 //y=2.08 //x2=34.155 //y2=2.22
cc_3527 ( N_D_c_4575_n N_RN_c_5881_n ) capacitor c=2.3323e-19 //x=33.02 \
 //y=1.915 //x2=34.155 //y2=2.22
cc_3528 ( N_D_c_4442_n N_RN_c_5882_n ) capacitor c=0.302834f //x=58.715 \
 //y=2.59 //x2=45.765 //y2=2.22
cc_3529 ( N_D_c_4442_n N_RN_c_5886_n ) capacitor c=0.026528f //x=58.715 \
 //y=2.59 //x2=42.295 //y2=2.22
cc_3530 ( N_D_c_4442_n N_RN_c_5887_n ) capacitor c=1.14541f //x=58.715 \
 //y=2.59 //x2=59.825 //y2=2.22
cc_3531 ( N_D_c_4450_n N_RN_c_5887_n ) capacitor c=0.021223f //x=58.83 \
 //y=2.08 //x2=59.825 //y2=2.22
cc_3532 ( N_D_c_4610_p N_RN_c_5887_n ) capacitor c=0.00583058f //x=58.92 \
 //y=1.915 //x2=59.825 //y2=2.22
cc_3533 ( N_D_c_4442_n N_RN_c_5898_n ) capacitor c=0.0265257f //x=58.715 \
 //y=2.59 //x2=45.995 //y2=2.22
cc_3534 ( N_D_c_4450_n N_RN_c_5907_n ) capacitor c=0.00165648f //x=58.83 \
 //y=2.08 //x2=60.055 //y2=2.22
cc_3535 ( N_D_c_4610_p N_RN_c_5907_n ) capacitor c=2.3323e-19 //x=58.92 \
 //y=1.915 //x2=60.055 //y2=2.22
cc_3536 ( N_D_c_4434_n N_RN_c_5913_n ) capacitor c=0.0221442f //x=32.815 \
 //y=2.59 //x2=8.14 //y2=2.08
cc_3537 ( N_D_c_4441_n N_RN_c_5913_n ) capacitor c=0.00128547f //x=7.145 \
 //y=2.59 //x2=8.14 //y2=2.08
cc_3538 ( N_D_c_4448_n N_RN_c_5913_n ) capacitor c=0.0443596f //x=7.03 \
 //y=2.08 //x2=8.14 //y2=2.08
cc_3539 ( N_D_c_4510_n N_RN_c_5913_n ) capacitor c=0.00223318f //x=7.12 \
 //y=1.915 //x2=8.14 //y2=2.08
cc_3540 ( N_D_c_4483_n N_RN_c_5913_n ) capacitor c=0.00142741f //x=7.03 \
 //y=4.7 //x2=8.14 //y2=2.08
cc_3541 ( N_D_c_4434_n N_RN_c_5914_n ) capacitor c=0.0236632f //x=32.815 \
 //y=2.59 //x2=16.28 //y2=2.08
cc_3542 ( N_D_c_4434_n N_RN_c_5915_n ) capacitor c=0.025687f //x=32.815 \
 //y=2.59 //x2=19.98 //y2=2.08
cc_3543 ( N_D_c_4442_n N_RN_c_5916_n ) capacitor c=0.0198038f //x=58.715 \
 //y=2.59 //x2=34.04 //y2=2.08
cc_3544 ( N_D_c_4538_n N_RN_c_5916_n ) capacitor c=0.00128547f //x=33.045 \
 //y=2.59 //x2=34.04 //y2=2.08
cc_3545 ( N_D_c_4449_n N_RN_c_5916_n ) capacitor c=0.0413732f //x=32.93 \
 //y=2.08 //x2=34.04 //y2=2.08
cc_3546 ( N_D_c_4575_n N_RN_c_5916_n ) capacitor c=0.00203728f //x=33.02 \
 //y=1.915 //x2=34.04 //y2=2.08
cc_3547 ( N_D_c_4547_n N_RN_c_5916_n ) capacitor c=0.00142741f //x=32.93 \
 //y=4.7 //x2=34.04 //y2=2.08
cc_3548 ( N_D_c_4442_n N_RN_c_5917_n ) capacitor c=0.0198038f //x=58.715 \
 //y=2.59 //x2=42.18 //y2=2.08
cc_3549 ( N_D_c_4442_n N_RN_c_5918_n ) capacitor c=0.0208419f //x=58.715 \
 //y=2.59 //x2=45.88 //y2=2.08
cc_3550 ( N_D_c_4442_n N_RN_c_5919_n ) capacitor c=0.00575746f //x=58.715 \
 //y=2.59 //x2=59.94 //y2=2.08
cc_3551 ( N_D_c_4450_n N_RN_c_5919_n ) capacitor c=0.0422177f //x=58.83 \
 //y=2.08 //x2=59.94 //y2=2.08
cc_3552 ( N_D_c_4610_p N_RN_c_5919_n ) capacitor c=0.00203728f //x=58.92 \
 //y=1.915 //x2=59.94 //y2=2.08
cc_3553 ( N_D_c_4599_p N_RN_c_5919_n ) capacitor c=0.00142741f //x=58.83 \
 //y=4.7 //x2=59.94 //y2=2.08
cc_3554 ( N_D_M62_noxref_g N_RN_M64_noxref_g ) capacitor c=0.0101598f //x=7 \
 //y=6.02 //x2=7.88 //y2=6.02
cc_3555 ( N_D_M63_noxref_g N_RN_M64_noxref_g ) capacitor c=0.0602553f //x=7.44 \
 //y=6.02 //x2=7.88 //y2=6.02
cc_3556 ( N_D_M63_noxref_g N_RN_M65_noxref_g ) capacitor c=0.0101598f //x=7.44 \
 //y=6.02 //x2=8.32 //y2=6.02
cc_3557 ( N_D_M94_noxref_g N_RN_M96_noxref_g ) capacitor c=0.0101598f //x=32.9 \
 //y=6.02 //x2=33.78 //y2=6.02
cc_3558 ( N_D_M95_noxref_g N_RN_M96_noxref_g ) capacitor c=0.0602553f \
 //x=33.34 //y=6.02 //x2=33.78 //y2=6.02
cc_3559 ( N_D_M95_noxref_g N_RN_M97_noxref_g ) capacitor c=0.0101598f \
 //x=33.34 //y=6.02 //x2=34.22 //y2=6.02
cc_3560 ( N_D_M126_noxref_g N_RN_M128_noxref_g ) capacitor c=0.0101598f \
 //x=58.8 //y=6.02 //x2=59.68 //y2=6.02
cc_3561 ( N_D_M127_noxref_g N_RN_M128_noxref_g ) capacitor c=0.0602553f \
 //x=59.24 //y=6.02 //x2=59.68 //y2=6.02
cc_3562 ( N_D_M127_noxref_g N_RN_M129_noxref_g ) capacitor c=0.0101598f \
 //x=59.24 //y=6.02 //x2=60.12 //y2=6.02
cc_3563 ( N_D_c_4507_n N_RN_c_5988_n ) capacitor c=0.00456962f //x=7.12 \
 //y=0.91 //x2=8.13 //y2=0.915
cc_3564 ( N_D_c_4508_n N_RN_c_5989_n ) capacitor c=0.00438372f //x=7.12 \
 //y=1.22 //x2=8.13 //y2=1.26
cc_3565 ( N_D_c_4509_n N_RN_c_5990_n ) capacitor c=0.00438372f //x=7.12 \
 //y=1.45 //x2=8.13 //y2=1.57
cc_3566 ( N_D_c_4572_n N_RN_c_6109_n ) capacitor c=0.00456962f //x=33.02 \
 //y=0.91 //x2=34.03 //y2=0.915
cc_3567 ( N_D_c_4573_n N_RN_c_6110_n ) capacitor c=0.00438372f //x=33.02 \
 //y=1.22 //x2=34.03 //y2=1.26
cc_3568 ( N_D_c_4574_n N_RN_c_6111_n ) capacitor c=0.00438372f //x=33.02 \
 //y=1.45 //x2=34.03 //y2=1.57
cc_3569 ( N_D_c_4621_p N_RN_c_6268_n ) capacitor c=0.00456962f //x=58.92 \
 //y=0.91 //x2=59.93 //y2=0.915
cc_3570 ( N_D_c_4623_p N_RN_c_6269_n ) capacitor c=0.00438372f //x=58.92 \
 //y=1.22 //x2=59.93 //y2=1.26
cc_3571 ( N_D_c_4624_p N_RN_c_6270_n ) capacitor c=0.00438372f //x=58.92 \
 //y=1.45 //x2=59.93 //y2=1.57
cc_3572 ( N_D_c_4448_n N_RN_c_5997_n ) capacitor c=0.00209043f //x=7.03 \
 //y=2.08 //x2=8.14 //y2=2.08
cc_3573 ( N_D_c_4510_n N_RN_c_5997_n ) capacitor c=0.00881982f //x=7.12 \
 //y=1.915 //x2=8.14 //y2=2.08
cc_3574 ( N_D_c_4510_n N_RN_c_5998_n ) capacitor c=0.00438372f //x=7.12 \
 //y=1.915 //x2=8.14 //y2=1.915
cc_3575 ( N_D_c_4448_n N_RN_c_6000_n ) capacitor c=0.00219458f //x=7.03 \
 //y=2.08 //x2=8.14 //y2=4.7
cc_3576 ( N_D_c_4482_n N_RN_c_6000_n ) capacitor c=0.0611812f //x=7.365 \
 //y=4.79 //x2=8.14 //y2=4.7
cc_3577 ( N_D_c_4483_n N_RN_c_6000_n ) capacitor c=0.00487508f //x=7.03 \
 //y=4.7 //x2=8.14 //y2=4.7
cc_3578 ( N_D_c_4449_n N_RN_c_6118_n ) capacitor c=0.00201097f //x=32.93 \
 //y=2.08 //x2=34.04 //y2=2.08
cc_3579 ( N_D_c_4575_n N_RN_c_6118_n ) capacitor c=0.00828003f //x=33.02 \
 //y=1.915 //x2=34.04 //y2=2.08
cc_3580 ( N_D_c_4575_n N_RN_c_6119_n ) capacitor c=0.00438372f //x=33.02 \
 //y=1.915 //x2=34.04 //y2=1.915
cc_3581 ( N_D_c_4449_n N_RN_c_6121_n ) capacitor c=0.00219458f //x=32.93 \
 //y=2.08 //x2=34.04 //y2=4.7
cc_3582 ( N_D_c_4546_n N_RN_c_6121_n ) capacitor c=0.0611812f //x=33.265 \
 //y=4.79 //x2=34.04 //y2=4.7
cc_3583 ( N_D_c_4547_n N_RN_c_6121_n ) capacitor c=0.00487508f //x=32.93 \
 //y=4.7 //x2=34.04 //y2=4.7
cc_3584 ( N_D_c_4450_n N_RN_c_6283_n ) capacitor c=0.00201097f //x=58.83 \
 //y=2.08 //x2=59.94 //y2=2.08
cc_3585 ( N_D_c_4610_p N_RN_c_6283_n ) capacitor c=0.00828003f //x=58.92 \
 //y=1.915 //x2=59.94 //y2=2.08
cc_3586 ( N_D_c_4610_p N_RN_c_6285_n ) capacitor c=0.00438372f //x=58.92 \
 //y=1.915 //x2=59.94 //y2=1.915
cc_3587 ( N_D_c_4450_n N_RN_c_6286_n ) capacitor c=0.00219458f //x=58.83 \
 //y=2.08 //x2=59.94 //y2=4.7
cc_3588 ( N_D_c_4598_p N_RN_c_6286_n ) capacitor c=0.0611812f //x=59.165 \
 //y=4.79 //x2=59.94 //y2=4.7
cc_3589 ( N_D_c_4599_p N_RN_c_6286_n ) capacitor c=0.00487508f //x=58.83 \
 //y=4.7 //x2=59.94 //y2=4.7
cc_3590 ( N_D_c_4450_n N_noxref_16_c_6831_n ) capacitor c=0.0190126f //x=58.83 \
 //y=2.08 //x2=63.155 //y2=4.07
cc_3591 ( N_D_c_4442_n N_noxref_16_c_6801_n ) capacitor c=0.0188253f \
 //x=58.715 //y=2.59 //x2=52.91 //y2=2.08
cc_3592 ( N_D_c_4442_n N_noxref_17_c_7491_n ) capacitor c=0.0295716f \
 //x=58.715 //y=2.59 //x2=50.945 //y2=3.33
cc_3593 ( N_D_c_4442_n N_noxref_17_c_7495_n ) capacitor c=9.8111e-19 \
 //x=58.715 //y=2.59 //x2=47.105 //y2=3.33
cc_3594 ( N_D_c_4442_n N_noxref_17_c_7362_n ) capacitor c=0.0302604f \
 //x=58.715 //y=2.59 //x2=55.015 //y2=3.33
cc_3595 ( N_D_c_4442_n N_noxref_17_c_7529_n ) capacitor c=5.75258e-19 \
 //x=58.715 //y=2.59 //x2=51.175 //y2=3.33
cc_3596 ( N_D_c_4442_n N_noxref_17_c_7559_n ) capacitor c=0.0284903f \
 //x=58.715 //y=2.59 //x2=60.565 //y2=3.33
cc_3597 ( N_D_c_4450_n N_noxref_17_c_7559_n ) capacitor c=0.0190562f //x=58.83 \
 //y=2.08 //x2=60.565 //y2=3.33
cc_3598 ( N_D_c_4442_n N_noxref_17_c_7561_n ) capacitor c=6.6144e-19 \
 //x=58.715 //y=2.59 //x2=55.245 //y2=3.33
cc_3599 ( N_D_c_4442_n N_noxref_17_c_7301_n ) capacitor c=0.0179628f \
 //x=58.715 //y=2.59 //x2=46.99 //y2=2.08
cc_3600 ( N_D_c_4442_n N_noxref_17_c_7303_n ) capacitor c=0.0165961f \
 //x=58.715 //y=2.59 //x2=51.06 //y2=3.33
cc_3601 ( N_D_c_4442_n N_noxref_17_c_7304_n ) capacitor c=0.0179628f \
 //x=58.715 //y=2.59 //x2=55.13 //y2=2.08
cc_3602 ( N_D_c_4450_n N_noxref_17_c_7385_n ) capacitor c=0.0146f //x=58.83 \
 //y=2.08 //x2=58.935 //y2=5.155
cc_3603 ( N_D_M126_noxref_g N_noxref_17_c_7385_n ) capacitor c=0.0165266f \
 //x=58.8 //y=6.02 //x2=58.935 //y2=5.155
cc_3604 ( N_D_c_4599_p N_noxref_17_c_7385_n ) capacitor c=0.00322054f \
 //x=58.83 //y=4.7 //x2=58.935 //y2=5.155
cc_3605 ( N_D_M127_noxref_g N_noxref_17_c_7391_n ) capacitor c=0.01736f \
 //x=59.24 //y=6.02 //x2=59.815 //y2=5.155
cc_3606 ( N_D_c_4450_n N_noxref_17_c_7399_n ) capacitor c=0.00252523f \
 //x=58.83 //y=2.08 //x2=60.68 //y2=3.33
cc_3607 ( N_D_c_4598_p N_noxref_17_c_7570_n ) capacitor c=0.00426767f \
 //x=59.165 //y=4.79 //x2=59.02 //y2=5.155
cc_3608 ( N_D_M126_noxref_g N_noxref_17_M126_noxref_d ) capacitor c=0.0180032f \
 //x=58.8 //y=6.02 //x2=58.875 //y2=5.02
cc_3609 ( N_D_M127_noxref_g N_noxref_17_M126_noxref_d ) capacitor c=0.0180032f \
 //x=59.24 //y=6.02 //x2=58.875 //y2=5.02
cc_3610 ( N_D_c_4434_n N_noxref_20_c_8515_n ) capacitor c=0.334584f //x=32.815 \
 //y=2.59 //x2=25.045 //y2=2.96
cc_3611 ( N_D_c_4434_n N_noxref_20_c_8606_n ) capacitor c=0.0290442f \
 //x=32.815 //y=2.59 //x2=21.205 //y2=2.96
cc_3612 ( N_D_c_4434_n N_noxref_20_c_8516_n ) capacitor c=0.659576f //x=32.815 \
 //y=2.59 //x2=83.505 //y2=2.96
cc_3613 ( N_D_c_4442_n N_noxref_20_c_8516_n ) capacitor c=2.2789f //x=58.715 \
 //y=2.59 //x2=83.505 //y2=2.96
cc_3614 ( N_D_c_4538_n N_noxref_20_c_8516_n ) capacitor c=0.0265456f \
 //x=33.045 //y=2.59 //x2=83.505 //y2=2.96
cc_3615 ( N_D_c_4449_n N_noxref_20_c_8516_n ) capacitor c=0.0208701f //x=32.93 \
 //y=2.08 //x2=83.505 //y2=2.96
cc_3616 ( N_D_c_4450_n N_noxref_20_c_8516_n ) capacitor c=0.0208701f //x=58.83 \
 //y=2.08 //x2=83.505 //y2=2.96
cc_3617 ( N_D_c_4434_n N_noxref_20_c_8608_n ) capacitor c=0.0265752f \
 //x=32.815 //y=2.59 //x2=25.275 //y2=2.96
cc_3618 ( N_D_c_4434_n N_noxref_20_c_8538_n ) capacitor c=0.0197974f \
 //x=32.815 //y=2.59 //x2=21.09 //y2=2.08
cc_3619 ( N_D_c_4434_n N_noxref_20_c_8540_n ) capacitor c=0.0184306f \
 //x=32.815 //y=2.59 //x2=25.16 //y2=2.96
cc_3620 ( N_D_c_4502_n N_noxref_25_c_9371_n ) capacitor c=0.0167228f //x=6.595 \
 //y=0.91 //x2=7.255 //y2=0.54
cc_3621 ( N_D_c_4507_n N_noxref_25_c_9371_n ) capacitor c=0.00534519f //x=7.12 \
 //y=0.91 //x2=7.255 //y2=0.54
cc_3622 ( N_D_c_4434_n N_noxref_25_c_9381_n ) capacitor c=0.0029635f \
 //x=32.815 //y=2.59 //x2=7.255 //y2=1.59
cc_3623 ( N_D_c_4441_n N_noxref_25_c_9381_n ) capacitor c=0.00236045f \
 //x=7.145 //y=2.59 //x2=7.255 //y2=1.59
cc_3624 ( N_D_c_4448_n N_noxref_25_c_9381_n ) capacitor c=0.0120444f //x=7.03 \
 //y=2.08 //x2=7.255 //y2=1.59
cc_3625 ( N_D_c_4505_n N_noxref_25_c_9381_n ) capacitor c=0.0153476f //x=6.595 \
 //y=1.22 //x2=7.255 //y2=1.59
cc_3626 ( N_D_c_4510_n N_noxref_25_c_9381_n ) capacitor c=0.0219169f //x=7.12 \
 //y=1.915 //x2=7.255 //y2=1.59
cc_3627 ( N_D_c_4434_n N_noxref_25_M3_noxref_s ) capacitor c=0.0041843f \
 //x=32.815 //y=2.59 //x2=5.265 //y2=0.375
cc_3628 ( N_D_c_4502_n N_noxref_25_M3_noxref_s ) capacitor c=0.00798959f \
 //x=6.595 //y=0.91 //x2=5.265 //y2=0.375
cc_3629 ( N_D_c_4509_n N_noxref_25_M3_noxref_s ) capacitor c=0.00212176f \
 //x=7.12 //y=1.45 //x2=5.265 //y2=0.375
cc_3630 ( N_D_c_4510_n N_noxref_25_M3_noxref_s ) capacitor c=0.00298115f \
 //x=7.12 //y=1.915 //x2=5.265 //y2=0.375
cc_3631 ( N_D_c_4434_n N_noxref_26_c_9416_n ) capacitor c=0.00494691f \
 //x=32.815 //y=2.59 //x2=7.825 //y2=0.995
cc_3632 ( N_D_c_4749_p N_noxref_26_c_9416_n ) capacitor c=2.14837e-19 \
 //x=6.965 //y=0.755 //x2=7.825 //y2=0.995
cc_3633 ( N_D_c_4507_n N_noxref_26_c_9416_n ) capacitor c=0.00123426f //x=7.12 \
 //y=0.91 //x2=7.825 //y2=0.995
cc_3634 ( N_D_c_4508_n N_noxref_26_c_9416_n ) capacitor c=0.0129288f //x=7.12 \
 //y=1.22 //x2=7.825 //y2=0.995
cc_3635 ( N_D_c_4509_n N_noxref_26_c_9416_n ) capacitor c=0.00142359f //x=7.12 \
 //y=1.45 //x2=7.825 //y2=0.995
cc_3636 ( N_D_c_4502_n N_noxref_26_M4_noxref_d ) capacitor c=0.00223875f \
 //x=6.595 //y=0.91 //x2=6.67 //y2=0.91
cc_3637 ( N_D_c_4505_n N_noxref_26_M4_noxref_d ) capacitor c=0.00262485f \
 //x=6.595 //y=1.22 //x2=6.67 //y2=0.91
cc_3638 ( N_D_c_4749_p N_noxref_26_M4_noxref_d ) capacitor c=0.00220746f \
 //x=6.965 //y=0.755 //x2=6.67 //y2=0.91
cc_3639 ( N_D_c_4756_p N_noxref_26_M4_noxref_d ) capacitor c=0.00194798f \
 //x=6.965 //y=1.375 //x2=6.67 //y2=0.91
cc_3640 ( N_D_c_4507_n N_noxref_26_M4_noxref_d ) capacitor c=0.00198465f \
 //x=7.12 //y=0.91 //x2=6.67 //y2=0.91
cc_3641 ( N_D_c_4508_n N_noxref_26_M4_noxref_d ) capacitor c=0.00128384f \
 //x=7.12 //y=1.22 //x2=6.67 //y2=0.91
cc_3642 ( N_D_c_4434_n N_noxref_26_M5_noxref_s ) capacitor c=0.00448771f \
 //x=32.815 //y=2.59 //x2=7.775 //y2=0.375
cc_3643 ( N_D_c_4507_n N_noxref_26_M5_noxref_s ) capacitor c=7.21316e-19 \
 //x=7.12 //y=0.91 //x2=7.775 //y2=0.375
cc_3644 ( N_D_c_4508_n N_noxref_26_M5_noxref_s ) capacitor c=0.00348171f \
 //x=7.12 //y=1.22 //x2=7.775 //y2=0.375
cc_3645 ( N_D_c_4567_n N_noxref_35_c_9885_n ) capacitor c=0.0167228f \
 //x=32.495 //y=0.91 //x2=33.155 //y2=0.54
cc_3646 ( N_D_c_4572_n N_noxref_35_c_9885_n ) capacitor c=0.00534519f \
 //x=33.02 //y=0.91 //x2=33.155 //y2=0.54
cc_3647 ( N_D_c_4449_n N_noxref_35_c_9908_n ) capacitor c=0.0120267f //x=32.93 \
 //y=2.08 //x2=33.155 //y2=1.59
cc_3648 ( N_D_c_4570_n N_noxref_35_c_9908_n ) capacitor c=0.0157358f \
 //x=32.495 //y=1.22 //x2=33.155 //y2=1.59
cc_3649 ( N_D_c_4575_n N_noxref_35_c_9908_n ) capacitor c=0.021347f //x=33.02 \
 //y=1.915 //x2=33.155 //y2=1.59
cc_3650 ( N_D_c_4567_n N_noxref_35_M19_noxref_s ) capacitor c=0.00798959f \
 //x=32.495 //y=0.91 //x2=31.165 //y2=0.375
cc_3651 ( N_D_c_4574_n N_noxref_35_M19_noxref_s ) capacitor c=0.00212176f \
 //x=33.02 //y=1.45 //x2=31.165 //y2=0.375
cc_3652 ( N_D_c_4575_n N_noxref_35_M19_noxref_s ) capacitor c=0.00298115f \
 //x=33.02 //y=1.915 //x2=31.165 //y2=0.375
cc_3653 ( N_D_c_4770_p N_noxref_36_c_9927_n ) capacitor c=2.14837e-19 \
 //x=32.865 //y=0.755 //x2=33.725 //y2=0.995
cc_3654 ( N_D_c_4572_n N_noxref_36_c_9927_n ) capacitor c=0.00123426f \
 //x=33.02 //y=0.91 //x2=33.725 //y2=0.995
cc_3655 ( N_D_c_4573_n N_noxref_36_c_9927_n ) capacitor c=0.0129288f //x=33.02 \
 //y=1.22 //x2=33.725 //y2=0.995
cc_3656 ( N_D_c_4574_n N_noxref_36_c_9927_n ) capacitor c=0.00142359f \
 //x=33.02 //y=1.45 //x2=33.725 //y2=0.995
cc_3657 ( N_D_c_4567_n N_noxref_36_M20_noxref_d ) capacitor c=0.00223875f \
 //x=32.495 //y=0.91 //x2=32.57 //y2=0.91
cc_3658 ( N_D_c_4570_n N_noxref_36_M20_noxref_d ) capacitor c=0.00262485f \
 //x=32.495 //y=1.22 //x2=32.57 //y2=0.91
cc_3659 ( N_D_c_4770_p N_noxref_36_M20_noxref_d ) capacitor c=0.00220746f \
 //x=32.865 //y=0.755 //x2=32.57 //y2=0.91
cc_3660 ( N_D_c_4777_p N_noxref_36_M20_noxref_d ) capacitor c=0.00194798f \
 //x=32.865 //y=1.375 //x2=32.57 //y2=0.91
cc_3661 ( N_D_c_4572_n N_noxref_36_M20_noxref_d ) capacitor c=0.00198465f \
 //x=33.02 //y=0.91 //x2=32.57 //y2=0.91
cc_3662 ( N_D_c_4573_n N_noxref_36_M20_noxref_d ) capacitor c=0.00128384f \
 //x=33.02 //y=1.22 //x2=32.57 //y2=0.91
cc_3663 ( N_D_c_4572_n N_noxref_36_M21_noxref_s ) capacitor c=7.21316e-19 \
 //x=33.02 //y=0.91 //x2=33.675 //y2=0.375
cc_3664 ( N_D_c_4573_n N_noxref_36_M21_noxref_s ) capacitor c=0.00348171f \
 //x=33.02 //y=1.22 //x2=33.675 //y2=0.375
cc_3665 ( N_D_c_4615_p N_noxref_45_c_10396_n ) capacitor c=0.0167228f \
 //x=58.395 //y=0.91 //x2=59.055 //y2=0.54
cc_3666 ( N_D_c_4621_p N_noxref_45_c_10396_n ) capacitor c=0.00534519f \
 //x=58.92 //y=0.91 //x2=59.055 //y2=0.54
cc_3667 ( N_D_c_4450_n N_noxref_45_c_10406_n ) capacitor c=0.0117694f \
 //x=58.83 //y=2.08 //x2=59.055 //y2=1.59
cc_3668 ( N_D_c_4617_p N_noxref_45_c_10406_n ) capacitor c=0.0157358f \
 //x=58.395 //y=1.22 //x2=59.055 //y2=1.59
cc_3669 ( N_D_c_4610_p N_noxref_45_c_10406_n ) capacitor c=0.021347f //x=58.92 \
 //y=1.915 //x2=59.055 //y2=1.59
cc_3670 ( N_D_c_4615_p N_noxref_45_M35_noxref_s ) capacitor c=0.00798959f \
 //x=58.395 //y=0.91 //x2=57.065 //y2=0.375
cc_3671 ( N_D_c_4624_p N_noxref_45_M35_noxref_s ) capacitor c=0.00212176f \
 //x=58.92 //y=1.45 //x2=57.065 //y2=0.375
cc_3672 ( N_D_c_4610_p N_noxref_45_M35_noxref_s ) capacitor c=0.00298115f \
 //x=58.92 //y=1.915 //x2=57.065 //y2=0.375
cc_3673 ( N_D_c_4790_p N_noxref_46_c_10438_n ) capacitor c=2.14837e-19 \
 //x=58.765 //y=0.755 //x2=59.625 //y2=0.995
cc_3674 ( N_D_c_4621_p N_noxref_46_c_10438_n ) capacitor c=0.00123426f \
 //x=58.92 //y=0.91 //x2=59.625 //y2=0.995
cc_3675 ( N_D_c_4623_p N_noxref_46_c_10438_n ) capacitor c=0.0129288f \
 //x=58.92 //y=1.22 //x2=59.625 //y2=0.995
cc_3676 ( N_D_c_4624_p N_noxref_46_c_10438_n ) capacitor c=0.00142359f \
 //x=58.92 //y=1.45 //x2=59.625 //y2=0.995
cc_3677 ( N_D_c_4615_p N_noxref_46_M36_noxref_d ) capacitor c=0.00223875f \
 //x=58.395 //y=0.91 //x2=58.47 //y2=0.91
cc_3678 ( N_D_c_4617_p N_noxref_46_M36_noxref_d ) capacitor c=0.00262485f \
 //x=58.395 //y=1.22 //x2=58.47 //y2=0.91
cc_3679 ( N_D_c_4790_p N_noxref_46_M36_noxref_d ) capacitor c=0.00220746f \
 //x=58.765 //y=0.755 //x2=58.47 //y2=0.91
cc_3680 ( N_D_c_4797_p N_noxref_46_M36_noxref_d ) capacitor c=0.00194798f \
 //x=58.765 //y=1.375 //x2=58.47 //y2=0.91
cc_3681 ( N_D_c_4621_p N_noxref_46_M36_noxref_d ) capacitor c=0.00198465f \
 //x=58.92 //y=0.91 //x2=58.47 //y2=0.91
cc_3682 ( N_D_c_4623_p N_noxref_46_M36_noxref_d ) capacitor c=0.00128384f \
 //x=58.92 //y=1.22 //x2=58.47 //y2=0.91
cc_3683 ( N_D_c_4621_p N_noxref_46_M37_noxref_s ) capacitor c=7.21316e-19 \
 //x=58.92 //y=0.91 //x2=59.575 //y2=0.375
cc_3684 ( N_D_c_4623_p N_noxref_46_M37_noxref_s ) capacitor c=0.00348171f \
 //x=58.92 //y=1.22 //x2=59.575 //y2=0.375
cc_3685 ( N_CLK_c_4880_n N_noxref_14_c_5684_n ) capacitor c=0.00910993f \
 //x=66.855 //y=4.44 //x2=57.605 //y2=3.7
cc_3686 ( N_CLK_c_4880_n N_noxref_14_c_5685_n ) capacitor c=7.95009e-19 \
 //x=66.855 //y=4.44 //x2=55.985 //y2=3.7
cc_3687 ( N_CLK_c_4880_n N_noxref_14_c_5659_n ) capacitor c=0.06678f \
 //x=66.855 //y=4.44 //x2=70.555 //y2=3.7
cc_3688 ( N_CLK_c_4807_n N_noxref_14_c_5659_n ) capacitor c=0.0190398f \
 //x=66.97 //y=2.08 //x2=70.555 //y2=3.7
cc_3689 ( N_CLK_c_4880_n N_noxref_14_c_5660_n ) capacitor c=6.59178e-19 \
 //x=66.855 //y=4.44 //x2=57.835 //y2=3.7
cc_3690 ( N_CLK_c_4897_n N_noxref_14_c_5611_n ) capacitor c=0.00241768f \
 //x=54.135 //y=4.44 //x2=54.125 //y2=5.155
cc_3691 ( N_CLK_c_4806_n N_noxref_14_c_5611_n ) capacitor c=0.014564f \
 //x=54.02 //y=2.08 //x2=54.125 //y2=5.155
cc_3692 ( N_CLK_M120_noxref_g N_noxref_14_c_5611_n ) capacitor c=0.016514f \
 //x=53.99 //y=6.02 //x2=54.125 //y2=5.155
cc_3693 ( N_CLK_c_5242_p N_noxref_14_c_5611_n ) capacitor c=0.00322046f \
 //x=54.02 //y=4.7 //x2=54.125 //y2=5.155
cc_3694 ( N_CLK_c_4862_n N_noxref_14_c_5615_n ) capacitor c=0.0219114f \
 //x=53.905 //y=4.44 //x2=53.415 //y2=5.155
cc_3695 ( N_CLK_M121_noxref_g N_noxref_14_c_5617_n ) capacitor c=0.01736f \
 //x=54.43 //y=6.02 //x2=55.005 //y2=5.155
cc_3696 ( N_CLK_c_4880_n N_noxref_14_c_5621_n ) capacitor c=0.0183122f \
 //x=66.855 //y=4.44 //x2=55.785 //y2=5.155
cc_3697 ( N_CLK_c_4880_n N_noxref_14_c_5625_n ) capacitor c=0.0210274f \
 //x=66.855 //y=4.44 //x2=55.87 //y2=3.7
cc_3698 ( N_CLK_c_4806_n N_noxref_14_c_5625_n ) capacitor c=0.00246013f \
 //x=54.02 //y=2.08 //x2=55.87 //y2=3.7
cc_3699 ( N_CLK_c_4880_n N_noxref_14_c_5588_n ) capacitor c=0.0208709f \
 //x=66.855 //y=4.44 //x2=57.72 //y2=2.08
cc_3700 ( N_CLK_c_4880_n N_noxref_14_c_5699_n ) capacitor c=0.0311227f \
 //x=66.855 //y=4.44 //x2=54.21 //y2=5.155
cc_3701 ( N_CLK_c_5250_p N_noxref_14_c_5699_n ) capacitor c=0.00426767f \
 //x=54.355 //y=4.79 //x2=54.21 //y2=5.155
cc_3702 ( N_CLK_c_4880_n N_noxref_14_c_5640_n ) capacitor c=0.0166984f \
 //x=66.855 //y=4.44 //x2=57.995 //y2=4.79
cc_3703 ( N_CLK_M120_noxref_g N_noxref_14_M120_noxref_d ) capacitor \
 c=0.0180032f //x=53.99 //y=6.02 //x2=54.065 //y2=5.02
cc_3704 ( N_CLK_M121_noxref_g N_noxref_14_M120_noxref_d ) capacitor \
 c=0.0180032f //x=54.43 //y=6.02 //x2=54.065 //y2=5.02
cc_3705 ( N_CLK_c_4803_n N_RN_c_5846_n ) capacitor c=0.0193884f //x=15.17 \
 //y=2.08 //x2=16.165 //y2=2.22
cc_3706 ( N_CLK_c_4984_n N_RN_c_5846_n ) capacitor c=0.00583058f //x=15.26 \
 //y=1.915 //x2=16.165 //y2=2.22
cc_3707 ( N_CLK_c_4803_n N_RN_c_5860_n ) capacitor c=0.00165648f //x=15.17 \
 //y=2.08 //x2=16.395 //y2=2.22
cc_3708 ( N_CLK_c_4984_n N_RN_c_5860_n ) capacitor c=2.3323e-19 //x=15.26 \
 //y=1.915 //x2=16.395 //y2=2.22
cc_3709 ( N_CLK_c_4804_n N_RN_c_5861_n ) capacitor c=0.0193884f //x=28.12 \
 //y=2.08 //x2=33.925 //y2=2.22
cc_3710 ( N_CLK_c_5097_n N_RN_c_5861_n ) capacitor c=0.00583058f //x=28.21 \
 //y=1.915 //x2=33.925 //y2=2.22
cc_3711 ( N_CLK_c_4805_n N_RN_c_5873_n ) capacitor c=0.0193884f //x=41.07 \
 //y=2.08 //x2=42.065 //y2=2.22
cc_3712 ( N_CLK_c_5126_n N_RN_c_5873_n ) capacitor c=0.00583058f //x=41.16 \
 //y=1.915 //x2=42.065 //y2=2.22
cc_3713 ( N_CLK_c_4805_n N_RN_c_5886_n ) capacitor c=0.00165648f //x=41.07 \
 //y=2.08 //x2=42.295 //y2=2.22
cc_3714 ( N_CLK_c_5126_n N_RN_c_5886_n ) capacitor c=2.3323e-19 //x=41.16 \
 //y=1.915 //x2=42.295 //y2=2.22
cc_3715 ( N_CLK_c_4806_n N_RN_c_5887_n ) capacitor c=0.0193884f //x=54.02 \
 //y=2.08 //x2=59.825 //y2=2.22
cc_3716 ( N_CLK_c_5265_p N_RN_c_5887_n ) capacitor c=0.00583058f //x=54.11 \
 //y=1.915 //x2=59.825 //y2=2.22
cc_3717 ( N_CLK_c_4807_n N_RN_c_5899_n ) capacitor c=0.021729f //x=66.97 \
 //y=2.08 //x2=67.965 //y2=2.22
cc_3718 ( N_CLK_c_5267_p N_RN_c_5899_n ) capacitor c=0.00583058f //x=67.06 \
 //y=1.915 //x2=67.965 //y2=2.22
cc_3719 ( N_CLK_c_4807_n N_RN_c_5912_n ) capacitor c=0.00165648f //x=66.97 \
 //y=2.08 //x2=68.195 //y2=2.22
cc_3720 ( N_CLK_c_5267_p N_RN_c_5912_n ) capacitor c=2.3323e-19 //x=67.06 \
 //y=1.915 //x2=68.195 //y2=2.22
cc_3721 ( N_CLK_c_4808_n N_RN_c_5913_n ) capacitor c=0.0200057f //x=15.055 \
 //y=4.44 //x2=8.14 //y2=2.08
cc_3722 ( N_CLK_c_4826_n N_RN_c_5914_n ) capacitor c=0.0200057f //x=28.005 \
 //y=4.44 //x2=16.28 //y2=2.08
cc_3723 ( N_CLK_c_4843_n N_RN_c_5914_n ) capacitor c=0.00153281f //x=15.285 \
 //y=4.44 //x2=16.28 //y2=2.08
cc_3724 ( N_CLK_c_4803_n N_RN_c_5914_n ) capacitor c=0.0459525f //x=15.17 \
 //y=2.08 //x2=16.28 //y2=2.08
cc_3725 ( N_CLK_c_4984_n N_RN_c_5914_n ) capacitor c=0.00203728f //x=15.26 \
 //y=1.915 //x2=16.28 //y2=2.08
cc_3726 ( N_CLK_c_4986_n N_RN_c_5914_n ) capacitor c=0.00142741f //x=15.17 \
 //y=4.7 //x2=16.28 //y2=2.08
cc_3727 ( N_CLK_c_4826_n N_RN_c_5915_n ) capacitor c=0.0210462f //x=28.005 \
 //y=4.44 //x2=19.98 //y2=2.08
cc_3728 ( N_CLK_c_4844_n N_RN_c_5916_n ) capacitor c=0.0200057f //x=40.955 \
 //y=4.44 //x2=34.04 //y2=2.08
cc_3729 ( N_CLK_c_4862_n N_RN_c_5917_n ) capacitor c=0.0200057f //x=53.905 \
 //y=4.44 //x2=42.18 //y2=2.08
cc_3730 ( N_CLK_c_4879_n N_RN_c_5917_n ) capacitor c=0.00153281f //x=41.185 \
 //y=4.44 //x2=42.18 //y2=2.08
cc_3731 ( N_CLK_c_4805_n N_RN_c_5917_n ) capacitor c=0.0435729f //x=41.07 \
 //y=2.08 //x2=42.18 //y2=2.08
cc_3732 ( N_CLK_c_5126_n N_RN_c_5917_n ) capacitor c=0.00203728f //x=41.16 \
 //y=1.915 //x2=42.18 //y2=2.08
cc_3733 ( N_CLK_c_5128_n N_RN_c_5917_n ) capacitor c=0.00142741f //x=41.07 \
 //y=4.7 //x2=42.18 //y2=2.08
cc_3734 ( N_CLK_c_4862_n N_RN_c_5918_n ) capacitor c=0.0210462f //x=53.905 \
 //y=4.44 //x2=45.88 //y2=2.08
cc_3735 ( N_CLK_c_4880_n N_RN_c_5919_n ) capacitor c=0.0200057f //x=66.855 \
 //y=4.44 //x2=59.94 //y2=2.08
cc_3736 ( N_CLK_c_4880_n N_RN_c_5920_n ) capacitor c=0.00551083f //x=66.855 \
 //y=4.44 //x2=68.08 //y2=2.08
cc_3737 ( N_CLK_c_4807_n N_RN_c_5920_n ) capacitor c=0.0446428f //x=66.97 \
 //y=2.08 //x2=68.08 //y2=2.08
cc_3738 ( N_CLK_c_5267_p N_RN_c_5920_n ) capacitor c=0.00203728f //x=67.06 \
 //y=1.915 //x2=68.08 //y2=2.08
cc_3739 ( N_CLK_c_5288_p N_RN_c_5920_n ) capacitor c=0.00142741f //x=66.97 \
 //y=4.7 //x2=68.08 //y2=2.08
cc_3740 ( N_CLK_M72_noxref_g N_RN_M74_noxref_g ) capacitor c=0.0101598f \
 //x=15.14 //y=6.02 //x2=16.02 //y2=6.02
cc_3741 ( N_CLK_M73_noxref_g N_RN_M74_noxref_g ) capacitor c=0.0602553f \
 //x=15.58 //y=6.02 //x2=16.02 //y2=6.02
cc_3742 ( N_CLK_M73_noxref_g N_RN_M75_noxref_g ) capacitor c=0.0101598f \
 //x=15.58 //y=6.02 //x2=16.46 //y2=6.02
cc_3743 ( N_CLK_M104_noxref_g N_RN_M106_noxref_g ) capacitor c=0.0101598f \
 //x=41.04 //y=6.02 //x2=41.92 //y2=6.02
cc_3744 ( N_CLK_M105_noxref_g N_RN_M106_noxref_g ) capacitor c=0.0602553f \
 //x=41.48 //y=6.02 //x2=41.92 //y2=6.02
cc_3745 ( N_CLK_M105_noxref_g N_RN_M107_noxref_g ) capacitor c=0.0101598f \
 //x=41.48 //y=6.02 //x2=42.36 //y2=6.02
cc_3746 ( N_CLK_M136_noxref_g N_RN_M138_noxref_g ) capacitor c=0.0101598f \
 //x=66.94 //y=6.02 //x2=67.82 //y2=6.02
cc_3747 ( N_CLK_M137_noxref_g N_RN_M138_noxref_g ) capacitor c=0.0602553f \
 //x=67.38 //y=6.02 //x2=67.82 //y2=6.02
cc_3748 ( N_CLK_M137_noxref_g N_RN_M139_noxref_g ) capacitor c=0.0101598f \
 //x=67.38 //y=6.02 //x2=68.26 //y2=6.02
cc_3749 ( N_CLK_c_4981_n N_RN_c_6075_n ) capacitor c=0.00456962f //x=15.26 \
 //y=0.91 //x2=16.27 //y2=0.915
cc_3750 ( N_CLK_c_4982_n N_RN_c_6076_n ) capacitor c=0.00438372f //x=15.26 \
 //y=1.22 //x2=16.27 //y2=1.26
cc_3751 ( N_CLK_c_4983_n N_RN_c_6077_n ) capacitor c=0.00438372f //x=15.26 \
 //y=1.45 //x2=16.27 //y2=1.57
cc_3752 ( N_CLK_c_4826_n N_RN_c_6084_n ) capacitor c=0.0085986f //x=28.005 \
 //y=4.44 //x2=20.315 //y2=4.79
cc_3753 ( N_CLK_c_5123_n N_RN_c_6196_n ) capacitor c=0.00456962f //x=41.16 \
 //y=0.91 //x2=42.17 //y2=0.915
cc_3754 ( N_CLK_c_5124_n N_RN_c_6197_n ) capacitor c=0.00438372f //x=41.16 \
 //y=1.22 //x2=42.17 //y2=1.26
cc_3755 ( N_CLK_c_5125_n N_RN_c_6198_n ) capacitor c=0.00438372f //x=41.16 \
 //y=1.45 //x2=42.17 //y2=1.57
cc_3756 ( N_CLK_c_4862_n N_RN_c_6172_n ) capacitor c=0.0085986f //x=53.905 \
 //y=4.44 //x2=46.215 //y2=4.79
cc_3757 ( N_CLK_c_5306_p N_RN_c_6341_n ) capacitor c=0.00456962f //x=67.06 \
 //y=0.91 //x2=68.07 //y2=0.915
cc_3758 ( N_CLK_c_5307_p N_RN_c_6342_n ) capacitor c=0.00438372f //x=67.06 \
 //y=1.22 //x2=68.07 //y2=1.26
cc_3759 ( N_CLK_c_5308_p N_RN_c_6343_n ) capacitor c=0.00438372f //x=67.06 \
 //y=1.45 //x2=68.07 //y2=1.57
cc_3760 ( N_CLK_c_4808_n N_RN_c_6000_n ) capacitor c=0.0111881f //x=15.055 \
 //y=4.44 //x2=8.14 //y2=4.7
cc_3761 ( N_CLK_c_4803_n N_RN_c_6085_n ) capacitor c=0.00201097f //x=15.17 \
 //y=2.08 //x2=16.28 //y2=2.08
cc_3762 ( N_CLK_c_4984_n N_RN_c_6085_n ) capacitor c=0.00828003f //x=15.26 \
 //y=1.915 //x2=16.28 //y2=2.08
cc_3763 ( N_CLK_c_4984_n N_RN_c_6086_n ) capacitor c=0.00438372f //x=15.26 \
 //y=1.915 //x2=16.28 //y2=1.915
cc_3764 ( N_CLK_c_4826_n N_RN_c_6088_n ) capacitor c=0.0111881f //x=28.005 \
 //y=4.44 //x2=16.28 //y2=4.7
cc_3765 ( N_CLK_c_4803_n N_RN_c_6088_n ) capacitor c=0.00218014f //x=15.17 \
 //y=2.08 //x2=16.28 //y2=4.7
cc_3766 ( N_CLK_c_5070_n N_RN_c_6088_n ) capacitor c=0.0611812f //x=15.505 \
 //y=4.79 //x2=16.28 //y2=4.7
cc_3767 ( N_CLK_c_4986_n N_RN_c_6088_n ) capacitor c=0.00487508f //x=15.17 \
 //y=4.7 //x2=16.28 //y2=4.7
cc_3768 ( N_CLK_c_4826_n N_RN_c_6039_n ) capacitor c=0.00293313f //x=28.005 \
 //y=4.44 //x2=19.98 //y2=4.7
cc_3769 ( N_CLK_c_4844_n N_RN_c_6121_n ) capacitor c=0.0111881f //x=40.955 \
 //y=4.44 //x2=34.04 //y2=4.7
cc_3770 ( N_CLK_c_4805_n N_RN_c_6205_n ) capacitor c=0.00201097f //x=41.07 \
 //y=2.08 //x2=42.18 //y2=2.08
cc_3771 ( N_CLK_c_5126_n N_RN_c_6205_n ) capacitor c=0.00828003f //x=41.16 \
 //y=1.915 //x2=42.18 //y2=2.08
cc_3772 ( N_CLK_c_5126_n N_RN_c_6206_n ) capacitor c=0.00438372f //x=41.16 \
 //y=1.915 //x2=42.18 //y2=1.915
cc_3773 ( N_CLK_c_4862_n N_RN_c_6208_n ) capacitor c=0.0111881f //x=53.905 \
 //y=4.44 //x2=42.18 //y2=4.7
cc_3774 ( N_CLK_c_4805_n N_RN_c_6208_n ) capacitor c=0.00218014f //x=41.07 \
 //y=2.08 //x2=42.18 //y2=4.7
cc_3775 ( N_CLK_c_5215_n N_RN_c_6208_n ) capacitor c=0.0611812f //x=41.405 \
 //y=4.79 //x2=42.18 //y2=4.7
cc_3776 ( N_CLK_c_5128_n N_RN_c_6208_n ) capacitor c=0.00487508f //x=41.07 \
 //y=4.7 //x2=42.18 //y2=4.7
cc_3777 ( N_CLK_c_4862_n N_RN_c_6159_n ) capacitor c=0.00293313f //x=53.905 \
 //y=4.44 //x2=45.88 //y2=4.7
cc_3778 ( N_CLK_c_4880_n N_RN_c_6286_n ) capacitor c=0.0111881f //x=66.855 \
 //y=4.44 //x2=59.94 //y2=4.7
cc_3779 ( N_CLK_c_4807_n N_RN_c_6363_n ) capacitor c=0.00201097f //x=66.97 \
 //y=2.08 //x2=68.08 //y2=2.08
cc_3780 ( N_CLK_c_5267_p N_RN_c_6363_n ) capacitor c=0.00828003f //x=67.06 \
 //y=1.915 //x2=68.08 //y2=2.08
cc_3781 ( N_CLK_c_5267_p N_RN_c_6365_n ) capacitor c=0.00438372f //x=67.06 \
 //y=1.915 //x2=68.08 //y2=1.915
cc_3782 ( N_CLK_c_4807_n N_RN_c_6366_n ) capacitor c=0.00218014f //x=66.97 \
 //y=2.08 //x2=68.08 //y2=4.7
cc_3783 ( N_CLK_c_5332_p N_RN_c_6366_n ) capacitor c=0.0611812f //x=67.305 \
 //y=4.79 //x2=68.08 //y2=4.7
cc_3784 ( N_CLK_c_5288_p N_RN_c_6366_n ) capacitor c=0.00487508f //x=66.97 \
 //y=4.7 //x2=68.08 //y2=4.7
cc_3785 ( N_CLK_c_4862_n N_noxref_16_c_6831_n ) capacitor c=0.076217f \
 //x=53.905 //y=4.44 //x2=63.155 //y2=4.07
cc_3786 ( N_CLK_c_4880_n N_noxref_16_c_6831_n ) capacitor c=0.784553f \
 //x=66.855 //y=4.44 //x2=63.155 //y2=4.07
cc_3787 ( N_CLK_c_4897_n N_noxref_16_c_6831_n ) capacitor c=0.026534f \
 //x=54.135 //y=4.44 //x2=63.155 //y2=4.07
cc_3788 ( N_CLK_c_4806_n N_noxref_16_c_6831_n ) capacitor c=0.0231929f \
 //x=54.02 //y=2.08 //x2=63.155 //y2=4.07
cc_3789 ( N_CLK_c_4862_n N_noxref_16_c_6833_n ) capacitor c=0.0290178f \
 //x=53.905 //y=4.44 //x2=53.025 //y2=4.07
cc_3790 ( N_CLK_c_4806_n N_noxref_16_c_6833_n ) capacitor c=0.00128547f \
 //x=54.02 //y=2.08 //x2=53.025 //y2=4.07
cc_3791 ( N_CLK_c_4880_n N_noxref_16_c_6834_n ) capacitor c=0.331988f \
 //x=66.855 //y=4.44 //x2=68.705 //y2=4.07
cc_3792 ( N_CLK_c_4807_n N_noxref_16_c_6834_n ) capacitor c=0.0208526f \
 //x=66.97 //y=2.08 //x2=68.705 //y2=4.07
cc_3793 ( N_CLK_c_5332_p N_noxref_16_c_6834_n ) capacitor c=0.00660387f \
 //x=67.305 //y=4.79 //x2=68.705 //y2=4.07
cc_3794 ( N_CLK_c_4880_n N_noxref_16_c_6962_n ) capacitor c=0.0263375f \
 //x=66.855 //y=4.44 //x2=63.385 //y2=4.07
cc_3795 ( N_CLK_c_4862_n N_noxref_16_c_6801_n ) capacitor c=0.0227055f \
 //x=53.905 //y=4.44 //x2=52.91 //y2=2.08
cc_3796 ( N_CLK_c_4897_n N_noxref_16_c_6801_n ) capacitor c=0.00153281f \
 //x=54.135 //y=4.44 //x2=52.91 //y2=2.08
cc_3797 ( N_CLK_c_4806_n N_noxref_16_c_6801_n ) capacitor c=0.0434907f \
 //x=54.02 //y=2.08 //x2=52.91 //y2=2.08
cc_3798 ( N_CLK_c_5265_p N_noxref_16_c_6801_n ) capacitor c=0.00203769f \
 //x=54.11 //y=1.915 //x2=52.91 //y2=2.08
cc_3799 ( N_CLK_c_5242_p N_noxref_16_c_6801_n ) capacitor c=0.00183762f \
 //x=54.02 //y=4.7 //x2=52.91 //y2=2.08
cc_3800 ( N_CLK_c_4880_n N_noxref_16_c_6968_n ) capacitor c=0.0016972f \
 //x=66.855 //y=4.44 //x2=63.27 //y2=4.535
cc_3801 ( N_CLK_c_4880_n N_noxref_16_c_6802_n ) capacitor c=0.0207534f \
 //x=66.855 //y=4.44 //x2=63.27 //y2=2.08
cc_3802 ( N_CLK_c_4880_n N_noxref_16_c_6863_n ) capacitor c=0.00241768f \
 //x=66.855 //y=4.44 //x2=67.075 //y2=5.155
cc_3803 ( N_CLK_c_4807_n N_noxref_16_c_6863_n ) capacitor c=0.014564f \
 //x=66.97 //y=2.08 //x2=67.075 //y2=5.155
cc_3804 ( N_CLK_M136_noxref_g N_noxref_16_c_6863_n ) capacitor c=0.016514f \
 //x=66.94 //y=6.02 //x2=67.075 //y2=5.155
cc_3805 ( N_CLK_c_5288_p N_noxref_16_c_6863_n ) capacitor c=0.00322046f \
 //x=66.97 //y=4.7 //x2=67.075 //y2=5.155
cc_3806 ( N_CLK_c_4880_n N_noxref_16_c_6867_n ) capacitor c=0.0219114f \
 //x=66.855 //y=4.44 //x2=66.365 //y2=5.155
cc_3807 ( N_CLK_M137_noxref_g N_noxref_16_c_6869_n ) capacitor c=0.0184045f \
 //x=67.38 //y=6.02 //x2=67.955 //y2=5.155
cc_3808 ( N_CLK_c_4807_n N_noxref_16_c_6877_n ) capacitor c=0.0026631f \
 //x=66.97 //y=2.08 //x2=68.82 //y2=4.07
cc_3809 ( N_CLK_c_4880_n N_noxref_16_c_6977_n ) capacitor c=0.00101864f \
 //x=66.855 //y=4.44 //x2=67.16 //y2=5.155
cc_3810 ( N_CLK_c_5332_p N_noxref_16_c_6977_n ) capacitor c=0.00427771f \
 //x=67.305 //y=4.79 //x2=67.16 //y2=5.155
cc_3811 ( N_CLK_M120_noxref_g N_noxref_16_M118_noxref_g ) capacitor \
 c=0.0105869f //x=53.99 //y=6.02 //x2=53.11 //y2=6.02
cc_3812 ( N_CLK_M120_noxref_g N_noxref_16_M119_noxref_g ) capacitor c=0.10632f \
 //x=53.99 //y=6.02 //x2=53.55 //y2=6.02
cc_3813 ( N_CLK_M121_noxref_g N_noxref_16_M119_noxref_g ) capacitor \
 c=0.0101598f //x=54.43 //y=6.02 //x2=53.55 //y2=6.02
cc_3814 ( N_CLK_c_5363_p N_noxref_16_c_6809_n ) capacitor c=5.72482e-19 \
 //x=53.585 //y=0.91 //x2=52.61 //y2=0.875
cc_3815 ( N_CLK_c_5363_p N_noxref_16_c_6811_n ) capacitor c=0.00149976f \
 //x=53.585 //y=0.91 //x2=52.61 //y2=1.22
cc_3816 ( N_CLK_c_5365_p N_noxref_16_c_6812_n ) capacitor c=0.00111227f \
 //x=53.585 //y=1.22 //x2=52.61 //y2=1.53
cc_3817 ( N_CLK_c_4806_n N_noxref_16_c_6813_n ) capacitor c=0.00210802f \
 //x=54.02 //y=2.08 //x2=52.61 //y2=1.915
cc_3818 ( N_CLK_c_5265_p N_noxref_16_c_6813_n ) capacitor c=0.00834532f \
 //x=54.11 //y=1.915 //x2=52.61 //y2=1.915
cc_3819 ( N_CLK_c_5363_p N_noxref_16_c_6816_n ) capacitor c=0.0160123f \
 //x=53.585 //y=0.91 //x2=53.14 //y2=0.875
cc_3820 ( N_CLK_c_5369_p N_noxref_16_c_6816_n ) capacitor c=0.00103227f \
 //x=54.11 //y=0.91 //x2=53.14 //y2=0.875
cc_3821 ( N_CLK_c_5365_p N_noxref_16_c_6818_n ) capacitor c=0.0124075f \
 //x=53.585 //y=1.22 //x2=53.14 //y2=1.22
cc_3822 ( N_CLK_c_5371_p N_noxref_16_c_6818_n ) capacitor c=0.0010154f \
 //x=54.11 //y=1.22 //x2=53.14 //y2=1.22
cc_3823 ( N_CLK_c_5372_p N_noxref_16_c_6818_n ) capacitor c=9.23422e-19 \
 //x=54.11 //y=1.45 //x2=53.14 //y2=1.22
cc_3824 ( N_CLK_c_4806_n N_noxref_16_c_6992_n ) capacitor c=0.00147352f \
 //x=54.02 //y=2.08 //x2=53.475 //y2=4.79
cc_3825 ( N_CLK_c_5242_p N_noxref_16_c_6992_n ) capacitor c=0.0168581f \
 //x=54.02 //y=4.7 //x2=53.475 //y2=4.79
cc_3826 ( N_CLK_c_4862_n N_noxref_16_c_6916_n ) capacitor c=0.0166959f \
 //x=53.905 //y=4.44 //x2=53.185 //y2=4.79
cc_3827 ( N_CLK_c_4806_n N_noxref_16_c_6916_n ) capacitor c=0.00141297f \
 //x=54.02 //y=2.08 //x2=53.185 //y2=4.79
cc_3828 ( N_CLK_c_5242_p N_noxref_16_c_6916_n ) capacitor c=0.00484466f \
 //x=54.02 //y=4.7 //x2=53.185 //y2=4.79
cc_3829 ( N_CLK_c_4880_n N_noxref_16_c_6997_n ) capacitor c=0.00960248f \
 //x=66.855 //y=4.44 //x2=63.675 //y2=4.79
cc_3830 ( N_CLK_c_4880_n N_noxref_16_c_6998_n ) capacitor c=0.00203982f \
 //x=66.855 //y=4.44 //x2=63.3 //y2=4.7
cc_3831 ( N_CLK_M136_noxref_g N_noxref_16_M136_noxref_d ) capacitor \
 c=0.0180032f //x=66.94 //y=6.02 //x2=67.015 //y2=5.02
cc_3832 ( N_CLK_M137_noxref_g N_noxref_16_M136_noxref_d ) capacitor \
 c=0.0180032f //x=67.38 //y=6.02 //x2=67.015 //y2=5.02
cc_3833 ( N_CLK_c_4862_n N_noxref_17_c_7491_n ) capacitor c=0.0213591f \
 //x=53.905 //y=4.44 //x2=50.945 //y2=3.33
cc_3834 ( N_CLK_c_4862_n N_noxref_17_c_7495_n ) capacitor c=4.49102e-19 \
 //x=53.905 //y=4.44 //x2=47.105 //y2=3.33
cc_3835 ( N_CLK_c_4862_n N_noxref_17_c_7362_n ) capacitor c=0.0551577f \
 //x=53.905 //y=4.44 //x2=55.015 //y2=3.33
cc_3836 ( N_CLK_c_4880_n N_noxref_17_c_7362_n ) capacitor c=0.00681804f \
 //x=66.855 //y=4.44 //x2=55.015 //y2=3.33
cc_3837 ( N_CLK_c_4897_n N_noxref_17_c_7362_n ) capacitor c=5.01525e-19 \
 //x=54.135 //y=4.44 //x2=55.015 //y2=3.33
cc_3838 ( N_CLK_c_4806_n N_noxref_17_c_7362_n ) capacitor c=0.0213922f \
 //x=54.02 //y=2.08 //x2=55.015 //y2=3.33
cc_3839 ( N_CLK_c_4862_n N_noxref_17_c_7529_n ) capacitor c=0.00691318f \
 //x=53.905 //y=4.44 //x2=51.175 //y2=3.33
cc_3840 ( N_CLK_c_4880_n N_noxref_17_c_7559_n ) capacitor c=0.00360213f \
 //x=66.855 //y=4.44 //x2=60.565 //y2=3.33
cc_3841 ( N_CLK_c_4880_n N_noxref_17_c_7561_n ) capacitor c=3.0365e-19 \
 //x=66.855 //y=4.44 //x2=55.245 //y2=3.33
cc_3842 ( N_CLK_c_4806_n N_noxref_17_c_7561_n ) capacitor c=8.4254e-19 \
 //x=54.02 //y=2.08 //x2=55.245 //y2=3.33
cc_3843 ( N_CLK_c_4807_n N_noxref_17_c_7583_n ) capacitor c=0.0190562f \
 //x=66.97 //y=2.08 //x2=78.325 //y2=3.33
cc_3844 ( N_CLK_c_4807_n N_noxref_17_c_7584_n ) capacitor c=9.95819e-19 \
 //x=66.97 //y=2.08 //x2=65.975 //y2=3.33
cc_3845 ( N_CLK_c_4862_n N_noxref_17_c_7301_n ) capacitor c=0.0200057f \
 //x=53.905 //y=4.44 //x2=46.99 //y2=2.08
cc_3846 ( N_CLK_c_4862_n N_noxref_17_c_7373_n ) capacitor c=0.0185677f \
 //x=53.905 //y=4.44 //x2=50.495 //y2=5.2
cc_3847 ( N_CLK_c_4862_n N_noxref_17_c_7377_n ) capacitor c=0.018142f \
 //x=53.905 //y=4.44 //x2=49.785 //y2=5.2
cc_3848 ( N_CLK_c_4862_n N_noxref_17_c_7303_n ) capacitor c=0.0247848f \
 //x=53.905 //y=4.44 //x2=51.06 //y2=3.33
cc_3849 ( N_CLK_c_4806_n N_noxref_17_c_7303_n ) capacitor c=5.2263e-19 \
 //x=54.02 //y=2.08 //x2=51.06 //y2=3.33
cc_3850 ( N_CLK_c_4880_n N_noxref_17_c_7304_n ) capacitor c=0.0200057f \
 //x=66.855 //y=4.44 //x2=55.13 //y2=2.08
cc_3851 ( N_CLK_c_4897_n N_noxref_17_c_7304_n ) capacitor c=0.00153281f \
 //x=54.135 //y=4.44 //x2=55.13 //y2=2.08
cc_3852 ( N_CLK_c_4806_n N_noxref_17_c_7304_n ) capacitor c=0.0435157f \
 //x=54.02 //y=2.08 //x2=55.13 //y2=2.08
cc_3853 ( N_CLK_c_5265_p N_noxref_17_c_7304_n ) capacitor c=0.00205895f \
 //x=54.11 //y=1.915 //x2=55.13 //y2=2.08
cc_3854 ( N_CLK_c_5242_p N_noxref_17_c_7304_n ) capacitor c=0.00142741f \
 //x=54.02 //y=4.7 //x2=55.13 //y2=2.08
cc_3855 ( N_CLK_c_4880_n N_noxref_17_c_7385_n ) capacitor c=0.0322189f \
 //x=66.855 //y=4.44 //x2=58.935 //y2=5.155
cc_3856 ( N_CLK_c_4880_n N_noxref_17_c_7389_n ) capacitor c=0.0230136f \
 //x=66.855 //y=4.44 //x2=58.225 //y2=5.155
cc_3857 ( N_CLK_c_4880_n N_noxref_17_c_7395_n ) capacitor c=0.0183122f \
 //x=66.855 //y=4.44 //x2=60.595 //y2=5.155
cc_3858 ( N_CLK_c_4880_n N_noxref_17_c_7399_n ) capacitor c=0.0210274f \
 //x=66.855 //y=4.44 //x2=60.68 //y2=3.33
cc_3859 ( N_CLK_c_4880_n N_noxref_17_c_7306_n ) capacitor c=0.0198304f \
 //x=66.855 //y=4.44 //x2=62.53 //y2=2.08
cc_3860 ( N_CLK_c_4880_n N_noxref_17_c_7403_n ) capacitor c=0.0185297f \
 //x=66.855 //y=4.44 //x2=63.445 //y2=5.2
cc_3861 ( N_CLK_c_4880_n N_noxref_17_c_7407_n ) capacitor c=0.0181237f \
 //x=66.855 //y=4.44 //x2=62.735 //y2=5.2
cc_3862 ( N_CLK_c_4880_n N_noxref_17_c_7308_n ) capacitor c=0.0208321f \
 //x=66.855 //y=4.44 //x2=64.01 //y2=3.33
cc_3863 ( N_CLK_c_4807_n N_noxref_17_c_7308_n ) capacitor c=3.3533e-19 \
 //x=66.97 //y=2.08 //x2=64.01 //y2=3.33
cc_3864 ( N_CLK_c_4880_n N_noxref_17_c_7309_n ) capacitor c=0.0224037f \
 //x=66.855 //y=4.44 //x2=65.86 //y2=2.08
cc_3865 ( N_CLK_c_4807_n N_noxref_17_c_7309_n ) capacitor c=0.0437387f \
 //x=66.97 //y=2.08 //x2=65.86 //y2=2.08
cc_3866 ( N_CLK_c_5267_p N_noxref_17_c_7309_n ) capacitor c=0.00203769f \
 //x=67.06 //y=1.915 //x2=65.86 //y2=2.08
cc_3867 ( N_CLK_c_5288_p N_noxref_17_c_7309_n ) capacitor c=0.00183762f \
 //x=66.97 //y=4.7 //x2=65.86 //y2=2.08
cc_3868 ( N_CLK_M120_noxref_g N_noxref_17_M122_noxref_g ) capacitor \
 c=0.0101598f //x=53.99 //y=6.02 //x2=54.87 //y2=6.02
cc_3869 ( N_CLK_M121_noxref_g N_noxref_17_M122_noxref_g ) capacitor \
 c=0.0602553f //x=54.43 //y=6.02 //x2=54.87 //y2=6.02
cc_3870 ( N_CLK_M121_noxref_g N_noxref_17_M123_noxref_g ) capacitor \
 c=0.0101598f //x=54.43 //y=6.02 //x2=55.31 //y2=6.02
cc_3871 ( N_CLK_M136_noxref_g N_noxref_17_M134_noxref_g ) capacitor \
 c=0.0105869f //x=66.94 //y=6.02 //x2=66.06 //y2=6.02
cc_3872 ( N_CLK_M136_noxref_g N_noxref_17_M135_noxref_g ) capacitor c=0.10632f \
 //x=66.94 //y=6.02 //x2=66.5 //y2=6.02
cc_3873 ( N_CLK_M137_noxref_g N_noxref_17_M135_noxref_g ) capacitor \
 c=0.0101598f //x=67.38 //y=6.02 //x2=66.5 //y2=6.02
cc_3874 ( N_CLK_c_5369_p N_noxref_17_c_7614_n ) capacitor c=0.00456962f \
 //x=54.11 //y=0.91 //x2=55.12 //y2=0.915
cc_3875 ( N_CLK_c_5371_p N_noxref_17_c_7615_n ) capacitor c=0.00438372f \
 //x=54.11 //y=1.22 //x2=55.12 //y2=1.26
cc_3876 ( N_CLK_c_5372_p N_noxref_17_c_7616_n ) capacitor c=0.00438372f \
 //x=54.11 //y=1.45 //x2=55.12 //y2=1.57
cc_3877 ( N_CLK_c_5426_p N_noxref_17_c_7325_n ) capacitor c=5.72482e-19 \
 //x=66.535 //y=0.91 //x2=65.56 //y2=0.875
cc_3878 ( N_CLK_c_5426_p N_noxref_17_c_7327_n ) capacitor c=0.00149976f \
 //x=66.535 //y=0.91 //x2=65.56 //y2=1.22
cc_3879 ( N_CLK_c_5428_p N_noxref_17_c_7328_n ) capacitor c=0.00111227f \
 //x=66.535 //y=1.22 //x2=65.56 //y2=1.53
cc_3880 ( N_CLK_c_4807_n N_noxref_17_c_7329_n ) capacitor c=0.00210802f \
 //x=66.97 //y=2.08 //x2=65.56 //y2=1.915
cc_3881 ( N_CLK_c_5267_p N_noxref_17_c_7329_n ) capacitor c=0.00834532f \
 //x=67.06 //y=1.915 //x2=65.56 //y2=1.915
cc_3882 ( N_CLK_c_5426_p N_noxref_17_c_7332_n ) capacitor c=0.0160123f \
 //x=66.535 //y=0.91 //x2=66.09 //y2=0.875
cc_3883 ( N_CLK_c_5306_p N_noxref_17_c_7332_n ) capacitor c=0.00103227f \
 //x=67.06 //y=0.91 //x2=66.09 //y2=0.875
cc_3884 ( N_CLK_c_5428_p N_noxref_17_c_7334_n ) capacitor c=0.0124075f \
 //x=66.535 //y=1.22 //x2=66.09 //y2=1.22
cc_3885 ( N_CLK_c_5307_p N_noxref_17_c_7334_n ) capacitor c=0.0010154f \
 //x=67.06 //y=1.22 //x2=66.09 //y2=1.22
cc_3886 ( N_CLK_c_5308_p N_noxref_17_c_7334_n ) capacitor c=9.23422e-19 \
 //x=67.06 //y=1.45 //x2=66.09 //y2=1.22
cc_3887 ( N_CLK_c_4807_n N_noxref_17_c_7627_n ) capacitor c=0.00147352f \
 //x=66.97 //y=2.08 //x2=66.425 //y2=4.79
cc_3888 ( N_CLK_c_5288_p N_noxref_17_c_7627_n ) capacitor c=0.0168581f \
 //x=66.97 //y=4.7 //x2=66.425 //y2=4.79
cc_3889 ( N_CLK_c_4880_n N_noxref_17_c_7447_n ) capacitor c=0.0168539f \
 //x=66.855 //y=4.44 //x2=66.135 //y2=4.79
cc_3890 ( N_CLK_c_4807_n N_noxref_17_c_7447_n ) capacitor c=0.00141297f \
 //x=66.97 //y=2.08 //x2=66.135 //y2=4.79
cc_3891 ( N_CLK_c_5288_p N_noxref_17_c_7447_n ) capacitor c=0.00484466f \
 //x=66.97 //y=4.7 //x2=66.135 //y2=4.79
cc_3892 ( N_CLK_c_4862_n N_noxref_17_c_7522_n ) capacitor c=0.0111881f \
 //x=53.905 //y=4.44 //x2=46.99 //y2=4.7
cc_3893 ( N_CLK_c_4806_n N_noxref_17_c_7633_n ) capacitor c=0.00201097f \
 //x=54.02 //y=2.08 //x2=55.13 //y2=2.08
cc_3894 ( N_CLK_c_5265_p N_noxref_17_c_7633_n ) capacitor c=0.00828003f \
 //x=54.11 //y=1.915 //x2=55.13 //y2=2.08
cc_3895 ( N_CLK_c_5265_p N_noxref_17_c_7635_n ) capacitor c=0.00438372f \
 //x=54.11 //y=1.915 //x2=55.13 //y2=1.915
cc_3896 ( N_CLK_c_4880_n N_noxref_17_c_7636_n ) capacitor c=0.0111881f \
 //x=66.855 //y=4.44 //x2=55.13 //y2=4.7
cc_3897 ( N_CLK_c_4806_n N_noxref_17_c_7636_n ) capacitor c=0.00218014f \
 //x=54.02 //y=2.08 //x2=55.13 //y2=4.7
cc_3898 ( N_CLK_c_5250_p N_noxref_17_c_7636_n ) capacitor c=0.0611812f \
 //x=54.355 //y=4.79 //x2=55.13 //y2=4.7
cc_3899 ( N_CLK_c_5242_p N_noxref_17_c_7636_n ) capacitor c=0.00487508f \
 //x=54.02 //y=4.7 //x2=55.13 //y2=4.7
cc_3900 ( N_CLK_c_4880_n N_noxref_17_c_7451_n ) capacitor c=0.0107057f \
 //x=66.855 //y=4.44 //x2=62.53 //y2=4.7
cc_3901 ( N_CLK_c_4826_n N_noxref_20_c_8515_n ) capacitor c=0.0237816f \
 //x=28.005 //y=4.44 //x2=25.045 //y2=2.96
cc_3902 ( N_CLK_c_4826_n N_noxref_20_c_8606_n ) capacitor c=3.65189e-19 \
 //x=28.005 //y=4.44 //x2=21.205 //y2=2.96
cc_3903 ( N_CLK_c_4826_n N_noxref_20_c_8516_n ) capacitor c=0.0422962f \
 //x=28.005 //y=4.44 //x2=83.505 //y2=2.96
cc_3904 ( N_CLK_c_4844_n N_noxref_20_c_8516_n ) capacitor c=0.00594004f \
 //x=40.955 //y=4.44 //x2=83.505 //y2=2.96
cc_3905 ( N_CLK_c_4861_n N_noxref_20_c_8516_n ) capacitor c=4.4954e-19 \
 //x=28.235 //y=4.44 //x2=83.505 //y2=2.96
cc_3906 ( N_CLK_c_4862_n N_noxref_20_c_8516_n ) capacitor c=0.0214843f \
 //x=53.905 //y=4.44 //x2=83.505 //y2=2.96
cc_3907 ( N_CLK_c_4804_n N_noxref_20_c_8516_n ) capacitor c=0.0228892f \
 //x=28.12 //y=2.08 //x2=83.505 //y2=2.96
cc_3908 ( N_CLK_c_4805_n N_noxref_20_c_8516_n ) capacitor c=0.0213717f \
 //x=41.07 //y=2.08 //x2=83.505 //y2=2.96
cc_3909 ( N_CLK_c_4806_n N_noxref_20_c_8516_n ) capacitor c=0.0190322f \
 //x=54.02 //y=2.08 //x2=83.505 //y2=2.96
cc_3910 ( N_CLK_c_4807_n N_noxref_20_c_8516_n ) capacitor c=0.021326f \
 //x=66.97 //y=2.08 //x2=83.505 //y2=2.96
cc_3911 ( N_CLK_c_4826_n N_noxref_20_c_8608_n ) capacitor c=0.00454388f \
 //x=28.005 //y=4.44 //x2=25.275 //y2=2.96
cc_3912 ( N_CLK_c_4826_n N_noxref_20_c_8538_n ) capacitor c=0.0200057f \
 //x=28.005 //y=4.44 //x2=21.09 //y2=2.08
cc_3913 ( N_CLK_c_4826_n N_noxref_20_c_8560_n ) capacitor c=0.0185677f \
 //x=28.005 //y=4.44 //x2=24.595 //y2=5.2
cc_3914 ( N_CLK_c_4826_n N_noxref_20_c_8564_n ) capacitor c=0.0181237f \
 //x=28.005 //y=4.44 //x2=23.885 //y2=5.2
cc_3915 ( N_CLK_c_4826_n N_noxref_20_c_8540_n ) capacitor c=0.0257082f \
 //x=28.005 //y=4.44 //x2=25.16 //y2=2.96
cc_3916 ( N_CLK_c_4804_n N_noxref_20_c_8540_n ) capacitor c=5.89489e-19 \
 //x=28.12 //y=2.08 //x2=25.16 //y2=2.96
cc_3917 ( N_CLK_c_4826_n N_noxref_20_c_8650_n ) capacitor c=0.0111881f \
 //x=28.005 //y=4.44 //x2=21.09 //y2=4.7
cc_3918 ( N_CLK_c_5060_n N_noxref_23_c_9273_n ) capacitor c=0.0167228f \
 //x=1.785 //y=0.91 //x2=2.445 //y2=0.54
cc_3919 ( N_CLK_c_4952_n N_noxref_23_c_9273_n ) capacitor c=0.00534519f \
 //x=2.31 //y=0.91 //x2=2.445 //y2=0.54
cc_3920 ( N_CLK_c_4802_n N_noxref_23_c_9290_n ) capacitor c=0.012357f //x=2.22 \
 //y=2.08 //x2=2.445 //y2=1.59
cc_3921 ( N_CLK_c_5063_n N_noxref_23_c_9290_n ) capacitor c=0.0153476f \
 //x=1.785 //y=1.22 //x2=2.445 //y2=1.59
cc_3922 ( N_CLK_c_4955_n N_noxref_23_c_9290_n ) capacitor c=0.0230663f \
 //x=2.31 //y=1.915 //x2=2.445 //y2=1.59
cc_3923 ( N_CLK_c_5060_n N_noxref_23_M0_noxref_s ) capacitor c=0.00798959f \
 //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_3924 ( N_CLK_c_4954_n N_noxref_23_M0_noxref_s ) capacitor c=0.00212176f \
 //x=2.31 //y=1.45 //x2=0.455 //y2=0.375
cc_3925 ( N_CLK_c_4955_n N_noxref_23_M0_noxref_s ) capacitor c=0.00298115f \
 //x=2.31 //y=1.915 //x2=0.455 //y2=0.375
cc_3926 ( N_CLK_c_5475_p N_noxref_24_c_9312_n ) capacitor c=2.14837e-19 \
 //x=2.155 //y=0.755 //x2=3.015 //y2=0.995
cc_3927 ( N_CLK_c_4952_n N_noxref_24_c_9312_n ) capacitor c=0.00123426f \
 //x=2.31 //y=0.91 //x2=3.015 //y2=0.995
cc_3928 ( N_CLK_c_4953_n N_noxref_24_c_9312_n ) capacitor c=0.0129288f \
 //x=2.31 //y=1.22 //x2=3.015 //y2=0.995
cc_3929 ( N_CLK_c_4954_n N_noxref_24_c_9312_n ) capacitor c=0.00142359f \
 //x=2.31 //y=1.45 //x2=3.015 //y2=0.995
cc_3930 ( N_CLK_c_5060_n N_noxref_24_M1_noxref_d ) capacitor c=0.00223875f \
 //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_3931 ( N_CLK_c_5063_n N_noxref_24_M1_noxref_d ) capacitor c=0.00262485f \
 //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_3932 ( N_CLK_c_5475_p N_noxref_24_M1_noxref_d ) capacitor c=0.00220746f \
 //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_3933 ( N_CLK_c_5482_p N_noxref_24_M1_noxref_d ) capacitor c=0.00194798f \
 //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_3934 ( N_CLK_c_4952_n N_noxref_24_M1_noxref_d ) capacitor c=0.00198465f \
 //x=2.31 //y=0.91 //x2=1.86 //y2=0.91
cc_3935 ( N_CLK_c_4953_n N_noxref_24_M1_noxref_d ) capacitor c=0.00128384f \
 //x=2.31 //y=1.22 //x2=1.86 //y2=0.91
cc_3936 ( N_CLK_c_4952_n N_noxref_24_M2_noxref_s ) capacitor c=7.21316e-19 \
 //x=2.31 //y=0.91 //x2=2.965 //y2=0.375
cc_3937 ( N_CLK_c_4953_n N_noxref_24_M2_noxref_s ) capacitor c=0.00348171f \
 //x=2.31 //y=1.22 //x2=2.965 //y2=0.375
cc_3938 ( N_CLK_c_4976_n N_noxref_28_c_9527_n ) capacitor c=0.0167228f \
 //x=14.735 //y=0.91 //x2=15.395 //y2=0.54
cc_3939 ( N_CLK_c_4981_n N_noxref_28_c_9527_n ) capacitor c=0.00534519f \
 //x=15.26 //y=0.91 //x2=15.395 //y2=0.54
cc_3940 ( N_CLK_c_4803_n N_noxref_28_c_9550_n ) capacitor c=0.0117694f \
 //x=15.17 //y=2.08 //x2=15.395 //y2=1.59
cc_3941 ( N_CLK_c_4979_n N_noxref_28_c_9550_n ) capacitor c=0.0157358f \
 //x=14.735 //y=1.22 //x2=15.395 //y2=1.59
cc_3942 ( N_CLK_c_4984_n N_noxref_28_c_9550_n ) capacitor c=0.021347f \
 //x=15.26 //y=1.915 //x2=15.395 //y2=1.59
cc_3943 ( N_CLK_c_4976_n N_noxref_28_M8_noxref_s ) capacitor c=0.00798959f \
 //x=14.735 //y=0.91 //x2=13.405 //y2=0.375
cc_3944 ( N_CLK_c_4983_n N_noxref_28_M8_noxref_s ) capacitor c=0.00212176f \
 //x=15.26 //y=1.45 //x2=13.405 //y2=0.375
cc_3945 ( N_CLK_c_4984_n N_noxref_28_M8_noxref_s ) capacitor c=0.00298115f \
 //x=15.26 //y=1.915 //x2=13.405 //y2=0.375
cc_3946 ( N_CLK_c_5495_p N_noxref_29_c_9569_n ) capacitor c=2.14837e-19 \
 //x=15.105 //y=0.755 //x2=15.965 //y2=0.995
cc_3947 ( N_CLK_c_4981_n N_noxref_29_c_9569_n ) capacitor c=0.00123426f \
 //x=15.26 //y=0.91 //x2=15.965 //y2=0.995
cc_3948 ( N_CLK_c_4982_n N_noxref_29_c_9569_n ) capacitor c=0.0129288f \
 //x=15.26 //y=1.22 //x2=15.965 //y2=0.995
cc_3949 ( N_CLK_c_4983_n N_noxref_29_c_9569_n ) capacitor c=0.00142359f \
 //x=15.26 //y=1.45 //x2=15.965 //y2=0.995
cc_3950 ( N_CLK_c_4976_n N_noxref_29_M9_noxref_d ) capacitor c=0.00223875f \
 //x=14.735 //y=0.91 //x2=14.81 //y2=0.91
cc_3951 ( N_CLK_c_4979_n N_noxref_29_M9_noxref_d ) capacitor c=0.00262485f \
 //x=14.735 //y=1.22 //x2=14.81 //y2=0.91
cc_3952 ( N_CLK_c_5495_p N_noxref_29_M9_noxref_d ) capacitor c=0.00220746f \
 //x=15.105 //y=0.755 //x2=14.81 //y2=0.91
cc_3953 ( N_CLK_c_5502_p N_noxref_29_M9_noxref_d ) capacitor c=0.00194798f \
 //x=15.105 //y=1.375 //x2=14.81 //y2=0.91
cc_3954 ( N_CLK_c_4981_n N_noxref_29_M9_noxref_d ) capacitor c=0.00198465f \
 //x=15.26 //y=0.91 //x2=14.81 //y2=0.91
cc_3955 ( N_CLK_c_4982_n N_noxref_29_M9_noxref_d ) capacitor c=0.00128384f \
 //x=15.26 //y=1.22 //x2=14.81 //y2=0.91
cc_3956 ( N_CLK_c_4981_n N_noxref_29_M10_noxref_s ) capacitor c=7.21316e-19 \
 //x=15.26 //y=0.91 //x2=15.915 //y2=0.375
cc_3957 ( N_CLK_c_4982_n N_noxref_29_M10_noxref_s ) capacitor c=0.00348171f \
 //x=15.26 //y=1.22 //x2=15.915 //y2=0.375
cc_3958 ( N_CLK_c_5205_n N_noxref_33_c_9784_n ) capacitor c=0.0167228f \
 //x=27.685 //y=0.91 //x2=28.345 //y2=0.54
cc_3959 ( N_CLK_c_5094_n N_noxref_33_c_9784_n ) capacitor c=0.00534519f \
 //x=28.21 //y=0.91 //x2=28.345 //y2=0.54
cc_3960 ( N_CLK_c_4804_n N_noxref_33_c_9805_n ) capacitor c=0.0117694f \
 //x=28.12 //y=2.08 //x2=28.345 //y2=1.59
cc_3961 ( N_CLK_c_5208_n N_noxref_33_c_9805_n ) capacitor c=0.0157358f \
 //x=27.685 //y=1.22 //x2=28.345 //y2=1.59
cc_3962 ( N_CLK_c_5097_n N_noxref_33_c_9805_n ) capacitor c=0.021347f \
 //x=28.21 //y=1.915 //x2=28.345 //y2=1.59
cc_3963 ( N_CLK_c_5205_n N_noxref_33_M16_noxref_s ) capacitor c=0.00798959f \
 //x=27.685 //y=0.91 //x2=26.355 //y2=0.375
cc_3964 ( N_CLK_c_5096_n N_noxref_33_M16_noxref_s ) capacitor c=0.00212176f \
 //x=28.21 //y=1.45 //x2=26.355 //y2=0.375
cc_3965 ( N_CLK_c_5097_n N_noxref_33_M16_noxref_s ) capacitor c=0.00298115f \
 //x=28.21 //y=1.915 //x2=26.355 //y2=0.375
cc_3966 ( N_CLK_c_5515_p N_noxref_34_c_9826_n ) capacitor c=2.14837e-19 \
 //x=28.055 //y=0.755 //x2=28.915 //y2=0.995
cc_3967 ( N_CLK_c_5094_n N_noxref_34_c_9826_n ) capacitor c=0.00123426f \
 //x=28.21 //y=0.91 //x2=28.915 //y2=0.995
cc_3968 ( N_CLK_c_5095_n N_noxref_34_c_9826_n ) capacitor c=0.0129288f \
 //x=28.21 //y=1.22 //x2=28.915 //y2=0.995
cc_3969 ( N_CLK_c_5096_n N_noxref_34_c_9826_n ) capacitor c=0.00142359f \
 //x=28.21 //y=1.45 //x2=28.915 //y2=0.995
cc_3970 ( N_CLK_c_5205_n N_noxref_34_M17_noxref_d ) capacitor c=0.00223875f \
 //x=27.685 //y=0.91 //x2=27.76 //y2=0.91
cc_3971 ( N_CLK_c_5208_n N_noxref_34_M17_noxref_d ) capacitor c=0.00262485f \
 //x=27.685 //y=1.22 //x2=27.76 //y2=0.91
cc_3972 ( N_CLK_c_5515_p N_noxref_34_M17_noxref_d ) capacitor c=0.00220746f \
 //x=28.055 //y=0.755 //x2=27.76 //y2=0.91
cc_3973 ( N_CLK_c_5522_p N_noxref_34_M17_noxref_d ) capacitor c=0.00194798f \
 //x=28.055 //y=1.375 //x2=27.76 //y2=0.91
cc_3974 ( N_CLK_c_5094_n N_noxref_34_M17_noxref_d ) capacitor c=0.00198465f \
 //x=28.21 //y=0.91 //x2=27.76 //y2=0.91
cc_3975 ( N_CLK_c_5095_n N_noxref_34_M17_noxref_d ) capacitor c=0.00128384f \
 //x=28.21 //y=1.22 //x2=27.76 //y2=0.91
cc_3976 ( N_CLK_c_5094_n N_noxref_34_M18_noxref_s ) capacitor c=7.21316e-19 \
 //x=28.21 //y=0.91 //x2=28.865 //y2=0.375
cc_3977 ( N_CLK_c_5095_n N_noxref_34_M18_noxref_s ) capacitor c=0.00348171f \
 //x=28.21 //y=1.22 //x2=28.865 //y2=0.375
cc_3978 ( N_CLK_c_5118_n N_noxref_38_c_10038_n ) capacitor c=0.0167228f \
 //x=40.635 //y=0.91 //x2=41.295 //y2=0.54
cc_3979 ( N_CLK_c_5123_n N_noxref_38_c_10038_n ) capacitor c=0.00534519f \
 //x=41.16 //y=0.91 //x2=41.295 //y2=0.54
cc_3980 ( N_CLK_c_4805_n N_noxref_38_c_10061_n ) capacitor c=0.0117694f \
 //x=41.07 //y=2.08 //x2=41.295 //y2=1.59
cc_3981 ( N_CLK_c_5121_n N_noxref_38_c_10061_n ) capacitor c=0.0157358f \
 //x=40.635 //y=1.22 //x2=41.295 //y2=1.59
cc_3982 ( N_CLK_c_5126_n N_noxref_38_c_10061_n ) capacitor c=0.021347f \
 //x=41.16 //y=1.915 //x2=41.295 //y2=1.59
cc_3983 ( N_CLK_c_5118_n N_noxref_38_M24_noxref_s ) capacitor c=0.00798959f \
 //x=40.635 //y=0.91 //x2=39.305 //y2=0.375
cc_3984 ( N_CLK_c_5125_n N_noxref_38_M24_noxref_s ) capacitor c=0.00212176f \
 //x=41.16 //y=1.45 //x2=39.305 //y2=0.375
cc_3985 ( N_CLK_c_5126_n N_noxref_38_M24_noxref_s ) capacitor c=0.00298115f \
 //x=41.16 //y=1.915 //x2=39.305 //y2=0.375
cc_3986 ( N_CLK_c_5535_p N_noxref_39_c_10080_n ) capacitor c=2.14837e-19 \
 //x=41.005 //y=0.755 //x2=41.865 //y2=0.995
cc_3987 ( N_CLK_c_5123_n N_noxref_39_c_10080_n ) capacitor c=0.00123426f \
 //x=41.16 //y=0.91 //x2=41.865 //y2=0.995
cc_3988 ( N_CLK_c_5124_n N_noxref_39_c_10080_n ) capacitor c=0.0129288f \
 //x=41.16 //y=1.22 //x2=41.865 //y2=0.995
cc_3989 ( N_CLK_c_5125_n N_noxref_39_c_10080_n ) capacitor c=0.00142359f \
 //x=41.16 //y=1.45 //x2=41.865 //y2=0.995
cc_3990 ( N_CLK_c_5118_n N_noxref_39_M25_noxref_d ) capacitor c=0.00223875f \
 //x=40.635 //y=0.91 //x2=40.71 //y2=0.91
cc_3991 ( N_CLK_c_5121_n N_noxref_39_M25_noxref_d ) capacitor c=0.00262485f \
 //x=40.635 //y=1.22 //x2=40.71 //y2=0.91
cc_3992 ( N_CLK_c_5535_p N_noxref_39_M25_noxref_d ) capacitor c=0.00220746f \
 //x=41.005 //y=0.755 //x2=40.71 //y2=0.91
cc_3993 ( N_CLK_c_5542_p N_noxref_39_M25_noxref_d ) capacitor c=0.00194798f \
 //x=41.005 //y=1.375 //x2=40.71 //y2=0.91
cc_3994 ( N_CLK_c_5123_n N_noxref_39_M25_noxref_d ) capacitor c=0.00198465f \
 //x=41.16 //y=0.91 //x2=40.71 //y2=0.91
cc_3995 ( N_CLK_c_5124_n N_noxref_39_M25_noxref_d ) capacitor c=0.00128384f \
 //x=41.16 //y=1.22 //x2=40.71 //y2=0.91
cc_3996 ( N_CLK_c_5123_n N_noxref_39_M26_noxref_s ) capacitor c=7.21316e-19 \
 //x=41.16 //y=0.91 //x2=41.815 //y2=0.375
cc_3997 ( N_CLK_c_5124_n N_noxref_39_M26_noxref_s ) capacitor c=0.00348171f \
 //x=41.16 //y=1.22 //x2=41.815 //y2=0.375
cc_3998 ( N_CLK_c_5363_p N_noxref_43_c_10295_n ) capacitor c=0.0167228f \
 //x=53.585 //y=0.91 //x2=54.245 //y2=0.54
cc_3999 ( N_CLK_c_5369_p N_noxref_43_c_10295_n ) capacitor c=0.00534519f \
 //x=54.11 //y=0.91 //x2=54.245 //y2=0.54
cc_4000 ( N_CLK_c_4806_n N_noxref_43_c_10305_n ) capacitor c=0.0117694f \
 //x=54.02 //y=2.08 //x2=54.245 //y2=1.59
cc_4001 ( N_CLK_c_5365_p N_noxref_43_c_10305_n ) capacitor c=0.0157358f \
 //x=53.585 //y=1.22 //x2=54.245 //y2=1.59
cc_4002 ( N_CLK_c_5265_p N_noxref_43_c_10305_n ) capacitor c=0.021347f \
 //x=54.11 //y=1.915 //x2=54.245 //y2=1.59
cc_4003 ( N_CLK_c_5363_p N_noxref_43_M32_noxref_s ) capacitor c=0.00798959f \
 //x=53.585 //y=0.91 //x2=52.255 //y2=0.375
cc_4004 ( N_CLK_c_5372_p N_noxref_43_M32_noxref_s ) capacitor c=0.00212176f \
 //x=54.11 //y=1.45 //x2=52.255 //y2=0.375
cc_4005 ( N_CLK_c_5265_p N_noxref_43_M32_noxref_s ) capacitor c=0.00298115f \
 //x=54.11 //y=1.915 //x2=52.255 //y2=0.375
cc_4006 ( N_CLK_c_5555_p N_noxref_44_c_10337_n ) capacitor c=2.14837e-19 \
 //x=53.955 //y=0.755 //x2=54.815 //y2=0.995
cc_4007 ( N_CLK_c_5369_p N_noxref_44_c_10337_n ) capacitor c=0.00123426f \
 //x=54.11 //y=0.91 //x2=54.815 //y2=0.995
cc_4008 ( N_CLK_c_5371_p N_noxref_44_c_10337_n ) capacitor c=0.0129288f \
 //x=54.11 //y=1.22 //x2=54.815 //y2=0.995
cc_4009 ( N_CLK_c_5372_p N_noxref_44_c_10337_n ) capacitor c=0.00142359f \
 //x=54.11 //y=1.45 //x2=54.815 //y2=0.995
cc_4010 ( N_CLK_c_5363_p N_noxref_44_M33_noxref_d ) capacitor c=0.00223875f \
 //x=53.585 //y=0.91 //x2=53.66 //y2=0.91
cc_4011 ( N_CLK_c_5365_p N_noxref_44_M33_noxref_d ) capacitor c=0.00262485f \
 //x=53.585 //y=1.22 //x2=53.66 //y2=0.91
cc_4012 ( N_CLK_c_5555_p N_noxref_44_M33_noxref_d ) capacitor c=0.00220746f \
 //x=53.955 //y=0.755 //x2=53.66 //y2=0.91
cc_4013 ( N_CLK_c_5562_p N_noxref_44_M33_noxref_d ) capacitor c=0.00194798f \
 //x=53.955 //y=1.375 //x2=53.66 //y2=0.91
cc_4014 ( N_CLK_c_5369_p N_noxref_44_M33_noxref_d ) capacitor c=0.00198465f \
 //x=54.11 //y=0.91 //x2=53.66 //y2=0.91
cc_4015 ( N_CLK_c_5371_p N_noxref_44_M33_noxref_d ) capacitor c=0.00128384f \
 //x=54.11 //y=1.22 //x2=53.66 //y2=0.91
cc_4016 ( N_CLK_c_5369_p N_noxref_44_M34_noxref_s ) capacitor c=7.21316e-19 \
 //x=54.11 //y=0.91 //x2=54.765 //y2=0.375
cc_4017 ( N_CLK_c_5371_p N_noxref_44_M34_noxref_s ) capacitor c=0.00348171f \
 //x=54.11 //y=1.22 //x2=54.765 //y2=0.375
cc_4018 ( N_CLK_c_5426_p N_noxref_48_c_10549_n ) capacitor c=0.0167228f \
 //x=66.535 //y=0.91 //x2=67.195 //y2=0.54
cc_4019 ( N_CLK_c_5306_p N_noxref_48_c_10549_n ) capacitor c=0.00534519f \
 //x=67.06 //y=0.91 //x2=67.195 //y2=0.54
cc_4020 ( N_CLK_c_4807_n N_noxref_48_c_10559_n ) capacitor c=0.0117694f \
 //x=66.97 //y=2.08 //x2=67.195 //y2=1.59
cc_4021 ( N_CLK_c_5428_p N_noxref_48_c_10559_n ) capacitor c=0.0157358f \
 //x=66.535 //y=1.22 //x2=67.195 //y2=1.59
cc_4022 ( N_CLK_c_5267_p N_noxref_48_c_10559_n ) capacitor c=0.021347f \
 //x=67.06 //y=1.915 //x2=67.195 //y2=1.59
cc_4023 ( N_CLK_c_5426_p N_noxref_48_M40_noxref_s ) capacitor c=0.00798959f \
 //x=66.535 //y=0.91 //x2=65.205 //y2=0.375
cc_4024 ( N_CLK_c_5308_p N_noxref_48_M40_noxref_s ) capacitor c=0.00212176f \
 //x=67.06 //y=1.45 //x2=65.205 //y2=0.375
cc_4025 ( N_CLK_c_5267_p N_noxref_48_M40_noxref_s ) capacitor c=0.00298115f \
 //x=67.06 //y=1.915 //x2=65.205 //y2=0.375
cc_4026 ( N_CLK_c_5575_p N_noxref_49_c_10591_n ) capacitor c=2.14837e-19 \
 //x=66.905 //y=0.755 //x2=67.765 //y2=0.995
cc_4027 ( N_CLK_c_5306_p N_noxref_49_c_10591_n ) capacitor c=0.00123426f \
 //x=67.06 //y=0.91 //x2=67.765 //y2=0.995
cc_4028 ( N_CLK_c_5307_p N_noxref_49_c_10591_n ) capacitor c=0.0129288f \
 //x=67.06 //y=1.22 //x2=67.765 //y2=0.995
cc_4029 ( N_CLK_c_5308_p N_noxref_49_c_10591_n ) capacitor c=0.00142359f \
 //x=67.06 //y=1.45 //x2=67.765 //y2=0.995
cc_4030 ( N_CLK_c_5426_p N_noxref_49_M41_noxref_d ) capacitor c=0.00223875f \
 //x=66.535 //y=0.91 //x2=66.61 //y2=0.91
cc_4031 ( N_CLK_c_5428_p N_noxref_49_M41_noxref_d ) capacitor c=0.00262485f \
 //x=66.535 //y=1.22 //x2=66.61 //y2=0.91
cc_4032 ( N_CLK_c_5575_p N_noxref_49_M41_noxref_d ) capacitor c=0.00220746f \
 //x=66.905 //y=0.755 //x2=66.61 //y2=0.91
cc_4033 ( N_CLK_c_5582_p N_noxref_49_M41_noxref_d ) capacitor c=0.00194798f \
 //x=66.905 //y=1.375 //x2=66.61 //y2=0.91
cc_4034 ( N_CLK_c_5306_p N_noxref_49_M41_noxref_d ) capacitor c=0.00198465f \
 //x=67.06 //y=0.91 //x2=66.61 //y2=0.91
cc_4035 ( N_CLK_c_5307_p N_noxref_49_M41_noxref_d ) capacitor c=0.00128384f \
 //x=67.06 //y=1.22 //x2=66.61 //y2=0.91
cc_4036 ( N_CLK_c_5306_p N_noxref_49_M42_noxref_s ) capacitor c=7.21316e-19 \
 //x=67.06 //y=0.91 //x2=67.715 //y2=0.375
cc_4037 ( N_CLK_c_5307_p N_noxref_49_M42_noxref_s ) capacitor c=0.00348171f \
 //x=67.06 //y=1.22 //x2=67.715 //y2=0.375
cc_4038 ( N_noxref_14_c_5704_p N_RN_c_5887_n ) capacitor c=0.016327f //x=55.47 \
 //y=1.665 //x2=59.825 //y2=2.22
cc_4039 ( N_noxref_14_c_5625_n N_RN_c_5887_n ) capacitor c=0.0197307f \
 //x=55.87 //y=3.7 //x2=59.825 //y2=2.22
cc_4040 ( N_noxref_14_c_5588_n N_RN_c_5887_n ) capacitor c=0.0192695f \
 //x=57.72 //y=2.08 //x2=59.825 //y2=2.22
cc_4041 ( N_noxref_14_c_5594_n N_RN_c_5887_n ) capacitor c=0.011987f //x=57.42 \
 //y=1.915 //x2=59.825 //y2=2.22
cc_4042 ( N_noxref_14_c_5589_n N_RN_c_5908_n ) capacitor c=0.0226137f \
 //x=70.67 //y=2.08 //x2=71.665 //y2=2.22
cc_4043 ( N_noxref_14_c_5604_n N_RN_c_5908_n ) capacitor c=0.0121989f \
 //x=70.37 //y=1.915 //x2=71.665 //y2=2.22
cc_4044 ( N_noxref_14_c_5659_n N_RN_c_5919_n ) capacitor c=0.0179999f \
 //x=70.555 //y=3.7 //x2=59.94 //y2=2.08
cc_4045 ( N_noxref_14_c_5588_n N_RN_c_5919_n ) capacitor c=0.00108469f \
 //x=57.72 //y=2.08 //x2=59.94 //y2=2.08
cc_4046 ( N_noxref_14_c_5659_n N_RN_c_5920_n ) capacitor c=0.0179999f \
 //x=70.555 //y=3.7 //x2=68.08 //y2=2.08
cc_4047 ( N_noxref_14_c_5589_n N_RN_c_5920_n ) capacitor c=6.4547e-19 \
 //x=70.67 //y=2.08 //x2=68.08 //y2=2.08
cc_4048 ( N_noxref_14_c_5659_n N_RN_c_5921_n ) capacitor c=0.0027353f \
 //x=70.555 //y=3.7 //x2=71.78 //y2=2.08
cc_4049 ( N_noxref_14_c_5589_n N_RN_c_5921_n ) capacitor c=0.0475473f \
 //x=70.67 //y=2.08 //x2=71.78 //y2=2.08
cc_4050 ( N_noxref_14_c_5604_n N_RN_c_5921_n ) capacitor c=0.00208635f \
 //x=70.37 //y=1.915 //x2=71.78 //y2=2.08
cc_4051 ( N_noxref_14_c_5717_p N_RN_c_5921_n ) capacitor c=0.00147352f \
 //x=71.235 //y=4.79 //x2=71.78 //y2=2.08
cc_4052 ( N_noxref_14_c_5642_n N_RN_c_5921_n ) capacitor c=0.00142741f \
 //x=70.945 //y=4.79 //x2=71.78 //y2=2.08
cc_4053 ( N_noxref_14_M140_noxref_g N_RN_M142_noxref_g ) capacitor \
 c=0.0105869f //x=70.87 //y=6.02 //x2=71.75 //y2=6.02
cc_4054 ( N_noxref_14_M141_noxref_g N_RN_M142_noxref_g ) capacitor c=0.10632f \
 //x=71.31 //y=6.02 //x2=71.75 //y2=6.02
cc_4055 ( N_noxref_14_M141_noxref_g N_RN_M143_noxref_g ) capacitor \
 c=0.0101598f //x=71.31 //y=6.02 //x2=72.19 //y2=6.02
cc_4056 ( N_noxref_14_c_5600_n N_RN_c_6387_n ) capacitor c=5.72482e-19 \
 //x=70.37 //y=0.875 //x2=71.345 //y2=0.91
cc_4057 ( N_noxref_14_c_5602_n N_RN_c_6387_n ) capacitor c=0.00149976f \
 //x=70.37 //y=1.22 //x2=71.345 //y2=0.91
cc_4058 ( N_noxref_14_c_5607_n N_RN_c_6387_n ) capacitor c=0.0160123f //x=70.9 \
 //y=0.875 //x2=71.345 //y2=0.91
cc_4059 ( N_noxref_14_c_5603_n N_RN_c_6390_n ) capacitor c=0.00111227f \
 //x=70.37 //y=1.53 //x2=71.345 //y2=1.22
cc_4060 ( N_noxref_14_c_5609_n N_RN_c_6390_n ) capacitor c=0.0124075f //x=70.9 \
 //y=1.22 //x2=71.345 //y2=1.22
cc_4061 ( N_noxref_14_c_5607_n N_RN_c_6392_n ) capacitor c=0.00103227f \
 //x=70.9 //y=0.875 //x2=71.87 //y2=0.91
cc_4062 ( N_noxref_14_c_5609_n N_RN_c_6393_n ) capacitor c=0.0010154f //x=70.9 \
 //y=1.22 //x2=71.87 //y2=1.22
cc_4063 ( N_noxref_14_c_5609_n N_RN_c_6394_n ) capacitor c=9.23422e-19 \
 //x=70.9 //y=1.22 //x2=71.87 //y2=1.45
cc_4064 ( N_noxref_14_c_5589_n N_RN_c_6395_n ) capacitor c=0.00203769f \
 //x=70.67 //y=2.08 //x2=71.87 //y2=1.915
cc_4065 ( N_noxref_14_c_5604_n N_RN_c_6395_n ) capacitor c=0.00834532f \
 //x=70.37 //y=1.915 //x2=71.87 //y2=1.915
cc_4066 ( N_noxref_14_c_5589_n N_RN_c_6397_n ) capacitor c=0.00183762f \
 //x=70.67 //y=2.08 //x2=71.78 //y2=4.7
cc_4067 ( N_noxref_14_c_5717_p N_RN_c_6397_n ) capacitor c=0.0168581f \
 //x=71.235 //y=4.79 //x2=71.78 //y2=4.7
cc_4068 ( N_noxref_14_c_5642_n N_RN_c_6397_n ) capacitor c=0.00484466f \
 //x=70.945 //y=4.79 //x2=71.78 //y2=4.7
cc_4069 ( N_noxref_14_c_5684_n N_noxref_16_c_6831_n ) capacitor c=0.147447f \
 //x=57.605 //y=3.7 //x2=63.155 //y2=4.07
cc_4070 ( N_noxref_14_c_5685_n N_noxref_16_c_6831_n ) capacitor c=0.0294294f \
 //x=55.985 //y=3.7 //x2=63.155 //y2=4.07
cc_4071 ( N_noxref_14_c_5659_n N_noxref_16_c_6831_n ) capacitor c=0.467539f \
 //x=70.555 //y=3.7 //x2=63.155 //y2=4.07
cc_4072 ( N_noxref_14_c_5660_n N_noxref_16_c_6831_n ) capacitor c=0.0264476f \
 //x=57.835 //y=3.7 //x2=63.155 //y2=4.07
cc_4073 ( N_noxref_14_c_5625_n N_noxref_16_c_6831_n ) capacitor c=0.0200328f \
 //x=55.87 //y=3.7 //x2=63.155 //y2=4.07
cc_4074 ( N_noxref_14_c_5588_n N_noxref_16_c_6831_n ) capacitor c=0.0213516f \
 //x=57.72 //y=2.08 //x2=63.155 //y2=4.07
cc_4075 ( N_noxref_14_c_5659_n N_noxref_16_c_6834_n ) capacitor c=0.468066f \
 //x=70.555 //y=3.7 //x2=68.705 //y2=4.07
cc_4076 ( N_noxref_14_c_5659_n N_noxref_16_c_6962_n ) capacitor c=0.0267832f \
 //x=70.555 //y=3.7 //x2=63.385 //y2=4.07
cc_4077 ( N_noxref_14_c_5659_n N_noxref_16_c_6836_n ) capacitor c=0.176507f \
 //x=70.555 //y=3.7 //x2=73.515 //y2=4.07
cc_4078 ( N_noxref_14_c_5589_n N_noxref_16_c_6836_n ) capacitor c=0.0252746f \
 //x=70.67 //y=2.08 //x2=73.515 //y2=4.07
cc_4079 ( N_noxref_14_c_5642_n N_noxref_16_c_6836_n ) capacitor c=0.0115418f \
 //x=70.945 //y=4.79 //x2=73.515 //y2=4.07
cc_4080 ( N_noxref_14_c_5659_n N_noxref_16_c_6842_n ) capacitor c=0.0268461f \
 //x=70.555 //y=3.7 //x2=68.935 //y2=4.07
cc_4081 ( N_noxref_14_c_5589_n N_noxref_16_c_6842_n ) capacitor c=2.98083e-19 \
 //x=70.67 //y=2.08 //x2=68.935 //y2=4.07
cc_4082 ( N_noxref_14_c_5659_n N_noxref_16_c_6802_n ) capacitor c=0.0187965f \
 //x=70.555 //y=3.7 //x2=63.27 //y2=2.08
cc_4083 ( N_noxref_14_c_5659_n N_noxref_16_c_6877_n ) capacitor c=0.0212795f \
 //x=70.555 //y=3.7 //x2=68.82 //y2=4.07
cc_4084 ( N_noxref_14_c_5589_n N_noxref_16_c_6877_n ) capacitor c=0.0109598f \
 //x=70.67 //y=2.08 //x2=68.82 //y2=4.07
cc_4085 ( N_noxref_14_M141_noxref_g N_noxref_16_c_6878_n ) capacitor \
 c=0.0178794f //x=71.31 //y=6.02 //x2=71.885 //y2=5.155
cc_4086 ( N_noxref_14_M140_noxref_g N_noxref_16_c_6882_n ) capacitor \
 c=0.0213876f //x=70.87 //y=6.02 //x2=71.175 //y2=5.155
cc_4087 ( N_noxref_14_c_5717_p N_noxref_16_c_6882_n ) capacitor c=0.00429591f \
 //x=71.235 //y=4.79 //x2=71.175 //y2=5.155
cc_4088 ( N_noxref_14_c_5615_n N_noxref_16_M118_noxref_g ) capacitor \
 c=0.0213876f //x=53.415 //y=5.155 //x2=53.11 //y2=6.02
cc_4089 ( N_noxref_14_c_5611_n N_noxref_16_M119_noxref_g ) capacitor \
 c=0.0168349f //x=54.125 //y=5.155 //x2=53.55 //y2=6.02
cc_4090 ( N_noxref_14_M118_noxref_d N_noxref_16_M119_noxref_g ) capacitor \
 c=0.0180032f //x=53.185 //y=5.02 //x2=53.55 //y2=6.02
cc_4091 ( N_noxref_14_c_5615_n N_noxref_16_c_6992_n ) capacitor c=0.00428486f \
 //x=53.415 //y=5.155 //x2=53.475 //y2=4.79
cc_4092 ( N_noxref_14_M141_noxref_g N_noxref_16_M140_noxref_d ) capacitor \
 c=0.0180032f //x=71.31 //y=6.02 //x2=70.945 //y2=5.02
cc_4093 ( N_noxref_14_c_5684_n N_noxref_17_c_7559_n ) capacitor c=0.146539f \
 //x=57.605 //y=3.7 //x2=60.565 //y2=3.33
cc_4094 ( N_noxref_14_c_5685_n N_noxref_17_c_7559_n ) capacitor c=0.0294746f \
 //x=55.985 //y=3.7 //x2=60.565 //y2=3.33
cc_4095 ( N_noxref_14_c_5659_n N_noxref_17_c_7559_n ) capacitor c=0.238435f \
 //x=70.555 //y=3.7 //x2=60.565 //y2=3.33
cc_4096 ( N_noxref_14_c_5660_n N_noxref_17_c_7559_n ) capacitor c=0.0266966f \
 //x=57.835 //y=3.7 //x2=60.565 //y2=3.33
cc_4097 ( N_noxref_14_c_5625_n N_noxref_17_c_7559_n ) capacitor c=0.0206036f \
 //x=55.87 //y=3.7 //x2=60.565 //y2=3.33
cc_4098 ( N_noxref_14_c_5588_n N_noxref_17_c_7559_n ) capacitor c=0.0216412f \
 //x=57.72 //y=2.08 //x2=60.565 //y2=3.33
cc_4099 ( N_noxref_14_c_5625_n N_noxref_17_c_7561_n ) capacitor c=0.00179385f \
 //x=55.87 //y=3.7 //x2=55.245 //y2=3.33
cc_4100 ( N_noxref_14_c_5659_n N_noxref_17_c_7648_n ) capacitor c=0.146338f \
 //x=70.555 //y=3.7 //x2=62.415 //y2=3.33
cc_4101 ( N_noxref_14_c_5659_n N_noxref_17_c_7649_n ) capacitor c=0.0268386f \
 //x=70.555 //y=3.7 //x2=60.795 //y2=3.33
cc_4102 ( N_noxref_14_c_5659_n N_noxref_17_c_7650_n ) capacitor c=0.108749f \
 //x=70.555 //y=3.7 //x2=63.895 //y2=3.33
cc_4103 ( N_noxref_14_c_5659_n N_noxref_17_c_7651_n ) capacitor c=0.026764f \
 //x=70.555 //y=3.7 //x2=62.645 //y2=3.33
cc_4104 ( N_noxref_14_c_5659_n N_noxref_17_c_7652_n ) capacitor c=0.146498f \
 //x=70.555 //y=3.7 //x2=65.745 //y2=3.33
cc_4105 ( N_noxref_14_c_5659_n N_noxref_17_c_7653_n ) capacitor c=0.0267668f \
 //x=70.555 //y=3.7 //x2=64.125 //y2=3.33
cc_4106 ( N_noxref_14_c_5659_n N_noxref_17_c_7583_n ) capacitor c=0.433981f \
 //x=70.555 //y=3.7 //x2=78.325 //y2=3.33
cc_4107 ( N_noxref_14_c_5589_n N_noxref_17_c_7583_n ) capacitor c=0.021615f \
 //x=70.67 //y=2.08 //x2=78.325 //y2=3.33
cc_4108 ( N_noxref_14_c_5659_n N_noxref_17_c_7584_n ) capacitor c=0.0268338f \
 //x=70.555 //y=3.7 //x2=65.975 //y2=3.33
cc_4109 ( N_noxref_14_c_5615_n N_noxref_17_c_7303_n ) capacitor c=2.97874e-19 \
 //x=53.415 //y=5.155 //x2=51.06 //y2=3.33
cc_4110 ( N_noxref_14_c_5685_n N_noxref_17_c_7304_n ) capacitor c=0.00687545f \
 //x=55.985 //y=3.7 //x2=55.13 //y2=2.08
cc_4111 ( N_noxref_14_c_5625_n N_noxref_17_c_7304_n ) capacitor c=0.0760319f \
 //x=55.87 //y=3.7 //x2=55.13 //y2=2.08
cc_4112 ( N_noxref_14_c_5588_n N_noxref_17_c_7304_n ) capacitor c=8.46099e-19 \
 //x=57.72 //y=2.08 //x2=55.13 //y2=2.08
cc_4113 ( N_noxref_14_c_5779_p N_noxref_17_c_7304_n ) capacitor c=0.0171303f \
 //x=55.09 //y=5.155 //x2=55.13 //y2=2.08
cc_4114 ( N_noxref_14_M125_noxref_g N_noxref_17_c_7385_n ) capacitor \
 c=0.0168349f //x=58.36 //y=6.02 //x2=58.935 //y2=5.155
cc_4115 ( N_noxref_14_c_5621_n N_noxref_17_c_7389_n ) capacitor c=3.10026e-19 \
 //x=55.785 //y=5.155 //x2=58.225 //y2=5.155
cc_4116 ( N_noxref_14_M124_noxref_g N_noxref_17_c_7389_n ) capacitor \
 c=0.0213876f //x=57.92 //y=6.02 //x2=58.225 //y2=5.155
cc_4117 ( N_noxref_14_c_5680_n N_noxref_17_c_7389_n ) capacitor c=0.00428486f \
 //x=58.285 //y=4.79 //x2=58.225 //y2=5.155
cc_4118 ( N_noxref_14_c_5659_n N_noxref_17_c_7399_n ) capacitor c=0.0206044f \
 //x=70.555 //y=3.7 //x2=60.68 //y2=3.33
cc_4119 ( N_noxref_14_c_5659_n N_noxref_17_c_7306_n ) capacitor c=0.0205831f \
 //x=70.555 //y=3.7 //x2=62.53 //y2=2.08
cc_4120 ( N_noxref_14_c_5659_n N_noxref_17_c_7308_n ) capacitor c=0.0206034f \
 //x=70.555 //y=3.7 //x2=64.01 //y2=3.33
cc_4121 ( N_noxref_14_c_5659_n N_noxref_17_c_7309_n ) capacitor c=0.0216236f \
 //x=70.555 //y=3.7 //x2=65.86 //y2=2.08
cc_4122 ( N_noxref_14_c_5617_n N_noxref_17_M122_noxref_g ) capacitor \
 c=0.01736f //x=55.005 //y=5.155 //x2=54.87 //y2=6.02
cc_4123 ( N_noxref_14_M122_noxref_d N_noxref_17_M122_noxref_g ) capacitor \
 c=0.0180032f //x=54.945 //y=5.02 //x2=54.87 //y2=6.02
cc_4124 ( N_noxref_14_c_5621_n N_noxref_17_M123_noxref_g ) capacitor \
 c=0.0194981f //x=55.785 //y=5.155 //x2=55.31 //y2=6.02
cc_4125 ( N_noxref_14_M122_noxref_d N_noxref_17_M123_noxref_g ) capacitor \
 c=0.0194246f //x=54.945 //y=5.02 //x2=55.31 //y2=6.02
cc_4126 ( N_noxref_14_M34_noxref_d N_noxref_17_c_7614_n ) capacitor \
 c=0.00217566f //x=55.195 //y=0.915 //x2=55.12 //y2=0.915
cc_4127 ( N_noxref_14_M34_noxref_d N_noxref_17_c_7615_n ) capacitor \
 c=0.0034598f //x=55.195 //y=0.915 //x2=55.12 //y2=1.26
cc_4128 ( N_noxref_14_M34_noxref_d N_noxref_17_c_7616_n ) capacitor \
 c=0.00546784f //x=55.195 //y=0.915 //x2=55.12 //y2=1.57
cc_4129 ( N_noxref_14_M34_noxref_d N_noxref_17_c_7677_n ) capacitor \
 c=0.00241102f //x=55.195 //y=0.915 //x2=55.495 //y2=0.76
cc_4130 ( N_noxref_14_c_5587_n N_noxref_17_c_7678_n ) capacitor c=0.00371277f \
 //x=55.785 //y=1.665 //x2=55.495 //y2=1.415
cc_4131 ( N_noxref_14_M34_noxref_d N_noxref_17_c_7678_n ) capacitor \
 c=0.0138621f //x=55.195 //y=0.915 //x2=55.495 //y2=1.415
cc_4132 ( N_noxref_14_M34_noxref_d N_noxref_17_c_7680_n ) capacitor \
 c=0.00219619f //x=55.195 //y=0.915 //x2=55.65 //y2=0.915
cc_4133 ( N_noxref_14_c_5587_n N_noxref_17_c_7681_n ) capacitor c=0.00457401f \
 //x=55.785 //y=1.665 //x2=55.65 //y2=1.26
cc_4134 ( N_noxref_14_M34_noxref_d N_noxref_17_c_7681_n ) capacitor \
 c=0.00603828f //x=55.195 //y=0.915 //x2=55.65 //y2=1.26
cc_4135 ( N_noxref_14_c_5625_n N_noxref_17_c_7633_n ) capacitor c=0.00731987f \
 //x=55.87 //y=3.7 //x2=55.13 //y2=2.08
cc_4136 ( N_noxref_14_c_5625_n N_noxref_17_c_7635_n ) capacitor c=0.00283672f \
 //x=55.87 //y=3.7 //x2=55.13 //y2=1.915
cc_4137 ( N_noxref_14_M34_noxref_d N_noxref_17_c_7635_n ) capacitor \
 c=0.00661782f //x=55.195 //y=0.915 //x2=55.13 //y2=1.915
cc_4138 ( N_noxref_14_c_5621_n N_noxref_17_c_7636_n ) capacitor c=0.00201851f \
 //x=55.785 //y=5.155 //x2=55.13 //y2=4.7
cc_4139 ( N_noxref_14_c_5625_n N_noxref_17_c_7636_n ) capacitor c=0.013693f \
 //x=55.87 //y=3.7 //x2=55.13 //y2=4.7
cc_4140 ( N_noxref_14_c_5779_p N_noxref_17_c_7636_n ) capacitor c=0.00475601f \
 //x=55.09 //y=5.155 //x2=55.13 //y2=4.7
cc_4141 ( N_noxref_14_M125_noxref_g N_noxref_17_M124_noxref_d ) capacitor \
 c=0.0180032f //x=58.36 //y=6.02 //x2=57.995 //y2=5.02
cc_4142 ( N_noxref_14_c_5659_n N_noxref_18_c_8127_n ) capacitor c=0.00740361f \
 //x=70.555 //y=3.7 //x2=73.005 //y2=3.7
cc_4143 ( N_noxref_14_c_5589_n N_noxref_18_c_8065_n ) capacitor c=0.00104169f \
 //x=70.67 //y=2.08 //x2=72.89 //y2=2.08
cc_4144 ( N_noxref_14_c_5684_n N_noxref_20_c_8516_n ) capacitor c=0.0108826f \
 //x=57.605 //y=3.7 //x2=83.505 //y2=2.96
cc_4145 ( N_noxref_14_c_5685_n N_noxref_20_c_8516_n ) capacitor c=7.98411e-19 \
 //x=55.985 //y=3.7 //x2=83.505 //y2=2.96
cc_4146 ( N_noxref_14_c_5659_n N_noxref_20_c_8516_n ) capacitor c=0.096807f \
 //x=70.555 //y=3.7 //x2=83.505 //y2=2.96
cc_4147 ( N_noxref_14_c_5660_n N_noxref_20_c_8516_n ) capacitor c=5.46757e-19 \
 //x=57.835 //y=3.7 //x2=83.505 //y2=2.96
cc_4148 ( N_noxref_14_c_5625_n N_noxref_20_c_8516_n ) capacitor c=0.0187656f \
 //x=55.87 //y=3.7 //x2=83.505 //y2=2.96
cc_4149 ( N_noxref_14_c_5588_n N_noxref_20_c_8516_n ) capacitor c=0.0197816f \
 //x=57.72 //y=2.08 //x2=83.505 //y2=2.96
cc_4150 ( N_noxref_14_c_5589_n N_noxref_20_c_8516_n ) capacitor c=0.0220492f \
 //x=70.67 //y=2.08 //x2=83.505 //y2=2.96
cc_4151 ( N_noxref_14_M34_noxref_d N_noxref_43_M32_noxref_s ) capacitor \
 c=0.00309936f //x=55.195 //y=0.915 //x2=52.255 //y2=0.375
cc_4152 ( N_noxref_14_c_5587_n N_noxref_44_c_10342_n ) capacitor c=0.00457167f \
 //x=55.785 //y=1.665 //x2=55.785 //y2=0.54
cc_4153 ( N_noxref_14_M34_noxref_d N_noxref_44_c_10342_n ) capacitor \
 c=0.0115903f //x=55.195 //y=0.915 //x2=55.785 //y2=0.54
cc_4154 ( N_noxref_14_c_5704_p N_noxref_44_c_10364_n ) capacitor c=0.0200405f \
 //x=55.47 //y=1.665 //x2=54.9 //y2=0.995
cc_4155 ( N_noxref_14_M34_noxref_d N_noxref_44_M33_noxref_d ) capacitor \
 c=5.27807e-19 //x=55.195 //y=0.915 //x2=53.66 //y2=0.91
cc_4156 ( N_noxref_14_c_5587_n N_noxref_44_M34_noxref_s ) capacitor \
 c=0.0196084f //x=55.785 //y=1.665 //x2=54.765 //y2=0.375
cc_4157 ( N_noxref_14_M34_noxref_d N_noxref_44_M34_noxref_s ) capacitor \
 c=0.0426368f //x=55.195 //y=0.915 //x2=54.765 //y2=0.375
cc_4158 ( N_noxref_14_c_5587_n N_noxref_45_c_10412_n ) capacitor c=3.84569e-19 \
 //x=55.785 //y=1.665 //x2=57.2 //y2=1.505
cc_4159 ( N_noxref_14_c_5594_n N_noxref_45_c_10412_n ) capacitor c=0.0034165f \
 //x=57.42 //y=1.915 //x2=57.2 //y2=1.505
cc_4160 ( N_noxref_14_c_5588_n N_noxref_45_c_10389_n ) capacitor c=0.0115578f \
 //x=57.72 //y=2.08 //x2=58.085 //y2=1.59
cc_4161 ( N_noxref_14_c_5593_n N_noxref_45_c_10389_n ) capacitor c=0.00697148f \
 //x=57.42 //y=1.53 //x2=58.085 //y2=1.59
cc_4162 ( N_noxref_14_c_5594_n N_noxref_45_c_10389_n ) capacitor c=0.0204849f \
 //x=57.42 //y=1.915 //x2=58.085 //y2=1.59
cc_4163 ( N_noxref_14_c_5596_n N_noxref_45_c_10389_n ) capacitor c=0.00610316f \
 //x=57.795 //y=1.375 //x2=58.085 //y2=1.59
cc_4164 ( N_noxref_14_c_5599_n N_noxref_45_c_10389_n ) capacitor c=0.00698822f \
 //x=57.95 //y=1.22 //x2=58.085 //y2=1.59
cc_4165 ( N_noxref_14_c_5590_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.0327271f //x=57.42 //y=0.875 //x2=57.065 //y2=0.375
cc_4166 ( N_noxref_14_c_5593_n N_noxref_45_M35_noxref_s ) capacitor \
 c=7.99997e-19 //x=57.42 //y=1.53 //x2=57.065 //y2=0.375
cc_4167 ( N_noxref_14_c_5594_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.00122123f //x=57.42 //y=1.915 //x2=57.065 //y2=0.375
cc_4168 ( N_noxref_14_c_5597_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.0121427f //x=57.95 //y=0.875 //x2=57.065 //y2=0.375
cc_4169 ( N_noxref_14_M34_noxref_d N_noxref_45_M35_noxref_s ) capacitor \
 c=2.55333e-19 //x=55.195 //y=0.915 //x2=57.065 //y2=0.375
cc_4170 ( N_noxref_14_c_5604_n N_noxref_50_c_10659_n ) capacitor c=0.0034165f \
 //x=70.37 //y=1.915 //x2=70.15 //y2=1.505
cc_4171 ( N_noxref_14_c_5589_n N_noxref_50_c_10644_n ) capacitor c=0.0115578f \
 //x=70.67 //y=2.08 //x2=71.035 //y2=1.59
cc_4172 ( N_noxref_14_c_5603_n N_noxref_50_c_10644_n ) capacitor c=0.00697148f \
 //x=70.37 //y=1.53 //x2=71.035 //y2=1.59
cc_4173 ( N_noxref_14_c_5604_n N_noxref_50_c_10644_n ) capacitor c=0.0204849f \
 //x=70.37 //y=1.915 //x2=71.035 //y2=1.59
cc_4174 ( N_noxref_14_c_5606_n N_noxref_50_c_10644_n ) capacitor c=0.00610316f \
 //x=70.745 //y=1.375 //x2=71.035 //y2=1.59
cc_4175 ( N_noxref_14_c_5609_n N_noxref_50_c_10644_n ) capacitor c=0.00698822f \
 //x=70.9 //y=1.22 //x2=71.035 //y2=1.59
cc_4176 ( N_noxref_14_c_5600_n N_noxref_50_M43_noxref_s ) capacitor \
 c=0.0327271f //x=70.37 //y=0.875 //x2=70.015 //y2=0.375
cc_4177 ( N_noxref_14_c_5603_n N_noxref_50_M43_noxref_s ) capacitor \
 c=7.99997e-19 //x=70.37 //y=1.53 //x2=70.015 //y2=0.375
cc_4178 ( N_noxref_14_c_5604_n N_noxref_50_M43_noxref_s ) capacitor \
 c=0.00122123f //x=70.37 //y=1.915 //x2=70.015 //y2=0.375
cc_4179 ( N_noxref_14_c_5607_n N_noxref_50_M43_noxref_s ) capacitor \
 c=0.0121427f //x=70.9 //y=0.875 //x2=70.015 //y2=0.375
cc_4180 ( N_RN_c_5919_n N_noxref_16_c_6831_n ) capacitor c=0.0179722f \
 //x=59.94 //y=2.08 //x2=63.155 //y2=4.07
cc_4181 ( N_RN_c_5920_n N_noxref_16_c_6834_n ) capacitor c=0.0219145f \
 //x=68.08 //y=2.08 //x2=68.705 //y2=4.07
cc_4182 ( N_RN_c_6366_n N_noxref_16_c_6834_n ) capacitor c=0.00881004f \
 //x=68.08 //y=4.7 //x2=68.705 //y2=4.07
cc_4183 ( N_RN_c_5921_n N_noxref_16_c_6836_n ) capacitor c=0.0252951f \
 //x=71.78 //y=2.08 //x2=73.515 //y2=4.07
cc_4184 ( N_RN_c_6404_p N_noxref_16_c_6836_n ) capacitor c=0.00495688f \
 //x=72.115 //y=4.79 //x2=73.515 //y2=4.07
cc_4185 ( N_RN_c_6397_n N_noxref_16_c_6836_n ) capacitor c=0.0018068f \
 //x=71.78 //y=4.7 //x2=73.515 //y2=4.07
cc_4186 ( N_RN_c_5920_n N_noxref_16_c_6842_n ) capacitor c=0.00179385f \
 //x=68.08 //y=2.08 //x2=68.935 //y2=4.07
cc_4187 ( N_RN_c_5887_n N_noxref_16_c_6801_n ) capacitor c=0.0192695f \
 //x=59.825 //y=2.22 //x2=52.91 //y2=2.08
cc_4188 ( N_RN_c_5899_n N_noxref_16_c_6802_n ) capacitor c=0.0201924f \
 //x=67.965 //y=2.22 //x2=63.27 //y2=2.08
cc_4189 ( N_RN_M138_noxref_g N_noxref_16_c_6869_n ) capacitor c=0.0184045f \
 //x=67.82 //y=6.02 //x2=67.955 //y2=5.155
cc_4190 ( N_RN_M139_noxref_g N_noxref_16_c_6873_n ) capacitor c=0.0205426f \
 //x=68.26 //y=6.02 //x2=68.735 //y2=5.155
cc_4191 ( N_RN_c_6366_n N_noxref_16_c_6873_n ) capacitor c=0.00201851f \
 //x=68.08 //y=4.7 //x2=68.735 //y2=5.155
cc_4192 ( N_RN_c_6412_p N_noxref_16_c_6804_n ) capacitor c=0.00371277f \
 //x=68.445 //y=1.415 //x2=68.735 //y2=1.665
cc_4193 ( N_RN_c_6413_p N_noxref_16_c_6804_n ) capacitor c=0.00457401f \
 //x=68.6 //y=1.26 //x2=68.735 //y2=1.665
cc_4194 ( N_RN_c_5908_n N_noxref_16_c_7039_n ) capacitor c=0.016327f \
 //x=71.665 //y=2.22 //x2=68.42 //y2=1.665
cc_4195 ( N_RN_c_5908_n N_noxref_16_c_6877_n ) capacitor c=0.0220713f \
 //x=71.665 //y=2.22 //x2=68.82 //y2=4.07
cc_4196 ( N_RN_c_5912_n N_noxref_16_c_6877_n ) capacitor c=0.0012045f \
 //x=68.195 //y=2.22 //x2=68.82 //y2=4.07
cc_4197 ( N_RN_c_5920_n N_noxref_16_c_6877_n ) capacitor c=0.0800391f \
 //x=68.08 //y=2.08 //x2=68.82 //y2=4.07
cc_4198 ( N_RN_c_5921_n N_noxref_16_c_6877_n ) capacitor c=5.69417e-19 \
 //x=71.78 //y=2.08 //x2=68.82 //y2=4.07
cc_4199 ( N_RN_c_6363_n N_noxref_16_c_6877_n ) capacitor c=0.00709342f \
 //x=68.08 //y=2.08 //x2=68.82 //y2=4.07
cc_4200 ( N_RN_c_6365_n N_noxref_16_c_6877_n ) capacitor c=0.00283672f \
 //x=68.08 //y=1.915 //x2=68.82 //y2=4.07
cc_4201 ( N_RN_c_6366_n N_noxref_16_c_6877_n ) capacitor c=0.013693f //x=68.08 \
 //y=4.7 //x2=68.82 //y2=4.07
cc_4202 ( N_RN_c_5921_n N_noxref_16_c_6878_n ) capacitor c=0.0146836f \
 //x=71.78 //y=2.08 //x2=71.885 //y2=5.155
cc_4203 ( N_RN_M142_noxref_g N_noxref_16_c_6878_n ) capacitor c=0.0166659f \
 //x=71.75 //y=6.02 //x2=71.885 //y2=5.155
cc_4204 ( N_RN_c_6397_n N_noxref_16_c_6878_n ) capacitor c=0.00322396f \
 //x=71.78 //y=4.7 //x2=71.885 //y2=5.155
cc_4205 ( N_RN_M143_noxref_g N_noxref_16_c_6884_n ) capacitor c=0.0184045f \
 //x=72.19 //y=6.02 //x2=72.765 //y2=5.155
cc_4206 ( N_RN_c_5921_n N_noxref_16_c_6892_n ) capacitor c=0.00296344f \
 //x=71.78 //y=2.08 //x2=73.63 //y2=4.07
cc_4207 ( N_RN_c_5920_n N_noxref_16_c_7052_n ) capacitor c=0.0174995f \
 //x=68.08 //y=2.08 //x2=68.04 //y2=5.155
cc_4208 ( N_RN_c_6366_n N_noxref_16_c_7052_n ) capacitor c=0.00475729f \
 //x=68.08 //y=4.7 //x2=68.04 //y2=5.155
cc_4209 ( N_RN_c_6404_p N_noxref_16_c_7054_n ) capacitor c=0.00427862f \
 //x=72.115 //y=4.79 //x2=71.97 //y2=5.155
cc_4210 ( N_RN_c_5887_n N_noxref_16_c_6813_n ) capacitor c=0.011987f \
 //x=59.825 //y=2.22 //x2=52.61 //y2=1.915
cc_4211 ( N_RN_c_5899_n N_noxref_16_c_7056_n ) capacitor c=3.11115e-19 \
 //x=67.965 //y=2.22 //x2=63.68 //y2=1.405
cc_4212 ( N_RN_c_5899_n N_noxref_16_c_7057_n ) capacitor c=0.00570799f \
 //x=67.965 //y=2.22 //x2=63.27 //y2=2.08
cc_4213 ( N_RN_c_6341_n N_noxref_16_M42_noxref_d ) capacitor c=0.00217566f \
 //x=68.07 //y=0.915 //x2=68.145 //y2=0.915
cc_4214 ( N_RN_c_6342_n N_noxref_16_M42_noxref_d ) capacitor c=0.0034598f \
 //x=68.07 //y=1.26 //x2=68.145 //y2=0.915
cc_4215 ( N_RN_c_6343_n N_noxref_16_M42_noxref_d ) capacitor c=0.00546784f \
 //x=68.07 //y=1.57 //x2=68.145 //y2=0.915
cc_4216 ( N_RN_c_6436_p N_noxref_16_M42_noxref_d ) capacitor c=0.00241102f \
 //x=68.445 //y=0.76 //x2=68.145 //y2=0.915
cc_4217 ( N_RN_c_6412_p N_noxref_16_M42_noxref_d ) capacitor c=0.0138621f \
 //x=68.445 //y=1.415 //x2=68.145 //y2=0.915
cc_4218 ( N_RN_c_6438_p N_noxref_16_M42_noxref_d ) capacitor c=0.00219619f \
 //x=68.6 //y=0.915 //x2=68.145 //y2=0.915
cc_4219 ( N_RN_c_6413_p N_noxref_16_M42_noxref_d ) capacitor c=0.00603828f \
 //x=68.6 //y=1.26 //x2=68.145 //y2=0.915
cc_4220 ( N_RN_c_6365_n N_noxref_16_M42_noxref_d ) capacitor c=0.00661782f \
 //x=68.08 //y=1.915 //x2=68.145 //y2=0.915
cc_4221 ( N_RN_M138_noxref_g N_noxref_16_M138_noxref_d ) capacitor \
 c=0.0180032f //x=67.82 //y=6.02 //x2=67.895 //y2=5.02
cc_4222 ( N_RN_M139_noxref_g N_noxref_16_M138_noxref_d ) capacitor \
 c=0.0194246f //x=68.26 //y=6.02 //x2=67.895 //y2=5.02
cc_4223 ( N_RN_M142_noxref_g N_noxref_16_M142_noxref_d ) capacitor \
 c=0.0180032f //x=71.75 //y=6.02 //x2=71.825 //y2=5.02
cc_4224 ( N_RN_M143_noxref_g N_noxref_16_M142_noxref_d ) capacitor \
 c=0.0180032f //x=72.19 //y=6.02 //x2=71.825 //y2=5.02
cc_4225 ( N_RN_c_5918_n N_noxref_17_c_7495_n ) capacitor c=0.00526349f \
 //x=45.88 //y=2.08 //x2=47.105 //y2=3.33
cc_4226 ( N_RN_c_5887_n N_noxref_17_c_7559_n ) capacitor c=0.0057225f \
 //x=59.825 //y=2.22 //x2=60.565 //y2=3.33
cc_4227 ( N_RN_c_5899_n N_noxref_17_c_7559_n ) capacitor c=0.00397775f \
 //x=67.965 //y=2.22 //x2=60.565 //y2=3.33
cc_4228 ( N_RN_c_5907_n N_noxref_17_c_7559_n ) capacitor c=4.86139e-19 \
 //x=60.055 //y=2.22 //x2=60.565 //y2=3.33
cc_4229 ( N_RN_c_5919_n N_noxref_17_c_7559_n ) capacitor c=0.0180187f \
 //x=59.94 //y=2.08 //x2=60.565 //y2=3.33
cc_4230 ( N_RN_c_5899_n N_noxref_17_c_7648_n ) capacitor c=0.00953758f \
 //x=67.965 //y=2.22 //x2=62.415 //y2=3.33
cc_4231 ( N_RN_c_5899_n N_noxref_17_c_7649_n ) capacitor c=4.49298e-19 \
 //x=67.965 //y=2.22 //x2=60.795 //y2=3.33
cc_4232 ( N_RN_c_5919_n N_noxref_17_c_7649_n ) capacitor c=0.00131333f \
 //x=59.94 //y=2.08 //x2=60.795 //y2=3.33
cc_4233 ( N_RN_c_5899_n N_noxref_17_c_7650_n ) capacitor c=0.00843676f \
 //x=67.965 //y=2.22 //x2=63.895 //y2=3.33
cc_4234 ( N_RN_c_5899_n N_noxref_17_c_7651_n ) capacitor c=4.44019e-19 \
 //x=67.965 //y=2.22 //x2=62.645 //y2=3.33
cc_4235 ( N_RN_c_5899_n N_noxref_17_c_7652_n ) capacitor c=0.0092367f \
 //x=67.965 //y=2.22 //x2=65.745 //y2=3.33
cc_4236 ( N_RN_c_5899_n N_noxref_17_c_7653_n ) capacitor c=4.47816e-19 \
 //x=67.965 //y=2.22 //x2=64.125 //y2=3.33
cc_4237 ( N_RN_c_5899_n N_noxref_17_c_7583_n ) capacitor c=0.0138575f \
 //x=67.965 //y=2.22 //x2=78.325 //y2=3.33
cc_4238 ( N_RN_c_5908_n N_noxref_17_c_7583_n ) capacitor c=0.0212638f \
 //x=71.665 //y=2.22 //x2=78.325 //y2=3.33
cc_4239 ( N_RN_c_5912_n N_noxref_17_c_7583_n ) capacitor c=4.86139e-19 \
 //x=68.195 //y=2.22 //x2=78.325 //y2=3.33
cc_4240 ( N_RN_c_5920_n N_noxref_17_c_7583_n ) capacitor c=0.0180187f \
 //x=68.08 //y=2.08 //x2=78.325 //y2=3.33
cc_4241 ( N_RN_c_5921_n N_noxref_17_c_7583_n ) capacitor c=0.0213922f \
 //x=71.78 //y=2.08 //x2=78.325 //y2=3.33
cc_4242 ( N_RN_c_5899_n N_noxref_17_c_7584_n ) capacitor c=4.26867e-19 \
 //x=67.965 //y=2.22 //x2=65.975 //y2=3.33
cc_4243 ( N_RN_c_5887_n N_noxref_17_c_7301_n ) capacitor c=0.0186201f \
 //x=59.825 //y=2.22 //x2=46.99 //y2=2.08
cc_4244 ( N_RN_c_5898_n N_noxref_17_c_7301_n ) capacitor c=0.00165648f \
 //x=45.995 //y=2.22 //x2=46.99 //y2=2.08
cc_4245 ( N_RN_c_5918_n N_noxref_17_c_7301_n ) capacitor c=0.044193f //x=45.88 \
 //y=2.08 //x2=46.99 //y2=2.08
cc_4246 ( N_RN_c_6157_n N_noxref_17_c_7301_n ) capacitor c=0.00205895f \
 //x=45.97 //y=1.915 //x2=46.99 //y2=2.08
cc_4247 ( N_RN_c_6159_n N_noxref_17_c_7301_n ) capacitor c=0.00142741f \
 //x=45.88 //y=4.7 //x2=46.99 //y2=2.08
cc_4248 ( N_RN_c_5887_n N_noxref_17_c_7713_n ) capacitor c=0.0146822f \
 //x=59.825 //y=2.22 //x2=50.705 //y2=1.655
cc_4249 ( N_RN_c_5887_n N_noxref_17_c_7303_n ) capacitor c=0.0199049f \
 //x=59.825 //y=2.22 //x2=51.06 //y2=3.33
cc_4250 ( N_RN_c_5887_n N_noxref_17_c_7304_n ) capacitor c=0.0186201f \
 //x=59.825 //y=2.22 //x2=55.13 //y2=2.08
cc_4251 ( N_RN_M128_noxref_g N_noxref_17_c_7391_n ) capacitor c=0.01736f \
 //x=59.68 //y=6.02 //x2=59.815 //y2=5.155
cc_4252 ( N_RN_M129_noxref_g N_noxref_17_c_7395_n ) capacitor c=0.0194981f \
 //x=60.12 //y=6.02 //x2=60.595 //y2=5.155
cc_4253 ( N_RN_c_6286_n N_noxref_17_c_7395_n ) capacitor c=0.00201851f \
 //x=59.94 //y=4.7 //x2=60.595 //y2=5.155
cc_4254 ( N_RN_c_6474_p N_noxref_17_c_7305_n ) capacitor c=0.00371277f \
 //x=60.305 //y=1.415 //x2=60.595 //y2=1.665
cc_4255 ( N_RN_c_6475_p N_noxref_17_c_7305_n ) capacitor c=0.00457401f \
 //x=60.46 //y=1.26 //x2=60.595 //y2=1.665
cc_4256 ( N_RN_c_5899_n N_noxref_17_c_7721_n ) capacitor c=0.016327f \
 //x=67.965 //y=2.22 //x2=60.28 //y2=1.665
cc_4257 ( N_RN_c_5899_n N_noxref_17_c_7399_n ) capacitor c=0.0220713f \
 //x=67.965 //y=2.22 //x2=60.68 //y2=3.33
cc_4258 ( N_RN_c_5907_n N_noxref_17_c_7399_n ) capacitor c=0.00184436f \
 //x=60.055 //y=2.22 //x2=60.68 //y2=3.33
cc_4259 ( N_RN_c_5919_n N_noxref_17_c_7399_n ) capacitor c=0.0775087f \
 //x=59.94 //y=2.08 //x2=60.68 //y2=3.33
cc_4260 ( N_RN_c_6283_n N_noxref_17_c_7399_n ) capacitor c=0.00709342f \
 //x=59.94 //y=2.08 //x2=60.68 //y2=3.33
cc_4261 ( N_RN_c_6285_n N_noxref_17_c_7399_n ) capacitor c=0.00283672f \
 //x=59.94 //y=1.915 //x2=60.68 //y2=3.33
cc_4262 ( N_RN_c_6286_n N_noxref_17_c_7399_n ) capacitor c=0.013844f //x=59.94 \
 //y=4.7 //x2=60.68 //y2=3.33
cc_4263 ( N_RN_c_5899_n N_noxref_17_c_7306_n ) capacitor c=0.0208418f \
 //x=67.965 //y=2.22 //x2=62.53 //y2=2.08
cc_4264 ( N_RN_c_5919_n N_noxref_17_c_7306_n ) capacitor c=6.23409e-19 \
 //x=59.94 //y=2.08 //x2=62.53 //y2=2.08
cc_4265 ( N_RN_c_5899_n N_noxref_17_c_7730_n ) capacitor c=0.0146822f \
 //x=67.965 //y=2.22 //x2=63.655 //y2=1.655
cc_4266 ( N_RN_c_5899_n N_noxref_17_c_7308_n ) capacitor c=0.0222456f \
 //x=67.965 //y=2.22 //x2=64.01 //y2=3.33
cc_4267 ( N_RN_c_5899_n N_noxref_17_c_7309_n ) capacitor c=0.0216101f \
 //x=67.965 //y=2.22 //x2=65.86 //y2=2.08
cc_4268 ( N_RN_c_5920_n N_noxref_17_c_7309_n ) capacitor c=0.00115753f \
 //x=68.08 //y=2.08 //x2=65.86 //y2=2.08
cc_4269 ( N_RN_c_5919_n N_noxref_17_c_7734_n ) capacitor c=0.0171303f \
 //x=59.94 //y=2.08 //x2=59.9 //y2=5.155
cc_4270 ( N_RN_c_6286_n N_noxref_17_c_7734_n ) capacitor c=0.00475601f \
 //x=59.94 //y=4.7 //x2=59.9 //y2=5.155
cc_4271 ( N_RN_M110_noxref_g N_noxref_17_M112_noxref_g ) capacitor \
 c=0.0101598f //x=45.85 //y=6.02 //x2=46.73 //y2=6.02
cc_4272 ( N_RN_M111_noxref_g N_noxref_17_M112_noxref_g ) capacitor \
 c=0.0602553f //x=46.29 //y=6.02 //x2=46.73 //y2=6.02
cc_4273 ( N_RN_M111_noxref_g N_noxref_17_M113_noxref_g ) capacitor \
 c=0.0101598f //x=46.29 //y=6.02 //x2=47.17 //y2=6.02
cc_4274 ( N_RN_c_6154_n N_noxref_17_c_7510_n ) capacitor c=0.00456962f \
 //x=45.97 //y=0.91 //x2=46.98 //y2=0.915
cc_4275 ( N_RN_c_6155_n N_noxref_17_c_7511_n ) capacitor c=0.00438372f \
 //x=45.97 //y=1.22 //x2=46.98 //y2=1.26
cc_4276 ( N_RN_c_6156_n N_noxref_17_c_7512_n ) capacitor c=0.00438372f \
 //x=45.97 //y=1.45 //x2=46.98 //y2=1.57
cc_4277 ( N_RN_c_5887_n N_noxref_17_c_7514_n ) capacitor c=3.13485e-19 \
 //x=59.825 //y=2.22 //x2=47.355 //y2=1.415
cc_4278 ( N_RN_c_5887_n N_noxref_17_c_7678_n ) capacitor c=3.13485e-19 \
 //x=59.825 //y=2.22 //x2=55.495 //y2=1.415
cc_4279 ( N_RN_c_5899_n N_noxref_17_c_7319_n ) capacitor c=0.00894156f \
 //x=67.965 //y=2.22 //x2=62.335 //y2=1.915
cc_4280 ( N_RN_c_5899_n N_noxref_17_c_7329_n ) capacitor c=0.011987f \
 //x=67.965 //y=2.22 //x2=65.56 //y2=1.915
cc_4281 ( N_RN_c_5887_n N_noxref_17_c_7519_n ) capacitor c=0.00584491f \
 //x=59.825 //y=2.22 //x2=46.99 //y2=2.08
cc_4282 ( N_RN_c_5898_n N_noxref_17_c_7519_n ) capacitor c=2.3323e-19 \
 //x=45.995 //y=2.22 //x2=46.99 //y2=2.08
cc_4283 ( N_RN_c_5918_n N_noxref_17_c_7519_n ) capacitor c=0.0019893f \
 //x=45.88 //y=2.08 //x2=46.99 //y2=2.08
cc_4284 ( N_RN_c_6157_n N_noxref_17_c_7519_n ) capacitor c=0.00828003f \
 //x=45.97 //y=1.915 //x2=46.99 //y2=2.08
cc_4285 ( N_RN_c_6157_n N_noxref_17_c_7520_n ) capacitor c=0.00438372f \
 //x=45.97 //y=1.915 //x2=46.99 //y2=1.915
cc_4286 ( N_RN_c_5918_n N_noxref_17_c_7522_n ) capacitor c=0.00219458f \
 //x=45.88 //y=2.08 //x2=46.99 //y2=4.7
cc_4287 ( N_RN_c_6172_n N_noxref_17_c_7522_n ) capacitor c=0.0611812f \
 //x=46.215 //y=4.79 //x2=46.99 //y2=4.7
cc_4288 ( N_RN_c_6159_n N_noxref_17_c_7522_n ) capacitor c=0.00487508f \
 //x=45.88 //y=4.7 //x2=46.99 //y2=4.7
cc_4289 ( N_RN_c_5887_n N_noxref_17_c_7633_n ) capacitor c=0.00584491f \
 //x=59.825 //y=2.22 //x2=55.13 //y2=2.08
cc_4290 ( N_RN_c_6268_n N_noxref_17_M37_noxref_d ) capacitor c=0.00217566f \
 //x=59.93 //y=0.915 //x2=60.005 //y2=0.915
cc_4291 ( N_RN_c_6269_n N_noxref_17_M37_noxref_d ) capacitor c=0.0034598f \
 //x=59.93 //y=1.26 //x2=60.005 //y2=0.915
cc_4292 ( N_RN_c_6270_n N_noxref_17_M37_noxref_d ) capacitor c=0.00546784f \
 //x=59.93 //y=1.57 //x2=60.005 //y2=0.915
cc_4293 ( N_RN_c_6513_p N_noxref_17_M37_noxref_d ) capacitor c=0.00241102f \
 //x=60.305 //y=0.76 //x2=60.005 //y2=0.915
cc_4294 ( N_RN_c_6474_p N_noxref_17_M37_noxref_d ) capacitor c=0.0138621f \
 //x=60.305 //y=1.415 //x2=60.005 //y2=0.915
cc_4295 ( N_RN_c_6515_p N_noxref_17_M37_noxref_d ) capacitor c=0.00219619f \
 //x=60.46 //y=0.915 //x2=60.005 //y2=0.915
cc_4296 ( N_RN_c_6475_p N_noxref_17_M37_noxref_d ) capacitor c=0.00603828f \
 //x=60.46 //y=1.26 //x2=60.005 //y2=0.915
cc_4297 ( N_RN_c_6285_n N_noxref_17_M37_noxref_d ) capacitor c=0.00661782f \
 //x=59.94 //y=1.915 //x2=60.005 //y2=0.915
cc_4298 ( N_RN_M128_noxref_g N_noxref_17_M128_noxref_d ) capacitor \
 c=0.0180032f //x=59.68 //y=6.02 //x2=59.755 //y2=5.02
cc_4299 ( N_RN_M129_noxref_g N_noxref_17_M128_noxref_d ) capacitor \
 c=0.0194246f //x=60.12 //y=6.02 //x2=59.755 //y2=5.02
cc_4300 ( N_RN_c_5921_n N_noxref_18_c_8127_n ) capacitor c=0.0027353f \
 //x=71.78 //y=2.08 //x2=73.005 //y2=3.7
cc_4301 ( N_RN_c_5908_n N_noxref_18_c_8065_n ) capacitor c=0.00558344f \
 //x=71.665 //y=2.22 //x2=72.89 //y2=2.08
cc_4302 ( N_RN_c_5921_n N_noxref_18_c_8065_n ) capacitor c=0.0482297f \
 //x=71.78 //y=2.08 //x2=72.89 //y2=2.08
cc_4303 ( N_RN_c_6395_n N_noxref_18_c_8065_n ) capacitor c=0.00213841f \
 //x=71.87 //y=1.915 //x2=72.89 //y2=2.08
cc_4304 ( N_RN_c_6397_n N_noxref_18_c_8065_n ) capacitor c=0.00142741f \
 //x=71.78 //y=4.7 //x2=72.89 //y2=2.08
cc_4305 ( N_RN_M142_noxref_g N_noxref_18_M144_noxref_g ) capacitor \
 c=0.0101598f //x=71.75 //y=6.02 //x2=72.63 //y2=6.02
cc_4306 ( N_RN_M143_noxref_g N_noxref_18_M144_noxref_g ) capacitor \
 c=0.0602553f //x=72.19 //y=6.02 //x2=72.63 //y2=6.02
cc_4307 ( N_RN_M143_noxref_g N_noxref_18_M145_noxref_g ) capacitor \
 c=0.0101598f //x=72.19 //y=6.02 //x2=73.07 //y2=6.02
cc_4308 ( N_RN_c_6392_n N_noxref_18_c_8137_n ) capacitor c=0.00456962f \
 //x=71.87 //y=0.91 //x2=72.88 //y2=0.915
cc_4309 ( N_RN_c_6393_n N_noxref_18_c_8138_n ) capacitor c=0.00438372f \
 //x=71.87 //y=1.22 //x2=72.88 //y2=1.26
cc_4310 ( N_RN_c_6394_n N_noxref_18_c_8139_n ) capacitor c=0.00438372f \
 //x=71.87 //y=1.45 //x2=72.88 //y2=1.57
cc_4311 ( N_RN_c_5908_n N_noxref_18_c_8140_n ) capacitor c=0.00341397f \
 //x=71.665 //y=2.22 //x2=72.89 //y2=2.08
cc_4312 ( N_RN_c_5921_n N_noxref_18_c_8140_n ) capacitor c=0.0021852f \
 //x=71.78 //y=2.08 //x2=72.89 //y2=2.08
cc_4313 ( N_RN_c_6395_n N_noxref_18_c_8140_n ) capacitor c=0.00896806f \
 //x=71.87 //y=1.915 //x2=72.89 //y2=2.08
cc_4314 ( N_RN_c_6395_n N_noxref_18_c_8143_n ) capacitor c=0.00438372f \
 //x=71.87 //y=1.915 //x2=72.89 //y2=1.915
cc_4315 ( N_RN_c_5921_n N_noxref_18_c_8144_n ) capacitor c=0.00219458f \
 //x=71.78 //y=2.08 //x2=72.89 //y2=4.7
cc_4316 ( N_RN_c_6404_p N_noxref_18_c_8144_n ) capacitor c=0.0611812f \
 //x=72.115 //y=4.79 //x2=72.89 //y2=4.7
cc_4317 ( N_RN_c_6397_n N_noxref_18_c_8144_n ) capacitor c=0.00487508f \
 //x=71.78 //y=4.7 //x2=72.89 //y2=4.7
cc_4318 ( N_RN_c_5861_n N_noxref_20_c_8515_n ) capacitor c=0.0293706f \
 //x=33.925 //y=2.22 //x2=25.045 //y2=2.96
cc_4319 ( N_RN_c_5861_n N_noxref_20_c_8606_n ) capacitor c=9.7414e-19 \
 //x=33.925 //y=2.22 //x2=21.205 //y2=2.96
cc_4320 ( N_RN_c_5915_n N_noxref_20_c_8606_n ) capacitor c=0.00526349f \
 //x=19.98 //y=2.08 //x2=21.205 //y2=2.96
cc_4321 ( N_RN_c_5861_n N_noxref_20_c_8516_n ) capacitor c=0.0666921f \
 //x=33.925 //y=2.22 //x2=83.505 //y2=2.96
cc_4322 ( N_RN_c_5873_n N_noxref_20_c_8516_n ) capacitor c=0.0599768f \
 //x=42.065 //y=2.22 //x2=83.505 //y2=2.96
cc_4323 ( N_RN_c_5881_n N_noxref_20_c_8516_n ) capacitor c=6.59215e-19 \
 //x=34.155 //y=2.22 //x2=83.505 //y2=2.96
cc_4324 ( N_RN_c_5882_n N_noxref_20_c_8516_n ) capacitor c=0.0260426f \
 //x=45.765 //y=2.22 //x2=83.505 //y2=2.96
cc_4325 ( N_RN_c_5886_n N_noxref_20_c_8516_n ) capacitor c=6.59215e-19 \
 //x=42.295 //y=2.22 //x2=83.505 //y2=2.96
cc_4326 ( N_RN_c_5887_n N_noxref_20_c_8516_n ) capacitor c=0.129549f \
 //x=59.825 //y=2.22 //x2=83.505 //y2=2.96
cc_4327 ( N_RN_c_5898_n N_noxref_20_c_8516_n ) capacitor c=6.59215e-19 \
 //x=45.995 //y=2.22 //x2=83.505 //y2=2.96
cc_4328 ( N_RN_c_5899_n N_noxref_20_c_8516_n ) capacitor c=0.332655f \
 //x=67.965 //y=2.22 //x2=83.505 //y2=2.96
cc_4329 ( N_RN_c_5907_n N_noxref_20_c_8516_n ) capacitor c=0.0120222f \
 //x=60.055 //y=2.22 //x2=83.505 //y2=2.96
cc_4330 ( N_RN_c_5908_n N_noxref_20_c_8516_n ) capacitor c=0.16049f //x=71.665 \
 //y=2.22 //x2=83.505 //y2=2.96
cc_4331 ( N_RN_c_5912_n N_noxref_20_c_8516_n ) capacitor c=0.0120222f \
 //x=68.195 //y=2.22 //x2=83.505 //y2=2.96
cc_4332 ( N_RN_c_5916_n N_noxref_20_c_8516_n ) capacitor c=0.0179917f \
 //x=34.04 //y=2.08 //x2=83.505 //y2=2.96
cc_4333 ( N_RN_c_5917_n N_noxref_20_c_8516_n ) capacitor c=0.0203312f \
 //x=42.18 //y=2.08 //x2=83.505 //y2=2.96
cc_4334 ( N_RN_c_5918_n N_noxref_20_c_8516_n ) capacitor c=0.0228892f \
 //x=45.88 //y=2.08 //x2=83.505 //y2=2.96
cc_4335 ( N_RN_c_5919_n N_noxref_20_c_8516_n ) capacitor c=0.0206071f \
 //x=59.94 //y=2.08 //x2=83.505 //y2=2.96
cc_4336 ( N_RN_c_5920_n N_noxref_20_c_8516_n ) capacitor c=0.0206071f \
 //x=68.08 //y=2.08 //x2=83.505 //y2=2.96
cc_4337 ( N_RN_c_5921_n N_noxref_20_c_8516_n ) capacitor c=0.0216476f \
 //x=71.78 //y=2.08 //x2=83.505 //y2=2.96
cc_4338 ( N_RN_c_6395_n N_noxref_20_c_8516_n ) capacitor c=4.10467e-19 \
 //x=71.87 //y=1.915 //x2=83.505 //y2=2.96
cc_4339 ( N_RN_c_5861_n N_noxref_20_c_8608_n ) capacitor c=5.71765e-19 \
 //x=33.925 //y=2.22 //x2=25.275 //y2=2.96
cc_4340 ( N_RN_c_5861_n N_noxref_20_c_8538_n ) capacitor c=0.0186201f \
 //x=33.925 //y=2.22 //x2=21.09 //y2=2.08
cc_4341 ( N_RN_c_5872_n N_noxref_20_c_8538_n ) capacitor c=0.00165648f \
 //x=20.095 //y=2.22 //x2=21.09 //y2=2.08
cc_4342 ( N_RN_c_5915_n N_noxref_20_c_8538_n ) capacitor c=0.046799f //x=19.98 \
 //y=2.08 //x2=21.09 //y2=2.08
cc_4343 ( N_RN_c_6037_n N_noxref_20_c_8538_n ) capacitor c=0.00205895f \
 //x=20.07 //y=1.915 //x2=21.09 //y2=2.08
cc_4344 ( N_RN_c_6039_n N_noxref_20_c_8538_n ) capacitor c=0.00142741f \
 //x=19.98 //y=4.7 //x2=21.09 //y2=2.08
cc_4345 ( N_RN_c_5861_n N_noxref_20_c_8761_n ) capacitor c=0.0146822f \
 //x=33.925 //y=2.22 //x2=24.805 //y2=1.655
cc_4346 ( N_RN_c_5861_n N_noxref_20_c_8540_n ) capacitor c=0.0199049f \
 //x=33.925 //y=2.22 //x2=25.16 //y2=2.96
cc_4347 ( N_RN_M78_noxref_g N_noxref_20_M80_noxref_g ) capacitor c=0.0101598f \
 //x=19.95 //y=6.02 //x2=20.83 //y2=6.02
cc_4348 ( N_RN_M79_noxref_g N_noxref_20_M80_noxref_g ) capacitor c=0.0602553f \
 //x=20.39 //y=6.02 //x2=20.83 //y2=6.02
cc_4349 ( N_RN_M79_noxref_g N_noxref_20_M81_noxref_g ) capacitor c=0.0101598f \
 //x=20.39 //y=6.02 //x2=21.27 //y2=6.02
cc_4350 ( N_RN_c_6034_n N_noxref_20_c_8638_n ) capacitor c=0.00456962f \
 //x=20.07 //y=0.91 //x2=21.08 //y2=0.915
cc_4351 ( N_RN_c_6035_n N_noxref_20_c_8639_n ) capacitor c=0.00438372f \
 //x=20.07 //y=1.22 //x2=21.08 //y2=1.26
cc_4352 ( N_RN_c_6036_n N_noxref_20_c_8640_n ) capacitor c=0.00438372f \
 //x=20.07 //y=1.45 //x2=21.08 //y2=1.57
cc_4353 ( N_RN_c_5861_n N_noxref_20_c_8642_n ) capacitor c=3.13485e-19 \
 //x=33.925 //y=2.22 //x2=21.455 //y2=1.415
cc_4354 ( N_RN_c_5861_n N_noxref_20_c_8647_n ) capacitor c=0.00584491f \
 //x=33.925 //y=2.22 //x2=21.09 //y2=2.08
cc_4355 ( N_RN_c_5872_n N_noxref_20_c_8647_n ) capacitor c=2.3323e-19 \
 //x=20.095 //y=2.22 //x2=21.09 //y2=2.08
cc_4356 ( N_RN_c_5915_n N_noxref_20_c_8647_n ) capacitor c=0.0019893f \
 //x=19.98 //y=2.08 //x2=21.09 //y2=2.08
cc_4357 ( N_RN_c_6037_n N_noxref_20_c_8647_n ) capacitor c=0.00828003f \
 //x=20.07 //y=1.915 //x2=21.09 //y2=2.08
cc_4358 ( N_RN_c_6037_n N_noxref_20_c_8648_n ) capacitor c=0.00438372f \
 //x=20.07 //y=1.915 //x2=21.09 //y2=1.915
cc_4359 ( N_RN_c_5915_n N_noxref_20_c_8650_n ) capacitor c=0.00219458f \
 //x=19.98 //y=2.08 //x2=21.09 //y2=4.7
cc_4360 ( N_RN_c_6084_n N_noxref_20_c_8650_n ) capacitor c=0.0611812f \
 //x=20.315 //y=4.79 //x2=21.09 //y2=4.7
cc_4361 ( N_RN_c_6039_n N_noxref_20_c_8650_n ) capacitor c=0.00487508f \
 //x=19.98 //y=4.7 //x2=21.09 //y2=4.7
cc_4362 ( N_RN_c_5846_n N_noxref_26_c_9421_n ) capacitor c=7.41833e-19 \
 //x=16.165 //y=2.22 //x2=8.795 //y2=0.54
cc_4363 ( N_RN_c_5854_n N_noxref_26_c_9421_n ) capacitor c=7.4531e-19 \
 //x=8.255 //y=2.22 //x2=8.795 //y2=0.54
cc_4364 ( N_RN_c_5913_n N_noxref_26_c_9421_n ) capacitor c=0.00204178f \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_4365 ( N_RN_c_5988_n N_noxref_26_c_9421_n ) capacitor c=0.0194423f //x=8.13 \
 //y=0.915 //x2=8.795 //y2=0.54
cc_4366 ( N_RN_c_5994_n N_noxref_26_c_9421_n ) capacitor c=0.00656458f \
 //x=8.66 //y=0.915 //x2=8.795 //y2=0.54
cc_4367 ( N_RN_c_5997_n N_noxref_26_c_9421_n ) capacitor c=2.20712e-19 \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_4368 ( N_RN_c_5989_n N_noxref_26_c_9431_n ) capacitor c=0.00538829f \
 //x=8.13 //y=1.26 //x2=7.91 //y2=0.995
cc_4369 ( N_RN_c_5988_n N_noxref_26_M5_noxref_s ) capacitor c=0.00538829f \
 //x=8.13 //y=0.915 //x2=7.775 //y2=0.375
cc_4370 ( N_RN_c_5990_n N_noxref_26_M5_noxref_s ) capacitor c=0.00538829f \
 //x=8.13 //y=1.57 //x2=7.775 //y2=0.375
cc_4371 ( N_RN_c_5994_n N_noxref_26_M5_noxref_s ) capacitor c=0.0143002f \
 //x=8.66 //y=0.915 //x2=7.775 //y2=0.375
cc_4372 ( N_RN_c_5995_n N_noxref_26_M5_noxref_s ) capacitor c=0.00290153f \
 //x=8.66 //y=1.26 //x2=7.775 //y2=0.375
cc_4373 ( N_RN_c_5846_n N_noxref_27_c_9487_n ) capacitor c=0.00635755f \
 //x=16.165 //y=2.22 //x2=10.315 //y2=1.495
cc_4374 ( N_RN_c_5846_n N_noxref_27_c_9469_n ) capacitor c=0.0223494f \
 //x=16.165 //y=2.22 //x2=11.2 //y2=1.58
cc_4375 ( N_RN_c_5846_n N_noxref_27_c_9476_n ) capacitor c=0.00649228f \
 //x=16.165 //y=2.22 //x2=11.285 //y2=1.495
cc_4376 ( N_RN_c_5846_n N_noxref_27_c_9477_n ) capacitor c=0.00178534f \
 //x=16.165 //y=2.22 //x2=12.17 //y2=0.53
cc_4377 ( N_RN_c_5846_n N_noxref_27_M6_noxref_s ) capacitor c=0.00113237f \
 //x=16.165 //y=2.22 //x2=10.18 //y2=0.365
cc_4378 ( N_RN_c_5846_n N_noxref_28_c_9535_n ) capacitor c=0.00642985f \
 //x=16.165 //y=2.22 //x2=13.54 //y2=1.505
cc_4379 ( N_RN_c_5846_n N_noxref_28_c_9520_n ) capacitor c=0.0225733f \
 //x=16.165 //y=2.22 //x2=14.425 //y2=1.59
cc_4380 ( N_RN_c_5846_n N_noxref_28_c_9550_n ) capacitor c=0.0203655f \
 //x=16.165 //y=2.22 //x2=15.395 //y2=1.59
cc_4381 ( N_RN_c_5846_n N_noxref_28_M8_noxref_s ) capacitor c=0.012425f \
 //x=16.165 //y=2.22 //x2=13.405 //y2=0.375
cc_4382 ( N_RN_c_5846_n N_noxref_29_c_9569_n ) capacitor c=0.00657782f \
 //x=16.165 //y=2.22 //x2=15.965 //y2=0.995
cc_4383 ( N_RN_c_5856_n N_noxref_29_c_9574_n ) capacitor c=7.41833e-19 \
 //x=19.865 //y=2.22 //x2=16.935 //y2=0.54
cc_4384 ( N_RN_c_5860_n N_noxref_29_c_9574_n ) capacitor c=7.4531e-19 \
 //x=16.395 //y=2.22 //x2=16.935 //y2=0.54
cc_4385 ( N_RN_c_5914_n N_noxref_29_c_9574_n ) capacitor c=0.00204178f \
 //x=16.28 //y=2.08 //x2=16.935 //y2=0.54
cc_4386 ( N_RN_c_6075_n N_noxref_29_c_9574_n ) capacitor c=0.0194423f \
 //x=16.27 //y=0.915 //x2=16.935 //y2=0.54
cc_4387 ( N_RN_c_6081_n N_noxref_29_c_9574_n ) capacitor c=0.00656458f \
 //x=16.8 //y=0.915 //x2=16.935 //y2=0.54
cc_4388 ( N_RN_c_6085_n N_noxref_29_c_9574_n ) capacitor c=2.20712e-19 \
 //x=16.28 //y=2.08 //x2=16.935 //y2=0.54
cc_4389 ( N_RN_c_6076_n N_noxref_29_c_9584_n ) capacitor c=0.00538829f \
 //x=16.27 //y=1.26 //x2=16.05 //y2=0.995
cc_4390 ( N_RN_c_5846_n N_noxref_29_M10_noxref_s ) capacitor c=0.00642985f \
 //x=16.165 //y=2.22 //x2=15.915 //y2=0.375
cc_4391 ( N_RN_c_6075_n N_noxref_29_M10_noxref_s ) capacitor c=0.00538829f \
 //x=16.27 //y=0.915 //x2=15.915 //y2=0.375
cc_4392 ( N_RN_c_6077_n N_noxref_29_M10_noxref_s ) capacitor c=0.00538829f \
 //x=16.27 //y=1.57 //x2=15.915 //y2=0.375
cc_4393 ( N_RN_c_6081_n N_noxref_29_M10_noxref_s ) capacitor c=0.0143002f \
 //x=16.8 //y=0.915 //x2=15.915 //y2=0.375
cc_4394 ( N_RN_c_6082_n N_noxref_29_M10_noxref_s ) capacitor c=0.00290153f \
 //x=16.8 //y=1.26 //x2=15.915 //y2=0.375
cc_4395 ( N_RN_c_5856_n N_noxref_30_c_9637_n ) capacitor c=0.00642985f \
 //x=19.865 //y=2.22 //x2=18.35 //y2=1.505
cc_4396 ( N_RN_c_5856_n N_noxref_30_c_9622_n ) capacitor c=0.0225733f \
 //x=19.865 //y=2.22 //x2=19.235 //y2=1.59
cc_4397 ( N_RN_c_6029_n N_noxref_30_c_9629_n ) capacitor c=0.0167228f \
 //x=19.545 //y=0.91 //x2=20.205 //y2=0.54
cc_4398 ( N_RN_c_6034_n N_noxref_30_c_9629_n ) capacitor c=0.00534519f \
 //x=20.07 //y=0.91 //x2=20.205 //y2=0.54
cc_4399 ( N_RN_c_5856_n N_noxref_30_c_9654_n ) capacitor c=0.0139868f \
 //x=19.865 //y=2.22 //x2=20.205 //y2=1.59
cc_4400 ( N_RN_c_5861_n N_noxref_30_c_9654_n ) capacitor c=0.00387656f \
 //x=33.925 //y=2.22 //x2=20.205 //y2=1.59
cc_4401 ( N_RN_c_5872_n N_noxref_30_c_9654_n ) capacitor c=0.00251375f \
 //x=20.095 //y=2.22 //x2=20.205 //y2=1.59
cc_4402 ( N_RN_c_5915_n N_noxref_30_c_9654_n ) capacitor c=0.0119919f \
 //x=19.98 //y=2.08 //x2=20.205 //y2=1.59
cc_4403 ( N_RN_c_6032_n N_noxref_30_c_9654_n ) capacitor c=0.0157358f \
 //x=19.545 //y=1.22 //x2=20.205 //y2=1.59
cc_4404 ( N_RN_c_6037_n N_noxref_30_c_9654_n ) capacitor c=0.0213278f \
 //x=20.07 //y=1.915 //x2=20.205 //y2=1.59
cc_4405 ( N_RN_c_5856_n N_noxref_30_M11_noxref_s ) capacitor c=0.00642985f \
 //x=19.865 //y=2.22 //x2=18.215 //y2=0.375
cc_4406 ( N_RN_c_5861_n N_noxref_30_M11_noxref_s ) capacitor c=0.00599513f \
 //x=33.925 //y=2.22 //x2=18.215 //y2=0.375
cc_4407 ( N_RN_c_6029_n N_noxref_30_M11_noxref_s ) capacitor c=0.00798959f \
 //x=19.545 //y=0.91 //x2=18.215 //y2=0.375
cc_4408 ( N_RN_c_6036_n N_noxref_30_M11_noxref_s ) capacitor c=0.00212176f \
 //x=20.07 //y=1.45 //x2=18.215 //y2=0.375
cc_4409 ( N_RN_c_6037_n N_noxref_30_M11_noxref_s ) capacitor c=0.00298115f \
 //x=20.07 //y=1.915 //x2=18.215 //y2=0.375
cc_4410 ( N_RN_c_5861_n N_noxref_31_c_9674_n ) capacitor c=0.00657782f \
 //x=33.925 //y=2.22 //x2=20.775 //y2=0.995
cc_4411 ( N_RN_c_6631_p N_noxref_31_c_9674_n ) capacitor c=2.14837e-19 \
 //x=19.915 //y=0.755 //x2=20.775 //y2=0.995
cc_4412 ( N_RN_c_6034_n N_noxref_31_c_9674_n ) capacitor c=0.00123426f \
 //x=20.07 //y=0.91 //x2=20.775 //y2=0.995
cc_4413 ( N_RN_c_6035_n N_noxref_31_c_9674_n ) capacitor c=0.0129288f \
 //x=20.07 //y=1.22 //x2=20.775 //y2=0.995
cc_4414 ( N_RN_c_6036_n N_noxref_31_c_9674_n ) capacitor c=0.00142359f \
 //x=20.07 //y=1.45 //x2=20.775 //y2=0.995
cc_4415 ( N_RN_c_5861_n N_noxref_31_c_9679_n ) capacitor c=0.00147946f \
 //x=33.925 //y=2.22 //x2=21.745 //y2=0.54
cc_4416 ( N_RN_c_6029_n N_noxref_31_M12_noxref_d ) capacitor c=0.00223875f \
 //x=19.545 //y=0.91 //x2=19.62 //y2=0.91
cc_4417 ( N_RN_c_6032_n N_noxref_31_M12_noxref_d ) capacitor c=0.00262485f \
 //x=19.545 //y=1.22 //x2=19.62 //y2=0.91
cc_4418 ( N_RN_c_6631_p N_noxref_31_M12_noxref_d ) capacitor c=0.00220746f \
 //x=19.915 //y=0.755 //x2=19.62 //y2=0.91
cc_4419 ( N_RN_c_6639_p N_noxref_31_M12_noxref_d ) capacitor c=0.00194798f \
 //x=19.915 //y=1.375 //x2=19.62 //y2=0.91
cc_4420 ( N_RN_c_6034_n N_noxref_31_M12_noxref_d ) capacitor c=0.00198465f \
 //x=20.07 //y=0.91 //x2=19.62 //y2=0.91
cc_4421 ( N_RN_c_6035_n N_noxref_31_M12_noxref_d ) capacitor c=0.00128384f \
 //x=20.07 //y=1.22 //x2=19.62 //y2=0.91
cc_4422 ( N_RN_c_5861_n N_noxref_31_M13_noxref_s ) capacitor c=0.00642985f \
 //x=33.925 //y=2.22 //x2=20.725 //y2=0.375
cc_4423 ( N_RN_c_6034_n N_noxref_31_M13_noxref_s ) capacitor c=7.21316e-19 \
 //x=20.07 //y=0.91 //x2=20.725 //y2=0.375
cc_4424 ( N_RN_c_6035_n N_noxref_31_M13_noxref_s ) capacitor c=0.00348171f \
 //x=20.07 //y=1.22 //x2=20.725 //y2=0.375
cc_4425 ( N_RN_c_5861_n N_noxref_32_c_9744_n ) capacitor c=0.00635755f \
 //x=33.925 //y=2.22 //x2=23.265 //y2=1.495
cc_4426 ( N_RN_c_5861_n N_noxref_32_c_9726_n ) capacitor c=0.0223494f \
 //x=33.925 //y=2.22 //x2=24.15 //y2=1.58
cc_4427 ( N_RN_c_5861_n N_noxref_32_c_9733_n ) capacitor c=0.00649228f \
 //x=33.925 //y=2.22 //x2=24.235 //y2=1.495
cc_4428 ( N_RN_c_5861_n N_noxref_32_c_9734_n ) capacitor c=0.00178534f \
 //x=33.925 //y=2.22 //x2=25.12 //y2=0.53
cc_4429 ( N_RN_c_5861_n N_noxref_32_M14_noxref_s ) capacitor c=0.00113237f \
 //x=33.925 //y=2.22 //x2=23.13 //y2=0.365
cc_4430 ( N_RN_c_5861_n N_noxref_33_c_9793_n ) capacitor c=0.00642985f \
 //x=33.925 //y=2.22 //x2=26.49 //y2=1.505
cc_4431 ( N_RN_c_5861_n N_noxref_33_c_9777_n ) capacitor c=0.0225733f \
 //x=33.925 //y=2.22 //x2=27.375 //y2=1.59
cc_4432 ( N_RN_c_5861_n N_noxref_33_c_9805_n ) capacitor c=0.0203655f \
 //x=33.925 //y=2.22 //x2=28.345 //y2=1.59
cc_4433 ( N_RN_c_5861_n N_noxref_33_M16_noxref_s ) capacitor c=0.012425f \
 //x=33.925 //y=2.22 //x2=26.355 //y2=0.375
cc_4434 ( N_RN_c_5861_n N_noxref_34_c_9826_n ) capacitor c=0.00657782f \
 //x=33.925 //y=2.22 //x2=28.915 //y2=0.995
cc_4435 ( N_RN_c_5861_n N_noxref_34_c_9831_n ) capacitor c=0.00147946f \
 //x=33.925 //y=2.22 //x2=29.885 //y2=0.54
cc_4436 ( N_RN_c_5861_n N_noxref_34_M18_noxref_s ) capacitor c=0.00642985f \
 //x=33.925 //y=2.22 //x2=28.865 //y2=0.375
cc_4437 ( N_RN_c_5861_n N_noxref_35_c_9894_n ) capacitor c=0.00642985f \
 //x=33.925 //y=2.22 //x2=31.3 //y2=1.505
cc_4438 ( N_RN_c_5861_n N_noxref_35_c_9878_n ) capacitor c=0.0225733f \
 //x=33.925 //y=2.22 //x2=32.185 //y2=1.59
cc_4439 ( N_RN_c_5861_n N_noxref_35_c_9908_n ) capacitor c=0.0203655f \
 //x=33.925 //y=2.22 //x2=33.155 //y2=1.59
cc_4440 ( N_RN_c_5861_n N_noxref_35_M19_noxref_s ) capacitor c=0.012425f \
 //x=33.925 //y=2.22 //x2=31.165 //y2=0.375
cc_4441 ( N_RN_c_5861_n N_noxref_36_c_9927_n ) capacitor c=0.00657782f \
 //x=33.925 //y=2.22 //x2=33.725 //y2=0.995
cc_4442 ( N_RN_c_5873_n N_noxref_36_c_9932_n ) capacitor c=7.41833e-19 \
 //x=42.065 //y=2.22 //x2=34.695 //y2=0.54
cc_4443 ( N_RN_c_5881_n N_noxref_36_c_9932_n ) capacitor c=7.4531e-19 \
 //x=34.155 //y=2.22 //x2=34.695 //y2=0.54
cc_4444 ( N_RN_c_5916_n N_noxref_36_c_9932_n ) capacitor c=0.00204178f \
 //x=34.04 //y=2.08 //x2=34.695 //y2=0.54
cc_4445 ( N_RN_c_6109_n N_noxref_36_c_9932_n ) capacitor c=0.0194423f \
 //x=34.03 //y=0.915 //x2=34.695 //y2=0.54
cc_4446 ( N_RN_c_6115_n N_noxref_36_c_9932_n ) capacitor c=0.00656458f \
 //x=34.56 //y=0.915 //x2=34.695 //y2=0.54
cc_4447 ( N_RN_c_6118_n N_noxref_36_c_9932_n ) capacitor c=2.20712e-19 \
 //x=34.04 //y=2.08 //x2=34.695 //y2=0.54
cc_4448 ( N_RN_c_6110_n N_noxref_36_c_9942_n ) capacitor c=0.00538829f \
 //x=34.03 //y=1.26 //x2=33.81 //y2=0.995
cc_4449 ( N_RN_c_5861_n N_noxref_36_M21_noxref_s ) capacitor c=0.00642985f \
 //x=33.925 //y=2.22 //x2=33.675 //y2=0.375
cc_4450 ( N_RN_c_6109_n N_noxref_36_M21_noxref_s ) capacitor c=0.00538829f \
 //x=34.03 //y=0.915 //x2=33.675 //y2=0.375
cc_4451 ( N_RN_c_6111_n N_noxref_36_M21_noxref_s ) capacitor c=0.00538829f \
 //x=34.03 //y=1.57 //x2=33.675 //y2=0.375
cc_4452 ( N_RN_c_6115_n N_noxref_36_M21_noxref_s ) capacitor c=0.0143002f \
 //x=34.56 //y=0.915 //x2=33.675 //y2=0.375
cc_4453 ( N_RN_c_6116_n N_noxref_36_M21_noxref_s ) capacitor c=0.00290153f \
 //x=34.56 //y=1.26 //x2=33.675 //y2=0.375
cc_4454 ( N_RN_c_5873_n N_noxref_37_c_9998_n ) capacitor c=0.00635755f \
 //x=42.065 //y=2.22 //x2=36.215 //y2=1.495
cc_4455 ( N_RN_c_5873_n N_noxref_37_c_9980_n ) capacitor c=0.0223494f \
 //x=42.065 //y=2.22 //x2=37.1 //y2=1.58
cc_4456 ( N_RN_c_5873_n N_noxref_37_c_9987_n ) capacitor c=0.00649228f \
 //x=42.065 //y=2.22 //x2=37.185 //y2=1.495
cc_4457 ( N_RN_c_5873_n N_noxref_37_c_9988_n ) capacitor c=0.00178534f \
 //x=42.065 //y=2.22 //x2=38.07 //y2=0.53
cc_4458 ( N_RN_c_5873_n N_noxref_37_M22_noxref_s ) capacitor c=0.00113237f \
 //x=42.065 //y=2.22 //x2=36.08 //y2=0.365
cc_4459 ( N_RN_c_5873_n N_noxref_38_c_10046_n ) capacitor c=0.00642985f \
 //x=42.065 //y=2.22 //x2=39.44 //y2=1.505
cc_4460 ( N_RN_c_5873_n N_noxref_38_c_10031_n ) capacitor c=0.0225733f \
 //x=42.065 //y=2.22 //x2=40.325 //y2=1.59
cc_4461 ( N_RN_c_5873_n N_noxref_38_c_10061_n ) capacitor c=0.0203655f \
 //x=42.065 //y=2.22 //x2=41.295 //y2=1.59
cc_4462 ( N_RN_c_5873_n N_noxref_38_M24_noxref_s ) capacitor c=0.012425f \
 //x=42.065 //y=2.22 //x2=39.305 //y2=0.375
cc_4463 ( N_RN_c_5873_n N_noxref_39_c_10080_n ) capacitor c=0.00657782f \
 //x=42.065 //y=2.22 //x2=41.865 //y2=0.995
cc_4464 ( N_RN_c_5882_n N_noxref_39_c_10085_n ) capacitor c=7.41833e-19 \
 //x=45.765 //y=2.22 //x2=42.835 //y2=0.54
cc_4465 ( N_RN_c_5886_n N_noxref_39_c_10085_n ) capacitor c=7.4531e-19 \
 //x=42.295 //y=2.22 //x2=42.835 //y2=0.54
cc_4466 ( N_RN_c_5917_n N_noxref_39_c_10085_n ) capacitor c=0.00204178f \
 //x=42.18 //y=2.08 //x2=42.835 //y2=0.54
cc_4467 ( N_RN_c_6196_n N_noxref_39_c_10085_n ) capacitor c=0.0194423f \
 //x=42.17 //y=0.915 //x2=42.835 //y2=0.54
cc_4468 ( N_RN_c_6202_n N_noxref_39_c_10085_n ) capacitor c=0.00656458f \
 //x=42.7 //y=0.915 //x2=42.835 //y2=0.54
cc_4469 ( N_RN_c_6205_n N_noxref_39_c_10085_n ) capacitor c=2.20712e-19 \
 //x=42.18 //y=2.08 //x2=42.835 //y2=0.54
cc_4470 ( N_RN_c_6197_n N_noxref_39_c_10095_n ) capacitor c=0.00538829f \
 //x=42.17 //y=1.26 //x2=41.95 //y2=0.995
cc_4471 ( N_RN_c_5873_n N_noxref_39_M26_noxref_s ) capacitor c=0.00642985f \
 //x=42.065 //y=2.22 //x2=41.815 //y2=0.375
cc_4472 ( N_RN_c_6196_n N_noxref_39_M26_noxref_s ) capacitor c=0.00538829f \
 //x=42.17 //y=0.915 //x2=41.815 //y2=0.375
cc_4473 ( N_RN_c_6198_n N_noxref_39_M26_noxref_s ) capacitor c=0.00538829f \
 //x=42.17 //y=1.57 //x2=41.815 //y2=0.375
cc_4474 ( N_RN_c_6202_n N_noxref_39_M26_noxref_s ) capacitor c=0.0143002f \
 //x=42.7 //y=0.915 //x2=41.815 //y2=0.375
cc_4475 ( N_RN_c_6203_n N_noxref_39_M26_noxref_s ) capacitor c=0.00290153f \
 //x=42.7 //y=1.26 //x2=41.815 //y2=0.375
cc_4476 ( N_RN_c_5882_n N_noxref_40_c_10148_n ) capacitor c=0.00642985f \
 //x=45.765 //y=2.22 //x2=44.25 //y2=1.505
cc_4477 ( N_RN_c_5882_n N_noxref_40_c_10133_n ) capacitor c=0.0225733f \
 //x=45.765 //y=2.22 //x2=45.135 //y2=1.59
cc_4478 ( N_RN_c_6149_n N_noxref_40_c_10140_n ) capacitor c=0.0167228f \
 //x=45.445 //y=0.91 //x2=46.105 //y2=0.54
cc_4479 ( N_RN_c_6154_n N_noxref_40_c_10140_n ) capacitor c=0.00534519f \
 //x=45.97 //y=0.91 //x2=46.105 //y2=0.54
cc_4480 ( N_RN_c_5882_n N_noxref_40_c_10165_n ) capacitor c=0.0139868f \
 //x=45.765 //y=2.22 //x2=46.105 //y2=1.59
cc_4481 ( N_RN_c_5887_n N_noxref_40_c_10165_n ) capacitor c=0.00387656f \
 //x=59.825 //y=2.22 //x2=46.105 //y2=1.59
cc_4482 ( N_RN_c_5898_n N_noxref_40_c_10165_n ) capacitor c=0.00251375f \
 //x=45.995 //y=2.22 //x2=46.105 //y2=1.59
cc_4483 ( N_RN_c_5918_n N_noxref_40_c_10165_n ) capacitor c=0.011736f \
 //x=45.88 //y=2.08 //x2=46.105 //y2=1.59
cc_4484 ( N_RN_c_6152_n N_noxref_40_c_10165_n ) capacitor c=0.0157358f \
 //x=45.445 //y=1.22 //x2=46.105 //y2=1.59
cc_4485 ( N_RN_c_6157_n N_noxref_40_c_10165_n ) capacitor c=0.0213278f \
 //x=45.97 //y=1.915 //x2=46.105 //y2=1.59
cc_4486 ( N_RN_c_5882_n N_noxref_40_M27_noxref_s ) capacitor c=0.00642985f \
 //x=45.765 //y=2.22 //x2=44.115 //y2=0.375
cc_4487 ( N_RN_c_5887_n N_noxref_40_M27_noxref_s ) capacitor c=0.00599513f \
 //x=59.825 //y=2.22 //x2=44.115 //y2=0.375
cc_4488 ( N_RN_c_6149_n N_noxref_40_M27_noxref_s ) capacitor c=0.00798959f \
 //x=45.445 //y=0.91 //x2=44.115 //y2=0.375
cc_4489 ( N_RN_c_6156_n N_noxref_40_M27_noxref_s ) capacitor c=0.00212176f \
 //x=45.97 //y=1.45 //x2=44.115 //y2=0.375
cc_4490 ( N_RN_c_6157_n N_noxref_40_M27_noxref_s ) capacitor c=0.00298115f \
 //x=45.97 //y=1.915 //x2=44.115 //y2=0.375
cc_4491 ( N_RN_c_5887_n N_noxref_41_c_10185_n ) capacitor c=0.00657782f \
 //x=59.825 //y=2.22 //x2=46.675 //y2=0.995
cc_4492 ( N_RN_c_6712_p N_noxref_41_c_10185_n ) capacitor c=2.14837e-19 \
 //x=45.815 //y=0.755 //x2=46.675 //y2=0.995
cc_4493 ( N_RN_c_6154_n N_noxref_41_c_10185_n ) capacitor c=0.00123426f \
 //x=45.97 //y=0.91 //x2=46.675 //y2=0.995
cc_4494 ( N_RN_c_6155_n N_noxref_41_c_10185_n ) capacitor c=0.0129288f \
 //x=45.97 //y=1.22 //x2=46.675 //y2=0.995
cc_4495 ( N_RN_c_6156_n N_noxref_41_c_10185_n ) capacitor c=0.00142359f \
 //x=45.97 //y=1.45 //x2=46.675 //y2=0.995
cc_4496 ( N_RN_c_5887_n N_noxref_41_c_10190_n ) capacitor c=0.00147946f \
 //x=59.825 //y=2.22 //x2=47.645 //y2=0.54
cc_4497 ( N_RN_c_6149_n N_noxref_41_M28_noxref_d ) capacitor c=0.00223875f \
 //x=45.445 //y=0.91 //x2=45.52 //y2=0.91
cc_4498 ( N_RN_c_6152_n N_noxref_41_M28_noxref_d ) capacitor c=0.00262485f \
 //x=45.445 //y=1.22 //x2=45.52 //y2=0.91
cc_4499 ( N_RN_c_6712_p N_noxref_41_M28_noxref_d ) capacitor c=0.00220746f \
 //x=45.815 //y=0.755 //x2=45.52 //y2=0.91
cc_4500 ( N_RN_c_6720_p N_noxref_41_M28_noxref_d ) capacitor c=0.00194798f \
 //x=45.815 //y=1.375 //x2=45.52 //y2=0.91
cc_4501 ( N_RN_c_6154_n N_noxref_41_M28_noxref_d ) capacitor c=0.00198465f \
 //x=45.97 //y=0.91 //x2=45.52 //y2=0.91
cc_4502 ( N_RN_c_6155_n N_noxref_41_M28_noxref_d ) capacitor c=0.00128384f \
 //x=45.97 //y=1.22 //x2=45.52 //y2=0.91
cc_4503 ( N_RN_c_5887_n N_noxref_41_M29_noxref_s ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=46.625 //y2=0.375
cc_4504 ( N_RN_c_6154_n N_noxref_41_M29_noxref_s ) capacitor c=7.21316e-19 \
 //x=45.97 //y=0.91 //x2=46.625 //y2=0.375
cc_4505 ( N_RN_c_6155_n N_noxref_41_M29_noxref_s ) capacitor c=0.00348171f \
 //x=45.97 //y=1.22 //x2=46.625 //y2=0.375
cc_4506 ( N_RN_c_5887_n N_noxref_42_c_10255_n ) capacitor c=0.00635755f \
 //x=59.825 //y=2.22 //x2=49.165 //y2=1.495
cc_4507 ( N_RN_c_5887_n N_noxref_42_c_10237_n ) capacitor c=0.0223494f \
 //x=59.825 //y=2.22 //x2=50.05 //y2=1.58
cc_4508 ( N_RN_c_5887_n N_noxref_42_c_10244_n ) capacitor c=0.00649228f \
 //x=59.825 //y=2.22 //x2=50.135 //y2=1.495
cc_4509 ( N_RN_c_5887_n N_noxref_42_c_10245_n ) capacitor c=0.00178534f \
 //x=59.825 //y=2.22 //x2=51.02 //y2=0.53
cc_4510 ( N_RN_c_5887_n N_noxref_42_M30_noxref_s ) capacitor c=0.00113237f \
 //x=59.825 //y=2.22 //x2=49.03 //y2=0.365
cc_4511 ( N_RN_c_5887_n N_noxref_43_c_10312_n ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=52.39 //y2=1.505
cc_4512 ( N_RN_c_5887_n N_noxref_43_c_10288_n ) capacitor c=0.0225733f \
 //x=59.825 //y=2.22 //x2=53.275 //y2=1.59
cc_4513 ( N_RN_c_5887_n N_noxref_43_c_10305_n ) capacitor c=0.0203655f \
 //x=59.825 //y=2.22 //x2=54.245 //y2=1.59
cc_4514 ( N_RN_c_5887_n N_noxref_43_M32_noxref_s ) capacitor c=0.012425f \
 //x=59.825 //y=2.22 //x2=52.255 //y2=0.375
cc_4515 ( N_RN_c_5887_n N_noxref_44_c_10337_n ) capacitor c=0.00657782f \
 //x=59.825 //y=2.22 //x2=54.815 //y2=0.995
cc_4516 ( N_RN_c_5887_n N_noxref_44_c_10342_n ) capacitor c=0.00147946f \
 //x=59.825 //y=2.22 //x2=55.785 //y2=0.54
cc_4517 ( N_RN_c_5887_n N_noxref_44_M34_noxref_s ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=54.765 //y2=0.375
cc_4518 ( N_RN_c_5887_n N_noxref_45_c_10412_n ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=57.2 //y2=1.505
cc_4519 ( N_RN_c_5887_n N_noxref_45_c_10389_n ) capacitor c=0.0225733f \
 //x=59.825 //y=2.22 //x2=58.085 //y2=1.59
cc_4520 ( N_RN_c_5887_n N_noxref_45_c_10406_n ) capacitor c=0.0203655f \
 //x=59.825 //y=2.22 //x2=59.055 //y2=1.59
cc_4521 ( N_RN_c_5887_n N_noxref_45_M35_noxref_s ) capacitor c=0.012425f \
 //x=59.825 //y=2.22 //x2=57.065 //y2=0.375
cc_4522 ( N_RN_c_5887_n N_noxref_46_c_10438_n ) capacitor c=0.00657782f \
 //x=59.825 //y=2.22 //x2=59.625 //y2=0.995
cc_4523 ( N_RN_c_5899_n N_noxref_46_c_10443_n ) capacitor c=7.41833e-19 \
 //x=67.965 //y=2.22 //x2=60.595 //y2=0.54
cc_4524 ( N_RN_c_5907_n N_noxref_46_c_10443_n ) capacitor c=7.4531e-19 \
 //x=60.055 //y=2.22 //x2=60.595 //y2=0.54
cc_4525 ( N_RN_c_5919_n N_noxref_46_c_10443_n ) capacitor c=0.00204178f \
 //x=59.94 //y=2.08 //x2=60.595 //y2=0.54
cc_4526 ( N_RN_c_6268_n N_noxref_46_c_10443_n ) capacitor c=0.0194423f \
 //x=59.93 //y=0.915 //x2=60.595 //y2=0.54
cc_4527 ( N_RN_c_6515_p N_noxref_46_c_10443_n ) capacitor c=0.00656458f \
 //x=60.46 //y=0.915 //x2=60.595 //y2=0.54
cc_4528 ( N_RN_c_6283_n N_noxref_46_c_10443_n ) capacitor c=2.20712e-19 \
 //x=59.94 //y=2.08 //x2=60.595 //y2=0.54
cc_4529 ( N_RN_c_6269_n N_noxref_46_c_10470_n ) capacitor c=0.00538829f \
 //x=59.93 //y=1.26 //x2=59.71 //y2=0.995
cc_4530 ( N_RN_c_5887_n N_noxref_46_M37_noxref_s ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=59.575 //y2=0.375
cc_4531 ( N_RN_c_6268_n N_noxref_46_M37_noxref_s ) capacitor c=0.00538829f \
 //x=59.93 //y=0.915 //x2=59.575 //y2=0.375
cc_4532 ( N_RN_c_6270_n N_noxref_46_M37_noxref_s ) capacitor c=0.00538829f \
 //x=59.93 //y=1.57 //x2=59.575 //y2=0.375
cc_4533 ( N_RN_c_6515_p N_noxref_46_M37_noxref_s ) capacitor c=0.0143002f \
 //x=60.46 //y=0.915 //x2=59.575 //y2=0.375
cc_4534 ( N_RN_c_6475_p N_noxref_46_M37_noxref_s ) capacitor c=0.00290153f \
 //x=60.46 //y=1.26 //x2=59.575 //y2=0.375
cc_4535 ( N_RN_c_5899_n N_noxref_47_c_10509_n ) capacitor c=0.00635755f \
 //x=67.965 //y=2.22 //x2=62.115 //y2=1.495
cc_4536 ( N_RN_c_5899_n N_noxref_47_c_10491_n ) capacitor c=0.0223494f \
 //x=67.965 //y=2.22 //x2=63 //y2=1.58
cc_4537 ( N_RN_c_5899_n N_noxref_47_c_10498_n ) capacitor c=0.00649228f \
 //x=67.965 //y=2.22 //x2=63.085 //y2=1.495
cc_4538 ( N_RN_c_5899_n N_noxref_47_c_10499_n ) capacitor c=0.00178534f \
 //x=67.965 //y=2.22 //x2=63.97 //y2=0.53
cc_4539 ( N_RN_c_5899_n N_noxref_47_M38_noxref_s ) capacitor c=0.00113237f \
 //x=67.965 //y=2.22 //x2=61.98 //y2=0.365
cc_4540 ( N_RN_c_5899_n N_noxref_48_c_10565_n ) capacitor c=0.00642985f \
 //x=67.965 //y=2.22 //x2=65.34 //y2=1.505
cc_4541 ( N_RN_c_5899_n N_noxref_48_c_10542_n ) capacitor c=0.0225733f \
 //x=67.965 //y=2.22 //x2=66.225 //y2=1.59
cc_4542 ( N_RN_c_5899_n N_noxref_48_c_10559_n ) capacitor c=0.0203655f \
 //x=67.965 //y=2.22 //x2=67.195 //y2=1.59
cc_4543 ( N_RN_c_5899_n N_noxref_48_M40_noxref_s ) capacitor c=0.012425f \
 //x=67.965 //y=2.22 //x2=65.205 //y2=0.375
cc_4544 ( N_RN_c_5899_n N_noxref_49_c_10591_n ) capacitor c=0.00657782f \
 //x=67.965 //y=2.22 //x2=67.765 //y2=0.995
cc_4545 ( N_RN_c_5908_n N_noxref_49_c_10596_n ) capacitor c=7.41833e-19 \
 //x=71.665 //y=2.22 //x2=68.735 //y2=0.54
cc_4546 ( N_RN_c_5912_n N_noxref_49_c_10596_n ) capacitor c=7.4531e-19 \
 //x=68.195 //y=2.22 //x2=68.735 //y2=0.54
cc_4547 ( N_RN_c_5920_n N_noxref_49_c_10596_n ) capacitor c=0.00204178f \
 //x=68.08 //y=2.08 //x2=68.735 //y2=0.54
cc_4548 ( N_RN_c_6341_n N_noxref_49_c_10596_n ) capacitor c=0.0194423f \
 //x=68.07 //y=0.915 //x2=68.735 //y2=0.54
cc_4549 ( N_RN_c_6438_p N_noxref_49_c_10596_n ) capacitor c=0.00656458f \
 //x=68.6 //y=0.915 //x2=68.735 //y2=0.54
cc_4550 ( N_RN_c_6363_n N_noxref_49_c_10596_n ) capacitor c=2.20712e-19 \
 //x=68.08 //y=2.08 //x2=68.735 //y2=0.54
cc_4551 ( N_RN_c_6342_n N_noxref_49_c_10623_n ) capacitor c=0.00538829f \
 //x=68.07 //y=1.26 //x2=67.85 //y2=0.995
cc_4552 ( N_RN_c_5899_n N_noxref_49_M42_noxref_s ) capacitor c=0.00642985f \
 //x=67.965 //y=2.22 //x2=67.715 //y2=0.375
cc_4553 ( N_RN_c_6341_n N_noxref_49_M42_noxref_s ) capacitor c=0.00538829f \
 //x=68.07 //y=0.915 //x2=67.715 //y2=0.375
cc_4554 ( N_RN_c_6343_n N_noxref_49_M42_noxref_s ) capacitor c=0.00538829f \
 //x=68.07 //y=1.57 //x2=67.715 //y2=0.375
cc_4555 ( N_RN_c_6438_p N_noxref_49_M42_noxref_s ) capacitor c=0.0143002f \
 //x=68.6 //y=0.915 //x2=67.715 //y2=0.375
cc_4556 ( N_RN_c_6413_p N_noxref_49_M42_noxref_s ) capacitor c=0.00290153f \
 //x=68.6 //y=1.26 //x2=67.715 //y2=0.375
cc_4557 ( N_RN_c_5908_n N_noxref_50_c_10659_n ) capacitor c=0.00642985f \
 //x=71.665 //y=2.22 //x2=70.15 //y2=1.505
cc_4558 ( N_RN_c_5908_n N_noxref_50_c_10644_n ) capacitor c=0.0225733f \
 //x=71.665 //y=2.22 //x2=71.035 //y2=1.59
cc_4559 ( N_RN_c_6387_n N_noxref_50_c_10651_n ) capacitor c=0.0167228f \
 //x=71.345 //y=0.91 //x2=72.005 //y2=0.54
cc_4560 ( N_RN_c_6392_n N_noxref_50_c_10651_n ) capacitor c=0.00534519f \
 //x=71.87 //y=0.91 //x2=72.005 //y2=0.54
cc_4561 ( N_RN_c_5908_n N_noxref_50_c_10673_n ) capacitor c=0.0178105f \
 //x=71.665 //y=2.22 //x2=72.005 //y2=1.59
cc_4562 ( N_RN_c_5921_n N_noxref_50_c_10673_n ) capacitor c=0.0119919f \
 //x=71.78 //y=2.08 //x2=72.005 //y2=1.59
cc_4563 ( N_RN_c_6390_n N_noxref_50_c_10673_n ) capacitor c=0.0157358f \
 //x=71.345 //y=1.22 //x2=72.005 //y2=1.59
cc_4564 ( N_RN_c_6395_n N_noxref_50_c_10673_n ) capacitor c=0.0215856f \
 //x=71.87 //y=1.915 //x2=72.005 //y2=1.59
cc_4565 ( N_RN_c_5908_n N_noxref_50_M43_noxref_s ) capacitor c=0.00642985f \
 //x=71.665 //y=2.22 //x2=70.015 //y2=0.375
cc_4566 ( N_RN_c_6387_n N_noxref_50_M43_noxref_s ) capacitor c=0.00798959f \
 //x=71.345 //y=0.91 //x2=70.015 //y2=0.375
cc_4567 ( N_RN_c_6394_n N_noxref_50_M43_noxref_s ) capacitor c=0.00212176f \
 //x=71.87 //y=1.45 //x2=70.015 //y2=0.375
cc_4568 ( N_RN_c_6395_n N_noxref_50_M43_noxref_s ) capacitor c=0.00298115f \
 //x=71.87 //y=1.915 //x2=70.015 //y2=0.375
cc_4569 ( N_RN_c_6789_p N_noxref_51_c_10695_n ) capacitor c=2.14837e-19 \
 //x=71.715 //y=0.755 //x2=72.575 //y2=0.995
cc_4570 ( N_RN_c_6392_n N_noxref_51_c_10695_n ) capacitor c=0.00123426f \
 //x=71.87 //y=0.91 //x2=72.575 //y2=0.995
cc_4571 ( N_RN_c_6393_n N_noxref_51_c_10695_n ) capacitor c=0.0129288f \
 //x=71.87 //y=1.22 //x2=72.575 //y2=0.995
cc_4572 ( N_RN_c_6394_n N_noxref_51_c_10695_n ) capacitor c=0.00142359f \
 //x=71.87 //y=1.45 //x2=72.575 //y2=0.995
cc_4573 ( N_RN_c_6387_n N_noxref_51_M44_noxref_d ) capacitor c=0.00223875f \
 //x=71.345 //y=0.91 //x2=71.42 //y2=0.91
cc_4574 ( N_RN_c_6390_n N_noxref_51_M44_noxref_d ) capacitor c=0.00262485f \
 //x=71.345 //y=1.22 //x2=71.42 //y2=0.91
cc_4575 ( N_RN_c_6789_p N_noxref_51_M44_noxref_d ) capacitor c=0.00220746f \
 //x=71.715 //y=0.755 //x2=71.42 //y2=0.91
cc_4576 ( N_RN_c_6796_p N_noxref_51_M44_noxref_d ) capacitor c=0.00194798f \
 //x=71.715 //y=1.375 //x2=71.42 //y2=0.91
cc_4577 ( N_RN_c_6392_n N_noxref_51_M44_noxref_d ) capacitor c=0.00198465f \
 //x=71.87 //y=0.91 //x2=71.42 //y2=0.91
cc_4578 ( N_RN_c_6393_n N_noxref_51_M44_noxref_d ) capacitor c=0.00128384f \
 //x=71.87 //y=1.22 //x2=71.42 //y2=0.91
cc_4579 ( N_RN_c_6392_n N_noxref_51_M45_noxref_s ) capacitor c=7.21316e-19 \
 //x=71.87 //y=0.91 //x2=72.525 //y2=0.375
cc_4580 ( N_RN_c_6393_n N_noxref_51_M45_noxref_s ) capacitor c=0.00348171f \
 //x=71.87 //y=1.22 //x2=72.525 //y2=0.375
cc_4581 ( N_noxref_16_c_6831_n N_noxref_17_c_7362_n ) capacitor c=0.0838118f \
 //x=63.155 //y=4.07 //x2=55.015 //y2=3.33
cc_4582 ( N_noxref_16_c_6833_n N_noxref_17_c_7362_n ) capacitor c=0.0134837f \
 //x=53.025 //y=4.07 //x2=55.015 //y2=3.33
cc_4583 ( N_noxref_16_c_6801_n N_noxref_17_c_7362_n ) capacitor c=0.0224361f \
 //x=52.91 //y=2.08 //x2=55.015 //y2=3.33
cc_4584 ( N_noxref_16_c_6801_n N_noxref_17_c_7529_n ) capacitor c=4.54066e-19 \
 //x=52.91 //y=2.08 //x2=51.175 //y2=3.33
cc_4585 ( N_noxref_16_c_6831_n N_noxref_17_c_7559_n ) capacitor c=0.0558554f \
 //x=63.155 //y=4.07 //x2=60.565 //y2=3.33
cc_4586 ( N_noxref_16_c_6831_n N_noxref_17_c_7561_n ) capacitor c=0.0122198f \
 //x=63.155 //y=4.07 //x2=55.245 //y2=3.33
cc_4587 ( N_noxref_16_c_6831_n N_noxref_17_c_7648_n ) capacitor c=0.0100907f \
 //x=63.155 //y=4.07 //x2=62.415 //y2=3.33
cc_4588 ( N_noxref_16_c_6831_n N_noxref_17_c_7649_n ) capacitor c=4.80262e-19 \
 //x=63.155 //y=4.07 //x2=60.795 //y2=3.33
cc_4589 ( N_noxref_16_c_6831_n N_noxref_17_c_7650_n ) capacitor c=0.00539136f \
 //x=63.155 //y=4.07 //x2=63.895 //y2=3.33
cc_4590 ( N_noxref_16_c_6834_n N_noxref_17_c_7650_n ) capacitor c=0.00509378f \
 //x=68.705 //y=4.07 //x2=63.895 //y2=3.33
cc_4591 ( N_noxref_16_c_6962_n N_noxref_17_c_7650_n ) capacitor c=5.18288e-19 \
 //x=63.385 //y=4.07 //x2=63.895 //y2=3.33
cc_4592 ( N_noxref_16_c_6802_n N_noxref_17_c_7650_n ) capacitor c=0.0169786f \
 //x=63.27 //y=2.08 //x2=63.895 //y2=3.33
cc_4593 ( N_noxref_16_c_6831_n N_noxref_17_c_7651_n ) capacitor c=5.70482e-19 \
 //x=63.155 //y=4.07 //x2=62.645 //y2=3.33
cc_4594 ( N_noxref_16_c_6802_n N_noxref_17_c_7651_n ) capacitor c=7.76154e-19 \
 //x=63.27 //y=2.08 //x2=62.645 //y2=3.33
cc_4595 ( N_noxref_16_c_6834_n N_noxref_17_c_7652_n ) capacitor c=0.00994749f \
 //x=68.705 //y=4.07 //x2=65.745 //y2=3.33
cc_4596 ( N_noxref_16_c_6834_n N_noxref_17_c_7653_n ) capacitor c=5.70661e-19 \
 //x=68.705 //y=4.07 //x2=64.125 //y2=3.33
cc_4597 ( N_noxref_16_c_6802_n N_noxref_17_c_7653_n ) capacitor c=7.76154e-19 \
 //x=63.27 //y=2.08 //x2=64.125 //y2=3.33
cc_4598 ( N_noxref_16_c_6834_n N_noxref_17_c_7583_n ) capacitor c=0.0242164f \
 //x=68.705 //y=4.07 //x2=78.325 //y2=3.33
cc_4599 ( N_noxref_16_c_6836_n N_noxref_17_c_7583_n ) capacitor c=0.0977797f \
 //x=73.515 //y=4.07 //x2=78.325 //y2=3.33
cc_4600 ( N_noxref_16_c_6842_n N_noxref_17_c_7583_n ) capacitor c=4.80451e-19 \
 //x=68.935 //y=4.07 //x2=78.325 //y2=3.33
cc_4601 ( N_noxref_16_c_6845_n N_noxref_17_c_7583_n ) capacitor c=0.0100877f \
 //x=75.365 //y=4.07 //x2=78.325 //y2=3.33
cc_4602 ( N_noxref_16_c_6851_n N_noxref_17_c_7583_n ) capacitor c=4.80451e-19 \
 //x=73.745 //y=4.07 //x2=78.325 //y2=3.33
cc_4603 ( N_noxref_16_c_6854_n N_noxref_17_c_7583_n ) capacitor c=0.00613746f \
 //x=76.105 //y=4.07 //x2=78.325 //y2=3.33
cc_4604 ( N_noxref_16_c_6855_n N_noxref_17_c_7583_n ) capacitor c=5.77052e-19 \
 //x=75.595 //y=4.07 //x2=78.325 //y2=3.33
cc_4605 ( N_noxref_16_c_6877_n N_noxref_17_c_7583_n ) capacitor c=0.0187428f \
 //x=68.82 //y=4.07 //x2=78.325 //y2=3.33
cc_4606 ( N_noxref_16_c_6892_n N_noxref_17_c_7583_n ) capacitor c=0.018769f \
 //x=73.63 //y=4.07 //x2=78.325 //y2=3.33
cc_4607 ( N_noxref_16_c_6806_n N_noxref_17_c_7583_n ) capacitor c=0.0187666f \
 //x=75.48 //y=2.08 //x2=78.325 //y2=3.33
cc_4608 ( N_noxref_16_c_6807_n N_noxref_17_c_7583_n ) capacitor c=0.0169803f \
 //x=76.22 //y=2.08 //x2=78.325 //y2=3.33
cc_4609 ( N_noxref_16_c_6834_n N_noxref_17_c_7584_n ) capacitor c=5.3905e-19 \
 //x=68.705 //y=4.07 //x2=65.975 //y2=3.33
cc_4610 ( N_noxref_16_c_6833_n N_noxref_17_c_7303_n ) capacitor c=0.00103915f \
 //x=53.025 //y=4.07 //x2=51.06 //y2=3.33
cc_4611 ( N_noxref_16_c_6801_n N_noxref_17_c_7303_n ) capacitor c=0.0129951f \
 //x=52.91 //y=2.08 //x2=51.06 //y2=3.33
cc_4612 ( N_noxref_16_c_6831_n N_noxref_17_c_7304_n ) capacitor c=0.0206302f \
 //x=63.155 //y=4.07 //x2=55.13 //y2=2.08
cc_4613 ( N_noxref_16_c_6801_n N_noxref_17_c_7304_n ) capacitor c=0.0011415f \
 //x=52.91 //y=2.08 //x2=55.13 //y2=2.08
cc_4614 ( N_noxref_16_c_6831_n N_noxref_17_c_7399_n ) capacitor c=0.0181982f \
 //x=63.155 //y=4.07 //x2=60.68 //y2=3.33
cc_4615 ( N_noxref_16_c_6802_n N_noxref_17_c_7399_n ) capacitor c=5.85299e-19 \
 //x=63.27 //y=2.08 //x2=60.68 //y2=3.33
cc_4616 ( N_noxref_16_c_6831_n N_noxref_17_c_7306_n ) capacitor c=0.0184765f \
 //x=63.155 //y=4.07 //x2=62.53 //y2=2.08
cc_4617 ( N_noxref_16_c_6962_n N_noxref_17_c_7306_n ) capacitor c=0.00179385f \
 //x=63.385 //y=4.07 //x2=62.53 //y2=2.08
cc_4618 ( N_noxref_16_c_6968_n N_noxref_17_c_7306_n ) capacitor c=0.00400249f \
 //x=63.27 //y=4.535 //x2=62.53 //y2=2.08
cc_4619 ( N_noxref_16_c_6802_n N_noxref_17_c_7306_n ) capacitor c=0.0735279f \
 //x=63.27 //y=2.08 //x2=62.53 //y2=2.08
cc_4620 ( N_noxref_16_c_7057_n N_noxref_17_c_7306_n ) capacitor c=0.00282278f \
 //x=63.27 //y=2.08 //x2=62.53 //y2=2.08
cc_4621 ( N_noxref_16_c_6998_n N_noxref_17_c_7306_n ) capacitor c=0.00344981f \
 //x=63.3 //y=4.7 //x2=62.53 //y2=2.08
cc_4622 ( N_noxref_16_c_6968_n N_noxref_17_c_7403_n ) capacitor c=0.0127164f \
 //x=63.27 //y=4.535 //x2=63.445 //y2=5.2
cc_4623 ( N_noxref_16_M132_noxref_g N_noxref_17_c_7403_n ) capacitor \
 c=0.0166421f //x=63.31 //y=6.02 //x2=63.445 //y2=5.2
cc_4624 ( N_noxref_16_c_6998_n N_noxref_17_c_7403_n ) capacitor c=0.00346527f \
 //x=63.3 //y=4.7 //x2=63.445 //y2=5.2
cc_4625 ( N_noxref_16_M133_noxref_g N_noxref_17_c_7409_n ) capacitor \
 c=0.018922f //x=63.75 //y=6.02 //x2=63.925 //y2=5.2
cc_4626 ( N_noxref_16_c_7056_n N_noxref_17_c_7307_n ) capacitor c=0.00371277f \
 //x=63.68 //y=1.405 //x2=63.925 //y2=1.655
cc_4627 ( N_noxref_16_c_7116_p N_noxref_17_c_7307_n ) capacitor c=0.00457401f \
 //x=63.835 //y=1.25 //x2=63.925 //y2=1.655
cc_4628 ( N_noxref_16_c_6834_n N_noxref_17_c_7308_n ) capacitor c=0.0181936f \
 //x=68.705 //y=4.07 //x2=64.01 //y2=3.33
cc_4629 ( N_noxref_16_c_6962_n N_noxref_17_c_7308_n ) capacitor c=0.00179385f \
 //x=63.385 //y=4.07 //x2=64.01 //y2=3.33
cc_4630 ( N_noxref_16_c_6968_n N_noxref_17_c_7308_n ) capacitor c=0.0101115f \
 //x=63.27 //y=4.535 //x2=64.01 //y2=3.33
cc_4631 ( N_noxref_16_c_6802_n N_noxref_17_c_7308_n ) capacitor c=0.0685501f \
 //x=63.27 //y=2.08 //x2=64.01 //y2=3.33
cc_4632 ( N_noxref_16_c_6867_n N_noxref_17_c_7308_n ) capacitor c=2.97874e-19 \
 //x=66.365 //y=5.155 //x2=64.01 //y2=3.33
cc_4633 ( N_noxref_16_c_6997_n N_noxref_17_c_7308_n ) capacitor c=0.0142673f \
 //x=63.675 //y=4.79 //x2=64.01 //y2=3.33
cc_4634 ( N_noxref_16_c_7057_n N_noxref_17_c_7308_n ) capacitor c=0.00731987f \
 //x=63.27 //y=2.08 //x2=64.01 //y2=3.33
cc_4635 ( N_noxref_16_c_7124_p N_noxref_17_c_7308_n ) capacitor c=0.00306024f \
 //x=63.27 //y=1.915 //x2=64.01 //y2=3.33
cc_4636 ( N_noxref_16_c_6998_n N_noxref_17_c_7308_n ) capacitor c=0.00517969f \
 //x=63.3 //y=4.7 //x2=64.01 //y2=3.33
cc_4637 ( N_noxref_16_c_6834_n N_noxref_17_c_7309_n ) capacitor c=0.019517f \
 //x=68.705 //y=4.07 //x2=65.86 //y2=2.08
cc_4638 ( N_noxref_16_c_6802_n N_noxref_17_c_7309_n ) capacitor c=5.85299e-19 \
 //x=63.27 //y=2.08 //x2=65.86 //y2=2.08
cc_4639 ( N_noxref_16_c_6807_n N_noxref_17_c_7310_n ) capacitor c=8.49976e-19 \
 //x=76.22 //y=2.08 //x2=78.44 //y2=2.08
cc_4640 ( N_noxref_16_c_6997_n N_noxref_17_c_7824_n ) capacitor c=0.00407665f \
 //x=63.675 //y=4.79 //x2=63.53 //y2=5.2
cc_4641 ( N_noxref_16_M132_noxref_g N_noxref_17_M130_noxref_g ) capacitor \
 c=0.0104611f //x=63.31 //y=6.02 //x2=62.43 //y2=6.02
cc_4642 ( N_noxref_16_M132_noxref_g N_noxref_17_M131_noxref_g ) capacitor \
 c=0.106811f //x=63.31 //y=6.02 //x2=62.87 //y2=6.02
cc_4643 ( N_noxref_16_M133_noxref_g N_noxref_17_M131_noxref_g ) capacitor \
 c=0.0100341f //x=63.75 //y=6.02 //x2=62.87 //y2=6.02
cc_4644 ( N_noxref_16_c_6867_n N_noxref_17_M134_noxref_g ) capacitor \
 c=0.0213876f //x=66.365 //y=5.155 //x2=66.06 //y2=6.02
cc_4645 ( N_noxref_16_c_6863_n N_noxref_17_M135_noxref_g ) capacitor \
 c=0.0168349f //x=67.075 //y=5.155 //x2=66.5 //y2=6.02
cc_4646 ( N_noxref_16_M134_noxref_d N_noxref_17_M135_noxref_g ) capacitor \
 c=0.0180032f //x=66.135 //y=5.02 //x2=66.5 //y2=6.02
cc_4647 ( N_noxref_16_c_7136_p N_noxref_17_c_7315_n ) capacitor c=4.86506e-19 \
 //x=63.305 //y=0.905 //x2=62.335 //y2=0.865
cc_4648 ( N_noxref_16_c_7136_p N_noxref_17_c_7317_n ) capacitor c=0.00152104f \
 //x=63.305 //y=0.905 //x2=62.335 //y2=1.21
cc_4649 ( N_noxref_16_c_7138_p N_noxref_17_c_7318_n ) capacitor c=0.00109982f \
 //x=63.305 //y=1.25 //x2=62.335 //y2=1.52
cc_4650 ( N_noxref_16_c_7139_p N_noxref_17_c_7318_n ) capacitor c=9.57794e-19 \
 //x=63.305 //y=1.56 //x2=62.335 //y2=1.52
cc_4651 ( N_noxref_16_c_6802_n N_noxref_17_c_7319_n ) capacitor c=0.00284029f \
 //x=63.27 //y=2.08 //x2=62.335 //y2=1.915
cc_4652 ( N_noxref_16_c_7139_p N_noxref_17_c_7319_n ) capacitor c=0.00662747f \
 //x=63.305 //y=1.56 //x2=62.335 //y2=1.915
cc_4653 ( N_noxref_16_c_7057_n N_noxref_17_c_7319_n ) capacitor c=0.0172771f \
 //x=63.27 //y=2.08 //x2=62.335 //y2=1.915
cc_4654 ( N_noxref_16_c_7136_p N_noxref_17_c_7322_n ) capacitor c=0.0151475f \
 //x=63.305 //y=0.905 //x2=62.865 //y2=0.865
cc_4655 ( N_noxref_16_c_7144_p N_noxref_17_c_7322_n ) capacitor c=0.00124821f \
 //x=63.835 //y=0.905 //x2=62.865 //y2=0.865
cc_4656 ( N_noxref_16_c_7138_p N_noxref_17_c_7324_n ) capacitor c=0.0111064f \
 //x=63.305 //y=1.25 //x2=62.865 //y2=1.21
cc_4657 ( N_noxref_16_c_7139_p N_noxref_17_c_7324_n ) capacitor c=0.00862358f \
 //x=63.305 //y=1.56 //x2=62.865 //y2=1.21
cc_4658 ( N_noxref_16_c_7116_p N_noxref_17_c_7324_n ) capacitor c=0.00200715f \
 //x=63.835 //y=1.25 //x2=62.865 //y2=1.21
cc_4659 ( N_noxref_16_c_6867_n N_noxref_17_c_7627_n ) capacitor c=0.00428486f \
 //x=66.365 //y=5.155 //x2=66.425 //y2=4.79
cc_4660 ( N_noxref_16_c_6968_n N_noxref_17_c_7451_n ) capacitor c=0.00417994f \
 //x=63.27 //y=4.535 //x2=62.53 //y2=4.7
cc_4661 ( N_noxref_16_c_6998_n N_noxref_17_c_7451_n ) capacitor c=0.0293367f \
 //x=63.3 //y=4.7 //x2=62.53 //y2=4.7
cc_4662 ( N_noxref_16_c_7136_p N_noxref_17_M39_noxref_d ) capacitor \
 c=0.00217566f //x=63.305 //y=0.905 //x2=63.38 //y2=0.905
cc_4663 ( N_noxref_16_c_7138_p N_noxref_17_M39_noxref_d ) capacitor \
 c=0.0034598f //x=63.305 //y=1.25 //x2=63.38 //y2=0.905
cc_4664 ( N_noxref_16_c_7139_p N_noxref_17_M39_noxref_d ) capacitor \
 c=0.00669531f //x=63.305 //y=1.56 //x2=63.38 //y2=0.905
cc_4665 ( N_noxref_16_c_7154_p N_noxref_17_M39_noxref_d ) capacitor \
 c=0.00241102f //x=63.68 //y=0.75 //x2=63.38 //y2=0.905
cc_4666 ( N_noxref_16_c_7056_n N_noxref_17_M39_noxref_d ) capacitor \
 c=0.0137169f //x=63.68 //y=1.405 //x2=63.38 //y2=0.905
cc_4667 ( N_noxref_16_c_7144_p N_noxref_17_M39_noxref_d ) capacitor \
 c=0.00132245f //x=63.835 //y=0.905 //x2=63.38 //y2=0.905
cc_4668 ( N_noxref_16_c_7116_p N_noxref_17_M39_noxref_d ) capacitor \
 c=0.00566463f //x=63.835 //y=1.25 //x2=63.38 //y2=0.905
cc_4669 ( N_noxref_16_c_7124_p N_noxref_17_M39_noxref_d ) capacitor \
 c=0.00660593f //x=63.27 //y=1.915 //x2=63.38 //y2=0.905
cc_4670 ( N_noxref_16_M132_noxref_g N_noxref_17_M132_noxref_d ) capacitor \
 c=0.0173476f //x=63.31 //y=6.02 //x2=63.385 //y2=5.02
cc_4671 ( N_noxref_16_M133_noxref_g N_noxref_17_M132_noxref_d ) capacitor \
 c=0.0179769f //x=63.75 //y=6.02 //x2=63.385 //y2=5.02
cc_4672 ( N_noxref_16_c_6836_n N_noxref_18_c_8076_n ) capacitor c=0.0445797f \
 //x=73.515 //y=4.07 //x2=76.845 //y2=3.7
cc_4673 ( N_noxref_16_c_6845_n N_noxref_18_c_8076_n ) capacitor c=0.14702f \
 //x=75.365 //y=4.07 //x2=76.845 //y2=3.7
cc_4674 ( N_noxref_16_c_6851_n N_noxref_18_c_8076_n ) capacitor c=0.0268461f \
 //x=73.745 //y=4.07 //x2=76.845 //y2=3.7
cc_4675 ( N_noxref_16_c_6854_n N_noxref_18_c_8076_n ) capacitor c=0.0739186f \
 //x=76.105 //y=4.07 //x2=76.845 //y2=3.7
cc_4676 ( N_noxref_16_c_6855_n N_noxref_18_c_8076_n ) capacitor c=0.0265532f \
 //x=75.595 //y=4.07 //x2=76.845 //y2=3.7
cc_4677 ( N_noxref_16_c_6892_n N_noxref_18_c_8076_n ) capacitor c=0.0206044f \
 //x=73.63 //y=4.07 //x2=76.845 //y2=3.7
cc_4678 ( N_noxref_16_c_6806_n N_noxref_18_c_8076_n ) capacitor c=0.020561f \
 //x=75.48 //y=2.08 //x2=76.845 //y2=3.7
cc_4679 ( N_noxref_16_c_6807_n N_noxref_18_c_8076_n ) capacitor c=0.0187982f \
 //x=76.22 //y=2.08 //x2=76.845 //y2=3.7
cc_4680 ( N_noxref_16_c_7169_p N_noxref_18_c_8076_n ) capacitor c=0.00624857f \
 //x=76.625 //y=4.79 //x2=76.845 //y2=3.7
cc_4681 ( N_noxref_16_c_7170_p N_noxref_18_c_8076_n ) capacitor c=2.85902e-19 \
 //x=76.25 //y=4.7 //x2=76.845 //y2=3.7
cc_4682 ( N_noxref_16_c_6836_n N_noxref_18_c_8127_n ) capacitor c=0.0292842f \
 //x=73.515 //y=4.07 //x2=73.005 //y2=3.7
cc_4683 ( N_noxref_16_c_6892_n N_noxref_18_c_8127_n ) capacitor c=0.00117715f \
 //x=73.63 //y=4.07 //x2=73.005 //y2=3.7
cc_4684 ( N_noxref_16_c_6807_n N_noxref_18_c_8079_n ) capacitor c=0.00117715f \
 //x=76.22 //y=2.08 //x2=77.075 //y2=3.7
cc_4685 ( N_noxref_16_c_6854_n N_noxref_18_c_8085_n ) capacitor c=0.00480721f \
 //x=76.105 //y=4.07 //x2=79.665 //y2=4.07
cc_4686 ( N_noxref_16_c_6836_n N_noxref_18_c_8065_n ) capacitor c=0.0237491f \
 //x=73.515 //y=4.07 //x2=72.89 //y2=2.08
cc_4687 ( N_noxref_16_c_6851_n N_noxref_18_c_8065_n ) capacitor c=0.00131333f \
 //x=73.745 //y=4.07 //x2=72.89 //y2=2.08
cc_4688 ( N_noxref_16_c_6892_n N_noxref_18_c_8065_n ) capacitor c=0.0824281f \
 //x=73.63 //y=4.07 //x2=72.89 //y2=2.08
cc_4689 ( N_noxref_16_c_6806_n N_noxref_18_c_8065_n ) capacitor c=5.57926e-19 \
 //x=75.48 //y=2.08 //x2=72.89 //y2=2.08
cc_4690 ( N_noxref_16_c_7179_p N_noxref_18_c_8065_n ) capacitor c=0.0168082f \
 //x=72.85 //y=5.155 //x2=72.89 //y2=2.08
cc_4691 ( N_noxref_16_c_6854_n N_noxref_18_c_8087_n ) capacitor c=0.00208151f \
 //x=76.105 //y=4.07 //x2=76.395 //y2=5.2
cc_4692 ( N_noxref_16_c_7181_p N_noxref_18_c_8087_n ) capacitor c=0.0129794f \
 //x=76.22 //y=4.535 //x2=76.395 //y2=5.2
cc_4693 ( N_noxref_16_M147_noxref_g N_noxref_18_c_8087_n ) capacitor \
 c=0.0179814f //x=75.82 //y=6.02 //x2=76.395 //y2=5.2
cc_4694 ( N_noxref_16_M148_noxref_g N_noxref_18_c_8087_n ) capacitor \
 c=0.0166421f //x=76.26 //y=6.02 //x2=76.395 //y2=5.2
cc_4695 ( N_noxref_16_c_7170_p N_noxref_18_c_8087_n ) capacitor c=0.00346627f \
 //x=76.25 //y=4.7 //x2=76.395 //y2=5.2
cc_4696 ( N_noxref_16_c_6854_n N_noxref_18_c_8091_n ) capacitor c=0.0124916f \
 //x=76.105 //y=4.07 //x2=75.685 //y2=5.2
cc_4697 ( N_noxref_16_c_6855_n N_noxref_18_c_8091_n ) capacitor c=7.54159e-19 \
 //x=75.595 //y=4.07 //x2=75.685 //y2=5.2
cc_4698 ( N_noxref_16_c_6806_n N_noxref_18_c_8091_n ) capacitor c=0.00529872f \
 //x=75.48 //y=2.08 //x2=75.685 //y2=5.2
cc_4699 ( N_noxref_16_M146_noxref_g N_noxref_18_c_8091_n ) capacitor \
 c=0.0177326f //x=75.38 //y=6.02 //x2=75.685 //y2=5.2
cc_4700 ( N_noxref_16_c_6918_n N_noxref_18_c_8091_n ) capacitor c=0.00582217f \
 //x=75.48 //y=4.7 //x2=75.685 //y2=5.2
cc_4701 ( N_noxref_16_M149_noxref_g N_noxref_18_c_8093_n ) capacitor \
 c=0.0206783f //x=76.7 //y=6.02 //x2=76.875 //y2=5.2
cc_4702 ( N_noxref_16_c_7191_p N_noxref_18_c_8066_n ) capacitor c=0.00359704f \
 //x=76.63 //y=1.405 //x2=76.875 //y2=1.655
cc_4703 ( N_noxref_16_c_7192_p N_noxref_18_c_8066_n ) capacitor c=0.00457401f \
 //x=76.785 //y=1.25 //x2=76.875 //y2=1.655
cc_4704 ( N_noxref_16_c_6854_n N_noxref_18_c_8067_n ) capacitor c=0.00465962f \
 //x=76.105 //y=4.07 //x2=76.96 //y2=3.7
cc_4705 ( N_noxref_16_c_6892_n N_noxref_18_c_8067_n ) capacitor c=3.52729e-19 \
 //x=73.63 //y=4.07 //x2=76.96 //y2=3.7
cc_4706 ( N_noxref_16_c_6806_n N_noxref_18_c_8067_n ) capacitor c=0.00377558f \
 //x=75.48 //y=2.08 //x2=76.96 //y2=3.7
cc_4707 ( N_noxref_16_c_7181_p N_noxref_18_c_8067_n ) capacitor c=0.0101197f \
 //x=76.22 //y=4.535 //x2=76.96 //y2=3.7
cc_4708 ( N_noxref_16_c_6807_n N_noxref_18_c_8067_n ) capacitor c=0.074114f \
 //x=76.22 //y=2.08 //x2=76.96 //y2=3.7
cc_4709 ( N_noxref_16_c_7169_p N_noxref_18_c_8067_n ) capacitor c=0.0142673f \
 //x=76.625 //y=4.79 //x2=76.96 //y2=3.7
cc_4710 ( N_noxref_16_c_7199_p N_noxref_18_c_8067_n ) capacitor c=0.00877984f \
 //x=76.22 //y=2.08 //x2=76.96 //y2=3.7
cc_4711 ( N_noxref_16_c_7200_p N_noxref_18_c_8067_n ) capacitor c=0.00306024f \
 //x=76.22 //y=1.915 //x2=76.96 //y2=3.7
cc_4712 ( N_noxref_16_c_7170_p N_noxref_18_c_8067_n ) capacitor c=0.00517969f \
 //x=76.25 //y=4.7 //x2=76.96 //y2=3.7
cc_4713 ( N_noxref_16_c_7169_p N_noxref_18_c_8188_n ) capacitor c=0.00421574f \
 //x=76.625 //y=4.79 //x2=76.48 //y2=5.2
cc_4714 ( N_noxref_16_c_6884_n N_noxref_18_M144_noxref_g ) capacitor \
 c=0.0184045f //x=72.765 //y=5.155 //x2=72.63 //y2=6.02
cc_4715 ( N_noxref_16_M144_noxref_d N_noxref_18_M144_noxref_g ) capacitor \
 c=0.0180032f //x=72.705 //y=5.02 //x2=72.63 //y2=6.02
cc_4716 ( N_noxref_16_c_6888_n N_noxref_18_M145_noxref_g ) capacitor \
 c=0.0205426f //x=73.545 //y=5.155 //x2=73.07 //y2=6.02
cc_4717 ( N_noxref_16_M144_noxref_d N_noxref_18_M145_noxref_g ) capacitor \
 c=0.0194246f //x=72.705 //y=5.02 //x2=73.07 //y2=6.02
cc_4718 ( N_noxref_16_M45_noxref_d N_noxref_18_c_8137_n ) capacitor \
 c=0.00217566f //x=72.955 //y=0.915 //x2=72.88 //y2=0.915
cc_4719 ( N_noxref_16_M45_noxref_d N_noxref_18_c_8138_n ) capacitor \
 c=0.0034598f //x=72.955 //y=0.915 //x2=72.88 //y2=1.26
cc_4720 ( N_noxref_16_M45_noxref_d N_noxref_18_c_8139_n ) capacitor \
 c=0.00544291f //x=72.955 //y=0.915 //x2=72.88 //y2=1.57
cc_4721 ( N_noxref_16_M45_noxref_d N_noxref_18_c_8196_n ) capacitor \
 c=0.00241102f //x=72.955 //y=0.915 //x2=73.255 //y2=0.76
cc_4722 ( N_noxref_16_c_6805_n N_noxref_18_c_8197_n ) capacitor c=0.00359704f \
 //x=73.545 //y=1.665 //x2=73.255 //y2=1.415
cc_4723 ( N_noxref_16_M45_noxref_d N_noxref_18_c_8197_n ) capacitor \
 c=0.0140297f //x=72.955 //y=0.915 //x2=73.255 //y2=1.415
cc_4724 ( N_noxref_16_M45_noxref_d N_noxref_18_c_8199_n ) capacitor \
 c=0.00219619f //x=72.955 //y=0.915 //x2=73.41 //y2=0.915
cc_4725 ( N_noxref_16_c_6805_n N_noxref_18_c_8200_n ) capacitor c=0.00457401f \
 //x=73.545 //y=1.665 //x2=73.41 //y2=1.26
cc_4726 ( N_noxref_16_M45_noxref_d N_noxref_18_c_8200_n ) capacitor \
 c=0.00603828f //x=72.955 //y=0.915 //x2=73.41 //y2=1.26
cc_4727 ( N_noxref_16_c_6892_n N_noxref_18_c_8140_n ) capacitor c=0.00772308f \
 //x=73.63 //y=4.07 //x2=72.89 //y2=2.08
cc_4728 ( N_noxref_16_c_6892_n N_noxref_18_c_8143_n ) capacitor c=0.00283672f \
 //x=73.63 //y=4.07 //x2=72.89 //y2=1.915
cc_4729 ( N_noxref_16_M45_noxref_d N_noxref_18_c_8143_n ) capacitor \
 c=0.00661782f //x=72.955 //y=0.915 //x2=72.89 //y2=1.915
cc_4730 ( N_noxref_16_c_6836_n N_noxref_18_c_8144_n ) capacitor c=0.00775263f \
 //x=73.515 //y=4.07 //x2=72.89 //y2=4.7
cc_4731 ( N_noxref_16_c_6888_n N_noxref_18_c_8144_n ) capacitor c=0.00201851f \
 //x=73.545 //y=5.155 //x2=72.89 //y2=4.7
cc_4732 ( N_noxref_16_c_6892_n N_noxref_18_c_8144_n ) capacitor c=0.013844f \
 //x=73.63 //y=4.07 //x2=72.89 //y2=4.7
cc_4733 ( N_noxref_16_c_7179_p N_noxref_18_c_8144_n ) capacitor c=0.00475729f \
 //x=72.85 //y=5.155 //x2=72.89 //y2=4.7
cc_4734 ( N_noxref_16_c_7223_p N_noxref_18_M47_noxref_d ) capacitor \
 c=0.00217566f //x=76.255 //y=0.905 //x2=76.33 //y2=0.905
cc_4735 ( N_noxref_16_c_7224_p N_noxref_18_M47_noxref_d ) capacitor \
 c=0.0034598f //x=76.255 //y=1.25 //x2=76.33 //y2=0.905
cc_4736 ( N_noxref_16_c_7225_p N_noxref_18_M47_noxref_d ) capacitor \
 c=0.0065582f //x=76.255 //y=1.56 //x2=76.33 //y2=0.905
cc_4737 ( N_noxref_16_c_7226_p N_noxref_18_M47_noxref_d ) capacitor \
 c=0.00241102f //x=76.63 //y=0.75 //x2=76.33 //y2=0.905
cc_4738 ( N_noxref_16_c_7191_p N_noxref_18_M47_noxref_d ) capacitor \
 c=0.0138845f //x=76.63 //y=1.405 //x2=76.33 //y2=0.905
cc_4739 ( N_noxref_16_c_7228_p N_noxref_18_M47_noxref_d ) capacitor \
 c=0.00132245f //x=76.785 //y=0.905 //x2=76.33 //y2=0.905
cc_4740 ( N_noxref_16_c_7192_p N_noxref_18_M47_noxref_d ) capacitor \
 c=0.00566463f //x=76.785 //y=1.25 //x2=76.33 //y2=0.905
cc_4741 ( N_noxref_16_c_7200_p N_noxref_18_M47_noxref_d ) capacitor \
 c=0.00660593f //x=76.22 //y=1.915 //x2=76.33 //y2=0.905
cc_4742 ( N_noxref_16_M147_noxref_g N_noxref_18_M146_noxref_d ) capacitor \
 c=0.0173476f //x=75.82 //y=6.02 //x2=75.455 //y2=5.02
cc_4743 ( N_noxref_16_M148_noxref_g N_noxref_18_M148_noxref_d ) capacitor \
 c=0.0173477f //x=76.26 //y=6.02 //x2=76.335 //y2=5.02
cc_4744 ( N_noxref_16_M149_noxref_g N_noxref_18_M148_noxref_d ) capacitor \
 c=0.0179769f //x=76.7 //y=6.02 //x2=76.335 //y2=5.02
cc_4745 ( N_noxref_16_c_6831_n N_noxref_20_c_8516_n ) capacitor c=0.0176477f \
 //x=63.155 //y=4.07 //x2=83.505 //y2=2.96
cc_4746 ( N_noxref_16_c_6833_n N_noxref_20_c_8516_n ) capacitor c=5.11078e-19 \
 //x=53.025 //y=4.07 //x2=83.505 //y2=2.96
cc_4747 ( N_noxref_16_c_6836_n N_noxref_20_c_8516_n ) capacitor c=0.0132553f \
 //x=73.515 //y=4.07 //x2=83.505 //y2=2.96
cc_4748 ( N_noxref_16_c_6801_n N_noxref_20_c_8516_n ) capacitor c=0.0197554f \
 //x=52.91 //y=2.08 //x2=83.505 //y2=2.96
cc_4749 ( N_noxref_16_c_6802_n N_noxref_20_c_8516_n ) capacitor c=0.0192451f \
 //x=63.27 //y=2.08 //x2=83.505 //y2=2.96
cc_4750 ( N_noxref_16_c_6877_n N_noxref_20_c_8516_n ) capacitor c=0.0210712f \
 //x=68.82 //y=4.07 //x2=83.505 //y2=2.96
cc_4751 ( N_noxref_16_c_7240_p N_noxref_20_c_8516_n ) capacitor c=0.00838703f \
 //x=73.23 //y=1.665 //x2=83.505 //y2=2.96
cc_4752 ( N_noxref_16_c_6892_n N_noxref_20_c_8516_n ) capacitor c=0.0238173f \
 //x=73.63 //y=4.07 //x2=83.505 //y2=2.96
cc_4753 ( N_noxref_16_c_6806_n N_noxref_20_c_8516_n ) capacitor c=0.0231982f \
 //x=75.48 //y=2.08 //x2=83.505 //y2=2.96
cc_4754 ( N_noxref_16_c_6807_n N_noxref_20_c_8516_n ) capacitor c=0.0214083f \
 //x=76.22 //y=2.08 //x2=83.505 //y2=2.96
cc_4755 ( N_noxref_16_c_6823_n N_noxref_20_c_8516_n ) capacitor c=0.00425556f \
 //x=75.285 //y=1.915 //x2=83.505 //y2=2.96
cc_4756 ( N_noxref_16_c_7199_p N_noxref_20_c_8516_n ) capacitor c=0.00172252f \
 //x=76.22 //y=2.08 //x2=83.505 //y2=2.96
cc_4757 ( N_noxref_16_c_6813_n N_noxref_43_c_10312_n ) capacitor c=0.0034165f \
 //x=52.61 //y=1.915 //x2=52.39 //y2=1.505
cc_4758 ( N_noxref_16_c_6801_n N_noxref_43_c_10288_n ) capacitor c=0.0115578f \
 //x=52.91 //y=2.08 //x2=53.275 //y2=1.59
cc_4759 ( N_noxref_16_c_6812_n N_noxref_43_c_10288_n ) capacitor c=0.00697148f \
 //x=52.61 //y=1.53 //x2=53.275 //y2=1.59
cc_4760 ( N_noxref_16_c_6813_n N_noxref_43_c_10288_n ) capacitor c=0.0204849f \
 //x=52.61 //y=1.915 //x2=53.275 //y2=1.59
cc_4761 ( N_noxref_16_c_6815_n N_noxref_43_c_10288_n ) capacitor c=0.00610316f \
 //x=52.985 //y=1.375 //x2=53.275 //y2=1.59
cc_4762 ( N_noxref_16_c_6818_n N_noxref_43_c_10288_n ) capacitor c=0.00698822f \
 //x=53.14 //y=1.22 //x2=53.275 //y2=1.59
cc_4763 ( N_noxref_16_c_6809_n N_noxref_43_M32_noxref_s ) capacitor \
 c=0.0327271f //x=52.61 //y=0.875 //x2=52.255 //y2=0.375
cc_4764 ( N_noxref_16_c_6812_n N_noxref_43_M32_noxref_s ) capacitor \
 c=7.99997e-19 //x=52.61 //y=1.53 //x2=52.255 //y2=0.375
cc_4765 ( N_noxref_16_c_6813_n N_noxref_43_M32_noxref_s ) capacitor \
 c=0.00122123f //x=52.61 //y=1.915 //x2=52.255 //y2=0.375
cc_4766 ( N_noxref_16_c_6816_n N_noxref_43_M32_noxref_s ) capacitor \
 c=0.0121427f //x=53.14 //y=0.875 //x2=52.255 //y2=0.375
cc_4767 ( N_noxref_16_c_7139_p N_noxref_47_c_10498_n ) capacitor c=0.00623646f \
 //x=63.305 //y=1.56 //x2=63.085 //y2=1.495
cc_4768 ( N_noxref_16_c_7057_n N_noxref_47_c_10498_n ) capacitor c=0.00173579f \
 //x=63.27 //y=2.08 //x2=63.085 //y2=1.495
cc_4769 ( N_noxref_16_c_6802_n N_noxref_47_c_10499_n ) capacitor c=0.00156605f \
 //x=63.27 //y=2.08 //x2=63.97 //y2=0.53
cc_4770 ( N_noxref_16_c_7136_p N_noxref_47_c_10499_n ) capacitor c=0.0188655f \
 //x=63.305 //y=0.905 //x2=63.97 //y2=0.53
cc_4771 ( N_noxref_16_c_7144_p N_noxref_47_c_10499_n ) capacitor c=0.00656458f \
 //x=63.835 //y=0.905 //x2=63.97 //y2=0.53
cc_4772 ( N_noxref_16_c_7057_n N_noxref_47_c_10499_n ) capacitor c=2.1838e-19 \
 //x=63.27 //y=2.08 //x2=63.97 //y2=0.53
cc_4773 ( N_noxref_16_c_7136_p N_noxref_47_M38_noxref_s ) capacitor \
 c=0.00623646f //x=63.305 //y=0.905 //x2=61.98 //y2=0.365
cc_4774 ( N_noxref_16_c_7144_p N_noxref_47_M38_noxref_s ) capacitor \
 c=0.0143002f //x=63.835 //y=0.905 //x2=61.98 //y2=0.365
cc_4775 ( N_noxref_16_c_7116_p N_noxref_47_M38_noxref_s ) capacitor \
 c=0.00290153f //x=63.835 //y=1.25 //x2=61.98 //y2=0.365
cc_4776 ( N_noxref_16_M42_noxref_d N_noxref_48_M40_noxref_s ) capacitor \
 c=0.00309936f //x=68.145 //y=0.915 //x2=65.205 //y2=0.375
cc_4777 ( N_noxref_16_c_6804_n N_noxref_49_c_10596_n ) capacitor c=0.00457167f \
 //x=68.735 //y=1.665 //x2=68.735 //y2=0.54
cc_4778 ( N_noxref_16_M42_noxref_d N_noxref_49_c_10596_n ) capacitor \
 c=0.0115903f //x=68.145 //y=0.915 //x2=68.735 //y2=0.54
cc_4779 ( N_noxref_16_c_7039_n N_noxref_49_c_10623_n ) capacitor c=0.0200405f \
 //x=68.42 //y=1.665 //x2=67.85 //y2=0.995
cc_4780 ( N_noxref_16_M42_noxref_d N_noxref_49_M41_noxref_d ) capacitor \
 c=5.27807e-19 //x=68.145 //y=0.915 //x2=66.61 //y2=0.91
cc_4781 ( N_noxref_16_c_6804_n N_noxref_49_M42_noxref_s ) capacitor \
 c=0.0196084f //x=68.735 //y=1.665 //x2=67.715 //y2=0.375
cc_4782 ( N_noxref_16_M42_noxref_d N_noxref_49_M42_noxref_s ) capacitor \
 c=0.0426368f //x=68.145 //y=0.915 //x2=67.715 //y2=0.375
cc_4783 ( N_noxref_16_c_6804_n N_noxref_50_c_10659_n ) capacitor c=3.84569e-19 \
 //x=68.735 //y=1.665 //x2=70.15 //y2=1.505
cc_4784 ( N_noxref_16_M42_noxref_d N_noxref_50_M43_noxref_s ) capacitor \
 c=2.55333e-19 //x=68.145 //y=0.915 //x2=70.015 //y2=0.375
cc_4785 ( N_noxref_16_M45_noxref_d N_noxref_50_M43_noxref_s ) capacitor \
 c=0.00309936f //x=72.955 //y=0.915 //x2=70.015 //y2=0.375
cc_4786 ( N_noxref_16_c_6805_n N_noxref_51_c_10700_n ) capacitor c=0.00464291f \
 //x=73.545 //y=1.665 //x2=73.545 //y2=0.54
cc_4787 ( N_noxref_16_M45_noxref_d N_noxref_51_c_10700_n ) capacitor \
 c=0.0117407f //x=72.955 //y=0.915 //x2=73.545 //y2=0.54
cc_4788 ( N_noxref_16_c_7240_p N_noxref_51_c_10722_n ) capacitor c=0.020048f \
 //x=73.23 //y=1.665 //x2=72.66 //y2=0.995
cc_4789 ( N_noxref_16_M45_noxref_d N_noxref_51_M44_noxref_d ) capacitor \
 c=5.27807e-19 //x=72.955 //y=0.915 //x2=71.42 //y2=0.91
cc_4790 ( N_noxref_16_c_6805_n N_noxref_51_M45_noxref_s ) capacitor \
 c=0.0205269f //x=73.545 //y=1.665 //x2=72.525 //y2=0.375
cc_4791 ( N_noxref_16_M45_noxref_d N_noxref_51_M45_noxref_s ) capacitor \
 c=0.0426444f //x=72.955 //y=0.915 //x2=72.525 //y2=0.375
cc_4792 ( N_noxref_16_c_6805_n N_noxref_52_c_10765_n ) capacitor c=3.04182e-19 \
 //x=73.545 //y=1.665 //x2=75.065 //y2=1.495
cc_4793 ( N_noxref_16_c_6823_n N_noxref_52_c_10765_n ) capacitor c=0.0034165f \
 //x=75.285 //y=1.915 //x2=75.065 //y2=1.495
cc_4794 ( N_noxref_16_c_6806_n N_noxref_52_c_10747_n ) capacitor c=0.0115894f \
 //x=75.48 //y=2.08 //x2=75.95 //y2=1.58
cc_4795 ( N_noxref_16_c_6822_n N_noxref_52_c_10747_n ) capacitor c=0.00703567f \
 //x=75.285 //y=1.52 //x2=75.95 //y2=1.58
cc_4796 ( N_noxref_16_c_6823_n N_noxref_52_c_10747_n ) capacitor c=0.01939f \
 //x=75.285 //y=1.915 //x2=75.95 //y2=1.58
cc_4797 ( N_noxref_16_c_6825_n N_noxref_52_c_10747_n ) capacitor c=0.00780629f \
 //x=75.66 //y=1.365 //x2=75.95 //y2=1.58
cc_4798 ( N_noxref_16_c_6828_n N_noxref_52_c_10747_n ) capacitor c=0.00339872f \
 //x=75.815 //y=1.21 //x2=75.95 //y2=1.58
cc_4799 ( N_noxref_16_c_6823_n N_noxref_52_c_10754_n ) capacitor c=6.71402e-19 \
 //x=75.285 //y=1.915 //x2=76.035 //y2=1.495
cc_4800 ( N_noxref_16_c_7225_p N_noxref_52_c_10754_n ) capacitor c=0.00623646f \
 //x=76.255 //y=1.56 //x2=76.035 //y2=1.495
cc_4801 ( N_noxref_16_c_7199_p N_noxref_52_c_10754_n ) capacitor c=0.00174428f \
 //x=76.22 //y=2.08 //x2=76.035 //y2=1.495
cc_4802 ( N_noxref_16_c_6807_n N_noxref_52_c_10755_n ) capacitor c=0.00159235f \
 //x=76.22 //y=2.08 //x2=76.92 //y2=0.53
cc_4803 ( N_noxref_16_c_7223_p N_noxref_52_c_10755_n ) capacitor c=0.0188655f \
 //x=76.255 //y=0.905 //x2=76.92 //y2=0.53
cc_4804 ( N_noxref_16_c_7228_p N_noxref_52_c_10755_n ) capacitor c=0.00656458f \
 //x=76.785 //y=0.905 //x2=76.92 //y2=0.53
cc_4805 ( N_noxref_16_c_7199_p N_noxref_52_c_10755_n ) capacitor c=2.1838e-19 \
 //x=76.22 //y=2.08 //x2=76.92 //y2=0.53
cc_4806 ( N_noxref_16_c_6819_n N_noxref_52_M46_noxref_s ) capacitor \
 c=0.0327502f //x=75.285 //y=0.865 //x2=74.93 //y2=0.365
cc_4807 ( N_noxref_16_c_6822_n N_noxref_52_M46_noxref_s ) capacitor \
 c=3.48408e-19 //x=75.285 //y=1.52 //x2=74.93 //y2=0.365
cc_4808 ( N_noxref_16_c_6826_n N_noxref_52_M46_noxref_s ) capacitor \
 c=0.0120759f //x=75.815 //y=0.865 //x2=74.93 //y2=0.365
cc_4809 ( N_noxref_16_c_7223_p N_noxref_52_M46_noxref_s ) capacitor \
 c=0.00623646f //x=76.255 //y=0.905 //x2=74.93 //y2=0.365
cc_4810 ( N_noxref_16_c_7228_p N_noxref_52_M46_noxref_s ) capacitor \
 c=0.0143002f //x=76.785 //y=0.905 //x2=74.93 //y2=0.365
cc_4811 ( N_noxref_16_c_7192_p N_noxref_52_M46_noxref_s ) capacitor \
 c=0.00290153f //x=76.785 //y=1.25 //x2=74.93 //y2=0.365
cc_4812 ( N_noxref_17_c_7583_n N_noxref_18_c_8076_n ) capacitor c=0.33882f \
 //x=78.325 //y=3.33 //x2=76.845 //y2=3.7
cc_4813 ( N_noxref_17_c_7583_n N_noxref_18_c_8127_n ) capacitor c=0.029444f \
 //x=78.325 //y=3.33 //x2=73.005 //y2=3.7
cc_4814 ( N_noxref_17_c_7583_n N_noxref_18_c_8077_n ) capacitor c=0.142709f \
 //x=78.325 //y=3.33 //x2=79.435 //y2=3.7
cc_4815 ( N_noxref_17_c_7363_n N_noxref_18_c_8077_n ) capacitor c=0.0367508f \
 //x=82.025 //y=4.44 //x2=79.435 //y2=3.7
cc_4816 ( N_noxref_17_c_7368_n N_noxref_18_c_8077_n ) capacitor c=0.0133548f \
 //x=78.555 //y=4.44 //x2=79.435 //y2=3.7
cc_4817 ( N_noxref_17_c_7310_n N_noxref_18_c_8077_n ) capacitor c=0.0247053f \
 //x=78.44 //y=2.08 //x2=79.435 //y2=3.7
cc_4818 ( N_noxref_17_c_7313_n N_noxref_18_c_8077_n ) capacitor c=0.00144897f \
 //x=82.14 //y=2.08 //x2=79.435 //y2=3.7
cc_4819 ( N_noxref_17_c_7583_n N_noxref_18_c_8079_n ) capacitor c=0.0266742f \
 //x=78.325 //y=3.33 //x2=77.075 //y2=3.7
cc_4820 ( N_noxref_17_c_7310_n N_noxref_18_c_8079_n ) capacitor c=5.11371e-19 \
 //x=78.44 //y=2.08 //x2=77.075 //y2=3.7
cc_4821 ( N_noxref_17_c_7363_n N_noxref_18_c_8064_n ) capacitor c=0.23799f \
 //x=82.025 //y=4.44 //x2=86.095 //y2=4.07
cc_4822 ( N_noxref_17_c_7313_n N_noxref_18_c_8064_n ) capacitor c=0.0258036f \
 //x=82.14 //y=2.08 //x2=86.095 //y2=4.07
cc_4823 ( N_noxref_17_c_7452_n N_noxref_18_c_8064_n ) capacitor c=0.00381677f \
 //x=82.14 //y=4.705 //x2=86.095 //y2=4.07
cc_4824 ( N_noxref_17_c_7363_n N_noxref_18_c_8085_n ) capacitor c=0.0289488f \
 //x=82.025 //y=4.44 //x2=79.665 //y2=4.07
cc_4825 ( N_noxref_17_c_7310_n N_noxref_18_c_8085_n ) capacitor c=0.0032662f \
 //x=78.44 //y=2.08 //x2=79.665 //y2=4.07
cc_4826 ( N_noxref_17_c_7583_n N_noxref_18_c_8065_n ) capacitor c=0.0198536f \
 //x=78.325 //y=3.33 //x2=72.89 //y2=2.08
cc_4827 ( N_noxref_17_c_7583_n N_noxref_18_c_8067_n ) capacitor c=0.0212814f \
 //x=78.325 //y=3.33 //x2=76.96 //y2=3.7
cc_4828 ( N_noxref_17_c_7310_n N_noxref_18_c_8067_n ) capacitor c=0.016365f \
 //x=78.44 //y=2.08 //x2=76.96 //y2=3.7
cc_4829 ( N_noxref_17_c_7363_n N_noxref_18_c_8099_n ) capacitor c=0.00210648f \
 //x=82.025 //y=4.44 //x2=79.55 //y2=4.54
cc_4830 ( N_noxref_17_c_7310_n N_noxref_18_c_8099_n ) capacitor c=0.00227044f \
 //x=78.44 //y=2.08 //x2=79.55 //y2=4.54
cc_4831 ( N_noxref_17_c_7875_p N_noxref_18_c_8099_n ) capacitor c=0.00155256f \
 //x=79.075 //y=4.795 //x2=79.55 //y2=4.54
cc_4832 ( N_noxref_17_c_7449_n N_noxref_18_c_8099_n ) capacitor c=0.00180548f \
 //x=78.785 //y=4.795 //x2=79.55 //y2=4.54
cc_4833 ( N_noxref_17_c_7583_n N_noxref_18_c_8068_n ) capacitor c=0.00431181f \
 //x=78.325 //y=3.33 //x2=79.55 //y2=2.08
cc_4834 ( N_noxref_17_c_7363_n N_noxref_18_c_8068_n ) capacitor c=0.0232321f \
 //x=82.025 //y=4.44 //x2=79.55 //y2=2.08
cc_4835 ( N_noxref_17_c_7368_n N_noxref_18_c_8068_n ) capacitor c=9.10428e-19 \
 //x=78.555 //y=4.44 //x2=79.55 //y2=2.08
cc_4836 ( N_noxref_17_c_7310_n N_noxref_18_c_8068_n ) capacitor c=0.0455851f \
 //x=78.44 //y=2.08 //x2=79.55 //y2=2.08
cc_4837 ( N_noxref_17_c_7313_n N_noxref_18_c_8068_n ) capacitor c=0.00873163f \
 //x=82.14 //y=2.08 //x2=79.55 //y2=2.08
cc_4838 ( N_noxref_17_c_7354_n N_noxref_18_c_8068_n ) capacitor c=0.00236728f \
 //x=78.44 //y=2.08 //x2=79.55 //y2=2.08
cc_4839 ( N_noxref_17_M150_noxref_g N_noxref_18_M152_noxref_g ) capacitor \
 c=0.010584f //x=78.71 //y=6.025 //x2=79.59 //y2=6.025
cc_4840 ( N_noxref_17_M151_noxref_g N_noxref_18_M152_noxref_g ) capacitor \
 c=0.106414f //x=79.15 //y=6.025 //x2=79.59 //y2=6.025
cc_4841 ( N_noxref_17_M151_noxref_g N_noxref_18_M153_noxref_g ) capacitor \
 c=0.0102479f //x=79.15 //y=6.025 //x2=80.03 //y2=6.025
cc_4842 ( N_noxref_17_c_7335_n N_noxref_18_c_8250_n ) capacitor c=4.86506e-19 \
 //x=78.615 //y=0.865 //x2=79.585 //y2=0.905
cc_4843 ( N_noxref_17_c_7337_n N_noxref_18_c_8250_n ) capacitor c=0.00152104f \
 //x=78.615 //y=1.21 //x2=79.585 //y2=0.905
cc_4844 ( N_noxref_17_c_7342_n N_noxref_18_c_8250_n ) capacitor c=0.0151475f \
 //x=79.145 //y=0.865 //x2=79.585 //y2=0.905
cc_4845 ( N_noxref_17_c_7338_n N_noxref_18_c_8253_n ) capacitor c=0.00109982f \
 //x=78.615 //y=1.52 //x2=79.585 //y2=1.25
cc_4846 ( N_noxref_17_c_7344_n N_noxref_18_c_8253_n ) capacitor c=0.0111064f \
 //x=79.145 //y=1.21 //x2=79.585 //y2=1.25
cc_4847 ( N_noxref_17_c_7338_n N_noxref_18_c_8255_n ) capacitor c=0.00179029f \
 //x=78.615 //y=1.52 //x2=79.585 //y2=1.56
cc_4848 ( N_noxref_17_c_7339_n N_noxref_18_c_8255_n ) capacitor c=0.00662747f \
 //x=78.615 //y=1.915 //x2=79.585 //y2=1.56
cc_4849 ( N_noxref_17_c_7344_n N_noxref_18_c_8255_n ) capacitor c=0.00862358f \
 //x=79.145 //y=1.21 //x2=79.585 //y2=1.56
cc_4850 ( N_noxref_17_c_7363_n N_noxref_18_c_8114_n ) capacitor c=0.0069773f \
 //x=82.025 //y=4.44 //x2=79.955 //y2=4.795
cc_4851 ( N_noxref_17_c_7342_n N_noxref_18_c_8259_n ) capacitor c=0.00124846f \
 //x=79.145 //y=0.865 //x2=80.115 //y2=0.905
cc_4852 ( N_noxref_17_c_7344_n N_noxref_18_c_8260_n ) capacitor c=0.00168739f \
 //x=79.145 //y=1.21 //x2=80.115 //y2=1.25
cc_4853 ( N_noxref_17_c_7310_n N_noxref_18_c_8072_n ) capacitor c=0.00224607f \
 //x=78.44 //y=2.08 //x2=79.55 //y2=2.08
cc_4854 ( N_noxref_17_c_7354_n N_noxref_18_c_8072_n ) capacitor c=0.00942627f \
 //x=78.44 //y=2.08 //x2=79.55 //y2=2.08
cc_4855 ( N_noxref_17_c_7363_n N_noxref_18_c_8115_n ) capacitor c=0.0014023f \
 //x=82.025 //y=4.44 //x2=79.59 //y2=4.705
cc_4856 ( N_noxref_17_c_7310_n N_noxref_18_c_8115_n ) capacitor c=0.00228787f \
 //x=78.44 //y=2.08 //x2=79.59 //y2=4.705
cc_4857 ( N_noxref_17_c_7875_p N_noxref_18_c_8115_n ) capacitor c=0.0201611f \
 //x=79.075 //y=4.795 //x2=79.59 //y2=4.705
cc_4858 ( N_noxref_17_c_7449_n N_noxref_18_c_8115_n ) capacitor c=0.00447195f \
 //x=78.785 //y=4.795 //x2=79.59 //y2=4.705
cc_4859 ( N_noxref_17_c_7363_n N_noxref_19_c_8424_n ) capacitor c=0.0856654f \
 //x=82.025 //y=4.44 //x2=81.695 //y2=5.21
cc_4860 ( N_noxref_17_M154_noxref_g N_noxref_19_c_8424_n ) capacitor \
 c=0.00503498f //x=82.03 //y=6.025 //x2=81.695 //y2=5.21
cc_4861 ( N_noxref_17_c_7363_n N_noxref_19_c_8430_n ) capacitor c=0.0130311f \
 //x=82.025 //y=4.44 //x2=79.925 //y2=5.21
cc_4862 ( N_noxref_17_c_7363_n N_noxref_19_c_8435_n ) capacitor c=0.00145992f \
 //x=82.025 //y=4.44 //x2=79.725 //y2=5.21
cc_4863 ( N_noxref_17_M151_noxref_g N_noxref_19_c_8435_n ) capacitor \
 c=0.0169795f //x=79.15 //y=6.025 //x2=79.725 //y2=5.21
cc_4864 ( N_noxref_17_c_7363_n N_noxref_19_c_8439_n ) capacitor c=0.0197096f \
 //x=82.025 //y=4.44 //x2=79.015 //y2=5.21
cc_4865 ( N_noxref_17_M150_noxref_g N_noxref_19_c_8439_n ) capacitor \
 c=0.0172236f //x=78.71 //y=6.025 //x2=79.015 //y2=5.21
cc_4866 ( N_noxref_17_c_7875_p N_noxref_19_c_8439_n ) capacitor c=0.00405363f \
 //x=79.075 //y=4.795 //x2=79.015 //y2=5.21
cc_4867 ( N_noxref_17_c_7363_n N_noxref_19_c_8441_n ) capacitor c=0.00467548f \
 //x=82.025 //y=4.44 //x2=79.81 //y2=5.295
cc_4868 ( N_noxref_17_c_7363_n N_noxref_19_c_8444_n ) capacitor c=0.00439121f \
 //x=82.025 //y=4.44 //x2=81.81 //y2=5.21
cc_4869 ( N_noxref_17_M154_noxref_g N_noxref_19_c_8444_n ) capacitor \
 c=0.0481665f //x=82.03 //y=6.025 //x2=81.81 //y2=5.21
cc_4870 ( N_noxref_17_c_7363_n N_noxref_19_c_8470_n ) capacitor c=0.00249667f \
 //x=82.025 //y=4.44 //x2=82.605 //y2=6.91
cc_4871 ( N_noxref_17_c_7313_n N_noxref_19_c_8470_n ) capacitor c=8.81369e-19 \
 //x=82.14 //y=2.08 //x2=82.605 //y2=6.91
cc_4872 ( N_noxref_17_M154_noxref_g N_noxref_19_c_8470_n ) capacitor \
 c=0.0163949f //x=82.03 //y=6.025 //x2=82.605 //y2=6.91
cc_4873 ( N_noxref_17_M155_noxref_g N_noxref_19_c_8470_n ) capacitor \
 c=0.0150104f //x=82.47 //y=6.025 //x2=82.605 //y2=6.91
cc_4874 ( N_noxref_17_M151_noxref_g N_noxref_19_M150_noxref_d ) capacitor \
 c=0.0169879f //x=79.15 //y=6.025 //x2=78.785 //y2=5.025
cc_4875 ( N_noxref_17_M155_noxref_g N_noxref_19_M155_noxref_d ) capacitor \
 c=0.0130327f //x=82.47 //y=6.025 //x2=82.545 //y2=5.025
cc_4876 ( N_noxref_17_c_7491_n N_noxref_20_c_8516_n ) capacitor c=0.336622f \
 //x=50.945 //y=3.33 //x2=83.505 //y2=2.96
cc_4877 ( N_noxref_17_c_7495_n N_noxref_20_c_8516_n ) capacitor c=0.0291389f \
 //x=47.105 //y=3.33 //x2=83.505 //y2=2.96
cc_4878 ( N_noxref_17_c_7362_n N_noxref_20_c_8516_n ) capacitor c=0.338403f \
 //x=55.015 //y=3.33 //x2=83.505 //y2=2.96
cc_4879 ( N_noxref_17_c_7529_n N_noxref_20_c_8516_n ) capacitor c=0.0266415f \
 //x=51.175 //y=3.33 //x2=83.505 //y2=2.96
cc_4880 ( N_noxref_17_c_7559_n N_noxref_20_c_8516_n ) capacitor c=0.466581f \
 //x=60.565 //y=3.33 //x2=83.505 //y2=2.96
cc_4881 ( N_noxref_17_c_7561_n N_noxref_20_c_8516_n ) capacitor c=0.0264915f \
 //x=55.245 //y=3.33 //x2=83.505 //y2=2.96
cc_4882 ( N_noxref_17_c_7648_n N_noxref_20_c_8516_n ) capacitor c=0.144314f \
 //x=62.415 //y=3.33 //x2=83.505 //y2=2.96
cc_4883 ( N_noxref_17_c_7649_n N_noxref_20_c_8516_n ) capacitor c=0.0266688f \
 //x=60.795 //y=3.33 //x2=83.505 //y2=2.96
cc_4884 ( N_noxref_17_c_7650_n N_noxref_20_c_8516_n ) capacitor c=0.108685f \
 //x=63.895 //y=3.33 //x2=83.505 //y2=2.96
cc_4885 ( N_noxref_17_c_7651_n N_noxref_20_c_8516_n ) capacitor c=0.0265703f \
 //x=62.645 //y=3.33 //x2=83.505 //y2=2.96
cc_4886 ( N_noxref_17_c_7652_n N_noxref_20_c_8516_n ) capacitor c=0.14468f \
 //x=65.745 //y=3.33 //x2=83.505 //y2=2.96
cc_4887 ( N_noxref_17_c_7653_n N_noxref_20_c_8516_n ) capacitor c=0.0266415f \
 //x=64.125 //y=3.33 //x2=83.505 //y2=2.96
cc_4888 ( N_noxref_17_c_7583_n N_noxref_20_c_8516_n ) capacitor c=1.11237f \
 //x=78.325 //y=3.33 //x2=83.505 //y2=2.96
cc_4889 ( N_noxref_17_c_7584_n N_noxref_20_c_8516_n ) capacitor c=0.0265971f \
 //x=65.975 //y=3.33 //x2=83.505 //y2=2.96
cc_4890 ( N_noxref_17_c_7363_n N_noxref_20_c_8516_n ) capacitor c=0.0132753f \
 //x=82.025 //y=4.44 //x2=83.505 //y2=2.96
cc_4891 ( N_noxref_17_c_7301_n N_noxref_20_c_8516_n ) capacitor c=0.0198264f \
 //x=46.99 //y=2.08 //x2=83.505 //y2=2.96
cc_4892 ( N_noxref_17_c_7303_n N_noxref_20_c_8516_n ) capacitor c=0.0205752f \
 //x=51.06 //y=3.33 //x2=83.505 //y2=2.96
cc_4893 ( N_noxref_17_c_7304_n N_noxref_20_c_8516_n ) capacitor c=0.0198264f \
 //x=55.13 //y=2.08 //x2=83.505 //y2=2.96
cc_4894 ( N_noxref_17_c_7399_n N_noxref_20_c_8516_n ) capacitor c=0.0229319f \
 //x=60.68 //y=3.33 //x2=83.505 //y2=2.96
cc_4895 ( N_noxref_17_c_7306_n N_noxref_20_c_8516_n ) capacitor c=0.0228696f \
 //x=62.53 //y=2.08 //x2=83.505 //y2=2.96
cc_4896 ( N_noxref_17_c_7308_n N_noxref_20_c_8516_n ) capacitor c=0.0229357f \
 //x=64.01 //y=3.33 //x2=83.505 //y2=2.96
cc_4897 ( N_noxref_17_c_7309_n N_noxref_20_c_8516_n ) capacitor c=0.02391f \
 //x=65.86 //y=2.08 //x2=83.505 //y2=2.96
cc_4898 ( N_noxref_17_c_7310_n N_noxref_20_c_8516_n ) capacitor c=0.0258141f \
 //x=78.44 //y=2.08 //x2=83.505 //y2=2.96
cc_4899 ( N_noxref_17_c_7313_n N_noxref_20_c_8516_n ) capacitor c=0.0289771f \
 //x=82.14 //y=2.08 //x2=83.505 //y2=2.96
cc_4900 ( N_noxref_17_c_7348_n N_noxref_20_c_8516_n ) capacitor c=0.00383621f \
 //x=81.945 //y=1.915 //x2=83.505 //y2=2.96
cc_4901 ( N_noxref_17_c_7354_n N_noxref_20_c_8516_n ) capacitor c=0.00409269f \
 //x=78.44 //y=2.08 //x2=83.505 //y2=2.96
cc_4902 ( N_noxref_17_c_7313_n N_noxref_20_c_8537_n ) capacitor c=0.00622935f \
 //x=82.14 //y=2.08 //x2=83.735 //y2=2.08
cc_4903 ( N_noxref_17_c_7363_n N_noxref_20_c_8541_n ) capacitor c=0.00408068f \
 //x=82.025 //y=4.44 //x2=83.62 //y2=2.08
cc_4904 ( N_noxref_17_c_7313_n N_noxref_20_c_8541_n ) capacitor c=0.0343626f \
 //x=82.14 //y=2.08 //x2=83.62 //y2=2.08
cc_4905 ( N_noxref_17_c_7348_n N_noxref_20_c_8541_n ) capacitor c=2.35599e-19 \
 //x=81.945 //y=1.915 //x2=83.62 //y2=2.08
cc_4906 ( N_noxref_17_c_7452_n N_noxref_20_c_8541_n ) capacitor c=2.35599e-19 \
 //x=82.14 //y=4.705 //x2=83.62 //y2=2.08
cc_4907 ( N_noxref_17_c_7313_n N_noxref_20_c_8543_n ) capacitor c=5.76627e-19 \
 //x=82.14 //y=2.08 //x2=85.1 //y2=2.08
cc_4908 ( N_noxref_17_M154_noxref_g N_noxref_20_M156_noxref_g ) capacitor \
 c=0.009459f //x=82.03 //y=6.025 //x2=82.91 //y2=6.025
cc_4909 ( N_noxref_17_M155_noxref_g N_noxref_20_M156_noxref_g ) capacitor \
 c=0.0626756f //x=82.47 //y=6.025 //x2=82.91 //y2=6.025
cc_4910 ( N_noxref_17_M155_noxref_g N_noxref_20_M157_noxref_g ) capacitor \
 c=0.00899012f //x=82.47 //y=6.025 //x2=83.35 //y2=6.025
cc_4911 ( N_noxref_17_c_7345_n N_noxref_20_c_8825_n ) capacitor c=4.86506e-19 \
 //x=81.945 //y=0.865 //x2=82.915 //y2=0.905
cc_4912 ( N_noxref_17_c_7347_n N_noxref_20_c_8825_n ) capacitor c=0.00101233f \
 //x=81.945 //y=1.21 //x2=82.915 //y2=0.905
cc_4913 ( N_noxref_17_c_7351_n N_noxref_20_c_8825_n ) capacitor c=0.0168844f \
 //x=82.475 //y=0.865 //x2=82.915 //y2=0.905
cc_4914 ( N_noxref_17_c_7958_p N_noxref_20_c_8828_n ) capacitor c=7.88071e-19 \
 //x=81.945 //y=1.52 //x2=82.915 //y2=1.25
cc_4915 ( N_noxref_17_c_7353_n N_noxref_20_c_8828_n ) capacitor c=0.0168218f \
 //x=82.475 //y=1.21 //x2=82.915 //y2=1.25
cc_4916 ( N_noxref_17_c_7313_n N_noxref_20_c_8830_n ) capacitor c=9.39431e-19 \
 //x=82.14 //y=2.08 //x2=82.985 //y2=4.795
cc_4917 ( N_noxref_17_c_7452_n N_noxref_20_c_8830_n ) capacitor c=0.0634092f \
 //x=82.14 //y=4.705 //x2=82.985 //y2=4.795
cc_4918 ( N_noxref_17_c_7313_n N_noxref_20_c_8584_n ) capacitor c=2.35599e-19 \
 //x=82.14 //y=2.08 //x2=83.35 //y2=4.87
cc_4919 ( N_noxref_17_c_7452_n N_noxref_20_c_8584_n ) capacitor c=5.35364e-19 \
 //x=82.14 //y=4.705 //x2=83.35 //y2=4.87
cc_4920 ( N_noxref_17_c_7351_n N_noxref_20_c_8834_n ) capacitor c=0.00124821f \
 //x=82.475 //y=0.865 //x2=83.445 //y2=0.905
cc_4921 ( N_noxref_17_c_7353_n N_noxref_20_c_8835_n ) capacitor c=8.19575e-19 \
 //x=82.475 //y=1.21 //x2=83.445 //y2=1.25
cc_4922 ( N_noxref_17_c_7353_n N_noxref_20_c_8836_n ) capacitor c=3.60397e-19 \
 //x=82.475 //y=1.21 //x2=83.445 //y2=1.56
cc_4923 ( N_noxref_17_c_7348_n N_noxref_20_c_8544_n ) capacitor c=4.61972e-19 \
 //x=81.945 //y=1.915 //x2=83.445 //y2=1.915
cc_4924 ( N_noxref_17_M155_noxref_g N_noxref_21_c_9023_n ) capacitor \
 c=0.0179287f //x=82.47 //y=6.025 //x2=83.045 //y2=5.21
cc_4925 ( N_noxref_17_c_7363_n N_noxref_21_c_9014_n ) capacitor c=0.0021588f \
 //x=82.025 //y=4.44 //x2=82.335 //y2=5.21
cc_4926 ( N_noxref_17_c_7313_n N_noxref_21_c_9014_n ) capacitor c=0.0056513f \
 //x=82.14 //y=2.08 //x2=82.335 //y2=5.21
cc_4927 ( N_noxref_17_M154_noxref_g N_noxref_21_c_9014_n ) capacitor \
 c=0.0132827f //x=82.03 //y=6.025 //x2=82.335 //y2=5.21
cc_4928 ( N_noxref_17_c_7452_n N_noxref_21_c_9014_n ) capacitor c=0.00554802f \
 //x=82.14 //y=4.705 //x2=82.335 //y2=5.21
cc_4929 ( N_noxref_17_M155_noxref_g N_noxref_21_M154_noxref_d ) capacitor \
 c=0.0130327f //x=82.47 //y=6.025 //x2=82.105 //y2=5.025
cc_4930 ( N_noxref_17_c_7347_n N_QN_c_9097_n ) capacitor c=0.00500281f \
 //x=81.945 //y=1.21 //x2=83.065 //y2=1.18
cc_4931 ( N_noxref_17_c_7958_p N_QN_c_9097_n ) capacitor c=0.00342096f \
 //x=81.945 //y=1.52 //x2=83.065 //y2=1.18
cc_4932 ( N_noxref_17_c_7349_n N_QN_c_9097_n ) capacitor c=4.02408e-19 \
 //x=82.32 //y=0.71 //x2=83.065 //y2=1.18
cc_4933 ( N_noxref_17_c_7350_n N_QN_c_9097_n ) capacitor c=0.0032199f \
 //x=82.32 //y=1.365 //x2=83.065 //y2=1.18
cc_4934 ( N_noxref_17_c_7353_n N_QN_c_9097_n ) capacitor c=0.00735559f \
 //x=82.475 //y=1.21 //x2=83.065 //y2=1.18
cc_4935 ( N_noxref_17_c_7301_n N_noxref_41_c_10190_n ) capacitor c=0.00204385f \
 //x=46.99 //y=2.08 //x2=47.645 //y2=0.54
cc_4936 ( N_noxref_17_c_7510_n N_noxref_41_c_10190_n ) capacitor c=0.0194423f \
 //x=46.98 //y=0.915 //x2=47.645 //y2=0.54
cc_4937 ( N_noxref_17_c_7516_n N_noxref_41_c_10190_n ) capacitor c=0.00656458f \
 //x=47.51 //y=0.915 //x2=47.645 //y2=0.54
cc_4938 ( N_noxref_17_c_7519_n N_noxref_41_c_10190_n ) capacitor c=2.20712e-19 \
 //x=46.99 //y=2.08 //x2=47.645 //y2=0.54
cc_4939 ( N_noxref_17_c_7511_n N_noxref_41_c_10200_n ) capacitor c=0.00538829f \
 //x=46.98 //y=1.26 //x2=46.76 //y2=0.995
cc_4940 ( N_noxref_17_c_7510_n N_noxref_41_M29_noxref_s ) capacitor \
 c=0.00538829f //x=46.98 //y=0.915 //x2=46.625 //y2=0.375
cc_4941 ( N_noxref_17_c_7512_n N_noxref_41_M29_noxref_s ) capacitor \
 c=0.00538829f //x=46.98 //y=1.57 //x2=46.625 //y2=0.375
cc_4942 ( N_noxref_17_c_7516_n N_noxref_41_M29_noxref_s ) capacitor \
 c=0.0143002f //x=47.51 //y=0.915 //x2=46.625 //y2=0.375
cc_4943 ( N_noxref_17_c_7517_n N_noxref_41_M29_noxref_s ) capacitor \
 c=0.00290153f //x=47.51 //y=1.26 //x2=46.625 //y2=0.375
cc_4944 ( N_noxref_17_c_7713_n N_noxref_42_c_10255_n ) capacitor c=3.15806e-19 \
 //x=50.705 //y=1.655 //x2=49.165 //y2=1.495
cc_4945 ( N_noxref_17_c_7713_n N_noxref_42_c_10244_n ) capacitor c=0.020324f \
 //x=50.705 //y=1.655 //x2=50.135 //y2=1.495
cc_4946 ( N_noxref_17_c_7302_n N_noxref_42_c_10245_n ) capacitor c=0.00457164f \
 //x=50.975 //y=1.655 //x2=51.02 //y2=0.53
cc_4947 ( N_noxref_17_M31_noxref_d N_noxref_42_c_10245_n ) capacitor \
 c=0.0115831f //x=50.43 //y=0.905 //x2=51.02 //y2=0.53
cc_4948 ( N_noxref_17_c_7302_n N_noxref_42_M30_noxref_s ) capacitor \
 c=0.013435f //x=50.975 //y=1.655 //x2=49.03 //y2=0.365
cc_4949 ( N_noxref_17_M31_noxref_d N_noxref_42_M30_noxref_s ) capacitor \
 c=0.0439476f //x=50.43 //y=0.905 //x2=49.03 //y2=0.365
cc_4950 ( N_noxref_17_c_7302_n N_noxref_43_c_10312_n ) capacitor c=4.08644e-19 \
 //x=50.975 //y=1.655 //x2=52.39 //y2=1.505
cc_4951 ( N_noxref_17_M31_noxref_d N_noxref_43_M32_noxref_s ) capacitor \
 c=2.53688e-19 //x=50.43 //y=0.905 //x2=52.255 //y2=0.375
cc_4952 ( N_noxref_17_c_7304_n N_noxref_44_c_10342_n ) capacitor c=0.00204385f \
 //x=55.13 //y=2.08 //x2=55.785 //y2=0.54
cc_4953 ( N_noxref_17_c_7614_n N_noxref_44_c_10342_n ) capacitor c=0.0194423f \
 //x=55.12 //y=0.915 //x2=55.785 //y2=0.54
cc_4954 ( N_noxref_17_c_7680_n N_noxref_44_c_10342_n ) capacitor c=0.00656458f \
 //x=55.65 //y=0.915 //x2=55.785 //y2=0.54
cc_4955 ( N_noxref_17_c_7633_n N_noxref_44_c_10342_n ) capacitor c=2.20712e-19 \
 //x=55.13 //y=2.08 //x2=55.785 //y2=0.54
cc_4956 ( N_noxref_17_c_7615_n N_noxref_44_c_10364_n ) capacitor c=0.00538829f \
 //x=55.12 //y=1.26 //x2=54.9 //y2=0.995
cc_4957 ( N_noxref_17_c_7614_n N_noxref_44_M34_noxref_s ) capacitor \
 c=0.00538829f //x=55.12 //y=0.915 //x2=54.765 //y2=0.375
cc_4958 ( N_noxref_17_c_7616_n N_noxref_44_M34_noxref_s ) capacitor \
 c=0.00538829f //x=55.12 //y=1.57 //x2=54.765 //y2=0.375
cc_4959 ( N_noxref_17_c_7680_n N_noxref_44_M34_noxref_s ) capacitor \
 c=0.0143002f //x=55.65 //y=0.915 //x2=54.765 //y2=0.375
cc_4960 ( N_noxref_17_c_7681_n N_noxref_44_M34_noxref_s ) capacitor \
 c=0.00290153f //x=55.65 //y=1.26 //x2=54.765 //y2=0.375
cc_4961 ( N_noxref_17_M37_noxref_d N_noxref_45_M35_noxref_s ) capacitor \
 c=0.00309936f //x=60.005 //y=0.915 //x2=57.065 //y2=0.375
cc_4962 ( N_noxref_17_c_7305_n N_noxref_46_c_10443_n ) capacitor c=0.00457167f \
 //x=60.595 //y=1.665 //x2=60.595 //y2=0.54
cc_4963 ( N_noxref_17_M37_noxref_d N_noxref_46_c_10443_n ) capacitor \
 c=0.0115903f //x=60.005 //y=0.915 //x2=60.595 //y2=0.54
cc_4964 ( N_noxref_17_c_7721_n N_noxref_46_c_10470_n ) capacitor c=0.020048f \
 //x=60.28 //y=1.665 //x2=59.71 //y2=0.995
cc_4965 ( N_noxref_17_M37_noxref_d N_noxref_46_M36_noxref_d ) capacitor \
 c=5.27807e-19 //x=60.005 //y=0.915 //x2=58.47 //y2=0.91
cc_4966 ( N_noxref_17_c_7305_n N_noxref_46_M37_noxref_s ) capacitor \
 c=0.0196084f //x=60.595 //y=1.665 //x2=59.575 //y2=0.375
cc_4967 ( N_noxref_17_M37_noxref_d N_noxref_46_M37_noxref_s ) capacitor \
 c=0.0426444f //x=60.005 //y=0.915 //x2=59.575 //y2=0.375
cc_4968 ( N_noxref_17_c_7305_n N_noxref_47_c_10509_n ) capacitor c=3.04182e-19 \
 //x=60.595 //y=1.665 //x2=62.115 //y2=1.495
cc_4969 ( N_noxref_17_c_7730_n N_noxref_47_c_10509_n ) capacitor c=3.15806e-19 \
 //x=63.655 //y=1.655 //x2=62.115 //y2=1.495
cc_4970 ( N_noxref_17_c_7319_n N_noxref_47_c_10509_n ) capacitor c=0.0034165f \
 //x=62.335 //y=1.915 //x2=62.115 //y2=1.495
cc_4971 ( N_noxref_17_c_7306_n N_noxref_47_c_10491_n ) capacitor c=0.011618f \
 //x=62.53 //y=2.08 //x2=63 //y2=1.58
cc_4972 ( N_noxref_17_c_7318_n N_noxref_47_c_10491_n ) capacitor c=0.00696403f \
 //x=62.335 //y=1.52 //x2=63 //y2=1.58
cc_4973 ( N_noxref_17_c_7319_n N_noxref_47_c_10491_n ) capacitor c=0.0174694f \
 //x=62.335 //y=1.915 //x2=63 //y2=1.58
cc_4974 ( N_noxref_17_c_7321_n N_noxref_47_c_10491_n ) capacitor c=0.00776811f \
 //x=62.71 //y=1.365 //x2=63 //y2=1.58
cc_4975 ( N_noxref_17_c_7324_n N_noxref_47_c_10491_n ) capacitor c=0.00339872f \
 //x=62.865 //y=1.21 //x2=63 //y2=1.58
cc_4976 ( N_noxref_17_c_7730_n N_noxref_47_c_10498_n ) capacitor c=0.020324f \
 //x=63.655 //y=1.655 //x2=63.085 //y2=1.495
cc_4977 ( N_noxref_17_c_7319_n N_noxref_47_c_10498_n ) capacitor c=6.71402e-19 \
 //x=62.335 //y=1.915 //x2=63.085 //y2=1.495
cc_4978 ( N_noxref_17_c_7307_n N_noxref_47_c_10499_n ) capacitor c=0.00457164f \
 //x=63.925 //y=1.655 //x2=63.97 //y2=0.53
cc_4979 ( N_noxref_17_M39_noxref_d N_noxref_47_c_10499_n ) capacitor \
 c=0.0115831f //x=63.38 //y=0.905 //x2=63.97 //y2=0.53
cc_4980 ( N_noxref_17_c_7307_n N_noxref_47_M38_noxref_s ) capacitor \
 c=0.013435f //x=63.925 //y=1.655 //x2=61.98 //y2=0.365
cc_4981 ( N_noxref_17_c_7315_n N_noxref_47_M38_noxref_s ) capacitor \
 c=0.0327502f //x=62.335 //y=0.865 //x2=61.98 //y2=0.365
cc_4982 ( N_noxref_17_c_7318_n N_noxref_47_M38_noxref_s ) capacitor \
 c=3.48408e-19 //x=62.335 //y=1.52 //x2=61.98 //y2=0.365
cc_4983 ( N_noxref_17_c_7322_n N_noxref_47_M38_noxref_s ) capacitor \
 c=0.0120759f //x=62.865 //y=0.865 //x2=61.98 //y2=0.365
cc_4984 ( N_noxref_17_M39_noxref_d N_noxref_47_M38_noxref_s ) capacitor \
 c=0.0439476f //x=63.38 //y=0.905 //x2=61.98 //y2=0.365
cc_4985 ( N_noxref_17_c_7307_n N_noxref_48_c_10565_n ) capacitor c=4.08644e-19 \
 //x=63.925 //y=1.655 //x2=65.34 //y2=1.505
cc_4986 ( N_noxref_17_c_7329_n N_noxref_48_c_10565_n ) capacitor c=0.0034165f \
 //x=65.56 //y=1.915 //x2=65.34 //y2=1.505
cc_4987 ( N_noxref_17_c_7309_n N_noxref_48_c_10542_n ) capacitor c=0.0115578f \
 //x=65.86 //y=2.08 //x2=66.225 //y2=1.59
cc_4988 ( N_noxref_17_c_7328_n N_noxref_48_c_10542_n ) capacitor c=0.00697148f \
 //x=65.56 //y=1.53 //x2=66.225 //y2=1.59
cc_4989 ( N_noxref_17_c_7329_n N_noxref_48_c_10542_n ) capacitor c=0.0204849f \
 //x=65.56 //y=1.915 //x2=66.225 //y2=1.59
cc_4990 ( N_noxref_17_c_7331_n N_noxref_48_c_10542_n ) capacitor c=0.00610316f \
 //x=65.935 //y=1.375 //x2=66.225 //y2=1.59
cc_4991 ( N_noxref_17_c_7334_n N_noxref_48_c_10542_n ) capacitor c=0.00698822f \
 //x=66.09 //y=1.22 //x2=66.225 //y2=1.59
cc_4992 ( N_noxref_17_c_7325_n N_noxref_48_M40_noxref_s ) capacitor \
 c=0.0327271f //x=65.56 //y=0.875 //x2=65.205 //y2=0.375
cc_4993 ( N_noxref_17_c_7328_n N_noxref_48_M40_noxref_s ) capacitor \
 c=7.99997e-19 //x=65.56 //y=1.53 //x2=65.205 //y2=0.375
cc_4994 ( N_noxref_17_c_7329_n N_noxref_48_M40_noxref_s ) capacitor \
 c=0.00122123f //x=65.56 //y=1.915 //x2=65.205 //y2=0.375
cc_4995 ( N_noxref_17_c_7332_n N_noxref_48_M40_noxref_s ) capacitor \
 c=0.0121427f //x=66.09 //y=0.875 //x2=65.205 //y2=0.375
cc_4996 ( N_noxref_17_M39_noxref_d N_noxref_48_M40_noxref_s ) capacitor \
 c=2.53688e-19 //x=63.38 //y=0.905 //x2=65.205 //y2=0.375
cc_4997 ( N_noxref_17_c_7310_n N_noxref_53_c_10816_n ) capacitor c=0.0160451f \
 //x=78.44 //y=2.08 //x2=78.395 //y2=1.495
cc_4998 ( N_noxref_17_c_7339_n N_noxref_53_c_10816_n ) capacitor c=0.0034165f \
 //x=78.615 //y=1.915 //x2=78.395 //y2=1.495
cc_4999 ( N_noxref_17_c_7354_n N_noxref_53_c_10816_n ) capacitor c=0.00781973f \
 //x=78.44 //y=2.08 //x2=78.395 //y2=1.495
cc_5000 ( N_noxref_17_c_7310_n N_noxref_53_c_10798_n ) capacitor c=0.00513915f \
 //x=78.44 //y=2.08 //x2=79.28 //y2=1.58
cc_5001 ( N_noxref_17_c_7338_n N_noxref_53_c_10798_n ) capacitor c=0.00720513f \
 //x=78.615 //y=1.52 //x2=79.28 //y2=1.58
cc_5002 ( N_noxref_17_c_7339_n N_noxref_53_c_10798_n ) capacitor c=0.0140339f \
 //x=78.615 //y=1.915 //x2=79.28 //y2=1.58
cc_5003 ( N_noxref_17_c_7341_n N_noxref_53_c_10798_n ) capacitor c=0.0100869f \
 //x=78.99 //y=1.365 //x2=79.28 //y2=1.58
cc_5004 ( N_noxref_17_c_7344_n N_noxref_53_c_10798_n ) capacitor c=0.00339872f \
 //x=79.145 //y=1.21 //x2=79.28 //y2=1.58
cc_5005 ( N_noxref_17_c_7354_n N_noxref_53_c_10798_n ) capacitor c=0.00324565f \
 //x=78.44 //y=2.08 //x2=79.28 //y2=1.58
cc_5006 ( N_noxref_17_c_7339_n N_noxref_53_c_10805_n ) capacitor c=6.71402e-19 \
 //x=78.615 //y=1.915 //x2=79.365 //y2=1.495
cc_5007 ( N_noxref_17_c_7335_n N_noxref_53_M48_noxref_s ) capacitor \
 c=0.0326001f //x=78.615 //y=0.865 //x2=78.26 //y2=0.365
cc_5008 ( N_noxref_17_c_7338_n N_noxref_53_M48_noxref_s ) capacitor \
 c=0.00110192f //x=78.615 //y=1.52 //x2=78.26 //y2=0.365
cc_5009 ( N_noxref_17_c_7342_n N_noxref_53_M48_noxref_s ) capacitor \
 c=0.0120759f //x=79.145 //y=0.865 //x2=78.26 //y2=0.365
cc_5010 ( N_noxref_17_c_7348_n N_noxref_54_c_10872_n ) capacitor c=0.0034165f \
 //x=81.945 //y=1.915 //x2=81.725 //y2=1.495
cc_5011 ( N_noxref_17_c_7313_n N_noxref_54_c_10855_n ) capacitor c=0.011159f \
 //x=82.14 //y=2.08 //x2=82.61 //y2=1.58
cc_5012 ( N_noxref_17_c_7958_p N_noxref_54_c_10855_n ) capacitor c=0.00598984f \
 //x=81.945 //y=1.52 //x2=82.61 //y2=1.58
cc_5013 ( N_noxref_17_c_7348_n N_noxref_54_c_10855_n ) capacitor c=0.0197952f \
 //x=81.945 //y=1.915 //x2=82.61 //y2=1.58
cc_5014 ( N_noxref_17_c_7350_n N_noxref_54_c_10855_n ) capacitor c=0.00767729f \
 //x=82.32 //y=1.365 //x2=82.61 //y2=1.58
cc_5015 ( N_noxref_17_c_7353_n N_noxref_54_c_10855_n ) capacitor c=0.0059368f \
 //x=82.475 //y=1.21 //x2=82.61 //y2=1.58
cc_5016 ( N_noxref_17_c_7348_n N_noxref_54_c_10861_n ) capacitor c=0.00122123f \
 //x=81.945 //y=1.915 //x2=82.695 //y2=1.495
cc_5017 ( N_noxref_17_c_7345_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.0312776f //x=81.945 //y=0.865 //x2=81.59 //y2=0.365
cc_5018 ( N_noxref_17_c_7958_p N_noxref_54_M50_noxref_s ) capacitor \
 c=3.48408e-19 //x=81.945 //y=1.52 //x2=81.59 //y2=0.365
cc_5019 ( N_noxref_17_c_7351_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.0132463f //x=82.475 //y=0.865 //x2=81.59 //y2=0.365
cc_5020 ( N_noxref_18_c_8064_n N_noxref_19_c_8424_n ) capacitor c=0.00923886f \
 //x=86.095 //y=4.07 //x2=81.695 //y2=5.21
cc_5021 ( N_noxref_18_M153_noxref_g N_noxref_19_c_8424_n ) capacitor \
 c=0.0104371f //x=80.03 //y=6.025 //x2=81.695 //y2=5.21
cc_5022 ( N_noxref_18_c_8064_n N_noxref_19_c_8430_n ) capacitor c=0.00122833f \
 //x=86.095 //y=4.07 //x2=79.925 //y2=5.21
cc_5023 ( N_noxref_18_M152_noxref_g N_noxref_19_c_8430_n ) capacitor \
 c=0.0010118f //x=79.59 //y=6.025 //x2=79.925 //y2=5.21
cc_5024 ( N_noxref_18_M153_noxref_g N_noxref_19_c_8430_n ) capacitor \
 c=8.30848e-19 //x=80.03 //y=6.025 //x2=79.925 //y2=5.21
cc_5025 ( N_noxref_18_c_8099_n N_noxref_19_c_8435_n ) capacitor c=0.0126743f \
 //x=79.55 //y=4.54 //x2=79.725 //y2=5.21
cc_5026 ( N_noxref_18_M152_noxref_g N_noxref_19_c_8435_n ) capacitor \
 c=0.0161605f //x=79.59 //y=6.025 //x2=79.725 //y2=5.21
cc_5027 ( N_noxref_18_c_8115_n N_noxref_19_c_8435_n ) capacitor c=0.00307538f \
 //x=79.59 //y=4.705 //x2=79.725 //y2=5.21
cc_5028 ( N_noxref_18_M152_noxref_g N_noxref_19_c_8441_n ) capacitor \
 c=0.00226657f //x=79.59 //y=6.025 //x2=79.81 //y2=5.295
cc_5029 ( N_noxref_18_M153_noxref_g N_noxref_19_c_8441_n ) capacitor \
 c=0.0197448f //x=80.03 //y=6.025 //x2=79.81 //y2=5.295
cc_5030 ( N_noxref_18_c_8114_n N_noxref_19_c_8441_n ) capacitor c=0.00458101f \
 //x=79.955 //y=4.795 //x2=79.81 //y2=5.295
cc_5031 ( N_noxref_18_M152_noxref_g N_noxref_19_M152_noxref_d ) capacitor \
 c=0.016914f //x=79.59 //y=6.025 //x2=79.665 //y2=5.025
cc_5032 ( N_noxref_18_c_8076_n N_noxref_20_c_8516_n ) capacitor c=0.0288894f \
 //x=76.845 //y=3.7 //x2=83.505 //y2=2.96
cc_5033 ( N_noxref_18_c_8127_n N_noxref_20_c_8516_n ) capacitor c=8.32553e-19 \
 //x=73.005 //y=3.7 //x2=83.505 //y2=2.96
cc_5034 ( N_noxref_18_c_8077_n N_noxref_20_c_8516_n ) capacitor c=0.0586541f \
 //x=79.435 //y=3.7 //x2=83.505 //y2=2.96
cc_5035 ( N_noxref_18_c_8079_n N_noxref_20_c_8516_n ) capacitor c=5.76918e-19 \
 //x=77.075 //y=3.7 //x2=83.505 //y2=2.96
cc_5036 ( N_noxref_18_c_8064_n N_noxref_20_c_8516_n ) capacitor c=0.123045f \
 //x=86.095 //y=4.07 //x2=83.505 //y2=2.96
cc_5037 ( N_noxref_18_c_8085_n N_noxref_20_c_8516_n ) capacitor c=6.10859e-19 \
 //x=79.665 //y=4.07 //x2=83.505 //y2=2.96
cc_5038 ( N_noxref_18_c_8065_n N_noxref_20_c_8516_n ) capacitor c=0.022447f \
 //x=72.89 //y=2.08 //x2=83.505 //y2=2.96
cc_5039 ( N_noxref_18_c_8286_p N_noxref_20_c_8516_n ) capacitor c=0.00745069f \
 //x=76.605 //y=1.655 //x2=83.505 //y2=2.96
cc_5040 ( N_noxref_18_c_8067_n N_noxref_20_c_8516_n ) capacitor c=0.0236021f \
 //x=76.96 //y=3.7 //x2=83.505 //y2=2.96
cc_5041 ( N_noxref_18_c_8068_n N_noxref_20_c_8516_n ) capacitor c=0.0270235f \
 //x=79.55 //y=2.08 //x2=83.505 //y2=2.96
cc_5042 ( N_noxref_18_c_8140_n N_noxref_20_c_8516_n ) capacitor c=0.0018311f \
 //x=72.89 //y=2.08 //x2=83.505 //y2=2.96
cc_5043 ( N_noxref_18_c_8072_n N_noxref_20_c_8516_n ) capacitor c=0.00172252f \
 //x=79.55 //y=2.08 //x2=83.505 //y2=2.96
cc_5044 ( N_noxref_18_c_8064_n N_noxref_20_c_8536_n ) capacitor c=0.0234111f \
 //x=86.095 //y=4.07 //x2=84.985 //y2=2.08
cc_5045 ( N_noxref_18_c_8070_n N_noxref_20_c_8536_n ) capacitor c=0.00668632f \
 //x=86.21 //y=2.08 //x2=84.985 //y2=2.08
cc_5046 ( N_noxref_18_c_8293_p N_noxref_20_c_8536_n ) capacitor c=0.00319611f \
 //x=86.21 //y=2.08 //x2=84.985 //y2=2.08
cc_5047 ( N_noxref_18_c_8064_n N_noxref_20_c_8541_n ) capacitor c=0.0261405f \
 //x=86.095 //y=4.07 //x2=83.62 //y2=2.08
cc_5048 ( N_noxref_18_c_8070_n N_noxref_20_c_8541_n ) capacitor c=7.56813e-19 \
 //x=86.21 //y=2.08 //x2=83.62 //y2=2.08
cc_5049 ( N_noxref_18_c_8064_n N_noxref_20_c_8543_n ) capacitor c=0.0285749f \
 //x=86.095 //y=4.07 //x2=85.1 //y2=2.08
cc_5050 ( N_noxref_18_c_8070_n N_noxref_20_c_8543_n ) capacitor c=0.0538261f \
 //x=86.21 //y=2.08 //x2=85.1 //y2=2.08
cc_5051 ( N_noxref_18_c_8293_p N_noxref_20_c_8543_n ) capacitor c=0.00207994f \
 //x=86.21 //y=2.08 //x2=85.1 //y2=2.08
cc_5052 ( N_noxref_18_c_8299_p N_noxref_20_c_8543_n ) capacitor c=0.00196222f \
 //x=86.23 //y=4.705 //x2=85.1 //y2=2.08
cc_5053 ( N_noxref_18_M160_noxref_g N_noxref_20_M158_noxref_g ) capacitor \
 c=0.00932631f //x=86.25 //y=6.025 //x2=85.37 //y2=6.025
cc_5054 ( N_noxref_18_M160_noxref_g N_noxref_20_M159_noxref_g ) capacitor \
 c=0.110179f //x=86.25 //y=6.025 //x2=85.81 //y2=6.025
cc_5055 ( N_noxref_18_M161_noxref_g N_noxref_20_M159_noxref_g ) capacitor \
 c=0.00876656f //x=86.69 //y=6.025 //x2=85.81 //y2=6.025
cc_5056 ( N_noxref_18_c_8064_n N_noxref_20_c_8830_n ) capacitor c=0.00791694f \
 //x=86.095 //y=4.07 //x2=82.985 //y2=4.795
cc_5057 ( N_noxref_18_c_8064_n N_noxref_20_c_8584_n ) capacitor c=0.0014567f \
 //x=86.095 //y=4.07 //x2=83.35 //y2=4.87
cc_5058 ( N_noxref_18_c_8305_p N_noxref_20_c_8545_n ) capacitor c=4.86506e-19 \
 //x=86.245 //y=0.905 //x2=85.275 //y2=0.865
cc_5059 ( N_noxref_18_c_8305_p N_noxref_20_c_8547_n ) capacitor c=0.00101233f \
 //x=86.245 //y=0.905 //x2=85.275 //y2=1.21
cc_5060 ( N_noxref_18_c_8307_p N_noxref_20_c_8866_n ) capacitor c=0.00257836f \
 //x=86.245 //y=1.56 //x2=85.275 //y2=1.52
cc_5061 ( N_noxref_18_c_8307_p N_noxref_20_c_8548_n ) capacitor c=0.00662747f \
 //x=86.245 //y=1.56 //x2=85.275 //y2=1.915
cc_5062 ( N_noxref_18_c_8309_p N_noxref_20_c_8868_n ) capacitor c=0.00168516f \
 //x=86.23 //y=4.705 //x2=85.735 //y2=4.795
cc_5063 ( N_noxref_18_c_8299_p N_noxref_20_c_8868_n ) capacitor c=0.0225854f \
 //x=86.23 //y=4.705 //x2=85.735 //y2=4.795
cc_5064 ( N_noxref_18_c_8064_n N_noxref_20_c_8585_n ) capacitor c=0.0117386f \
 //x=86.095 //y=4.07 //x2=85.445 //y2=4.795
cc_5065 ( N_noxref_18_c_8309_p N_noxref_20_c_8585_n ) capacitor c=0.00143876f \
 //x=86.23 //y=4.705 //x2=85.445 //y2=4.795
cc_5066 ( N_noxref_18_c_8299_p N_noxref_20_c_8585_n ) capacitor c=0.00469886f \
 //x=86.23 //y=4.705 //x2=85.445 //y2=4.795
cc_5067 ( N_noxref_18_c_8305_p N_noxref_20_c_8551_n ) capacitor c=0.0161138f \
 //x=86.245 //y=0.905 //x2=85.805 //y2=0.865
cc_5068 ( N_noxref_18_c_8315_p N_noxref_20_c_8551_n ) capacitor c=0.00130607f \
 //x=86.775 //y=0.905 //x2=85.805 //y2=0.865
cc_5069 ( N_noxref_18_c_8316_p N_noxref_20_c_8553_n ) capacitor c=0.0120728f \
 //x=86.245 //y=1.255 //x2=85.805 //y2=1.21
cc_5070 ( N_noxref_18_c_8307_p N_noxref_20_c_8553_n ) capacitor c=0.00862358f \
 //x=86.245 //y=1.56 //x2=85.805 //y2=1.21
cc_5071 ( N_noxref_18_c_8318_p N_noxref_20_c_8553_n ) capacitor c=4.4593e-19 \
 //x=86.62 //y=1.405 //x2=85.805 //y2=1.21
cc_5072 ( N_noxref_18_c_8319_p N_noxref_20_c_8553_n ) capacitor c=0.00111855f \
 //x=86.775 //y=1.255 //x2=85.805 //y2=1.21
cc_5073 ( N_noxref_18_c_8070_n N_noxref_20_c_8554_n ) capacitor c=0.00218919f \
 //x=86.21 //y=2.08 //x2=85.1 //y2=2.08
cc_5074 ( N_noxref_18_c_8293_p N_noxref_20_c_8554_n ) capacitor c=0.00908973f \
 //x=86.21 //y=2.08 //x2=85.1 //y2=2.08
cc_5075 ( N_noxref_18_c_8064_n N_noxref_21_c_9008_n ) capacitor c=0.0535575f \
 //x=86.095 //y=4.07 //x2=85.035 //y2=5.21
cc_5076 ( N_noxref_18_c_8064_n N_noxref_21_c_9012_n ) capacitor c=0.008149f \
 //x=86.095 //y=4.07 //x2=83.245 //y2=5.21
cc_5077 ( N_noxref_18_c_8064_n N_noxref_21_c_9023_n ) capacitor c=3.2507e-19 \
 //x=86.095 //y=4.07 //x2=83.045 //y2=5.21
cc_5078 ( N_noxref_18_c_8064_n N_noxref_21_c_9014_n ) capacitor c=0.0181202f \
 //x=86.095 //y=4.07 //x2=82.335 //y2=5.21
cc_5079 ( N_noxref_18_c_8064_n N_noxref_21_c_9015_n ) capacitor c=0.00337443f \
 //x=86.095 //y=4.07 //x2=83.13 //y2=5.295
cc_5080 ( N_noxref_18_c_8064_n N_noxref_21_c_9016_n ) capacitor c=0.0011253f \
 //x=86.095 //y=4.07 //x2=85.15 //y2=5.21
cc_5081 ( N_noxref_18_c_8064_n N_noxref_21_c_9035_n ) capacitor c=0.00358031f \
 //x=86.095 //y=4.07 //x2=85.945 //y2=6.91
cc_5082 ( N_noxref_18_M160_noxref_g N_noxref_21_c_9036_n ) capacitor \
 c=0.0150104f //x=86.25 //y=6.025 //x2=86.825 //y2=6.91
cc_5083 ( N_noxref_18_M161_noxref_g N_noxref_21_c_9036_n ) capacitor \
 c=0.0163361f //x=86.69 //y=6.025 //x2=86.825 //y2=6.91
cc_5084 ( N_noxref_18_M160_noxref_g N_noxref_21_M159_noxref_d ) capacitor \
 c=0.0130327f //x=86.25 //y=6.025 //x2=85.885 //y2=5.025
cc_5085 ( N_noxref_18_M161_noxref_g N_noxref_21_M161_noxref_d ) capacitor \
 c=0.0351101f //x=86.69 //y=6.025 //x2=86.765 //y2=5.025
cc_5086 ( N_noxref_18_c_8064_n N_QN_c_9097_n ) capacitor c=0.00322521f \
 //x=86.095 //y=4.07 //x2=83.065 //y2=1.18
cc_5087 ( N_noxref_18_c_8259_n N_QN_c_9097_n ) capacitor c=4.67724e-19 \
 //x=80.115 //y=0.905 //x2=83.065 //y2=1.18
cc_5088 ( N_noxref_18_c_8260_n N_QN_c_9097_n ) capacitor c=0.00732681f \
 //x=80.115 //y=1.25 //x2=83.065 //y2=1.18
cc_5089 ( N_noxref_18_c_8064_n N_QN_c_9104_n ) capacitor c=4.20225e-19 \
 //x=86.095 //y=4.07 //x2=79.965 //y2=1.18
cc_5090 ( N_noxref_18_c_8250_n N_QN_c_9104_n ) capacitor c=3.66947e-19 \
 //x=79.585 //y=0.905 //x2=79.965 //y2=1.18
cc_5091 ( N_noxref_18_c_8253_n N_QN_c_9104_n ) capacitor c=0.00353233f \
 //x=79.585 //y=1.25 //x2=79.965 //y2=1.18
cc_5092 ( N_noxref_18_c_8255_n N_QN_c_9104_n ) capacitor c=0.00289074f \
 //x=79.585 //y=1.56 //x2=79.965 //y2=1.18
cc_5093 ( N_noxref_18_c_8340_p N_QN_c_9104_n ) capacitor c=4.06815e-19 \
 //x=79.96 //y=0.75 //x2=79.965 //y2=1.18
cc_5094 ( N_noxref_18_c_8341_p N_QN_c_9104_n ) capacitor c=7.42023e-19 \
 //x=79.96 //y=1.405 //x2=79.965 //y2=1.18
cc_5095 ( N_noxref_18_c_8260_n N_QN_c_9104_n ) capacitor c=0.00133904f \
 //x=80.115 //y=1.25 //x2=79.965 //y2=1.18
cc_5096 ( N_noxref_18_c_8064_n N_QN_c_9105_n ) capacitor c=0.0113709f \
 //x=86.095 //y=4.07 //x2=86.395 //y2=1.18
cc_5097 ( N_noxref_18_c_8070_n N_QN_c_9105_n ) capacitor c=0.00449159f \
 //x=86.21 //y=2.08 //x2=86.395 //y2=1.18
cc_5098 ( N_noxref_18_c_8305_p N_QN_c_9105_n ) capacitor c=6.33948e-19 \
 //x=86.245 //y=0.905 //x2=86.395 //y2=1.18
cc_5099 ( N_noxref_18_c_8316_p N_QN_c_9105_n ) capacitor c=0.0043333f \
 //x=86.245 //y=1.255 //x2=86.395 //y2=1.18
cc_5100 ( N_noxref_18_c_8307_p N_QN_c_9105_n ) capacitor c=0.0040799f \
 //x=86.245 //y=1.56 //x2=86.395 //y2=1.18
cc_5101 ( N_noxref_18_c_8348_p N_QN_c_9105_n ) capacitor c=4.52813e-19 \
 //x=86.62 //y=0.75 //x2=86.395 //y2=1.18
cc_5102 ( N_noxref_18_c_8318_p N_QN_c_9105_n ) capacitor c=0.00296491f \
 //x=86.62 //y=1.405 //x2=86.395 //y2=1.18
cc_5103 ( N_noxref_18_c_8315_p N_QN_c_9105_n ) capacitor c=2.65983e-19 \
 //x=86.775 //y=0.905 //x2=86.395 //y2=1.18
cc_5104 ( N_noxref_18_c_8319_p N_QN_c_9105_n ) capacitor c=0.00362989f \
 //x=86.775 //y=1.255 //x2=86.395 //y2=1.18
cc_5105 ( N_noxref_18_c_8293_p N_QN_c_9105_n ) capacitor c=5.89141e-19 \
 //x=86.21 //y=2.08 //x2=86.395 //y2=1.18
cc_5106 ( N_noxref_18_c_8064_n N_QN_c_9111_n ) capacitor c=3.74512e-19 \
 //x=86.095 //y=4.07 //x2=83.295 //y2=1.18
cc_5107 ( N_noxref_18_c_8064_n QN ) capacitor c=0.00642908f //x=86.095 \
 //y=4.07 //x2=86.95 //y2=2.22
cc_5108 ( N_noxref_18_c_8070_n QN ) capacitor c=0.0816497f //x=86.21 //y=2.08 \
 //x2=86.95 //y2=2.22
cc_5109 ( N_noxref_18_c_8309_p QN ) capacitor c=0.00998395f //x=86.23 \
 //y=4.705 //x2=86.95 //y2=2.22
cc_5110 ( N_noxref_18_c_8357_p QN ) capacitor c=0.0143966f //x=86.615 \
 //y=4.795 //x2=86.95 //y2=2.22
cc_5111 ( N_noxref_18_c_8293_p QN ) capacitor c=0.00704374f //x=86.21 //y=2.08 \
 //x2=86.95 //y2=2.22
cc_5112 ( N_noxref_18_c_8359_p QN ) capacitor c=0.0033061f //x=86.21 //y=1.915 \
 //x2=86.95 //y2=2.22
cc_5113 ( N_noxref_18_c_8299_p QN ) capacitor c=0.00526987f //x=86.23 \
 //y=4.705 //x2=86.95 //y2=2.22
cc_5114 ( N_noxref_18_c_8064_n N_QN_c_9164_n ) capacitor c=0.00154966f \
 //x=86.095 //y=4.07 //x2=86.385 //y2=5.21
cc_5115 ( N_noxref_18_c_8309_p N_QN_c_9164_n ) capacitor c=0.0128151f \
 //x=86.23 //y=4.705 //x2=86.385 //y2=5.21
cc_5116 ( N_noxref_18_M160_noxref_g N_QN_c_9164_n ) capacitor c=0.0167296f \
 //x=86.25 //y=6.025 //x2=86.385 //y2=5.21
cc_5117 ( N_noxref_18_c_8299_p N_QN_c_9164_n ) capacitor c=0.00368327f \
 //x=86.23 //y=4.705 //x2=86.385 //y2=5.21
cc_5118 ( N_noxref_18_c_8064_n N_QN_c_9126_n ) capacitor c=0.0138451f \
 //x=86.095 //y=4.07 //x2=85.675 //y2=5.21
cc_5119 ( N_noxref_18_M161_noxref_g N_QN_c_9127_n ) capacitor c=0.0222938f \
 //x=86.69 //y=6.025 //x2=86.865 //y2=5.21
cc_5120 ( N_noxref_18_c_8318_p N_QN_c_9113_n ) capacitor c=0.00810194f \
 //x=86.62 //y=1.405 //x2=86.865 //y2=1.645
cc_5121 ( N_noxref_18_c_8359_p N_QN_c_9171_n ) capacitor c=0.00671029f \
 //x=86.21 //y=1.915 //x2=86.595 //y2=1.645
cc_5122 ( N_noxref_18_c_8357_p N_QN_c_9172_n ) capacitor c=0.00410596f \
 //x=86.615 //y=4.795 //x2=86.47 //y2=5.21
cc_5123 ( N_noxref_18_c_8250_n N_QN_M49_noxref_d ) capacitor c=0.00218556f \
 //x=79.585 //y=0.905 //x2=79.66 //y2=0.905
cc_5124 ( N_noxref_18_c_8253_n N_QN_M49_noxref_d ) capacitor c=0.00327871f \
 //x=79.585 //y=1.25 //x2=79.66 //y2=0.905
cc_5125 ( N_noxref_18_c_8255_n N_QN_M49_noxref_d ) capacitor c=0.00292542f \
 //x=79.585 //y=1.56 //x2=79.66 //y2=0.905
cc_5126 ( N_noxref_18_c_8340_p N_QN_M49_noxref_d ) capacitor c=0.00235569f \
 //x=79.96 //y=0.75 //x2=79.66 //y2=0.905
cc_5127 ( N_noxref_18_c_8341_p N_QN_M49_noxref_d ) capacitor c=0.00613695f \
 //x=79.96 //y=1.405 //x2=79.66 //y2=0.905
cc_5128 ( N_noxref_18_c_8259_n N_QN_M49_noxref_d ) capacitor c=0.00131413f \
 //x=80.115 //y=0.905 //x2=79.66 //y2=0.905
cc_5129 ( N_noxref_18_c_8260_n N_QN_M49_noxref_d ) capacitor c=0.00676348f \
 //x=80.115 //y=1.25 //x2=79.66 //y2=0.905
cc_5130 ( N_noxref_18_c_8305_p N_QN_M53_noxref_d ) capacitor c=0.00226395f \
 //x=86.245 //y=0.905 //x2=86.32 //y2=0.905
cc_5131 ( N_noxref_18_c_8316_p N_QN_M53_noxref_d ) capacitor c=0.004517f \
 //x=86.245 //y=1.255 //x2=86.32 //y2=0.905
cc_5132 ( N_noxref_18_c_8307_p N_QN_M53_noxref_d ) capacitor c=0.00655125f \
 //x=86.245 //y=1.56 //x2=86.32 //y2=0.905
cc_5133 ( N_noxref_18_c_8348_p N_QN_M53_noxref_d ) capacitor c=0.00241003f \
 //x=86.62 //y=0.75 //x2=86.32 //y2=0.905
cc_5134 ( N_noxref_18_c_8318_p N_QN_M53_noxref_d ) capacitor c=0.0159024f \
 //x=86.62 //y=1.405 //x2=86.32 //y2=0.905
cc_5135 ( N_noxref_18_c_8315_p N_QN_M53_noxref_d ) capacitor c=0.00132831f \
 //x=86.775 //y=0.905 //x2=86.32 //y2=0.905
cc_5136 ( N_noxref_18_c_8319_p N_QN_M53_noxref_d ) capacitor c=0.00330743f \
 //x=86.775 //y=1.255 //x2=86.32 //y2=0.905
cc_5137 ( N_noxref_18_M160_noxref_g N_QN_M160_noxref_d ) capacitor \
 c=0.0130327f //x=86.25 //y=6.025 //x2=86.325 //y2=5.025
cc_5138 ( N_noxref_18_M161_noxref_g N_QN_M160_noxref_d ) capacitor \
 c=0.0136385f //x=86.69 //y=6.025 //x2=86.325 //y2=5.025
cc_5139 ( N_noxref_18_c_8065_n N_noxref_51_c_10700_n ) capacitor c=0.00207733f \
 //x=72.89 //y=2.08 //x2=73.545 //y2=0.54
cc_5140 ( N_noxref_18_c_8137_n N_noxref_51_c_10700_n ) capacitor c=0.0194423f \
 //x=72.88 //y=0.915 //x2=73.545 //y2=0.54
cc_5141 ( N_noxref_18_c_8199_n N_noxref_51_c_10700_n ) capacitor c=0.00656458f \
 //x=73.41 //y=0.915 //x2=73.545 //y2=0.54
cc_5142 ( N_noxref_18_c_8140_n N_noxref_51_c_10700_n ) capacitor c=2.20712e-19 \
 //x=72.89 //y=2.08 //x2=73.545 //y2=0.54
cc_5143 ( N_noxref_18_c_8138_n N_noxref_51_c_10722_n ) capacitor c=0.00538829f \
 //x=72.88 //y=1.26 //x2=72.66 //y2=0.995
cc_5144 ( N_noxref_18_c_8137_n N_noxref_51_M45_noxref_s ) capacitor \
 c=0.00538829f //x=72.88 //y=0.915 //x2=72.525 //y2=0.375
cc_5145 ( N_noxref_18_c_8139_n N_noxref_51_M45_noxref_s ) capacitor \
 c=0.00538829f //x=72.88 //y=1.57 //x2=72.525 //y2=0.375
cc_5146 ( N_noxref_18_c_8199_n N_noxref_51_M45_noxref_s ) capacitor \
 c=0.0143002f //x=73.41 //y=0.915 //x2=72.525 //y2=0.375
cc_5147 ( N_noxref_18_c_8200_n N_noxref_51_M45_noxref_s ) capacitor \
 c=0.00290153f //x=73.41 //y=1.26 //x2=72.525 //y2=0.375
cc_5148 ( N_noxref_18_c_8286_p N_noxref_52_c_10765_n ) capacitor c=3.15806e-19 \
 //x=76.605 //y=1.655 //x2=75.065 //y2=1.495
cc_5149 ( N_noxref_18_c_8286_p N_noxref_52_c_10754_n ) capacitor c=0.020324f \
 //x=76.605 //y=1.655 //x2=76.035 //y2=1.495
cc_5150 ( N_noxref_18_c_8066_n N_noxref_52_c_10755_n ) capacitor c=0.00464204f \
 //x=76.875 //y=1.655 //x2=76.92 //y2=0.53
cc_5151 ( N_noxref_18_M47_noxref_d N_noxref_52_c_10755_n ) capacitor \
 c=0.0117318f //x=76.33 //y=0.905 //x2=76.92 //y2=0.53
cc_5152 ( N_noxref_18_c_8066_n N_noxref_52_M46_noxref_s ) capacitor \
 c=0.0140283f //x=76.875 //y=1.655 //x2=74.93 //y2=0.365
cc_5153 ( N_noxref_18_M47_noxref_d N_noxref_52_M46_noxref_s ) capacitor \
 c=0.0439149f //x=76.33 //y=0.905 //x2=74.93 //y2=0.365
cc_5154 ( N_noxref_18_c_8066_n N_noxref_53_c_10816_n ) capacitor c=3.22188e-19 \
 //x=76.875 //y=1.655 //x2=78.395 //y2=1.495
cc_5155 ( N_noxref_18_c_8255_n N_noxref_53_c_10805_n ) capacitor c=0.00746306f \
 //x=79.585 //y=1.56 //x2=79.365 //y2=1.495
cc_5156 ( N_noxref_18_c_8072_n N_noxref_53_c_10805_n ) capacitor c=0.00174428f \
 //x=79.55 //y=2.08 //x2=79.365 //y2=1.495
cc_5157 ( N_noxref_18_c_8068_n N_noxref_53_c_10806_n ) capacitor c=0.00159234f \
 //x=79.55 //y=2.08 //x2=80.25 //y2=0.53
cc_5158 ( N_noxref_18_c_8250_n N_noxref_53_c_10806_n ) capacitor c=0.0200006f \
 //x=79.585 //y=0.905 //x2=80.25 //y2=0.53
cc_5159 ( N_noxref_18_c_8259_n N_noxref_53_c_10806_n ) capacitor c=0.00825432f \
 //x=80.115 //y=0.905 //x2=80.25 //y2=0.53
cc_5160 ( N_noxref_18_c_8072_n N_noxref_53_c_10806_n ) capacitor c=2.1838e-19 \
 //x=79.55 //y=2.08 //x2=80.25 //y2=0.53
cc_5161 ( N_noxref_18_c_8250_n N_noxref_53_M48_noxref_s ) capacitor \
 c=0.00746306f //x=79.585 //y=0.905 //x2=78.26 //y2=0.365
cc_5162 ( N_noxref_18_c_8255_n N_noxref_53_M48_noxref_s ) capacitor \
 c=0.00211573f //x=79.585 //y=1.56 //x2=78.26 //y2=0.365
cc_5163 ( N_noxref_18_c_8259_n N_noxref_53_M48_noxref_s ) capacitor \
 c=0.0133026f //x=80.115 //y=0.905 //x2=78.26 //y2=0.365
cc_5164 ( N_noxref_18_c_8260_n N_noxref_53_M48_noxref_s ) capacitor \
 c=0.00793126f //x=80.115 //y=1.25 //x2=78.26 //y2=0.365
cc_5165 ( N_noxref_18_c_8412_p N_noxref_53_M48_noxref_s ) capacitor \
 c=0.00392195f //x=79.55 //y=1.915 //x2=78.26 //y2=0.365
cc_5166 ( N_noxref_18_c_8064_n N_noxref_55_c_10910_n ) capacitor c=0.00631223f \
 //x=86.095 //y=4.07 //x2=85.94 //y2=1.58
cc_5167 ( N_noxref_18_c_8064_n N_noxref_55_c_10916_n ) capacitor c=0.00108825f \
 //x=86.095 //y=4.07 //x2=86.025 //y2=1.495
cc_5168 ( N_noxref_18_c_8307_p N_noxref_55_c_10916_n ) capacitor c=0.00698471f \
 //x=86.245 //y=1.56 //x2=86.025 //y2=1.495
cc_5169 ( N_noxref_18_c_8293_p N_noxref_55_c_10916_n ) capacitor c=0.00171785f \
 //x=86.21 //y=2.08 //x2=86.025 //y2=1.495
cc_5170 ( N_noxref_18_c_8070_n N_noxref_55_c_10917_n ) capacitor c=0.00118117f \
 //x=86.21 //y=2.08 //x2=86.91 //y2=0.53
cc_5171 ( N_noxref_18_c_8305_p N_noxref_55_c_10917_n ) capacitor c=0.0191024f \
 //x=86.245 //y=0.905 //x2=86.91 //y2=0.53
cc_5172 ( N_noxref_18_c_8315_p N_noxref_55_c_10917_n ) capacitor c=0.00655165f \
 //x=86.775 //y=0.905 //x2=86.91 //y2=0.53
cc_5173 ( N_noxref_18_c_8293_p N_noxref_55_c_10917_n ) capacitor c=2.1838e-19 \
 //x=86.21 //y=2.08 //x2=86.91 //y2=0.53
cc_5174 ( N_noxref_18_c_8305_p N_noxref_55_M52_noxref_s ) capacitor \
 c=0.00698471f //x=86.245 //y=0.905 //x2=84.92 //y2=0.365
cc_5175 ( N_noxref_18_c_8318_p N_noxref_55_M52_noxref_s ) capacitor \
 c=0.00316186f //x=86.62 //y=1.405 //x2=84.92 //y2=0.365
cc_5176 ( N_noxref_18_c_8315_p N_noxref_55_M52_noxref_s ) capacitor \
 c=0.0142835f //x=86.775 //y=0.905 //x2=84.92 //y2=0.365
cc_5177 ( N_noxref_19_M157_noxref_d N_noxref_20_c_8541_n ) capacitor \
 c=0.00496677f //x=83.425 //y=5.025 //x2=83.62 //y2=2.08
cc_5178 ( N_noxref_19_c_8489_p N_noxref_20_M156_noxref_g ) capacitor \
 c=0.0150104f //x=83.485 //y=6.91 //x2=82.91 //y2=6.025
cc_5179 ( N_noxref_19_M155_noxref_d N_noxref_20_M156_noxref_g ) capacitor \
 c=0.0130327f //x=82.545 //y=5.025 //x2=82.91 //y2=6.025
cc_5180 ( N_noxref_19_c_8489_p N_noxref_20_M157_noxref_g ) capacitor \
 c=0.0155183f //x=83.485 //y=6.91 //x2=83.35 //y2=6.025
cc_5181 ( N_noxref_19_M157_noxref_d N_noxref_20_M157_noxref_g ) capacitor \
 c=0.0398886f //x=83.425 //y=5.025 //x2=83.35 //y2=6.025
cc_5182 ( N_noxref_19_M157_noxref_d N_noxref_20_c_8584_n ) capacitor \
 c=0.00411435f //x=83.425 //y=5.025 //x2=83.35 //y2=4.87
cc_5183 ( N_noxref_19_c_8489_p N_noxref_21_c_9008_n ) capacitor c=0.00546043f \
 //x=83.485 //y=6.91 //x2=85.035 //y2=5.21
cc_5184 ( N_noxref_19_M157_noxref_d N_noxref_21_c_9008_n ) capacitor \
 c=0.00675852f //x=83.425 //y=5.025 //x2=85.035 //y2=5.21
cc_5185 ( N_noxref_19_c_8424_n N_noxref_21_c_9012_n ) capacitor c=0.0086908f \
 //x=81.695 //y=5.21 //x2=83.245 //y2=5.21
cc_5186 ( N_noxref_19_c_8489_p N_noxref_21_c_9012_n ) capacitor c=9.39989e-19 \
 //x=83.485 //y=6.91 //x2=83.245 //y2=5.21
cc_5187 ( N_noxref_19_c_8470_n N_noxref_21_c_9023_n ) capacitor c=0.00102709f \
 //x=82.605 //y=6.91 //x2=83.045 //y2=5.21
cc_5188 ( N_noxref_19_c_8489_p N_noxref_21_c_9023_n ) capacitor c=9.89472e-19 \
 //x=83.485 //y=6.91 //x2=83.045 //y2=5.21
cc_5189 ( N_noxref_19_M155_noxref_d N_noxref_21_c_9023_n ) capacitor \
 c=0.0124612f //x=82.545 //y=5.025 //x2=83.045 //y2=5.21
cc_5190 ( N_noxref_19_c_8424_n N_noxref_21_c_9014_n ) capacitor c=0.00638395f \
 //x=81.695 //y=5.21 //x2=82.335 //y2=5.21
cc_5191 ( N_noxref_19_c_8444_n N_noxref_21_c_9014_n ) capacitor c=0.0682565f \
 //x=81.81 //y=5.21 //x2=82.335 //y2=5.21
cc_5192 ( N_noxref_19_c_8444_n N_noxref_21_c_9015_n ) capacitor c=9.46973e-19 \
 //x=81.81 //y=5.21 //x2=83.13 //y2=5.295
cc_5193 ( N_noxref_19_M157_noxref_d N_noxref_21_c_9016_n ) capacitor \
 c=0.001104f //x=83.425 //y=5.025 //x2=85.15 //y2=5.21
cc_5194 ( N_noxref_19_c_8489_p N_noxref_21_c_9018_n ) capacitor c=0.001104f \
 //x=83.485 //y=6.91 //x2=85.235 //y2=6.91
cc_5195 ( N_noxref_19_c_8424_n N_noxref_21_M154_noxref_d ) capacitor \
 c=4.76678e-19 //x=81.695 //y=5.21 //x2=82.105 //y2=5.025
cc_5196 ( N_noxref_19_c_8470_n N_noxref_21_M154_noxref_d ) capacitor \
 c=0.0115421f //x=82.605 //y=6.91 //x2=82.105 //y2=5.025
cc_5197 ( N_noxref_19_M155_noxref_d N_noxref_21_M154_noxref_d ) capacitor \
 c=0.0458293f //x=82.545 //y=5.025 //x2=82.105 //y2=5.025
cc_5198 ( N_noxref_19_M157_noxref_d N_noxref_21_M154_noxref_d ) capacitor \
 c=7.47391e-19 //x=83.425 //y=5.025 //x2=82.105 //y2=5.025
cc_5199 ( N_noxref_19_c_8444_n N_noxref_21_M156_noxref_d ) capacitor \
 c=9.55e-19 //x=81.81 //y=5.21 //x2=82.985 //y2=5.025
cc_5200 ( N_noxref_19_c_8489_p N_noxref_21_M156_noxref_d ) capacitor \
 c=0.0115693f //x=83.485 //y=6.91 //x2=82.985 //y2=5.025
cc_5201 ( N_noxref_19_M155_noxref_d N_noxref_21_M156_noxref_d ) capacitor \
 c=0.0458293f //x=82.545 //y=5.025 //x2=82.985 //y2=5.025
cc_5202 ( N_noxref_19_M157_noxref_d N_noxref_21_M156_noxref_d ) capacitor \
 c=0.0550393f //x=83.425 //y=5.025 //x2=82.985 //y2=5.025
cc_5203 ( N_noxref_19_c_8444_n N_noxref_54_c_10872_n ) capacitor c=0.00109479f \
 //x=81.81 //y=5.21 //x2=81.725 //y2=1.495
cc_5204 ( N_noxref_20_c_8516_n N_noxref_21_c_9008_n ) capacitor c=7.38711e-19 \
 //x=83.505 //y=2.96 //x2=85.035 //y2=5.21
cc_5205 ( N_noxref_20_c_8536_n N_noxref_21_c_9008_n ) capacitor c=5.48246e-19 \
 //x=84.985 //y=2.08 //x2=85.035 //y2=5.21
cc_5206 ( N_noxref_20_c_8541_n N_noxref_21_c_9008_n ) capacitor c=0.00419026f \
 //x=83.62 //y=2.08 //x2=85.035 //y2=5.21
cc_5207 ( N_noxref_20_c_8543_n N_noxref_21_c_9008_n ) capacitor c=0.0031527f \
 //x=85.1 //y=2.08 //x2=85.035 //y2=5.21
cc_5208 ( N_noxref_20_M157_noxref_g N_noxref_21_c_9008_n ) capacitor \
 c=0.0109874f //x=83.35 //y=6.025 //x2=85.035 //y2=5.21
cc_5209 ( N_noxref_20_M158_noxref_g N_noxref_21_c_9008_n ) capacitor \
 c=0.00645933f //x=85.37 //y=6.025 //x2=85.035 //y2=5.21
cc_5210 ( N_noxref_20_c_8584_n N_noxref_21_c_9008_n ) capacitor c=0.00270424f \
 //x=83.35 //y=4.87 //x2=85.035 //y2=5.21
cc_5211 ( N_noxref_20_c_8585_n N_noxref_21_c_9008_n ) capacitor c=0.00176728f \
 //x=85.445 //y=4.795 //x2=85.035 //y2=5.21
cc_5212 ( N_noxref_20_c_8516_n N_noxref_21_c_9012_n ) capacitor c=3.75024e-19 \
 //x=83.505 //y=2.96 //x2=83.245 //y2=5.21
cc_5213 ( N_noxref_20_M156_noxref_g N_noxref_21_c_9012_n ) capacitor \
 c=6.87102e-19 //x=82.91 //y=6.025 //x2=83.245 //y2=5.21
cc_5214 ( N_noxref_20_M157_noxref_g N_noxref_21_c_9012_n ) capacitor \
 c=8.33934e-19 //x=83.35 //y=6.025 //x2=83.245 //y2=5.21
cc_5215 ( N_noxref_20_M156_noxref_g N_noxref_21_c_9023_n ) capacitor \
 c=0.0179287f //x=82.91 //y=6.025 //x2=83.045 //y2=5.21
cc_5216 ( N_noxref_20_M156_noxref_g N_noxref_21_c_9015_n ) capacitor \
 c=0.0019882f //x=82.91 //y=6.025 //x2=83.13 //y2=5.295
cc_5217 ( N_noxref_20_M157_noxref_g N_noxref_21_c_9015_n ) capacitor \
 c=0.0159381f //x=83.35 //y=6.025 //x2=83.13 //y2=5.295
cc_5218 ( N_noxref_20_c_8901_p N_noxref_21_c_9015_n ) capacitor c=0.00456817f \
 //x=83.275 //y=4.795 //x2=83.13 //y2=5.295
cc_5219 ( N_noxref_20_c_8543_n N_noxref_21_c_9016_n ) capacitor c=0.0183146f \
 //x=85.1 //y=2.08 //x2=85.15 //y2=5.21
cc_5220 ( N_noxref_20_M158_noxref_g N_noxref_21_c_9016_n ) capacitor \
 c=0.0484795f //x=85.37 //y=6.025 //x2=85.15 //y2=5.21
cc_5221 ( N_noxref_20_c_8585_n N_noxref_21_c_9016_n ) capacitor c=0.0078825f \
 //x=85.445 //y=4.795 //x2=85.15 //y2=5.21
cc_5222 ( N_noxref_20_M158_noxref_g N_noxref_21_c_9035_n ) capacitor \
 c=0.0164606f //x=85.37 //y=6.025 //x2=85.945 //y2=6.91
cc_5223 ( N_noxref_20_M159_noxref_g N_noxref_21_c_9035_n ) capacitor \
 c=0.0150104f //x=85.81 //y=6.025 //x2=85.945 //y2=6.91
cc_5224 ( N_noxref_20_M156_noxref_g N_noxref_21_M156_noxref_d ) capacitor \
 c=0.0129738f //x=82.91 //y=6.025 //x2=82.985 //y2=5.025
cc_5225 ( N_noxref_20_M159_noxref_g N_noxref_21_M159_noxref_d ) capacitor \
 c=0.0130327f //x=85.81 //y=6.025 //x2=85.885 //y2=5.025
cc_5226 ( N_noxref_20_c_8516_n N_QN_c_9097_n ) capacitor c=0.0489549f \
 //x=83.505 //y=2.96 //x2=83.065 //y2=1.18
cc_5227 ( N_noxref_20_c_8825_n N_QN_c_9097_n ) capacitor c=5.17481e-19 \
 //x=82.915 //y=0.905 //x2=83.065 //y2=1.18
cc_5228 ( N_noxref_20_c_8828_n N_QN_c_9097_n ) capacitor c=0.00609699f \
 //x=82.915 //y=1.25 //x2=83.065 //y2=1.18
cc_5229 ( N_noxref_20_c_8516_n N_QN_c_9104_n ) capacitor c=0.00467724f \
 //x=83.505 //y=2.96 //x2=79.965 //y2=1.18
cc_5230 ( N_noxref_20_c_8516_n N_QN_c_9105_n ) capacitor c=0.00337366f \
 //x=83.505 //y=2.96 //x2=86.395 //y2=1.18
cc_5231 ( N_noxref_20_c_8536_n N_QN_c_9105_n ) capacitor c=0.053129f \
 //x=84.985 //y=2.08 //x2=86.395 //y2=1.18
cc_5232 ( N_noxref_20_c_8537_n N_QN_c_9105_n ) capacitor c=0.0102038f \
 //x=83.735 //y=2.08 //x2=86.395 //y2=1.18
cc_5233 ( N_noxref_20_c_8541_n N_QN_c_9105_n ) capacitor c=0.00189559f \
 //x=83.62 //y=2.08 //x2=86.395 //y2=1.18
cc_5234 ( N_noxref_20_c_8543_n N_QN_c_9105_n ) capacitor c=0.00134607f \
 //x=85.1 //y=2.08 //x2=86.395 //y2=1.18
cc_5235 ( N_noxref_20_c_8834_n N_QN_c_9105_n ) capacitor c=4.67724e-19 \
 //x=83.445 //y=0.905 //x2=86.395 //y2=1.18
cc_5236 ( N_noxref_20_c_8835_n N_QN_c_9105_n ) capacitor c=0.00591245f \
 //x=83.445 //y=1.25 //x2=86.395 //y2=1.18
cc_5237 ( N_noxref_20_c_8836_n N_QN_c_9105_n ) capacitor c=0.00326119f \
 //x=83.445 //y=1.56 //x2=86.395 //y2=1.18
cc_5238 ( N_noxref_20_c_8544_n N_QN_c_9105_n ) capacitor c=2.04565e-19 \
 //x=83.445 //y=1.915 //x2=86.395 //y2=1.18
cc_5239 ( N_noxref_20_c_8547_n N_QN_c_9105_n ) capacitor c=0.00500281f \
 //x=85.275 //y=1.21 //x2=86.395 //y2=1.18
cc_5240 ( N_noxref_20_c_8866_n N_QN_c_9105_n ) capacitor c=0.00361177f \
 //x=85.275 //y=1.52 //x2=86.395 //y2=1.18
cc_5241 ( N_noxref_20_c_8549_n N_QN_c_9105_n ) capacitor c=4.02408e-19 \
 //x=85.65 //y=0.71 //x2=86.395 //y2=1.18
cc_5242 ( N_noxref_20_c_8550_n N_QN_c_9105_n ) capacitor c=0.0036677f \
 //x=85.65 //y=1.365 //x2=86.395 //y2=1.18
cc_5243 ( N_noxref_20_c_8553_n N_QN_c_9105_n ) capacitor c=0.00776505f \
 //x=85.805 //y=1.21 //x2=86.395 //y2=1.18
cc_5244 ( N_noxref_20_c_8516_n N_QN_c_9111_n ) capacitor c=0.00413336f \
 //x=83.505 //y=2.96 //x2=83.295 //y2=1.18
cc_5245 ( N_noxref_20_c_8828_n N_QN_c_9111_n ) capacitor c=0.0015439f \
 //x=82.915 //y=1.25 //x2=83.295 //y2=1.18
cc_5246 ( N_noxref_20_c_8929_p N_QN_c_9111_n ) capacitor c=4.52813e-19 \
 //x=83.29 //y=0.75 //x2=83.295 //y2=1.18
cc_5247 ( N_noxref_20_c_8930_p N_QN_c_9111_n ) capacitor c=7.42023e-19 \
 //x=83.29 //y=1.405 //x2=83.295 //y2=1.18
cc_5248 ( N_noxref_20_c_8835_n N_QN_c_9111_n ) capacitor c=4.79299e-19 \
 //x=83.445 //y=1.25 //x2=83.295 //y2=1.18
cc_5249 ( N_noxref_20_c_8836_n N_QN_c_9111_n ) capacitor c=9.64184e-19 \
 //x=83.445 //y=1.56 //x2=83.295 //y2=1.18
cc_5250 ( N_noxref_20_c_8543_n QN ) capacitor c=0.00370801f //x=85.1 //y=2.08 \
 //x2=86.95 //y2=2.22
cc_5251 ( N_noxref_20_M159_noxref_g N_QN_c_9164_n ) capacitor c=0.0179287f \
 //x=85.81 //y=6.025 //x2=86.385 //y2=5.21
cc_5252 ( N_noxref_20_M158_noxref_g N_QN_c_9126_n ) capacitor c=0.0132916f \
 //x=85.37 //y=6.025 //x2=85.675 //y2=5.21
cc_5253 ( N_noxref_20_c_8868_n N_QN_c_9126_n ) capacitor c=0.00405122f \
 //x=85.735 //y=4.795 //x2=85.675 //y2=5.21
cc_5254 ( N_noxref_20_c_8516_n N_QN_M49_noxref_d ) capacitor c=0.00446326f \
 //x=83.505 //y=2.96 //x2=79.66 //y2=0.905
cc_5255 ( N_noxref_20_c_8516_n N_QN_M51_noxref_d ) capacitor c=0.00446423f \
 //x=83.505 //y=2.96 //x2=82.99 //y2=0.905
cc_5256 ( N_noxref_20_c_8825_n N_QN_M51_noxref_d ) capacitor c=0.00217566f \
 //x=82.915 //y=0.905 //x2=82.99 //y2=0.905
cc_5257 ( N_noxref_20_c_8828_n N_QN_M51_noxref_d ) capacitor c=0.00711747f \
 //x=82.915 //y=1.25 //x2=82.99 //y2=0.905
cc_5258 ( N_noxref_20_c_8929_p N_QN_M51_noxref_d ) capacitor c=0.00234223f \
 //x=83.29 //y=0.75 //x2=82.99 //y2=0.905
cc_5259 ( N_noxref_20_c_8930_p N_QN_M51_noxref_d ) capacitor c=0.00602848f \
 //x=83.29 //y=1.405 //x2=82.99 //y2=0.905
cc_5260 ( N_noxref_20_c_8834_n N_QN_M51_noxref_d ) capacitor c=0.00132245f \
 //x=83.445 //y=0.905 //x2=82.99 //y2=0.905
cc_5261 ( N_noxref_20_c_8835_n N_QN_M51_noxref_d ) capacitor c=0.004434f \
 //x=83.445 //y=1.25 //x2=82.99 //y2=0.905
cc_5262 ( N_noxref_20_c_8836_n N_QN_M51_noxref_d ) capacitor c=0.00270197f \
 //x=83.445 //y=1.56 //x2=82.99 //y2=0.905
cc_5263 ( N_noxref_20_M159_noxref_g N_QN_M158_noxref_d ) capacitor \
 c=0.0130327f //x=85.81 //y=6.025 //x2=85.445 //y2=5.025
cc_5264 ( N_noxref_20_c_8538_n N_noxref_31_c_9679_n ) capacitor c=0.00204385f \
 //x=21.09 //y=2.08 //x2=21.745 //y2=0.54
cc_5265 ( N_noxref_20_c_8638_n N_noxref_31_c_9679_n ) capacitor c=0.0194423f \
 //x=21.08 //y=0.915 //x2=21.745 //y2=0.54
cc_5266 ( N_noxref_20_c_8644_n N_noxref_31_c_9679_n ) capacitor c=0.00656458f \
 //x=21.61 //y=0.915 //x2=21.745 //y2=0.54
cc_5267 ( N_noxref_20_c_8647_n N_noxref_31_c_9679_n ) capacitor c=2.20712e-19 \
 //x=21.09 //y=2.08 //x2=21.745 //y2=0.54
cc_5268 ( N_noxref_20_c_8639_n N_noxref_31_c_9689_n ) capacitor c=0.00538829f \
 //x=21.08 //y=1.26 //x2=20.86 //y2=0.995
cc_5269 ( N_noxref_20_c_8638_n N_noxref_31_M13_noxref_s ) capacitor \
 c=0.00538829f //x=21.08 //y=0.915 //x2=20.725 //y2=0.375
cc_5270 ( N_noxref_20_c_8640_n N_noxref_31_M13_noxref_s ) capacitor \
 c=0.00538829f //x=21.08 //y=1.57 //x2=20.725 //y2=0.375
cc_5271 ( N_noxref_20_c_8644_n N_noxref_31_M13_noxref_s ) capacitor \
 c=0.0143002f //x=21.61 //y=0.915 //x2=20.725 //y2=0.375
cc_5272 ( N_noxref_20_c_8645_n N_noxref_31_M13_noxref_s ) capacitor \
 c=0.00290153f //x=21.61 //y=1.26 //x2=20.725 //y2=0.375
cc_5273 ( N_noxref_20_c_8761_n N_noxref_32_c_9744_n ) capacitor c=3.15806e-19 \
 //x=24.805 //y=1.655 //x2=23.265 //y2=1.495
cc_5274 ( N_noxref_20_c_8761_n N_noxref_32_c_9733_n ) capacitor c=0.020324f \
 //x=24.805 //y=1.655 //x2=24.235 //y2=1.495
cc_5275 ( N_noxref_20_c_8539_n N_noxref_32_c_9734_n ) capacitor c=0.00457164f \
 //x=25.075 //y=1.655 //x2=25.12 //y2=0.53
cc_5276 ( N_noxref_20_M15_noxref_d N_noxref_32_c_9734_n ) capacitor \
 c=0.0115831f //x=24.53 //y=0.905 //x2=25.12 //y2=0.53
cc_5277 ( N_noxref_20_c_8539_n N_noxref_32_M14_noxref_s ) capacitor \
 c=0.013435f //x=25.075 //y=1.655 //x2=23.13 //y2=0.365
cc_5278 ( N_noxref_20_M15_noxref_d N_noxref_32_M14_noxref_s ) capacitor \
 c=0.0439476f //x=24.53 //y=0.905 //x2=23.13 //y2=0.365
cc_5279 ( N_noxref_20_c_8539_n N_noxref_33_c_9793_n ) capacitor c=4.08644e-19 \
 //x=25.075 //y=1.655 //x2=26.49 //y2=1.505
cc_5280 ( N_noxref_20_M15_noxref_d N_noxref_33_M16_noxref_s ) capacitor \
 c=2.53688e-19 //x=24.53 //y=0.905 //x2=26.355 //y2=0.375
cc_5281 ( N_noxref_20_c_8516_n N_noxref_50_c_10673_n ) capacitor c=0.00152987f \
 //x=83.505 //y=2.96 //x2=72.005 //y2=1.59
cc_5282 ( N_noxref_20_c_8516_n N_noxref_50_M43_noxref_s ) capacitor \
 c=0.00302917f //x=83.505 //y=2.96 //x2=70.015 //y2=0.375
cc_5283 ( N_noxref_20_c_8516_n N_noxref_51_c_10695_n ) capacitor c=0.00383675f \
 //x=83.505 //y=2.96 //x2=72.575 //y2=0.995
cc_5284 ( N_noxref_20_c_8516_n N_noxref_51_c_10700_n ) capacitor c=6.69632e-19 \
 //x=83.505 //y=2.96 //x2=73.545 //y2=0.54
cc_5285 ( N_noxref_20_c_8516_n N_noxref_51_M45_noxref_s ) capacitor \
 c=0.00324882f //x=83.505 //y=2.96 //x2=72.525 //y2=0.375
cc_5286 ( N_noxref_20_c_8516_n N_noxref_52_c_10765_n ) capacitor c=0.00321948f \
 //x=83.505 //y=2.96 //x2=75.065 //y2=1.495
cc_5287 ( N_noxref_20_c_8516_n N_noxref_52_c_10747_n ) capacitor c=0.0126836f \
 //x=83.505 //y=2.96 //x2=75.95 //y2=1.58
cc_5288 ( N_noxref_20_c_8516_n N_noxref_52_c_10754_n ) capacitor c=0.00321948f \
 //x=83.505 //y=2.96 //x2=76.035 //y2=1.495
cc_5289 ( N_noxref_20_c_8516_n N_noxref_52_c_10755_n ) capacitor c=9.10579e-19 \
 //x=83.505 //y=2.96 //x2=76.92 //y2=0.53
cc_5290 ( N_noxref_20_c_8516_n N_noxref_52_M46_noxref_s ) capacitor \
 c=6.20367e-19 //x=83.505 //y=2.96 //x2=74.93 //y2=0.365
cc_5291 ( N_noxref_20_c_8516_n N_noxref_53_c_10816_n ) capacitor c=8.52215e-19 \
 //x=83.505 //y=2.96 //x2=78.395 //y2=1.495
cc_5292 ( N_noxref_20_c_8516_n N_noxref_53_c_10798_n ) capacitor c=0.0139765f \
 //x=83.505 //y=2.96 //x2=79.28 //y2=1.58
cc_5293 ( N_noxref_20_c_8516_n N_noxref_53_c_10805_n ) capacitor c=0.00321948f \
 //x=83.505 //y=2.96 //x2=79.365 //y2=1.495
cc_5294 ( N_noxref_20_c_8516_n N_noxref_53_c_10806_n ) capacitor c=4.76383e-19 \
 //x=83.505 //y=2.96 //x2=80.25 //y2=0.53
cc_5295 ( N_noxref_20_c_8516_n N_noxref_53_M48_noxref_s ) capacitor \
 c=0.00285734f //x=83.505 //y=2.96 //x2=78.26 //y2=0.365
cc_5296 ( N_noxref_20_c_8516_n N_noxref_54_c_10872_n ) capacitor c=0.00256304f \
 //x=83.505 //y=2.96 //x2=81.725 //y2=1.495
cc_5297 ( N_noxref_20_c_8516_n N_noxref_54_c_10855_n ) capacitor c=0.0114954f \
 //x=83.505 //y=2.96 //x2=82.61 //y2=1.58
cc_5298 ( N_noxref_20_c_8516_n N_noxref_54_c_10861_n ) capacitor c=0.00285734f \
 //x=83.505 //y=2.96 //x2=82.695 //y2=1.495
cc_5299 ( N_noxref_20_c_8544_n N_noxref_54_c_10861_n ) capacitor c=0.0028747f \
 //x=83.445 //y=1.915 //x2=82.695 //y2=1.495
cc_5300 ( N_noxref_20_c_8825_n N_noxref_54_c_10862_n ) capacitor c=0.021566f \
 //x=82.915 //y=0.905 //x2=83.58 //y2=0.53
cc_5301 ( N_noxref_20_c_8834_n N_noxref_54_c_10862_n ) capacitor c=0.00781103f \
 //x=83.445 //y=0.905 //x2=83.58 //y2=0.53
cc_5302 ( N_noxref_20_c_8536_n N_noxref_54_M50_noxref_s ) capacitor \
 c=5.34178e-19 //x=84.985 //y=2.08 //x2=81.59 //y2=0.365
cc_5303 ( N_noxref_20_c_8537_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.00116116f //x=83.735 //y=2.08 //x2=81.59 //y2=0.365
cc_5304 ( N_noxref_20_c_8541_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.016698f //x=83.62 //y=2.08 //x2=81.59 //y2=0.365
cc_5305 ( N_noxref_20_c_8825_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.0064603f //x=82.915 //y=0.905 //x2=81.59 //y2=0.365
cc_5306 ( N_noxref_20_c_8828_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.00602248f //x=82.915 //y=1.25 //x2=81.59 //y2=0.365
cc_5307 ( N_noxref_20_c_8834_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.0321601f //x=83.445 //y=0.905 //x2=81.59 //y2=0.365
cc_5308 ( N_noxref_20_c_8836_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.00239072f //x=83.445 //y=1.56 //x2=81.59 //y2=0.365
cc_5309 ( N_noxref_20_c_8544_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.00784558f //x=83.445 //y=1.915 //x2=81.59 //y2=0.365
cc_5310 ( N_noxref_20_c_8536_n N_noxref_55_c_10937_n ) capacitor c=0.00169534f \
 //x=84.985 //y=2.08 //x2=85.055 //y2=1.495
cc_5311 ( N_noxref_20_c_8543_n N_noxref_55_c_10937_n ) capacitor c=0.016698f \
 //x=85.1 //y=2.08 //x2=85.055 //y2=1.495
cc_5312 ( N_noxref_20_c_8548_n N_noxref_55_c_10937_n ) capacitor c=0.0034165f \
 //x=85.275 //y=1.915 //x2=85.055 //y2=1.495
cc_5313 ( N_noxref_20_c_8554_n N_noxref_55_c_10937_n ) capacitor c=0.00531095f \
 //x=85.1 //y=2.08 //x2=85.055 //y2=1.495
cc_5314 ( N_noxref_20_c_8536_n N_noxref_55_c_10910_n ) capacitor c=0.00222439f \
 //x=84.985 //y=2.08 //x2=85.94 //y2=1.58
cc_5315 ( N_noxref_20_c_8543_n N_noxref_55_c_10910_n ) capacitor c=0.00587616f \
 //x=85.1 //y=2.08 //x2=85.94 //y2=1.58
cc_5316 ( N_noxref_20_c_8866_n N_noxref_55_c_10910_n ) capacitor c=0.0061593f \
 //x=85.275 //y=1.52 //x2=85.94 //y2=1.58
cc_5317 ( N_noxref_20_c_8548_n N_noxref_55_c_10910_n ) capacitor c=0.0142098f \
 //x=85.275 //y=1.915 //x2=85.94 //y2=1.58
cc_5318 ( N_noxref_20_c_8550_n N_noxref_55_c_10910_n ) capacitor c=0.00991953f \
 //x=85.65 //y=1.365 //x2=85.94 //y2=1.58
cc_5319 ( N_noxref_20_c_8553_n N_noxref_55_c_10910_n ) capacitor c=0.00339872f \
 //x=85.805 //y=1.21 //x2=85.94 //y2=1.58
cc_5320 ( N_noxref_20_c_8554_n N_noxref_55_c_10910_n ) capacitor c=0.00147967f \
 //x=85.1 //y=2.08 //x2=85.94 //y2=1.58
cc_5321 ( N_noxref_20_c_8548_n N_noxref_55_c_10916_n ) capacitor c=6.71402e-19 \
 //x=85.275 //y=1.915 //x2=86.025 //y2=1.495
cc_5322 ( N_noxref_20_c_8545_n N_noxref_55_M52_noxref_s ) capacitor \
 c=0.0314164f //x=85.275 //y=0.865 //x2=84.92 //y2=0.365
cc_5323 ( N_noxref_20_c_8866_n N_noxref_55_M52_noxref_s ) capacitor \
 c=0.00110192f //x=85.275 //y=1.52 //x2=84.92 //y2=0.365
cc_5324 ( N_noxref_20_c_8551_n N_noxref_55_M52_noxref_s ) capacitor \
 c=0.0132463f //x=85.805 //y=0.865 //x2=84.92 //y2=0.365
cc_5325 ( N_noxref_21_c_9016_n QN ) capacitor c=3.02032e-19 //x=85.15 //y=5.21 \
 //x2=86.95 //y2=2.22
cc_5326 ( N_noxref_21_c_9035_n N_QN_c_9164_n ) capacitor c=0.00102709f \
 //x=85.945 //y=6.91 //x2=86.385 //y2=5.21
cc_5327 ( N_noxref_21_c_9036_n N_QN_c_9164_n ) capacitor c=0.00101874f \
 //x=86.825 //y=6.91 //x2=86.385 //y2=5.21
cc_5328 ( N_noxref_21_M159_noxref_d N_QN_c_9164_n ) capacitor c=0.012404f \
 //x=85.885 //y=5.025 //x2=86.385 //y2=5.21
cc_5329 ( N_noxref_21_c_9008_n N_QN_c_9126_n ) capacitor c=0.00602307f \
 //x=85.035 //y=5.21 //x2=85.675 //y2=5.21
cc_5330 ( N_noxref_21_c_9016_n N_QN_c_9126_n ) capacitor c=0.0683084f \
 //x=85.15 //y=5.21 //x2=85.675 //y2=5.21
cc_5331 ( N_noxref_21_c_9036_n N_QN_c_9127_n ) capacitor c=0.00173777f \
 //x=86.825 //y=6.91 //x2=86.865 //y2=5.21
cc_5332 ( N_noxref_21_M161_noxref_d N_QN_c_9127_n ) capacitor c=0.0159033f \
 //x=86.765 //y=5.025 //x2=86.865 //y2=5.21
cc_5333 ( N_noxref_21_c_9008_n N_QN_M158_noxref_d ) capacitor c=8.04912e-19 \
 //x=85.035 //y=5.21 //x2=85.445 //y2=5.025
cc_5334 ( N_noxref_21_c_9035_n N_QN_M158_noxref_d ) capacitor c=0.0117542f \
 //x=85.945 //y=6.91 //x2=85.445 //y2=5.025
cc_5335 ( N_noxref_21_M159_noxref_d N_QN_M158_noxref_d ) capacitor \
 c=0.0458293f //x=85.885 //y=5.025 //x2=85.445 //y2=5.025
cc_5336 ( N_noxref_21_c_9016_n N_QN_M160_noxref_d ) capacitor c=9.91979e-19 \
 //x=85.15 //y=5.21 //x2=86.325 //y2=5.025
cc_5337 ( N_noxref_21_c_9036_n N_QN_M160_noxref_d ) capacitor c=0.0118172f \
 //x=86.825 //y=6.91 //x2=86.325 //y2=5.025
cc_5338 ( N_noxref_21_M159_noxref_d N_QN_M160_noxref_d ) capacitor \
 c=0.0458293f //x=85.885 //y=5.025 //x2=86.325 //y2=5.025
cc_5339 ( N_noxref_21_M161_noxref_d N_QN_M160_noxref_d ) capacitor \
 c=0.0458293f //x=86.765 //y=5.025 //x2=86.325 //y2=5.025
cc_5340 ( N_QN_c_9097_n N_noxref_53_c_10806_n ) capacitor c=0.00641749f \
 //x=83.065 //y=1.18 //x2=80.25 //y2=0.53
cc_5341 ( N_QN_c_9104_n N_noxref_53_c_10806_n ) capacitor c=0.00219859f \
 //x=79.965 //y=1.18 //x2=80.25 //y2=0.53
cc_5342 ( N_QN_M49_noxref_d N_noxref_53_c_10806_n ) capacitor c=0.0136817f \
 //x=79.66 //y=0.905 //x2=80.25 //y2=0.53
cc_5343 ( N_QN_c_9097_n N_noxref_53_M48_noxref_s ) capacitor c=0.0207977f \
 //x=83.065 //y=1.18 //x2=78.26 //y2=0.365
cc_5344 ( N_QN_c_9104_n N_noxref_53_M48_noxref_s ) capacitor c=0.00804471f \
 //x=79.965 //y=1.18 //x2=78.26 //y2=0.365
cc_5345 ( N_QN_M49_noxref_d N_noxref_53_M48_noxref_s ) capacitor c=0.0458734f \
 //x=79.66 //y=0.905 //x2=78.26 //y2=0.365
cc_5346 ( N_QN_c_9097_n N_noxref_54_c_10855_n ) capacitor c=0.0224452f \
 //x=83.065 //y=1.18 //x2=82.61 //y2=1.58
cc_5347 ( N_QN_c_9097_n N_noxref_54_c_10862_n ) capacitor c=0.00641749f \
 //x=83.065 //y=1.18 //x2=83.58 //y2=0.53
cc_5348 ( N_QN_c_9105_n N_noxref_54_c_10862_n ) capacitor c=0.00641749f \
 //x=86.395 //y=1.18 //x2=83.58 //y2=0.53
cc_5349 ( N_QN_c_9111_n N_noxref_54_c_10862_n ) capacitor c=0.0015838f \
 //x=83.295 //y=1.18 //x2=83.58 //y2=0.53
cc_5350 ( N_QN_M51_noxref_d N_noxref_54_c_10862_n ) capacitor c=0.0130616f \
 //x=82.99 //y=0.905 //x2=83.58 //y2=0.53
cc_5351 ( N_QN_c_9097_n N_noxref_54_M50_noxref_s ) capacitor c=0.0443893f \
 //x=83.065 //y=1.18 //x2=81.59 //y2=0.365
cc_5352 ( N_QN_c_9105_n N_noxref_54_M50_noxref_s ) capacitor c=0.019112f \
 //x=86.395 //y=1.18 //x2=81.59 //y2=0.365
cc_5353 ( N_QN_c_9111_n N_noxref_54_M50_noxref_s ) capacitor c=0.00279707f \
 //x=83.295 //y=1.18 //x2=81.59 //y2=0.365
cc_5354 ( N_QN_M51_noxref_d N_noxref_54_M50_noxref_s ) capacitor c=0.0444718f \
 //x=82.99 //y=0.905 //x2=81.59 //y2=0.365
cc_5355 ( N_QN_c_9171_n N_noxref_55_c_10937_n ) capacitor c=2.73698e-19 \
 //x=86.595 //y=1.645 //x2=85.055 //y2=1.495
cc_5356 ( N_QN_c_9105_n N_noxref_55_c_10910_n ) capacitor c=0.0234642f \
 //x=86.395 //y=1.18 //x2=85.94 //y2=1.58
cc_5357 ( N_QN_c_9171_n N_noxref_55_c_10916_n ) capacitor c=0.0195484f \
 //x=86.595 //y=1.645 //x2=86.025 //y2=1.495
cc_5358 ( N_QN_c_9105_n N_noxref_55_c_10917_n ) capacitor c=0.0069137f \
 //x=86.395 //y=1.18 //x2=86.91 //y2=0.53
cc_5359 ( N_QN_c_9113_n N_noxref_55_c_10917_n ) capacitor c=0.00458011f \
 //x=86.865 //y=1.645 //x2=86.91 //y2=0.53
cc_5360 ( N_QN_M53_noxref_d N_noxref_55_c_10917_n ) capacitor c=0.0132979f \
 //x=86.32 //y=0.905 //x2=86.91 //y2=0.53
cc_5361 ( N_QN_c_9105_n N_noxref_55_M52_noxref_s ) capacitor c=0.0513705f \
 //x=86.395 //y=1.18 //x2=84.92 //y2=0.365
cc_5362 ( N_QN_c_9113_n N_noxref_55_M52_noxref_s ) capacitor c=0.0155576f \
 //x=86.865 //y=1.645 //x2=84.92 //y2=0.365
cc_5363 ( N_QN_M53_noxref_d N_noxref_55_M52_noxref_s ) capacitor c=0.0438441f \
 //x=86.32 //y=0.905 //x2=84.92 //y2=0.365
cc_5364 ( N_noxref_23_c_9273_n N_noxref_24_c_9312_n ) capacitor c=0.0136048f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_5365 ( N_noxref_23_c_9290_n N_noxref_24_c_9312_n ) capacitor c=0.0102225f \
 //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_5366 ( N_noxref_23_M0_noxref_s N_noxref_24_c_9312_n ) capacitor \
 c=0.0228676f //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_5367 ( N_noxref_23_M0_noxref_s N_noxref_24_c_9314_n ) capacitor \
 c=0.0180035f //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_5368 ( N_noxref_23_c_9273_n N_noxref_24_M1_noxref_d ) capacitor \
 c=0.0129526f //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_5369 ( N_noxref_23_c_9290_n N_noxref_24_M1_noxref_d ) capacitor \
 c=0.00908243f //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_5370 ( N_noxref_23_M0_noxref_s N_noxref_24_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_5371 ( N_noxref_23_M0_noxref_s N_noxref_24_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_5372 ( N_noxref_24_c_9319_n N_noxref_25_M3_noxref_s ) capacitor \
 c=0.00191848f //x=4.07 //y=0.625 //x2=5.265 //y2=0.375
cc_5373 ( N_noxref_25_c_9371_n N_noxref_26_c_9416_n ) capacitor c=0.013301f \
 //x=7.255 //y=0.54 //x2=7.825 //y2=0.995
cc_5374 ( N_noxref_25_c_9381_n N_noxref_26_c_9416_n ) capacitor c=0.0100026f \
 //x=7.255 //y=1.59 //x2=7.825 //y2=0.995
cc_5375 ( N_noxref_25_M3_noxref_s N_noxref_26_c_9416_n ) capacitor \
 c=0.0224457f //x=5.265 //y=0.375 //x2=7.825 //y2=0.995
cc_5376 ( N_noxref_25_M3_noxref_s N_noxref_26_c_9418_n ) capacitor \
 c=0.0180035f //x=5.265 //y=0.375 //x2=7.91 //y2=0.625
cc_5377 ( N_noxref_25_c_9371_n N_noxref_26_M4_noxref_d ) capacitor \
 c=0.0128591f //x=7.255 //y=0.54 //x2=6.67 //y2=0.91
cc_5378 ( N_noxref_25_c_9381_n N_noxref_26_M4_noxref_d ) capacitor \
 c=0.00891456f //x=7.255 //y=1.59 //x2=6.67 //y2=0.91
cc_5379 ( N_noxref_25_M3_noxref_s N_noxref_26_M4_noxref_d ) capacitor \
 c=0.0159202f //x=5.265 //y=0.375 //x2=6.67 //y2=0.91
cc_5380 ( N_noxref_25_M3_noxref_s N_noxref_26_M5_noxref_s ) capacitor \
 c=0.0213553f //x=5.265 //y=0.375 //x2=7.775 //y2=0.375
cc_5381 ( N_noxref_26_c_9423_n N_noxref_27_M6_noxref_s ) capacitor \
 c=0.00164795f //x=8.88 //y=0.625 //x2=10.18 //y2=0.365
cc_5382 ( N_noxref_27_c_9479_n N_noxref_28_M8_noxref_s ) capacitor \
 c=0.00199452f //x=12.255 //y=0.615 //x2=13.405 //y2=0.375
cc_5383 ( N_noxref_28_c_9527_n N_noxref_29_c_9569_n ) capacitor c=0.0131877f \
 //x=15.395 //y=0.54 //x2=15.965 //y2=0.995
cc_5384 ( N_noxref_28_c_9550_n N_noxref_29_c_9569_n ) capacitor c=0.00981707f \
 //x=15.395 //y=1.59 //x2=15.965 //y2=0.995
cc_5385 ( N_noxref_28_M8_noxref_s N_noxref_29_c_9569_n ) capacitor \
 c=0.0221661f //x=13.405 //y=0.375 //x2=15.965 //y2=0.995
cc_5386 ( N_noxref_28_M8_noxref_s N_noxref_29_c_9571_n ) capacitor \
 c=0.0180035f //x=13.405 //y=0.375 //x2=16.05 //y2=0.625
cc_5387 ( N_noxref_28_c_9527_n N_noxref_29_M9_noxref_d ) capacitor \
 c=0.0127191f //x=15.395 //y=0.54 //x2=14.81 //y2=0.91
cc_5388 ( N_noxref_28_c_9550_n N_noxref_29_M9_noxref_d ) capacitor \
 c=0.00861161f //x=15.395 //y=1.59 //x2=14.81 //y2=0.91
cc_5389 ( N_noxref_28_M8_noxref_s N_noxref_29_M9_noxref_d ) capacitor \
 c=0.0159202f //x=13.405 //y=0.375 //x2=14.81 //y2=0.91
cc_5390 ( N_noxref_28_M8_noxref_s N_noxref_29_M10_noxref_s ) capacitor \
 c=0.0213553f //x=13.405 //y=0.375 //x2=15.915 //y2=0.375
cc_5391 ( N_noxref_29_c_9576_n N_noxref_30_M11_noxref_s ) capacitor \
 c=0.00191848f //x=17.02 //y=0.625 //x2=18.215 //y2=0.375
cc_5392 ( N_noxref_30_c_9629_n N_noxref_31_c_9674_n ) capacitor c=0.0131801f \
 //x=20.205 //y=0.54 //x2=20.775 //y2=0.995
cc_5393 ( N_noxref_30_c_9654_n N_noxref_31_c_9674_n ) capacitor c=0.00980353f \
 //x=20.205 //y=1.59 //x2=20.775 //y2=0.995
cc_5394 ( N_noxref_30_M11_noxref_s N_noxref_31_c_9674_n ) capacitor \
 c=0.0221661f //x=18.215 //y=0.375 //x2=20.775 //y2=0.995
cc_5395 ( N_noxref_30_M11_noxref_s N_noxref_31_c_9676_n ) capacitor \
 c=0.0180035f //x=18.215 //y=0.375 //x2=20.86 //y2=0.625
cc_5396 ( N_noxref_30_c_9629_n N_noxref_31_M12_noxref_d ) capacitor \
 c=0.0127176f //x=20.205 //y=0.54 //x2=19.62 //y2=0.91
cc_5397 ( N_noxref_30_c_9654_n N_noxref_31_M12_noxref_d ) capacitor \
 c=0.0086073f //x=20.205 //y=1.59 //x2=19.62 //y2=0.91
cc_5398 ( N_noxref_30_M11_noxref_s N_noxref_31_M12_noxref_d ) capacitor \
 c=0.0159202f //x=18.215 //y=0.375 //x2=19.62 //y2=0.91
cc_5399 ( N_noxref_30_M11_noxref_s N_noxref_31_M13_noxref_s ) capacitor \
 c=0.0213553f //x=18.215 //y=0.375 //x2=20.725 //y2=0.375
cc_5400 ( N_noxref_31_c_9681_n N_noxref_32_M14_noxref_s ) capacitor \
 c=0.00164795f //x=21.83 //y=0.625 //x2=23.13 //y2=0.365
cc_5401 ( N_noxref_32_c_9736_n N_noxref_33_M16_noxref_s ) capacitor \
 c=0.00199452f //x=25.205 //y=0.615 //x2=26.355 //y2=0.375
cc_5402 ( N_noxref_33_c_9784_n N_noxref_34_c_9826_n ) capacitor c=0.0131877f \
 //x=28.345 //y=0.54 //x2=28.915 //y2=0.995
cc_5403 ( N_noxref_33_c_9805_n N_noxref_34_c_9826_n ) capacitor c=0.00981707f \
 //x=28.345 //y=1.59 //x2=28.915 //y2=0.995
cc_5404 ( N_noxref_33_M16_noxref_s N_noxref_34_c_9826_n ) capacitor \
 c=0.0221661f //x=26.355 //y=0.375 //x2=28.915 //y2=0.995
cc_5405 ( N_noxref_33_M16_noxref_s N_noxref_34_c_9828_n ) capacitor \
 c=0.0180035f //x=26.355 //y=0.375 //x2=29 //y2=0.625
cc_5406 ( N_noxref_33_c_9784_n N_noxref_34_M17_noxref_d ) capacitor \
 c=0.0127191f //x=28.345 //y=0.54 //x2=27.76 //y2=0.91
cc_5407 ( N_noxref_33_c_9805_n N_noxref_34_M17_noxref_d ) capacitor \
 c=0.00861161f //x=28.345 //y=1.59 //x2=27.76 //y2=0.91
cc_5408 ( N_noxref_33_M16_noxref_s N_noxref_34_M17_noxref_d ) capacitor \
 c=0.0159202f //x=26.355 //y=0.375 //x2=27.76 //y2=0.91
cc_5409 ( N_noxref_33_M16_noxref_s N_noxref_34_M18_noxref_s ) capacitor \
 c=0.0213553f //x=26.355 //y=0.375 //x2=28.865 //y2=0.375
cc_5410 ( N_noxref_34_c_9833_n N_noxref_35_M19_noxref_s ) capacitor \
 c=0.00191848f //x=29.97 //y=0.625 //x2=31.165 //y2=0.375
cc_5411 ( N_noxref_35_c_9885_n N_noxref_36_c_9927_n ) capacitor c=0.0131877f \
 //x=33.155 //y=0.54 //x2=33.725 //y2=0.995
cc_5412 ( N_noxref_35_c_9908_n N_noxref_36_c_9927_n ) capacitor c=0.00981707f \
 //x=33.155 //y=1.59 //x2=33.725 //y2=0.995
cc_5413 ( N_noxref_35_M19_noxref_s N_noxref_36_c_9927_n ) capacitor \
 c=0.0221661f //x=31.165 //y=0.375 //x2=33.725 //y2=0.995
cc_5414 ( N_noxref_35_M19_noxref_s N_noxref_36_c_9929_n ) capacitor \
 c=0.0180035f //x=31.165 //y=0.375 //x2=33.81 //y2=0.625
cc_5415 ( N_noxref_35_c_9885_n N_noxref_36_M20_noxref_d ) capacitor \
 c=0.0127191f //x=33.155 //y=0.54 //x2=32.57 //y2=0.91
cc_5416 ( N_noxref_35_c_9908_n N_noxref_36_M20_noxref_d ) capacitor \
 c=0.00861161f //x=33.155 //y=1.59 //x2=32.57 //y2=0.91
cc_5417 ( N_noxref_35_M19_noxref_s N_noxref_36_M20_noxref_d ) capacitor \
 c=0.0159202f //x=31.165 //y=0.375 //x2=32.57 //y2=0.91
cc_5418 ( N_noxref_35_M19_noxref_s N_noxref_36_M21_noxref_s ) capacitor \
 c=0.0213553f //x=31.165 //y=0.375 //x2=33.675 //y2=0.375
cc_5419 ( N_noxref_36_c_9934_n N_noxref_37_M22_noxref_s ) capacitor \
 c=0.00164795f //x=34.78 //y=0.625 //x2=36.08 //y2=0.365
cc_5420 ( N_noxref_37_c_9990_n N_noxref_38_M24_noxref_s ) capacitor \
 c=0.00199452f //x=38.155 //y=0.615 //x2=39.305 //y2=0.375
cc_5421 ( N_noxref_38_c_10038_n N_noxref_39_c_10080_n ) capacitor c=0.0131877f \
 //x=41.295 //y=0.54 //x2=41.865 //y2=0.995
cc_5422 ( N_noxref_38_c_10061_n N_noxref_39_c_10080_n ) capacitor \
 c=0.00981707f //x=41.295 //y=1.59 //x2=41.865 //y2=0.995
cc_5423 ( N_noxref_38_M24_noxref_s N_noxref_39_c_10080_n ) capacitor \
 c=0.0221661f //x=39.305 //y=0.375 //x2=41.865 //y2=0.995
cc_5424 ( N_noxref_38_M24_noxref_s N_noxref_39_c_10082_n ) capacitor \
 c=0.0180035f //x=39.305 //y=0.375 //x2=41.95 //y2=0.625
cc_5425 ( N_noxref_38_c_10038_n N_noxref_39_M25_noxref_d ) capacitor \
 c=0.0127191f //x=41.295 //y=0.54 //x2=40.71 //y2=0.91
cc_5426 ( N_noxref_38_c_10061_n N_noxref_39_M25_noxref_d ) capacitor \
 c=0.00861161f //x=41.295 //y=1.59 //x2=40.71 //y2=0.91
cc_5427 ( N_noxref_38_M24_noxref_s N_noxref_39_M25_noxref_d ) capacitor \
 c=0.0159202f //x=39.305 //y=0.375 //x2=40.71 //y2=0.91
cc_5428 ( N_noxref_38_M24_noxref_s N_noxref_39_M26_noxref_s ) capacitor \
 c=0.0213553f //x=39.305 //y=0.375 //x2=41.815 //y2=0.375
cc_5429 ( N_noxref_39_c_10087_n N_noxref_40_M27_noxref_s ) capacitor \
 c=0.00191848f //x=42.92 //y=0.625 //x2=44.115 //y2=0.375
cc_5430 ( N_noxref_40_c_10140_n N_noxref_41_c_10185_n ) capacitor c=0.0131801f \
 //x=46.105 //y=0.54 //x2=46.675 //y2=0.995
cc_5431 ( N_noxref_40_c_10165_n N_noxref_41_c_10185_n ) capacitor \
 c=0.00980353f //x=46.105 //y=1.59 //x2=46.675 //y2=0.995
cc_5432 ( N_noxref_40_M27_noxref_s N_noxref_41_c_10185_n ) capacitor \
 c=0.0221661f //x=44.115 //y=0.375 //x2=46.675 //y2=0.995
cc_5433 ( N_noxref_40_M27_noxref_s N_noxref_41_c_10187_n ) capacitor \
 c=0.0180035f //x=44.115 //y=0.375 //x2=46.76 //y2=0.625
cc_5434 ( N_noxref_40_c_10140_n N_noxref_41_M28_noxref_d ) capacitor \
 c=0.0127176f //x=46.105 //y=0.54 //x2=45.52 //y2=0.91
cc_5435 ( N_noxref_40_c_10165_n N_noxref_41_M28_noxref_d ) capacitor \
 c=0.0086073f //x=46.105 //y=1.59 //x2=45.52 //y2=0.91
cc_5436 ( N_noxref_40_M27_noxref_s N_noxref_41_M28_noxref_d ) capacitor \
 c=0.0159202f //x=44.115 //y=0.375 //x2=45.52 //y2=0.91
cc_5437 ( N_noxref_40_M27_noxref_s N_noxref_41_M29_noxref_s ) capacitor \
 c=0.0213553f //x=44.115 //y=0.375 //x2=46.625 //y2=0.375
cc_5438 ( N_noxref_41_c_10192_n N_noxref_42_M30_noxref_s ) capacitor \
 c=0.00164795f //x=47.73 //y=0.625 //x2=49.03 //y2=0.365
cc_5439 ( N_noxref_42_c_10247_n N_noxref_43_M32_noxref_s ) capacitor \
 c=0.00199452f //x=51.105 //y=0.615 //x2=52.255 //y2=0.375
cc_5440 ( N_noxref_43_c_10295_n N_noxref_44_c_10337_n ) capacitor c=0.0131877f \
 //x=54.245 //y=0.54 //x2=54.815 //y2=0.995
cc_5441 ( N_noxref_43_c_10305_n N_noxref_44_c_10337_n ) capacitor \
 c=0.00981707f //x=54.245 //y=1.59 //x2=54.815 //y2=0.995
cc_5442 ( N_noxref_43_M32_noxref_s N_noxref_44_c_10337_n ) capacitor \
 c=0.0221661f //x=52.255 //y=0.375 //x2=54.815 //y2=0.995
cc_5443 ( N_noxref_43_M32_noxref_s N_noxref_44_c_10339_n ) capacitor \
 c=0.0180035f //x=52.255 //y=0.375 //x2=54.9 //y2=0.625
cc_5444 ( N_noxref_43_c_10295_n N_noxref_44_M33_noxref_d ) capacitor \
 c=0.0127191f //x=54.245 //y=0.54 //x2=53.66 //y2=0.91
cc_5445 ( N_noxref_43_c_10305_n N_noxref_44_M33_noxref_d ) capacitor \
 c=0.00861161f //x=54.245 //y=1.59 //x2=53.66 //y2=0.91
cc_5446 ( N_noxref_43_M32_noxref_s N_noxref_44_M33_noxref_d ) capacitor \
 c=0.0159202f //x=52.255 //y=0.375 //x2=53.66 //y2=0.91
cc_5447 ( N_noxref_43_M32_noxref_s N_noxref_44_M34_noxref_s ) capacitor \
 c=0.0213553f //x=52.255 //y=0.375 //x2=54.765 //y2=0.375
cc_5448 ( N_noxref_44_c_10344_n N_noxref_45_M35_noxref_s ) capacitor \
 c=0.00191848f //x=55.87 //y=0.625 //x2=57.065 //y2=0.375
cc_5449 ( N_noxref_45_c_10396_n N_noxref_46_c_10438_n ) capacitor c=0.0131877f \
 //x=59.055 //y=0.54 //x2=59.625 //y2=0.995
cc_5450 ( N_noxref_45_c_10406_n N_noxref_46_c_10438_n ) capacitor \
 c=0.00981707f //x=59.055 //y=1.59 //x2=59.625 //y2=0.995
cc_5451 ( N_noxref_45_M35_noxref_s N_noxref_46_c_10438_n ) capacitor \
 c=0.0221661f //x=57.065 //y=0.375 //x2=59.625 //y2=0.995
cc_5452 ( N_noxref_45_M35_noxref_s N_noxref_46_c_10440_n ) capacitor \
 c=0.0180035f //x=57.065 //y=0.375 //x2=59.71 //y2=0.625
cc_5453 ( N_noxref_45_c_10396_n N_noxref_46_M36_noxref_d ) capacitor \
 c=0.0127191f //x=59.055 //y=0.54 //x2=58.47 //y2=0.91
cc_5454 ( N_noxref_45_c_10406_n N_noxref_46_M36_noxref_d ) capacitor \
 c=0.00861161f //x=59.055 //y=1.59 //x2=58.47 //y2=0.91
cc_5455 ( N_noxref_45_M35_noxref_s N_noxref_46_M36_noxref_d ) capacitor \
 c=0.0159202f //x=57.065 //y=0.375 //x2=58.47 //y2=0.91
cc_5456 ( N_noxref_45_M35_noxref_s N_noxref_46_M37_noxref_s ) capacitor \
 c=0.0213553f //x=57.065 //y=0.375 //x2=59.575 //y2=0.375
cc_5457 ( N_noxref_46_c_10445_n N_noxref_47_M38_noxref_s ) capacitor \
 c=0.00164795f //x=60.68 //y=0.625 //x2=61.98 //y2=0.365
cc_5458 ( N_noxref_47_c_10501_n N_noxref_48_M40_noxref_s ) capacitor \
 c=0.00199452f //x=64.055 //y=0.615 //x2=65.205 //y2=0.375
cc_5459 ( N_noxref_48_c_10549_n N_noxref_49_c_10591_n ) capacitor c=0.0131877f \
 //x=67.195 //y=0.54 //x2=67.765 //y2=0.995
cc_5460 ( N_noxref_48_c_10559_n N_noxref_49_c_10591_n ) capacitor \
 c=0.00981707f //x=67.195 //y=1.59 //x2=67.765 //y2=0.995
cc_5461 ( N_noxref_48_M40_noxref_s N_noxref_49_c_10591_n ) capacitor \
 c=0.0221661f //x=65.205 //y=0.375 //x2=67.765 //y2=0.995
cc_5462 ( N_noxref_48_M40_noxref_s N_noxref_49_c_10593_n ) capacitor \
 c=0.0180035f //x=65.205 //y=0.375 //x2=67.85 //y2=0.625
cc_5463 ( N_noxref_48_c_10549_n N_noxref_49_M41_noxref_d ) capacitor \
 c=0.0127191f //x=67.195 //y=0.54 //x2=66.61 //y2=0.91
cc_5464 ( N_noxref_48_c_10559_n N_noxref_49_M41_noxref_d ) capacitor \
 c=0.00861161f //x=67.195 //y=1.59 //x2=66.61 //y2=0.91
cc_5465 ( N_noxref_48_M40_noxref_s N_noxref_49_M41_noxref_d ) capacitor \
 c=0.0159202f //x=65.205 //y=0.375 //x2=66.61 //y2=0.91
cc_5466 ( N_noxref_48_M40_noxref_s N_noxref_49_M42_noxref_s ) capacitor \
 c=0.0213553f //x=65.205 //y=0.375 //x2=67.715 //y2=0.375
cc_5467 ( N_noxref_49_c_10598_n N_noxref_50_M43_noxref_s ) capacitor \
 c=0.00191848f //x=68.82 //y=0.625 //x2=70.015 //y2=0.375
cc_5468 ( N_noxref_50_c_10651_n N_noxref_51_c_10695_n ) capacitor c=0.0132328f \
 //x=72.005 //y=0.54 //x2=72.575 //y2=0.995
cc_5469 ( N_noxref_50_c_10673_n N_noxref_51_c_10695_n ) capacitor \
 c=0.00988406f //x=72.005 //y=1.59 //x2=72.575 //y2=0.995
cc_5470 ( N_noxref_50_M43_noxref_s N_noxref_51_c_10695_n ) capacitor \
 c=0.0226274f //x=70.015 //y=0.375 //x2=72.575 //y2=0.995
cc_5471 ( N_noxref_50_M43_noxref_s N_noxref_51_c_10697_n ) capacitor \
 c=0.0180035f //x=70.015 //y=0.375 //x2=72.66 //y2=0.625
cc_5472 ( N_noxref_50_c_10651_n N_noxref_51_M44_noxref_d ) capacitor \
 c=0.0127176f //x=72.005 //y=0.54 //x2=71.42 //y2=0.91
cc_5473 ( N_noxref_50_c_10673_n N_noxref_51_M44_noxref_d ) capacitor \
 c=0.0086073f //x=72.005 //y=1.59 //x2=71.42 //y2=0.91
cc_5474 ( N_noxref_50_M43_noxref_s N_noxref_51_M44_noxref_d ) capacitor \
 c=0.0159202f //x=70.015 //y=0.375 //x2=71.42 //y2=0.91
cc_5475 ( N_noxref_50_M43_noxref_s N_noxref_51_M45_noxref_s ) capacitor \
 c=0.0213553f //x=70.015 //y=0.375 //x2=72.525 //y2=0.375
cc_5476 ( N_noxref_51_c_10702_n N_noxref_52_M46_noxref_s ) capacitor \
 c=0.00164795f //x=73.63 //y=0.625 //x2=74.93 //y2=0.365
cc_5477 ( N_noxref_52_c_10757_n N_noxref_53_M48_noxref_s ) capacitor \
 c=0.00205929f //x=77.005 //y=0.615 //x2=78.26 //y2=0.365
cc_5478 ( N_noxref_53_M48_noxref_s N_noxref_54_c_10872_n ) capacitor \
 c=0.0011299f //x=78.26 //y=0.365 //x2=81.725 //y2=1.495
cc_5479 ( N_noxref_53_c_10808_n N_noxref_54_M50_noxref_s ) capacitor \
 c=0.0011299f //x=80.335 //y=0.615 //x2=81.59 //y2=0.365
cc_5480 ( N_noxref_54_M50_noxref_s N_noxref_55_c_10937_n ) capacitor \
 c=0.0011299f //x=81.59 //y=0.365 //x2=85.055 //y2=1.495
cc_5481 ( N_noxref_54_c_10864_n N_noxref_55_M52_noxref_s ) capacitor \
 c=0.0011299f //x=83.665 //y=0.615 //x2=84.92 //y2=0.365
