* SPICE3 file created from VOTERN3X1.ext - technology: sky130A

.subckt VOTERN3X1 YN A B C VDD GND
X0 GND B votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X1 GND B votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X2 GND C votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X3 votern3x1_pcell_0/a_805_1331# B VDD VDD pshort w=2 l=0.15
X4 YN C votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X5 votern3x1_pcell_0/a_805_1331# A VDD VDD pshort w=2 l=0.15
X6 votern3x1_pcell_0/a_893_1059# C votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X7 votern3x1_pcell_0/a_893_1059# B votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X8 YN C votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X9 YN A votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X10 YN A votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X11 YN A votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
C0 VDD GND 18.63fF
.ends
