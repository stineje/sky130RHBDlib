magic
tech sky130A
magscale 1 2
timestamp 1670370157
<< error_s >>
rect 198 296 214 312
rect 392 296 408 312
rect 586 296 602 312
rect 1147 297 1163 313
rect 274 266 304 296
rect 468 266 498 296
rect 662 266 692 296
rect 1223 267 1253 297
rect 198 250 214 266
rect 258 250 274 266
rect 393 252 408 266
rect 392 251 408 252
rect 452 252 467 266
rect 587 252 602 266
rect 452 251 468 252
rect 586 251 602 252
rect 646 252 661 266
rect 646 251 662 252
rect 1147 251 1163 267
rect 1207 251 1223 267
rect 391 250 392 251
rect 468 250 469 251
rect 585 250 586 251
rect 662 250 663 251
rect 198 165 214 181
rect 258 165 274 181
rect 392 165 408 181
rect 452 165 468 181
rect 586 165 602 181
rect 646 165 662 181
rect 1147 166 1163 182
rect 1207 166 1223 182
rect 168 135 198 165
rect 274 135 304 165
rect 362 135 392 165
rect 468 135 498 165
rect 556 135 586 165
rect 662 135 692 165
rect 1117 136 1147 166
rect 1223 136 1253 166
<< locali >>
rect 205 871 239 905
rect 353 871 387 905
rect 575 871 609 905
rect 1241 871 1275 905
rect 205 797 239 831
rect 353 797 387 831
rect 575 797 609 831
rect 1241 797 1275 831
rect 205 723 239 757
rect 353 723 387 757
rect 575 723 609 757
rect 1241 723 1275 757
rect 205 649 239 683
rect 353 649 387 683
rect 575 649 609 683
rect 1241 649 1275 683
rect 205 575 239 609
rect 353 575 387 609
rect 575 575 609 609
rect 1241 575 1275 609
rect 205 501 239 535
rect 353 501 387 535
rect 575 501 609 535
rect 1241 501 1275 535
rect 205 427 239 461
rect 353 427 387 461
rect 575 427 609 461
rect 1241 427 1275 461
use or3x1_pcell  or3x1_pcell_0 pcells
timestamp 1670369097
transform 1 0 296 0 1 0
box -383 -34 1197 1550
<< labels >>
rlabel locali 1241 427 1275 461 1 Y
port 1 nsew signal output
rlabel locali 1241 501 1275 535 1 Y
port 1 nsew signal output
rlabel locali 1241 575 1275 609 1 Y
port 1 nsew signal output
rlabel locali 1241 649 1275 683 1 Y
port 1 nsew signal output
rlabel locali 1241 723 1275 757 1 Y
port 1 nsew signal output
rlabel locali 1241 797 1275 831 1 Y
port 1 nsew signal output
rlabel locali 1241 871 1275 905 1 Y
port 1 nsew signal output
rlabel locali 205 871 239 905 1 A
port 2 nsew signal input
rlabel locali 205 797 239 831 1 A
port 2 nsew signal input
rlabel locali 205 723 239 757 1 A
port 2 nsew signal input
rlabel locali 205 649 239 683 1 A
port 2 nsew signal input
rlabel locali 205 575 239 609 1 A
port 2 nsew signal input
rlabel locali 205 501 239 535 1 A
port 2 nsew signal input
rlabel locali 205 427 239 461 1 A
port 2 nsew signal input
rlabel locali 353 871 387 905 1 B
port 3 nsew signal input
rlabel locali 353 797 387 831 1 B
port 3 nsew signal input
rlabel locali 353 723 387 757 1 B
port 3 nsew signal input
rlabel locali 353 649 387 683 1 B
port 3 nsew signal input
rlabel locali 353 575 387 609 1 B
port 3 nsew signal input
rlabel locali 353 501 387 535 1 B
port 3 nsew signal input
rlabel locali 353 427 387 461 1 B
port 3 nsew signal input
rlabel locali 575 871 609 905 1 C
port 4 nsew signal output
rlabel locali 575 797 609 831 1 C
port 4 nsew signal input
rlabel locali 575 723 609 757 1 C
port 4 nsew signal input
rlabel locali 575 649 609 683 1 C
port 4 nsew signal input
rlabel locali 575 575 609 609 1 C
port 4 nsew signal input
rlabel locali 575 501 609 535 1 C
port 4 nsew signal input
rlabel locali 575 427 609 461 1 C
port 4 nsew signal input
rlabel space -34 1446 1440 1514 1 VDD
port 5 nsew power bidirectional abutment
rlabel space -34 -34 1440 34 1 GND
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1406 1480
string LEFclass CORE
string LEFsite unitrh
string LEFsymmetry X Y R90
<< end >>
