* SPICE3 file created from VOTERN3X1.ext - technology: sky130A

.subckt VOTERN3X1 YN A B C VDD GND
X0 GND B a_112_73 GND nshort w=3 l=0.15
X1 GND C a_1444_73 GND nshort w=3 l=0.15
X2 YN A a_1444_73 GND nshort w=3 l=0.15
X3 YN A a_881_1005 VDD pshort w=2 l=0.15 M=2
X4 VDD B a_217_1005 VDD pshort w=2 l=0.15 M=2
X5 a_881_1005 C a_217_1005 VDD pshort w=2 l=0.15 M=2
X6 VDD A a_217_1005 VDD pshort w=2 l=0.15 M=2
X7 YN A a_112_73 GND nshort w=3 l=0.15
X8 a_881_1005 B a_217_1005 VDD pshort w=2 l=0.15 M=2
X9 a_881_1005 C YN VDD pshort w=2 l=0.15 M=2
X10 YN C a_778_73 GND nshort w=3 l=0.15
X11 GND B a_778_73 GND nshort w=3 l=0.15
C0 VDD GND 5.10fF
.ends
