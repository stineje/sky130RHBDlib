magic
tech sky130A
magscale 1 2
timestamp 1648739814
<< metal1 >>
rect 426 945 2981 979
rect 241 871 4901 905
rect 867 797 3782 831
rect 689 723 2174 757
rect 2461 723 2785 757
rect 1607 501 3963 535
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 222 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 666 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 444 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 814 0 -1 814
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_1
timestamp 1648064657
transform 1 0 962 0 1 0
box -84 0 1046 1575
use nand3x1_pcell  nand3x1_pcell_0
timestamp 1648064657
transform 1 0 0 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 1628 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform -1 0 1184 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 2146 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform -1 0 1776 0 -1 740
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_0
timestamp 1648064633
transform 1 0 1924 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform 1 0 2812 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform -1 0 2442 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform 1 0 2294 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 3034 0 1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform -1 0 3256 0 -1 518
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_3
timestamp 1648064657
transform 1 0 2590 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 3774 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform 1 0 3404 0 1 888
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_1
timestamp 1648064633
transform 1 0 4514 0 1 0
box -84 0 750 1575
use li1_M1_contact  li1_M1_contact_18
timestamp 1648061256
transform 1 0 3996 0 1 518
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_4
timestamp 1648064657
transform 1 0 3552 0 1 0
box -84 0 1046 1575
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform 1 0 4884 0 1 888
box -53 -33 29 33
<< end >>
