* SPICE3 file created from VOTERN3X1.ext - technology: sky130A

.subckt VOTERN3X1 YN A B C VDD VSS
X0 YN A a_881_1051 VDD sky130_fd_pr__pfet_01v8 ad=0.00116 pd=9.16 as=0 ps=0 w=2 l=0.15 M=2
X1 VDD B a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0.00168 pd=1.368 as=0 ps=0 w=2 l=0.15 M=2
X2 a_881_1051 C a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X3 VSS B a_778_101 VSS sky130_fd_pr__nfet_01v8 ad=0.005373 pd=4.71 as=0 ps=0 w=3 l=0.15
X4 VSS B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X5 VSS C a_1444_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X6 VDD A a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X7 a_881_1051 B a_217_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X8 a_881_1051 C YN VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X9 YN A a_1444_101 VSS sky130_fd_pr__nfet_01v8 ad=0.005373 pd=4.72 as=0 ps=0 w=3 l=0.15
X10 YN A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X11 YN C a_778_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 VDD a_217_1051 3.12f
C1 VDD VSS 4.20f
.ends
