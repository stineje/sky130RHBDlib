* NGSPICE file created from INVX1.ext - technology: sky130A

.subckt INVX1 Y A VPWR VGND
X0 Y A VGND VGND sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=1.1408p ps=8.1u L=0.15 W=3
X1 VPWR A Y VPWR sky130_fd_pr__pfet_01v8 ad=1.1p pd=9.1u as=5.8p ps=4.58u L=0.15 W=2 M=2
C0 Y VPWR 1.04fF
C1 A VPWR 0.38fF
C2 Y A 0.28fF
.ends
