* SPICE3 file created from DFFRNX1.ext - technology: sky130A

.subckt DFFRNX1 Q QN D CLK RN GND
X0 GND dffrnx1_pcell_0/m1_241_797# dffrnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 dffrnx1_pcell_0/m1_867_723# dffrnx1_pcell_0/m1_689_649# dffrnx1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X2 dffrnx1_pcell_0/nand3x1_pcell_0/li_393_182# CLK dffrnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X3 VDD dffrnx1_pcell_0/m1_241_797# dffrnx1_pcell_0/m1_867_723# VDD pshort w=2 l=0.15
X4 VDD CLK dffrnx1_pcell_0/m1_867_723# VDD pshort w=2 l=0.15
X5 VDD dffrnx1_pcell_0/m1_689_649# dffrnx1_pcell_0/m1_867_723# VDD pshort w=2 l=0.15
X6 GND dffrnx1_pcell_0/m1_867_723# dffrnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X7 dffrnx1_pcell_0/m1_689_649# RN dffrnx1_pcell_0/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X8 dffrnx1_pcell_0/nand3x1_pcell_1/li_393_182# D dffrnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X9 VDD dffrnx1_pcell_0/m1_867_723# dffrnx1_pcell_0/m1_689_649# VDD pshort w=2 l=0.15
X10 VDD D dffrnx1_pcell_0/m1_689_649# VDD pshort w=2 l=0.15
X11 VDD RN dffrnx1_pcell_0/m1_689_649# VDD pshort w=2 l=0.15
X12 GND dffrnx1_pcell_0/m1_2461_649# dffrnx1_pcell_0/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X13 dffrnx1_pcell_0/m1_241_797# RN dffrnx1_pcell_0/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X14 dffrnx1_pcell_0/nand3x1_pcell_3/li_393_182# CLK dffrnx1_pcell_0/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X15 VDD dffrnx1_pcell_0/m1_2461_649# dffrnx1_pcell_0/m1_241_797# VDD pshort w=2 l=0.15
X16 VDD CLK dffrnx1_pcell_0/m1_241_797# VDD pshort w=2 l=0.15
X17 VDD RN dffrnx1_pcell_0/m1_241_797# VDD pshort w=2 l=0.15
X18 GND dffrnx1_pcell_0/m1_867_723# dffrnx1_pcell_0/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X19 QN Q dffrnx1_pcell_0/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X20 dffrnx1_pcell_0/nand3x1_pcell_4/li_393_182# RN dffrnx1_pcell_0/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X21 VDD dffrnx1_pcell_0/m1_867_723# QN VDD pshort w=2 l=0.15
X22 VDD RN QN VDD pshort w=2 l=0.15
X23 VDD Q QN VDD pshort w=2 l=0.15
X24 GND dffrnx1_pcell_0/m1_689_649# dffrnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X25 dffrnx1_pcell_0/m1_2461_649# dffrnx1_pcell_0/m1_241_797# dffrnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X26 VDD dffrnx1_pcell_0/m1_689_649# dffrnx1_pcell_0/m1_2461_649# VDD pshort w=2 l=0.15
X27 VDD dffrnx1_pcell_0/m1_241_797# dffrnx1_pcell_0/m1_2461_649# VDD pshort w=2 l=0.15
X28 GND QN dffrnx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X29 Q dffrnx1_pcell_0/m1_241_797# dffrnx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X30 VDD QN Q VDD pshort w=2 l=0.15
X31 VDD dffrnx1_pcell_0/m1_241_797# Q VDD pshort w=2 l=0.15
C0 VDD dffrnx1_pcell_0/m1_241_797# 2.82fF
.ends
