magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -66 377 1506 897
<< pwell >>
rect 53 43 1433 317
rect -26 -43 1466 43
<< locali >>
rect 255 441 321 689
rect 567 441 633 689
rect 879 441 945 689
rect 1191 441 1257 689
rect 255 407 1422 441
rect 62 316 1352 363
rect 239 279 1245 280
rect 1388 279 1422 407
rect 239 246 1422 279
rect 239 146 281 246
rect 551 146 593 246
rect 863 146 905 246
rect 1183 245 1422 246
rect 1183 146 1313 245
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1440 831
rect 19 729 1405 759
rect 53 695 91 729
rect 125 695 163 729
rect 197 725 355 729
rect 19 489 197 695
rect 389 695 427 729
rect 461 695 499 729
rect 533 725 667 729
rect 355 477 533 695
rect 701 695 739 729
rect 773 695 811 729
rect 845 725 979 729
rect 667 477 845 695
rect 1013 695 1051 729
rect 1085 695 1123 729
rect 1157 725 1291 729
rect 979 477 1157 695
rect 1325 695 1371 729
rect 1291 477 1405 695
rect 19 110 197 277
rect 315 110 517 209
rect 627 110 829 209
rect 939 110 1149 209
rect 1347 110 1421 209
rect 19 76 91 110
rect 125 76 163 110
rect 197 76 235 110
rect 269 76 307 110
rect 341 76 379 110
rect 413 76 451 110
rect 485 76 523 110
rect 557 76 595 110
rect 629 76 667 110
rect 701 76 739 110
rect 773 76 811 110
rect 845 76 883 110
rect 917 76 955 110
rect 989 76 1027 110
rect 1061 76 1099 110
rect 1133 76 1171 110
rect 1205 76 1243 110
rect 1277 76 1315 110
rect 1349 76 1387 110
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 19 695 53 729
rect 91 695 125 729
rect 163 695 197 729
rect 355 695 389 729
rect 427 695 461 729
rect 499 695 533 729
rect 667 695 701 729
rect 739 695 773 729
rect 811 695 845 729
rect 979 695 1013 729
rect 1051 695 1085 729
rect 1123 695 1157 729
rect 1291 695 1325 729
rect 1371 695 1405 729
rect 91 76 125 110
rect 163 76 197 110
rect 235 76 269 110
rect 307 76 341 110
rect 379 76 413 110
rect 451 76 485 110
rect 523 76 557 110
rect 595 76 629 110
rect 667 76 701 110
rect 739 76 773 110
rect 811 76 845 110
rect 883 76 917 110
rect 955 76 989 110
rect 1027 76 1061 110
rect 1099 76 1133 110
rect 1171 76 1205 110
rect 1243 76 1277 110
rect 1315 76 1349 110
rect 1387 76 1421 110
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
<< metal1 >>
rect 0 831 1440 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1440 831
rect 0 791 1440 797
rect 0 729 1440 763
rect 0 695 19 729
rect 53 695 91 729
rect 125 695 163 729
rect 197 695 355 729
rect 389 695 427 729
rect 461 695 499 729
rect 533 695 667 729
rect 701 695 739 729
rect 773 695 811 729
rect 845 695 979 729
rect 1013 695 1051 729
rect 1085 695 1123 729
rect 1157 695 1291 729
rect 1325 695 1371 729
rect 1405 695 1440 729
rect 0 689 1440 695
rect 0 110 1440 125
rect 0 76 91 110
rect 125 76 163 110
rect 197 76 235 110
rect 269 76 307 110
rect 341 76 379 110
rect 413 76 451 110
rect 485 76 523 110
rect 557 76 595 110
rect 629 76 667 110
rect 701 76 739 110
rect 773 76 811 110
rect 845 76 883 110
rect 917 76 955 110
rect 989 76 1027 110
rect 1061 76 1099 110
rect 1133 76 1171 110
rect 1205 76 1243 110
rect 1277 76 1315 110
rect 1349 76 1387 110
rect 1421 76 1440 110
rect 0 51 1440 76
rect 0 17 1440 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1440 17
rect 0 -23 1440 -17
<< labels >>
rlabel locali s 62 316 1352 363 6 A
port 1 nsew signal input
rlabel metal1 s 0 51 1440 125 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 -23 1440 23 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s -26 -43 1466 43 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 53 43 1433 317 6 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 791 1440 837 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -66 377 1506 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 1440 763 6 VPWR
port 5 nsew power bidirectional
rlabel locali s 1183 146 1313 245 6 Y
port 6 nsew signal output
rlabel locali s 1183 245 1422 246 6 Y
port 6 nsew signal output
rlabel locali s 863 146 905 246 6 Y
port 6 nsew signal output
rlabel locali s 551 146 593 246 6 Y
port 6 nsew signal output
rlabel locali s 239 146 281 246 6 Y
port 6 nsew signal output
rlabel locali s 239 246 1422 279 6 Y
port 6 nsew signal output
rlabel locali s 1388 279 1422 407 6 Y
port 6 nsew signal output
rlabel locali s 239 279 1245 280 6 Y
port 6 nsew signal output
rlabel locali s 255 407 1422 441 6 Y
port 6 nsew signal output
rlabel locali s 1191 441 1257 689 6 Y
port 6 nsew signal output
rlabel locali s 879 441 945 689 6 Y
port 6 nsew signal output
rlabel locali s 567 441 633 689 6 Y
port 6 nsew signal output
rlabel locali s 255 441 321 689 6 Y
port 6 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 1440 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 59604
string GDS_START 42586
<< end >>
