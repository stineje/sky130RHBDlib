magic
tech sky130A
magscale 1 2
timestamp 1653605740
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 205 871 239 905
rect 1093 871 1127 905
rect 2943 871 2977 905
rect 5977 871 6011 905
rect 7827 871 7861 905
rect 10861 871 10895 905
rect 12711 871 12745 905
rect 16929 871 16963 905
rect 205 797 239 831
rect 4349 797 4383 831
rect 5089 797 5123 831
rect 9973 797 10007 831
rect 16929 797 16963 831
rect 205 723 239 757
rect 1093 723 1127 757
rect 5089 723 5123 757
rect 5977 723 6011 757
rect 9973 723 10007 757
rect 10861 723 10895 757
rect 16929 723 16963 757
rect 205 649 239 683
rect 1093 649 1127 683
rect 2055 649 2089 683
rect 2943 649 2977 683
rect 16929 649 16963 683
rect 205 575 239 609
rect 5089 575 5123 609
rect 9973 575 10007 609
rect 16929 575 16963 609
rect 205 501 239 535
rect 2055 501 2089 535
rect 2943 501 2977 535
rect 4349 501 4383 535
rect 5089 501 5123 535
rect 7827 501 7861 535
rect 11823 501 11857 535
rect 12711 501 12745 535
rect 16929 501 16963 535
rect 1093 427 1127 461
rect 2055 427 2089 461
rect 4349 427 4383 461
rect 6939 427 6973 461
rect 9233 427 9267 461
rect 11823 427 11857 461
rect 14117 427 14151 461
rect 16929 427 16963 461
<< metal1 >>
rect -34 1446 17128 1514
rect 13561 945 13878 979
rect 1163 871 2907 905
rect 2989 871 5965 905
rect 6047 871 7791 905
rect 7873 871 10849 905
rect 10931 871 12675 905
rect 13413 871 15028 905
rect 3813 797 4132 831
rect 8522 797 9567 831
rect 3606 649 15819 683
rect 275 575 5077 609
rect 5159 575 9937 609
rect 10121 575 14969 609
rect 10121 535 10155 575
rect 8629 501 8975 535
rect 9639 501 10155 535
rect 2106 427 4343 461
rect 4389 427 6933 461
rect 6979 427 9227 461
rect 9273 427 11817 461
rect 11863 427 14111 461
rect -34 -34 17128 34
use li1_M1_contact  li1_M1_contact_18 pcells
timestamp 1648061256
transform 1 0 4144 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 3774 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform -1 0 222 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform -1 0 4736 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_20
timestamp 1648061256
transform -1 0 3626 0 -1 666
box -53 -33 29 33
use dffsnx1_pcell  dffsnx1_pcell_0 pcells
timestamp 1652396184
transform 1 0 0 0 1 0
box -87 -34 4971 1550
use dffsnx1_pcell  dffsnx1_pcell_1
timestamp 1652396184
transform 1 0 4884 0 1 0
box -87 -34 4971 1550
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 9620 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform 1 0 9620 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 8510 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 1 0 9028 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 8658 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 9990 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 5106 0 -1 592
box -53 -33 29 33
use dffsnx1_pcell  dffsnx1_pcell_2
timestamp 1652396184
transform 1 0 9768 0 1 0
box -87 -34 4971 1550
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform 1 0 15022 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 13542 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 13912 0 1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform 1 0 14504 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 13394 0 -1 888
box -53 -33 29 33
use voter3x1_pcell  voter3x1_pcell_0 pcells
timestamp 1652393968
transform 1 0 14652 0 1 0
box -87 -34 2529 1550
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform 1 0 15836 0 -1 666
box -53 -33 29 33
<< labels >>
rlabel locali 16929 797 16963 831 1 Q
port 1 nsew signal output
rlabel locali 16929 723 16963 757 1 Q
port 1 nsew signal output
rlabel locali 16929 649 16963 683 1 Q
port 1 nsew signal output
rlabel locali 16929 575 16963 609 1 Q
port 1 nsew signal output
rlabel locali 16929 501 16963 535 1 Q
port 1 nsew signal output
rlabel locali 16929 427 16963 461 1 Q
port 1 nsew signal output
rlabel locali 16929 871 16963 905 1 Q
port 1 nsew signal output
rlabel locali 5089 575 5123 609 1 D
port 2 nsew signal input
rlabel locali 5089 501 5123 535 1 D
port 2 nsew signal input
rlabel locali 5089 723 5123 757 1 D
port 2 nsew signal input
rlabel locali 5089 797 5123 831 1 D
port 2 nsew signal input
rlabel locali 9973 575 10007 609 1 D
port 2 nsew signal input
rlabel locali 9973 723 10007 757 1 D
port 2 nsew signal input
rlabel locali 9973 797 10007 831 1 D
port 2 nsew signal input
rlabel locali 205 575 239 609 1 D
port 2 nsew signal input
rlabel locali 205 649 239 683 1 D
port 2 nsew signal input
rlabel locali 205 723 239 757 1 D
port 2 nsew signal input
rlabel locali 205 797 239 831 1 D
port 2 nsew signal input
rlabel locali 205 871 239 905 1 D
port 2 nsew signal input
rlabel locali 205 501 239 535 1 D
port 2 nsew signal input
rlabel locali 1093 871 1127 905 1 CLK
port 3 nsew signal input
rlabel locali 1093 723 1127 757 1 CLK
port 3 nsew signal input
rlabel locali 1093 649 1127 683 1 CLK
port 3 nsew signal input
rlabel locali 1093 427 1127 461 1 CLK
port 3 nsew signal input
rlabel locali 2943 649 2977 683 1 CLK
port 3 nsew signal input
rlabel locali 2943 871 2977 905 1 CLK
port 3 nsew signal input
rlabel locali 2943 501 2977 535 1 CLK
port 3 nsew signal input
rlabel locali 5977 871 6011 905 1 CLK
port 3 nsew signal input
rlabel locali 7827 871 7861 905 1 CLK
port 3 nsew signal input
rlabel locali 7827 501 7861 535 1 CLK
port 3 nsew signal input
rlabel locali 5977 723 6011 757 1 CLK
port 3 nsew signal input
rlabel locali 10861 871 10895 905 1 CLK
port 3 nsew signal input
rlabel locali 12711 871 12745 905 1 CLK
port 3 nsew signal input
rlabel locali 12711 501 12745 535 1 CLK
port 3 nsew signal input
rlabel locali 10861 723 10895 757 1 CLK
port 3 nsew signal input
rlabel locali 2055 427 2089 461 1 SN
port 4 nsew signal input
rlabel locali 2055 501 2089 535 1 SN
port 4 nsew signal input
rlabel locali 2055 649 2089 683 1 SN
port 4 nsew signal input
rlabel locali 4349 427 4383 461 1 SN
port 4 nsew signal input
rlabel locali 4349 501 4383 535 1 SN
port 4 nsew signal input
rlabel locali 4349 797 4383 831 1 SN
port 4 nsew signal input
rlabel locali 6939 427 6973 461 1 SN
port 4 nsew signal input
rlabel locali 11823 427 11857 461 1 SN
port 4 nsew signal input
rlabel locali 11823 501 11857 535 1 SN
port 4 nsew signal input
rlabel locali 14117 427 14151 461 1 SN
port 4 nsew signal input
rlabel metal1 -34 1446 17128 1514 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 -34 -34 17128 34 1 GND
port 6 nsew ground bidirectional abutment
<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 17094 1480
string LEFsymmetry X Y R90
<< end >>
