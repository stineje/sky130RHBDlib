* SPICE3 file created from TIELO.ext - technology: sky130A

.subckt TIELO YN VDD GND
X0 YN a_155_381# GND GND nshort w=3 l=0.15
X1 VDD a_155_381# a_155_381# VDD pshort w=2 l=0.15
C0 VDD GND 2.23fF
.ends
