* SPICE3 file created from TMRDFFSNQX1.ext - technology: sky130A

.subckt TMRDFFSNQX1 Q D CLK SN VPB VNB
M1000 VPB.t67 CLK a_5227_383.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_15533_1005.t6 a_3599_383.t7 a_15044_181.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VNB D a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=4.9019p pd=41.07u as=0p ps=0u
M1003 a_3599_383.t4 SN VPB.t76 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VNB a_343_383.t11 a_3368_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1005 VNB a_9985_1004.t8 a_11487_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t61 CLK a_11033_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t13 a_8357_1004.t5 a_8483_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_5227_383.t4 CLK VPB.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_14869_1005.t6 a_3599_383.t8 a_15533_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t52 D a_217_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPB.t86 a_1265_943.t5 a_1905_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t53 D a_5101_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_9985_1004.t4 a_10111_383.t7 VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPB.t26 a_5101_1004.t5 a_6789_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_15533_1005.t1 a_8483_383.t7 a_15044_181.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_6789_1004.t4 a_6149_943.t6 VPB.t38 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t83 a_11033_943.t6 a_11673_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_3599_383.t5 a_1265_943.t6 VPB.t90 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_13241_1004.t1 a_10111_383.t9 VPB.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VNB D a_9880_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1905_1004.t1 a_217_1004.t6 VPB.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t7 a_11673_1004.t7 a_11033_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_14869_1005.t4 a_13367_383.t7 a_15533_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPB.t95 a_343_383.t7 a_217_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPB.t48 a_5227_383.t7 a_5101_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_11673_1004.t5 a_11033_943.t7 VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPB.t23 a_217_1004.t7 a_343_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPB.t0 a_15044_181.t7 a_16835_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB.t31 a_13241_1004.t6 a_13367_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_3473_1004.t3 a_3599_383.t10 VPB.t82 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_10111_383.t3 CLK VPB.t60 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 VNB a_217_1004.t10 a_757_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_5227_383.t3 a_6149_943.t7 VPB.t41 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPB.t28 a_11033_943.t9 a_10111_383.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_13241_1004.t4 a_13367_383.t8 VPB.t94 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPB.t46 a_5227_383.t9 a_8357_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VNB a_1905_1004.t7 a_2702_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_6149_943.t3 CLK VPB.t65 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_14869_1005.t1 a_13367_383.t10 VPB.t44 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 VNB a_10111_383.t10 a_13136_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPB.t42 a_6149_943.t8 a_8483_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_13367_383.t2 a_13241_1004.t7 VPB.t49 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 VNB a_5227_383.t8 a_8252_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1044 VNB a_8357_1004.t7 a_8897_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPB.t21 a_8483_383.t8 a_14869_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPB.t63 CLK a_343_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_3473_1004.t1 a_343_383.t9 VPB.t57 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 VPB.t20 a_1905_1004.t8 a_1265_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_8483_383.t6 SN VPB.t72 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 VPB.t79 SN a_13367_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_10111_383.t0 a_9985_1004.t5 VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 a_15533_1005.t7 a_13367_383.t11 a_14869_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 VPB.t8 a_10111_383.t11 a_9985_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 VNB a_13367_383.t9 a_14764_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1055 VPB.t70 SN a_11673_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_6149_943.t0 a_6789_1004.t7 VPB.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 VPB.t56 a_3473_1004.t6 a_3599_383.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 VPB.t19 a_1265_943.t8 a_3599_383.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 VNB a_217_1004.t5 a_1719_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1060 VPB.t85 a_1265_943.t9 a_343_383.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 a_8483_383.t0 a_8357_1004.t6 VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 VPB.t32 a_11033_943.t10 a_13367_383.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 VPB.t91 a_5101_1004.t8 a_5227_383.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_8483_383.t2 a_6149_943.t9 VPB.t39 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 a_15533_1005.t4 a_3599_383.t13 a_14869_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_217_1004.t1 D VPB.t54 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1067 VPB.t50 D a_9985_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_1905_1004.t5 a_1265_943.t10 VPB.t89 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_6789_1004.t0 a_5101_1004.t9 VPB.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 VPB.t2 a_9985_1004.t7 a_11673_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_15044_181.t2 a_8483_383.t10 a_15533_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 VPB.t74 SN a_3599_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 VPB.t78 SN a_6789_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 VNB a_6789_1004.t8 a_7586_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1075 VNB a_3599_383.t12 a_16096_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1076 VNB D a_4996_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1077 a_11033_943.t0 a_11673_1004.t8 VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 VNB a_13241_1004.t5 a_13781_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1079 a_1905_1004.t3 SN VPB.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_5101_1004.t1 a_5227_383.t10 VPB.t47 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 a_217_1004.t0 a_343_383.t10 VPB.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 VNB a_5101_1004.t6 a_5641_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_6789_1004.t5 SN VPB.t77 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_16835_182.t0 a_15044_181.t9 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_15044_181.t5 a_3599_383.t14 a_15533_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 VPB.t25 a_9985_1004.t9 a_10111_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 VPB.t10 a_8483_383.t12 a_8357_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_343_383.t0 a_217_1004.t8 VPB.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 VPB.t37 a_6149_943.t11 a_6789_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 VPB.t9 a_10111_383.t12 a_13241_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 a_10111_383.t5 a_11033_943.t11 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 a_8357_1004.t3 a_5227_383.t11 VPB.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 VPB.t14 a_217_1004.t9 a_1905_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 VPB.t33 a_6789_1004.t9 a_6149_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 a_11033_943.t3 CLK VPB.t58 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 a_5101_1004.t3 D VPB.t51 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_343_383.t2 CLK VPB.t69 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_14869_1005.t2 a_8483_383.t13 VPB.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 VNB a_5101_1004.t7 a_6603_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_9985_1004.t0 D VPB.t55 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 a_13367_383.t0 SN VPB.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_1265_943.t4 a_1905_1004.t9 VPB.t87 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 VPB.t88 a_3599_383.t15 a_3473_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 VNB a_3473_1004.t5 a_4013_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1105 VPB.t59 CLK a_10111_383.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 a_11673_1004.t2 SN VPB.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 VPB.t68 CLK a_1265_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 VPB.t40 a_6149_943.t12 a_5227_383.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 VPB.t93 a_13367_383.t14 a_13241_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 VNB a_11673_1004.t9 a_12470_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1111 a_8357_1004.t2 a_8483_383.t14 VPB.t43 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1112 a_3599_383.t6 a_3473_1004.t7 VPB.t92 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 VPB.t64 CLK a_6149_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1114 VPB.t35 a_13367_383.t15 a_14869_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 VNB a_9985_1004.t6 a_10525_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1116 VNB a_13367_383.t13 a_15430_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_343_383.t5 a_1265_943.t13 VPB.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 VPB.t36 a_343_383.t12 a_3473_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_5227_383.t0 a_5101_1004.t10 VPB.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 VPB.t80 SN a_8483_383.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 a_13367_383.t5 a_11033_943.t13 VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 a_1265_943.t2 CLK VPB.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 VPB.t81 SN a_1905_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1124 a_11673_1004.t0 a_9985_1004.t10 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB D 0.24fF
C1 VPB CLK 3.26fF
C2 VPB SN 0.30fF
C3 D CLK 1.75fF
C4 D SN 3.39fF
C5 CLK SN 0.41fF
R0 a_6149_943.n6 a_6149_943.t6 454.685
R1 a_6149_943.n8 a_6149_943.t7 454.685
R2 a_6149_943.n4 a_6149_943.t9 454.685
R3 a_6149_943.n6 a_6149_943.t11 428.979
R4 a_6149_943.n8 a_6149_943.t12 428.979
R5 a_6149_943.n4 a_6149_943.t8 428.979
R6 a_6149_943.n7 a_6149_943.t5 248.006
R7 a_6149_943.n9 a_6149_943.t13 248.006
R8 a_6149_943.n5 a_6149_943.t10 248.006
R9 a_6149_943.n14 a_6149_943.n12 220.639
R10 a_6149_943.n12 a_6149_943.n3 135.994
R11 a_6149_943.n7 a_6149_943.n6 81.941
R12 a_6149_943.n9 a_6149_943.n8 81.941
R13 a_6149_943.n5 a_6149_943.n4 81.941
R14 a_6149_943.n11 a_6149_943.n5 81.396
R15 a_6149_943.n10 a_6149_943.n9 79.491
R16 a_6149_943.n3 a_6149_943.n2 76.002
R17 a_6149_943.n10 a_6149_943.n7 76
R18 a_6149_943.n12 a_6149_943.n11 76
R19 a_6149_943.n14 a_6149_943.n13 30
R20 a_6149_943.n15 a_6149_943.n0 24.383
R21 a_6149_943.n15 a_6149_943.n14 23.684
R22 a_6149_943.n1 a_6149_943.t2 14.282
R23 a_6149_943.n1 a_6149_943.t3 14.282
R24 a_6149_943.n2 a_6149_943.t1 14.282
R25 a_6149_943.n2 a_6149_943.t0 14.282
R26 a_6149_943.n3 a_6149_943.n1 12.85
R27 a_6149_943.n11 a_6149_943.n10 2.947
R28 a_6884_182.n13 a_6884_182.n6 82.852
R29 a_6884_182.t0 a_6884_182.n1 46.91
R30 a_6884_182.n10 a_6884_182.n8 34.805
R31 a_6884_182.n10 a_6884_182.n9 32.622
R32 a_6884_182.t0 a_6884_182.n13 32.417
R33 a_6884_182.n6 a_6884_182.n5 27.2
R34 a_6884_182.n4 a_6884_182.n3 23.498
R35 a_6884_182.n6 a_6884_182.n4 22.4
R36 a_6884_182.n12 a_6884_182.n10 19.017
R37 a_6884_182.n1 a_6884_182.n0 17.006
R38 a_6884_182.t0 a_6884_182.n2 8.137
R39 a_6884_182.n8 a_6884_182.n7 7.5
R40 a_6884_182.n12 a_6884_182.n11 7.5
R41 a_6884_182.n13 a_6884_182.n12 1.435
R42 a_6789_1004.n5 a_6789_1004.t9 480.392
R43 a_6789_1004.n5 a_6789_1004.t7 403.272
R44 a_6789_1004.n7 a_6789_1004.n4 233.952
R45 a_6789_1004.n6 a_6789_1004.t8 213.869
R46 a_6789_1004.n6 a_6789_1004.n5 161.6
R47 a_6789_1004.n7 a_6789_1004.n6 153.315
R48 a_6789_1004.n9 a_6789_1004.n7 150.014
R49 a_6789_1004.n3 a_6789_1004.n2 79.232
R50 a_6789_1004.n4 a_6789_1004.n3 63.152
R51 a_6789_1004.n4 a_6789_1004.n0 16.08
R52 a_6789_1004.n3 a_6789_1004.n1 16.08
R53 a_6789_1004.n9 a_6789_1004.n8 15.218
R54 a_6789_1004.n0 a_6789_1004.t3 14.282
R55 a_6789_1004.n0 a_6789_1004.t4 14.282
R56 a_6789_1004.n1 a_6789_1004.t6 14.282
R57 a_6789_1004.n1 a_6789_1004.t5 14.282
R58 a_6789_1004.n2 a_6789_1004.t1 14.282
R59 a_6789_1004.n2 a_6789_1004.t0 14.282
R60 a_6789_1004.n10 a_6789_1004.n9 12.014
R61 a_5227_383.n6 a_5227_383.t9 480.392
R62 a_5227_383.n8 a_5227_383.t7 472.359
R63 a_5227_383.n6 a_5227_383.t11 403.272
R64 a_5227_383.n8 a_5227_383.t10 384.527
R65 a_5227_383.n7 a_5227_383.t8 320.08
R66 a_5227_383.n9 a_5227_383.t12 277.772
R67 a_5227_383.n13 a_5227_383.n11 249.364
R68 a_5227_383.n11 a_5227_383.n5 127.401
R69 a_5227_383.n10 a_5227_383.n7 83.304
R70 a_5227_383.n10 a_5227_383.n9 80.032
R71 a_5227_383.n4 a_5227_383.n3 79.232
R72 a_5227_383.n11 a_5227_383.n10 76
R73 a_5227_383.n9 a_5227_383.n8 67.001
R74 a_5227_383.n5 a_5227_383.n4 63.152
R75 a_5227_383.n7 a_5227_383.n6 55.388
R76 a_5227_383.n13 a_5227_383.n12 30
R77 a_5227_383.n14 a_5227_383.n0 24.383
R78 a_5227_383.n14 a_5227_383.n13 23.684
R79 a_5227_383.n5 a_5227_383.n1 16.08
R80 a_5227_383.n4 a_5227_383.n2 16.08
R81 a_5227_383.n1 a_5227_383.t2 14.282
R82 a_5227_383.n1 a_5227_383.t3 14.282
R83 a_5227_383.n2 a_5227_383.t5 14.282
R84 a_5227_383.n2 a_5227_383.t4 14.282
R85 a_5227_383.n3 a_5227_383.t6 14.282
R86 a_5227_383.n3 a_5227_383.t0 14.282
R87 VPB VPB.n1549 126.832
R88 VPB.n49 VPB.n47 94.117
R89 VPB.n1485 VPB.n1483 94.117
R90 VPB.n1402 VPB.n1400 94.117
R91 VPB.n1339 VPB.n1337 94.117
R92 VPB.n1276 VPB.n1274 94.117
R93 VPB.n1193 VPB.n1191 94.117
R94 VPB.n1130 VPB.n1128 94.117
R95 VPB.n1047 VPB.n1045 94.117
R96 VPB.n964 VPB.n962 94.117
R97 VPB.n901 VPB.n899 94.117
R98 VPB.n134 VPB.n132 94.117
R99 VPB.n819 VPB.n817 94.117
R100 VPB.n756 VPB.n754 94.117
R101 VPB.n673 VPB.n671 94.117
R102 VPB.n590 VPB.n588 94.117
R103 VPB.n527 VPB.n525 94.117
R104 VPB.n464 VPB.n462 94.117
R105 VPB.n381 VPB.n379 94.117
R106 VPB.n318 VPB.n316 94.117
R107 VPB.n263 VPB.n261 94.117
R108 VPB.n208 VPB.n206 91.036
R109 VPB.n394 VPB.n393 80.104
R110 VPB.n603 VPB.n602 80.104
R111 VPB.n686 VPB.n685 80.104
R112 VPB.n832 VPB.n831 80.104
R113 VPB.n977 VPB.n976 80.104
R114 VPB.n1060 VPB.n1059 80.104
R115 VPB.n1206 VPB.n1205 80.104
R116 VPB.n1415 VPB.n1414 80.104
R117 VPB.n1498 VPB.n1497 80.104
R118 VPB.n169 VPB.n163 76.136
R119 VPB.n169 VPB.n168 76
R120 VPB.n173 VPB.n172 76
R121 VPB.n179 VPB.n178 76
R122 VPB.n183 VPB.n182 76
R123 VPB.n210 VPB.n209 76
R124 VPB.n214 VPB.n213 76
R125 VPB.n218 VPB.n217 76
R126 VPB.n222 VPB.n221 76
R127 VPB.n226 VPB.n225 76
R128 VPB.n230 VPB.n229 76
R129 VPB.n234 VPB.n233 76
R130 VPB.n238 VPB.n237 76
R131 VPB.n265 VPB.n264 76
R132 VPB.n269 VPB.n268 76
R133 VPB.n273 VPB.n272 76
R134 VPB.n277 VPB.n276 76
R135 VPB.n281 VPB.n280 76
R136 VPB.n285 VPB.n284 76
R137 VPB.n289 VPB.n288 76
R138 VPB.n293 VPB.n292 76
R139 VPB.n320 VPB.n319 76
R140 VPB.n325 VPB.n324 76
R141 VPB.n330 VPB.n329 76
R142 VPB.n337 VPB.n336 76
R143 VPB.n342 VPB.n341 76
R144 VPB.n347 VPB.n346 76
R145 VPB.n352 VPB.n351 76
R146 VPB.n356 VPB.n355 76
R147 VPB.n383 VPB.n382 76
R148 VPB.n387 VPB.n386 76
R149 VPB.n392 VPB.n391 76
R150 VPB.n397 VPB.n396 76
R151 VPB.n404 VPB.n403 76
R152 VPB.n409 VPB.n408 76
R153 VPB.n414 VPB.n413 76
R154 VPB.n421 VPB.n420 76
R155 VPB.n426 VPB.n425 76
R156 VPB.n431 VPB.n430 76
R157 VPB.n435 VPB.n434 76
R158 VPB.n439 VPB.n438 76
R159 VPB.n466 VPB.n465 76
R160 VPB.n471 VPB.n470 76
R161 VPB.n476 VPB.n475 76
R162 VPB.n483 VPB.n482 76
R163 VPB.n488 VPB.n487 76
R164 VPB.n493 VPB.n492 76
R165 VPB.n498 VPB.n497 76
R166 VPB.n502 VPB.n501 76
R167 VPB.n529 VPB.n528 76
R168 VPB.n534 VPB.n533 76
R169 VPB.n539 VPB.n538 76
R170 VPB.n546 VPB.n545 76
R171 VPB.n551 VPB.n550 76
R172 VPB.n556 VPB.n555 76
R173 VPB.n561 VPB.n560 76
R174 VPB.n565 VPB.n564 76
R175 VPB.n592 VPB.n591 76
R176 VPB.n596 VPB.n595 76
R177 VPB.n601 VPB.n600 76
R178 VPB.n606 VPB.n605 76
R179 VPB.n613 VPB.n612 76
R180 VPB.n618 VPB.n617 76
R181 VPB.n623 VPB.n622 76
R182 VPB.n630 VPB.n629 76
R183 VPB.n635 VPB.n634 76
R184 VPB.n640 VPB.n639 76
R185 VPB.n644 VPB.n643 76
R186 VPB.n648 VPB.n647 76
R187 VPB.n675 VPB.n674 76
R188 VPB.n679 VPB.n678 76
R189 VPB.n684 VPB.n683 76
R190 VPB.n689 VPB.n688 76
R191 VPB.n696 VPB.n695 76
R192 VPB.n701 VPB.n700 76
R193 VPB.n706 VPB.n705 76
R194 VPB.n713 VPB.n712 76
R195 VPB.n718 VPB.n717 76
R196 VPB.n723 VPB.n722 76
R197 VPB.n727 VPB.n726 76
R198 VPB.n731 VPB.n730 76
R199 VPB.n758 VPB.n757 76
R200 VPB.n763 VPB.n762 76
R201 VPB.n768 VPB.n767 76
R202 VPB.n775 VPB.n774 76
R203 VPB.n780 VPB.n779 76
R204 VPB.n785 VPB.n784 76
R205 VPB.n790 VPB.n789 76
R206 VPB.n794 VPB.n793 76
R207 VPB.n821 VPB.n820 76
R208 VPB.n825 VPB.n824 76
R209 VPB.n830 VPB.n829 76
R210 VPB.n835 VPB.n834 76
R211 VPB.n850 VPB.n846 76
R212 VPB.n857 VPB.n856 76
R213 VPB.n862 VPB.n861 76
R214 VPB.n867 VPB.n866 76
R215 VPB.n872 VPB.n871 76
R216 VPB.n876 VPB.n875 76
R217 VPB.n903 VPB.n902 76
R218 VPB.n908 VPB.n907 76
R219 VPB.n913 VPB.n912 76
R220 VPB.n920 VPB.n919 76
R221 VPB.n925 VPB.n924 76
R222 VPB.n930 VPB.n929 76
R223 VPB.n935 VPB.n934 76
R224 VPB.n939 VPB.n938 76
R225 VPB.n966 VPB.n965 76
R226 VPB.n970 VPB.n969 76
R227 VPB.n975 VPB.n974 76
R228 VPB.n980 VPB.n979 76
R229 VPB.n987 VPB.n986 76
R230 VPB.n992 VPB.n991 76
R231 VPB.n997 VPB.n996 76
R232 VPB.n1004 VPB.n1003 76
R233 VPB.n1009 VPB.n1008 76
R234 VPB.n1014 VPB.n1013 76
R235 VPB.n1018 VPB.n1017 76
R236 VPB.n1022 VPB.n1021 76
R237 VPB.n1049 VPB.n1048 76
R238 VPB.n1053 VPB.n1052 76
R239 VPB.n1058 VPB.n1057 76
R240 VPB.n1063 VPB.n1062 76
R241 VPB.n1070 VPB.n1069 76
R242 VPB.n1075 VPB.n1074 76
R243 VPB.n1080 VPB.n1079 76
R244 VPB.n1087 VPB.n1086 76
R245 VPB.n1092 VPB.n1091 76
R246 VPB.n1097 VPB.n1096 76
R247 VPB.n1101 VPB.n1100 76
R248 VPB.n1105 VPB.n1104 76
R249 VPB.n1132 VPB.n1131 76
R250 VPB.n1137 VPB.n1136 76
R251 VPB.n1142 VPB.n1141 76
R252 VPB.n1149 VPB.n1148 76
R253 VPB.n1154 VPB.n1153 76
R254 VPB.n1159 VPB.n1158 76
R255 VPB.n1164 VPB.n1163 76
R256 VPB.n1168 VPB.n1167 76
R257 VPB.n1195 VPB.n1194 76
R258 VPB.n1199 VPB.n1198 76
R259 VPB.n1204 VPB.n1203 76
R260 VPB.n1209 VPB.n1208 76
R261 VPB.n1216 VPB.n1215 76
R262 VPB.n1221 VPB.n1220 76
R263 VPB.n1226 VPB.n1225 76
R264 VPB.n1233 VPB.n1232 76
R265 VPB.n1238 VPB.n1237 76
R266 VPB.n1243 VPB.n1242 76
R267 VPB.n1247 VPB.n1246 76
R268 VPB.n1251 VPB.n1250 76
R269 VPB.n1278 VPB.n1277 76
R270 VPB.n1283 VPB.n1282 76
R271 VPB.n1288 VPB.n1287 76
R272 VPB.n1295 VPB.n1294 76
R273 VPB.n1300 VPB.n1299 76
R274 VPB.n1305 VPB.n1304 76
R275 VPB.n1310 VPB.n1309 76
R276 VPB.n1314 VPB.n1313 76
R277 VPB.n1341 VPB.n1340 76
R278 VPB.n1346 VPB.n1345 76
R279 VPB.n1351 VPB.n1350 76
R280 VPB.n1358 VPB.n1357 76
R281 VPB.n1363 VPB.n1362 76
R282 VPB.n1368 VPB.n1367 76
R283 VPB.n1373 VPB.n1372 76
R284 VPB.n1377 VPB.n1376 76
R285 VPB.n1404 VPB.n1403 76
R286 VPB.n1408 VPB.n1407 76
R287 VPB.n1413 VPB.n1412 76
R288 VPB.n1418 VPB.n1417 76
R289 VPB.n1425 VPB.n1424 76
R290 VPB.n1430 VPB.n1429 76
R291 VPB.n1435 VPB.n1434 76
R292 VPB.n1442 VPB.n1441 76
R293 VPB.n1447 VPB.n1446 76
R294 VPB.n1452 VPB.n1451 76
R295 VPB.n1456 VPB.n1455 76
R296 VPB.n1460 VPB.n1459 76
R297 VPB.n1487 VPB.n1486 76
R298 VPB.n1491 VPB.n1490 76
R299 VPB.n1496 VPB.n1495 76
R300 VPB.n1501 VPB.n1500 76
R301 VPB.n1508 VPB.n1507 76
R302 VPB.n1513 VPB.n1512 76
R303 VPB.n1518 VPB.n1517 76
R304 VPB.n1525 VPB.n1524 76
R305 VPB.n1530 VPB.n1529 76
R306 VPB.n1542 VPB.n1541 76
R307 VPB.n423 VPB.n422 75.654
R308 VPB.n632 VPB.n631 75.654
R309 VPB.n715 VPB.n714 75.654
R310 VPB.n118 VPB.n117 75.654
R311 VPB.n1006 VPB.n1005 75.654
R312 VPB.n1089 VPB.n1088 75.654
R313 VPB.n1235 VPB.n1234 75.654
R314 VPB.n1444 VPB.n1443 75.654
R315 VPB.n1527 VPB.n1526 75.654
R316 VPB.n176 VPB.n175 68.979
R317 VPB.n166 VPB.n165 64.528
R318 VPB.n21 VPB.n20 61.764
R319 VPB.n1467 VPB.n1466 61.764
R320 VPB.n1384 VPB.n1383 61.764
R321 VPB.n1321 VPB.n1320 61.764
R322 VPB.n1258 VPB.n1257 61.764
R323 VPB.n1175 VPB.n1174 61.764
R324 VPB.n1112 VPB.n1111 61.764
R325 VPB.n1029 VPB.n1028 61.764
R326 VPB.n946 VPB.n945 61.764
R327 VPB.n883 VPB.n882 61.764
R328 VPB.n82 VPB.n81 61.764
R329 VPB.n801 VPB.n800 61.764
R330 VPB.n738 VPB.n737 61.764
R331 VPB.n655 VPB.n654 61.764
R332 VPB.n572 VPB.n571 61.764
R333 VPB.n509 VPB.n508 61.764
R334 VPB.n446 VPB.n445 61.764
R335 VPB.n363 VPB.n362 61.764
R336 VPB.n300 VPB.n299 61.764
R337 VPB.n245 VPB.n244 61.764
R338 VPB.n190 VPB.n189 61.764
R339 VPB.n348 VPB.t44 55.465
R340 VPB.n321 VPB.t21 55.465
R341 VPB.n72 VPB.t54 55.106
R342 VPB.n39 VPB.t84 55.106
R343 VPB.n1448 VPB.t29 55.106
R344 VPB.n1369 VPB.t87 55.106
R345 VPB.n1306 VPB.t57 55.106
R346 VPB.n1239 VPB.t92 55.106
R347 VPB.n1160 VPB.t51 55.106
R348 VPB.n1093 VPB.t16 55.106
R349 VPB.n1010 VPB.t24 55.106
R350 VPB.n931 VPB.t34 55.106
R351 VPB.n868 VPB.t45 55.106
R352 VPB.n124 VPB.t11 55.106
R353 VPB.n786 VPB.t55 55.106
R354 VPB.n719 VPB.t3 55.106
R355 VPB.n636 VPB.t1 55.106
R356 VPB.n557 VPB.t4 55.106
R357 VPB.n494 VPB.t15 55.106
R358 VPB.n427 VPB.t49 55.106
R359 VPB.n174 VPB.t6 55.106
R360 VPB.n164 VPB.t0 55.106
R361 VPB.n54 VPB.t95 55.106
R362 VPB.n1492 VPB.t85 55.106
R363 VPB.n1409 VPB.t86 55.106
R364 VPB.n1342 VPB.t68 55.106
R365 VPB.n1279 VPB.t88 55.106
R366 VPB.n1200 VPB.t19 55.106
R367 VPB.n1133 VPB.t48 55.106
R368 VPB.n1054 VPB.t40 55.106
R369 VPB.n971 VPB.t37 55.106
R370 VPB.n904 VPB.t64 55.106
R371 VPB.n139 VPB.t10 55.106
R372 VPB.n826 VPB.t42 55.106
R373 VPB.n759 VPB.t8 55.106
R374 VPB.n680 VPB.t28 55.106
R375 VPB.n597 VPB.t83 55.106
R376 VPB.n530 VPB.t61 55.106
R377 VPB.n467 VPB.t93 55.106
R378 VPB.n388 VPB.t32 55.106
R379 VPB.n327 VPB.n326 48.952
R380 VPB.n401 VPB.n400 48.952
R381 VPB.n473 VPB.n472 48.952
R382 VPB.n536 VPB.n535 48.952
R383 VPB.n610 VPB.n609 48.952
R384 VPB.n693 VPB.n692 48.952
R385 VPB.n765 VPB.n764 48.952
R386 VPB.n100 VPB.n99 48.952
R387 VPB.n848 VPB.n847 48.952
R388 VPB.n910 VPB.n909 48.952
R389 VPB.n984 VPB.n983 48.952
R390 VPB.n1067 VPB.n1066 48.952
R391 VPB.n1139 VPB.n1138 48.952
R392 VPB.n1213 VPB.n1212 48.952
R393 VPB.n1285 VPB.n1284 48.952
R394 VPB.n1348 VPB.n1347 48.952
R395 VPB.n1422 VPB.n1421 48.952
R396 VPB.n1505 VPB.n1504 48.952
R397 VPB.n56 VPB.n55 48.952
R398 VPB.n344 VPB.n343 44.502
R399 VPB.n418 VPB.n417 44.502
R400 VPB.n490 VPB.n489 44.502
R401 VPB.n553 VPB.n552 44.502
R402 VPB.n627 VPB.n626 44.502
R403 VPB.n710 VPB.n709 44.502
R404 VPB.n782 VPB.n781 44.502
R405 VPB.n114 VPB.n113 44.502
R406 VPB.n864 VPB.n863 44.502
R407 VPB.n927 VPB.n926 44.502
R408 VPB.n1001 VPB.n1000 44.502
R409 VPB.n1084 VPB.n1083 44.502
R410 VPB.n1156 VPB.n1155 44.502
R411 VPB.n1230 VPB.n1229 44.502
R412 VPB.n1302 VPB.n1301 44.502
R413 VPB.n1365 VPB.n1364 44.502
R414 VPB.n1439 VPB.n1438 44.502
R415 VPB.n1522 VPB.n1521 44.502
R416 VPB.n69 VPB.n68 44.502
R417 VPB.n332 VPB.n331 41.183
R418 VPB.n63 VPB.n14 40.824
R419 VPB.n1520 VPB.n1519 40.824
R420 VPB.n1503 VPB.n1502 40.824
R421 VPB.n1437 VPB.n1436 40.824
R422 VPB.n1420 VPB.n1419 40.824
R423 VPB.n1353 VPB.n1352 40.824
R424 VPB.n1290 VPB.n1289 40.824
R425 VPB.n1228 VPB.n1227 40.824
R426 VPB.n1211 VPB.n1210 40.824
R427 VPB.n1144 VPB.n1143 40.824
R428 VPB.n1082 VPB.n1081 40.824
R429 VPB.n1065 VPB.n1064 40.824
R430 VPB.n999 VPB.n998 40.824
R431 VPB.n982 VPB.n981 40.824
R432 VPB.n915 VPB.n914 40.824
R433 VPB.n852 VPB.n851 40.824
R434 VPB.n112 VPB.n97 40.824
R435 VPB.n103 VPB.n98 40.824
R436 VPB.n770 VPB.n769 40.824
R437 VPB.n708 VPB.n707 40.824
R438 VPB.n691 VPB.n690 40.824
R439 VPB.n625 VPB.n624 40.824
R440 VPB.n608 VPB.n607 40.824
R441 VPB.n541 VPB.n540 40.824
R442 VPB.n478 VPB.n477 40.824
R443 VPB.n416 VPB.n415 40.824
R444 VPB.n399 VPB.n398 40.824
R445 VPB.n1546 VPB.n1542 20.452
R446 VPB.n163 VPB.n160 20.452
R447 VPB.n334 VPB.n333 17.801
R448 VPB.n406 VPB.n405 17.801
R449 VPB.n480 VPB.n479 17.801
R450 VPB.n543 VPB.n542 17.801
R451 VPB.n615 VPB.n614 17.801
R452 VPB.n698 VPB.n697 17.801
R453 VPB.n772 VPB.n771 17.801
R454 VPB.n105 VPB.n104 17.801
R455 VPB.n854 VPB.n853 17.801
R456 VPB.n917 VPB.n916 17.801
R457 VPB.n989 VPB.n988 17.801
R458 VPB.n1072 VPB.n1071 17.801
R459 VPB.n1146 VPB.n1145 17.801
R460 VPB.n1218 VPB.n1217 17.801
R461 VPB.n1292 VPB.n1291 17.801
R462 VPB.n1355 VPB.n1354 17.801
R463 VPB.n1427 VPB.n1426 17.801
R464 VPB.n1510 VPB.n1509 17.801
R465 VPB.n60 VPB.n59 17.801
R466 VPB.n14 VPB.t30 14.282
R467 VPB.n14 VPB.t52 14.282
R468 VPB.n1519 VPB.t69 14.282
R469 VPB.n1519 VPB.t23 14.282
R470 VPB.n1502 VPB.t22 14.282
R471 VPB.n1502 VPB.t63 14.282
R472 VPB.n1436 VPB.t73 14.282
R473 VPB.n1436 VPB.t14 14.282
R474 VPB.n1419 VPB.t89 14.282
R475 VPB.n1419 VPB.t81 14.282
R476 VPB.n1352 VPB.t62 14.282
R477 VPB.n1352 VPB.t20 14.282
R478 VPB.n1289 VPB.t82 14.282
R479 VPB.n1289 VPB.t36 14.282
R480 VPB.n1227 VPB.t76 14.282
R481 VPB.n1227 VPB.t56 14.282
R482 VPB.n1210 VPB.t90 14.282
R483 VPB.n1210 VPB.t74 14.282
R484 VPB.n1143 VPB.t47 14.282
R485 VPB.n1143 VPB.t53 14.282
R486 VPB.n1081 VPB.t66 14.282
R487 VPB.n1081 VPB.t91 14.282
R488 VPB.n1064 VPB.t41 14.282
R489 VPB.n1064 VPB.t67 14.282
R490 VPB.n998 VPB.t77 14.282
R491 VPB.n998 VPB.t26 14.282
R492 VPB.n981 VPB.t38 14.282
R493 VPB.n981 VPB.t78 14.282
R494 VPB.n914 VPB.t65 14.282
R495 VPB.n914 VPB.t33 14.282
R496 VPB.n851 VPB.t43 14.282
R497 VPB.n851 VPB.t46 14.282
R498 VPB.n97 VPB.t72 14.282
R499 VPB.n97 VPB.t13 14.282
R500 VPB.n98 VPB.t39 14.282
R501 VPB.n98 VPB.t80 14.282
R502 VPB.n769 VPB.t17 14.282
R503 VPB.n769 VPB.t50 14.282
R504 VPB.n707 VPB.t60 14.282
R505 VPB.n707 VPB.t25 14.282
R506 VPB.n690 VPB.t12 14.282
R507 VPB.n690 VPB.t59 14.282
R508 VPB.n624 VPB.t71 14.282
R509 VPB.n624 VPB.t2 14.282
R510 VPB.n607 VPB.t5 14.282
R511 VPB.n607 VPB.t70 14.282
R512 VPB.n540 VPB.t58 14.282
R513 VPB.n540 VPB.t7 14.282
R514 VPB.n477 VPB.t94 14.282
R515 VPB.n477 VPB.t9 14.282
R516 VPB.n415 VPB.t75 14.282
R517 VPB.n415 VPB.t31 14.282
R518 VPB.n398 VPB.t18 14.282
R519 VPB.n398 VPB.t79 14.282
R520 VPB.n331 VPB.t27 14.282
R521 VPB.n331 VPB.t35 14.282
R522 VPB.n163 VPB.n162 13.653
R523 VPB.n162 VPB.n161 13.653
R524 VPB.n168 VPB.n167 13.653
R525 VPB.n167 VPB.n166 13.653
R526 VPB.n172 VPB.n171 13.653
R527 VPB.n171 VPB.n170 13.653
R528 VPB.n178 VPB.n177 13.653
R529 VPB.n177 VPB.n176 13.653
R530 VPB.n182 VPB.n181 13.653
R531 VPB.n181 VPB.n180 13.653
R532 VPB.n209 VPB.n208 13.653
R533 VPB.n208 VPB.n207 13.653
R534 VPB.n213 VPB.n212 13.653
R535 VPB.n212 VPB.n211 13.653
R536 VPB.n217 VPB.n216 13.653
R537 VPB.n216 VPB.n215 13.653
R538 VPB.n221 VPB.n220 13.653
R539 VPB.n220 VPB.n219 13.653
R540 VPB.n225 VPB.n224 13.653
R541 VPB.n224 VPB.n223 13.653
R542 VPB.n229 VPB.n228 13.653
R543 VPB.n228 VPB.n227 13.653
R544 VPB.n233 VPB.n232 13.653
R545 VPB.n232 VPB.n231 13.653
R546 VPB.n237 VPB.n236 13.653
R547 VPB.n236 VPB.n235 13.653
R548 VPB.n264 VPB.n263 13.653
R549 VPB.n263 VPB.n262 13.653
R550 VPB.n268 VPB.n267 13.653
R551 VPB.n267 VPB.n266 13.653
R552 VPB.n272 VPB.n271 13.653
R553 VPB.n271 VPB.n270 13.653
R554 VPB.n276 VPB.n275 13.653
R555 VPB.n275 VPB.n274 13.653
R556 VPB.n280 VPB.n279 13.653
R557 VPB.n279 VPB.n278 13.653
R558 VPB.n284 VPB.n283 13.653
R559 VPB.n283 VPB.n282 13.653
R560 VPB.n288 VPB.n287 13.653
R561 VPB.n287 VPB.n286 13.653
R562 VPB.n292 VPB.n291 13.653
R563 VPB.n291 VPB.n290 13.653
R564 VPB.n319 VPB.n318 13.653
R565 VPB.n318 VPB.n317 13.653
R566 VPB.n324 VPB.n323 13.653
R567 VPB.n323 VPB.n322 13.653
R568 VPB.n329 VPB.n328 13.653
R569 VPB.n328 VPB.n327 13.653
R570 VPB.n336 VPB.n335 13.653
R571 VPB.n335 VPB.n334 13.653
R572 VPB.n341 VPB.n340 13.653
R573 VPB.n340 VPB.n339 13.653
R574 VPB.n346 VPB.n345 13.653
R575 VPB.n345 VPB.n344 13.653
R576 VPB.n351 VPB.n350 13.653
R577 VPB.n350 VPB.n349 13.653
R578 VPB.n355 VPB.n354 13.653
R579 VPB.n354 VPB.n353 13.653
R580 VPB.n382 VPB.n381 13.653
R581 VPB.n381 VPB.n380 13.653
R582 VPB.n386 VPB.n385 13.653
R583 VPB.n385 VPB.n384 13.653
R584 VPB.n391 VPB.n390 13.653
R585 VPB.n390 VPB.n389 13.653
R586 VPB.n396 VPB.n395 13.653
R587 VPB.n395 VPB.n394 13.653
R588 VPB.n403 VPB.n402 13.653
R589 VPB.n402 VPB.n401 13.653
R590 VPB.n408 VPB.n407 13.653
R591 VPB.n407 VPB.n406 13.653
R592 VPB.n413 VPB.n412 13.653
R593 VPB.n412 VPB.n411 13.653
R594 VPB.n420 VPB.n419 13.653
R595 VPB.n419 VPB.n418 13.653
R596 VPB.n425 VPB.n424 13.653
R597 VPB.n424 VPB.n423 13.653
R598 VPB.n430 VPB.n429 13.653
R599 VPB.n429 VPB.n428 13.653
R600 VPB.n434 VPB.n433 13.653
R601 VPB.n433 VPB.n432 13.653
R602 VPB.n438 VPB.n437 13.653
R603 VPB.n437 VPB.n436 13.653
R604 VPB.n465 VPB.n464 13.653
R605 VPB.n464 VPB.n463 13.653
R606 VPB.n470 VPB.n469 13.653
R607 VPB.n469 VPB.n468 13.653
R608 VPB.n475 VPB.n474 13.653
R609 VPB.n474 VPB.n473 13.653
R610 VPB.n482 VPB.n481 13.653
R611 VPB.n481 VPB.n480 13.653
R612 VPB.n487 VPB.n486 13.653
R613 VPB.n486 VPB.n485 13.653
R614 VPB.n492 VPB.n491 13.653
R615 VPB.n491 VPB.n490 13.653
R616 VPB.n497 VPB.n496 13.653
R617 VPB.n496 VPB.n495 13.653
R618 VPB.n501 VPB.n500 13.653
R619 VPB.n500 VPB.n499 13.653
R620 VPB.n528 VPB.n527 13.653
R621 VPB.n527 VPB.n526 13.653
R622 VPB.n533 VPB.n532 13.653
R623 VPB.n532 VPB.n531 13.653
R624 VPB.n538 VPB.n537 13.653
R625 VPB.n537 VPB.n536 13.653
R626 VPB.n545 VPB.n544 13.653
R627 VPB.n544 VPB.n543 13.653
R628 VPB.n550 VPB.n549 13.653
R629 VPB.n549 VPB.n548 13.653
R630 VPB.n555 VPB.n554 13.653
R631 VPB.n554 VPB.n553 13.653
R632 VPB.n560 VPB.n559 13.653
R633 VPB.n559 VPB.n558 13.653
R634 VPB.n564 VPB.n563 13.653
R635 VPB.n563 VPB.n562 13.653
R636 VPB.n591 VPB.n590 13.653
R637 VPB.n590 VPB.n589 13.653
R638 VPB.n595 VPB.n594 13.653
R639 VPB.n594 VPB.n593 13.653
R640 VPB.n600 VPB.n599 13.653
R641 VPB.n599 VPB.n598 13.653
R642 VPB.n605 VPB.n604 13.653
R643 VPB.n604 VPB.n603 13.653
R644 VPB.n612 VPB.n611 13.653
R645 VPB.n611 VPB.n610 13.653
R646 VPB.n617 VPB.n616 13.653
R647 VPB.n616 VPB.n615 13.653
R648 VPB.n622 VPB.n621 13.653
R649 VPB.n621 VPB.n620 13.653
R650 VPB.n629 VPB.n628 13.653
R651 VPB.n628 VPB.n627 13.653
R652 VPB.n634 VPB.n633 13.653
R653 VPB.n633 VPB.n632 13.653
R654 VPB.n639 VPB.n638 13.653
R655 VPB.n638 VPB.n637 13.653
R656 VPB.n643 VPB.n642 13.653
R657 VPB.n642 VPB.n641 13.653
R658 VPB.n647 VPB.n646 13.653
R659 VPB.n646 VPB.n645 13.653
R660 VPB.n674 VPB.n673 13.653
R661 VPB.n673 VPB.n672 13.653
R662 VPB.n678 VPB.n677 13.653
R663 VPB.n677 VPB.n676 13.653
R664 VPB.n683 VPB.n682 13.653
R665 VPB.n682 VPB.n681 13.653
R666 VPB.n688 VPB.n687 13.653
R667 VPB.n687 VPB.n686 13.653
R668 VPB.n695 VPB.n694 13.653
R669 VPB.n694 VPB.n693 13.653
R670 VPB.n700 VPB.n699 13.653
R671 VPB.n699 VPB.n698 13.653
R672 VPB.n705 VPB.n704 13.653
R673 VPB.n704 VPB.n703 13.653
R674 VPB.n712 VPB.n711 13.653
R675 VPB.n711 VPB.n710 13.653
R676 VPB.n717 VPB.n716 13.653
R677 VPB.n716 VPB.n715 13.653
R678 VPB.n722 VPB.n721 13.653
R679 VPB.n721 VPB.n720 13.653
R680 VPB.n726 VPB.n725 13.653
R681 VPB.n725 VPB.n724 13.653
R682 VPB.n730 VPB.n729 13.653
R683 VPB.n729 VPB.n728 13.653
R684 VPB.n757 VPB.n756 13.653
R685 VPB.n756 VPB.n755 13.653
R686 VPB.n762 VPB.n761 13.653
R687 VPB.n761 VPB.n760 13.653
R688 VPB.n767 VPB.n766 13.653
R689 VPB.n766 VPB.n765 13.653
R690 VPB.n774 VPB.n773 13.653
R691 VPB.n773 VPB.n772 13.653
R692 VPB.n779 VPB.n778 13.653
R693 VPB.n778 VPB.n777 13.653
R694 VPB.n784 VPB.n783 13.653
R695 VPB.n783 VPB.n782 13.653
R696 VPB.n789 VPB.n788 13.653
R697 VPB.n788 VPB.n787 13.653
R698 VPB.n793 VPB.n792 13.653
R699 VPB.n792 VPB.n791 13.653
R700 VPB.n820 VPB.n819 13.653
R701 VPB.n819 VPB.n818 13.653
R702 VPB.n824 VPB.n823 13.653
R703 VPB.n823 VPB.n822 13.653
R704 VPB.n829 VPB.n828 13.653
R705 VPB.n828 VPB.n827 13.653
R706 VPB.n834 VPB.n833 13.653
R707 VPB.n833 VPB.n832 13.653
R708 VPB.n102 VPB.n101 13.653
R709 VPB.n101 VPB.n100 13.653
R710 VPB.n107 VPB.n106 13.653
R711 VPB.n106 VPB.n105 13.653
R712 VPB.n111 VPB.n110 13.653
R713 VPB.n110 VPB.n109 13.653
R714 VPB.n116 VPB.n115 13.653
R715 VPB.n115 VPB.n114 13.653
R716 VPB.n120 VPB.n119 13.653
R717 VPB.n119 VPB.n118 13.653
R718 VPB.n123 VPB.n122 13.653
R719 VPB.n122 VPB.n121 13.653
R720 VPB.n127 VPB.n126 13.653
R721 VPB.n126 VPB.n125 13.653
R722 VPB.n130 VPB.n129 13.653
R723 VPB.n129 VPB.n128 13.653
R724 VPB.n135 VPB.n134 13.653
R725 VPB.n134 VPB.n133 13.653
R726 VPB.n138 VPB.n137 13.653
R727 VPB.n137 VPB.n136 13.653
R728 VPB.n850 VPB.n849 13.653
R729 VPB.n849 VPB.n848 13.653
R730 VPB.n856 VPB.n855 13.653
R731 VPB.n855 VPB.n854 13.653
R732 VPB.n861 VPB.n860 13.653
R733 VPB.n860 VPB.n859 13.653
R734 VPB.n866 VPB.n865 13.653
R735 VPB.n865 VPB.n864 13.653
R736 VPB.n871 VPB.n870 13.653
R737 VPB.n870 VPB.n869 13.653
R738 VPB.n875 VPB.n874 13.653
R739 VPB.n874 VPB.n873 13.653
R740 VPB.n902 VPB.n901 13.653
R741 VPB.n901 VPB.n900 13.653
R742 VPB.n907 VPB.n906 13.653
R743 VPB.n906 VPB.n905 13.653
R744 VPB.n912 VPB.n911 13.653
R745 VPB.n911 VPB.n910 13.653
R746 VPB.n919 VPB.n918 13.653
R747 VPB.n918 VPB.n917 13.653
R748 VPB.n924 VPB.n923 13.653
R749 VPB.n923 VPB.n922 13.653
R750 VPB.n929 VPB.n928 13.653
R751 VPB.n928 VPB.n927 13.653
R752 VPB.n934 VPB.n933 13.653
R753 VPB.n933 VPB.n932 13.653
R754 VPB.n938 VPB.n937 13.653
R755 VPB.n937 VPB.n936 13.653
R756 VPB.n965 VPB.n964 13.653
R757 VPB.n964 VPB.n963 13.653
R758 VPB.n969 VPB.n968 13.653
R759 VPB.n968 VPB.n967 13.653
R760 VPB.n974 VPB.n973 13.653
R761 VPB.n973 VPB.n972 13.653
R762 VPB.n979 VPB.n978 13.653
R763 VPB.n978 VPB.n977 13.653
R764 VPB.n986 VPB.n985 13.653
R765 VPB.n985 VPB.n984 13.653
R766 VPB.n991 VPB.n990 13.653
R767 VPB.n990 VPB.n989 13.653
R768 VPB.n996 VPB.n995 13.653
R769 VPB.n995 VPB.n994 13.653
R770 VPB.n1003 VPB.n1002 13.653
R771 VPB.n1002 VPB.n1001 13.653
R772 VPB.n1008 VPB.n1007 13.653
R773 VPB.n1007 VPB.n1006 13.653
R774 VPB.n1013 VPB.n1012 13.653
R775 VPB.n1012 VPB.n1011 13.653
R776 VPB.n1017 VPB.n1016 13.653
R777 VPB.n1016 VPB.n1015 13.653
R778 VPB.n1021 VPB.n1020 13.653
R779 VPB.n1020 VPB.n1019 13.653
R780 VPB.n1048 VPB.n1047 13.653
R781 VPB.n1047 VPB.n1046 13.653
R782 VPB.n1052 VPB.n1051 13.653
R783 VPB.n1051 VPB.n1050 13.653
R784 VPB.n1057 VPB.n1056 13.653
R785 VPB.n1056 VPB.n1055 13.653
R786 VPB.n1062 VPB.n1061 13.653
R787 VPB.n1061 VPB.n1060 13.653
R788 VPB.n1069 VPB.n1068 13.653
R789 VPB.n1068 VPB.n1067 13.653
R790 VPB.n1074 VPB.n1073 13.653
R791 VPB.n1073 VPB.n1072 13.653
R792 VPB.n1079 VPB.n1078 13.653
R793 VPB.n1078 VPB.n1077 13.653
R794 VPB.n1086 VPB.n1085 13.653
R795 VPB.n1085 VPB.n1084 13.653
R796 VPB.n1091 VPB.n1090 13.653
R797 VPB.n1090 VPB.n1089 13.653
R798 VPB.n1096 VPB.n1095 13.653
R799 VPB.n1095 VPB.n1094 13.653
R800 VPB.n1100 VPB.n1099 13.653
R801 VPB.n1099 VPB.n1098 13.653
R802 VPB.n1104 VPB.n1103 13.653
R803 VPB.n1103 VPB.n1102 13.653
R804 VPB.n1131 VPB.n1130 13.653
R805 VPB.n1130 VPB.n1129 13.653
R806 VPB.n1136 VPB.n1135 13.653
R807 VPB.n1135 VPB.n1134 13.653
R808 VPB.n1141 VPB.n1140 13.653
R809 VPB.n1140 VPB.n1139 13.653
R810 VPB.n1148 VPB.n1147 13.653
R811 VPB.n1147 VPB.n1146 13.653
R812 VPB.n1153 VPB.n1152 13.653
R813 VPB.n1152 VPB.n1151 13.653
R814 VPB.n1158 VPB.n1157 13.653
R815 VPB.n1157 VPB.n1156 13.653
R816 VPB.n1163 VPB.n1162 13.653
R817 VPB.n1162 VPB.n1161 13.653
R818 VPB.n1167 VPB.n1166 13.653
R819 VPB.n1166 VPB.n1165 13.653
R820 VPB.n1194 VPB.n1193 13.653
R821 VPB.n1193 VPB.n1192 13.653
R822 VPB.n1198 VPB.n1197 13.653
R823 VPB.n1197 VPB.n1196 13.653
R824 VPB.n1203 VPB.n1202 13.653
R825 VPB.n1202 VPB.n1201 13.653
R826 VPB.n1208 VPB.n1207 13.653
R827 VPB.n1207 VPB.n1206 13.653
R828 VPB.n1215 VPB.n1214 13.653
R829 VPB.n1214 VPB.n1213 13.653
R830 VPB.n1220 VPB.n1219 13.653
R831 VPB.n1219 VPB.n1218 13.653
R832 VPB.n1225 VPB.n1224 13.653
R833 VPB.n1224 VPB.n1223 13.653
R834 VPB.n1232 VPB.n1231 13.653
R835 VPB.n1231 VPB.n1230 13.653
R836 VPB.n1237 VPB.n1236 13.653
R837 VPB.n1236 VPB.n1235 13.653
R838 VPB.n1242 VPB.n1241 13.653
R839 VPB.n1241 VPB.n1240 13.653
R840 VPB.n1246 VPB.n1245 13.653
R841 VPB.n1245 VPB.n1244 13.653
R842 VPB.n1250 VPB.n1249 13.653
R843 VPB.n1249 VPB.n1248 13.653
R844 VPB.n1277 VPB.n1276 13.653
R845 VPB.n1276 VPB.n1275 13.653
R846 VPB.n1282 VPB.n1281 13.653
R847 VPB.n1281 VPB.n1280 13.653
R848 VPB.n1287 VPB.n1286 13.653
R849 VPB.n1286 VPB.n1285 13.653
R850 VPB.n1294 VPB.n1293 13.653
R851 VPB.n1293 VPB.n1292 13.653
R852 VPB.n1299 VPB.n1298 13.653
R853 VPB.n1298 VPB.n1297 13.653
R854 VPB.n1304 VPB.n1303 13.653
R855 VPB.n1303 VPB.n1302 13.653
R856 VPB.n1309 VPB.n1308 13.653
R857 VPB.n1308 VPB.n1307 13.653
R858 VPB.n1313 VPB.n1312 13.653
R859 VPB.n1312 VPB.n1311 13.653
R860 VPB.n1340 VPB.n1339 13.653
R861 VPB.n1339 VPB.n1338 13.653
R862 VPB.n1345 VPB.n1344 13.653
R863 VPB.n1344 VPB.n1343 13.653
R864 VPB.n1350 VPB.n1349 13.653
R865 VPB.n1349 VPB.n1348 13.653
R866 VPB.n1357 VPB.n1356 13.653
R867 VPB.n1356 VPB.n1355 13.653
R868 VPB.n1362 VPB.n1361 13.653
R869 VPB.n1361 VPB.n1360 13.653
R870 VPB.n1367 VPB.n1366 13.653
R871 VPB.n1366 VPB.n1365 13.653
R872 VPB.n1372 VPB.n1371 13.653
R873 VPB.n1371 VPB.n1370 13.653
R874 VPB.n1376 VPB.n1375 13.653
R875 VPB.n1375 VPB.n1374 13.653
R876 VPB.n1403 VPB.n1402 13.653
R877 VPB.n1402 VPB.n1401 13.653
R878 VPB.n1407 VPB.n1406 13.653
R879 VPB.n1406 VPB.n1405 13.653
R880 VPB.n1412 VPB.n1411 13.653
R881 VPB.n1411 VPB.n1410 13.653
R882 VPB.n1417 VPB.n1416 13.653
R883 VPB.n1416 VPB.n1415 13.653
R884 VPB.n1424 VPB.n1423 13.653
R885 VPB.n1423 VPB.n1422 13.653
R886 VPB.n1429 VPB.n1428 13.653
R887 VPB.n1428 VPB.n1427 13.653
R888 VPB.n1434 VPB.n1433 13.653
R889 VPB.n1433 VPB.n1432 13.653
R890 VPB.n1441 VPB.n1440 13.653
R891 VPB.n1440 VPB.n1439 13.653
R892 VPB.n1446 VPB.n1445 13.653
R893 VPB.n1445 VPB.n1444 13.653
R894 VPB.n1451 VPB.n1450 13.653
R895 VPB.n1450 VPB.n1449 13.653
R896 VPB.n1455 VPB.n1454 13.653
R897 VPB.n1454 VPB.n1453 13.653
R898 VPB.n1459 VPB.n1458 13.653
R899 VPB.n1458 VPB.n1457 13.653
R900 VPB.n1486 VPB.n1485 13.653
R901 VPB.n1485 VPB.n1484 13.653
R902 VPB.n1490 VPB.n1489 13.653
R903 VPB.n1489 VPB.n1488 13.653
R904 VPB.n1495 VPB.n1494 13.653
R905 VPB.n1494 VPB.n1493 13.653
R906 VPB.n1500 VPB.n1499 13.653
R907 VPB.n1499 VPB.n1498 13.653
R908 VPB.n1507 VPB.n1506 13.653
R909 VPB.n1506 VPB.n1505 13.653
R910 VPB.n1512 VPB.n1511 13.653
R911 VPB.n1511 VPB.n1510 13.653
R912 VPB.n1517 VPB.n1516 13.653
R913 VPB.n1516 VPB.n1515 13.653
R914 VPB.n1524 VPB.n1523 13.653
R915 VPB.n1523 VPB.n1522 13.653
R916 VPB.n1529 VPB.n1528 13.653
R917 VPB.n1528 VPB.n1527 13.653
R918 VPB.n38 VPB.n37 13.653
R919 VPB.n37 VPB.n36 13.653
R920 VPB.n42 VPB.n41 13.653
R921 VPB.n41 VPB.n40 13.653
R922 VPB.n45 VPB.n44 13.653
R923 VPB.n44 VPB.n43 13.653
R924 VPB.n50 VPB.n49 13.653
R925 VPB.n49 VPB.n48 13.653
R926 VPB.n53 VPB.n52 13.653
R927 VPB.n52 VPB.n51 13.653
R928 VPB.n58 VPB.n57 13.653
R929 VPB.n57 VPB.n56 13.653
R930 VPB.n62 VPB.n61 13.653
R931 VPB.n61 VPB.n60 13.653
R932 VPB.n67 VPB.n66 13.653
R933 VPB.n66 VPB.n65 13.653
R934 VPB.n71 VPB.n70 13.653
R935 VPB.n70 VPB.n69 13.653
R936 VPB.n75 VPB.n74 13.653
R937 VPB.n74 VPB.n73 13.653
R938 VPB.n1542 VPB.n0 13.653
R939 VPB VPB.n0 13.653
R940 VPB.n339 VPB.n338 13.35
R941 VPB.n411 VPB.n410 13.35
R942 VPB.n485 VPB.n484 13.35
R943 VPB.n548 VPB.n547 13.35
R944 VPB.n620 VPB.n619 13.35
R945 VPB.n703 VPB.n702 13.35
R946 VPB.n777 VPB.n776 13.35
R947 VPB.n109 VPB.n108 13.35
R948 VPB.n859 VPB.n858 13.35
R949 VPB.n922 VPB.n921 13.35
R950 VPB.n994 VPB.n993 13.35
R951 VPB.n1077 VPB.n1076 13.35
R952 VPB.n1151 VPB.n1150 13.35
R953 VPB.n1223 VPB.n1222 13.35
R954 VPB.n1297 VPB.n1296 13.35
R955 VPB.n1360 VPB.n1359 13.35
R956 VPB.n1432 VPB.n1431 13.35
R957 VPB.n1515 VPB.n1514 13.35
R958 VPB.n65 VPB.n64 13.35
R959 VPB.n1546 VPB.n1545 13.276
R960 VPB.n1545 VPB.n1543 13.276
R961 VPB.n35 VPB.n17 13.276
R962 VPB.n17 VPB.n15 13.276
R963 VPB.n1481 VPB.n1463 13.276
R964 VPB.n1463 VPB.n1461 13.276
R965 VPB.n1398 VPB.n1380 13.276
R966 VPB.n1380 VPB.n1378 13.276
R967 VPB.n1335 VPB.n1317 13.276
R968 VPB.n1317 VPB.n1315 13.276
R969 VPB.n1272 VPB.n1254 13.276
R970 VPB.n1254 VPB.n1252 13.276
R971 VPB.n1189 VPB.n1171 13.276
R972 VPB.n1171 VPB.n1169 13.276
R973 VPB.n1126 VPB.n1108 13.276
R974 VPB.n1108 VPB.n1106 13.276
R975 VPB.n1043 VPB.n1025 13.276
R976 VPB.n1025 VPB.n1023 13.276
R977 VPB.n960 VPB.n942 13.276
R978 VPB.n942 VPB.n940 13.276
R979 VPB.n897 VPB.n879 13.276
R980 VPB.n879 VPB.n877 13.276
R981 VPB.n96 VPB.n78 13.276
R982 VPB.n78 VPB.n76 13.276
R983 VPB.n815 VPB.n797 13.276
R984 VPB.n797 VPB.n795 13.276
R985 VPB.n752 VPB.n734 13.276
R986 VPB.n734 VPB.n732 13.276
R987 VPB.n669 VPB.n651 13.276
R988 VPB.n651 VPB.n649 13.276
R989 VPB.n586 VPB.n568 13.276
R990 VPB.n568 VPB.n566 13.276
R991 VPB.n523 VPB.n505 13.276
R992 VPB.n505 VPB.n503 13.276
R993 VPB.n460 VPB.n442 13.276
R994 VPB.n442 VPB.n440 13.276
R995 VPB.n377 VPB.n359 13.276
R996 VPB.n359 VPB.n357 13.276
R997 VPB.n314 VPB.n296 13.276
R998 VPB.n296 VPB.n294 13.276
R999 VPB.n259 VPB.n241 13.276
R1000 VPB.n241 VPB.n239 13.276
R1001 VPB.n204 VPB.n186 13.276
R1002 VPB.n186 VPB.n184 13.276
R1003 VPB.n209 VPB.n205 13.276
R1004 VPB.n264 VPB.n260 13.276
R1005 VPB.n319 VPB.n315 13.276
R1006 VPB.n382 VPB.n378 13.276
R1007 VPB.n465 VPB.n461 13.276
R1008 VPB.n528 VPB.n524 13.276
R1009 VPB.n591 VPB.n587 13.276
R1010 VPB.n674 VPB.n670 13.276
R1011 VPB.n757 VPB.n753 13.276
R1012 VPB.n820 VPB.n816 13.276
R1013 VPB.n111 VPB.n107 13.276
R1014 VPB.n120 VPB.n116 13.276
R1015 VPB.n123 VPB.n120 13.276
R1016 VPB.n130 VPB.n127 13.276
R1017 VPB.n131 VPB.n130 13.276
R1018 VPB.n135 VPB.n131 13.276
R1019 VPB.n138 VPB.n135 13.276
R1020 VPB.n856 VPB.n850 13.276
R1021 VPB.n902 VPB.n898 13.276
R1022 VPB.n965 VPB.n961 13.276
R1023 VPB.n1048 VPB.n1044 13.276
R1024 VPB.n1131 VPB.n1127 13.276
R1025 VPB.n1194 VPB.n1190 13.276
R1026 VPB.n1277 VPB.n1273 13.276
R1027 VPB.n1340 VPB.n1336 13.276
R1028 VPB.n1403 VPB.n1399 13.276
R1029 VPB.n1486 VPB.n1482 13.276
R1030 VPB.n45 VPB.n42 13.276
R1031 VPB.n46 VPB.n45 13.276
R1032 VPB.n50 VPB.n46 13.276
R1033 VPB.n53 VPB.n50 13.276
R1034 VPB.n62 VPB.n58 13.276
R1035 VPB.n71 VPB.n67 13.276
R1036 VPB.n1542 VPB.n75 13.276
R1037 VPB.n160 VPB.n142 13.276
R1038 VPB.n142 VPB.n140 13.276
R1039 VPB.n147 VPB.n145 12.796
R1040 VPB.n147 VPB.n146 12.564
R1041 VPB.n127 VPB.n124 12.558
R1042 VPB.n42 VPB.n39 12.558
R1043 VPB.n153 VPB.n152 12.198
R1044 VPB.n155 VPB.n154 12.198
R1045 VPB.n153 VPB.n150 12.198
R1046 VPB.n850 VPB.n139 11.841
R1047 VPB.n58 VPB.n54 11.841
R1048 VPB.n72 VPB.n71 11.482
R1049 VPB.n107 VPB.n103 9.329
R1050 VPB.n112 VPB.n111 8.97
R1051 VPB.n160 VPB.n159 7.5
R1052 VPB.n145 VPB.n144 7.5
R1053 VPB.n152 VPB.n151 7.5
R1054 VPB.n150 VPB.n149 7.5
R1055 VPB.n142 VPB.n141 7.5
R1056 VPB.n157 VPB.n143 7.5
R1057 VPB.n186 VPB.n185 7.5
R1058 VPB.n199 VPB.n198 7.5
R1059 VPB.n193 VPB.n192 7.5
R1060 VPB.n195 VPB.n194 7.5
R1061 VPB.n188 VPB.n187 7.5
R1062 VPB.n204 VPB.n203 7.5
R1063 VPB.n241 VPB.n240 7.5
R1064 VPB.n254 VPB.n253 7.5
R1065 VPB.n248 VPB.n247 7.5
R1066 VPB.n250 VPB.n249 7.5
R1067 VPB.n243 VPB.n242 7.5
R1068 VPB.n259 VPB.n258 7.5
R1069 VPB.n296 VPB.n295 7.5
R1070 VPB.n309 VPB.n308 7.5
R1071 VPB.n303 VPB.n302 7.5
R1072 VPB.n305 VPB.n304 7.5
R1073 VPB.n298 VPB.n297 7.5
R1074 VPB.n314 VPB.n313 7.5
R1075 VPB.n359 VPB.n358 7.5
R1076 VPB.n372 VPB.n371 7.5
R1077 VPB.n366 VPB.n365 7.5
R1078 VPB.n368 VPB.n367 7.5
R1079 VPB.n361 VPB.n360 7.5
R1080 VPB.n377 VPB.n376 7.5
R1081 VPB.n442 VPB.n441 7.5
R1082 VPB.n455 VPB.n454 7.5
R1083 VPB.n449 VPB.n448 7.5
R1084 VPB.n451 VPB.n450 7.5
R1085 VPB.n444 VPB.n443 7.5
R1086 VPB.n460 VPB.n459 7.5
R1087 VPB.n505 VPB.n504 7.5
R1088 VPB.n518 VPB.n517 7.5
R1089 VPB.n512 VPB.n511 7.5
R1090 VPB.n514 VPB.n513 7.5
R1091 VPB.n507 VPB.n506 7.5
R1092 VPB.n523 VPB.n522 7.5
R1093 VPB.n568 VPB.n567 7.5
R1094 VPB.n581 VPB.n580 7.5
R1095 VPB.n575 VPB.n574 7.5
R1096 VPB.n577 VPB.n576 7.5
R1097 VPB.n570 VPB.n569 7.5
R1098 VPB.n586 VPB.n585 7.5
R1099 VPB.n651 VPB.n650 7.5
R1100 VPB.n664 VPB.n663 7.5
R1101 VPB.n658 VPB.n657 7.5
R1102 VPB.n660 VPB.n659 7.5
R1103 VPB.n653 VPB.n652 7.5
R1104 VPB.n669 VPB.n668 7.5
R1105 VPB.n734 VPB.n733 7.5
R1106 VPB.n747 VPB.n746 7.5
R1107 VPB.n741 VPB.n740 7.5
R1108 VPB.n743 VPB.n742 7.5
R1109 VPB.n736 VPB.n735 7.5
R1110 VPB.n752 VPB.n751 7.5
R1111 VPB.n797 VPB.n796 7.5
R1112 VPB.n810 VPB.n809 7.5
R1113 VPB.n804 VPB.n803 7.5
R1114 VPB.n806 VPB.n805 7.5
R1115 VPB.n799 VPB.n798 7.5
R1116 VPB.n815 VPB.n814 7.5
R1117 VPB.n78 VPB.n77 7.5
R1118 VPB.n91 VPB.n90 7.5
R1119 VPB.n85 VPB.n84 7.5
R1120 VPB.n87 VPB.n86 7.5
R1121 VPB.n80 VPB.n79 7.5
R1122 VPB.n96 VPB.n95 7.5
R1123 VPB.n879 VPB.n878 7.5
R1124 VPB.n892 VPB.n891 7.5
R1125 VPB.n886 VPB.n885 7.5
R1126 VPB.n888 VPB.n887 7.5
R1127 VPB.n881 VPB.n880 7.5
R1128 VPB.n897 VPB.n896 7.5
R1129 VPB.n942 VPB.n941 7.5
R1130 VPB.n955 VPB.n954 7.5
R1131 VPB.n949 VPB.n948 7.5
R1132 VPB.n951 VPB.n950 7.5
R1133 VPB.n944 VPB.n943 7.5
R1134 VPB.n960 VPB.n959 7.5
R1135 VPB.n1025 VPB.n1024 7.5
R1136 VPB.n1038 VPB.n1037 7.5
R1137 VPB.n1032 VPB.n1031 7.5
R1138 VPB.n1034 VPB.n1033 7.5
R1139 VPB.n1027 VPB.n1026 7.5
R1140 VPB.n1043 VPB.n1042 7.5
R1141 VPB.n1108 VPB.n1107 7.5
R1142 VPB.n1121 VPB.n1120 7.5
R1143 VPB.n1115 VPB.n1114 7.5
R1144 VPB.n1117 VPB.n1116 7.5
R1145 VPB.n1110 VPB.n1109 7.5
R1146 VPB.n1126 VPB.n1125 7.5
R1147 VPB.n1171 VPB.n1170 7.5
R1148 VPB.n1184 VPB.n1183 7.5
R1149 VPB.n1178 VPB.n1177 7.5
R1150 VPB.n1180 VPB.n1179 7.5
R1151 VPB.n1173 VPB.n1172 7.5
R1152 VPB.n1189 VPB.n1188 7.5
R1153 VPB.n1254 VPB.n1253 7.5
R1154 VPB.n1267 VPB.n1266 7.5
R1155 VPB.n1261 VPB.n1260 7.5
R1156 VPB.n1263 VPB.n1262 7.5
R1157 VPB.n1256 VPB.n1255 7.5
R1158 VPB.n1272 VPB.n1271 7.5
R1159 VPB.n1317 VPB.n1316 7.5
R1160 VPB.n1330 VPB.n1329 7.5
R1161 VPB.n1324 VPB.n1323 7.5
R1162 VPB.n1326 VPB.n1325 7.5
R1163 VPB.n1319 VPB.n1318 7.5
R1164 VPB.n1335 VPB.n1334 7.5
R1165 VPB.n1380 VPB.n1379 7.5
R1166 VPB.n1393 VPB.n1392 7.5
R1167 VPB.n1387 VPB.n1386 7.5
R1168 VPB.n1389 VPB.n1388 7.5
R1169 VPB.n1382 VPB.n1381 7.5
R1170 VPB.n1398 VPB.n1397 7.5
R1171 VPB.n1463 VPB.n1462 7.5
R1172 VPB.n1476 VPB.n1475 7.5
R1173 VPB.n1470 VPB.n1469 7.5
R1174 VPB.n1472 VPB.n1471 7.5
R1175 VPB.n1465 VPB.n1464 7.5
R1176 VPB.n1481 VPB.n1480 7.5
R1177 VPB.n17 VPB.n16 7.5
R1178 VPB.n30 VPB.n29 7.5
R1179 VPB.n24 VPB.n23 7.5
R1180 VPB.n26 VPB.n25 7.5
R1181 VPB.n19 VPB.n18 7.5
R1182 VPB.n35 VPB.n34 7.5
R1183 VPB.n1545 VPB.n1544 7.5
R1184 VPB.n12 VPB.n11 7.5
R1185 VPB.n6 VPB.n5 7.5
R1186 VPB.n8 VPB.n7 7.5
R1187 VPB.n2 VPB.n1 7.5
R1188 VPB.n1547 VPB.n1546 7.5
R1189 VPB.n46 VPB.n35 7.176
R1190 VPB.n1482 VPB.n1481 7.176
R1191 VPB.n1399 VPB.n1398 7.176
R1192 VPB.n1336 VPB.n1335 7.176
R1193 VPB.n1273 VPB.n1272 7.176
R1194 VPB.n1190 VPB.n1189 7.176
R1195 VPB.n1127 VPB.n1126 7.176
R1196 VPB.n1044 VPB.n1043 7.176
R1197 VPB.n961 VPB.n960 7.176
R1198 VPB.n898 VPB.n897 7.176
R1199 VPB.n131 VPB.n96 7.176
R1200 VPB.n816 VPB.n815 7.176
R1201 VPB.n753 VPB.n752 7.176
R1202 VPB.n670 VPB.n669 7.176
R1203 VPB.n587 VPB.n586 7.176
R1204 VPB.n524 VPB.n523 7.176
R1205 VPB.n461 VPB.n460 7.176
R1206 VPB.n378 VPB.n377 7.176
R1207 VPB.n315 VPB.n314 7.176
R1208 VPB.n260 VPB.n259 7.176
R1209 VPB.n205 VPB.n204 7.176
R1210 VPB.n67 VPB.n63 6.817
R1211 VPB.n200 VPB.n197 6.729
R1212 VPB.n196 VPB.n193 6.729
R1213 VPB.n191 VPB.n188 6.729
R1214 VPB.n255 VPB.n252 6.729
R1215 VPB.n251 VPB.n248 6.729
R1216 VPB.n246 VPB.n243 6.729
R1217 VPB.n310 VPB.n307 6.729
R1218 VPB.n306 VPB.n303 6.729
R1219 VPB.n301 VPB.n298 6.729
R1220 VPB.n373 VPB.n370 6.729
R1221 VPB.n369 VPB.n366 6.729
R1222 VPB.n364 VPB.n361 6.729
R1223 VPB.n456 VPB.n453 6.729
R1224 VPB.n452 VPB.n449 6.729
R1225 VPB.n447 VPB.n444 6.729
R1226 VPB.n519 VPB.n516 6.729
R1227 VPB.n515 VPB.n512 6.729
R1228 VPB.n510 VPB.n507 6.729
R1229 VPB.n582 VPB.n579 6.729
R1230 VPB.n578 VPB.n575 6.729
R1231 VPB.n573 VPB.n570 6.729
R1232 VPB.n665 VPB.n662 6.729
R1233 VPB.n661 VPB.n658 6.729
R1234 VPB.n656 VPB.n653 6.729
R1235 VPB.n748 VPB.n745 6.729
R1236 VPB.n744 VPB.n741 6.729
R1237 VPB.n739 VPB.n736 6.729
R1238 VPB.n811 VPB.n808 6.729
R1239 VPB.n807 VPB.n804 6.729
R1240 VPB.n802 VPB.n799 6.729
R1241 VPB.n92 VPB.n89 6.729
R1242 VPB.n88 VPB.n85 6.729
R1243 VPB.n83 VPB.n80 6.729
R1244 VPB.n893 VPB.n890 6.729
R1245 VPB.n889 VPB.n886 6.729
R1246 VPB.n884 VPB.n881 6.729
R1247 VPB.n956 VPB.n953 6.729
R1248 VPB.n952 VPB.n949 6.729
R1249 VPB.n947 VPB.n944 6.729
R1250 VPB.n1039 VPB.n1036 6.729
R1251 VPB.n1035 VPB.n1032 6.729
R1252 VPB.n1030 VPB.n1027 6.729
R1253 VPB.n1122 VPB.n1119 6.729
R1254 VPB.n1118 VPB.n1115 6.729
R1255 VPB.n1113 VPB.n1110 6.729
R1256 VPB.n1185 VPB.n1182 6.729
R1257 VPB.n1181 VPB.n1178 6.729
R1258 VPB.n1176 VPB.n1173 6.729
R1259 VPB.n1268 VPB.n1265 6.729
R1260 VPB.n1264 VPB.n1261 6.729
R1261 VPB.n1259 VPB.n1256 6.729
R1262 VPB.n1331 VPB.n1328 6.729
R1263 VPB.n1327 VPB.n1324 6.729
R1264 VPB.n1322 VPB.n1319 6.729
R1265 VPB.n1394 VPB.n1391 6.729
R1266 VPB.n1390 VPB.n1387 6.729
R1267 VPB.n1385 VPB.n1382 6.729
R1268 VPB.n1477 VPB.n1474 6.729
R1269 VPB.n1473 VPB.n1470 6.729
R1270 VPB.n1468 VPB.n1465 6.729
R1271 VPB.n31 VPB.n28 6.729
R1272 VPB.n27 VPB.n24 6.729
R1273 VPB.n22 VPB.n19 6.729
R1274 VPB.n13 VPB.n10 6.729
R1275 VPB.n9 VPB.n6 6.729
R1276 VPB.n4 VPB.n2 6.729
R1277 VPB.n191 VPB.n190 6.728
R1278 VPB.n196 VPB.n195 6.728
R1279 VPB.n200 VPB.n199 6.728
R1280 VPB.n203 VPB.n202 6.728
R1281 VPB.n246 VPB.n245 6.728
R1282 VPB.n251 VPB.n250 6.728
R1283 VPB.n255 VPB.n254 6.728
R1284 VPB.n258 VPB.n257 6.728
R1285 VPB.n301 VPB.n300 6.728
R1286 VPB.n306 VPB.n305 6.728
R1287 VPB.n310 VPB.n309 6.728
R1288 VPB.n313 VPB.n312 6.728
R1289 VPB.n364 VPB.n363 6.728
R1290 VPB.n369 VPB.n368 6.728
R1291 VPB.n373 VPB.n372 6.728
R1292 VPB.n376 VPB.n375 6.728
R1293 VPB.n447 VPB.n446 6.728
R1294 VPB.n452 VPB.n451 6.728
R1295 VPB.n456 VPB.n455 6.728
R1296 VPB.n459 VPB.n458 6.728
R1297 VPB.n510 VPB.n509 6.728
R1298 VPB.n515 VPB.n514 6.728
R1299 VPB.n519 VPB.n518 6.728
R1300 VPB.n522 VPB.n521 6.728
R1301 VPB.n573 VPB.n572 6.728
R1302 VPB.n578 VPB.n577 6.728
R1303 VPB.n582 VPB.n581 6.728
R1304 VPB.n585 VPB.n584 6.728
R1305 VPB.n656 VPB.n655 6.728
R1306 VPB.n661 VPB.n660 6.728
R1307 VPB.n665 VPB.n664 6.728
R1308 VPB.n668 VPB.n667 6.728
R1309 VPB.n739 VPB.n738 6.728
R1310 VPB.n744 VPB.n743 6.728
R1311 VPB.n748 VPB.n747 6.728
R1312 VPB.n751 VPB.n750 6.728
R1313 VPB.n802 VPB.n801 6.728
R1314 VPB.n807 VPB.n806 6.728
R1315 VPB.n811 VPB.n810 6.728
R1316 VPB.n814 VPB.n813 6.728
R1317 VPB.n83 VPB.n82 6.728
R1318 VPB.n88 VPB.n87 6.728
R1319 VPB.n92 VPB.n91 6.728
R1320 VPB.n95 VPB.n94 6.728
R1321 VPB.n884 VPB.n883 6.728
R1322 VPB.n889 VPB.n888 6.728
R1323 VPB.n893 VPB.n892 6.728
R1324 VPB.n896 VPB.n895 6.728
R1325 VPB.n947 VPB.n946 6.728
R1326 VPB.n952 VPB.n951 6.728
R1327 VPB.n956 VPB.n955 6.728
R1328 VPB.n959 VPB.n958 6.728
R1329 VPB.n1030 VPB.n1029 6.728
R1330 VPB.n1035 VPB.n1034 6.728
R1331 VPB.n1039 VPB.n1038 6.728
R1332 VPB.n1042 VPB.n1041 6.728
R1333 VPB.n1113 VPB.n1112 6.728
R1334 VPB.n1118 VPB.n1117 6.728
R1335 VPB.n1122 VPB.n1121 6.728
R1336 VPB.n1125 VPB.n1124 6.728
R1337 VPB.n1176 VPB.n1175 6.728
R1338 VPB.n1181 VPB.n1180 6.728
R1339 VPB.n1185 VPB.n1184 6.728
R1340 VPB.n1188 VPB.n1187 6.728
R1341 VPB.n1259 VPB.n1258 6.728
R1342 VPB.n1264 VPB.n1263 6.728
R1343 VPB.n1268 VPB.n1267 6.728
R1344 VPB.n1271 VPB.n1270 6.728
R1345 VPB.n1322 VPB.n1321 6.728
R1346 VPB.n1327 VPB.n1326 6.728
R1347 VPB.n1331 VPB.n1330 6.728
R1348 VPB.n1334 VPB.n1333 6.728
R1349 VPB.n1385 VPB.n1384 6.728
R1350 VPB.n1390 VPB.n1389 6.728
R1351 VPB.n1394 VPB.n1393 6.728
R1352 VPB.n1397 VPB.n1396 6.728
R1353 VPB.n1468 VPB.n1467 6.728
R1354 VPB.n1473 VPB.n1472 6.728
R1355 VPB.n1477 VPB.n1476 6.728
R1356 VPB.n1480 VPB.n1479 6.728
R1357 VPB.n22 VPB.n21 6.728
R1358 VPB.n27 VPB.n26 6.728
R1359 VPB.n31 VPB.n30 6.728
R1360 VPB.n34 VPB.n33 6.728
R1361 VPB.n4 VPB.n3 6.728
R1362 VPB.n9 VPB.n8 6.728
R1363 VPB.n13 VPB.n12 6.728
R1364 VPB.n1548 VPB.n1547 6.728
R1365 VPB.n336 VPB.n332 6.458
R1366 VPB.n482 VPB.n478 6.458
R1367 VPB.n545 VPB.n541 6.458
R1368 VPB.n774 VPB.n770 6.458
R1369 VPB.n856 VPB.n852 6.458
R1370 VPB.n919 VPB.n915 6.458
R1371 VPB.n1148 VPB.n1144 6.458
R1372 VPB.n1294 VPB.n1290 6.458
R1373 VPB.n1357 VPB.n1353 6.458
R1374 VPB.n63 VPB.n62 6.458
R1375 VPB.n159 VPB.n158 6.398
R1376 VPB.n420 VPB.n416 4.305
R1377 VPB.n629 VPB.n625 4.305
R1378 VPB.n712 VPB.n708 4.305
R1379 VPB.n116 VPB.n112 4.305
R1380 VPB.n1003 VPB.n999 4.305
R1381 VPB.n1086 VPB.n1082 4.305
R1382 VPB.n1232 VPB.n1228 4.305
R1383 VPB.n1441 VPB.n1437 4.305
R1384 VPB.n1524 VPB.n1520 4.305
R1385 VPB.n403 VPB.n399 3.947
R1386 VPB.n612 VPB.n608 3.947
R1387 VPB.n695 VPB.n691 3.947
R1388 VPB.n103 VPB.n102 3.947
R1389 VPB.n986 VPB.n982 3.947
R1390 VPB.n1069 VPB.n1065 3.947
R1391 VPB.n1215 VPB.n1211 3.947
R1392 VPB.n1424 VPB.n1420 3.947
R1393 VPB.n1507 VPB.n1503 3.947
R1394 VPB.n168 VPB.n164 2.691
R1395 VPB.n178 VPB.n174 2.332
R1396 VPB.n351 VPB.n348 1.794
R1397 VPB.n497 VPB.n494 1.794
R1398 VPB.n560 VPB.n557 1.794
R1399 VPB.n789 VPB.n786 1.794
R1400 VPB.n871 VPB.n868 1.794
R1401 VPB.n934 VPB.n931 1.794
R1402 VPB.n1163 VPB.n1160 1.794
R1403 VPB.n1309 VPB.n1306 1.794
R1404 VPB.n1372 VPB.n1369 1.794
R1405 VPB.n75 VPB.n72 1.794
R1406 VPB.n324 VPB.n321 1.435
R1407 VPB.n470 VPB.n467 1.435
R1408 VPB.n533 VPB.n530 1.435
R1409 VPB.n762 VPB.n759 1.435
R1410 VPB.n139 VPB.n138 1.435
R1411 VPB.n907 VPB.n904 1.435
R1412 VPB.n1136 VPB.n1133 1.435
R1413 VPB.n1282 VPB.n1279 1.435
R1414 VPB.n1345 VPB.n1342 1.435
R1415 VPB.n54 VPB.n53 1.435
R1416 VPB.n157 VPB.n148 1.402
R1417 VPB.n157 VPB.n153 1.402
R1418 VPB.n157 VPB.n155 1.402
R1419 VPB.n157 VPB.n156 1.402
R1420 VPB.n391 VPB.n388 1.076
R1421 VPB.n600 VPB.n597 1.076
R1422 VPB.n683 VPB.n680 1.076
R1423 VPB.n829 VPB.n826 1.076
R1424 VPB.n974 VPB.n971 1.076
R1425 VPB.n1057 VPB.n1054 1.076
R1426 VPB.n1203 VPB.n1200 1.076
R1427 VPB.n1412 VPB.n1409 1.076
R1428 VPB.n1495 VPB.n1492 1.076
R1429 VPB.n158 VPB.n157 0.735
R1430 VPB.n157 VPB.n147 0.735
R1431 VPB.n430 VPB.n427 0.717
R1432 VPB.n639 VPB.n636 0.717
R1433 VPB.n722 VPB.n719 0.717
R1434 VPB.n124 VPB.n123 0.717
R1435 VPB.n1013 VPB.n1010 0.717
R1436 VPB.n1096 VPB.n1093 0.717
R1437 VPB.n1242 VPB.n1239 0.717
R1438 VPB.n1451 VPB.n1448 0.717
R1439 VPB.n39 VPB.n38 0.717
R1440 VPB.n201 VPB.n200 0.387
R1441 VPB.n201 VPB.n196 0.387
R1442 VPB.n201 VPB.n191 0.387
R1443 VPB.n202 VPB.n201 0.387
R1444 VPB.n256 VPB.n255 0.387
R1445 VPB.n256 VPB.n251 0.387
R1446 VPB.n256 VPB.n246 0.387
R1447 VPB.n257 VPB.n256 0.387
R1448 VPB.n311 VPB.n310 0.387
R1449 VPB.n311 VPB.n306 0.387
R1450 VPB.n311 VPB.n301 0.387
R1451 VPB.n312 VPB.n311 0.387
R1452 VPB.n374 VPB.n373 0.387
R1453 VPB.n374 VPB.n369 0.387
R1454 VPB.n374 VPB.n364 0.387
R1455 VPB.n375 VPB.n374 0.387
R1456 VPB.n457 VPB.n456 0.387
R1457 VPB.n457 VPB.n452 0.387
R1458 VPB.n457 VPB.n447 0.387
R1459 VPB.n458 VPB.n457 0.387
R1460 VPB.n520 VPB.n519 0.387
R1461 VPB.n520 VPB.n515 0.387
R1462 VPB.n520 VPB.n510 0.387
R1463 VPB.n521 VPB.n520 0.387
R1464 VPB.n583 VPB.n582 0.387
R1465 VPB.n583 VPB.n578 0.387
R1466 VPB.n583 VPB.n573 0.387
R1467 VPB.n584 VPB.n583 0.387
R1468 VPB.n666 VPB.n665 0.387
R1469 VPB.n666 VPB.n661 0.387
R1470 VPB.n666 VPB.n656 0.387
R1471 VPB.n667 VPB.n666 0.387
R1472 VPB.n749 VPB.n748 0.387
R1473 VPB.n749 VPB.n744 0.387
R1474 VPB.n749 VPB.n739 0.387
R1475 VPB.n750 VPB.n749 0.387
R1476 VPB.n812 VPB.n811 0.387
R1477 VPB.n812 VPB.n807 0.387
R1478 VPB.n812 VPB.n802 0.387
R1479 VPB.n813 VPB.n812 0.387
R1480 VPB.n93 VPB.n92 0.387
R1481 VPB.n93 VPB.n88 0.387
R1482 VPB.n93 VPB.n83 0.387
R1483 VPB.n94 VPB.n93 0.387
R1484 VPB.n894 VPB.n893 0.387
R1485 VPB.n894 VPB.n889 0.387
R1486 VPB.n894 VPB.n884 0.387
R1487 VPB.n895 VPB.n894 0.387
R1488 VPB.n957 VPB.n956 0.387
R1489 VPB.n957 VPB.n952 0.387
R1490 VPB.n957 VPB.n947 0.387
R1491 VPB.n958 VPB.n957 0.387
R1492 VPB.n1040 VPB.n1039 0.387
R1493 VPB.n1040 VPB.n1035 0.387
R1494 VPB.n1040 VPB.n1030 0.387
R1495 VPB.n1041 VPB.n1040 0.387
R1496 VPB.n1123 VPB.n1122 0.387
R1497 VPB.n1123 VPB.n1118 0.387
R1498 VPB.n1123 VPB.n1113 0.387
R1499 VPB.n1124 VPB.n1123 0.387
R1500 VPB.n1186 VPB.n1185 0.387
R1501 VPB.n1186 VPB.n1181 0.387
R1502 VPB.n1186 VPB.n1176 0.387
R1503 VPB.n1187 VPB.n1186 0.387
R1504 VPB.n1269 VPB.n1268 0.387
R1505 VPB.n1269 VPB.n1264 0.387
R1506 VPB.n1269 VPB.n1259 0.387
R1507 VPB.n1270 VPB.n1269 0.387
R1508 VPB.n1332 VPB.n1331 0.387
R1509 VPB.n1332 VPB.n1327 0.387
R1510 VPB.n1332 VPB.n1322 0.387
R1511 VPB.n1333 VPB.n1332 0.387
R1512 VPB.n1395 VPB.n1394 0.387
R1513 VPB.n1395 VPB.n1390 0.387
R1514 VPB.n1395 VPB.n1385 0.387
R1515 VPB.n1396 VPB.n1395 0.387
R1516 VPB.n1478 VPB.n1477 0.387
R1517 VPB.n1478 VPB.n1473 0.387
R1518 VPB.n1478 VPB.n1468 0.387
R1519 VPB.n1479 VPB.n1478 0.387
R1520 VPB.n32 VPB.n31 0.387
R1521 VPB.n32 VPB.n27 0.387
R1522 VPB.n32 VPB.n22 0.387
R1523 VPB.n33 VPB.n32 0.387
R1524 VPB.n1549 VPB.n13 0.387
R1525 VPB.n1549 VPB.n9 0.387
R1526 VPB.n1549 VPB.n4 0.387
R1527 VPB.n1549 VPB.n1548 0.387
R1528 VPB.n210 VPB.n183 0.272
R1529 VPB.n265 VPB.n238 0.272
R1530 VPB.n320 VPB.n293 0.272
R1531 VPB.n383 VPB.n356 0.272
R1532 VPB.n466 VPB.n439 0.272
R1533 VPB.n529 VPB.n502 0.272
R1534 VPB.n592 VPB.n565 0.272
R1535 VPB.n675 VPB.n648 0.272
R1536 VPB.n758 VPB.n731 0.272
R1537 VPB.n821 VPB.n794 0.272
R1538 VPB.n844 VPB.n843 0.272
R1539 VPB.n903 VPB.n876 0.272
R1540 VPB.n966 VPB.n939 0.272
R1541 VPB.n1049 VPB.n1022 0.272
R1542 VPB.n1132 VPB.n1105 0.272
R1543 VPB.n1195 VPB.n1168 0.272
R1544 VPB.n1278 VPB.n1251 0.272
R1545 VPB.n1341 VPB.n1314 0.272
R1546 VPB.n1404 VPB.n1377 0.272
R1547 VPB.n1487 VPB.n1460 0.272
R1548 VPB.n1534 VPB.n1533 0.272
R1549 VPB.n1541 VPB 0.198
R1550 VPB.n173 VPB.n169 0.136
R1551 VPB.n179 VPB.n173 0.136
R1552 VPB.n183 VPB.n179 0.136
R1553 VPB.n214 VPB.n210 0.136
R1554 VPB.n218 VPB.n214 0.136
R1555 VPB.n222 VPB.n218 0.136
R1556 VPB.n226 VPB.n222 0.136
R1557 VPB.n230 VPB.n226 0.136
R1558 VPB.n234 VPB.n230 0.136
R1559 VPB.n238 VPB.n234 0.136
R1560 VPB.n269 VPB.n265 0.136
R1561 VPB.n273 VPB.n269 0.136
R1562 VPB.n277 VPB.n273 0.136
R1563 VPB.n281 VPB.n277 0.136
R1564 VPB.n285 VPB.n281 0.136
R1565 VPB.n289 VPB.n285 0.136
R1566 VPB.n293 VPB.n289 0.136
R1567 VPB.n325 VPB.n320 0.136
R1568 VPB.n330 VPB.n325 0.136
R1569 VPB.n337 VPB.n330 0.136
R1570 VPB.n342 VPB.n337 0.136
R1571 VPB.n347 VPB.n342 0.136
R1572 VPB.n352 VPB.n347 0.136
R1573 VPB.n356 VPB.n352 0.136
R1574 VPB.n387 VPB.n383 0.136
R1575 VPB.n392 VPB.n387 0.136
R1576 VPB.n397 VPB.n392 0.136
R1577 VPB.n404 VPB.n397 0.136
R1578 VPB.n409 VPB.n404 0.136
R1579 VPB.n414 VPB.n409 0.136
R1580 VPB.n421 VPB.n414 0.136
R1581 VPB.n426 VPB.n421 0.136
R1582 VPB.n431 VPB.n426 0.136
R1583 VPB.n435 VPB.n431 0.136
R1584 VPB.n439 VPB.n435 0.136
R1585 VPB.n471 VPB.n466 0.136
R1586 VPB.n476 VPB.n471 0.136
R1587 VPB.n483 VPB.n476 0.136
R1588 VPB.n488 VPB.n483 0.136
R1589 VPB.n493 VPB.n488 0.136
R1590 VPB.n498 VPB.n493 0.136
R1591 VPB.n502 VPB.n498 0.136
R1592 VPB.n534 VPB.n529 0.136
R1593 VPB.n539 VPB.n534 0.136
R1594 VPB.n546 VPB.n539 0.136
R1595 VPB.n551 VPB.n546 0.136
R1596 VPB.n556 VPB.n551 0.136
R1597 VPB.n561 VPB.n556 0.136
R1598 VPB.n565 VPB.n561 0.136
R1599 VPB.n596 VPB.n592 0.136
R1600 VPB.n601 VPB.n596 0.136
R1601 VPB.n606 VPB.n601 0.136
R1602 VPB.n613 VPB.n606 0.136
R1603 VPB.n618 VPB.n613 0.136
R1604 VPB.n623 VPB.n618 0.136
R1605 VPB.n630 VPB.n623 0.136
R1606 VPB.n635 VPB.n630 0.136
R1607 VPB.n640 VPB.n635 0.136
R1608 VPB.n644 VPB.n640 0.136
R1609 VPB.n648 VPB.n644 0.136
R1610 VPB.n679 VPB.n675 0.136
R1611 VPB.n684 VPB.n679 0.136
R1612 VPB.n689 VPB.n684 0.136
R1613 VPB.n696 VPB.n689 0.136
R1614 VPB.n701 VPB.n696 0.136
R1615 VPB.n706 VPB.n701 0.136
R1616 VPB.n713 VPB.n706 0.136
R1617 VPB.n718 VPB.n713 0.136
R1618 VPB.n723 VPB.n718 0.136
R1619 VPB.n727 VPB.n723 0.136
R1620 VPB.n731 VPB.n727 0.136
R1621 VPB.n763 VPB.n758 0.136
R1622 VPB.n768 VPB.n763 0.136
R1623 VPB.n775 VPB.n768 0.136
R1624 VPB.n780 VPB.n775 0.136
R1625 VPB.n785 VPB.n780 0.136
R1626 VPB.n790 VPB.n785 0.136
R1627 VPB.n794 VPB.n790 0.136
R1628 VPB.n825 VPB.n821 0.136
R1629 VPB.n830 VPB.n825 0.136
R1630 VPB.n835 VPB.n830 0.136
R1631 VPB.n836 VPB.n835 0.136
R1632 VPB.n837 VPB.n836 0.136
R1633 VPB.n838 VPB.n837 0.136
R1634 VPB.n839 VPB.n838 0.136
R1635 VPB.n840 VPB.n839 0.136
R1636 VPB.n841 VPB.n840 0.136
R1637 VPB.n842 VPB.n841 0.136
R1638 VPB.n843 VPB.n842 0.136
R1639 VPB.n845 VPB.n844 0.136
R1640 VPB.n846 VPB.n845 0.136
R1641 VPB.n862 VPB.n857 0.136
R1642 VPB.n867 VPB.n862 0.136
R1643 VPB.n872 VPB.n867 0.136
R1644 VPB.n876 VPB.n872 0.136
R1645 VPB.n908 VPB.n903 0.136
R1646 VPB.n913 VPB.n908 0.136
R1647 VPB.n920 VPB.n913 0.136
R1648 VPB.n925 VPB.n920 0.136
R1649 VPB.n930 VPB.n925 0.136
R1650 VPB.n935 VPB.n930 0.136
R1651 VPB.n939 VPB.n935 0.136
R1652 VPB.n970 VPB.n966 0.136
R1653 VPB.n975 VPB.n970 0.136
R1654 VPB.n980 VPB.n975 0.136
R1655 VPB.n987 VPB.n980 0.136
R1656 VPB.n992 VPB.n987 0.136
R1657 VPB.n997 VPB.n992 0.136
R1658 VPB.n1004 VPB.n997 0.136
R1659 VPB.n1009 VPB.n1004 0.136
R1660 VPB.n1014 VPB.n1009 0.136
R1661 VPB.n1018 VPB.n1014 0.136
R1662 VPB.n1022 VPB.n1018 0.136
R1663 VPB.n1053 VPB.n1049 0.136
R1664 VPB.n1058 VPB.n1053 0.136
R1665 VPB.n1063 VPB.n1058 0.136
R1666 VPB.n1070 VPB.n1063 0.136
R1667 VPB.n1075 VPB.n1070 0.136
R1668 VPB.n1080 VPB.n1075 0.136
R1669 VPB.n1087 VPB.n1080 0.136
R1670 VPB.n1092 VPB.n1087 0.136
R1671 VPB.n1097 VPB.n1092 0.136
R1672 VPB.n1101 VPB.n1097 0.136
R1673 VPB.n1105 VPB.n1101 0.136
R1674 VPB.n1137 VPB.n1132 0.136
R1675 VPB.n1142 VPB.n1137 0.136
R1676 VPB.n1149 VPB.n1142 0.136
R1677 VPB.n1154 VPB.n1149 0.136
R1678 VPB.n1159 VPB.n1154 0.136
R1679 VPB.n1164 VPB.n1159 0.136
R1680 VPB.n1168 VPB.n1164 0.136
R1681 VPB.n1199 VPB.n1195 0.136
R1682 VPB.n1204 VPB.n1199 0.136
R1683 VPB.n1209 VPB.n1204 0.136
R1684 VPB.n1216 VPB.n1209 0.136
R1685 VPB.n1221 VPB.n1216 0.136
R1686 VPB.n1226 VPB.n1221 0.136
R1687 VPB.n1233 VPB.n1226 0.136
R1688 VPB.n1238 VPB.n1233 0.136
R1689 VPB.n1243 VPB.n1238 0.136
R1690 VPB.n1247 VPB.n1243 0.136
R1691 VPB.n1251 VPB.n1247 0.136
R1692 VPB.n1283 VPB.n1278 0.136
R1693 VPB.n1288 VPB.n1283 0.136
R1694 VPB.n1295 VPB.n1288 0.136
R1695 VPB.n1300 VPB.n1295 0.136
R1696 VPB.n1305 VPB.n1300 0.136
R1697 VPB.n1310 VPB.n1305 0.136
R1698 VPB.n1314 VPB.n1310 0.136
R1699 VPB.n1346 VPB.n1341 0.136
R1700 VPB.n1351 VPB.n1346 0.136
R1701 VPB.n1358 VPB.n1351 0.136
R1702 VPB.n1363 VPB.n1358 0.136
R1703 VPB.n1368 VPB.n1363 0.136
R1704 VPB.n1373 VPB.n1368 0.136
R1705 VPB.n1377 VPB.n1373 0.136
R1706 VPB.n1408 VPB.n1404 0.136
R1707 VPB.n1413 VPB.n1408 0.136
R1708 VPB.n1418 VPB.n1413 0.136
R1709 VPB.n1425 VPB.n1418 0.136
R1710 VPB.n1430 VPB.n1425 0.136
R1711 VPB.n1435 VPB.n1430 0.136
R1712 VPB.n1442 VPB.n1435 0.136
R1713 VPB.n1447 VPB.n1442 0.136
R1714 VPB.n1452 VPB.n1447 0.136
R1715 VPB.n1456 VPB.n1452 0.136
R1716 VPB.n1460 VPB.n1456 0.136
R1717 VPB.n1491 VPB.n1487 0.136
R1718 VPB.n1496 VPB.n1491 0.136
R1719 VPB.n1501 VPB.n1496 0.136
R1720 VPB.n1508 VPB.n1501 0.136
R1721 VPB.n1513 VPB.n1508 0.136
R1722 VPB.n1518 VPB.n1513 0.136
R1723 VPB.n1525 VPB.n1518 0.136
R1724 VPB.n1530 VPB.n1525 0.136
R1725 VPB.n1531 VPB.n1530 0.136
R1726 VPB.n1532 VPB.n1531 0.136
R1727 VPB.n1533 VPB.n1532 0.136
R1728 VPB.n1535 VPB.n1534 0.136
R1729 VPB.n1536 VPB.n1535 0.136
R1730 VPB.n1537 VPB.n1536 0.136
R1731 VPB.n1538 VPB.n1537 0.136
R1732 VPB.n1539 VPB.n1538 0.136
R1733 VPB.n1540 VPB.n1539 0.136
R1734 VPB.n1541 VPB.n1540 0.136
R1735 VPB.n846 VPB 0.068
R1736 VPB.n857 VPB 0.068
R1737 a_3599_383.n7 a_3599_383.t7 512.525
R1738 a_3599_383.n6 a_3599_383.t13 512.525
R1739 a_3599_383.n11 a_3599_383.t15 472.359
R1740 a_3599_383.n11 a_3599_383.t10 384.527
R1741 a_3599_383.n7 a_3599_383.t14 371.139
R1742 a_3599_383.n6 a_3599_383.t8 371.139
R1743 a_3599_383.n8 a_3599_383.n7 258.98
R1744 a_3599_383.n12 a_3599_383.t11 224.666
R1745 a_3599_383.n16 a_3599_383.n14 196.598
R1746 a_3599_383.n14 a_3599_383.n5 180.846
R1747 a_3599_383.n8 a_3599_383.t12 176.995
R1748 a_3599_383.n9 a_3599_383.t9 170.569
R1749 a_3599_383.n10 a_3599_383.n6 169.274
R1750 a_3599_383.n9 a_3599_383.n8 153.043
R1751 a_3599_383.n12 a_3599_383.n11 120.107
R1752 a_3599_383.n13 a_3599_383.n10 116.763
R1753 a_3599_383.n10 a_3599_383.n9 89.705
R1754 a_3599_383.n13 a_3599_383.n12 80.035
R1755 a_3599_383.n4 a_3599_383.n3 79.232
R1756 a_3599_383.n14 a_3599_383.n13 76
R1757 a_3599_383.n5 a_3599_383.n4 63.152
R1758 a_3599_383.n17 a_3599_383.n0 55.263
R1759 a_3599_383.n16 a_3599_383.n15 30
R1760 a_3599_383.n17 a_3599_383.n16 23.684
R1761 a_3599_383.n5 a_3599_383.n1 16.08
R1762 a_3599_383.n4 a_3599_383.n2 16.08
R1763 a_3599_383.n1 a_3599_383.t0 14.282
R1764 a_3599_383.n1 a_3599_383.t5 14.282
R1765 a_3599_383.n2 a_3599_383.t3 14.282
R1766 a_3599_383.n2 a_3599_383.t4 14.282
R1767 a_3599_383.n3 a_3599_383.t2 14.282
R1768 a_3599_383.n3 a_3599_383.t6 14.282
R1769 a_15044_181.n4 a_15044_181.t7 512.525
R1770 a_15044_181.n4 a_15044_181.t9 371.139
R1771 a_15044_181.n5 a_15044_181.t8 273.368
R1772 a_15044_181.n16 a_15044_181.n6 226.775
R1773 a_15044_181.n6 a_15044_181.n5 153.043
R1774 a_15044_181.n6 a_15044_181.n3 110.158
R1775 a_15044_181.n15 a_15044_181.n14 105.802
R1776 a_15044_181.n5 a_15044_181.n4 105.194
R1777 a_15044_181.n15 a_15044_181.n10 96.417
R1778 a_15044_181.n16 a_15044_181.n15 78.403
R1779 a_15044_181.n3 a_15044_181.n2 75.271
R1780 a_15044_181.n19 a_15044_181.n0 55.263
R1781 a_15044_181.n10 a_15044_181.n9 30
R1782 a_15044_181.n18 a_15044_181.n17 30
R1783 a_15044_181.n19 a_15044_181.n18 25.263
R1784 a_15044_181.n8 a_15044_181.n7 24.383
R1785 a_15044_181.n12 a_15044_181.n11 24.383
R1786 a_15044_181.n10 a_15044_181.n8 23.684
R1787 a_15044_181.n18 a_15044_181.n16 20.417
R1788 a_15044_181.n1 a_15044_181.t3 14.282
R1789 a_15044_181.n1 a_15044_181.t2 14.282
R1790 a_15044_181.n2 a_15044_181.t4 14.282
R1791 a_15044_181.n2 a_15044_181.t5 14.282
R1792 a_15044_181.n14 a_15044_181.n13 13.452
R1793 a_15044_181.n3 a_15044_181.n1 12.119
R1794 a_15044_181.n14 a_15044_181.n12 10.62
R1795 a_15533_1005.n3 a_15533_1005.n2 196.002
R1796 a_15533_1005.n4 a_15533_1005.t1 89.553
R1797 a_15533_1005.n2 a_15533_1005.n1 75.271
R1798 a_15533_1005.n4 a_15533_1005.n3 75.214
R1799 a_15533_1005.n2 a_15533_1005.n0 36.52
R1800 a_15533_1005.n3 a_15533_1005.t5 14.338
R1801 a_15533_1005.n0 a_15533_1005.t3 14.282
R1802 a_15533_1005.n0 a_15533_1005.t4 14.282
R1803 a_15533_1005.n1 a_15533_1005.t2 14.282
R1804 a_15533_1005.n1 a_15533_1005.t7 14.282
R1805 a_15533_1005.n5 a_15533_1005.t0 14.282
R1806 a_15533_1005.t6 a_15533_1005.n5 14.282
R1807 a_15533_1005.n5 a_15533_1005.n4 12.122
R1808 a_11033_943.n6 a_11033_943.t7 454.685
R1809 a_11033_943.n8 a_11033_943.t11 454.685
R1810 a_11033_943.n4 a_11033_943.t13 454.685
R1811 a_11033_943.n6 a_11033_943.t6 428.979
R1812 a_11033_943.n8 a_11033_943.t9 428.979
R1813 a_11033_943.n4 a_11033_943.t10 428.979
R1814 a_11033_943.n7 a_11033_943.t8 248.006
R1815 a_11033_943.n9 a_11033_943.t5 248.006
R1816 a_11033_943.n5 a_11033_943.t12 248.006
R1817 a_11033_943.n14 a_11033_943.n12 220.639
R1818 a_11033_943.n12 a_11033_943.n3 135.994
R1819 a_11033_943.n7 a_11033_943.n6 81.941
R1820 a_11033_943.n9 a_11033_943.n8 81.941
R1821 a_11033_943.n5 a_11033_943.n4 81.941
R1822 a_11033_943.n11 a_11033_943.n5 81.396
R1823 a_11033_943.n10 a_11033_943.n9 79.491
R1824 a_11033_943.n3 a_11033_943.n2 76.002
R1825 a_11033_943.n10 a_11033_943.n7 76
R1826 a_11033_943.n12 a_11033_943.n11 76
R1827 a_11033_943.n14 a_11033_943.n13 30
R1828 a_11033_943.n15 a_11033_943.n0 24.383
R1829 a_11033_943.n15 a_11033_943.n14 23.684
R1830 a_11033_943.n1 a_11033_943.t4 14.282
R1831 a_11033_943.n1 a_11033_943.t3 14.282
R1832 a_11033_943.n2 a_11033_943.t1 14.282
R1833 a_11033_943.n2 a_11033_943.t0 14.282
R1834 a_11033_943.n3 a_11033_943.n1 12.85
R1835 a_11033_943.n11 a_11033_943.n10 2.947
R1836 a_8357_1004.n3 a_8357_1004.t5 512.525
R1837 a_8357_1004.n3 a_8357_1004.t6 371.139
R1838 a_8357_1004.n4 a_8357_1004.n3 225.866
R1839 a_8357_1004.n4 a_8357_1004.t7 218.057
R1840 a_8357_1004.n5 a_8357_1004.n2 215.652
R1841 a_8357_1004.n5 a_8357_1004.n4 153.315
R1842 a_8357_1004.n7 a_8357_1004.n5 147.503
R1843 a_8357_1004.n2 a_8357_1004.n1 76.002
R1844 a_8357_1004.n7 a_8357_1004.n6 15.218
R1845 a_8357_1004.n0 a_8357_1004.t0 14.282
R1846 a_8357_1004.n0 a_8357_1004.t2 14.282
R1847 a_8357_1004.n1 a_8357_1004.t4 14.282
R1848 a_8357_1004.n1 a_8357_1004.t3 14.282
R1849 a_8357_1004.n2 a_8357_1004.n0 12.85
R1850 a_8357_1004.n8 a_8357_1004.n7 12.014
R1851 a_8483_383.n10 a_8483_383.t7 475.572
R1852 a_8483_383.n6 a_8483_383.t12 472.359
R1853 a_8483_383.n9 a_8483_383.t8 469.145
R1854 a_8483_383.n6 a_8483_383.t14 384.527
R1855 a_8483_383.n10 a_8483_383.t10 384.527
R1856 a_8483_383.n9 a_8483_383.t13 384.527
R1857 a_8483_383.n7 a_8483_383.t11 277.772
R1858 a_8483_383.n11 a_8483_383.t15 277.772
R1859 a_8483_383.n13 a_8483_383.t9 198.113
R1860 a_8483_383.n14 a_8483_383.n13 171.961
R1861 a_8483_383.n12 a_8483_383.n11 156.851
R1862 a_8483_383.n8 a_8483_383.n7 156.035
R1863 a_8483_383.n16 a_8483_383.n14 143.492
R1864 a_8483_383.n8 a_8483_383.n5 127.74
R1865 a_8483_383.n14 a_8483_383.n8 106.211
R1866 a_8483_383.n13 a_8483_383.n12 79.658
R1867 a_8483_383.n4 a_8483_383.n3 79.232
R1868 a_8483_383.n11 a_8483_383.n10 67.889
R1869 a_8483_383.n7 a_8483_383.n6 67.001
R1870 a_8483_383.n12 a_8483_383.n9 66.88
R1871 a_8483_383.n5 a_8483_383.n4 63.152
R1872 a_8483_383.n16 a_8483_383.n15 30
R1873 a_8483_383.n17 a_8483_383.n0 24.383
R1874 a_8483_383.n17 a_8483_383.n16 23.684
R1875 a_8483_383.n5 a_8483_383.n1 16.08
R1876 a_8483_383.n4 a_8483_383.n2 16.08
R1877 a_8483_383.n1 a_8483_383.t3 14.282
R1878 a_8483_383.n1 a_8483_383.t2 14.282
R1879 a_8483_383.n2 a_8483_383.t5 14.282
R1880 a_8483_383.n2 a_8483_383.t6 14.282
R1881 a_8483_383.n3 a_8483_383.t1 14.282
R1882 a_8483_383.n3 a_8483_383.t0 14.282
R1883 a_9880_73.t0 a_9880_73.n1 93.333
R1884 a_9880_73.n4 a_9880_73.n2 55.07
R1885 a_9880_73.t0 a_9880_73.n0 8.137
R1886 a_9880_73.n4 a_9880_73.n3 4.619
R1887 a_9880_73.t0 a_9880_73.n4 0.071
R1888 VNB VNB.n1367 300.778
R1889 VNB.n184 VNB.n183 199.897
R1890 VNB.n243 VNB.n242 199.897
R1891 VNB.n302 VNB.n301 199.897
R1892 VNB.n354 VNB.n353 199.897
R1893 VNB.n429 VNB.n428 199.897
R1894 VNB.n481 VNB.n480 199.897
R1895 VNB.n540 VNB.n539 199.897
R1896 VNB.n608 VNB.n607 199.897
R1897 VNB.n676 VNB.n675 199.897
R1898 VNB.n728 VNB.n727 199.897
R1899 VNB.n73 VNB.n72 199.897
R1900 VNB.n805 VNB.n804 199.897
R1901 VNB.n864 VNB.n863 199.897
R1902 VNB.n932 VNB.n931 199.897
R1903 VNB.n1000 VNB.n999 199.897
R1904 VNB.n1059 VNB.n1058 199.897
R1905 VNB.n1127 VNB.n1126 199.897
R1906 VNB.n1179 VNB.n1178 199.897
R1907 VNB.n1231 VNB.n1230 199.897
R1908 VNB.n1299 VNB.n1298 199.897
R1909 VNB.n18 VNB.n17 199.897
R1910 VNB.n155 VNB.n154 158.304
R1911 VNB.n252 VNB.n250 154.509
R1912 VNB.n193 VNB.n191 154.509
R1913 VNB.n363 VNB.n361 154.509
R1914 VNB.n311 VNB.n309 154.509
R1915 VNB.n490 VNB.n488 154.509
R1916 VNB.n438 VNB.n436 154.509
R1917 VNB.n617 VNB.n615 154.509
R1918 VNB.n549 VNB.n547 154.509
R1919 VNB.n737 VNB.n735 154.509
R1920 VNB.n685 VNB.n683 154.509
R1921 VNB.n814 VNB.n812 154.509
R1922 VNB.n115 VNB.n113 154.509
R1923 VNB.n941 VNB.n939 154.509
R1924 VNB.n873 VNB.n871 154.509
R1925 VNB.n1068 VNB.n1066 154.509
R1926 VNB.n1009 VNB.n1007 154.509
R1927 VNB.n1188 VNB.n1186 154.509
R1928 VNB.n1136 VNB.n1134 154.509
R1929 VNB.n1308 VNB.n1306 154.509
R1930 VNB.n1240 VNB.n1238 154.509
R1931 VNB.n38 VNB.n36 154.509
R1932 VNB.n395 VNB.n394 147.75
R1933 VNB.n96 VNB.n95 147.75
R1934 VNB.n209 VNB.n208 121.366
R1935 VNB.n268 VNB.n267 121.366
R1936 VNB.n407 VNB.n404 121.366
R1937 VNB.n506 VNB.n505 121.366
R1938 VNB.n101 VNB.n99 121.366
R1939 VNB.n771 VNB.n770 121.366
R1940 VNB.n830 VNB.n829 121.366
R1941 VNB.n1025 VNB.n1024 121.366
R1942 VNB.n50 VNB.n49 121.366
R1943 VNB.n144 VNB.n143 105.536
R1944 VNB.n585 VNB.n584 85.559
R1945 VNB.n653 VNB.n652 85.559
R1946 VNB.n909 VNB.n908 85.559
R1947 VNB.n977 VNB.n976 85.559
R1948 VNB.n1104 VNB.n1103 85.559
R1949 VNB.n1276 VNB.n1275 85.559
R1950 VNB.n28 VNB.n24 85.559
R1951 VNB.n331 VNB.n330 84.842
R1952 VNB.n458 VNB.n457 84.842
R1953 VNB.n705 VNB.n704 84.842
R1954 VNB.n1156 VNB.n1155 84.842
R1955 VNB.n1208 VNB.n1207 84.842
R1956 VNB.n147 VNB.n137 76.136
R1957 VNB.n147 VNB.n146 76
R1958 VNB.n1354 VNB.n1353 76
R1959 VNB.n1342 VNB.n1341 76
R1960 VNB.n1338 VNB.n1337 76
R1961 VNB.n1334 VNB.n1333 76
R1962 VNB.n1330 VNB.n1329 76
R1963 VNB.n1326 VNB.n1325 76
R1964 VNB.n1322 VNB.n1321 76
R1965 VNB.n1318 VNB.n1317 76
R1966 VNB.n1314 VNB.n1313 76
R1967 VNB.n1310 VNB.n1309 76
R1968 VNB.n1288 VNB.n1287 76
R1969 VNB.n1284 VNB.n1283 76
R1970 VNB.n1280 VNB.n1279 76
R1971 VNB.n1274 VNB.n1273 76
R1972 VNB.n1270 VNB.n1269 76
R1973 VNB.n1266 VNB.n1265 76
R1974 VNB.n1262 VNB.n1261 76
R1975 VNB.n1258 VNB.n1257 76
R1976 VNB.n1254 VNB.n1253 76
R1977 VNB.n1250 VNB.n1249 76
R1978 VNB.n1246 VNB.n1245 76
R1979 VNB.n1242 VNB.n1241 76
R1980 VNB.n1220 VNB.n1219 76
R1981 VNB.n1216 VNB.n1215 76
R1982 VNB.n1212 VNB.n1211 76
R1983 VNB.n1206 VNB.n1205 76
R1984 VNB.n1202 VNB.n1201 76
R1985 VNB.n1198 VNB.n1197 76
R1986 VNB.n1194 VNB.n1193 76
R1987 VNB.n1190 VNB.n1189 76
R1988 VNB.n1168 VNB.n1167 76
R1989 VNB.n1164 VNB.n1163 76
R1990 VNB.n1160 VNB.n1159 76
R1991 VNB.n1154 VNB.n1153 76
R1992 VNB.n1150 VNB.n1149 76
R1993 VNB.n1146 VNB.n1145 76
R1994 VNB.n1142 VNB.n1141 76
R1995 VNB.n1138 VNB.n1137 76
R1996 VNB.n1116 VNB.n1115 76
R1997 VNB.n1112 VNB.n1111 76
R1998 VNB.n1108 VNB.n1107 76
R1999 VNB.n1102 VNB.n1101 76
R2000 VNB.n1098 VNB.n1097 76
R2001 VNB.n1094 VNB.n1093 76
R2002 VNB.n1090 VNB.n1089 76
R2003 VNB.n1086 VNB.n1085 76
R2004 VNB.n1082 VNB.n1081 76
R2005 VNB.n1078 VNB.n1077 76
R2006 VNB.n1074 VNB.n1073 76
R2007 VNB.n1070 VNB.n1069 76
R2008 VNB.n1048 VNB.n1047 76
R2009 VNB.n1044 VNB.n1043 76
R2010 VNB.n1040 VNB.n1039 76
R2011 VNB.n1029 VNB.n1028 76
R2012 VNB.n1023 VNB.n1022 76
R2013 VNB.n1019 VNB.n1018 76
R2014 VNB.n1015 VNB.n1014 76
R2015 VNB.n1011 VNB.n1010 76
R2016 VNB.n989 VNB.n988 76
R2017 VNB.n985 VNB.n984 76
R2018 VNB.n981 VNB.n980 76
R2019 VNB.n975 VNB.n974 76
R2020 VNB.n971 VNB.n970 76
R2021 VNB.n967 VNB.n966 76
R2022 VNB.n963 VNB.n962 76
R2023 VNB.n959 VNB.n958 76
R2024 VNB.n955 VNB.n954 76
R2025 VNB.n951 VNB.n950 76
R2026 VNB.n947 VNB.n946 76
R2027 VNB.n943 VNB.n942 76
R2028 VNB.n921 VNB.n920 76
R2029 VNB.n917 VNB.n916 76
R2030 VNB.n913 VNB.n912 76
R2031 VNB.n907 VNB.n906 76
R2032 VNB.n903 VNB.n902 76
R2033 VNB.n899 VNB.n898 76
R2034 VNB.n895 VNB.n894 76
R2035 VNB.n891 VNB.n890 76
R2036 VNB.n887 VNB.n886 76
R2037 VNB.n883 VNB.n882 76
R2038 VNB.n879 VNB.n878 76
R2039 VNB.n875 VNB.n874 76
R2040 VNB.n853 VNB.n852 76
R2041 VNB.n849 VNB.n848 76
R2042 VNB.n845 VNB.n844 76
R2043 VNB.n834 VNB.n833 76
R2044 VNB.n828 VNB.n827 76
R2045 VNB.n824 VNB.n823 76
R2046 VNB.n820 VNB.n819 76
R2047 VNB.n816 VNB.n815 76
R2048 VNB.n794 VNB.n793 76
R2049 VNB.n790 VNB.n789 76
R2050 VNB.n786 VNB.n785 76
R2051 VNB.n775 VNB.n774 76
R2052 VNB.n769 VNB.n768 76
R2053 VNB.n765 VNB.n762 76
R2054 VNB.n751 VNB.n750 76
R2055 VNB.n747 VNB.n746 76
R2056 VNB.n743 VNB.n742 76
R2057 VNB.n739 VNB.n738 76
R2058 VNB.n717 VNB.n716 76
R2059 VNB.n713 VNB.n712 76
R2060 VNB.n709 VNB.n708 76
R2061 VNB.n703 VNB.n702 76
R2062 VNB.n699 VNB.n698 76
R2063 VNB.n695 VNB.n694 76
R2064 VNB.n691 VNB.n690 76
R2065 VNB.n687 VNB.n686 76
R2066 VNB.n665 VNB.n664 76
R2067 VNB.n661 VNB.n660 76
R2068 VNB.n657 VNB.n656 76
R2069 VNB.n651 VNB.n650 76
R2070 VNB.n647 VNB.n646 76
R2071 VNB.n643 VNB.n642 76
R2072 VNB.n639 VNB.n638 76
R2073 VNB.n635 VNB.n634 76
R2074 VNB.n631 VNB.n630 76
R2075 VNB.n627 VNB.n626 76
R2076 VNB.n623 VNB.n622 76
R2077 VNB.n619 VNB.n618 76
R2078 VNB.n597 VNB.n596 76
R2079 VNB.n593 VNB.n592 76
R2080 VNB.n589 VNB.n588 76
R2081 VNB.n583 VNB.n582 76
R2082 VNB.n579 VNB.n578 76
R2083 VNB.n575 VNB.n574 76
R2084 VNB.n571 VNB.n570 76
R2085 VNB.n567 VNB.n566 76
R2086 VNB.n563 VNB.n562 76
R2087 VNB.n559 VNB.n558 76
R2088 VNB.n555 VNB.n554 76
R2089 VNB.n551 VNB.n550 76
R2090 VNB.n529 VNB.n528 76
R2091 VNB.n525 VNB.n524 76
R2092 VNB.n521 VNB.n520 76
R2093 VNB.n510 VNB.n509 76
R2094 VNB.n504 VNB.n503 76
R2095 VNB.n500 VNB.n499 76
R2096 VNB.n496 VNB.n495 76
R2097 VNB.n492 VNB.n491 76
R2098 VNB.n470 VNB.n469 76
R2099 VNB.n466 VNB.n465 76
R2100 VNB.n462 VNB.n461 76
R2101 VNB.n456 VNB.n455 76
R2102 VNB.n452 VNB.n451 76
R2103 VNB.n448 VNB.n447 76
R2104 VNB.n444 VNB.n443 76
R2105 VNB.n440 VNB.n439 76
R2106 VNB.n418 VNB.n417 76
R2107 VNB.n414 VNB.n413 76
R2108 VNB.n410 VNB.n409 76
R2109 VNB.n398 VNB.n397 76
R2110 VNB.n393 VNB.n392 76
R2111 VNB.n389 VNB.n388 76
R2112 VNB.n385 VNB.n384 76
R2113 VNB.n381 VNB.n380 76
R2114 VNB.n377 VNB.n376 76
R2115 VNB.n373 VNB.n372 76
R2116 VNB.n369 VNB.n368 76
R2117 VNB.n365 VNB.n364 76
R2118 VNB.n343 VNB.n342 76
R2119 VNB.n339 VNB.n338 76
R2120 VNB.n335 VNB.n334 76
R2121 VNB.n329 VNB.n328 76
R2122 VNB.n325 VNB.n324 76
R2123 VNB.n321 VNB.n320 76
R2124 VNB.n317 VNB.n316 76
R2125 VNB.n313 VNB.n312 76
R2126 VNB.n291 VNB.n290 76
R2127 VNB.n287 VNB.n286 76
R2128 VNB.n283 VNB.n282 76
R2129 VNB.n272 VNB.n271 76
R2130 VNB.n266 VNB.n265 76
R2131 VNB.n262 VNB.n261 76
R2132 VNB.n258 VNB.n257 76
R2133 VNB.n254 VNB.n253 76
R2134 VNB.n232 VNB.n231 76
R2135 VNB.n228 VNB.n227 76
R2136 VNB.n224 VNB.n223 76
R2137 VNB.n213 VNB.n212 76
R2138 VNB.n207 VNB.n206 76
R2139 VNB.n203 VNB.n202 76
R2140 VNB.n199 VNB.n198 76
R2141 VNB.n195 VNB.n194 76
R2142 VNB.n173 VNB.n172 76
R2143 VNB.n169 VNB.n168 76
R2144 VNB.n159 VNB.n158 76
R2145 VNB.n106 VNB.n105 73.875
R2146 VNB.n403 VNB.n402 64.552
R2147 VNB.n104 VNB.n82 64.552
R2148 VNB.n218 VNB.n217 63.835
R2149 VNB.n277 VNB.n276 63.835
R2150 VNB.n515 VNB.n514 63.835
R2151 VNB.n780 VNB.n779 63.835
R2152 VNB.n839 VNB.n838 63.835
R2153 VNB.n1034 VNB.n1033 63.835
R2154 VNB.n54 VNB.n7 63.835
R2155 VNB.n587 VNB.n586 41.971
R2156 VNB.n655 VNB.n654 41.971
R2157 VNB.n911 VNB.n910 41.971
R2158 VNB.n979 VNB.n978 41.971
R2159 VNB.n1106 VNB.n1105 41.971
R2160 VNB.n1278 VNB.n1277 41.971
R2161 VNB.n26 VNB.n25 41.971
R2162 VNB.n163 VNB.t21 39.412
R2163 VNB.n210 VNB.n209 36.937
R2164 VNB.n269 VNB.n268 36.937
R2165 VNB.n407 VNB.n406 36.937
R2166 VNB.n507 VNB.n506 36.937
R2167 VNB.n101 VNB.n100 36.937
R2168 VNB.n772 VNB.n771 36.937
R2169 VNB.n831 VNB.n830 36.937
R2170 VNB.n1026 VNB.n1025 36.937
R2171 VNB.n51 VNB.n50 36.937
R2172 VNB.n333 VNB.n332 36.678
R2173 VNB.n460 VNB.n459 36.678
R2174 VNB.n707 VNB.n706 36.678
R2175 VNB.n1158 VNB.n1157 36.678
R2176 VNB.n1210 VNB.n1209 36.678
R2177 VNB.n141 VNB.n140 35.01
R2178 VNB.n406 VNB.n405 29.844
R2179 VNB.n217 VNB.n216 28.421
R2180 VNB.n276 VNB.n275 28.421
R2181 VNB.n402 VNB.n401 28.421
R2182 VNB.n514 VNB.n513 28.421
R2183 VNB.n82 VNB.n81 28.421
R2184 VNB.n779 VNB.n778 28.421
R2185 VNB.n838 VNB.n837 28.421
R2186 VNB.n1033 VNB.n1032 28.421
R2187 VNB.n7 VNB.n6 28.421
R2188 VNB.n156 VNB.n153 27.855
R2189 VNB.n221 VNB.n220 27.855
R2190 VNB.n280 VNB.n279 27.855
R2191 VNB.n518 VNB.n517 27.855
R2192 VNB.n783 VNB.n782 27.855
R2193 VNB.n842 VNB.n841 27.855
R2194 VNB.n1037 VNB.n1036 27.855
R2195 VNB.n57 VNB.n56 27.855
R2196 VNB.n217 VNB.n215 25.263
R2197 VNB.n276 VNB.n274 25.263
R2198 VNB.n402 VNB.n400 25.263
R2199 VNB.n514 VNB.n512 25.263
R2200 VNB.n82 VNB.n80 25.263
R2201 VNB.n779 VNB.n777 25.263
R2202 VNB.n838 VNB.n836 25.263
R2203 VNB.n1033 VNB.n1031 25.263
R2204 VNB.n7 VNB.n5 25.263
R2205 VNB.n215 VNB.n214 24.383
R2206 VNB.n274 VNB.n273 24.383
R2207 VNB.n400 VNB.n399 24.383
R2208 VNB.n512 VNB.n511 24.383
R2209 VNB.n80 VNB.n79 24.383
R2210 VNB.n777 VNB.n776 24.383
R2211 VNB.n836 VNB.n835 24.383
R2212 VNB.n1031 VNB.n1030 24.383
R2213 VNB.n5 VNB.n4 24.383
R2214 VNB.n137 VNB.n134 20.452
R2215 VNB.n1355 VNB.n1354 20.452
R2216 VNB.n142 VNB.n141 20.094
R2217 VNB.n152 VNB.n151 20.094
R2218 VNB.n165 VNB.n164 20.094
R2219 VNB.n141 VNB.n139 19.017
R2220 VNB.n163 VNB.n162 17.185
R2221 VNB.n157 VNB.n156 16.721
R2222 VNB.n222 VNB.n221 16.721
R2223 VNB.n281 VNB.n280 16.721
R2224 VNB.n519 VNB.n518 16.721
R2225 VNB.n784 VNB.n783 16.721
R2226 VNB.n843 VNB.n842 16.721
R2227 VNB.n1038 VNB.n1037 16.721
R2228 VNB.n58 VNB.n57 16.721
R2229 VNB.n146 VNB.n145 13.653
R2230 VNB.n145 VNB.n144 13.653
R2231 VNB.n158 VNB.n157 13.653
R2232 VNB.n168 VNB.n167 13.653
R2233 VNB.n167 VNB.n166 13.653
R2234 VNB.n172 VNB.n171 13.653
R2235 VNB.n171 VNB.n170 13.653
R2236 VNB.n194 VNB.n193 13.653
R2237 VNB.n193 VNB.n192 13.653
R2238 VNB.n198 VNB.n197 13.653
R2239 VNB.n197 VNB.n196 13.653
R2240 VNB.n202 VNB.n201 13.653
R2241 VNB.n201 VNB.n200 13.653
R2242 VNB.n206 VNB.n205 13.653
R2243 VNB.n205 VNB.n204 13.653
R2244 VNB.n212 VNB.n211 13.653
R2245 VNB.n211 VNB.n210 13.653
R2246 VNB.n223 VNB.n222 13.653
R2247 VNB.n227 VNB.n226 13.653
R2248 VNB.n226 VNB.n225 13.653
R2249 VNB.n231 VNB.n230 13.653
R2250 VNB.n230 VNB.n229 13.653
R2251 VNB.n253 VNB.n252 13.653
R2252 VNB.n252 VNB.n251 13.653
R2253 VNB.n257 VNB.n256 13.653
R2254 VNB.n256 VNB.n255 13.653
R2255 VNB.n261 VNB.n260 13.653
R2256 VNB.n260 VNB.n259 13.653
R2257 VNB.n265 VNB.n264 13.653
R2258 VNB.n264 VNB.n263 13.653
R2259 VNB.n271 VNB.n270 13.653
R2260 VNB.n270 VNB.n269 13.653
R2261 VNB.n282 VNB.n281 13.653
R2262 VNB.n286 VNB.n285 13.653
R2263 VNB.n285 VNB.n284 13.653
R2264 VNB.n290 VNB.n289 13.653
R2265 VNB.n289 VNB.n288 13.653
R2266 VNB.n312 VNB.n311 13.653
R2267 VNB.n311 VNB.n310 13.653
R2268 VNB.n316 VNB.n315 13.653
R2269 VNB.n315 VNB.n314 13.653
R2270 VNB.n320 VNB.n319 13.653
R2271 VNB.n319 VNB.n318 13.653
R2272 VNB.n324 VNB.n323 13.653
R2273 VNB.n323 VNB.n322 13.653
R2274 VNB.n328 VNB.n327 13.653
R2275 VNB.n327 VNB.n326 13.653
R2276 VNB.n334 VNB.n333 13.653
R2277 VNB.n338 VNB.n337 13.653
R2278 VNB.n337 VNB.n336 13.653
R2279 VNB.n342 VNB.n341 13.653
R2280 VNB.n341 VNB.n340 13.653
R2281 VNB.n364 VNB.n363 13.653
R2282 VNB.n363 VNB.n362 13.653
R2283 VNB.n368 VNB.n367 13.653
R2284 VNB.n367 VNB.n366 13.653
R2285 VNB.n372 VNB.n371 13.653
R2286 VNB.n371 VNB.n370 13.653
R2287 VNB.n376 VNB.n375 13.653
R2288 VNB.n375 VNB.n374 13.653
R2289 VNB.n380 VNB.n379 13.653
R2290 VNB.n379 VNB.n378 13.653
R2291 VNB.n384 VNB.n383 13.653
R2292 VNB.n383 VNB.n382 13.653
R2293 VNB.n388 VNB.n387 13.653
R2294 VNB.n387 VNB.n386 13.653
R2295 VNB.n392 VNB.n391 13.653
R2296 VNB.n391 VNB.n390 13.653
R2297 VNB.n397 VNB.n396 13.653
R2298 VNB.n396 VNB.n395 13.653
R2299 VNB.n409 VNB.n408 13.653
R2300 VNB.n408 VNB.n407 13.653
R2301 VNB.n413 VNB.n412 13.653
R2302 VNB.n412 VNB.n411 13.653
R2303 VNB.n417 VNB.n416 13.653
R2304 VNB.n416 VNB.n415 13.653
R2305 VNB.n439 VNB.n438 13.653
R2306 VNB.n438 VNB.n437 13.653
R2307 VNB.n443 VNB.n442 13.653
R2308 VNB.n442 VNB.n441 13.653
R2309 VNB.n447 VNB.n446 13.653
R2310 VNB.n446 VNB.n445 13.653
R2311 VNB.n451 VNB.n450 13.653
R2312 VNB.n450 VNB.n449 13.653
R2313 VNB.n455 VNB.n454 13.653
R2314 VNB.n454 VNB.n453 13.653
R2315 VNB.n461 VNB.n460 13.653
R2316 VNB.n465 VNB.n464 13.653
R2317 VNB.n464 VNB.n463 13.653
R2318 VNB.n469 VNB.n468 13.653
R2319 VNB.n468 VNB.n467 13.653
R2320 VNB.n491 VNB.n490 13.653
R2321 VNB.n490 VNB.n489 13.653
R2322 VNB.n495 VNB.n494 13.653
R2323 VNB.n494 VNB.n493 13.653
R2324 VNB.n499 VNB.n498 13.653
R2325 VNB.n498 VNB.n497 13.653
R2326 VNB.n503 VNB.n502 13.653
R2327 VNB.n502 VNB.n501 13.653
R2328 VNB.n509 VNB.n508 13.653
R2329 VNB.n508 VNB.n507 13.653
R2330 VNB.n520 VNB.n519 13.653
R2331 VNB.n524 VNB.n523 13.653
R2332 VNB.n523 VNB.n522 13.653
R2333 VNB.n528 VNB.n527 13.653
R2334 VNB.n527 VNB.n526 13.653
R2335 VNB.n550 VNB.n549 13.653
R2336 VNB.n549 VNB.n548 13.653
R2337 VNB.n554 VNB.n553 13.653
R2338 VNB.n553 VNB.n552 13.653
R2339 VNB.n558 VNB.n557 13.653
R2340 VNB.n557 VNB.n556 13.653
R2341 VNB.n562 VNB.n561 13.653
R2342 VNB.n561 VNB.n560 13.653
R2343 VNB.n566 VNB.n565 13.653
R2344 VNB.n565 VNB.n564 13.653
R2345 VNB.n570 VNB.n569 13.653
R2346 VNB.n569 VNB.n568 13.653
R2347 VNB.n574 VNB.n573 13.653
R2348 VNB.n573 VNB.n572 13.653
R2349 VNB.n578 VNB.n577 13.653
R2350 VNB.n577 VNB.n576 13.653
R2351 VNB.n582 VNB.n581 13.653
R2352 VNB.n581 VNB.n580 13.653
R2353 VNB.n588 VNB.n587 13.653
R2354 VNB.n592 VNB.n591 13.653
R2355 VNB.n591 VNB.n590 13.653
R2356 VNB.n596 VNB.n595 13.653
R2357 VNB.n595 VNB.n594 13.653
R2358 VNB.n618 VNB.n617 13.653
R2359 VNB.n617 VNB.n616 13.653
R2360 VNB.n622 VNB.n621 13.653
R2361 VNB.n621 VNB.n620 13.653
R2362 VNB.n626 VNB.n625 13.653
R2363 VNB.n625 VNB.n624 13.653
R2364 VNB.n630 VNB.n629 13.653
R2365 VNB.n629 VNB.n628 13.653
R2366 VNB.n634 VNB.n633 13.653
R2367 VNB.n633 VNB.n632 13.653
R2368 VNB.n638 VNB.n637 13.653
R2369 VNB.n637 VNB.n636 13.653
R2370 VNB.n642 VNB.n641 13.653
R2371 VNB.n641 VNB.n640 13.653
R2372 VNB.n646 VNB.n645 13.653
R2373 VNB.n645 VNB.n644 13.653
R2374 VNB.n650 VNB.n649 13.653
R2375 VNB.n649 VNB.n648 13.653
R2376 VNB.n656 VNB.n655 13.653
R2377 VNB.n660 VNB.n659 13.653
R2378 VNB.n659 VNB.n658 13.653
R2379 VNB.n664 VNB.n663 13.653
R2380 VNB.n663 VNB.n662 13.653
R2381 VNB.n686 VNB.n685 13.653
R2382 VNB.n685 VNB.n684 13.653
R2383 VNB.n690 VNB.n689 13.653
R2384 VNB.n689 VNB.n688 13.653
R2385 VNB.n694 VNB.n693 13.653
R2386 VNB.n693 VNB.n692 13.653
R2387 VNB.n698 VNB.n697 13.653
R2388 VNB.n697 VNB.n696 13.653
R2389 VNB.n702 VNB.n701 13.653
R2390 VNB.n701 VNB.n700 13.653
R2391 VNB.n708 VNB.n707 13.653
R2392 VNB.n712 VNB.n711 13.653
R2393 VNB.n711 VNB.n710 13.653
R2394 VNB.n716 VNB.n715 13.653
R2395 VNB.n715 VNB.n714 13.653
R2396 VNB.n738 VNB.n737 13.653
R2397 VNB.n737 VNB.n736 13.653
R2398 VNB.n742 VNB.n741 13.653
R2399 VNB.n741 VNB.n740 13.653
R2400 VNB.n746 VNB.n745 13.653
R2401 VNB.n745 VNB.n744 13.653
R2402 VNB.n750 VNB.n749 13.653
R2403 VNB.n749 VNB.n748 13.653
R2404 VNB.n85 VNB.n84 13.653
R2405 VNB.n84 VNB.n83 13.653
R2406 VNB.n88 VNB.n87 13.653
R2407 VNB.n87 VNB.n86 13.653
R2408 VNB.n91 VNB.n90 13.653
R2409 VNB.n90 VNB.n89 13.653
R2410 VNB.n94 VNB.n93 13.653
R2411 VNB.n93 VNB.n92 13.653
R2412 VNB.n98 VNB.n97 13.653
R2413 VNB.n97 VNB.n96 13.653
R2414 VNB.n103 VNB.n102 13.653
R2415 VNB.n102 VNB.n101 13.653
R2416 VNB.n108 VNB.n107 13.653
R2417 VNB.n107 VNB.n106 13.653
R2418 VNB.n111 VNB.n110 13.653
R2419 VNB.n110 VNB.n109 13.653
R2420 VNB.n116 VNB.n115 13.653
R2421 VNB.n115 VNB.n114 13.653
R2422 VNB.n119 VNB.n118 13.653
R2423 VNB.n118 VNB.n117 13.653
R2424 VNB.n765 VNB.n764 13.653
R2425 VNB.n764 VNB.n763 13.653
R2426 VNB.n768 VNB.n767 13.653
R2427 VNB.n767 VNB.n766 13.653
R2428 VNB.n774 VNB.n773 13.653
R2429 VNB.n773 VNB.n772 13.653
R2430 VNB.n785 VNB.n784 13.653
R2431 VNB.n789 VNB.n788 13.653
R2432 VNB.n788 VNB.n787 13.653
R2433 VNB.n793 VNB.n792 13.653
R2434 VNB.n792 VNB.n791 13.653
R2435 VNB.n815 VNB.n814 13.653
R2436 VNB.n814 VNB.n813 13.653
R2437 VNB.n819 VNB.n818 13.653
R2438 VNB.n818 VNB.n817 13.653
R2439 VNB.n823 VNB.n822 13.653
R2440 VNB.n822 VNB.n821 13.653
R2441 VNB.n827 VNB.n826 13.653
R2442 VNB.n826 VNB.n825 13.653
R2443 VNB.n833 VNB.n832 13.653
R2444 VNB.n832 VNB.n831 13.653
R2445 VNB.n844 VNB.n843 13.653
R2446 VNB.n848 VNB.n847 13.653
R2447 VNB.n847 VNB.n846 13.653
R2448 VNB.n852 VNB.n851 13.653
R2449 VNB.n851 VNB.n850 13.653
R2450 VNB.n874 VNB.n873 13.653
R2451 VNB.n873 VNB.n872 13.653
R2452 VNB.n878 VNB.n877 13.653
R2453 VNB.n877 VNB.n876 13.653
R2454 VNB.n882 VNB.n881 13.653
R2455 VNB.n881 VNB.n880 13.653
R2456 VNB.n886 VNB.n885 13.653
R2457 VNB.n885 VNB.n884 13.653
R2458 VNB.n890 VNB.n889 13.653
R2459 VNB.n889 VNB.n888 13.653
R2460 VNB.n894 VNB.n893 13.653
R2461 VNB.n893 VNB.n892 13.653
R2462 VNB.n898 VNB.n897 13.653
R2463 VNB.n897 VNB.n896 13.653
R2464 VNB.n902 VNB.n901 13.653
R2465 VNB.n901 VNB.n900 13.653
R2466 VNB.n906 VNB.n905 13.653
R2467 VNB.n905 VNB.n904 13.653
R2468 VNB.n912 VNB.n911 13.653
R2469 VNB.n916 VNB.n915 13.653
R2470 VNB.n915 VNB.n914 13.653
R2471 VNB.n920 VNB.n919 13.653
R2472 VNB.n919 VNB.n918 13.653
R2473 VNB.n942 VNB.n941 13.653
R2474 VNB.n941 VNB.n940 13.653
R2475 VNB.n946 VNB.n945 13.653
R2476 VNB.n945 VNB.n944 13.653
R2477 VNB.n950 VNB.n949 13.653
R2478 VNB.n949 VNB.n948 13.653
R2479 VNB.n954 VNB.n953 13.653
R2480 VNB.n953 VNB.n952 13.653
R2481 VNB.n958 VNB.n957 13.653
R2482 VNB.n957 VNB.n956 13.653
R2483 VNB.n962 VNB.n961 13.653
R2484 VNB.n961 VNB.n960 13.653
R2485 VNB.n966 VNB.n965 13.653
R2486 VNB.n965 VNB.n964 13.653
R2487 VNB.n970 VNB.n969 13.653
R2488 VNB.n969 VNB.n968 13.653
R2489 VNB.n974 VNB.n973 13.653
R2490 VNB.n973 VNB.n972 13.653
R2491 VNB.n980 VNB.n979 13.653
R2492 VNB.n984 VNB.n983 13.653
R2493 VNB.n983 VNB.n982 13.653
R2494 VNB.n988 VNB.n987 13.653
R2495 VNB.n987 VNB.n986 13.653
R2496 VNB.n1010 VNB.n1009 13.653
R2497 VNB.n1009 VNB.n1008 13.653
R2498 VNB.n1014 VNB.n1013 13.653
R2499 VNB.n1013 VNB.n1012 13.653
R2500 VNB.n1018 VNB.n1017 13.653
R2501 VNB.n1017 VNB.n1016 13.653
R2502 VNB.n1022 VNB.n1021 13.653
R2503 VNB.n1021 VNB.n1020 13.653
R2504 VNB.n1028 VNB.n1027 13.653
R2505 VNB.n1027 VNB.n1026 13.653
R2506 VNB.n1039 VNB.n1038 13.653
R2507 VNB.n1043 VNB.n1042 13.653
R2508 VNB.n1042 VNB.n1041 13.653
R2509 VNB.n1047 VNB.n1046 13.653
R2510 VNB.n1046 VNB.n1045 13.653
R2511 VNB.n1069 VNB.n1068 13.653
R2512 VNB.n1068 VNB.n1067 13.653
R2513 VNB.n1073 VNB.n1072 13.653
R2514 VNB.n1072 VNB.n1071 13.653
R2515 VNB.n1077 VNB.n1076 13.653
R2516 VNB.n1076 VNB.n1075 13.653
R2517 VNB.n1081 VNB.n1080 13.653
R2518 VNB.n1080 VNB.n1079 13.653
R2519 VNB.n1085 VNB.n1084 13.653
R2520 VNB.n1084 VNB.n1083 13.653
R2521 VNB.n1089 VNB.n1088 13.653
R2522 VNB.n1088 VNB.n1087 13.653
R2523 VNB.n1093 VNB.n1092 13.653
R2524 VNB.n1092 VNB.n1091 13.653
R2525 VNB.n1097 VNB.n1096 13.653
R2526 VNB.n1096 VNB.n1095 13.653
R2527 VNB.n1101 VNB.n1100 13.653
R2528 VNB.n1100 VNB.n1099 13.653
R2529 VNB.n1107 VNB.n1106 13.653
R2530 VNB.n1111 VNB.n1110 13.653
R2531 VNB.n1110 VNB.n1109 13.653
R2532 VNB.n1115 VNB.n1114 13.653
R2533 VNB.n1114 VNB.n1113 13.653
R2534 VNB.n1137 VNB.n1136 13.653
R2535 VNB.n1136 VNB.n1135 13.653
R2536 VNB.n1141 VNB.n1140 13.653
R2537 VNB.n1140 VNB.n1139 13.653
R2538 VNB.n1145 VNB.n1144 13.653
R2539 VNB.n1144 VNB.n1143 13.653
R2540 VNB.n1149 VNB.n1148 13.653
R2541 VNB.n1148 VNB.n1147 13.653
R2542 VNB.n1153 VNB.n1152 13.653
R2543 VNB.n1152 VNB.n1151 13.653
R2544 VNB.n1159 VNB.n1158 13.653
R2545 VNB.n1163 VNB.n1162 13.653
R2546 VNB.n1162 VNB.n1161 13.653
R2547 VNB.n1167 VNB.n1166 13.653
R2548 VNB.n1166 VNB.n1165 13.653
R2549 VNB.n1189 VNB.n1188 13.653
R2550 VNB.n1188 VNB.n1187 13.653
R2551 VNB.n1193 VNB.n1192 13.653
R2552 VNB.n1192 VNB.n1191 13.653
R2553 VNB.n1197 VNB.n1196 13.653
R2554 VNB.n1196 VNB.n1195 13.653
R2555 VNB.n1201 VNB.n1200 13.653
R2556 VNB.n1200 VNB.n1199 13.653
R2557 VNB.n1205 VNB.n1204 13.653
R2558 VNB.n1204 VNB.n1203 13.653
R2559 VNB.n1211 VNB.n1210 13.653
R2560 VNB.n1215 VNB.n1214 13.653
R2561 VNB.n1214 VNB.n1213 13.653
R2562 VNB.n1219 VNB.n1218 13.653
R2563 VNB.n1218 VNB.n1217 13.653
R2564 VNB.n1241 VNB.n1240 13.653
R2565 VNB.n1240 VNB.n1239 13.653
R2566 VNB.n1245 VNB.n1244 13.653
R2567 VNB.n1244 VNB.n1243 13.653
R2568 VNB.n1249 VNB.n1248 13.653
R2569 VNB.n1248 VNB.n1247 13.653
R2570 VNB.n1253 VNB.n1252 13.653
R2571 VNB.n1252 VNB.n1251 13.653
R2572 VNB.n1257 VNB.n1256 13.653
R2573 VNB.n1256 VNB.n1255 13.653
R2574 VNB.n1261 VNB.n1260 13.653
R2575 VNB.n1260 VNB.n1259 13.653
R2576 VNB.n1265 VNB.n1264 13.653
R2577 VNB.n1264 VNB.n1263 13.653
R2578 VNB.n1269 VNB.n1268 13.653
R2579 VNB.n1268 VNB.n1267 13.653
R2580 VNB.n1273 VNB.n1272 13.653
R2581 VNB.n1272 VNB.n1271 13.653
R2582 VNB.n1279 VNB.n1278 13.653
R2583 VNB.n1283 VNB.n1282 13.653
R2584 VNB.n1282 VNB.n1281 13.653
R2585 VNB.n1287 VNB.n1286 13.653
R2586 VNB.n1286 VNB.n1285 13.653
R2587 VNB.n1309 VNB.n1308 13.653
R2588 VNB.n1308 VNB.n1307 13.653
R2589 VNB.n1313 VNB.n1312 13.653
R2590 VNB.n1312 VNB.n1311 13.653
R2591 VNB.n1317 VNB.n1316 13.653
R2592 VNB.n1316 VNB.n1315 13.653
R2593 VNB.n1321 VNB.n1320 13.653
R2594 VNB.n1320 VNB.n1319 13.653
R2595 VNB.n1325 VNB.n1324 13.653
R2596 VNB.n1324 VNB.n1323 13.653
R2597 VNB.n1329 VNB.n1328 13.653
R2598 VNB.n1328 VNB.n1327 13.653
R2599 VNB.n1333 VNB.n1332 13.653
R2600 VNB.n1332 VNB.n1331 13.653
R2601 VNB.n1337 VNB.n1336 13.653
R2602 VNB.n1336 VNB.n1335 13.653
R2603 VNB.n1341 VNB.n1340 13.653
R2604 VNB.n1340 VNB.n1339 13.653
R2605 VNB.n27 VNB.n26 13.653
R2606 VNB.n31 VNB.n30 13.653
R2607 VNB.n30 VNB.n29 13.653
R2608 VNB.n34 VNB.n33 13.653
R2609 VNB.n33 VNB.n32 13.653
R2610 VNB.n39 VNB.n38 13.653
R2611 VNB.n38 VNB.n37 13.653
R2612 VNB.n42 VNB.n41 13.653
R2613 VNB.n41 VNB.n40 13.653
R2614 VNB.n45 VNB.n44 13.653
R2615 VNB.n44 VNB.n43 13.653
R2616 VNB.n48 VNB.n47 13.653
R2617 VNB.n47 VNB.n46 13.653
R2618 VNB.n53 VNB.n52 13.653
R2619 VNB.n52 VNB.n51 13.653
R2620 VNB.n59 VNB.n58 13.653
R2621 VNB.n62 VNB.n61 13.653
R2622 VNB.n61 VNB.n60 13.653
R2623 VNB.n1354 VNB.n0 13.653
R2624 VNB VNB.n0 13.653
R2625 VNB.n137 VNB.n136 13.653
R2626 VNB.n136 VNB.n135 13.653
R2627 VNB.n1362 VNB.n1359 13.577
R2628 VNB.n122 VNB.n120 13.276
R2629 VNB.n134 VNB.n122 13.276
R2630 VNB.n176 VNB.n174 13.276
R2631 VNB.n189 VNB.n176 13.276
R2632 VNB.n235 VNB.n233 13.276
R2633 VNB.n248 VNB.n235 13.276
R2634 VNB.n294 VNB.n292 13.276
R2635 VNB.n307 VNB.n294 13.276
R2636 VNB.n346 VNB.n344 13.276
R2637 VNB.n359 VNB.n346 13.276
R2638 VNB.n421 VNB.n419 13.276
R2639 VNB.n434 VNB.n421 13.276
R2640 VNB.n473 VNB.n471 13.276
R2641 VNB.n486 VNB.n473 13.276
R2642 VNB.n532 VNB.n530 13.276
R2643 VNB.n545 VNB.n532 13.276
R2644 VNB.n600 VNB.n598 13.276
R2645 VNB.n613 VNB.n600 13.276
R2646 VNB.n668 VNB.n666 13.276
R2647 VNB.n681 VNB.n668 13.276
R2648 VNB.n720 VNB.n718 13.276
R2649 VNB.n733 VNB.n720 13.276
R2650 VNB.n65 VNB.n63 13.276
R2651 VNB.n78 VNB.n65 13.276
R2652 VNB.n797 VNB.n795 13.276
R2653 VNB.n810 VNB.n797 13.276
R2654 VNB.n856 VNB.n854 13.276
R2655 VNB.n869 VNB.n856 13.276
R2656 VNB.n924 VNB.n922 13.276
R2657 VNB.n937 VNB.n924 13.276
R2658 VNB.n992 VNB.n990 13.276
R2659 VNB.n1005 VNB.n992 13.276
R2660 VNB.n1051 VNB.n1049 13.276
R2661 VNB.n1064 VNB.n1051 13.276
R2662 VNB.n1119 VNB.n1117 13.276
R2663 VNB.n1132 VNB.n1119 13.276
R2664 VNB.n1171 VNB.n1169 13.276
R2665 VNB.n1184 VNB.n1171 13.276
R2666 VNB.n1223 VNB.n1221 13.276
R2667 VNB.n1236 VNB.n1223 13.276
R2668 VNB.n1291 VNB.n1289 13.276
R2669 VNB.n1304 VNB.n1291 13.276
R2670 VNB.n10 VNB.n8 13.276
R2671 VNB.n23 VNB.n10 13.276
R2672 VNB.n194 VNB.n190 13.276
R2673 VNB.n253 VNB.n249 13.276
R2674 VNB.n312 VNB.n308 13.276
R2675 VNB.n364 VNB.n360 13.276
R2676 VNB.n439 VNB.n435 13.276
R2677 VNB.n491 VNB.n487 13.276
R2678 VNB.n550 VNB.n546 13.276
R2679 VNB.n618 VNB.n614 13.276
R2680 VNB.n686 VNB.n682 13.276
R2681 VNB.n738 VNB.n734 13.276
R2682 VNB.n88 VNB.n85 13.276
R2683 VNB.n91 VNB.n88 13.276
R2684 VNB.n94 VNB.n91 13.276
R2685 VNB.n98 VNB.n94 13.276
R2686 VNB.n103 VNB.n98 13.276
R2687 VNB.n111 VNB.n108 13.276
R2688 VNB.n112 VNB.n111 13.276
R2689 VNB.n116 VNB.n112 13.276
R2690 VNB.n119 VNB.n116 13.276
R2691 VNB.n765 VNB.n119 13.276
R2692 VNB.n768 VNB.n765 13.276
R2693 VNB.n815 VNB.n811 13.276
R2694 VNB.n874 VNB.n870 13.276
R2695 VNB.n942 VNB.n938 13.276
R2696 VNB.n1010 VNB.n1006 13.276
R2697 VNB.n1069 VNB.n1065 13.276
R2698 VNB.n1137 VNB.n1133 13.276
R2699 VNB.n1189 VNB.n1185 13.276
R2700 VNB.n1241 VNB.n1237 13.276
R2701 VNB.n1309 VNB.n1305 13.276
R2702 VNB.n34 VNB.n31 13.276
R2703 VNB.n35 VNB.n34 13.276
R2704 VNB.n39 VNB.n35 13.276
R2705 VNB.n42 VNB.n39 13.276
R2706 VNB.n45 VNB.n42 13.276
R2707 VNB.n48 VNB.n45 13.276
R2708 VNB.n53 VNB.n48 13.276
R2709 VNB.n62 VNB.n59 13.276
R2710 VNB.n1354 VNB.n62 13.276
R2711 VNB.n3 VNB.n1 13.276
R2712 VNB.n1355 VNB.n3 13.276
R2713 VNB.n108 VNB.n104 12.02
R2714 VNB.n31 VNB.n28 12.02
R2715 VNB.n54 VNB.n53 10.764
R2716 VNB.n139 VNB.n138 7.5
R2717 VNB.n150 VNB.n149 7.5
R2718 VNB.n1364 VNB.n1363 7.5
R2719 VNB.n182 VNB.n181 7.5
R2720 VNB.n178 VNB.n177 7.5
R2721 VNB.n176 VNB.n175 7.5
R2722 VNB.n189 VNB.n188 7.5
R2723 VNB.n241 VNB.n240 7.5
R2724 VNB.n237 VNB.n236 7.5
R2725 VNB.n235 VNB.n234 7.5
R2726 VNB.n248 VNB.n247 7.5
R2727 VNB.n300 VNB.n299 7.5
R2728 VNB.n296 VNB.n295 7.5
R2729 VNB.n294 VNB.n293 7.5
R2730 VNB.n307 VNB.n306 7.5
R2731 VNB.n352 VNB.n351 7.5
R2732 VNB.n348 VNB.n347 7.5
R2733 VNB.n346 VNB.n345 7.5
R2734 VNB.n359 VNB.n358 7.5
R2735 VNB.n427 VNB.n426 7.5
R2736 VNB.n423 VNB.n422 7.5
R2737 VNB.n421 VNB.n420 7.5
R2738 VNB.n434 VNB.n433 7.5
R2739 VNB.n479 VNB.n478 7.5
R2740 VNB.n475 VNB.n474 7.5
R2741 VNB.n473 VNB.n472 7.5
R2742 VNB.n486 VNB.n485 7.5
R2743 VNB.n538 VNB.n537 7.5
R2744 VNB.n534 VNB.n533 7.5
R2745 VNB.n532 VNB.n531 7.5
R2746 VNB.n545 VNB.n544 7.5
R2747 VNB.n606 VNB.n605 7.5
R2748 VNB.n602 VNB.n601 7.5
R2749 VNB.n600 VNB.n599 7.5
R2750 VNB.n613 VNB.n612 7.5
R2751 VNB.n674 VNB.n673 7.5
R2752 VNB.n670 VNB.n669 7.5
R2753 VNB.n668 VNB.n667 7.5
R2754 VNB.n681 VNB.n680 7.5
R2755 VNB.n726 VNB.n725 7.5
R2756 VNB.n722 VNB.n721 7.5
R2757 VNB.n720 VNB.n719 7.5
R2758 VNB.n733 VNB.n732 7.5
R2759 VNB.n71 VNB.n70 7.5
R2760 VNB.n67 VNB.n66 7.5
R2761 VNB.n65 VNB.n64 7.5
R2762 VNB.n78 VNB.n77 7.5
R2763 VNB.n803 VNB.n802 7.5
R2764 VNB.n799 VNB.n798 7.5
R2765 VNB.n797 VNB.n796 7.5
R2766 VNB.n810 VNB.n809 7.5
R2767 VNB.n862 VNB.n861 7.5
R2768 VNB.n858 VNB.n857 7.5
R2769 VNB.n856 VNB.n855 7.5
R2770 VNB.n869 VNB.n868 7.5
R2771 VNB.n930 VNB.n929 7.5
R2772 VNB.n926 VNB.n925 7.5
R2773 VNB.n924 VNB.n923 7.5
R2774 VNB.n937 VNB.n936 7.5
R2775 VNB.n998 VNB.n997 7.5
R2776 VNB.n994 VNB.n993 7.5
R2777 VNB.n992 VNB.n991 7.5
R2778 VNB.n1005 VNB.n1004 7.5
R2779 VNB.n1057 VNB.n1056 7.5
R2780 VNB.n1053 VNB.n1052 7.5
R2781 VNB.n1051 VNB.n1050 7.5
R2782 VNB.n1064 VNB.n1063 7.5
R2783 VNB.n1125 VNB.n1124 7.5
R2784 VNB.n1121 VNB.n1120 7.5
R2785 VNB.n1119 VNB.n1118 7.5
R2786 VNB.n1132 VNB.n1131 7.5
R2787 VNB.n1177 VNB.n1176 7.5
R2788 VNB.n1173 VNB.n1172 7.5
R2789 VNB.n1171 VNB.n1170 7.5
R2790 VNB.n1184 VNB.n1183 7.5
R2791 VNB.n1229 VNB.n1228 7.5
R2792 VNB.n1225 VNB.n1224 7.5
R2793 VNB.n1223 VNB.n1222 7.5
R2794 VNB.n1236 VNB.n1235 7.5
R2795 VNB.n1297 VNB.n1296 7.5
R2796 VNB.n1293 VNB.n1292 7.5
R2797 VNB.n1291 VNB.n1290 7.5
R2798 VNB.n1304 VNB.n1303 7.5
R2799 VNB.n16 VNB.n15 7.5
R2800 VNB.n12 VNB.n11 7.5
R2801 VNB.n10 VNB.n9 7.5
R2802 VNB.n23 VNB.n22 7.5
R2803 VNB.n1356 VNB.n1355 7.5
R2804 VNB.n3 VNB.n2 7.5
R2805 VNB.n1361 VNB.n1360 7.5
R2806 VNB.n128 VNB.n127 7.5
R2807 VNB.n124 VNB.n123 7.5
R2808 VNB.n122 VNB.n121 7.5
R2809 VNB.n134 VNB.n133 7.5
R2810 VNB.n190 VNB.n189 7.176
R2811 VNB.n249 VNB.n248 7.176
R2812 VNB.n308 VNB.n307 7.176
R2813 VNB.n360 VNB.n359 7.176
R2814 VNB.n435 VNB.n434 7.176
R2815 VNB.n487 VNB.n486 7.176
R2816 VNB.n546 VNB.n545 7.176
R2817 VNB.n614 VNB.n613 7.176
R2818 VNB.n682 VNB.n681 7.176
R2819 VNB.n734 VNB.n733 7.176
R2820 VNB.n112 VNB.n78 7.176
R2821 VNB.n811 VNB.n810 7.176
R2822 VNB.n870 VNB.n869 7.176
R2823 VNB.n938 VNB.n937 7.176
R2824 VNB.n1006 VNB.n1005 7.176
R2825 VNB.n1065 VNB.n1064 7.176
R2826 VNB.n1133 VNB.n1132 7.176
R2827 VNB.n1185 VNB.n1184 7.176
R2828 VNB.n1237 VNB.n1236 7.176
R2829 VNB.n1305 VNB.n1304 7.176
R2830 VNB.n35 VNB.n23 7.176
R2831 VNB.n1366 VNB.n1364 7.011
R2832 VNB.n185 VNB.n182 7.011
R2833 VNB.n180 VNB.n178 7.011
R2834 VNB.n244 VNB.n241 7.011
R2835 VNB.n239 VNB.n237 7.011
R2836 VNB.n303 VNB.n300 7.011
R2837 VNB.n298 VNB.n296 7.011
R2838 VNB.n355 VNB.n352 7.011
R2839 VNB.n350 VNB.n348 7.011
R2840 VNB.n430 VNB.n427 7.011
R2841 VNB.n425 VNB.n423 7.011
R2842 VNB.n482 VNB.n479 7.011
R2843 VNB.n477 VNB.n475 7.011
R2844 VNB.n541 VNB.n538 7.011
R2845 VNB.n536 VNB.n534 7.011
R2846 VNB.n609 VNB.n606 7.011
R2847 VNB.n604 VNB.n602 7.011
R2848 VNB.n677 VNB.n674 7.011
R2849 VNB.n672 VNB.n670 7.011
R2850 VNB.n729 VNB.n726 7.011
R2851 VNB.n724 VNB.n722 7.011
R2852 VNB.n74 VNB.n71 7.011
R2853 VNB.n69 VNB.n67 7.011
R2854 VNB.n806 VNB.n803 7.011
R2855 VNB.n801 VNB.n799 7.011
R2856 VNB.n865 VNB.n862 7.011
R2857 VNB.n860 VNB.n858 7.011
R2858 VNB.n933 VNB.n930 7.011
R2859 VNB.n928 VNB.n926 7.011
R2860 VNB.n1001 VNB.n998 7.011
R2861 VNB.n996 VNB.n994 7.011
R2862 VNB.n1060 VNB.n1057 7.011
R2863 VNB.n1055 VNB.n1053 7.011
R2864 VNB.n1128 VNB.n1125 7.011
R2865 VNB.n1123 VNB.n1121 7.011
R2866 VNB.n1180 VNB.n1177 7.011
R2867 VNB.n1175 VNB.n1173 7.011
R2868 VNB.n1232 VNB.n1229 7.011
R2869 VNB.n1227 VNB.n1225 7.011
R2870 VNB.n1300 VNB.n1297 7.011
R2871 VNB.n1295 VNB.n1293 7.011
R2872 VNB.n19 VNB.n16 7.011
R2873 VNB.n14 VNB.n12 7.011
R2874 VNB.n130 VNB.n128 7.011
R2875 VNB.n126 VNB.n124 7.011
R2876 VNB.n188 VNB.n187 7.01
R2877 VNB.n180 VNB.n179 7.01
R2878 VNB.n185 VNB.n184 7.01
R2879 VNB.n247 VNB.n246 7.01
R2880 VNB.n239 VNB.n238 7.01
R2881 VNB.n244 VNB.n243 7.01
R2882 VNB.n306 VNB.n305 7.01
R2883 VNB.n298 VNB.n297 7.01
R2884 VNB.n303 VNB.n302 7.01
R2885 VNB.n358 VNB.n357 7.01
R2886 VNB.n350 VNB.n349 7.01
R2887 VNB.n355 VNB.n354 7.01
R2888 VNB.n433 VNB.n432 7.01
R2889 VNB.n425 VNB.n424 7.01
R2890 VNB.n430 VNB.n429 7.01
R2891 VNB.n485 VNB.n484 7.01
R2892 VNB.n477 VNB.n476 7.01
R2893 VNB.n482 VNB.n481 7.01
R2894 VNB.n544 VNB.n543 7.01
R2895 VNB.n536 VNB.n535 7.01
R2896 VNB.n541 VNB.n540 7.01
R2897 VNB.n612 VNB.n611 7.01
R2898 VNB.n604 VNB.n603 7.01
R2899 VNB.n609 VNB.n608 7.01
R2900 VNB.n680 VNB.n679 7.01
R2901 VNB.n672 VNB.n671 7.01
R2902 VNB.n677 VNB.n676 7.01
R2903 VNB.n732 VNB.n731 7.01
R2904 VNB.n724 VNB.n723 7.01
R2905 VNB.n729 VNB.n728 7.01
R2906 VNB.n77 VNB.n76 7.01
R2907 VNB.n69 VNB.n68 7.01
R2908 VNB.n74 VNB.n73 7.01
R2909 VNB.n809 VNB.n808 7.01
R2910 VNB.n801 VNB.n800 7.01
R2911 VNB.n806 VNB.n805 7.01
R2912 VNB.n868 VNB.n867 7.01
R2913 VNB.n860 VNB.n859 7.01
R2914 VNB.n865 VNB.n864 7.01
R2915 VNB.n936 VNB.n935 7.01
R2916 VNB.n928 VNB.n927 7.01
R2917 VNB.n933 VNB.n932 7.01
R2918 VNB.n1004 VNB.n1003 7.01
R2919 VNB.n996 VNB.n995 7.01
R2920 VNB.n1001 VNB.n1000 7.01
R2921 VNB.n1063 VNB.n1062 7.01
R2922 VNB.n1055 VNB.n1054 7.01
R2923 VNB.n1060 VNB.n1059 7.01
R2924 VNB.n1131 VNB.n1130 7.01
R2925 VNB.n1123 VNB.n1122 7.01
R2926 VNB.n1128 VNB.n1127 7.01
R2927 VNB.n1183 VNB.n1182 7.01
R2928 VNB.n1175 VNB.n1174 7.01
R2929 VNB.n1180 VNB.n1179 7.01
R2930 VNB.n1235 VNB.n1234 7.01
R2931 VNB.n1227 VNB.n1226 7.01
R2932 VNB.n1232 VNB.n1231 7.01
R2933 VNB.n1303 VNB.n1302 7.01
R2934 VNB.n1295 VNB.n1294 7.01
R2935 VNB.n1300 VNB.n1299 7.01
R2936 VNB.n22 VNB.n21 7.01
R2937 VNB.n14 VNB.n13 7.01
R2938 VNB.n19 VNB.n18 7.01
R2939 VNB.n133 VNB.n132 7.01
R2940 VNB.n126 VNB.n125 7.01
R2941 VNB.n130 VNB.n129 7.01
R2942 VNB.n1366 VNB.n1365 7.01
R2943 VNB.n1362 VNB.n1361 6.788
R2944 VNB.n1357 VNB.n1356 6.788
R2945 VNB.n164 VNB.n163 6.139
R2946 VNB.n161 VNB.n160 4.551
R2947 VNB.n146 VNB.n142 4.305
R2948 VNB.n168 VNB.n165 3.947
R2949 VNB.n223 VNB.n218 2.511
R2950 VNB.n282 VNB.n277 2.511
R2951 VNB.n334 VNB.n331 2.511
R2952 VNB.n461 VNB.n458 2.511
R2953 VNB.n520 VNB.n515 2.511
R2954 VNB.n708 VNB.n705 2.511
R2955 VNB.n785 VNB.n780 2.511
R2956 VNB.n844 VNB.n839 2.511
R2957 VNB.n1039 VNB.n1034 2.511
R2958 VNB.n1159 VNB.n1156 2.511
R2959 VNB.n1211 VNB.n1208 2.511
R2960 VNB.n59 VNB.n54 2.511
R2961 VNB.t21 VNB.n161 2.238
R2962 VNB.n156 VNB.n155 1.99
R2963 VNB.n221 VNB.n219 1.99
R2964 VNB.n280 VNB.n278 1.99
R2965 VNB.n518 VNB.n516 1.99
R2966 VNB.n783 VNB.n781 1.99
R2967 VNB.n842 VNB.n840 1.99
R2968 VNB.n1037 VNB.n1035 1.99
R2969 VNB.n57 VNB.n55 1.99
R2970 VNB.n149 VNB.n148 1.935
R2971 VNB.n409 VNB.n403 1.255
R2972 VNB.n588 VNB.n585 1.255
R2973 VNB.n656 VNB.n653 1.255
R2974 VNB.n104 VNB.n103 1.255
R2975 VNB.n912 VNB.n909 1.255
R2976 VNB.n980 VNB.n977 1.255
R2977 VNB.n1107 VNB.n1104 1.255
R2978 VNB.n1279 VNB.n1276 1.255
R2979 VNB.n28 VNB.n27 1.255
R2980 VNB.n1367 VNB.n1358 0.921
R2981 VNB.n1367 VNB.n1362 0.476
R2982 VNB.n1367 VNB.n1357 0.475
R2983 VNB.n151 VNB.n150 0.358
R2984 VNB.n195 VNB.n173 0.272
R2985 VNB.n254 VNB.n232 0.272
R2986 VNB.n313 VNB.n291 0.272
R2987 VNB.n365 VNB.n343 0.272
R2988 VNB.n440 VNB.n418 0.272
R2989 VNB.n492 VNB.n470 0.272
R2990 VNB.n551 VNB.n529 0.272
R2991 VNB.n619 VNB.n597 0.272
R2992 VNB.n687 VNB.n665 0.272
R2993 VNB.n739 VNB.n717 0.272
R2994 VNB.n760 VNB.n759 0.272
R2995 VNB.n816 VNB.n794 0.272
R2996 VNB.n875 VNB.n853 0.272
R2997 VNB.n943 VNB.n921 0.272
R2998 VNB.n1011 VNB.n989 0.272
R2999 VNB.n1070 VNB.n1048 0.272
R3000 VNB.n1138 VNB.n1116 0.272
R3001 VNB.n1190 VNB.n1168 0.272
R3002 VNB.n1242 VNB.n1220 0.272
R3003 VNB.n1310 VNB.n1288 0.272
R3004 VNB.n1346 VNB.n1345 0.272
R3005 VNB.n186 VNB.n180 0.246
R3006 VNB.n187 VNB.n186 0.246
R3007 VNB.n186 VNB.n185 0.246
R3008 VNB.n245 VNB.n239 0.246
R3009 VNB.n246 VNB.n245 0.246
R3010 VNB.n245 VNB.n244 0.246
R3011 VNB.n304 VNB.n298 0.246
R3012 VNB.n305 VNB.n304 0.246
R3013 VNB.n304 VNB.n303 0.246
R3014 VNB.n356 VNB.n350 0.246
R3015 VNB.n357 VNB.n356 0.246
R3016 VNB.n356 VNB.n355 0.246
R3017 VNB.n431 VNB.n425 0.246
R3018 VNB.n432 VNB.n431 0.246
R3019 VNB.n431 VNB.n430 0.246
R3020 VNB.n483 VNB.n477 0.246
R3021 VNB.n484 VNB.n483 0.246
R3022 VNB.n483 VNB.n482 0.246
R3023 VNB.n542 VNB.n536 0.246
R3024 VNB.n543 VNB.n542 0.246
R3025 VNB.n542 VNB.n541 0.246
R3026 VNB.n610 VNB.n604 0.246
R3027 VNB.n611 VNB.n610 0.246
R3028 VNB.n610 VNB.n609 0.246
R3029 VNB.n678 VNB.n672 0.246
R3030 VNB.n679 VNB.n678 0.246
R3031 VNB.n678 VNB.n677 0.246
R3032 VNB.n730 VNB.n724 0.246
R3033 VNB.n731 VNB.n730 0.246
R3034 VNB.n730 VNB.n729 0.246
R3035 VNB.n75 VNB.n69 0.246
R3036 VNB.n76 VNB.n75 0.246
R3037 VNB.n75 VNB.n74 0.246
R3038 VNB.n807 VNB.n801 0.246
R3039 VNB.n808 VNB.n807 0.246
R3040 VNB.n807 VNB.n806 0.246
R3041 VNB.n866 VNB.n860 0.246
R3042 VNB.n867 VNB.n866 0.246
R3043 VNB.n866 VNB.n865 0.246
R3044 VNB.n934 VNB.n928 0.246
R3045 VNB.n935 VNB.n934 0.246
R3046 VNB.n934 VNB.n933 0.246
R3047 VNB.n1002 VNB.n996 0.246
R3048 VNB.n1003 VNB.n1002 0.246
R3049 VNB.n1002 VNB.n1001 0.246
R3050 VNB.n1061 VNB.n1055 0.246
R3051 VNB.n1062 VNB.n1061 0.246
R3052 VNB.n1061 VNB.n1060 0.246
R3053 VNB.n1129 VNB.n1123 0.246
R3054 VNB.n1130 VNB.n1129 0.246
R3055 VNB.n1129 VNB.n1128 0.246
R3056 VNB.n1181 VNB.n1175 0.246
R3057 VNB.n1182 VNB.n1181 0.246
R3058 VNB.n1181 VNB.n1180 0.246
R3059 VNB.n1233 VNB.n1227 0.246
R3060 VNB.n1234 VNB.n1233 0.246
R3061 VNB.n1233 VNB.n1232 0.246
R3062 VNB.n1301 VNB.n1295 0.246
R3063 VNB.n1302 VNB.n1301 0.246
R3064 VNB.n1301 VNB.n1300 0.246
R3065 VNB.n20 VNB.n14 0.246
R3066 VNB.n21 VNB.n20 0.246
R3067 VNB.n20 VNB.n19 0.246
R3068 VNB.n131 VNB.n126 0.246
R3069 VNB.n132 VNB.n131 0.246
R3070 VNB.n131 VNB.n130 0.246
R3071 VNB.n1367 VNB.n1366 0.246
R3072 VNB.n1353 VNB 0.198
R3073 VNB.n158 VNB.n152 0.179
R3074 VNB.n159 VNB.n147 0.136
R3075 VNB.n169 VNB.n159 0.136
R3076 VNB.n173 VNB.n169 0.136
R3077 VNB.n199 VNB.n195 0.136
R3078 VNB.n203 VNB.n199 0.136
R3079 VNB.n207 VNB.n203 0.136
R3080 VNB.n213 VNB.n207 0.136
R3081 VNB.n224 VNB.n213 0.136
R3082 VNB.n228 VNB.n224 0.136
R3083 VNB.n232 VNB.n228 0.136
R3084 VNB.n258 VNB.n254 0.136
R3085 VNB.n262 VNB.n258 0.136
R3086 VNB.n266 VNB.n262 0.136
R3087 VNB.n272 VNB.n266 0.136
R3088 VNB.n283 VNB.n272 0.136
R3089 VNB.n287 VNB.n283 0.136
R3090 VNB.n291 VNB.n287 0.136
R3091 VNB.n317 VNB.n313 0.136
R3092 VNB.n321 VNB.n317 0.136
R3093 VNB.n325 VNB.n321 0.136
R3094 VNB.n329 VNB.n325 0.136
R3095 VNB.n335 VNB.n329 0.136
R3096 VNB.n339 VNB.n335 0.136
R3097 VNB.n343 VNB.n339 0.136
R3098 VNB.n369 VNB.n365 0.136
R3099 VNB.n373 VNB.n369 0.136
R3100 VNB.n377 VNB.n373 0.136
R3101 VNB.n381 VNB.n377 0.136
R3102 VNB.n385 VNB.n381 0.136
R3103 VNB.n389 VNB.n385 0.136
R3104 VNB.n393 VNB.n389 0.136
R3105 VNB.n398 VNB.n393 0.136
R3106 VNB.n410 VNB.n398 0.136
R3107 VNB.n414 VNB.n410 0.136
R3108 VNB.n418 VNB.n414 0.136
R3109 VNB.n444 VNB.n440 0.136
R3110 VNB.n448 VNB.n444 0.136
R3111 VNB.n452 VNB.n448 0.136
R3112 VNB.n456 VNB.n452 0.136
R3113 VNB.n462 VNB.n456 0.136
R3114 VNB.n466 VNB.n462 0.136
R3115 VNB.n470 VNB.n466 0.136
R3116 VNB.n496 VNB.n492 0.136
R3117 VNB.n500 VNB.n496 0.136
R3118 VNB.n504 VNB.n500 0.136
R3119 VNB.n510 VNB.n504 0.136
R3120 VNB.n521 VNB.n510 0.136
R3121 VNB.n525 VNB.n521 0.136
R3122 VNB.n529 VNB.n525 0.136
R3123 VNB.n555 VNB.n551 0.136
R3124 VNB.n559 VNB.n555 0.136
R3125 VNB.n563 VNB.n559 0.136
R3126 VNB.n567 VNB.n563 0.136
R3127 VNB.n571 VNB.n567 0.136
R3128 VNB.n575 VNB.n571 0.136
R3129 VNB.n579 VNB.n575 0.136
R3130 VNB.n583 VNB.n579 0.136
R3131 VNB.n589 VNB.n583 0.136
R3132 VNB.n593 VNB.n589 0.136
R3133 VNB.n597 VNB.n593 0.136
R3134 VNB.n623 VNB.n619 0.136
R3135 VNB.n627 VNB.n623 0.136
R3136 VNB.n631 VNB.n627 0.136
R3137 VNB.n635 VNB.n631 0.136
R3138 VNB.n639 VNB.n635 0.136
R3139 VNB.n643 VNB.n639 0.136
R3140 VNB.n647 VNB.n643 0.136
R3141 VNB.n651 VNB.n647 0.136
R3142 VNB.n657 VNB.n651 0.136
R3143 VNB.n661 VNB.n657 0.136
R3144 VNB.n665 VNB.n661 0.136
R3145 VNB.n691 VNB.n687 0.136
R3146 VNB.n695 VNB.n691 0.136
R3147 VNB.n699 VNB.n695 0.136
R3148 VNB.n703 VNB.n699 0.136
R3149 VNB.n709 VNB.n703 0.136
R3150 VNB.n713 VNB.n709 0.136
R3151 VNB.n717 VNB.n713 0.136
R3152 VNB.n743 VNB.n739 0.136
R3153 VNB.n747 VNB.n743 0.136
R3154 VNB.n751 VNB.n747 0.136
R3155 VNB.n752 VNB.n751 0.136
R3156 VNB.n753 VNB.n752 0.136
R3157 VNB.n754 VNB.n753 0.136
R3158 VNB.n755 VNB.n754 0.136
R3159 VNB.n756 VNB.n755 0.136
R3160 VNB.n757 VNB.n756 0.136
R3161 VNB.n758 VNB.n757 0.136
R3162 VNB.n759 VNB.n758 0.136
R3163 VNB.n761 VNB.n760 0.136
R3164 VNB.n762 VNB.n761 0.136
R3165 VNB.n775 VNB.n769 0.136
R3166 VNB.n786 VNB.n775 0.136
R3167 VNB.n790 VNB.n786 0.136
R3168 VNB.n794 VNB.n790 0.136
R3169 VNB.n820 VNB.n816 0.136
R3170 VNB.n824 VNB.n820 0.136
R3171 VNB.n828 VNB.n824 0.136
R3172 VNB.n834 VNB.n828 0.136
R3173 VNB.n845 VNB.n834 0.136
R3174 VNB.n849 VNB.n845 0.136
R3175 VNB.n853 VNB.n849 0.136
R3176 VNB.n879 VNB.n875 0.136
R3177 VNB.n883 VNB.n879 0.136
R3178 VNB.n887 VNB.n883 0.136
R3179 VNB.n891 VNB.n887 0.136
R3180 VNB.n895 VNB.n891 0.136
R3181 VNB.n899 VNB.n895 0.136
R3182 VNB.n903 VNB.n899 0.136
R3183 VNB.n907 VNB.n903 0.136
R3184 VNB.n913 VNB.n907 0.136
R3185 VNB.n917 VNB.n913 0.136
R3186 VNB.n921 VNB.n917 0.136
R3187 VNB.n947 VNB.n943 0.136
R3188 VNB.n951 VNB.n947 0.136
R3189 VNB.n955 VNB.n951 0.136
R3190 VNB.n959 VNB.n955 0.136
R3191 VNB.n963 VNB.n959 0.136
R3192 VNB.n967 VNB.n963 0.136
R3193 VNB.n971 VNB.n967 0.136
R3194 VNB.n975 VNB.n971 0.136
R3195 VNB.n981 VNB.n975 0.136
R3196 VNB.n985 VNB.n981 0.136
R3197 VNB.n989 VNB.n985 0.136
R3198 VNB.n1015 VNB.n1011 0.136
R3199 VNB.n1019 VNB.n1015 0.136
R3200 VNB.n1023 VNB.n1019 0.136
R3201 VNB.n1029 VNB.n1023 0.136
R3202 VNB.n1040 VNB.n1029 0.136
R3203 VNB.n1044 VNB.n1040 0.136
R3204 VNB.n1048 VNB.n1044 0.136
R3205 VNB.n1074 VNB.n1070 0.136
R3206 VNB.n1078 VNB.n1074 0.136
R3207 VNB.n1082 VNB.n1078 0.136
R3208 VNB.n1086 VNB.n1082 0.136
R3209 VNB.n1090 VNB.n1086 0.136
R3210 VNB.n1094 VNB.n1090 0.136
R3211 VNB.n1098 VNB.n1094 0.136
R3212 VNB.n1102 VNB.n1098 0.136
R3213 VNB.n1108 VNB.n1102 0.136
R3214 VNB.n1112 VNB.n1108 0.136
R3215 VNB.n1116 VNB.n1112 0.136
R3216 VNB.n1142 VNB.n1138 0.136
R3217 VNB.n1146 VNB.n1142 0.136
R3218 VNB.n1150 VNB.n1146 0.136
R3219 VNB.n1154 VNB.n1150 0.136
R3220 VNB.n1160 VNB.n1154 0.136
R3221 VNB.n1164 VNB.n1160 0.136
R3222 VNB.n1168 VNB.n1164 0.136
R3223 VNB.n1194 VNB.n1190 0.136
R3224 VNB.n1198 VNB.n1194 0.136
R3225 VNB.n1202 VNB.n1198 0.136
R3226 VNB.n1206 VNB.n1202 0.136
R3227 VNB.n1212 VNB.n1206 0.136
R3228 VNB.n1216 VNB.n1212 0.136
R3229 VNB.n1220 VNB.n1216 0.136
R3230 VNB.n1246 VNB.n1242 0.136
R3231 VNB.n1250 VNB.n1246 0.136
R3232 VNB.n1254 VNB.n1250 0.136
R3233 VNB.n1258 VNB.n1254 0.136
R3234 VNB.n1262 VNB.n1258 0.136
R3235 VNB.n1266 VNB.n1262 0.136
R3236 VNB.n1270 VNB.n1266 0.136
R3237 VNB.n1274 VNB.n1270 0.136
R3238 VNB.n1280 VNB.n1274 0.136
R3239 VNB.n1284 VNB.n1280 0.136
R3240 VNB.n1288 VNB.n1284 0.136
R3241 VNB.n1314 VNB.n1310 0.136
R3242 VNB.n1318 VNB.n1314 0.136
R3243 VNB.n1322 VNB.n1318 0.136
R3244 VNB.n1326 VNB.n1322 0.136
R3245 VNB.n1330 VNB.n1326 0.136
R3246 VNB.n1334 VNB.n1330 0.136
R3247 VNB.n1338 VNB.n1334 0.136
R3248 VNB.n1342 VNB.n1338 0.136
R3249 VNB.n1343 VNB.n1342 0.136
R3250 VNB.n1344 VNB.n1343 0.136
R3251 VNB.n1345 VNB.n1344 0.136
R3252 VNB.n1347 VNB.n1346 0.136
R3253 VNB.n1348 VNB.n1347 0.136
R3254 VNB.n1349 VNB.n1348 0.136
R3255 VNB.n1350 VNB.n1349 0.136
R3256 VNB.n1351 VNB.n1350 0.136
R3257 VNB.n1352 VNB.n1351 0.136
R3258 VNB.n1353 VNB.n1352 0.136
R3259 VNB.n762 VNB 0.068
R3260 VNB.n769 VNB 0.068
R3261 a_217_1004.n5 a_217_1004.t7 512.525
R3262 a_217_1004.n3 a_217_1004.t9 512.525
R3263 a_217_1004.n5 a_217_1004.t8 371.139
R3264 a_217_1004.n3 a_217_1004.t6 371.139
R3265 a_217_1004.n6 a_217_1004.n5 226.225
R3266 a_217_1004.n4 a_217_1004.n3 225.866
R3267 a_217_1004.n4 a_217_1004.t5 218.057
R3268 a_217_1004.n6 a_217_1004.t10 217.698
R3269 a_217_1004.n8 a_217_1004.n2 215.652
R3270 a_217_1004.n10 a_217_1004.n8 147.503
R3271 a_217_1004.n7 a_217_1004.n4 79.488
R3272 a_217_1004.n8 a_217_1004.n7 77.314
R3273 a_217_1004.n2 a_217_1004.n1 76.002
R3274 a_217_1004.n7 a_217_1004.n6 76
R3275 a_217_1004.n10 a_217_1004.n9 15.218
R3276 a_217_1004.n0 a_217_1004.t4 14.282
R3277 a_217_1004.n0 a_217_1004.t0 14.282
R3278 a_217_1004.n1 a_217_1004.t2 14.282
R3279 a_217_1004.n1 a_217_1004.t1 14.282
R3280 a_217_1004.n2 a_217_1004.n0 12.85
R3281 a_217_1004.n11 a_217_1004.n10 12.014
R3282 a_1719_75.n4 a_1719_75.n3 19.724
R3283 a_1719_75.t0 a_1719_75.n5 11.595
R3284 a_1719_75.t0 a_1719_75.n4 9.207
R3285 a_1719_75.n2 a_1719_75.n0 8.543
R3286 a_1719_75.t0 a_1719_75.n2 3.034
R3287 a_1719_75.n2 a_1719_75.n1 0.443
R3288 a_14869_1005.n4 a_14869_1005.n3 195.987
R3289 a_14869_1005.n2 a_14869_1005.t6 89.553
R3290 a_14869_1005.n4 a_14869_1005.n0 75.271
R3291 a_14869_1005.n3 a_14869_1005.n2 75.214
R3292 a_14869_1005.n5 a_14869_1005.n4 36.517
R3293 a_14869_1005.n3 a_14869_1005.t7 14.338
R3294 a_14869_1005.n1 a_14869_1005.t5 14.282
R3295 a_14869_1005.n1 a_14869_1005.t4 14.282
R3296 a_14869_1005.n0 a_14869_1005.t0 14.282
R3297 a_14869_1005.n0 a_14869_1005.t1 14.282
R3298 a_14869_1005.t3 a_14869_1005.n5 14.282
R3299 a_14869_1005.n5 a_14869_1005.t2 14.282
R3300 a_14869_1005.n2 a_14869_1005.n1 12.119
R3301 a_1265_943.n6 a_1265_943.t10 454.685
R3302 a_1265_943.n8 a_1265_943.t13 454.685
R3303 a_1265_943.n4 a_1265_943.t6 454.685
R3304 a_1265_943.n6 a_1265_943.t5 428.979
R3305 a_1265_943.n8 a_1265_943.t9 428.979
R3306 a_1265_943.n4 a_1265_943.t8 428.979
R3307 a_1265_943.n7 a_1265_943.t11 248.006
R3308 a_1265_943.n9 a_1265_943.t12 248.006
R3309 a_1265_943.n5 a_1265_943.t7 248.006
R3310 a_1265_943.n14 a_1265_943.n12 220.639
R3311 a_1265_943.n12 a_1265_943.n3 135.994
R3312 a_1265_943.n7 a_1265_943.n6 81.941
R3313 a_1265_943.n9 a_1265_943.n8 81.941
R3314 a_1265_943.n5 a_1265_943.n4 81.941
R3315 a_1265_943.n11 a_1265_943.n5 81.396
R3316 a_1265_943.n10 a_1265_943.n9 79.491
R3317 a_1265_943.n3 a_1265_943.n2 76.002
R3318 a_1265_943.n10 a_1265_943.n7 76
R3319 a_1265_943.n12 a_1265_943.n11 76
R3320 a_1265_943.n14 a_1265_943.n13 30
R3321 a_1265_943.n15 a_1265_943.n0 24.383
R3322 a_1265_943.n15 a_1265_943.n14 23.684
R3323 a_1265_943.n1 a_1265_943.t3 14.282
R3324 a_1265_943.n1 a_1265_943.t2 14.282
R3325 a_1265_943.n2 a_1265_943.t0 14.282
R3326 a_1265_943.n2 a_1265_943.t4 14.282
R3327 a_1265_943.n3 a_1265_943.n1 12.85
R3328 a_1265_943.n11 a_1265_943.n10 2.947
R3329 a_1905_1004.n6 a_1905_1004.t8 480.392
R3330 a_1905_1004.n6 a_1905_1004.t9 403.272
R3331 a_1905_1004.n8 a_1905_1004.n5 233.952
R3332 a_1905_1004.n7 a_1905_1004.t7 213.869
R3333 a_1905_1004.n7 a_1905_1004.n6 161.6
R3334 a_1905_1004.n8 a_1905_1004.n7 153.315
R3335 a_1905_1004.n10 a_1905_1004.n8 143.492
R3336 a_1905_1004.n4 a_1905_1004.n3 79.232
R3337 a_1905_1004.n5 a_1905_1004.n4 63.152
R3338 a_1905_1004.n10 a_1905_1004.n9 30
R3339 a_1905_1004.n11 a_1905_1004.n0 24.383
R3340 a_1905_1004.n11 a_1905_1004.n10 23.684
R3341 a_1905_1004.n5 a_1905_1004.n1 16.08
R3342 a_1905_1004.n4 a_1905_1004.n2 16.08
R3343 a_1905_1004.n1 a_1905_1004.t6 14.282
R3344 a_1905_1004.n1 a_1905_1004.t5 14.282
R3345 a_1905_1004.n2 a_1905_1004.t2 14.282
R3346 a_1905_1004.n2 a_1905_1004.t3 14.282
R3347 a_1905_1004.n3 a_1905_1004.t0 14.282
R3348 a_1905_1004.n3 a_1905_1004.t1 14.282
R3349 a_5101_1004.n6 a_5101_1004.t8 512.525
R3350 a_5101_1004.n4 a_5101_1004.t5 512.525
R3351 a_5101_1004.n6 a_5101_1004.t10 371.139
R3352 a_5101_1004.n4 a_5101_1004.t9 371.139
R3353 a_5101_1004.n7 a_5101_1004.n6 226.225
R3354 a_5101_1004.n5 a_5101_1004.n4 225.866
R3355 a_5101_1004.n5 a_5101_1004.t7 218.057
R3356 a_5101_1004.n7 a_5101_1004.t6 217.698
R3357 a_5101_1004.n9 a_5101_1004.n3 215.652
R3358 a_5101_1004.n11 a_5101_1004.n9 140.981
R3359 a_5101_1004.n8 a_5101_1004.n5 79.488
R3360 a_5101_1004.n9 a_5101_1004.n8 77.314
R3361 a_5101_1004.n3 a_5101_1004.n2 76.002
R3362 a_5101_1004.n8 a_5101_1004.n7 76
R3363 a_5101_1004.n11 a_5101_1004.n10 30
R3364 a_5101_1004.n12 a_5101_1004.n0 24.383
R3365 a_5101_1004.n12 a_5101_1004.n11 23.684
R3366 a_5101_1004.n1 a_5101_1004.t2 14.282
R3367 a_5101_1004.n1 a_5101_1004.t1 14.282
R3368 a_5101_1004.n2 a_5101_1004.t4 14.282
R3369 a_5101_1004.n2 a_5101_1004.t3 14.282
R3370 a_5101_1004.n3 a_5101_1004.n1 12.85
R3371 a_10111_383.n6 a_10111_383.t12 480.392
R3372 a_10111_383.n8 a_10111_383.t11 472.359
R3373 a_10111_383.n6 a_10111_383.t9 403.272
R3374 a_10111_383.n8 a_10111_383.t7 384.527
R3375 a_10111_383.n7 a_10111_383.t10 320.08
R3376 a_10111_383.n9 a_10111_383.t8 277.772
R3377 a_10111_383.n13 a_10111_383.n11 249.364
R3378 a_10111_383.n11 a_10111_383.n5 127.401
R3379 a_10111_383.n10 a_10111_383.n7 83.304
R3380 a_10111_383.n10 a_10111_383.n9 80.032
R3381 a_10111_383.n4 a_10111_383.n3 79.232
R3382 a_10111_383.n11 a_10111_383.n10 76
R3383 a_10111_383.n9 a_10111_383.n8 67.001
R3384 a_10111_383.n5 a_10111_383.n4 63.152
R3385 a_10111_383.n7 a_10111_383.n6 55.388
R3386 a_10111_383.n13 a_10111_383.n12 30
R3387 a_10111_383.n14 a_10111_383.n0 24.383
R3388 a_10111_383.n14 a_10111_383.n13 23.684
R3389 a_10111_383.n5 a_10111_383.n1 16.08
R3390 a_10111_383.n4 a_10111_383.n2 16.08
R3391 a_10111_383.n1 a_10111_383.t6 14.282
R3392 a_10111_383.n1 a_10111_383.t5 14.282
R3393 a_10111_383.n2 a_10111_383.t2 14.282
R3394 a_10111_383.n2 a_10111_383.t3 14.282
R3395 a_10111_383.n3 a_10111_383.t1 14.282
R3396 a_10111_383.n3 a_10111_383.t0 14.282
R3397 a_9985_1004.n5 a_9985_1004.t9 512.525
R3398 a_9985_1004.n3 a_9985_1004.t7 512.525
R3399 a_9985_1004.n5 a_9985_1004.t5 371.139
R3400 a_9985_1004.n3 a_9985_1004.t10 371.139
R3401 a_9985_1004.n6 a_9985_1004.n5 226.225
R3402 a_9985_1004.n4 a_9985_1004.n3 225.866
R3403 a_9985_1004.n4 a_9985_1004.t8 218.057
R3404 a_9985_1004.n6 a_9985_1004.t6 217.698
R3405 a_9985_1004.n8 a_9985_1004.n2 215.652
R3406 a_9985_1004.n10 a_9985_1004.n8 147.503
R3407 a_9985_1004.n7 a_9985_1004.n4 79.488
R3408 a_9985_1004.n8 a_9985_1004.n7 77.314
R3409 a_9985_1004.n2 a_9985_1004.n1 76.002
R3410 a_9985_1004.n7 a_9985_1004.n6 76
R3411 a_9985_1004.n10 a_9985_1004.n9 15.218
R3412 a_9985_1004.n0 a_9985_1004.t3 14.282
R3413 a_9985_1004.n0 a_9985_1004.t4 14.282
R3414 a_9985_1004.n1 a_9985_1004.t1 14.282
R3415 a_9985_1004.n1 a_9985_1004.t0 14.282
R3416 a_9985_1004.n2 a_9985_1004.n0 12.85
R3417 a_9985_1004.n11 a_9985_1004.n10 12.014
R3418 a_12470_73.n12 a_12470_73.n11 26.811
R3419 a_12470_73.n6 a_12470_73.n5 24.977
R3420 a_12470_73.n2 a_12470_73.n1 24.877
R3421 a_12470_73.t0 a_12470_73.n2 12.677
R3422 a_12470_73.t0 a_12470_73.n3 11.595
R3423 a_12470_73.t1 a_12470_73.n8 8.137
R3424 a_12470_73.t0 a_12470_73.n4 7.273
R3425 a_12470_73.t0 a_12470_73.n0 6.109
R3426 a_12470_73.t1 a_12470_73.n7 4.864
R3427 a_12470_73.t0 a_12470_73.n12 2.074
R3428 a_12470_73.n7 a_12470_73.n6 1.13
R3429 a_12470_73.n12 a_12470_73.t1 0.937
R3430 a_12470_73.t1 a_12470_73.n10 0.804
R3431 a_12470_73.n10 a_12470_73.n9 0.136
R3432 a_10806_182.n10 a_10806_182.n8 82.852
R3433 a_10806_182.n7 a_10806_182.n6 32.833
R3434 a_10806_182.n8 a_10806_182.t1 32.416
R3435 a_10806_182.n10 a_10806_182.n9 27.2
R3436 a_10806_182.n11 a_10806_182.n0 23.498
R3437 a_10806_182.n3 a_10806_182.n2 23.284
R3438 a_10806_182.n11 a_10806_182.n10 22.4
R3439 a_10806_182.n7 a_10806_182.n4 19.017
R3440 a_10806_182.n6 a_10806_182.n5 13.494
R3441 a_10806_182.t1 a_10806_182.n1 7.04
R3442 a_10806_182.t1 a_10806_182.n3 5.727
R3443 a_10806_182.n8 a_10806_182.n7 1.435
R3444 a_15430_73.n2 a_15430_73.n0 34.602
R3445 a_15430_73.n2 a_15430_73.n1 2.138
R3446 a_15430_73.t0 a_15430_73.n2 0.069
R3447 a_11673_1004.n6 a_11673_1004.t7 480.392
R3448 a_11673_1004.n6 a_11673_1004.t8 403.272
R3449 a_11673_1004.n8 a_11673_1004.n5 233.952
R3450 a_11673_1004.n7 a_11673_1004.t9 213.869
R3451 a_11673_1004.n7 a_11673_1004.n6 161.6
R3452 a_11673_1004.n8 a_11673_1004.n7 153.315
R3453 a_11673_1004.n10 a_11673_1004.n8 143.492
R3454 a_11673_1004.n4 a_11673_1004.n3 79.232
R3455 a_11673_1004.n5 a_11673_1004.n4 63.152
R3456 a_11673_1004.n10 a_11673_1004.n9 30
R3457 a_11673_1004.n11 a_11673_1004.n0 24.383
R3458 a_11673_1004.n11 a_11673_1004.n10 23.684
R3459 a_11673_1004.n5 a_11673_1004.n1 16.08
R3460 a_11673_1004.n4 a_11673_1004.n2 16.08
R3461 a_11673_1004.n1 a_11673_1004.t6 14.282
R3462 a_11673_1004.n1 a_11673_1004.t5 14.282
R3463 a_11673_1004.n2 a_11673_1004.t3 14.282
R3464 a_11673_1004.n2 a_11673_1004.t2 14.282
R3465 a_11673_1004.n3 a_11673_1004.t1 14.282
R3466 a_11673_1004.n3 a_11673_1004.t0 14.282
R3467 a_13781_75.n1 a_13781_75.n0 25.576
R3468 a_13781_75.n3 a_13781_75.n2 9.111
R3469 a_13781_75.n7 a_13781_75.n5 7.859
R3470 a_13781_75.t0 a_13781_75.n7 3.034
R3471 a_13781_75.n5 a_13781_75.n3 1.964
R3472 a_13781_75.n5 a_13781_75.n4 1.964
R3473 a_13781_75.t0 a_13781_75.n1 1.871
R3474 a_13781_75.n7 a_13781_75.n6 0.443
R3475 a_14062_182.n12 a_14062_182.n10 82.852
R3476 a_14062_182.n13 a_14062_182.n0 49.6
R3477 a_14062_182.t1 a_14062_182.n2 46.91
R3478 a_14062_182.n7 a_14062_182.n5 34.805
R3479 a_14062_182.n7 a_14062_182.n6 32.622
R3480 a_14062_182.n10 a_14062_182.t1 32.416
R3481 a_14062_182.n12 a_14062_182.n11 27.2
R3482 a_14062_182.n13 a_14062_182.n12 22.4
R3483 a_14062_182.n9 a_14062_182.n7 19.017
R3484 a_14062_182.n2 a_14062_182.n1 17.006
R3485 a_14062_182.n5 a_14062_182.n4 7.5
R3486 a_14062_182.n9 a_14062_182.n8 7.5
R3487 a_14062_182.t1 a_14062_182.n3 7.04
R3488 a_14062_182.n10 a_14062_182.n9 1.435
R3489 a_13241_1004.n3 a_13241_1004.t6 512.525
R3490 a_13241_1004.n3 a_13241_1004.t7 371.139
R3491 a_13241_1004.n4 a_13241_1004.t5 368.806
R3492 a_13241_1004.n7 a_13241_1004.n5 306.82
R3493 a_13241_1004.n5 a_13241_1004.n4 134.297
R3494 a_13241_1004.n2 a_13241_1004.n1 76.002
R3495 a_13241_1004.n4 a_13241_1004.n3 74.076
R3496 a_13241_1004.n5 a_13241_1004.n2 56.335
R3497 a_13241_1004.n7 a_13241_1004.n6 15.218
R3498 a_13241_1004.n0 a_13241_1004.t3 14.282
R3499 a_13241_1004.n0 a_13241_1004.t4 14.282
R3500 a_13241_1004.n1 a_13241_1004.t0 14.282
R3501 a_13241_1004.n1 a_13241_1004.t1 14.282
R3502 a_13241_1004.n2 a_13241_1004.n0 12.85
R3503 a_13241_1004.n8 a_13241_1004.n7 12.014
R3504 a_757_75.n4 a_757_75.n3 19.724
R3505 a_757_75.t0 a_757_75.n5 11.595
R3506 a_757_75.t0 a_757_75.n4 9.207
R3507 a_757_75.n2 a_757_75.n0 8.543
R3508 a_757_75.t0 a_757_75.n2 3.034
R3509 a_757_75.n2 a_757_75.n1 0.443
R3510 a_1038_182.n12 a_1038_182.n10 82.852
R3511 a_1038_182.n13 a_1038_182.n0 49.6
R3512 a_1038_182.t1 a_1038_182.n2 46.91
R3513 a_1038_182.n7 a_1038_182.n5 34.805
R3514 a_1038_182.n7 a_1038_182.n6 32.622
R3515 a_1038_182.n10 a_1038_182.t1 32.416
R3516 a_1038_182.n12 a_1038_182.n11 27.2
R3517 a_1038_182.n13 a_1038_182.n12 22.4
R3518 a_1038_182.n9 a_1038_182.n7 19.017
R3519 a_1038_182.n2 a_1038_182.n1 17.006
R3520 a_1038_182.n5 a_1038_182.n4 7.5
R3521 a_1038_182.n9 a_1038_182.n8 7.5
R3522 a_1038_182.t1 a_1038_182.n3 7.04
R3523 a_1038_182.n10 a_1038_182.n9 1.435
R3524 a_2702_73.n12 a_2702_73.n11 26.811
R3525 a_2702_73.n6 a_2702_73.n5 24.977
R3526 a_2702_73.n2 a_2702_73.n1 24.877
R3527 a_2702_73.t0 a_2702_73.n2 12.677
R3528 a_2702_73.t0 a_2702_73.n3 11.595
R3529 a_2702_73.t1 a_2702_73.n8 8.137
R3530 a_2702_73.t0 a_2702_73.n4 7.273
R3531 a_2702_73.t0 a_2702_73.n0 6.109
R3532 a_2702_73.t1 a_2702_73.n7 4.864
R3533 a_2702_73.t0 a_2702_73.n12 2.074
R3534 a_2702_73.n7 a_2702_73.n6 1.13
R3535 a_2702_73.n12 a_2702_73.t1 0.937
R3536 a_2702_73.t1 a_2702_73.n10 0.804
R3537 a_2702_73.n10 a_2702_73.n9 0.136
R3538 a_13367_383.n8 a_13367_383.t15 512.525
R3539 a_13367_383.n6 a_13367_383.t7 477.179
R3540 a_13367_383.n11 a_13367_383.t14 472.359
R3541 a_13367_383.n6 a_13367_383.t11 406.485
R3542 a_13367_383.n11 a_13367_383.t8 384.527
R3543 a_13367_383.n8 a_13367_383.t10 371.139
R3544 a_13367_383.n7 a_13367_383.t13 346.633
R3545 a_13367_383.n9 a_13367_383.t9 340.206
R3546 a_13367_383.n12 a_13367_383.t12 304.325
R3547 a_13367_383.n16 a_13367_383.n14 276.257
R3548 a_13367_383.n14 a_13367_383.n5 101.187
R3549 a_13367_383.n9 a_13367_383.n8 89.615
R3550 a_13367_383.n13 a_13367_383.n12 80.035
R3551 a_13367_383.n4 a_13367_383.n3 79.232
R3552 a_13367_383.n10 a_13367_383.n7 78.675
R3553 a_13367_383.n10 a_13367_383.n9 76
R3554 a_13367_383.n14 a_13367_383.n13 76
R3555 a_13367_383.n5 a_13367_383.n4 63.152
R3556 a_13367_383.n17 a_13367_383.n0 55.263
R3557 a_13367_383.n12 a_13367_383.n11 40.448
R3558 a_13367_383.n16 a_13367_383.n15 30
R3559 a_13367_383.n7 a_13367_383.n6 29.194
R3560 a_13367_383.n17 a_13367_383.n16 23.684
R3561 a_13367_383.n5 a_13367_383.n1 16.08
R3562 a_13367_383.n4 a_13367_383.n2 16.08
R3563 a_13367_383.n1 a_13367_383.t6 14.282
R3564 a_13367_383.n1 a_13367_383.t5 14.282
R3565 a_13367_383.n2 a_13367_383.t1 14.282
R3566 a_13367_383.n2 a_13367_383.t0 14.282
R3567 a_13367_383.n3 a_13367_383.t3 14.282
R3568 a_13367_383.n3 a_13367_383.t2 14.282
R3569 a_13367_383.n13 a_13367_383.n10 1.043
R3570 a_13136_73.t0 a_13136_73.n1 34.62
R3571 a_13136_73.t0 a_13136_73.n0 8.137
R3572 a_13136_73.t0 a_13136_73.n2 4.69
R3573 a_343_383.n6 a_343_383.t12 480.392
R3574 a_343_383.n8 a_343_383.t7 472.359
R3575 a_343_383.n6 a_343_383.t9 403.272
R3576 a_343_383.n8 a_343_383.t10 384.527
R3577 a_343_383.n7 a_343_383.t11 320.08
R3578 a_343_383.n9 a_343_383.t8 277.772
R3579 a_343_383.n13 a_343_383.n11 249.364
R3580 a_343_383.n11 a_343_383.n5 127.401
R3581 a_343_383.n10 a_343_383.n7 83.304
R3582 a_343_383.n10 a_343_383.n9 80.032
R3583 a_343_383.n4 a_343_383.n3 79.232
R3584 a_343_383.n11 a_343_383.n10 76
R3585 a_343_383.n9 a_343_383.n8 67.001
R3586 a_343_383.n5 a_343_383.n4 63.152
R3587 a_343_383.n7 a_343_383.n6 55.388
R3588 a_343_383.n14 a_343_383.n0 55.263
R3589 a_343_383.n13 a_343_383.n12 30
R3590 a_343_383.n14 a_343_383.n13 23.684
R3591 a_343_383.n5 a_343_383.n1 16.08
R3592 a_343_383.n4 a_343_383.n2 16.08
R3593 a_343_383.n1 a_343_383.t6 14.282
R3594 a_343_383.n1 a_343_383.t5 14.282
R3595 a_343_383.n2 a_343_383.t3 14.282
R3596 a_343_383.n2 a_343_383.t2 14.282
R3597 a_343_383.n3 a_343_383.t1 14.282
R3598 a_343_383.n3 a_343_383.t0 14.282
R3599 a_8252_73.n12 a_8252_73.n11 26.811
R3600 a_8252_73.n6 a_8252_73.n5 24.977
R3601 a_8252_73.n2 a_8252_73.n1 24.877
R3602 a_8252_73.t0 a_8252_73.n2 12.677
R3603 a_8252_73.t0 a_8252_73.n3 11.595
R3604 a_8252_73.t1 a_8252_73.n8 8.137
R3605 a_8252_73.t0 a_8252_73.n4 7.273
R3606 a_8252_73.t0 a_8252_73.n0 6.109
R3607 a_8252_73.t1 a_8252_73.n7 4.864
R3608 a_8252_73.t0 a_8252_73.n12 2.074
R3609 a_8252_73.n7 a_8252_73.n6 1.13
R3610 a_8252_73.n12 a_8252_73.t1 0.937
R3611 a_8252_73.t1 a_8252_73.n10 0.804
R3612 a_8252_73.n10 a_8252_73.n9 0.136
R3613 a_16835_182.n2 a_16835_182.n0 362.371
R3614 a_16835_182.n2 a_16835_182.n1 15.218
R3615 a_16835_182.n0 a_16835_182.t1 14.282
R3616 a_16835_182.n0 a_16835_182.t0 14.282
R3617 a_16835_182.n3 a_16835_182.n2 12.014
R3618 a_112_73.t0 a_112_73.n1 34.62
R3619 a_112_73.t0 a_112_73.n0 8.137
R3620 a_112_73.t0 a_112_73.n2 4.69
R3621 a_3473_1004.n4 a_3473_1004.t6 512.525
R3622 a_3473_1004.n4 a_3473_1004.t7 371.139
R3623 a_3473_1004.n5 a_3473_1004.t5 324.268
R3624 a_3473_1004.n8 a_3473_1004.n6 247.192
R3625 a_3473_1004.n6 a_3473_1004.n5 153.315
R3626 a_3473_1004.n5 a_3473_1004.n4 119.654
R3627 a_3473_1004.n6 a_3473_1004.n3 109.441
R3628 a_3473_1004.n3 a_3473_1004.n2 76.002
R3629 a_3473_1004.n8 a_3473_1004.n7 30
R3630 a_3473_1004.n9 a_3473_1004.n0 24.383
R3631 a_3473_1004.n9 a_3473_1004.n8 23.684
R3632 a_3473_1004.n1 a_3473_1004.t2 14.282
R3633 a_3473_1004.n1 a_3473_1004.t3 14.282
R3634 a_3473_1004.n2 a_3473_1004.t0 14.282
R3635 a_3473_1004.n2 a_3473_1004.t1 14.282
R3636 a_3473_1004.n3 a_3473_1004.n1 12.85
R3637 a_5641_75.n1 a_5641_75.n0 25.576
R3638 a_5641_75.n3 a_5641_75.n2 9.111
R3639 a_5641_75.n7 a_5641_75.n5 7.859
R3640 a_5641_75.t0 a_5641_75.n7 3.034
R3641 a_5641_75.n5 a_5641_75.n3 1.964
R3642 a_5641_75.n5 a_5641_75.n4 1.964
R3643 a_5641_75.t0 a_5641_75.n1 1.871
R3644 a_5641_75.n7 a_5641_75.n6 0.443
R3645 a_4294_182.n10 a_4294_182.n8 82.852
R3646 a_4294_182.n7 a_4294_182.n6 32.833
R3647 a_4294_182.n8 a_4294_182.t1 32.416
R3648 a_4294_182.n10 a_4294_182.n9 27.2
R3649 a_4294_182.n11 a_4294_182.n0 23.498
R3650 a_4294_182.n3 a_4294_182.n2 23.284
R3651 a_4294_182.n11 a_4294_182.n10 22.4
R3652 a_4294_182.n7 a_4294_182.n4 19.017
R3653 a_4294_182.n6 a_4294_182.n5 13.494
R3654 a_4294_182.t1 a_4294_182.n1 7.04
R3655 a_4294_182.t1 a_4294_182.n3 5.727
R3656 a_4294_182.n8 a_4294_182.n7 1.435
R3657 a_11768_182.n10 a_11768_182.n8 82.852
R3658 a_11768_182.n7 a_11768_182.n6 32.833
R3659 a_11768_182.n8 a_11768_182.t1 32.416
R3660 a_11768_182.n10 a_11768_182.n9 27.2
R3661 a_11768_182.n11 a_11768_182.n0 23.498
R3662 a_11768_182.n3 a_11768_182.n2 23.284
R3663 a_11768_182.n11 a_11768_182.n10 22.4
R3664 a_11768_182.n7 a_11768_182.n4 19.017
R3665 a_11768_182.n6 a_11768_182.n5 13.494
R3666 a_11768_182.t1 a_11768_182.n1 7.04
R3667 a_11768_182.t1 a_11768_182.n3 5.727
R3668 a_11768_182.n8 a_11768_182.n7 1.435
R3669 a_2000_182.n10 a_2000_182.n8 82.852
R3670 a_2000_182.n11 a_2000_182.n0 49.6
R3671 a_2000_182.n7 a_2000_182.n6 32.833
R3672 a_2000_182.n8 a_2000_182.t1 32.416
R3673 a_2000_182.n10 a_2000_182.n9 27.2
R3674 a_2000_182.n3 a_2000_182.n2 23.284
R3675 a_2000_182.n11 a_2000_182.n10 22.4
R3676 a_2000_182.n7 a_2000_182.n4 19.017
R3677 a_2000_182.n6 a_2000_182.n5 13.494
R3678 a_2000_182.t1 a_2000_182.n1 7.04
R3679 a_2000_182.t1 a_2000_182.n3 5.727
R3680 a_2000_182.n8 a_2000_182.n7 1.435
R3681 a_3368_73.n12 a_3368_73.n11 26.811
R3682 a_3368_73.n6 a_3368_73.n5 24.977
R3683 a_3368_73.n2 a_3368_73.n1 24.877
R3684 a_3368_73.t0 a_3368_73.n2 12.677
R3685 a_3368_73.t0 a_3368_73.n3 11.595
R3686 a_3368_73.t1 a_3368_73.n8 8.137
R3687 a_3368_73.t0 a_3368_73.n4 7.273
R3688 a_3368_73.t0 a_3368_73.n0 6.109
R3689 a_3368_73.t1 a_3368_73.n7 4.864
R3690 a_3368_73.t0 a_3368_73.n12 2.074
R3691 a_3368_73.n7 a_3368_73.n6 1.13
R3692 a_3368_73.n12 a_3368_73.t1 0.937
R3693 a_3368_73.t1 a_3368_73.n10 0.804
R3694 a_3368_73.n10 a_3368_73.n9 0.136
R3695 a_14764_73.n13 a_14764_73.n12 26.811
R3696 a_14764_73.n6 a_14764_73.n5 24.977
R3697 a_14764_73.n2 a_14764_73.n1 24.877
R3698 a_14764_73.t0 a_14764_73.n2 12.677
R3699 a_14764_73.t0 a_14764_73.n3 11.595
R3700 a_14764_73.n11 a_14764_73.n10 8.561
R3701 a_14764_73.t0 a_14764_73.n4 7.273
R3702 a_14764_73.n9 a_14764_73.n8 7.066
R3703 a_14764_73.t0 a_14764_73.n0 6.109
R3704 a_14764_73.t1 a_14764_73.n7 4.864
R3705 a_14764_73.t0 a_14764_73.n13 2.074
R3706 a_14764_73.n7 a_14764_73.n6 1.13
R3707 a_14764_73.t1 a_14764_73.n11 0.958
R3708 a_14764_73.n13 a_14764_73.t1 0.937
R3709 a_14764_73.t1 a_14764_73.n9 0.86
R3710 a_6603_75.n1 a_6603_75.n0 25.576
R3711 a_6603_75.n3 a_6603_75.n2 9.111
R3712 a_6603_75.n7 a_6603_75.n6 2.455
R3713 a_6603_75.n5 a_6603_75.n3 1.964
R3714 a_6603_75.n5 a_6603_75.n4 1.964
R3715 a_6603_75.t0 a_6603_75.n1 1.871
R3716 a_6603_75.n7 a_6603_75.n5 0.636
R3717 a_6603_75.t0 a_6603_75.n7 0.246
R3718 a_4013_75.n5 a_4013_75.n4 19.724
R3719 a_4013_75.t0 a_4013_75.n3 11.595
R3720 a_4013_75.t0 a_4013_75.n5 9.207
R3721 a_4013_75.n2 a_4013_75.n1 2.455
R3722 a_4013_75.n2 a_4013_75.n0 1.32
R3723 a_4013_75.t0 a_4013_75.n2 0.246
R3724 a_5922_182.n8 a_5922_182.n6 96.467
R3725 a_5922_182.n3 a_5922_182.n1 44.628
R3726 a_5922_182.t0 a_5922_182.n8 32.417
R3727 a_5922_182.n3 a_5922_182.n2 23.284
R3728 a_5922_182.n6 a_5922_182.n5 22.349
R3729 a_5922_182.t0 a_5922_182.n10 20.241
R3730 a_5922_182.n10 a_5922_182.n9 13.494
R3731 a_5922_182.n6 a_5922_182.n4 8.443
R3732 a_5922_182.t0 a_5922_182.n0 8.137
R3733 a_5922_182.t0 a_5922_182.n3 5.727
R3734 a_5922_182.n8 a_5922_182.n7 1.435
R3735 a_7586_73.n12 a_7586_73.n11 26.811
R3736 a_7586_73.n6 a_7586_73.n5 24.977
R3737 a_7586_73.n2 a_7586_73.n1 24.877
R3738 a_7586_73.t0 a_7586_73.n2 12.677
R3739 a_7586_73.t0 a_7586_73.n3 11.595
R3740 a_7586_73.t1 a_7586_73.n8 8.137
R3741 a_7586_73.t0 a_7586_73.n4 7.273
R3742 a_7586_73.t0 a_7586_73.n0 6.109
R3743 a_7586_73.t1 a_7586_73.n7 4.864
R3744 a_7586_73.t0 a_7586_73.n12 2.074
R3745 a_7586_73.n7 a_7586_73.n6 1.13
R3746 a_7586_73.n12 a_7586_73.t1 0.937
R3747 a_7586_73.t1 a_7586_73.n10 0.804
R3748 a_7586_73.n10 a_7586_73.n9 0.136
R3749 a_10525_75.n5 a_10525_75.n4 19.724
R3750 a_10525_75.t0 a_10525_75.n3 11.595
R3751 a_10525_75.t0 a_10525_75.n5 9.207
R3752 a_10525_75.n2 a_10525_75.n1 2.455
R3753 a_10525_75.n2 a_10525_75.n0 1.32
R3754 a_10525_75.t0 a_10525_75.n2 0.246
R3755 a_16096_73.t0 a_16096_73.n1 34.62
R3756 a_16096_73.t0 a_16096_73.n0 8.137
R3757 a_16096_73.t0 a_16096_73.n2 4.69
R3758 a_4996_73.t0 a_4996_73.n1 34.62
R3759 a_4996_73.t0 a_4996_73.n0 8.137
R3760 a_4996_73.t0 a_4996_73.n2 4.69
R3761 a_9178_182.n9 a_9178_182.n7 82.852
R3762 a_9178_182.n3 a_9178_182.n1 44.628
R3763 a_9178_182.t0 a_9178_182.n9 32.417
R3764 a_9178_182.n7 a_9178_182.n6 27.2
R3765 a_9178_182.n5 a_9178_182.n4 23.498
R3766 a_9178_182.n3 a_9178_182.n2 23.284
R3767 a_9178_182.n7 a_9178_182.n5 22.4
R3768 a_9178_182.t0 a_9178_182.n11 20.241
R3769 a_9178_182.n11 a_9178_182.n10 13.494
R3770 a_9178_182.t0 a_9178_182.n0 8.137
R3771 a_9178_182.t0 a_9178_182.n3 5.727
R3772 a_9178_182.n9 a_9178_182.n8 1.435
R3773 a_11487_75.n5 a_11487_75.n4 19.724
R3774 a_11487_75.t0 a_11487_75.n3 11.595
R3775 a_11487_75.t0 a_11487_75.n5 9.207
R3776 a_11487_75.n2 a_11487_75.n1 2.455
R3777 a_11487_75.n2 a_11487_75.n0 1.32
R3778 a_11487_75.t0 a_11487_75.n2 0.246
R3779 a_8897_75.n5 a_8897_75.n4 19.724
R3780 a_8897_75.t0 a_8897_75.n3 11.595
R3781 a_8897_75.t0 a_8897_75.n5 9.207
R3782 a_8897_75.n2 a_8897_75.n1 2.455
R3783 a_8897_75.n2 a_8897_75.n0 1.32
R3784 a_8897_75.t0 a_8897_75.n2 0.246
C6 VPB VNB 63.92fF
C7 a_8897_75.n0 VNB 0.10fF
C8 a_8897_75.n1 VNB 0.04fF
C9 a_8897_75.n2 VNB 0.03fF
C10 a_8897_75.n3 VNB 0.07fF
C11 a_8897_75.n4 VNB 0.08fF
C12 a_8897_75.n5 VNB 0.06fF
C13 a_11487_75.n0 VNB 0.10fF
C14 a_11487_75.n1 VNB 0.04fF
C15 a_11487_75.n2 VNB 0.03fF
C16 a_11487_75.n3 VNB 0.07fF
C17 a_11487_75.n4 VNB 0.08fF
C18 a_11487_75.n5 VNB 0.06fF
C19 a_9178_182.n0 VNB 0.07fF
C20 a_9178_182.n1 VNB 0.09fF
C21 a_9178_182.n2 VNB 0.13fF
C22 a_9178_182.n3 VNB 0.11fF
C23 a_9178_182.n4 VNB 0.02fF
C24 a_9178_182.n5 VNB 0.03fF
C25 a_9178_182.n6 VNB 0.02fF
C26 a_9178_182.n7 VNB 0.05fF
C27 a_9178_182.n8 VNB 0.03fF
C28 a_9178_182.n9 VNB 0.11fF
C29 a_9178_182.n10 VNB 0.06fF
C30 a_9178_182.n11 VNB 0.01fF
C31 a_9178_182.t0 VNB 0.33fF
C32 a_4996_73.n0 VNB 0.05fF
C33 a_4996_73.n1 VNB 0.12fF
C34 a_4996_73.n2 VNB 0.04fF
C35 a_16096_73.n0 VNB 0.06fF
C36 a_16096_73.n1 VNB 0.13fF
C37 a_16096_73.n2 VNB 0.04fF
C38 a_10525_75.n0 VNB 0.10fF
C39 a_10525_75.n1 VNB 0.04fF
C40 a_10525_75.n2 VNB 0.03fF
C41 a_10525_75.n3 VNB 0.07fF
C42 a_10525_75.n4 VNB 0.08fF
C43 a_10525_75.n5 VNB 0.06fF
C44 a_7586_73.n0 VNB 0.02fF
C45 a_7586_73.n1 VNB 0.10fF
C46 a_7586_73.n2 VNB 0.06fF
C47 a_7586_73.n3 VNB 0.06fF
C48 a_7586_73.n4 VNB 0.00fF
C49 a_7586_73.n5 VNB 0.04fF
C50 a_7586_73.n6 VNB 0.05fF
C51 a_7586_73.n7 VNB 0.02fF
C52 a_7586_73.n8 VNB 0.05fF
C53 a_7586_73.n9 VNB 0.08fF
C54 a_7586_73.n10 VNB 0.17fF
C55 a_7586_73.t1 VNB 0.23fF
C56 a_7586_73.n11 VNB 0.09fF
C57 a_7586_73.n12 VNB 0.00fF
C58 a_5922_182.n0 VNB 0.07fF
C59 a_5922_182.n1 VNB 0.09fF
C60 a_5922_182.n2 VNB 0.13fF
C61 a_5922_182.n3 VNB 0.11fF
C62 a_5922_182.n4 VNB 0.02fF
C63 a_5922_182.n5 VNB 0.03fF
C64 a_5922_182.n6 VNB 0.06fF
C65 a_5922_182.n7 VNB 0.03fF
C66 a_5922_182.n8 VNB 0.12fF
C67 a_5922_182.n9 VNB 0.06fF
C68 a_5922_182.n10 VNB 0.01fF
C69 a_5922_182.t0 VNB 0.33fF
C70 a_4013_75.n0 VNB 0.10fF
C71 a_4013_75.n1 VNB 0.04fF
C72 a_4013_75.n2 VNB 0.03fF
C73 a_4013_75.n3 VNB 0.07fF
C74 a_4013_75.n4 VNB 0.08fF
C75 a_4013_75.n5 VNB 0.06fF
C76 a_6603_75.n0 VNB 0.09fF
C77 a_6603_75.n1 VNB 0.10fF
C78 a_6603_75.n2 VNB 0.05fF
C79 a_6603_75.n3 VNB 0.03fF
C80 a_6603_75.n4 VNB 0.04fF
C81 a_6603_75.n5 VNB 0.03fF
C82 a_6603_75.n6 VNB 0.04fF
C83 a_14764_73.n0 VNB 0.02fF
C84 a_14764_73.n1 VNB 0.09fF
C85 a_14764_73.n2 VNB 0.05fF
C86 a_14764_73.n3 VNB 0.06fF
C87 a_14764_73.n4 VNB 0.00fF
C88 a_14764_73.n5 VNB 0.04fF
C89 a_14764_73.n6 VNB 0.05fF
C90 a_14764_73.n7 VNB 0.02fF
C91 a_14764_73.n8 VNB 0.05fF
C92 a_14764_73.n9 VNB 0.09fF
C93 a_14764_73.n10 VNB 0.21fF
C94 a_14764_73.n11 VNB 0.07fF
C95 a_14764_73.t1 VNB 0.14fF
C96 a_14764_73.n12 VNB 0.04fF
C97 a_14764_73.n13 VNB 0.00fF
C98 a_3368_73.n0 VNB 0.02fF
C99 a_3368_73.n1 VNB 0.10fF
C100 a_3368_73.n2 VNB 0.06fF
C101 a_3368_73.n3 VNB 0.06fF
C102 a_3368_73.n4 VNB 0.00fF
C103 a_3368_73.n5 VNB 0.04fF
C104 a_3368_73.n6 VNB 0.05fF
C105 a_3368_73.n7 VNB 0.02fF
C106 a_3368_73.n8 VNB 0.05fF
C107 a_3368_73.n9 VNB 0.08fF
C108 a_3368_73.n10 VNB 0.17fF
C109 a_3368_73.t1 VNB 0.23fF
C110 a_3368_73.n11 VNB 0.09fF
C111 a_3368_73.n12 VNB 0.00fF
C112 a_2000_182.n0 VNB 0.02fF
C113 a_2000_182.n1 VNB 0.09fF
C114 a_2000_182.n2 VNB 0.13fF
C115 a_2000_182.n3 VNB 0.11fF
C116 a_2000_182.t1 VNB 0.30fF
C117 a_2000_182.n4 VNB 0.09fF
C118 a_2000_182.n5 VNB 0.06fF
C119 a_2000_182.n6 VNB 0.01fF
C120 a_2000_182.n7 VNB 0.03fF
C121 a_2000_182.n8 VNB 0.11fF
C122 a_2000_182.n9 VNB 0.02fF
C123 a_2000_182.n10 VNB 0.05fF
C124 a_2000_182.n11 VNB 0.02fF
C125 a_11768_182.n0 VNB 0.02fF
C126 a_11768_182.n1 VNB 0.09fF
C127 a_11768_182.n2 VNB 0.13fF
C128 a_11768_182.n3 VNB 0.11fF
C129 a_11768_182.t1 VNB 0.30fF
C130 a_11768_182.n4 VNB 0.09fF
C131 a_11768_182.n5 VNB 0.06fF
C132 a_11768_182.n6 VNB 0.01fF
C133 a_11768_182.n7 VNB 0.03fF
C134 a_11768_182.n8 VNB 0.11fF
C135 a_11768_182.n9 VNB 0.02fF
C136 a_11768_182.n10 VNB 0.05fF
C137 a_11768_182.n11 VNB 0.03fF
C138 a_4294_182.n0 VNB 0.02fF
C139 a_4294_182.n1 VNB 0.09fF
C140 a_4294_182.n2 VNB 0.13fF
C141 a_4294_182.n3 VNB 0.11fF
C142 a_4294_182.t1 VNB 0.30fF
C143 a_4294_182.n4 VNB 0.09fF
C144 a_4294_182.n5 VNB 0.06fF
C145 a_4294_182.n6 VNB 0.01fF
C146 a_4294_182.n7 VNB 0.03fF
C147 a_4294_182.n8 VNB 0.11fF
C148 a_4294_182.n9 VNB 0.02fF
C149 a_4294_182.n10 VNB 0.05fF
C150 a_4294_182.n11 VNB 0.03fF
C151 a_5641_75.n0 VNB 0.09fF
C152 a_5641_75.n1 VNB 0.10fF
C153 a_5641_75.n2 VNB 0.05fF
C154 a_5641_75.n3 VNB 0.03fF
C155 a_5641_75.n4 VNB 0.04fF
C156 a_5641_75.n5 VNB 0.11fF
C157 a_5641_75.n6 VNB 0.04fF
C158 a_3473_1004.n0 VNB 0.04fF
C159 a_3473_1004.n1 VNB 0.58fF
C160 a_3473_1004.n2 VNB 0.69fF
C161 a_3473_1004.n3 VNB 0.28fF
C162 a_3473_1004.n4 VNB 0.31fF
C163 a_3473_1004.n5 VNB 0.72fF
C164 a_3473_1004.n6 VNB 0.65fF
C165 a_3473_1004.n7 VNB 0.04fF
C166 a_3473_1004.n8 VNB 0.38fF
C167 a_3473_1004.n9 VNB 0.06fF
C168 a_112_73.n0 VNB 0.05fF
C169 a_112_73.n1 VNB 0.12fF
C170 a_112_73.n2 VNB 0.04fF
C171 a_16835_182.n0 VNB 1.03fF
C172 a_16835_182.n1 VNB 0.09fF
C173 a_16835_182.n2 VNB 0.49fF
C174 a_16835_182.n3 VNB 0.05fF
C175 a_8252_73.n0 VNB 0.02fF
C176 a_8252_73.n1 VNB 0.10fF
C177 a_8252_73.n2 VNB 0.06fF
C178 a_8252_73.n3 VNB 0.06fF
C179 a_8252_73.n4 VNB 0.00fF
C180 a_8252_73.n5 VNB 0.04fF
C181 a_8252_73.n6 VNB 0.05fF
C182 a_8252_73.n7 VNB 0.02fF
C183 a_8252_73.n8 VNB 0.05fF
C184 a_8252_73.n9 VNB 0.08fF
C185 a_8252_73.n10 VNB 0.17fF
C186 a_8252_73.t1 VNB 0.23fF
C187 a_8252_73.n11 VNB 0.09fF
C188 a_8252_73.n12 VNB 0.00fF
C189 a_343_383.n0 VNB 0.06fF
C190 a_343_383.n1 VNB 0.76fF
C191 a_343_383.n2 VNB 0.76fF
C192 a_343_383.n3 VNB 0.89fF
C193 a_343_383.n4 VNB 0.28fF
C194 a_343_383.n5 VNB 0.36fF
C195 a_343_383.n6 VNB 0.46fF
C196 a_343_383.n7 VNB 0.66fF
C197 a_343_383.n8 VNB 0.41fF
C198 a_343_383.t8 VNB 0.81fF
C199 a_343_383.n9 VNB 0.56fF
C200 a_343_383.n10 VNB 3.54fF
C201 a_343_383.n11 VNB 0.63fF
C202 a_343_383.n12 VNB 0.06fF
C203 a_343_383.n13 VNB 0.49fF
C204 a_343_383.n14 VNB 0.06fF
C205 a_13136_73.n0 VNB 0.05fF
C206 a_13136_73.n1 VNB 0.12fF
C207 a_13136_73.n2 VNB 0.04fF
C208 a_13367_383.n0 VNB 0.04fF
C209 a_13367_383.n1 VNB 0.51fF
C210 a_13367_383.n2 VNB 0.51fF
C211 a_13367_383.n3 VNB 0.60fF
C212 a_13367_383.n4 VNB 0.19fF
C213 a_13367_383.n5 VNB 0.21fF
C214 a_13367_383.n6 VNB 0.28fF
C215 a_13367_383.n7 VNB 0.39fF
C216 a_13367_383.n8 VNB 0.25fF
C217 a_13367_383.n9 VNB 0.45fF
C218 a_13367_383.n10 VNB 0.72fF
C219 a_13367_383.n11 VNB 0.25fF
C220 a_13367_383.t12 VNB 0.57fF
C221 a_13367_383.n12 VNB 0.38fF
C222 a_13367_383.n13 VNB 0.99fF
C223 a_13367_383.n14 VNB 0.42fF
C224 a_13367_383.n15 VNB 0.04fF
C225 a_13367_383.n16 VNB 0.36fF
C226 a_13367_383.n17 VNB 0.04fF
C227 a_2702_73.n0 VNB 0.02fF
C228 a_2702_73.n1 VNB 0.10fF
C229 a_2702_73.n2 VNB 0.06fF
C230 a_2702_73.n3 VNB 0.06fF
C231 a_2702_73.n4 VNB 0.00fF
C232 a_2702_73.n5 VNB 0.04fF
C233 a_2702_73.n6 VNB 0.05fF
C234 a_2702_73.n7 VNB 0.02fF
C235 a_2702_73.n8 VNB 0.05fF
C236 a_2702_73.n9 VNB 0.08fF
C237 a_2702_73.n10 VNB 0.17fF
C238 a_2702_73.t1 VNB 0.23fF
C239 a_2702_73.n11 VNB 0.09fF
C240 a_2702_73.n12 VNB 0.00fF
C241 a_1038_182.n0 VNB 0.02fF
C242 a_1038_182.n1 VNB 0.07fF
C243 a_1038_182.n2 VNB 0.13fF
C244 a_1038_182.n3 VNB 0.09fF
C245 a_1038_182.t1 VNB 0.25fF
C246 a_1038_182.n4 VNB 0.05fF
C247 a_1038_182.n5 VNB 0.06fF
C248 a_1038_182.n6 VNB 0.07fF
C249 a_1038_182.n7 VNB 0.07fF
C250 a_1038_182.n8 VNB 0.03fF
C251 a_1038_182.n9 VNB 0.01fF
C252 a_1038_182.n10 VNB 0.11fF
C253 a_1038_182.n11 VNB 0.02fF
C254 a_1038_182.n12 VNB 0.05fF
C255 a_1038_182.n13 VNB 0.02fF
C256 a_757_75.n0 VNB 0.20fF
C257 a_757_75.n1 VNB 0.04fF
C258 a_757_75.n2 VNB 0.01fF
C259 a_757_75.n3 VNB 0.08fF
C260 a_757_75.n4 VNB 0.06fF
C261 a_757_75.n5 VNB 0.07fF
C262 a_13241_1004.n0 VNB 0.52fF
C263 a_13241_1004.n1 VNB 0.61fF
C264 a_13241_1004.n2 VNB 0.19fF
C265 a_13241_1004.n3 VNB 0.22fF
C266 a_13241_1004.n4 VNB 0.69fF
C267 a_13241_1004.n5 VNB 0.57fF
C268 a_13241_1004.n6 VNB 0.08fF
C269 a_13241_1004.n7 VNB 0.39fF
C270 a_13241_1004.n8 VNB 0.04fF
C271 a_14062_182.n0 VNB 0.02fF
C272 a_14062_182.n1 VNB 0.07fF
C273 a_14062_182.n2 VNB 0.13fF
C274 a_14062_182.n3 VNB 0.09fF
C275 a_14062_182.t1 VNB 0.25fF
C276 a_14062_182.n4 VNB 0.05fF
C277 a_14062_182.n5 VNB 0.06fF
C278 a_14062_182.n6 VNB 0.07fF
C279 a_14062_182.n7 VNB 0.07fF
C280 a_14062_182.n8 VNB 0.03fF
C281 a_14062_182.n9 VNB 0.01fF
C282 a_14062_182.n10 VNB 0.11fF
C283 a_14062_182.n11 VNB 0.02fF
C284 a_14062_182.n12 VNB 0.05fF
C285 a_14062_182.n13 VNB 0.02fF
C286 a_13781_75.n0 VNB 0.09fF
C287 a_13781_75.n1 VNB 0.10fF
C288 a_13781_75.n2 VNB 0.05fF
C289 a_13781_75.n3 VNB 0.03fF
C290 a_13781_75.n4 VNB 0.04fF
C291 a_13781_75.n5 VNB 0.11fF
C292 a_13781_75.n6 VNB 0.04fF
C293 a_11673_1004.n0 VNB 0.04fF
C294 a_11673_1004.n1 VNB 0.56fF
C295 a_11673_1004.n2 VNB 0.56fF
C296 a_11673_1004.n3 VNB 0.65fF
C297 a_11673_1004.n4 VNB 0.21fF
C298 a_11673_1004.n5 VNB 0.39fF
C299 a_11673_1004.n6 VNB 0.46fF
C300 a_11673_1004.n7 VNB 0.57fF
C301 a_11673_1004.n8 VNB 0.65fF
C302 a_11673_1004.n9 VNB 0.04fF
C303 a_11673_1004.n10 VNB 0.23fF
C304 a_11673_1004.n11 VNB 0.06fF
C305 a_15430_73.n0 VNB 0.13fF
C306 a_15430_73.n1 VNB 0.13fF
C307 a_15430_73.n2 VNB 0.14fF
C308 a_10806_182.n0 VNB 0.02fF
C309 a_10806_182.n1 VNB 0.09fF
C310 a_10806_182.n2 VNB 0.13fF
C311 a_10806_182.n3 VNB 0.11fF
C312 a_10806_182.t1 VNB 0.30fF
C313 a_10806_182.n4 VNB 0.09fF
C314 a_10806_182.n5 VNB 0.06fF
C315 a_10806_182.n6 VNB 0.01fF
C316 a_10806_182.n7 VNB 0.03fF
C317 a_10806_182.n8 VNB 0.11fF
C318 a_10806_182.n9 VNB 0.02fF
C319 a_10806_182.n10 VNB 0.05fF
C320 a_10806_182.n11 VNB 0.03fF
C321 a_12470_73.n0 VNB 0.02fF
C322 a_12470_73.n1 VNB 0.10fF
C323 a_12470_73.n2 VNB 0.06fF
C324 a_12470_73.n3 VNB 0.06fF
C325 a_12470_73.n4 VNB 0.00fF
C326 a_12470_73.n5 VNB 0.04fF
C327 a_12470_73.n6 VNB 0.05fF
C328 a_12470_73.n7 VNB 0.02fF
C329 a_12470_73.n8 VNB 0.05fF
C330 a_12470_73.n9 VNB 0.08fF
C331 a_12470_73.n10 VNB 0.17fF
C332 a_12470_73.t1 VNB 0.23fF
C333 a_12470_73.n11 VNB 0.09fF
C334 a_12470_73.n12 VNB 0.00fF
C335 a_9985_1004.n0 VNB 0.72fF
C336 a_9985_1004.n1 VNB 0.85fF
C337 a_9985_1004.n2 VNB 0.51fF
C338 a_9985_1004.n3 VNB 0.55fF
C339 a_9985_1004.n4 VNB 0.64fF
C340 a_9985_1004.n5 VNB 0.56fF
C341 a_9985_1004.n6 VNB 0.61fF
C342 a_9985_1004.n7 VNB 1.53fF
C343 a_9985_1004.n8 VNB 0.59fF
C344 a_9985_1004.n9 VNB 0.11fF
C345 a_9985_1004.n10 VNB 0.28fF
C346 a_9985_1004.n11 VNB 0.06fF
C347 a_10111_383.n0 VNB 0.06fF
C348 a_10111_383.n1 VNB 0.86fF
C349 a_10111_383.n2 VNB 0.86fF
C350 a_10111_383.n3 VNB 1.01fF
C351 a_10111_383.n4 VNB 0.32fF
C352 a_10111_383.n5 VNB 0.41fF
C353 a_10111_383.n6 VNB 0.52fF
C354 a_10111_383.n7 VNB 0.75fF
C355 a_10111_383.n8 VNB 0.46fF
C356 a_10111_383.t8 VNB 0.92fF
C357 a_10111_383.n9 VNB 0.64fF
C358 a_10111_383.n10 VNB 4.02fF
C359 a_10111_383.n11 VNB 0.72fF
C360 a_10111_383.n12 VNB 0.05fF
C361 a_10111_383.n13 VNB 0.55fF
C362 a_10111_383.n14 VNB 0.09fF
C363 a_5101_1004.n0 VNB 0.05fF
C364 a_5101_1004.n1 VNB 0.71fF
C365 a_5101_1004.n2 VNB 0.85fF
C366 a_5101_1004.n3 VNB 0.51fF
C367 a_5101_1004.n4 VNB 0.55fF
C368 a_5101_1004.n5 VNB 0.64fF
C369 a_5101_1004.n6 VNB 0.55fF
C370 a_5101_1004.n7 VNB 0.61fF
C371 a_5101_1004.n8 VNB 1.53fF
C372 a_5101_1004.n9 VNB 0.57fF
C373 a_5101_1004.n10 VNB 0.05fF
C374 a_5101_1004.n11 VNB 0.29fF
C375 a_5101_1004.n12 VNB 0.07fF
C376 a_1905_1004.n0 VNB 0.04fF
C377 a_1905_1004.n1 VNB 0.53fF
C378 a_1905_1004.n2 VNB 0.53fF
C379 a_1905_1004.n3 VNB 0.63fF
C380 a_1905_1004.n4 VNB 0.20fF
C381 a_1905_1004.n5 VNB 0.38fF
C382 a_1905_1004.n6 VNB 0.45fF
C383 a_1905_1004.n7 VNB 0.55fF
C384 a_1905_1004.n8 VNB 0.62fF
C385 a_1905_1004.n9 VNB 0.03fF
C386 a_1905_1004.n10 VNB 0.22fF
C387 a_1905_1004.n11 VNB 0.05fF
C388 a_1265_943.n0 VNB 0.06fF
C389 a_1265_943.n1 VNB 0.77fF
C390 a_1265_943.n2 VNB 0.91fF
C391 a_1265_943.n3 VNB 0.42fF
C392 a_1265_943.n4 VNB 0.52fF
C393 a_1265_943.t7 VNB 0.79fF
C394 a_1265_943.n5 VNB 0.59fF
C395 a_1265_943.n6 VNB 0.52fF
C396 a_1265_943.t11 VNB 0.79fF
C397 a_1265_943.n7 VNB 0.53fF
C398 a_1265_943.n8 VNB 0.52fF
C399 a_1265_943.t12 VNB 0.79fF
C400 a_1265_943.n9 VNB 0.55fF
C401 a_1265_943.n10 VNB 1.66fF
C402 a_1265_943.n11 VNB 2.24fF
C403 a_1265_943.n12 VNB 0.61fF
C404 a_1265_943.n13 VNB 0.05fF
C405 a_1265_943.n14 VNB 0.45fF
C406 a_1265_943.n15 VNB 0.08fF
C407 a_14869_1005.n0 VNB 0.41fF
C408 a_14869_1005.n1 VNB 0.33fF
C409 a_14869_1005.n2 VNB 0.23fF
C410 a_14869_1005.n3 VNB 0.63fF
C411 a_14869_1005.n4 VNB 0.28fF
C412 a_14869_1005.n5 VNB 0.37fF
C413 a_1719_75.n0 VNB 0.20fF
C414 a_1719_75.n1 VNB 0.04fF
C415 a_1719_75.n2 VNB 0.01fF
C416 a_1719_75.n3 VNB 0.08fF
C417 a_1719_75.n4 VNB 0.06fF
C418 a_1719_75.n5 VNB 0.07fF
C419 a_217_1004.n0 VNB 0.54fF
C420 a_217_1004.n1 VNB 0.64fF
C421 a_217_1004.n2 VNB 0.38fF
C422 a_217_1004.n3 VNB 0.42fF
C423 a_217_1004.n4 VNB 0.48fF
C424 a_217_1004.n5 VNB 0.42fF
C425 a_217_1004.n6 VNB 0.46fF
C426 a_217_1004.n7 VNB 1.15fF
C427 a_217_1004.n8 VNB 0.44fF
C428 a_217_1004.n9 VNB 0.08fF
C429 a_217_1004.n10 VNB 0.21fF
C430 a_217_1004.n11 VNB 0.05fF
C431 a_9880_73.n0 VNB 0.05fF
C432 a_9880_73.n1 VNB 0.02fF
C433 a_9880_73.n2 VNB 0.12fF
C434 a_9880_73.n3 VNB 0.04fF
C435 a_9880_73.n4 VNB 0.17fF
C436 a_8483_383.n0 VNB 0.08fF
C437 a_8483_383.n1 VNB 1.01fF
C438 a_8483_383.n2 VNB 1.01fF
C439 a_8483_383.n3 VNB 1.18fF
C440 a_8483_383.n4 VNB 0.37fF
C441 a_8483_383.n5 VNB 0.48fF
C442 a_8483_383.n6 VNB 0.54fF
C443 a_8483_383.t11 VNB 1.07fF
C444 a_8483_383.n7 VNB 1.60fF
C445 a_8483_383.n8 VNB 1.41fF
C446 a_8483_383.n9 VNB 0.54fF
C447 a_8483_383.n10 VNB 0.61fF
C448 a_8483_383.t15 VNB 1.07fF
C449 a_8483_383.n11 VNB 1.81fF
C450 a_8483_383.n12 VNB 1.38fF
C451 a_8483_383.t9 VNB 0.92fF
C452 a_8483_383.n13 VNB 4.79fF
C453 a_8483_383.n14 VNB 4.81fF
C454 a_8483_383.n15 VNB 0.06fF
C455 a_8483_383.n16 VNB 0.41fF
C456 a_8483_383.n17 VNB 0.10fF
C457 a_8357_1004.n0 VNB 0.60fF
C458 a_8357_1004.n1 VNB 0.71fF
C459 a_8357_1004.n2 VNB 0.43fF
C460 a_8357_1004.n3 VNB 0.46fF
C461 a_8357_1004.n4 VNB 0.71fF
C462 a_8357_1004.n5 VNB 0.69fF
C463 a_8357_1004.n6 VNB 0.09fF
C464 a_8357_1004.n7 VNB 0.23fF
C465 a_8357_1004.n8 VNB 0.05fF
C466 a_11033_943.n0 VNB 0.07fF
C467 a_11033_943.n1 VNB 0.88fF
C468 a_11033_943.n2 VNB 1.04fF
C469 a_11033_943.n3 VNB 0.48fF
C470 a_11033_943.n4 VNB 0.59fF
C471 a_11033_943.t12 VNB 0.90fF
C472 a_11033_943.n5 VNB 0.67fF
C473 a_11033_943.n6 VNB 0.59fF
C474 a_11033_943.t8 VNB 0.90fF
C475 a_11033_943.n7 VNB 0.60fF
C476 a_11033_943.n8 VNB 0.59fF
C477 a_11033_943.t5 VNB 0.90fF
C478 a_11033_943.n9 VNB 0.63fF
C479 a_11033_943.n10 VNB 1.89fF
C480 a_11033_943.n11 VNB 2.55fF
C481 a_11033_943.n12 VNB 0.69fF
C482 a_11033_943.n13 VNB 0.06fF
C483 a_11033_943.n14 VNB 0.51fF
C484 a_11033_943.n15 VNB 0.09fF
C485 a_15533_1005.n0 VNB 0.28fF
C486 a_15533_1005.n1 VNB 0.36fF
C487 a_15533_1005.n2 VNB 0.25fF
C488 a_15533_1005.n3 VNB 0.58fF
C489 a_15533_1005.n4 VNB 0.21fF
C490 a_15533_1005.n5 VNB 0.29fF
C491 a_15044_181.n0 VNB 0.05fF
C492 a_15044_181.n1 VNB 0.38fF
C493 a_15044_181.n2 VNB 0.46fF
C494 a_15044_181.n3 VNB 0.22fF
C495 a_15044_181.n4 VNB 0.24fF
C496 a_15044_181.t8 VNB 0.48fF
C497 a_15044_181.n5 VNB 0.49fF
C498 a_15044_181.n6 VNB 0.45fF
C499 a_15044_181.n7 VNB 0.03fF
C500 a_15044_181.n8 VNB 0.05fF
C501 a_15044_181.n9 VNB 0.03fF
C502 a_15044_181.n10 VNB 0.09fF
C503 a_15044_181.n11 VNB 0.03fF
C504 a_15044_181.n12 VNB 0.05fF
C505 a_15044_181.n13 VNB 0.02fF
C506 a_15044_181.n14 VNB 0.09fF
C507 a_15044_181.n15 VNB 0.98fF
C508 a_15044_181.n16 VNB 0.27fF
C509 a_15044_181.n17 VNB 0.02fF
C510 a_15044_181.n18 VNB 0.05fF
C511 a_15044_181.n19 VNB 0.04fF
C512 a_3599_383.n0 VNB 0.10fF
C513 a_3599_383.n1 VNB 1.27fF
C514 a_3599_383.n2 VNB 1.27fF
C515 a_3599_383.n3 VNB 1.49fF
C516 a_3599_383.n4 VNB 0.47fF
C517 a_3599_383.n5 VNB 0.75fF
C518 a_3599_383.n6 VNB 0.85fF
C519 a_3599_383.n7 VNB 1.10fF
C520 a_3599_383.n8 VNB 1.35fF
C521 a_3599_383.t9 VNB 1.03fF
C522 a_3599_383.n9 VNB 0.88fF
C523 a_3599_383.n10 VNB 4.46fF
C524 a_3599_383.n11 VNB 0.82fF
C525 a_3599_383.t11 VNB 1.21fF
C526 a_3599_383.n12 VNB 0.93fF
C527 a_3599_383.n13 VNB 19.81fF
C528 a_3599_383.n14 VNB 1.04fF
C529 a_3599_383.n15 VNB 0.10fF
C530 a_3599_383.n16 VNB 0.66fF
C531 a_3599_383.n17 VNB 0.11fF
C532 VPB.n0 VNB 0.03fF
C533 VPB.n1 VNB 0.04fF
C534 VPB.n2 VNB 0.02fF
C535 VPB.n3 VNB 0.14fF
C536 VPB.n5 VNB 0.02fF
C537 VPB.n6 VNB 0.02fF
C538 VPB.n7 VNB 0.02fF
C539 VPB.n8 VNB 0.02fF
C540 VPB.n10 VNB 0.02fF
C541 VPB.n11 VNB 0.02fF
C542 VPB.n12 VNB 0.02fF
C543 VPB.n14 VNB 0.10fF
C544 VPB.n15 VNB 0.02fF
C545 VPB.n16 VNB 0.02fF
C546 VPB.n17 VNB 0.02fF
C547 VPB.n18 VNB 0.04fF
C548 VPB.n19 VNB 0.02fF
C549 VPB.n20 VNB 0.25fF
C550 VPB.n21 VNB 0.04fF
C551 VPB.n23 VNB 0.02fF
C552 VPB.n24 VNB 0.02fF
C553 VPB.n25 VNB 0.02fF
C554 VPB.n26 VNB 0.02fF
C555 VPB.n28 VNB 0.02fF
C556 VPB.n29 VNB 0.02fF
C557 VPB.n30 VNB 0.02fF
C558 VPB.n32 VNB 0.28fF
C559 VPB.n34 VNB 0.03fF
C560 VPB.n35 VNB 0.02fF
C561 VPB.n36 VNB 0.21fF
C562 VPB.n37 VNB 0.02fF
C563 VPB.n38 VNB 0.01fF
C564 VPB.n39 VNB 0.06fF
C565 VPB.n40 VNB 0.28fF
C566 VPB.n41 VNB 0.02fF
C567 VPB.n42 VNB 0.02fF
C568 VPB.n43 VNB 0.28fF
C569 VPB.n44 VNB 0.01fF
C570 VPB.n45 VNB 0.02fF
C571 VPB.n46 VNB 0.03fF
C572 VPB.n47 VNB 0.03fF
C573 VPB.n48 VNB 0.28fF
C574 VPB.n49 VNB 0.01fF
C575 VPB.n50 VNB 0.02fF
C576 VPB.n51 VNB 0.23fF
C577 VPB.n52 VNB 0.02fF
C578 VPB.n53 VNB 0.01fF
C579 VPB.n54 VNB 0.05fF
C580 VPB.n55 VNB 0.14fF
C581 VPB.n56 VNB 0.16fF
C582 VPB.n57 VNB 0.02fF
C583 VPB.n58 VNB 0.02fF
C584 VPB.n59 VNB 0.14fF
C585 VPB.n60 VNB 0.15fF
C586 VPB.n61 VNB 0.02fF
C587 VPB.n62 VNB 0.02fF
C588 VPB.n63 VNB 0.02fF
C589 VPB.n64 VNB 0.14fF
C590 VPB.n65 VNB 0.15fF
C591 VPB.n66 VNB 0.02fF
C592 VPB.n67 VNB 0.02fF
C593 VPB.n68 VNB 0.14fF
C594 VPB.n69 VNB 0.16fF
C595 VPB.n70 VNB 0.02fF
C596 VPB.n71 VNB 0.02fF
C597 VPB.n72 VNB 0.06fF
C598 VPB.n73 VNB 0.24fF
C599 VPB.n74 VNB 0.02fF
C600 VPB.n75 VNB 0.01fF
C601 VPB.n76 VNB 0.02fF
C602 VPB.n77 VNB 0.02fF
C603 VPB.n78 VNB 0.02fF
C604 VPB.n79 VNB 0.04fF
C605 VPB.n80 VNB 0.02fF
C606 VPB.n81 VNB 0.24fF
C607 VPB.n82 VNB 0.04fF
C608 VPB.n84 VNB 0.02fF
C609 VPB.n85 VNB 0.02fF
C610 VPB.n86 VNB 0.02fF
C611 VPB.n87 VNB 0.02fF
C612 VPB.n89 VNB 0.02fF
C613 VPB.n90 VNB 0.02fF
C614 VPB.n91 VNB 0.02fF
C615 VPB.n93 VNB 0.28fF
C616 VPB.n95 VNB 0.03fF
C617 VPB.n96 VNB 0.02fF
C618 VPB.n97 VNB 0.10fF
C619 VPB.n98 VNB 0.10fF
C620 VPB.n99 VNB 0.14fF
C621 VPB.n100 VNB 0.16fF
C622 VPB.n101 VNB 0.02fF
C623 VPB.n102 VNB 0.02fF
C624 VPB.n103 VNB 0.02fF
C625 VPB.n104 VNB 0.14fF
C626 VPB.n105 VNB 0.15fF
C627 VPB.n106 VNB 0.02fF
C628 VPB.n107 VNB 0.02fF
C629 VPB.n108 VNB 0.14fF
C630 VPB.n109 VNB 0.15fF
C631 VPB.n110 VNB 0.02fF
C632 VPB.n111 VNB 0.02fF
C633 VPB.n112 VNB 0.02fF
C634 VPB.n113 VNB 0.14fF
C635 VPB.n114 VNB 0.16fF
C636 VPB.n115 VNB 0.02fF
C637 VPB.n116 VNB 0.02fF
C638 VPB.n117 VNB 0.14fF
C639 VPB.n118 VNB 0.16fF
C640 VPB.n119 VNB 0.02fF
C641 VPB.n120 VNB 0.02fF
C642 VPB.n121 VNB 0.21fF
C643 VPB.n122 VNB 0.02fF
C644 VPB.n123 VNB 0.01fF
C645 VPB.n124 VNB 0.06fF
C646 VPB.n125 VNB 0.28fF
C647 VPB.n126 VNB 0.02fF
C648 VPB.n127 VNB 0.02fF
C649 VPB.n128 VNB 0.28fF
C650 VPB.n129 VNB 0.01fF
C651 VPB.n130 VNB 0.02fF
C652 VPB.n131 VNB 0.03fF
C653 VPB.n132 VNB 0.03fF
C654 VPB.n133 VNB 0.28fF
C655 VPB.n134 VNB 0.01fF
C656 VPB.n135 VNB 0.02fF
C657 VPB.n136 VNB 0.23fF
C658 VPB.n137 VNB 0.02fF
C659 VPB.n138 VNB 0.01fF
C660 VPB.n139 VNB 0.05fF
C661 VPB.n140 VNB 0.02fF
C662 VPB.n141 VNB 0.02fF
C663 VPB.n142 VNB 0.02fF
C664 VPB.n143 VNB 0.11fF
C665 VPB.n144 VNB 0.03fF
C666 VPB.n145 VNB 0.02fF
C667 VPB.n146 VNB 0.05fF
C668 VPB.n147 VNB 0.01fF
C669 VPB.n149 VNB 0.02fF
C670 VPB.n150 VNB 0.02fF
C671 VPB.n151 VNB 0.02fF
C672 VPB.n152 VNB 0.02fF
C673 VPB.n154 VNB 0.02fF
C674 VPB.n157 VNB 0.46fF
C675 VPB.n159 VNB 0.04fF
C676 VPB.n160 VNB 0.04fF
C677 VPB.n161 VNB 0.28fF
C678 VPB.n162 VNB 0.03fF
C679 VPB.n163 VNB 0.03fF
C680 VPB.n164 VNB 0.06fF
C681 VPB.n165 VNB 0.14fF
C682 VPB.n166 VNB 0.19fF
C683 VPB.n167 VNB 0.02fF
C684 VPB.n168 VNB 0.01fF
C685 VPB.n169 VNB 0.07fF
C686 VPB.n170 VNB 0.16fF
C687 VPB.n171 VNB 0.02fF
C688 VPB.n172 VNB 0.02fF
C689 VPB.n173 VNB 0.02fF
C690 VPB.n174 VNB 0.06fF
C691 VPB.n175 VNB 0.14fF
C692 VPB.n176 VNB 0.20fF
C693 VPB.n177 VNB 0.02fF
C694 VPB.n178 VNB 0.01fF
C695 VPB.n179 VNB 0.02fF
C696 VPB.n180 VNB 0.28fF
C697 VPB.n181 VNB 0.01fF
C698 VPB.n182 VNB 0.02fF
C699 VPB.n183 VNB 0.04fF
C700 VPB.n184 VNB 0.02fF
C701 VPB.n185 VNB 0.02fF
C702 VPB.n186 VNB 0.02fF
C703 VPB.n187 VNB 0.04fF
C704 VPB.n188 VNB 0.02fF
C705 VPB.n189 VNB 0.17fF
C706 VPB.n190 VNB 0.04fF
C707 VPB.n192 VNB 0.02fF
C708 VPB.n193 VNB 0.02fF
C709 VPB.n194 VNB 0.02fF
C710 VPB.n195 VNB 0.02fF
C711 VPB.n197 VNB 0.02fF
C712 VPB.n198 VNB 0.02fF
C713 VPB.n199 VNB 0.02fF
C714 VPB.n201 VNB 0.28fF
C715 VPB.n203 VNB 0.03fF
C716 VPB.n204 VNB 0.02fF
C717 VPB.n205 VNB 0.03fF
C718 VPB.n206 VNB 0.03fF
C719 VPB.n207 VNB 0.28fF
C720 VPB.n208 VNB 0.01fF
C721 VPB.n209 VNB 0.02fF
C722 VPB.n210 VNB 0.04fF
C723 VPB.n211 VNB 0.28fF
C724 VPB.n212 VNB 0.02fF
C725 VPB.n213 VNB 0.02fF
C726 VPB.n214 VNB 0.02fF
C727 VPB.n215 VNB 0.28fF
C728 VPB.n216 VNB 0.02fF
C729 VPB.n217 VNB 0.02fF
C730 VPB.n218 VNB 0.02fF
C731 VPB.n219 VNB 0.28fF
C732 VPB.n220 VNB 0.02fF
C733 VPB.n221 VNB 0.02fF
C734 VPB.n222 VNB 0.02fF
C735 VPB.n223 VNB 0.28fF
C736 VPB.n224 VNB 0.02fF
C737 VPB.n225 VNB 0.02fF
C738 VPB.n226 VNB 0.02fF
C739 VPB.n227 VNB 0.28fF
C740 VPB.n228 VNB 0.02fF
C741 VPB.n229 VNB 0.02fF
C742 VPB.n230 VNB 0.02fF
C743 VPB.n231 VNB 0.28fF
C744 VPB.n232 VNB 0.02fF
C745 VPB.n233 VNB 0.02fF
C746 VPB.n234 VNB 0.02fF
C747 VPB.n235 VNB 0.28fF
C748 VPB.n236 VNB 0.01fF
C749 VPB.n237 VNB 0.02fF
C750 VPB.n238 VNB 0.04fF
C751 VPB.n239 VNB 0.02fF
C752 VPB.n240 VNB 0.02fF
C753 VPB.n241 VNB 0.02fF
C754 VPB.n242 VNB 0.04fF
C755 VPB.n243 VNB 0.02fF
C756 VPB.n244 VNB 0.20fF
C757 VPB.n245 VNB 0.04fF
C758 VPB.n247 VNB 0.02fF
C759 VPB.n248 VNB 0.02fF
C760 VPB.n249 VNB 0.02fF
C761 VPB.n250 VNB 0.02fF
C762 VPB.n252 VNB 0.02fF
C763 VPB.n253 VNB 0.02fF
C764 VPB.n254 VNB 0.02fF
C765 VPB.n256 VNB 0.28fF
C766 VPB.n258 VNB 0.03fF
C767 VPB.n259 VNB 0.02fF
C768 VPB.n260 VNB 0.03fF
C769 VPB.n261 VNB 0.03fF
C770 VPB.n262 VNB 0.28fF
C771 VPB.n263 VNB 0.01fF
C772 VPB.n264 VNB 0.02fF
C773 VPB.n265 VNB 0.04fF
C774 VPB.n266 VNB 0.28fF
C775 VPB.n267 VNB 0.02fF
C776 VPB.n268 VNB 0.02fF
C777 VPB.n269 VNB 0.02fF
C778 VPB.n270 VNB 0.28fF
C779 VPB.n271 VNB 0.02fF
C780 VPB.n272 VNB 0.02fF
C781 VPB.n273 VNB 0.02fF
C782 VPB.n274 VNB 0.28fF
C783 VPB.n275 VNB 0.02fF
C784 VPB.n276 VNB 0.02fF
C785 VPB.n277 VNB 0.02fF
C786 VPB.n278 VNB 0.28fF
C787 VPB.n279 VNB 0.02fF
C788 VPB.n280 VNB 0.02fF
C789 VPB.n281 VNB 0.02fF
C790 VPB.n282 VNB 0.28fF
C791 VPB.n283 VNB 0.02fF
C792 VPB.n284 VNB 0.02fF
C793 VPB.n285 VNB 0.02fF
C794 VPB.n286 VNB 0.28fF
C795 VPB.n287 VNB 0.02fF
C796 VPB.n288 VNB 0.02fF
C797 VPB.n289 VNB 0.02fF
C798 VPB.n290 VNB 0.28fF
C799 VPB.n291 VNB 0.01fF
C800 VPB.n292 VNB 0.02fF
C801 VPB.n293 VNB 0.04fF
C802 VPB.n294 VNB 0.02fF
C803 VPB.n295 VNB 0.02fF
C804 VPB.n296 VNB 0.02fF
C805 VPB.n297 VNB 0.04fF
C806 VPB.n298 VNB 0.02fF
C807 VPB.n299 VNB 0.20fF
C808 VPB.n300 VNB 0.04fF
C809 VPB.n302 VNB 0.02fF
C810 VPB.n303 VNB 0.02fF
C811 VPB.n304 VNB 0.02fF
C812 VPB.n305 VNB 0.02fF
C813 VPB.n307 VNB 0.02fF
C814 VPB.n308 VNB 0.02fF
C815 VPB.n309 VNB 0.02fF
C816 VPB.n311 VNB 0.28fF
C817 VPB.n313 VNB 0.03fF
C818 VPB.n314 VNB 0.02fF
C819 VPB.n315 VNB 0.03fF
C820 VPB.n316 VNB 0.03fF
C821 VPB.n317 VNB 0.28fF
C822 VPB.n318 VNB 0.01fF
C823 VPB.n319 VNB 0.02fF
C824 VPB.n320 VNB 0.04fF
C825 VPB.n321 VNB 0.06fF
C826 VPB.n322 VNB 0.23fF
C827 VPB.n323 VNB 0.02fF
C828 VPB.n324 VNB 0.01fF
C829 VPB.n325 VNB 0.02fF
C830 VPB.n326 VNB 0.14fF
C831 VPB.n327 VNB 0.16fF
C832 VPB.n328 VNB 0.02fF
C833 VPB.n329 VNB 0.02fF
C834 VPB.n330 VNB 0.02fF
C835 VPB.n331 VNB 0.10fF
C836 VPB.n332 VNB 0.02fF
C837 VPB.n333 VNB 0.14fF
C838 VPB.n334 VNB 0.15fF
C839 VPB.n335 VNB 0.02fF
C840 VPB.n336 VNB 0.02fF
C841 VPB.n337 VNB 0.02fF
C842 VPB.n338 VNB 0.14fF
C843 VPB.n339 VNB 0.15fF
C844 VPB.n340 VNB 0.02fF
C845 VPB.n341 VNB 0.02fF
C846 VPB.n342 VNB 0.02fF
C847 VPB.n343 VNB 0.14fF
C848 VPB.n344 VNB 0.16fF
C849 VPB.n345 VNB 0.02fF
C850 VPB.n346 VNB 0.02fF
C851 VPB.n347 VNB 0.02fF
C852 VPB.n348 VNB 0.06fF
C853 VPB.n349 VNB 0.24fF
C854 VPB.n350 VNB 0.02fF
C855 VPB.n351 VNB 0.01fF
C856 VPB.n352 VNB 0.02fF
C857 VPB.n353 VNB 0.28fF
C858 VPB.n354 VNB 0.01fF
C859 VPB.n355 VNB 0.02fF
C860 VPB.n356 VNB 0.04fF
C861 VPB.n357 VNB 0.02fF
C862 VPB.n358 VNB 0.02fF
C863 VPB.n359 VNB 0.02fF
C864 VPB.n360 VNB 0.04fF
C865 VPB.n361 VNB 0.02fF
C866 VPB.n362 VNB 0.24fF
C867 VPB.n363 VNB 0.04fF
C868 VPB.n365 VNB 0.02fF
C869 VPB.n366 VNB 0.02fF
C870 VPB.n367 VNB 0.02fF
C871 VPB.n368 VNB 0.02fF
C872 VPB.n370 VNB 0.02fF
C873 VPB.n371 VNB 0.02fF
C874 VPB.n372 VNB 0.02fF
C875 VPB.n374 VNB 0.28fF
C876 VPB.n376 VNB 0.03fF
C877 VPB.n377 VNB 0.02fF
C878 VPB.n378 VNB 0.03fF
C879 VPB.n379 VNB 0.03fF
C880 VPB.n380 VNB 0.28fF
C881 VPB.n381 VNB 0.01fF
C882 VPB.n382 VNB 0.02fF
C883 VPB.n383 VNB 0.04fF
C884 VPB.n384 VNB 0.28fF
C885 VPB.n385 VNB 0.02fF
C886 VPB.n386 VNB 0.02fF
C887 VPB.n387 VNB 0.02fF
C888 VPB.n388 VNB 0.05fF
C889 VPB.n389 VNB 0.21fF
C890 VPB.n390 VNB 0.02fF
C891 VPB.n391 VNB 0.01fF
C892 VPB.n392 VNB 0.02fF
C893 VPB.n393 VNB 0.14fF
C894 VPB.n394 VNB 0.16fF
C895 VPB.n395 VNB 0.02fF
C896 VPB.n396 VNB 0.02fF
C897 VPB.n397 VNB 0.02fF
C898 VPB.n398 VNB 0.10fF
C899 VPB.n399 VNB 0.02fF
C900 VPB.n400 VNB 0.14fF
C901 VPB.n401 VNB 0.16fF
C902 VPB.n402 VNB 0.02fF
C903 VPB.n403 VNB 0.02fF
C904 VPB.n404 VNB 0.02fF
C905 VPB.n405 VNB 0.14fF
C906 VPB.n406 VNB 0.15fF
C907 VPB.n407 VNB 0.02fF
C908 VPB.n408 VNB 0.02fF
C909 VPB.n409 VNB 0.02fF
C910 VPB.n410 VNB 0.14fF
C911 VPB.n411 VNB 0.15fF
C912 VPB.n412 VNB 0.02fF
C913 VPB.n413 VNB 0.02fF
C914 VPB.n414 VNB 0.02fF
C915 VPB.n415 VNB 0.10fF
C916 VPB.n416 VNB 0.02fF
C917 VPB.n417 VNB 0.14fF
C918 VPB.n418 VNB 0.16fF
C919 VPB.n419 VNB 0.02fF
C920 VPB.n420 VNB 0.02fF
C921 VPB.n421 VNB 0.02fF
C922 VPB.n422 VNB 0.14fF
C923 VPB.n423 VNB 0.16fF
C924 VPB.n424 VNB 0.02fF
C925 VPB.n425 VNB 0.02fF
C926 VPB.n426 VNB 0.02fF
C927 VPB.n427 VNB 0.06fF
C928 VPB.n428 VNB 0.21fF
C929 VPB.n429 VNB 0.02fF
C930 VPB.n430 VNB 0.01fF
C931 VPB.n431 VNB 0.02fF
C932 VPB.n432 VNB 0.28fF
C933 VPB.n433 VNB 0.02fF
C934 VPB.n434 VNB 0.02fF
C935 VPB.n435 VNB 0.02fF
C936 VPB.n436 VNB 0.28fF
C937 VPB.n437 VNB 0.01fF
C938 VPB.n438 VNB 0.02fF
C939 VPB.n439 VNB 0.04fF
C940 VPB.n440 VNB 0.02fF
C941 VPB.n441 VNB 0.02fF
C942 VPB.n442 VNB 0.02fF
C943 VPB.n443 VNB 0.04fF
C944 VPB.n444 VNB 0.02fF
C945 VPB.n445 VNB 0.24fF
C946 VPB.n446 VNB 0.04fF
C947 VPB.n448 VNB 0.02fF
C948 VPB.n449 VNB 0.02fF
C949 VPB.n450 VNB 0.02fF
C950 VPB.n451 VNB 0.02fF
C951 VPB.n453 VNB 0.02fF
C952 VPB.n454 VNB 0.02fF
C953 VPB.n455 VNB 0.02fF
C954 VPB.n457 VNB 0.28fF
C955 VPB.n459 VNB 0.03fF
C956 VPB.n460 VNB 0.02fF
C957 VPB.n461 VNB 0.03fF
C958 VPB.n462 VNB 0.03fF
C959 VPB.n463 VNB 0.28fF
C960 VPB.n464 VNB 0.01fF
C961 VPB.n465 VNB 0.02fF
C962 VPB.n466 VNB 0.04fF
C963 VPB.n467 VNB 0.05fF
C964 VPB.n468 VNB 0.23fF
C965 VPB.n469 VNB 0.02fF
C966 VPB.n470 VNB 0.01fF
C967 VPB.n471 VNB 0.02fF
C968 VPB.n472 VNB 0.14fF
C969 VPB.n473 VNB 0.16fF
C970 VPB.n474 VNB 0.02fF
C971 VPB.n475 VNB 0.02fF
C972 VPB.n476 VNB 0.02fF
C973 VPB.n477 VNB 0.10fF
C974 VPB.n478 VNB 0.02fF
C975 VPB.n479 VNB 0.14fF
C976 VPB.n480 VNB 0.15fF
C977 VPB.n481 VNB 0.02fF
C978 VPB.n482 VNB 0.02fF
C979 VPB.n483 VNB 0.02fF
C980 VPB.n484 VNB 0.14fF
C981 VPB.n485 VNB 0.15fF
C982 VPB.n486 VNB 0.02fF
C983 VPB.n487 VNB 0.02fF
C984 VPB.n488 VNB 0.02fF
C985 VPB.n489 VNB 0.14fF
C986 VPB.n490 VNB 0.16fF
C987 VPB.n491 VNB 0.02fF
C988 VPB.n492 VNB 0.02fF
C989 VPB.n493 VNB 0.02fF
C990 VPB.n494 VNB 0.06fF
C991 VPB.n495 VNB 0.24fF
C992 VPB.n496 VNB 0.02fF
C993 VPB.n497 VNB 0.01fF
C994 VPB.n498 VNB 0.02fF
C995 VPB.n499 VNB 0.28fF
C996 VPB.n500 VNB 0.01fF
C997 VPB.n501 VNB 0.02fF
C998 VPB.n502 VNB 0.04fF
C999 VPB.n503 VNB 0.02fF
C1000 VPB.n504 VNB 0.02fF
C1001 VPB.n505 VNB 0.02fF
C1002 VPB.n506 VNB 0.04fF
C1003 VPB.n507 VNB 0.02fF
C1004 VPB.n508 VNB 0.20fF
C1005 VPB.n509 VNB 0.04fF
C1006 VPB.n511 VNB 0.02fF
C1007 VPB.n512 VNB 0.02fF
C1008 VPB.n513 VNB 0.02fF
C1009 VPB.n514 VNB 0.02fF
C1010 VPB.n516 VNB 0.02fF
C1011 VPB.n517 VNB 0.02fF
C1012 VPB.n518 VNB 0.02fF
C1013 VPB.n520 VNB 0.28fF
C1014 VPB.n522 VNB 0.03fF
C1015 VPB.n523 VNB 0.02fF
C1016 VPB.n524 VNB 0.03fF
C1017 VPB.n525 VNB 0.03fF
C1018 VPB.n526 VNB 0.28fF
C1019 VPB.n527 VNB 0.01fF
C1020 VPB.n528 VNB 0.02fF
C1021 VPB.n529 VNB 0.04fF
C1022 VPB.n530 VNB 0.05fF
C1023 VPB.n531 VNB 0.23fF
C1024 VPB.n532 VNB 0.02fF
C1025 VPB.n533 VNB 0.01fF
C1026 VPB.n534 VNB 0.02fF
C1027 VPB.n535 VNB 0.14fF
C1028 VPB.n536 VNB 0.16fF
C1029 VPB.n537 VNB 0.02fF
C1030 VPB.n538 VNB 0.02fF
C1031 VPB.n539 VNB 0.02fF
C1032 VPB.n540 VNB 0.10fF
C1033 VPB.n541 VNB 0.02fF
C1034 VPB.n542 VNB 0.14fF
C1035 VPB.n543 VNB 0.15fF
C1036 VPB.n544 VNB 0.02fF
C1037 VPB.n545 VNB 0.02fF
C1038 VPB.n546 VNB 0.02fF
C1039 VPB.n547 VNB 0.14fF
C1040 VPB.n548 VNB 0.15fF
C1041 VPB.n549 VNB 0.02fF
C1042 VPB.n550 VNB 0.02fF
C1043 VPB.n551 VNB 0.02fF
C1044 VPB.n552 VNB 0.14fF
C1045 VPB.n553 VNB 0.16fF
C1046 VPB.n554 VNB 0.02fF
C1047 VPB.n555 VNB 0.02fF
C1048 VPB.n556 VNB 0.02fF
C1049 VPB.n557 VNB 0.06fF
C1050 VPB.n558 VNB 0.24fF
C1051 VPB.n559 VNB 0.02fF
C1052 VPB.n560 VNB 0.01fF
C1053 VPB.n561 VNB 0.02fF
C1054 VPB.n562 VNB 0.28fF
C1055 VPB.n563 VNB 0.01fF
C1056 VPB.n564 VNB 0.02fF
C1057 VPB.n565 VNB 0.04fF
C1058 VPB.n566 VNB 0.02fF
C1059 VPB.n567 VNB 0.02fF
C1060 VPB.n568 VNB 0.02fF
C1061 VPB.n569 VNB 0.04fF
C1062 VPB.n570 VNB 0.02fF
C1063 VPB.n571 VNB 0.24fF
C1064 VPB.n572 VNB 0.04fF
C1065 VPB.n574 VNB 0.02fF
C1066 VPB.n575 VNB 0.02fF
C1067 VPB.n576 VNB 0.02fF
C1068 VPB.n577 VNB 0.02fF
C1069 VPB.n579 VNB 0.02fF
C1070 VPB.n580 VNB 0.02fF
C1071 VPB.n581 VNB 0.02fF
C1072 VPB.n583 VNB 0.28fF
C1073 VPB.n585 VNB 0.03fF
C1074 VPB.n586 VNB 0.02fF
C1075 VPB.n587 VNB 0.03fF
C1076 VPB.n588 VNB 0.03fF
C1077 VPB.n589 VNB 0.28fF
C1078 VPB.n590 VNB 0.01fF
C1079 VPB.n591 VNB 0.02fF
C1080 VPB.n592 VNB 0.04fF
C1081 VPB.n593 VNB 0.28fF
C1082 VPB.n594 VNB 0.02fF
C1083 VPB.n595 VNB 0.02fF
C1084 VPB.n596 VNB 0.02fF
C1085 VPB.n597 VNB 0.05fF
C1086 VPB.n598 VNB 0.21fF
C1087 VPB.n599 VNB 0.02fF
C1088 VPB.n600 VNB 0.01fF
C1089 VPB.n601 VNB 0.02fF
C1090 VPB.n602 VNB 0.14fF
C1091 VPB.n603 VNB 0.16fF
C1092 VPB.n604 VNB 0.02fF
C1093 VPB.n605 VNB 0.02fF
C1094 VPB.n606 VNB 0.02fF
C1095 VPB.n607 VNB 0.10fF
C1096 VPB.n608 VNB 0.02fF
C1097 VPB.n609 VNB 0.14fF
C1098 VPB.n610 VNB 0.16fF
C1099 VPB.n611 VNB 0.02fF
C1100 VPB.n612 VNB 0.02fF
C1101 VPB.n613 VNB 0.02fF
C1102 VPB.n614 VNB 0.14fF
C1103 VPB.n615 VNB 0.15fF
C1104 VPB.n616 VNB 0.02fF
C1105 VPB.n617 VNB 0.02fF
C1106 VPB.n618 VNB 0.02fF
C1107 VPB.n619 VNB 0.14fF
C1108 VPB.n620 VNB 0.15fF
C1109 VPB.n621 VNB 0.02fF
C1110 VPB.n622 VNB 0.02fF
C1111 VPB.n623 VNB 0.02fF
C1112 VPB.n624 VNB 0.10fF
C1113 VPB.n625 VNB 0.02fF
C1114 VPB.n626 VNB 0.14fF
C1115 VPB.n627 VNB 0.16fF
C1116 VPB.n628 VNB 0.02fF
C1117 VPB.n629 VNB 0.02fF
C1118 VPB.n630 VNB 0.02fF
C1119 VPB.n631 VNB 0.14fF
C1120 VPB.n632 VNB 0.16fF
C1121 VPB.n633 VNB 0.02fF
C1122 VPB.n634 VNB 0.02fF
C1123 VPB.n635 VNB 0.02fF
C1124 VPB.n636 VNB 0.06fF
C1125 VPB.n637 VNB 0.21fF
C1126 VPB.n638 VNB 0.02fF
C1127 VPB.n639 VNB 0.01fF
C1128 VPB.n640 VNB 0.02fF
C1129 VPB.n641 VNB 0.28fF
C1130 VPB.n642 VNB 0.02fF
C1131 VPB.n643 VNB 0.02fF
C1132 VPB.n644 VNB 0.02fF
C1133 VPB.n645 VNB 0.28fF
C1134 VPB.n646 VNB 0.01fF
C1135 VPB.n647 VNB 0.02fF
C1136 VPB.n648 VNB 0.04fF
C1137 VPB.n649 VNB 0.02fF
C1138 VPB.n650 VNB 0.02fF
C1139 VPB.n651 VNB 0.02fF
C1140 VPB.n652 VNB 0.04fF
C1141 VPB.n653 VNB 0.02fF
C1142 VPB.n654 VNB 0.29fF
C1143 VPB.n655 VNB 0.04fF
C1144 VPB.n657 VNB 0.02fF
C1145 VPB.n658 VNB 0.02fF
C1146 VPB.n659 VNB 0.02fF
C1147 VPB.n660 VNB 0.02fF
C1148 VPB.n662 VNB 0.02fF
C1149 VPB.n663 VNB 0.02fF
C1150 VPB.n664 VNB 0.02fF
C1151 VPB.n666 VNB 0.28fF
C1152 VPB.n668 VNB 0.03fF
C1153 VPB.n669 VNB 0.02fF
C1154 VPB.n670 VNB 0.03fF
C1155 VPB.n671 VNB 0.03fF
C1156 VPB.n672 VNB 0.28fF
C1157 VPB.n673 VNB 0.01fF
C1158 VPB.n674 VNB 0.02fF
C1159 VPB.n675 VNB 0.04fF
C1160 VPB.n676 VNB 0.28fF
C1161 VPB.n677 VNB 0.02fF
C1162 VPB.n678 VNB 0.02fF
C1163 VPB.n679 VNB 0.02fF
C1164 VPB.n680 VNB 0.05fF
C1165 VPB.n681 VNB 0.21fF
C1166 VPB.n682 VNB 0.02fF
C1167 VPB.n683 VNB 0.01fF
C1168 VPB.n684 VNB 0.02fF
C1169 VPB.n685 VNB 0.14fF
C1170 VPB.n686 VNB 0.16fF
C1171 VPB.n687 VNB 0.02fF
C1172 VPB.n688 VNB 0.02fF
C1173 VPB.n689 VNB 0.02fF
C1174 VPB.n690 VNB 0.10fF
C1175 VPB.n691 VNB 0.02fF
C1176 VPB.n692 VNB 0.14fF
C1177 VPB.n693 VNB 0.16fF
C1178 VPB.n694 VNB 0.02fF
C1179 VPB.n695 VNB 0.02fF
C1180 VPB.n696 VNB 0.02fF
C1181 VPB.n697 VNB 0.14fF
C1182 VPB.n698 VNB 0.15fF
C1183 VPB.n699 VNB 0.02fF
C1184 VPB.n700 VNB 0.02fF
C1185 VPB.n701 VNB 0.02fF
C1186 VPB.n702 VNB 0.14fF
C1187 VPB.n703 VNB 0.15fF
C1188 VPB.n704 VNB 0.02fF
C1189 VPB.n705 VNB 0.02fF
C1190 VPB.n706 VNB 0.02fF
C1191 VPB.n707 VNB 0.10fF
C1192 VPB.n708 VNB 0.02fF
C1193 VPB.n709 VNB 0.14fF
C1194 VPB.n710 VNB 0.16fF
C1195 VPB.n711 VNB 0.02fF
C1196 VPB.n712 VNB 0.02fF
C1197 VPB.n713 VNB 0.02fF
C1198 VPB.n714 VNB 0.14fF
C1199 VPB.n715 VNB 0.16fF
C1200 VPB.n716 VNB 0.02fF
C1201 VPB.n717 VNB 0.02fF
C1202 VPB.n718 VNB 0.02fF
C1203 VPB.n719 VNB 0.06fF
C1204 VPB.n720 VNB 0.21fF
C1205 VPB.n721 VNB 0.02fF
C1206 VPB.n722 VNB 0.01fF
C1207 VPB.n723 VNB 0.02fF
C1208 VPB.n724 VNB 0.28fF
C1209 VPB.n725 VNB 0.02fF
C1210 VPB.n726 VNB 0.02fF
C1211 VPB.n727 VNB 0.02fF
C1212 VPB.n728 VNB 0.28fF
C1213 VPB.n729 VNB 0.01fF
C1214 VPB.n730 VNB 0.02fF
C1215 VPB.n731 VNB 0.04fF
C1216 VPB.n732 VNB 0.02fF
C1217 VPB.n733 VNB 0.02fF
C1218 VPB.n734 VNB 0.02fF
C1219 VPB.n735 VNB 0.04fF
C1220 VPB.n736 VNB 0.02fF
C1221 VPB.n737 VNB 0.24fF
C1222 VPB.n738 VNB 0.04fF
C1223 VPB.n740 VNB 0.02fF
C1224 VPB.n741 VNB 0.02fF
C1225 VPB.n742 VNB 0.02fF
C1226 VPB.n743 VNB 0.02fF
C1227 VPB.n745 VNB 0.02fF
C1228 VPB.n746 VNB 0.02fF
C1229 VPB.n747 VNB 0.02fF
C1230 VPB.n749 VNB 0.28fF
C1231 VPB.n751 VNB 0.03fF
C1232 VPB.n752 VNB 0.02fF
C1233 VPB.n753 VNB 0.03fF
C1234 VPB.n754 VNB 0.03fF
C1235 VPB.n755 VNB 0.28fF
C1236 VPB.n756 VNB 0.01fF
C1237 VPB.n757 VNB 0.02fF
C1238 VPB.n758 VNB 0.04fF
C1239 VPB.n759 VNB 0.05fF
C1240 VPB.n760 VNB 0.23fF
C1241 VPB.n761 VNB 0.02fF
C1242 VPB.n762 VNB 0.01fF
C1243 VPB.n763 VNB 0.02fF
C1244 VPB.n764 VNB 0.14fF
C1245 VPB.n765 VNB 0.16fF
C1246 VPB.n766 VNB 0.02fF
C1247 VPB.n767 VNB 0.02fF
C1248 VPB.n768 VNB 0.02fF
C1249 VPB.n769 VNB 0.10fF
C1250 VPB.n770 VNB 0.02fF
C1251 VPB.n771 VNB 0.14fF
C1252 VPB.n772 VNB 0.15fF
C1253 VPB.n773 VNB 0.02fF
C1254 VPB.n774 VNB 0.02fF
C1255 VPB.n775 VNB 0.02fF
C1256 VPB.n776 VNB 0.14fF
C1257 VPB.n777 VNB 0.15fF
C1258 VPB.n778 VNB 0.02fF
C1259 VPB.n779 VNB 0.02fF
C1260 VPB.n780 VNB 0.02fF
C1261 VPB.n781 VNB 0.14fF
C1262 VPB.n782 VNB 0.16fF
C1263 VPB.n783 VNB 0.02fF
C1264 VPB.n784 VNB 0.02fF
C1265 VPB.n785 VNB 0.02fF
C1266 VPB.n786 VNB 0.06fF
C1267 VPB.n787 VNB 0.24fF
C1268 VPB.n788 VNB 0.02fF
C1269 VPB.n789 VNB 0.01fF
C1270 VPB.n790 VNB 0.02fF
C1271 VPB.n791 VNB 0.28fF
C1272 VPB.n792 VNB 0.01fF
C1273 VPB.n793 VNB 0.02fF
C1274 VPB.n794 VNB 0.04fF
C1275 VPB.n795 VNB 0.02fF
C1276 VPB.n796 VNB 0.02fF
C1277 VPB.n797 VNB 0.02fF
C1278 VPB.n798 VNB 0.04fF
C1279 VPB.n799 VNB 0.02fF
C1280 VPB.n800 VNB 0.24fF
C1281 VPB.n801 VNB 0.04fF
C1282 VPB.n803 VNB 0.02fF
C1283 VPB.n804 VNB 0.02fF
C1284 VPB.n805 VNB 0.02fF
C1285 VPB.n806 VNB 0.02fF
C1286 VPB.n808 VNB 0.02fF
C1287 VPB.n809 VNB 0.02fF
C1288 VPB.n810 VNB 0.02fF
C1289 VPB.n812 VNB 0.28fF
C1290 VPB.n814 VNB 0.03fF
C1291 VPB.n815 VNB 0.02fF
C1292 VPB.n816 VNB 0.03fF
C1293 VPB.n817 VNB 0.03fF
C1294 VPB.n818 VNB 0.28fF
C1295 VPB.n819 VNB 0.01fF
C1296 VPB.n820 VNB 0.02fF
C1297 VPB.n821 VNB 0.04fF
C1298 VPB.n822 VNB 0.28fF
C1299 VPB.n823 VNB 0.02fF
C1300 VPB.n824 VNB 0.02fF
C1301 VPB.n825 VNB 0.02fF
C1302 VPB.n826 VNB 0.05fF
C1303 VPB.n827 VNB 0.21fF
C1304 VPB.n828 VNB 0.02fF
C1305 VPB.n829 VNB 0.01fF
C1306 VPB.n830 VNB 0.02fF
C1307 VPB.n831 VNB 0.14fF
C1308 VPB.n832 VNB 0.16fF
C1309 VPB.n833 VNB 0.02fF
C1310 VPB.n834 VNB 0.02fF
C1311 VPB.n835 VNB 0.02fF
C1312 VPB.n836 VNB 0.02fF
C1313 VPB.n837 VNB 0.02fF
C1314 VPB.n838 VNB 0.02fF
C1315 VPB.n839 VNB 0.02fF
C1316 VPB.n840 VNB 0.02fF
C1317 VPB.n841 VNB 0.02fF
C1318 VPB.n842 VNB 0.02fF
C1319 VPB.n843 VNB 0.04fF
C1320 VPB.n844 VNB 0.04fF
C1321 VPB.n845 VNB 0.02fF
C1322 VPB.n846 VNB 0.02fF
C1323 VPB.n847 VNB 0.14fF
C1324 VPB.n848 VNB 0.16fF
C1325 VPB.n849 VNB 0.02fF
C1326 VPB.n850 VNB 0.02fF
C1327 VPB.n851 VNB 0.10fF
C1328 VPB.n852 VNB 0.02fF
C1329 VPB.n853 VNB 0.14fF
C1330 VPB.n854 VNB 0.15fF
C1331 VPB.n855 VNB 0.02fF
C1332 VPB.n856 VNB 0.02fF
C1333 VPB.n857 VNB 0.02fF
C1334 VPB.n858 VNB 0.14fF
C1335 VPB.n859 VNB 0.15fF
C1336 VPB.n860 VNB 0.02fF
C1337 VPB.n861 VNB 0.02fF
C1338 VPB.n862 VNB 0.02fF
C1339 VPB.n863 VNB 0.14fF
C1340 VPB.n864 VNB 0.16fF
C1341 VPB.n865 VNB 0.02fF
C1342 VPB.n866 VNB 0.02fF
C1343 VPB.n867 VNB 0.02fF
C1344 VPB.n868 VNB 0.06fF
C1345 VPB.n869 VNB 0.24fF
C1346 VPB.n870 VNB 0.02fF
C1347 VPB.n871 VNB 0.01fF
C1348 VPB.n872 VNB 0.02fF
C1349 VPB.n873 VNB 0.28fF
C1350 VPB.n874 VNB 0.01fF
C1351 VPB.n875 VNB 0.02fF
C1352 VPB.n876 VNB 0.04fF
C1353 VPB.n877 VNB 0.02fF
C1354 VPB.n878 VNB 0.02fF
C1355 VPB.n879 VNB 0.02fF
C1356 VPB.n880 VNB 0.04fF
C1357 VPB.n881 VNB 0.02fF
C1358 VPB.n882 VNB 0.20fF
C1359 VPB.n883 VNB 0.04fF
C1360 VPB.n885 VNB 0.02fF
C1361 VPB.n886 VNB 0.02fF
C1362 VPB.n887 VNB 0.02fF
C1363 VPB.n888 VNB 0.02fF
C1364 VPB.n890 VNB 0.02fF
C1365 VPB.n891 VNB 0.02fF
C1366 VPB.n892 VNB 0.02fF
C1367 VPB.n894 VNB 0.28fF
C1368 VPB.n896 VNB 0.03fF
C1369 VPB.n897 VNB 0.02fF
C1370 VPB.n898 VNB 0.03fF
C1371 VPB.n899 VNB 0.03fF
C1372 VPB.n900 VNB 0.28fF
C1373 VPB.n901 VNB 0.01fF
C1374 VPB.n902 VNB 0.02fF
C1375 VPB.n903 VNB 0.04fF
C1376 VPB.n904 VNB 0.05fF
C1377 VPB.n905 VNB 0.23fF
C1378 VPB.n906 VNB 0.02fF
C1379 VPB.n907 VNB 0.01fF
C1380 VPB.n908 VNB 0.02fF
C1381 VPB.n909 VNB 0.14fF
C1382 VPB.n910 VNB 0.16fF
C1383 VPB.n911 VNB 0.02fF
C1384 VPB.n912 VNB 0.02fF
C1385 VPB.n913 VNB 0.02fF
C1386 VPB.n914 VNB 0.10fF
C1387 VPB.n915 VNB 0.02fF
C1388 VPB.n916 VNB 0.14fF
C1389 VPB.n917 VNB 0.15fF
C1390 VPB.n918 VNB 0.02fF
C1391 VPB.n919 VNB 0.02fF
C1392 VPB.n920 VNB 0.02fF
C1393 VPB.n921 VNB 0.14fF
C1394 VPB.n922 VNB 0.15fF
C1395 VPB.n923 VNB 0.02fF
C1396 VPB.n924 VNB 0.02fF
C1397 VPB.n925 VNB 0.02fF
C1398 VPB.n926 VNB 0.14fF
C1399 VPB.n927 VNB 0.16fF
C1400 VPB.n928 VNB 0.02fF
C1401 VPB.n929 VNB 0.02fF
C1402 VPB.n930 VNB 0.02fF
C1403 VPB.n931 VNB 0.06fF
C1404 VPB.n932 VNB 0.24fF
C1405 VPB.n933 VNB 0.02fF
C1406 VPB.n934 VNB 0.01fF
C1407 VPB.n935 VNB 0.02fF
C1408 VPB.n936 VNB 0.28fF
C1409 VPB.n937 VNB 0.01fF
C1410 VPB.n938 VNB 0.02fF
C1411 VPB.n939 VNB 0.04fF
C1412 VPB.n940 VNB 0.02fF
C1413 VPB.n941 VNB 0.02fF
C1414 VPB.n942 VNB 0.02fF
C1415 VPB.n943 VNB 0.04fF
C1416 VPB.n944 VNB 0.02fF
C1417 VPB.n945 VNB 0.24fF
C1418 VPB.n946 VNB 0.04fF
C1419 VPB.n948 VNB 0.02fF
C1420 VPB.n949 VNB 0.02fF
C1421 VPB.n950 VNB 0.02fF
C1422 VPB.n951 VNB 0.02fF
C1423 VPB.n953 VNB 0.02fF
C1424 VPB.n954 VNB 0.02fF
C1425 VPB.n955 VNB 0.02fF
C1426 VPB.n957 VNB 0.28fF
C1427 VPB.n959 VNB 0.03fF
C1428 VPB.n960 VNB 0.02fF
C1429 VPB.n961 VNB 0.03fF
C1430 VPB.n962 VNB 0.03fF
C1431 VPB.n963 VNB 0.28fF
C1432 VPB.n964 VNB 0.01fF
C1433 VPB.n965 VNB 0.02fF
C1434 VPB.n966 VNB 0.04fF
C1435 VPB.n967 VNB 0.28fF
C1436 VPB.n968 VNB 0.02fF
C1437 VPB.n969 VNB 0.02fF
C1438 VPB.n970 VNB 0.02fF
C1439 VPB.n971 VNB 0.05fF
C1440 VPB.n972 VNB 0.21fF
C1441 VPB.n973 VNB 0.02fF
C1442 VPB.n974 VNB 0.01fF
C1443 VPB.n975 VNB 0.02fF
C1444 VPB.n976 VNB 0.14fF
C1445 VPB.n977 VNB 0.16fF
C1446 VPB.n978 VNB 0.02fF
C1447 VPB.n979 VNB 0.02fF
C1448 VPB.n980 VNB 0.02fF
C1449 VPB.n981 VNB 0.10fF
C1450 VPB.n982 VNB 0.02fF
C1451 VPB.n983 VNB 0.14fF
C1452 VPB.n984 VNB 0.16fF
C1453 VPB.n985 VNB 0.02fF
C1454 VPB.n986 VNB 0.02fF
C1455 VPB.n987 VNB 0.02fF
C1456 VPB.n988 VNB 0.14fF
C1457 VPB.n989 VNB 0.15fF
C1458 VPB.n990 VNB 0.02fF
C1459 VPB.n991 VNB 0.02fF
C1460 VPB.n992 VNB 0.02fF
C1461 VPB.n993 VNB 0.14fF
C1462 VPB.n994 VNB 0.15fF
C1463 VPB.n995 VNB 0.02fF
C1464 VPB.n996 VNB 0.02fF
C1465 VPB.n997 VNB 0.02fF
C1466 VPB.n998 VNB 0.10fF
C1467 VPB.n999 VNB 0.02fF
C1468 VPB.n1000 VNB 0.14fF
C1469 VPB.n1001 VNB 0.16fF
C1470 VPB.n1002 VNB 0.02fF
C1471 VPB.n1003 VNB 0.02fF
C1472 VPB.n1004 VNB 0.02fF
C1473 VPB.n1005 VNB 0.14fF
C1474 VPB.n1006 VNB 0.16fF
C1475 VPB.n1007 VNB 0.02fF
C1476 VPB.n1008 VNB 0.02fF
C1477 VPB.n1009 VNB 0.02fF
C1478 VPB.n1010 VNB 0.06fF
C1479 VPB.n1011 VNB 0.21fF
C1480 VPB.n1012 VNB 0.02fF
C1481 VPB.n1013 VNB 0.01fF
C1482 VPB.n1014 VNB 0.02fF
C1483 VPB.n1015 VNB 0.28fF
C1484 VPB.n1016 VNB 0.02fF
C1485 VPB.n1017 VNB 0.02fF
C1486 VPB.n1018 VNB 0.02fF
C1487 VPB.n1019 VNB 0.28fF
C1488 VPB.n1020 VNB 0.01fF
C1489 VPB.n1021 VNB 0.02fF
C1490 VPB.n1022 VNB 0.04fF
C1491 VPB.n1023 VNB 0.02fF
C1492 VPB.n1024 VNB 0.02fF
C1493 VPB.n1025 VNB 0.02fF
C1494 VPB.n1026 VNB 0.04fF
C1495 VPB.n1027 VNB 0.02fF
C1496 VPB.n1028 VNB 0.29fF
C1497 VPB.n1029 VNB 0.04fF
C1498 VPB.n1031 VNB 0.02fF
C1499 VPB.n1032 VNB 0.02fF
C1500 VPB.n1033 VNB 0.02fF
C1501 VPB.n1034 VNB 0.02fF
C1502 VPB.n1036 VNB 0.02fF
C1503 VPB.n1037 VNB 0.02fF
C1504 VPB.n1038 VNB 0.02fF
C1505 VPB.n1040 VNB 0.28fF
C1506 VPB.n1042 VNB 0.03fF
C1507 VPB.n1043 VNB 0.02fF
C1508 VPB.n1044 VNB 0.03fF
C1509 VPB.n1045 VNB 0.03fF
C1510 VPB.n1046 VNB 0.28fF
C1511 VPB.n1047 VNB 0.01fF
C1512 VPB.n1048 VNB 0.02fF
C1513 VPB.n1049 VNB 0.04fF
C1514 VPB.n1050 VNB 0.28fF
C1515 VPB.n1051 VNB 0.02fF
C1516 VPB.n1052 VNB 0.02fF
C1517 VPB.n1053 VNB 0.02fF
C1518 VPB.n1054 VNB 0.05fF
C1519 VPB.n1055 VNB 0.21fF
C1520 VPB.n1056 VNB 0.02fF
C1521 VPB.n1057 VNB 0.01fF
C1522 VPB.n1058 VNB 0.02fF
C1523 VPB.n1059 VNB 0.14fF
C1524 VPB.n1060 VNB 0.16fF
C1525 VPB.n1061 VNB 0.02fF
C1526 VPB.n1062 VNB 0.02fF
C1527 VPB.n1063 VNB 0.02fF
C1528 VPB.n1064 VNB 0.10fF
C1529 VPB.n1065 VNB 0.02fF
C1530 VPB.n1066 VNB 0.14fF
C1531 VPB.n1067 VNB 0.16fF
C1532 VPB.n1068 VNB 0.02fF
C1533 VPB.n1069 VNB 0.02fF
C1534 VPB.n1070 VNB 0.02fF
C1535 VPB.n1071 VNB 0.14fF
C1536 VPB.n1072 VNB 0.15fF
C1537 VPB.n1073 VNB 0.02fF
C1538 VPB.n1074 VNB 0.02fF
C1539 VPB.n1075 VNB 0.02fF
C1540 VPB.n1076 VNB 0.14fF
C1541 VPB.n1077 VNB 0.15fF
C1542 VPB.n1078 VNB 0.02fF
C1543 VPB.n1079 VNB 0.02fF
C1544 VPB.n1080 VNB 0.02fF
C1545 VPB.n1081 VNB 0.10fF
C1546 VPB.n1082 VNB 0.02fF
C1547 VPB.n1083 VNB 0.14fF
C1548 VPB.n1084 VNB 0.16fF
C1549 VPB.n1085 VNB 0.02fF
C1550 VPB.n1086 VNB 0.02fF
C1551 VPB.n1087 VNB 0.02fF
C1552 VPB.n1088 VNB 0.14fF
C1553 VPB.n1089 VNB 0.16fF
C1554 VPB.n1090 VNB 0.02fF
C1555 VPB.n1091 VNB 0.02fF
C1556 VPB.n1092 VNB 0.02fF
C1557 VPB.n1093 VNB 0.06fF
C1558 VPB.n1094 VNB 0.21fF
C1559 VPB.n1095 VNB 0.02fF
C1560 VPB.n1096 VNB 0.01fF
C1561 VPB.n1097 VNB 0.02fF
C1562 VPB.n1098 VNB 0.28fF
C1563 VPB.n1099 VNB 0.02fF
C1564 VPB.n1100 VNB 0.02fF
C1565 VPB.n1101 VNB 0.02fF
C1566 VPB.n1102 VNB 0.28fF
C1567 VPB.n1103 VNB 0.01fF
C1568 VPB.n1104 VNB 0.02fF
C1569 VPB.n1105 VNB 0.04fF
C1570 VPB.n1106 VNB 0.02fF
C1571 VPB.n1107 VNB 0.02fF
C1572 VPB.n1108 VNB 0.02fF
C1573 VPB.n1109 VNB 0.04fF
C1574 VPB.n1110 VNB 0.02fF
C1575 VPB.n1111 VNB 0.24fF
C1576 VPB.n1112 VNB 0.04fF
C1577 VPB.n1114 VNB 0.02fF
C1578 VPB.n1115 VNB 0.02fF
C1579 VPB.n1116 VNB 0.02fF
C1580 VPB.n1117 VNB 0.02fF
C1581 VPB.n1119 VNB 0.02fF
C1582 VPB.n1120 VNB 0.02fF
C1583 VPB.n1121 VNB 0.02fF
C1584 VPB.n1123 VNB 0.28fF
C1585 VPB.n1125 VNB 0.03fF
C1586 VPB.n1126 VNB 0.02fF
C1587 VPB.n1127 VNB 0.03fF
C1588 VPB.n1128 VNB 0.03fF
C1589 VPB.n1129 VNB 0.28fF
C1590 VPB.n1130 VNB 0.01fF
C1591 VPB.n1131 VNB 0.02fF
C1592 VPB.n1132 VNB 0.04fF
C1593 VPB.n1133 VNB 0.05fF
C1594 VPB.n1134 VNB 0.23fF
C1595 VPB.n1135 VNB 0.02fF
C1596 VPB.n1136 VNB 0.01fF
C1597 VPB.n1137 VNB 0.02fF
C1598 VPB.n1138 VNB 0.14fF
C1599 VPB.n1139 VNB 0.16fF
C1600 VPB.n1140 VNB 0.02fF
C1601 VPB.n1141 VNB 0.02fF
C1602 VPB.n1142 VNB 0.02fF
C1603 VPB.n1143 VNB 0.10fF
C1604 VPB.n1144 VNB 0.02fF
C1605 VPB.n1145 VNB 0.14fF
C1606 VPB.n1146 VNB 0.15fF
C1607 VPB.n1147 VNB 0.02fF
C1608 VPB.n1148 VNB 0.02fF
C1609 VPB.n1149 VNB 0.02fF
C1610 VPB.n1150 VNB 0.14fF
C1611 VPB.n1151 VNB 0.15fF
C1612 VPB.n1152 VNB 0.02fF
C1613 VPB.n1153 VNB 0.02fF
C1614 VPB.n1154 VNB 0.02fF
C1615 VPB.n1155 VNB 0.14fF
C1616 VPB.n1156 VNB 0.16fF
C1617 VPB.n1157 VNB 0.02fF
C1618 VPB.n1158 VNB 0.02fF
C1619 VPB.n1159 VNB 0.02fF
C1620 VPB.n1160 VNB 0.06fF
C1621 VPB.n1161 VNB 0.24fF
C1622 VPB.n1162 VNB 0.02fF
C1623 VPB.n1163 VNB 0.01fF
C1624 VPB.n1164 VNB 0.02fF
C1625 VPB.n1165 VNB 0.28fF
C1626 VPB.n1166 VNB 0.01fF
C1627 VPB.n1167 VNB 0.02fF
C1628 VPB.n1168 VNB 0.04fF
C1629 VPB.n1169 VNB 0.02fF
C1630 VPB.n1170 VNB 0.02fF
C1631 VPB.n1171 VNB 0.02fF
C1632 VPB.n1172 VNB 0.04fF
C1633 VPB.n1173 VNB 0.02fF
C1634 VPB.n1174 VNB 0.24fF
C1635 VPB.n1175 VNB 0.04fF
C1636 VPB.n1177 VNB 0.02fF
C1637 VPB.n1178 VNB 0.02fF
C1638 VPB.n1179 VNB 0.02fF
C1639 VPB.n1180 VNB 0.02fF
C1640 VPB.n1182 VNB 0.02fF
C1641 VPB.n1183 VNB 0.02fF
C1642 VPB.n1184 VNB 0.02fF
C1643 VPB.n1186 VNB 0.28fF
C1644 VPB.n1188 VNB 0.03fF
C1645 VPB.n1189 VNB 0.02fF
C1646 VPB.n1190 VNB 0.03fF
C1647 VPB.n1191 VNB 0.03fF
C1648 VPB.n1192 VNB 0.28fF
C1649 VPB.n1193 VNB 0.01fF
C1650 VPB.n1194 VNB 0.02fF
C1651 VPB.n1195 VNB 0.04fF
C1652 VPB.n1196 VNB 0.28fF
C1653 VPB.n1197 VNB 0.02fF
C1654 VPB.n1198 VNB 0.02fF
C1655 VPB.n1199 VNB 0.02fF
C1656 VPB.n1200 VNB 0.05fF
C1657 VPB.n1201 VNB 0.21fF
C1658 VPB.n1202 VNB 0.02fF
C1659 VPB.n1203 VNB 0.01fF
C1660 VPB.n1204 VNB 0.02fF
C1661 VPB.n1205 VNB 0.14fF
C1662 VPB.n1206 VNB 0.16fF
C1663 VPB.n1207 VNB 0.02fF
C1664 VPB.n1208 VNB 0.02fF
C1665 VPB.n1209 VNB 0.02fF
C1666 VPB.n1210 VNB 0.10fF
C1667 VPB.n1211 VNB 0.02fF
C1668 VPB.n1212 VNB 0.14fF
C1669 VPB.n1213 VNB 0.16fF
C1670 VPB.n1214 VNB 0.02fF
C1671 VPB.n1215 VNB 0.02fF
C1672 VPB.n1216 VNB 0.02fF
C1673 VPB.n1217 VNB 0.14fF
C1674 VPB.n1218 VNB 0.15fF
C1675 VPB.n1219 VNB 0.02fF
C1676 VPB.n1220 VNB 0.02fF
C1677 VPB.n1221 VNB 0.02fF
C1678 VPB.n1222 VNB 0.14fF
C1679 VPB.n1223 VNB 0.15fF
C1680 VPB.n1224 VNB 0.02fF
C1681 VPB.n1225 VNB 0.02fF
C1682 VPB.n1226 VNB 0.02fF
C1683 VPB.n1227 VNB 0.10fF
C1684 VPB.n1228 VNB 0.02fF
C1685 VPB.n1229 VNB 0.14fF
C1686 VPB.n1230 VNB 0.16fF
C1687 VPB.n1231 VNB 0.02fF
C1688 VPB.n1232 VNB 0.02fF
C1689 VPB.n1233 VNB 0.02fF
C1690 VPB.n1234 VNB 0.14fF
C1691 VPB.n1235 VNB 0.16fF
C1692 VPB.n1236 VNB 0.02fF
C1693 VPB.n1237 VNB 0.02fF
C1694 VPB.n1238 VNB 0.02fF
C1695 VPB.n1239 VNB 0.06fF
C1696 VPB.n1240 VNB 0.21fF
C1697 VPB.n1241 VNB 0.02fF
C1698 VPB.n1242 VNB 0.01fF
C1699 VPB.n1243 VNB 0.02fF
C1700 VPB.n1244 VNB 0.28fF
C1701 VPB.n1245 VNB 0.02fF
C1702 VPB.n1246 VNB 0.02fF
C1703 VPB.n1247 VNB 0.02fF
C1704 VPB.n1248 VNB 0.28fF
C1705 VPB.n1249 VNB 0.01fF
C1706 VPB.n1250 VNB 0.02fF
C1707 VPB.n1251 VNB 0.04fF
C1708 VPB.n1252 VNB 0.02fF
C1709 VPB.n1253 VNB 0.02fF
C1710 VPB.n1254 VNB 0.02fF
C1711 VPB.n1255 VNB 0.04fF
C1712 VPB.n1256 VNB 0.02fF
C1713 VPB.n1257 VNB 0.24fF
C1714 VPB.n1258 VNB 0.04fF
C1715 VPB.n1260 VNB 0.02fF
C1716 VPB.n1261 VNB 0.02fF
C1717 VPB.n1262 VNB 0.02fF
C1718 VPB.n1263 VNB 0.02fF
C1719 VPB.n1265 VNB 0.02fF
C1720 VPB.n1266 VNB 0.02fF
C1721 VPB.n1267 VNB 0.02fF
C1722 VPB.n1269 VNB 0.28fF
C1723 VPB.n1271 VNB 0.03fF
C1724 VPB.n1272 VNB 0.02fF
C1725 VPB.n1273 VNB 0.03fF
C1726 VPB.n1274 VNB 0.03fF
C1727 VPB.n1275 VNB 0.28fF
C1728 VPB.n1276 VNB 0.01fF
C1729 VPB.n1277 VNB 0.02fF
C1730 VPB.n1278 VNB 0.04fF
C1731 VPB.n1279 VNB 0.05fF
C1732 VPB.n1280 VNB 0.23fF
C1733 VPB.n1281 VNB 0.02fF
C1734 VPB.n1282 VNB 0.01fF
C1735 VPB.n1283 VNB 0.02fF
C1736 VPB.n1284 VNB 0.14fF
C1737 VPB.n1285 VNB 0.16fF
C1738 VPB.n1286 VNB 0.02fF
C1739 VPB.n1287 VNB 0.02fF
C1740 VPB.n1288 VNB 0.02fF
C1741 VPB.n1289 VNB 0.10fF
C1742 VPB.n1290 VNB 0.02fF
C1743 VPB.n1291 VNB 0.14fF
C1744 VPB.n1292 VNB 0.15fF
C1745 VPB.n1293 VNB 0.02fF
C1746 VPB.n1294 VNB 0.02fF
C1747 VPB.n1295 VNB 0.02fF
C1748 VPB.n1296 VNB 0.14fF
C1749 VPB.n1297 VNB 0.15fF
C1750 VPB.n1298 VNB 0.02fF
C1751 VPB.n1299 VNB 0.02fF
C1752 VPB.n1300 VNB 0.02fF
C1753 VPB.n1301 VNB 0.14fF
C1754 VPB.n1302 VNB 0.16fF
C1755 VPB.n1303 VNB 0.02fF
C1756 VPB.n1304 VNB 0.02fF
C1757 VPB.n1305 VNB 0.02fF
C1758 VPB.n1306 VNB 0.06fF
C1759 VPB.n1307 VNB 0.24fF
C1760 VPB.n1308 VNB 0.02fF
C1761 VPB.n1309 VNB 0.01fF
C1762 VPB.n1310 VNB 0.02fF
C1763 VPB.n1311 VNB 0.28fF
C1764 VPB.n1312 VNB 0.01fF
C1765 VPB.n1313 VNB 0.02fF
C1766 VPB.n1314 VNB 0.04fF
C1767 VPB.n1315 VNB 0.02fF
C1768 VPB.n1316 VNB 0.02fF
C1769 VPB.n1317 VNB 0.02fF
C1770 VPB.n1318 VNB 0.04fF
C1771 VPB.n1319 VNB 0.02fF
C1772 VPB.n1320 VNB 0.20fF
C1773 VPB.n1321 VNB 0.04fF
C1774 VPB.n1323 VNB 0.02fF
C1775 VPB.n1324 VNB 0.02fF
C1776 VPB.n1325 VNB 0.02fF
C1777 VPB.n1326 VNB 0.02fF
C1778 VPB.n1328 VNB 0.02fF
C1779 VPB.n1329 VNB 0.02fF
C1780 VPB.n1330 VNB 0.02fF
C1781 VPB.n1332 VNB 0.28fF
C1782 VPB.n1334 VNB 0.03fF
C1783 VPB.n1335 VNB 0.02fF
C1784 VPB.n1336 VNB 0.03fF
C1785 VPB.n1337 VNB 0.03fF
C1786 VPB.n1338 VNB 0.28fF
C1787 VPB.n1339 VNB 0.01fF
C1788 VPB.n1340 VNB 0.02fF
C1789 VPB.n1341 VNB 0.04fF
C1790 VPB.n1342 VNB 0.05fF
C1791 VPB.n1343 VNB 0.23fF
C1792 VPB.n1344 VNB 0.02fF
C1793 VPB.n1345 VNB 0.01fF
C1794 VPB.n1346 VNB 0.02fF
C1795 VPB.n1347 VNB 0.14fF
C1796 VPB.n1348 VNB 0.16fF
C1797 VPB.n1349 VNB 0.02fF
C1798 VPB.n1350 VNB 0.02fF
C1799 VPB.n1351 VNB 0.02fF
C1800 VPB.n1352 VNB 0.10fF
C1801 VPB.n1353 VNB 0.02fF
C1802 VPB.n1354 VNB 0.14fF
C1803 VPB.n1355 VNB 0.15fF
C1804 VPB.n1356 VNB 0.02fF
C1805 VPB.n1357 VNB 0.02fF
C1806 VPB.n1358 VNB 0.02fF
C1807 VPB.n1359 VNB 0.14fF
C1808 VPB.n1360 VNB 0.15fF
C1809 VPB.n1361 VNB 0.02fF
C1810 VPB.n1362 VNB 0.02fF
C1811 VPB.n1363 VNB 0.02fF
C1812 VPB.n1364 VNB 0.14fF
C1813 VPB.n1365 VNB 0.16fF
C1814 VPB.n1366 VNB 0.02fF
C1815 VPB.n1367 VNB 0.02fF
C1816 VPB.n1368 VNB 0.02fF
C1817 VPB.n1369 VNB 0.06fF
C1818 VPB.n1370 VNB 0.24fF
C1819 VPB.n1371 VNB 0.02fF
C1820 VPB.n1372 VNB 0.01fF
C1821 VPB.n1373 VNB 0.02fF
C1822 VPB.n1374 VNB 0.28fF
C1823 VPB.n1375 VNB 0.01fF
C1824 VPB.n1376 VNB 0.02fF
C1825 VPB.n1377 VNB 0.04fF
C1826 VPB.n1378 VNB 0.02fF
C1827 VPB.n1379 VNB 0.02fF
C1828 VPB.n1380 VNB 0.02fF
C1829 VPB.n1381 VNB 0.04fF
C1830 VPB.n1382 VNB 0.02fF
C1831 VPB.n1383 VNB 0.24fF
C1832 VPB.n1384 VNB 0.04fF
C1833 VPB.n1386 VNB 0.02fF
C1834 VPB.n1387 VNB 0.02fF
C1835 VPB.n1388 VNB 0.02fF
C1836 VPB.n1389 VNB 0.02fF
C1837 VPB.n1391 VNB 0.02fF
C1838 VPB.n1392 VNB 0.02fF
C1839 VPB.n1393 VNB 0.02fF
C1840 VPB.n1395 VNB 0.28fF
C1841 VPB.n1397 VNB 0.03fF
C1842 VPB.n1398 VNB 0.02fF
C1843 VPB.n1399 VNB 0.03fF
C1844 VPB.n1400 VNB 0.03fF
C1845 VPB.n1401 VNB 0.28fF
C1846 VPB.n1402 VNB 0.01fF
C1847 VPB.n1403 VNB 0.02fF
C1848 VPB.n1404 VNB 0.04fF
C1849 VPB.n1405 VNB 0.28fF
C1850 VPB.n1406 VNB 0.02fF
C1851 VPB.n1407 VNB 0.02fF
C1852 VPB.n1408 VNB 0.02fF
C1853 VPB.n1409 VNB 0.05fF
C1854 VPB.n1410 VNB 0.21fF
C1855 VPB.n1411 VNB 0.02fF
C1856 VPB.n1412 VNB 0.01fF
C1857 VPB.n1413 VNB 0.02fF
C1858 VPB.n1414 VNB 0.14fF
C1859 VPB.n1415 VNB 0.16fF
C1860 VPB.n1416 VNB 0.02fF
C1861 VPB.n1417 VNB 0.02fF
C1862 VPB.n1418 VNB 0.02fF
C1863 VPB.n1419 VNB 0.10fF
C1864 VPB.n1420 VNB 0.02fF
C1865 VPB.n1421 VNB 0.14fF
C1866 VPB.n1422 VNB 0.16fF
C1867 VPB.n1423 VNB 0.02fF
C1868 VPB.n1424 VNB 0.02fF
C1869 VPB.n1425 VNB 0.02fF
C1870 VPB.n1426 VNB 0.14fF
C1871 VPB.n1427 VNB 0.15fF
C1872 VPB.n1428 VNB 0.02fF
C1873 VPB.n1429 VNB 0.02fF
C1874 VPB.n1430 VNB 0.02fF
C1875 VPB.n1431 VNB 0.14fF
C1876 VPB.n1432 VNB 0.15fF
C1877 VPB.n1433 VNB 0.02fF
C1878 VPB.n1434 VNB 0.02fF
C1879 VPB.n1435 VNB 0.02fF
C1880 VPB.n1436 VNB 0.10fF
C1881 VPB.n1437 VNB 0.02fF
C1882 VPB.n1438 VNB 0.14fF
C1883 VPB.n1439 VNB 0.16fF
C1884 VPB.n1440 VNB 0.02fF
C1885 VPB.n1441 VNB 0.02fF
C1886 VPB.n1442 VNB 0.02fF
C1887 VPB.n1443 VNB 0.14fF
C1888 VPB.n1444 VNB 0.16fF
C1889 VPB.n1445 VNB 0.02fF
C1890 VPB.n1446 VNB 0.02fF
C1891 VPB.n1447 VNB 0.02fF
C1892 VPB.n1448 VNB 0.06fF
C1893 VPB.n1449 VNB 0.21fF
C1894 VPB.n1450 VNB 0.02fF
C1895 VPB.n1451 VNB 0.01fF
C1896 VPB.n1452 VNB 0.02fF
C1897 VPB.n1453 VNB 0.28fF
C1898 VPB.n1454 VNB 0.02fF
C1899 VPB.n1455 VNB 0.02fF
C1900 VPB.n1456 VNB 0.02fF
C1901 VPB.n1457 VNB 0.28fF
C1902 VPB.n1458 VNB 0.01fF
C1903 VPB.n1459 VNB 0.02fF
C1904 VPB.n1460 VNB 0.04fF
C1905 VPB.n1461 VNB 0.02fF
C1906 VPB.n1462 VNB 0.02fF
C1907 VPB.n1463 VNB 0.02fF
C1908 VPB.n1464 VNB 0.04fF
C1909 VPB.n1465 VNB 0.02fF
C1910 VPB.n1466 VNB 0.29fF
C1911 VPB.n1467 VNB 0.04fF
C1912 VPB.n1469 VNB 0.02fF
C1913 VPB.n1470 VNB 0.02fF
C1914 VPB.n1471 VNB 0.02fF
C1915 VPB.n1472 VNB 0.02fF
C1916 VPB.n1474 VNB 0.02fF
C1917 VPB.n1475 VNB 0.02fF
C1918 VPB.n1476 VNB 0.02fF
C1919 VPB.n1478 VNB 0.28fF
C1920 VPB.n1480 VNB 0.03fF
C1921 VPB.n1481 VNB 0.02fF
C1922 VPB.n1482 VNB 0.03fF
C1923 VPB.n1483 VNB 0.03fF
C1924 VPB.n1484 VNB 0.28fF
C1925 VPB.n1485 VNB 0.01fF
C1926 VPB.n1486 VNB 0.02fF
C1927 VPB.n1487 VNB 0.04fF
C1928 VPB.n1488 VNB 0.28fF
C1929 VPB.n1489 VNB 0.02fF
C1930 VPB.n1490 VNB 0.02fF
C1931 VPB.n1491 VNB 0.02fF
C1932 VPB.n1492 VNB 0.05fF
C1933 VPB.n1493 VNB 0.21fF
C1934 VPB.n1494 VNB 0.02fF
C1935 VPB.n1495 VNB 0.01fF
C1936 VPB.n1496 VNB 0.02fF
C1937 VPB.n1497 VNB 0.14fF
C1938 VPB.n1498 VNB 0.16fF
C1939 VPB.n1499 VNB 0.02fF
C1940 VPB.n1500 VNB 0.02fF
C1941 VPB.n1501 VNB 0.02fF
C1942 VPB.n1502 VNB 0.10fF
C1943 VPB.n1503 VNB 0.02fF
C1944 VPB.n1504 VNB 0.14fF
C1945 VPB.n1505 VNB 0.16fF
C1946 VPB.n1506 VNB 0.02fF
C1947 VPB.n1507 VNB 0.02fF
C1948 VPB.n1508 VNB 0.02fF
C1949 VPB.n1509 VNB 0.14fF
C1950 VPB.n1510 VNB 0.15fF
C1951 VPB.n1511 VNB 0.02fF
C1952 VPB.n1512 VNB 0.02fF
C1953 VPB.n1513 VNB 0.02fF
C1954 VPB.n1514 VNB 0.14fF
C1955 VPB.n1515 VNB 0.15fF
C1956 VPB.n1516 VNB 0.02fF
C1957 VPB.n1517 VNB 0.02fF
C1958 VPB.n1518 VNB 0.02fF
C1959 VPB.n1519 VNB 0.10fF
C1960 VPB.n1520 VNB 0.02fF
C1961 VPB.n1521 VNB 0.14fF
C1962 VPB.n1522 VNB 0.16fF
C1963 VPB.n1523 VNB 0.02fF
C1964 VPB.n1524 VNB 0.02fF
C1965 VPB.n1525 VNB 0.02fF
C1966 VPB.n1526 VNB 0.14fF
C1967 VPB.n1527 VNB 0.16fF
C1968 VPB.n1528 VNB 0.02fF
C1969 VPB.n1529 VNB 0.02fF
C1970 VPB.n1530 VNB 0.02fF
C1971 VPB.n1531 VNB 0.02fF
C1972 VPB.n1532 VNB 0.02fF
C1973 VPB.n1533 VNB 0.04fF
C1974 VPB.n1534 VNB 0.04fF
C1975 VPB.n1535 VNB 0.02fF
C1976 VPB.n1536 VNB 0.02fF
C1977 VPB.n1537 VNB 0.02fF
C1978 VPB.n1538 VNB 0.02fF
C1979 VPB.n1539 VNB 0.02fF
C1980 VPB.n1540 VNB 0.02fF
C1981 VPB.n1541 VNB 0.03fF
C1982 VPB.n1542 VNB 0.04fF
C1983 VPB.n1543 VNB 0.02fF
C1984 VPB.n1544 VNB 0.02fF
C1985 VPB.n1545 VNB 0.02fF
C1986 VPB.n1546 VNB 0.04fF
C1987 VPB.n1547 VNB 0.04fF
C1988 VPB.n1549 VNB 0.43fF
C1989 a_5227_383.n0 VNB 0.07fF
C1990 a_5227_383.n1 VNB 0.90fF
C1991 a_5227_383.n2 VNB 0.90fF
C1992 a_5227_383.n3 VNB 1.05fF
C1993 a_5227_383.n4 VNB 0.33fF
C1994 a_5227_383.n5 VNB 0.43fF
C1995 a_5227_383.n6 VNB 0.54fF
C1996 a_5227_383.n7 VNB 0.78fF
C1997 a_5227_383.n8 VNB 0.48fF
C1998 a_5227_383.t12 VNB 0.95fF
C1999 a_5227_383.n9 VNB 0.67fF
C2000 a_5227_383.n10 VNB 4.19fF
C2001 a_5227_383.n11 VNB 0.74fF
C2002 a_5227_383.n12 VNB 0.06fF
C2003 a_5227_383.n13 VNB 0.58fF
C2004 a_5227_383.n14 VNB 0.09fF
C2005 a_6789_1004.n0 VNB 0.56fF
C2006 a_6789_1004.n1 VNB 0.56fF
C2007 a_6789_1004.n2 VNB 0.65fF
C2008 a_6789_1004.n3 VNB 0.21fF
C2009 a_6789_1004.n4 VNB 0.39fF
C2010 a_6789_1004.n5 VNB 0.46fF
C2011 a_6789_1004.n6 VNB 0.57fF
C2012 a_6789_1004.n7 VNB 0.66fF
C2013 a_6789_1004.n8 VNB 0.09fF
C2014 a_6789_1004.n9 VNB 0.22fF
C2015 a_6789_1004.n10 VNB 0.05fF
C2016 a_6884_182.n0 VNB 0.07fF
C2017 a_6884_182.n1 VNB 0.13fF
C2018 a_6884_182.n2 VNB 0.07fF
C2019 a_6884_182.n3 VNB 0.02fF
C2020 a_6884_182.n4 VNB 0.03fF
C2021 a_6884_182.n5 VNB 0.02fF
C2022 a_6884_182.n6 VNB 0.05fF
C2023 a_6884_182.n7 VNB 0.05fF
C2024 a_6884_182.n8 VNB 0.06fF
C2025 a_6884_182.n9 VNB 0.07fF
C2026 a_6884_182.n10 VNB 0.07fF
C2027 a_6884_182.n11 VNB 0.03fF
C2028 a_6884_182.n12 VNB 0.01fF
C2029 a_6884_182.n13 VNB 0.11fF
C2030 a_6884_182.t0 VNB 0.28fF
C2031 a_6149_943.n0 VNB 0.07fF
C2032 a_6149_943.n1 VNB 0.95fF
C2033 a_6149_943.n2 VNB 1.13fF
C2034 a_6149_943.n3 VNB 0.52fF
C2035 a_6149_943.n4 VNB 0.64fF
C2036 a_6149_943.t10 VNB 0.98fF
C2037 a_6149_943.n5 VNB 0.73fF
C2038 a_6149_943.n6 VNB 0.64fF
C2039 a_6149_943.t5 VNB 0.98fF
C2040 a_6149_943.n7 VNB 0.65fF
C2041 a_6149_943.n8 VNB 0.64fF
C2042 a_6149_943.t13 VNB 0.98fF
C2043 a_6149_943.n9 VNB 0.68fF
C2044 a_6149_943.n10 VNB 2.05fF
C2045 a_6149_943.n11 VNB 2.77fF
C2046 a_6149_943.n12 VNB 0.75fF
C2047 a_6149_943.n13 VNB 0.06fF
C2048 a_6149_943.n14 VNB 0.56fF
C2049 a_6149_943.n15 VNB 0.10fF
.ends
