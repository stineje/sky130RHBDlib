* SPICE3 file created from NAND3X1.ext - technology: sky130A

.subckt NAND3X1 Y A B C VDD GND
X0 VDD B Y VDD pshort w=2 l=0.15 M=2
X1 GND A a_91_75 GND nshort w=3 l=0.15
X2 VDD C Y VDD pshort w=2 l=0.15 M=2
X3 a_372_182 B a_91_75 GND nshort w=3 l=0.15
X4 Y A VDD VDD pshort w=2 l=0.15 M=2
X5 Y C a_372_182 GND nshort w=3 l=0.15
C0 VDD GND 2.67fF
.ends
