magic
tech sky130A
magscale 1 2
timestamp 1645210163
use sky130_fd_pr__hvdfl1sd2__example_55959141808488  sky130_fd_pr__hvdfl1sd2__example_55959141808488_0
timestamp 1645210163
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808488  sky130_fd_pr__hvdfl1sd2__example_55959141808488_1
timestamp 1645210163
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 29 128 29 0 FreeSans 300 0 0 0 D
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 8082524
string GDS_START 8081594
<< end >>
