* SPICE3 file created from TMRDFFSNRNQX1.ext - technology: sky130A

.subckt TMRDFFSNRNQX1 Q SN RN D CLK VPB VNB
M1000 a_4447_943.t3 SN VPB.t77 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VPB.t95 CLK a_6371_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_7333_943.t3 RN VPB.t51 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t47 D a_6049_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VNB a_6049_1004.t8 a_6825_75.t0 nshort w=-1.605u l=1.765u
+  ad=4.9019p pd=41.07u as=0p ps=0u
M1005 a_7973_1004.t3 SN VPB.t78 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_18197_1005.t3 a_10219_943.t7 a_17708_181.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t37 a_4447_943.t7 a_17533_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VNB a_4125_1004.t8 a_4901_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPB.t46 D a_277_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t43 D a_11821_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VNB a_4447_943.t15 a_17428_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t64 RN a_15669_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_599_943.t3 CLK VPB.t88 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPB.t57 RN a_9897_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPB.t97 CLK a_1561_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_11821_1004.t5 a_12143_943.t8 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t50 a_13105_943.t7 a_13745_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VNB D a_11635_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPB.t9 a_277_1004.t7 a_2201_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_7333_943.t6 CLK VPB.t86 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_10219_943.t1 SN VPB.t72 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t83 a_7333_943.t7 a_6371_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPB.t90 CLK a_12143_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPB.t108 a_17708_181.t7 Q.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_13105_943.t3 RN VPB.t68 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VNB a_6049_1004.t10 a_7787_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1027 VNB a_6371_943.t10 a_9711_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1028 VNB D a_5863_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB.t52 RN a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_6371_943.t6 a_6049_1004.t7 VPB.t107 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPB.t25 a_7973_1004.t7 a_7333_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPB.t112 a_9897_1004.t7 a_10219_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_17533_1005.t3 a_4447_943.t9 VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_12143_943.t5 CLK VPB.t87 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_599_943.t6 a_1561_943.t8 VPB.t104 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_15991_943.t0 a_15669_1004.t8 VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPB.t61 RN a_1561_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_9897_1004.t6 a_6371_943.t7 VPB.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VNB a_11821_1004.t9 a_12597_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_4125_1004.t3 a_599_943.t7 VPB.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPB.t80 SN a_2201_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VNB a_13745_1004.t9 a_14521_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_4125_1004.t5 a_4447_943.t10 VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 VNB a_9897_1004.t9 a_10673_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPB.t100 a_6371_943.t8 a_6049_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_18197_1005.t6 a_4447_943.t11 a_17533_1005.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_1561_943.t4 CLK VPB.t96 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 VNB a_7973_1004.t9 a_8749_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPB.t49 a_599_943.t8 a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 VNB D a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_13745_1004.t4 SN VPB.t69 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 a_17533_1005.t2 a_10219_943.t8 VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 Q a_17708_181.t8 VNB.t19 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1054 a_12143_943.t4 a_11821_1004.t7 VPB.t81 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 VPB.t6 a_13745_1004.t7 a_13105_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_15991_943.t3 SN VPB.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_15669_1004.t6 a_12143_943.t10 VPB.t82 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_4125_1004.t1 RN VPB.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 VNB a_11821_1004.t12 a_13559_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1060 VPB.t35 a_1561_943.t11 a_2201_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 VPB.t58 RN a_6049_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_7333_943.t1 a_7973_1004.t8 VPB.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_7973_1004.t5 a_7333_943.t10 VPB.t33 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_9897_1004.t1 a_10219_943.t11 VPB.t32 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 VPB.t105 a_13105_943.t8 a_15991_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 VNB a_12143_943.t7 a_15483_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_1561_943.t0 a_2201_1004.t8 VPB.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_18197_1005.t7 a_15991_943.t8 a_17533_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 VPB.t99 a_4125_1004.t7 a_4447_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_6371_943.t4 CLK VPB.t89 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 VPB.t93 CLK a_7333_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_6049_1004.t0 D VPB.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 a_17708_181.t3 a_10219_943.t12 a_18197_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 a_277_1004.t1 D VPB.t42 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 VPB.t92 CLK a_13105_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 a_15991_943.t6 a_13105_943.t10 VPB.t110 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 VNB a_15669_1004.t7 a_16445_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1078 VPB.t15 a_11821_1004.t8 a_13745_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 a_10219_943.t4 a_7333_943.t12 VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_15669_1004.t3 RN VPB.t63 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 VPB.t24 a_13105_943.t11 a_12143_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 VPB.t8 a_277_1004.t10 a_599_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_9897_1004.t3 RN VPB.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 VPB.t67 RN a_11821_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 VPB.t38 a_1561_943.t12 a_599_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_13745_1004.t0 a_13105_943.t12 VPB.t36 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 VPB.t74 SN a_4447_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_18197_1005.t4 a_15991_943.t9 a_17708_181.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 VPB.t102 a_15991_943.t10 a_15669_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 a_6371_943.t1 a_7333_943.t13 VPB.t26 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 Q.t0 a_17708_181.t9 VPB.t85 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 VPB.t55 RN a_7333_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 VPB.t73 SN a_7973_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_277_1004.t5 RN VPB.t53 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 a_11821_1004.t2 RN VPB.t54 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 VNB a_277_1004.t8 a_2015_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1097 VPB.t70 SN a_13745_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_10219_943.t6 a_9897_1004.t8 VPB.t113 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 VPB.t94 CLK a_599_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 VPB.t106 a_12143_943.t11 a_11821_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 a_1561_943.t1 RN VPB.t60 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 VPB.t22 a_1561_943.t13 a_4447_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_2201_1004.t3 SN VPB.t79 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 VPB.t65 RN a_4125_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 a_12143_943.t0 a_13105_943.t14 VPB.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VPB.t28 a_6049_1004.t9 a_7973_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 VPB.t62 RN a_13105_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 a_599_943.t4 a_277_1004.t11 VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 a_277_1004.t0 a_599_943.t10 VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_11821_1004.t0 D VPB.t44 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 VNB a_2201_1004.t7 a_2977_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1112 VNB a_15991_943.t12 a_18760_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1113 VNB a_4447_943.t12 a_18094_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1114 a_13105_943.t0 a_13745_1004.t8 VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 VPB.t48 a_15669_1004.t9 a_15991_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 VNB a_277_1004.t9 a_1053_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_7973_1004.t0 a_6049_1004.t11 VPB.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 VPB.t101 a_6371_943.t11 a_9897_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_2201_1004.t5 a_277_1004.t12 VPB.t40 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 VPB.t2 a_7333_943.t14 a_10219_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 a_2201_1004.t0 a_1561_943.t14 VPB.t103 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 VPB.t39 a_599_943.t12 a_4125_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 VPB.t31 a_4447_943.t13 a_4125_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1124 a_6049_1004.t2 RN VPB.t59 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1125 a_17533_1005.t5 a_4447_943.t14 a_18197_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1126 a_4447_943.t4 a_4125_1004.t9 VPB.t98 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1127 VPB.t27 a_6049_1004.t12 a_6371_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1128 a_4447_943.t6 a_1561_943.t15 VPB.t109 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1129 VNB a_599_943.t9 a_3939_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1130 a_15669_1004.t0 a_15991_943.t13 VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1131 VPB.t41 a_11821_1004.t10 a_12143_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1132 VPB.t29 a_10219_943.t14 a_17533_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1133 a_13105_943.t5 CLK VPB.t91 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1134 VPB.t76 SN a_15991_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1135 VPB.t71 SN a_10219_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1136 a_13745_1004.t5 a_11821_1004.t11 VPB.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1137 VPB.t12 a_12143_943.t12 a_15669_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1138 a_6049_1004.t4 a_6371_943.t12 VPB.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1139 VPB.t34 a_7333_943.t15 a_7973_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1140 VPB.t17 a_10219_943.t15 a_9897_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1141 VPB.t111 a_2201_1004.t9 a_1561_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1142 a_17708_181.t0 a_15991_943.t14 a_18197_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1143 a_17533_1005.t0 a_15991_943.t15 a_18197_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB Q 0.78fF
C1 VPB D 2.79fF
C2 VPB RN 0.48fF
C3 VPB SN 0.30fF
C4 VPB CLK 3.56fF
C5 D RN 2.37fF
C6 D SN 2.48fF
C7 D CLK 11.99fF
C8 RN SN 5.86fF
C9 RN CLK 1.03fF
C10 SN CLK 2.51fF
R0 VPB VPB.n1729 126.832
R1 VPB.n40 VPB.n38 94.117
R2 VPB.n1651 VPB.n1649 94.117
R3 VPB.n1568 VPB.n1566 94.117
R4 VPB.n1485 VPB.n1483 94.117
R5 VPB.n1402 VPB.n1400 94.117
R6 VPB.n1319 VPB.n1317 94.117
R7 VPB.n1236 VPB.n1234 94.117
R8 VPB.n1153 VPB.n1151 94.117
R9 VPB.n1070 VPB.n1068 94.117
R10 VPB.n987 VPB.n985 94.117
R11 VPB.n114 VPB.n112 94.117
R12 VPB.n884 VPB.n882 94.117
R13 VPB.n801 VPB.n799 94.117
R14 VPB.n718 VPB.n716 94.117
R15 VPB.n635 VPB.n633 94.117
R16 VPB.n552 VPB.n550 94.117
R17 VPB.n469 VPB.n467 94.117
R18 VPB.n386 VPB.n384 94.117
R19 VPB.n323 VPB.n321 94.117
R20 VPB.n268 VPB.n266 94.117
R21 VPB.n213 VPB.n211 91.036
R22 VPB.n399 VPB.n398 80.104
R23 VPB.n482 VPB.n481 80.104
R24 VPB.n565 VPB.n564 80.104
R25 VPB.n648 VPB.n647 80.104
R26 VPB.n731 VPB.n730 80.104
R27 VPB.n814 VPB.n813 80.104
R28 VPB.n897 VPB.n896 80.104
R29 VPB.n124 VPB.n123 80.104
R30 VPB.n1000 VPB.n999 80.104
R31 VPB.n1083 VPB.n1082 80.104
R32 VPB.n1166 VPB.n1165 80.104
R33 VPB.n1249 VPB.n1248 80.104
R34 VPB.n1332 VPB.n1331 80.104
R35 VPB.n1415 VPB.n1414 80.104
R36 VPB.n1498 VPB.n1497 80.104
R37 VPB.n1581 VPB.n1580 80.104
R38 VPB.n1664 VPB.n1663 80.104
R39 VPB.n50 VPB.n49 80.104
R40 VPB.n174 VPB.n168 76.136
R41 VPB.n174 VPB.n173 76
R42 VPB.n178 VPB.n177 76
R43 VPB.n184 VPB.n183 76
R44 VPB.n188 VPB.n187 76
R45 VPB.n215 VPB.n214 76
R46 VPB.n219 VPB.n218 76
R47 VPB.n223 VPB.n222 76
R48 VPB.n227 VPB.n226 76
R49 VPB.n231 VPB.n230 76
R50 VPB.n235 VPB.n234 76
R51 VPB.n239 VPB.n238 76
R52 VPB.n243 VPB.n242 76
R53 VPB.n270 VPB.n269 76
R54 VPB.n274 VPB.n273 76
R55 VPB.n278 VPB.n277 76
R56 VPB.n282 VPB.n281 76
R57 VPB.n286 VPB.n285 76
R58 VPB.n290 VPB.n289 76
R59 VPB.n294 VPB.n293 76
R60 VPB.n298 VPB.n297 76
R61 VPB.n325 VPB.n324 76
R62 VPB.n330 VPB.n329 76
R63 VPB.n335 VPB.n334 76
R64 VPB.n342 VPB.n341 76
R65 VPB.n347 VPB.n346 76
R66 VPB.n352 VPB.n351 76
R67 VPB.n357 VPB.n356 76
R68 VPB.n361 VPB.n360 76
R69 VPB.n388 VPB.n387 76
R70 VPB.n392 VPB.n391 76
R71 VPB.n397 VPB.n396 76
R72 VPB.n402 VPB.n401 76
R73 VPB.n409 VPB.n408 76
R74 VPB.n414 VPB.n413 76
R75 VPB.n419 VPB.n418 76
R76 VPB.n426 VPB.n425 76
R77 VPB.n431 VPB.n430 76
R78 VPB.n436 VPB.n435 76
R79 VPB.n440 VPB.n439 76
R80 VPB.n444 VPB.n443 76
R81 VPB.n471 VPB.n470 76
R82 VPB.n475 VPB.n474 76
R83 VPB.n480 VPB.n479 76
R84 VPB.n485 VPB.n484 76
R85 VPB.n492 VPB.n491 76
R86 VPB.n497 VPB.n496 76
R87 VPB.n502 VPB.n501 76
R88 VPB.n509 VPB.n508 76
R89 VPB.n514 VPB.n513 76
R90 VPB.n519 VPB.n518 76
R91 VPB.n523 VPB.n522 76
R92 VPB.n527 VPB.n526 76
R93 VPB.n554 VPB.n553 76
R94 VPB.n558 VPB.n557 76
R95 VPB.n563 VPB.n562 76
R96 VPB.n568 VPB.n567 76
R97 VPB.n575 VPB.n574 76
R98 VPB.n580 VPB.n579 76
R99 VPB.n585 VPB.n584 76
R100 VPB.n592 VPB.n591 76
R101 VPB.n597 VPB.n596 76
R102 VPB.n602 VPB.n601 76
R103 VPB.n606 VPB.n605 76
R104 VPB.n610 VPB.n609 76
R105 VPB.n637 VPB.n636 76
R106 VPB.n641 VPB.n640 76
R107 VPB.n646 VPB.n645 76
R108 VPB.n651 VPB.n650 76
R109 VPB.n658 VPB.n657 76
R110 VPB.n663 VPB.n662 76
R111 VPB.n668 VPB.n667 76
R112 VPB.n675 VPB.n674 76
R113 VPB.n680 VPB.n679 76
R114 VPB.n685 VPB.n684 76
R115 VPB.n689 VPB.n688 76
R116 VPB.n693 VPB.n692 76
R117 VPB.n720 VPB.n719 76
R118 VPB.n724 VPB.n723 76
R119 VPB.n729 VPB.n728 76
R120 VPB.n734 VPB.n733 76
R121 VPB.n741 VPB.n740 76
R122 VPB.n746 VPB.n745 76
R123 VPB.n751 VPB.n750 76
R124 VPB.n758 VPB.n757 76
R125 VPB.n763 VPB.n762 76
R126 VPB.n768 VPB.n767 76
R127 VPB.n772 VPB.n771 76
R128 VPB.n776 VPB.n775 76
R129 VPB.n803 VPB.n802 76
R130 VPB.n807 VPB.n806 76
R131 VPB.n812 VPB.n811 76
R132 VPB.n817 VPB.n816 76
R133 VPB.n824 VPB.n823 76
R134 VPB.n829 VPB.n828 76
R135 VPB.n834 VPB.n833 76
R136 VPB.n841 VPB.n840 76
R137 VPB.n846 VPB.n845 76
R138 VPB.n851 VPB.n850 76
R139 VPB.n855 VPB.n854 76
R140 VPB.n859 VPB.n858 76
R141 VPB.n886 VPB.n885 76
R142 VPB.n890 VPB.n889 76
R143 VPB.n895 VPB.n894 76
R144 VPB.n900 VPB.n899 76
R145 VPB.n907 VPB.n906 76
R146 VPB.n912 VPB.n911 76
R147 VPB.n917 VPB.n916 76
R148 VPB.n924 VPB.n923 76
R149 VPB.n929 VPB.n928 76
R150 VPB.n934 VPB.n933 76
R151 VPB.n949 VPB.n945 76
R152 VPB.n954 VPB.n953 76
R153 VPB.n958 VPB.n957 76
R154 VPB.n962 VPB.n961 76
R155 VPB.n989 VPB.n988 76
R156 VPB.n993 VPB.n992 76
R157 VPB.n998 VPB.n997 76
R158 VPB.n1003 VPB.n1002 76
R159 VPB.n1010 VPB.n1009 76
R160 VPB.n1015 VPB.n1014 76
R161 VPB.n1020 VPB.n1019 76
R162 VPB.n1027 VPB.n1026 76
R163 VPB.n1032 VPB.n1031 76
R164 VPB.n1037 VPB.n1036 76
R165 VPB.n1041 VPB.n1040 76
R166 VPB.n1045 VPB.n1044 76
R167 VPB.n1072 VPB.n1071 76
R168 VPB.n1076 VPB.n1075 76
R169 VPB.n1081 VPB.n1080 76
R170 VPB.n1086 VPB.n1085 76
R171 VPB.n1093 VPB.n1092 76
R172 VPB.n1098 VPB.n1097 76
R173 VPB.n1103 VPB.n1102 76
R174 VPB.n1110 VPB.n1109 76
R175 VPB.n1115 VPB.n1114 76
R176 VPB.n1120 VPB.n1119 76
R177 VPB.n1124 VPB.n1123 76
R178 VPB.n1128 VPB.n1127 76
R179 VPB.n1155 VPB.n1154 76
R180 VPB.n1159 VPB.n1158 76
R181 VPB.n1164 VPB.n1163 76
R182 VPB.n1169 VPB.n1168 76
R183 VPB.n1176 VPB.n1175 76
R184 VPB.n1181 VPB.n1180 76
R185 VPB.n1186 VPB.n1185 76
R186 VPB.n1193 VPB.n1192 76
R187 VPB.n1198 VPB.n1197 76
R188 VPB.n1203 VPB.n1202 76
R189 VPB.n1207 VPB.n1206 76
R190 VPB.n1211 VPB.n1210 76
R191 VPB.n1238 VPB.n1237 76
R192 VPB.n1242 VPB.n1241 76
R193 VPB.n1247 VPB.n1246 76
R194 VPB.n1252 VPB.n1251 76
R195 VPB.n1259 VPB.n1258 76
R196 VPB.n1264 VPB.n1263 76
R197 VPB.n1269 VPB.n1268 76
R198 VPB.n1276 VPB.n1275 76
R199 VPB.n1281 VPB.n1280 76
R200 VPB.n1286 VPB.n1285 76
R201 VPB.n1290 VPB.n1289 76
R202 VPB.n1294 VPB.n1293 76
R203 VPB.n1321 VPB.n1320 76
R204 VPB.n1325 VPB.n1324 76
R205 VPB.n1330 VPB.n1329 76
R206 VPB.n1335 VPB.n1334 76
R207 VPB.n1342 VPB.n1341 76
R208 VPB.n1347 VPB.n1346 76
R209 VPB.n1352 VPB.n1351 76
R210 VPB.n1359 VPB.n1358 76
R211 VPB.n1364 VPB.n1363 76
R212 VPB.n1369 VPB.n1368 76
R213 VPB.n1373 VPB.n1372 76
R214 VPB.n1377 VPB.n1376 76
R215 VPB.n1404 VPB.n1403 76
R216 VPB.n1408 VPB.n1407 76
R217 VPB.n1413 VPB.n1412 76
R218 VPB.n1418 VPB.n1417 76
R219 VPB.n1425 VPB.n1424 76
R220 VPB.n1430 VPB.n1429 76
R221 VPB.n1435 VPB.n1434 76
R222 VPB.n1442 VPB.n1441 76
R223 VPB.n1447 VPB.n1446 76
R224 VPB.n1452 VPB.n1451 76
R225 VPB.n1456 VPB.n1455 76
R226 VPB.n1460 VPB.n1459 76
R227 VPB.n1487 VPB.n1486 76
R228 VPB.n1491 VPB.n1490 76
R229 VPB.n1496 VPB.n1495 76
R230 VPB.n1501 VPB.n1500 76
R231 VPB.n1508 VPB.n1507 76
R232 VPB.n1513 VPB.n1512 76
R233 VPB.n1518 VPB.n1517 76
R234 VPB.n1525 VPB.n1524 76
R235 VPB.n1530 VPB.n1529 76
R236 VPB.n1535 VPB.n1534 76
R237 VPB.n1539 VPB.n1538 76
R238 VPB.n1543 VPB.n1542 76
R239 VPB.n1570 VPB.n1569 76
R240 VPB.n1574 VPB.n1573 76
R241 VPB.n1579 VPB.n1578 76
R242 VPB.n1584 VPB.n1583 76
R243 VPB.n1591 VPB.n1590 76
R244 VPB.n1596 VPB.n1595 76
R245 VPB.n1601 VPB.n1600 76
R246 VPB.n1608 VPB.n1607 76
R247 VPB.n1613 VPB.n1612 76
R248 VPB.n1618 VPB.n1617 76
R249 VPB.n1622 VPB.n1621 76
R250 VPB.n1626 VPB.n1625 76
R251 VPB.n1653 VPB.n1652 76
R252 VPB.n1657 VPB.n1656 76
R253 VPB.n1662 VPB.n1661 76
R254 VPB.n1667 VPB.n1666 76
R255 VPB.n1674 VPB.n1673 76
R256 VPB.n1679 VPB.n1678 76
R257 VPB.n1684 VPB.n1683 76
R258 VPB.n1691 VPB.n1690 76
R259 VPB.n1696 VPB.n1695 76
R260 VPB.n1701 VPB.n1700 76
R261 VPB.n1705 VPB.n1704 76
R262 VPB.n1709 VPB.n1708 76
R263 VPB.n1722 VPB.n1721 76
R264 VPB.n428 VPB.n427 75.654
R265 VPB.n511 VPB.n510 75.654
R266 VPB.n594 VPB.n593 75.654
R267 VPB.n677 VPB.n676 75.654
R268 VPB.n760 VPB.n759 75.654
R269 VPB.n843 VPB.n842 75.654
R270 VPB.n926 VPB.n925 75.654
R271 VPB.n947 VPB.n946 75.654
R272 VPB.n1029 VPB.n1028 75.654
R273 VPB.n1112 VPB.n1111 75.654
R274 VPB.n1195 VPB.n1194 75.654
R275 VPB.n1278 VPB.n1277 75.654
R276 VPB.n1361 VPB.n1360 75.654
R277 VPB.n1444 VPB.n1443 75.654
R278 VPB.n1527 VPB.n1526 75.654
R279 VPB.n1610 VPB.n1609 75.654
R280 VPB.n1693 VPB.n1692 75.654
R281 VPB.n72 VPB.n71 75.654
R282 VPB.n181 VPB.n180 68.979
R283 VPB.n171 VPB.n170 64.528
R284 VPB.n22 VPB.n21 61.764
R285 VPB.n1633 VPB.n1632 61.764
R286 VPB.n1550 VPB.n1549 61.764
R287 VPB.n1467 VPB.n1466 61.764
R288 VPB.n1384 VPB.n1383 61.764
R289 VPB.n1301 VPB.n1300 61.764
R290 VPB.n1218 VPB.n1217 61.764
R291 VPB.n1135 VPB.n1134 61.764
R292 VPB.n1052 VPB.n1051 61.764
R293 VPB.n969 VPB.n968 61.764
R294 VPB.n90 VPB.n89 61.764
R295 VPB.n866 VPB.n865 61.764
R296 VPB.n783 VPB.n782 61.764
R297 VPB.n700 VPB.n699 61.764
R298 VPB.n617 VPB.n616 61.764
R299 VPB.n534 VPB.n533 61.764
R300 VPB.n451 VPB.n450 61.764
R301 VPB.n368 VPB.n367 61.764
R302 VPB.n305 VPB.n304 61.764
R303 VPB.n250 VPB.n249 61.764
R304 VPB.n195 VPB.n194 61.764
R305 VPB.n353 VPB.t0 55.465
R306 VPB.n326 VPB.t29 55.465
R307 VPB.n78 VPB.t42 55.106
R308 VPB.n1697 VPB.t7 55.106
R309 VPB.n1614 VPB.t40 55.106
R310 VPB.n1531 VPB.t16 55.106
R311 VPB.n1448 VPB.t21 55.106
R312 VPB.n1365 VPB.t98 55.106
R313 VPB.n1282 VPB.t45 55.106
R314 VPB.n1199 VPB.t107 55.106
R315 VPB.n1116 VPB.t13 55.106
R316 VPB.n1033 VPB.t30 55.106
R317 VPB.n950 VPB.t19 55.106
R318 VPB.n930 VPB.t113 55.106
R319 VPB.n847 VPB.t44 55.106
R320 VPB.n764 VPB.t81 55.106
R321 VPB.n681 VPB.t10 55.106
R322 VPB.n598 VPB.t5 55.106
R323 VPB.n515 VPB.t82 55.106
R324 VPB.n432 VPB.t18 55.106
R325 VPB.n179 VPB.t85 55.106
R326 VPB.n169 VPB.t108 55.106
R327 VPB.n45 VPB.t49 55.106
R328 VPB.n1658 VPB.t38 55.106
R329 VPB.n1575 VPB.t35 55.106
R330 VPB.n1492 VPB.t61 55.106
R331 VPB.n1409 VPB.t31 55.106
R332 VPB.n1326 VPB.t22 55.106
R333 VPB.n1243 VPB.t100 55.106
R334 VPB.n1160 VPB.t83 55.106
R335 VPB.n1077 VPB.t34 55.106
R336 VPB.n994 VPB.t55 55.106
R337 VPB.n119 VPB.t17 55.106
R338 VPB.n891 VPB.t2 55.106
R339 VPB.n808 VPB.t106 55.106
R340 VPB.n725 VPB.t24 55.106
R341 VPB.n642 VPB.t50 55.106
R342 VPB.n559 VPB.t62 55.106
R343 VPB.n476 VPB.t102 55.106
R344 VPB.n393 VPB.t105 55.106
R345 VPB.n332 VPB.n331 48.952
R346 VPB.n406 VPB.n405 48.952
R347 VPB.n489 VPB.n488 48.952
R348 VPB.n572 VPB.n571 48.952
R349 VPB.n655 VPB.n654 48.952
R350 VPB.n738 VPB.n737 48.952
R351 VPB.n821 VPB.n820 48.952
R352 VPB.n904 VPB.n903 48.952
R353 VPB.n128 VPB.n127 48.952
R354 VPB.n1007 VPB.n1006 48.952
R355 VPB.n1090 VPB.n1089 48.952
R356 VPB.n1173 VPB.n1172 48.952
R357 VPB.n1256 VPB.n1255 48.952
R358 VPB.n1339 VPB.n1338 48.952
R359 VPB.n1422 VPB.n1421 48.952
R360 VPB.n1505 VPB.n1504 48.952
R361 VPB.n1588 VPB.n1587 48.952
R362 VPB.n1671 VPB.n1670 48.952
R363 VPB.n54 VPB.n53 48.952
R364 VPB.n349 VPB.n348 44.502
R365 VPB.n423 VPB.n422 44.502
R366 VPB.n506 VPB.n505 44.502
R367 VPB.n589 VPB.n588 44.502
R368 VPB.n672 VPB.n671 44.502
R369 VPB.n755 VPB.n754 44.502
R370 VPB.n838 VPB.n837 44.502
R371 VPB.n921 VPB.n920 44.502
R372 VPB.n142 VPB.n141 44.502
R373 VPB.n1024 VPB.n1023 44.502
R374 VPB.n1107 VPB.n1106 44.502
R375 VPB.n1190 VPB.n1189 44.502
R376 VPB.n1273 VPB.n1272 44.502
R377 VPB.n1356 VPB.n1355 44.502
R378 VPB.n1439 VPB.n1438 44.502
R379 VPB.n1522 VPB.n1521 44.502
R380 VPB.n1605 VPB.n1604 44.502
R381 VPB.n1688 VPB.n1687 44.502
R382 VPB.n68 VPB.n67 44.502
R383 VPB.n337 VPB.n336 41.183
R384 VPB.n66 VPB.n14 40.824
R385 VPB.n57 VPB.n15 40.824
R386 VPB.n1686 VPB.n1685 40.824
R387 VPB.n1669 VPB.n1668 40.824
R388 VPB.n1603 VPB.n1602 40.824
R389 VPB.n1586 VPB.n1585 40.824
R390 VPB.n1520 VPB.n1519 40.824
R391 VPB.n1503 VPB.n1502 40.824
R392 VPB.n1437 VPB.n1436 40.824
R393 VPB.n1420 VPB.n1419 40.824
R394 VPB.n1354 VPB.n1353 40.824
R395 VPB.n1337 VPB.n1336 40.824
R396 VPB.n1271 VPB.n1270 40.824
R397 VPB.n1254 VPB.n1253 40.824
R398 VPB.n1188 VPB.n1187 40.824
R399 VPB.n1171 VPB.n1170 40.824
R400 VPB.n1105 VPB.n1104 40.824
R401 VPB.n1088 VPB.n1087 40.824
R402 VPB.n1022 VPB.n1021 40.824
R403 VPB.n1005 VPB.n1004 40.824
R404 VPB.n140 VPB.n82 40.824
R405 VPB.n131 VPB.n83 40.824
R406 VPB.n919 VPB.n918 40.824
R407 VPB.n902 VPB.n901 40.824
R408 VPB.n836 VPB.n835 40.824
R409 VPB.n819 VPB.n818 40.824
R410 VPB.n753 VPB.n752 40.824
R411 VPB.n736 VPB.n735 40.824
R412 VPB.n670 VPB.n669 40.824
R413 VPB.n653 VPB.n652 40.824
R414 VPB.n587 VPB.n586 40.824
R415 VPB.n570 VPB.n569 40.824
R416 VPB.n504 VPB.n503 40.824
R417 VPB.n487 VPB.n486 40.824
R418 VPB.n421 VPB.n420 40.824
R419 VPB.n404 VPB.n403 40.824
R420 VPB.n1726 VPB.n1722 20.452
R421 VPB.n168 VPB.n165 20.452
R422 VPB.n339 VPB.n338 17.801
R423 VPB.n411 VPB.n410 17.801
R424 VPB.n494 VPB.n493 17.801
R425 VPB.n577 VPB.n576 17.801
R426 VPB.n660 VPB.n659 17.801
R427 VPB.n743 VPB.n742 17.801
R428 VPB.n826 VPB.n825 17.801
R429 VPB.n909 VPB.n908 17.801
R430 VPB.n133 VPB.n132 17.801
R431 VPB.n1012 VPB.n1011 17.801
R432 VPB.n1095 VPB.n1094 17.801
R433 VPB.n1178 VPB.n1177 17.801
R434 VPB.n1261 VPB.n1260 17.801
R435 VPB.n1344 VPB.n1343 17.801
R436 VPB.n1427 VPB.n1426 17.801
R437 VPB.n1510 VPB.n1509 17.801
R438 VPB.n1593 VPB.n1592 17.801
R439 VPB.n1676 VPB.n1675 17.801
R440 VPB.n59 VPB.n58 17.801
R441 VPB.n14 VPB.t53 14.282
R442 VPB.n14 VPB.t46 14.282
R443 VPB.n15 VPB.t20 14.282
R444 VPB.n15 VPB.t52 14.282
R445 VPB.n1685 VPB.t88 14.282
R446 VPB.n1685 VPB.t8 14.282
R447 VPB.n1668 VPB.t104 14.282
R448 VPB.n1668 VPB.t94 14.282
R449 VPB.n1602 VPB.t79 14.282
R450 VPB.n1602 VPB.t9 14.282
R451 VPB.n1585 VPB.t103 14.282
R452 VPB.n1585 VPB.t80 14.282
R453 VPB.n1519 VPB.t96 14.282
R454 VPB.n1519 VPB.t111 14.282
R455 VPB.n1502 VPB.t60 14.282
R456 VPB.n1502 VPB.t97 14.282
R457 VPB.n1436 VPB.t66 14.282
R458 VPB.n1436 VPB.t39 14.282
R459 VPB.n1419 VPB.t3 14.282
R460 VPB.n1419 VPB.t65 14.282
R461 VPB.n1353 VPB.t77 14.282
R462 VPB.n1353 VPB.t99 14.282
R463 VPB.n1336 VPB.t109 14.282
R464 VPB.n1336 VPB.t74 14.282
R465 VPB.n1270 VPB.t59 14.282
R466 VPB.n1270 VPB.t47 14.282
R467 VPB.n1253 VPB.t84 14.282
R468 VPB.n1253 VPB.t58 14.282
R469 VPB.n1187 VPB.t89 14.282
R470 VPB.n1187 VPB.t27 14.282
R471 VPB.n1170 VPB.t26 14.282
R472 VPB.n1170 VPB.t95 14.282
R473 VPB.n1104 VPB.t78 14.282
R474 VPB.n1104 VPB.t28 14.282
R475 VPB.n1087 VPB.t33 14.282
R476 VPB.n1087 VPB.t73 14.282
R477 VPB.n1021 VPB.t86 14.282
R478 VPB.n1021 VPB.t25 14.282
R479 VPB.n1004 VPB.t51 14.282
R480 VPB.n1004 VPB.t93 14.282
R481 VPB.n82 VPB.t56 14.282
R482 VPB.n82 VPB.t101 14.282
R483 VPB.n83 VPB.t32 14.282
R484 VPB.n83 VPB.t57 14.282
R485 VPB.n918 VPB.t72 14.282
R486 VPB.n918 VPB.t112 14.282
R487 VPB.n901 VPB.t11 14.282
R488 VPB.n901 VPB.t71 14.282
R489 VPB.n835 VPB.t54 14.282
R490 VPB.n835 VPB.t43 14.282
R491 VPB.n818 VPB.t1 14.282
R492 VPB.n818 VPB.t67 14.282
R493 VPB.n752 VPB.t87 14.282
R494 VPB.n752 VPB.t41 14.282
R495 VPB.n735 VPB.t23 14.282
R496 VPB.n735 VPB.t90 14.282
R497 VPB.n669 VPB.t69 14.282
R498 VPB.n669 VPB.t15 14.282
R499 VPB.n652 VPB.t36 14.282
R500 VPB.n652 VPB.t70 14.282
R501 VPB.n586 VPB.t91 14.282
R502 VPB.n586 VPB.t6 14.282
R503 VPB.n569 VPB.t68 14.282
R504 VPB.n569 VPB.t92 14.282
R505 VPB.n503 VPB.t63 14.282
R506 VPB.n503 VPB.t12 14.282
R507 VPB.n486 VPB.t4 14.282
R508 VPB.n486 VPB.t64 14.282
R509 VPB.n420 VPB.t75 14.282
R510 VPB.n420 VPB.t48 14.282
R511 VPB.n403 VPB.t110 14.282
R512 VPB.n403 VPB.t76 14.282
R513 VPB.n336 VPB.t14 14.282
R514 VPB.n336 VPB.t37 14.282
R515 VPB.n168 VPB.n167 13.653
R516 VPB.n167 VPB.n166 13.653
R517 VPB.n173 VPB.n172 13.653
R518 VPB.n172 VPB.n171 13.653
R519 VPB.n177 VPB.n176 13.653
R520 VPB.n176 VPB.n175 13.653
R521 VPB.n183 VPB.n182 13.653
R522 VPB.n182 VPB.n181 13.653
R523 VPB.n187 VPB.n186 13.653
R524 VPB.n186 VPB.n185 13.653
R525 VPB.n214 VPB.n213 13.653
R526 VPB.n213 VPB.n212 13.653
R527 VPB.n218 VPB.n217 13.653
R528 VPB.n217 VPB.n216 13.653
R529 VPB.n222 VPB.n221 13.653
R530 VPB.n221 VPB.n220 13.653
R531 VPB.n226 VPB.n225 13.653
R532 VPB.n225 VPB.n224 13.653
R533 VPB.n230 VPB.n229 13.653
R534 VPB.n229 VPB.n228 13.653
R535 VPB.n234 VPB.n233 13.653
R536 VPB.n233 VPB.n232 13.653
R537 VPB.n238 VPB.n237 13.653
R538 VPB.n237 VPB.n236 13.653
R539 VPB.n242 VPB.n241 13.653
R540 VPB.n241 VPB.n240 13.653
R541 VPB.n269 VPB.n268 13.653
R542 VPB.n268 VPB.n267 13.653
R543 VPB.n273 VPB.n272 13.653
R544 VPB.n272 VPB.n271 13.653
R545 VPB.n277 VPB.n276 13.653
R546 VPB.n276 VPB.n275 13.653
R547 VPB.n281 VPB.n280 13.653
R548 VPB.n280 VPB.n279 13.653
R549 VPB.n285 VPB.n284 13.653
R550 VPB.n284 VPB.n283 13.653
R551 VPB.n289 VPB.n288 13.653
R552 VPB.n288 VPB.n287 13.653
R553 VPB.n293 VPB.n292 13.653
R554 VPB.n292 VPB.n291 13.653
R555 VPB.n297 VPB.n296 13.653
R556 VPB.n296 VPB.n295 13.653
R557 VPB.n324 VPB.n323 13.653
R558 VPB.n323 VPB.n322 13.653
R559 VPB.n329 VPB.n328 13.653
R560 VPB.n328 VPB.n327 13.653
R561 VPB.n334 VPB.n333 13.653
R562 VPB.n333 VPB.n332 13.653
R563 VPB.n341 VPB.n340 13.653
R564 VPB.n340 VPB.n339 13.653
R565 VPB.n346 VPB.n345 13.653
R566 VPB.n345 VPB.n344 13.653
R567 VPB.n351 VPB.n350 13.653
R568 VPB.n350 VPB.n349 13.653
R569 VPB.n356 VPB.n355 13.653
R570 VPB.n355 VPB.n354 13.653
R571 VPB.n360 VPB.n359 13.653
R572 VPB.n359 VPB.n358 13.653
R573 VPB.n387 VPB.n386 13.653
R574 VPB.n386 VPB.n385 13.653
R575 VPB.n391 VPB.n390 13.653
R576 VPB.n390 VPB.n389 13.653
R577 VPB.n396 VPB.n395 13.653
R578 VPB.n395 VPB.n394 13.653
R579 VPB.n401 VPB.n400 13.653
R580 VPB.n400 VPB.n399 13.653
R581 VPB.n408 VPB.n407 13.653
R582 VPB.n407 VPB.n406 13.653
R583 VPB.n413 VPB.n412 13.653
R584 VPB.n412 VPB.n411 13.653
R585 VPB.n418 VPB.n417 13.653
R586 VPB.n417 VPB.n416 13.653
R587 VPB.n425 VPB.n424 13.653
R588 VPB.n424 VPB.n423 13.653
R589 VPB.n430 VPB.n429 13.653
R590 VPB.n429 VPB.n428 13.653
R591 VPB.n435 VPB.n434 13.653
R592 VPB.n434 VPB.n433 13.653
R593 VPB.n439 VPB.n438 13.653
R594 VPB.n438 VPB.n437 13.653
R595 VPB.n443 VPB.n442 13.653
R596 VPB.n442 VPB.n441 13.653
R597 VPB.n470 VPB.n469 13.653
R598 VPB.n469 VPB.n468 13.653
R599 VPB.n474 VPB.n473 13.653
R600 VPB.n473 VPB.n472 13.653
R601 VPB.n479 VPB.n478 13.653
R602 VPB.n478 VPB.n477 13.653
R603 VPB.n484 VPB.n483 13.653
R604 VPB.n483 VPB.n482 13.653
R605 VPB.n491 VPB.n490 13.653
R606 VPB.n490 VPB.n489 13.653
R607 VPB.n496 VPB.n495 13.653
R608 VPB.n495 VPB.n494 13.653
R609 VPB.n501 VPB.n500 13.653
R610 VPB.n500 VPB.n499 13.653
R611 VPB.n508 VPB.n507 13.653
R612 VPB.n507 VPB.n506 13.653
R613 VPB.n513 VPB.n512 13.653
R614 VPB.n512 VPB.n511 13.653
R615 VPB.n518 VPB.n517 13.653
R616 VPB.n517 VPB.n516 13.653
R617 VPB.n522 VPB.n521 13.653
R618 VPB.n521 VPB.n520 13.653
R619 VPB.n526 VPB.n525 13.653
R620 VPB.n525 VPB.n524 13.653
R621 VPB.n553 VPB.n552 13.653
R622 VPB.n552 VPB.n551 13.653
R623 VPB.n557 VPB.n556 13.653
R624 VPB.n556 VPB.n555 13.653
R625 VPB.n562 VPB.n561 13.653
R626 VPB.n561 VPB.n560 13.653
R627 VPB.n567 VPB.n566 13.653
R628 VPB.n566 VPB.n565 13.653
R629 VPB.n574 VPB.n573 13.653
R630 VPB.n573 VPB.n572 13.653
R631 VPB.n579 VPB.n578 13.653
R632 VPB.n578 VPB.n577 13.653
R633 VPB.n584 VPB.n583 13.653
R634 VPB.n583 VPB.n582 13.653
R635 VPB.n591 VPB.n590 13.653
R636 VPB.n590 VPB.n589 13.653
R637 VPB.n596 VPB.n595 13.653
R638 VPB.n595 VPB.n594 13.653
R639 VPB.n601 VPB.n600 13.653
R640 VPB.n600 VPB.n599 13.653
R641 VPB.n605 VPB.n604 13.653
R642 VPB.n604 VPB.n603 13.653
R643 VPB.n609 VPB.n608 13.653
R644 VPB.n608 VPB.n607 13.653
R645 VPB.n636 VPB.n635 13.653
R646 VPB.n635 VPB.n634 13.653
R647 VPB.n640 VPB.n639 13.653
R648 VPB.n639 VPB.n638 13.653
R649 VPB.n645 VPB.n644 13.653
R650 VPB.n644 VPB.n643 13.653
R651 VPB.n650 VPB.n649 13.653
R652 VPB.n649 VPB.n648 13.653
R653 VPB.n657 VPB.n656 13.653
R654 VPB.n656 VPB.n655 13.653
R655 VPB.n662 VPB.n661 13.653
R656 VPB.n661 VPB.n660 13.653
R657 VPB.n667 VPB.n666 13.653
R658 VPB.n666 VPB.n665 13.653
R659 VPB.n674 VPB.n673 13.653
R660 VPB.n673 VPB.n672 13.653
R661 VPB.n679 VPB.n678 13.653
R662 VPB.n678 VPB.n677 13.653
R663 VPB.n684 VPB.n683 13.653
R664 VPB.n683 VPB.n682 13.653
R665 VPB.n688 VPB.n687 13.653
R666 VPB.n687 VPB.n686 13.653
R667 VPB.n692 VPB.n691 13.653
R668 VPB.n691 VPB.n690 13.653
R669 VPB.n719 VPB.n718 13.653
R670 VPB.n718 VPB.n717 13.653
R671 VPB.n723 VPB.n722 13.653
R672 VPB.n722 VPB.n721 13.653
R673 VPB.n728 VPB.n727 13.653
R674 VPB.n727 VPB.n726 13.653
R675 VPB.n733 VPB.n732 13.653
R676 VPB.n732 VPB.n731 13.653
R677 VPB.n740 VPB.n739 13.653
R678 VPB.n739 VPB.n738 13.653
R679 VPB.n745 VPB.n744 13.653
R680 VPB.n744 VPB.n743 13.653
R681 VPB.n750 VPB.n749 13.653
R682 VPB.n749 VPB.n748 13.653
R683 VPB.n757 VPB.n756 13.653
R684 VPB.n756 VPB.n755 13.653
R685 VPB.n762 VPB.n761 13.653
R686 VPB.n761 VPB.n760 13.653
R687 VPB.n767 VPB.n766 13.653
R688 VPB.n766 VPB.n765 13.653
R689 VPB.n771 VPB.n770 13.653
R690 VPB.n770 VPB.n769 13.653
R691 VPB.n775 VPB.n774 13.653
R692 VPB.n774 VPB.n773 13.653
R693 VPB.n802 VPB.n801 13.653
R694 VPB.n801 VPB.n800 13.653
R695 VPB.n806 VPB.n805 13.653
R696 VPB.n805 VPB.n804 13.653
R697 VPB.n811 VPB.n810 13.653
R698 VPB.n810 VPB.n809 13.653
R699 VPB.n816 VPB.n815 13.653
R700 VPB.n815 VPB.n814 13.653
R701 VPB.n823 VPB.n822 13.653
R702 VPB.n822 VPB.n821 13.653
R703 VPB.n828 VPB.n827 13.653
R704 VPB.n827 VPB.n826 13.653
R705 VPB.n833 VPB.n832 13.653
R706 VPB.n832 VPB.n831 13.653
R707 VPB.n840 VPB.n839 13.653
R708 VPB.n839 VPB.n838 13.653
R709 VPB.n845 VPB.n844 13.653
R710 VPB.n844 VPB.n843 13.653
R711 VPB.n850 VPB.n849 13.653
R712 VPB.n849 VPB.n848 13.653
R713 VPB.n854 VPB.n853 13.653
R714 VPB.n853 VPB.n852 13.653
R715 VPB.n858 VPB.n857 13.653
R716 VPB.n857 VPB.n856 13.653
R717 VPB.n885 VPB.n884 13.653
R718 VPB.n884 VPB.n883 13.653
R719 VPB.n889 VPB.n888 13.653
R720 VPB.n888 VPB.n887 13.653
R721 VPB.n894 VPB.n893 13.653
R722 VPB.n893 VPB.n892 13.653
R723 VPB.n899 VPB.n898 13.653
R724 VPB.n898 VPB.n897 13.653
R725 VPB.n906 VPB.n905 13.653
R726 VPB.n905 VPB.n904 13.653
R727 VPB.n911 VPB.n910 13.653
R728 VPB.n910 VPB.n909 13.653
R729 VPB.n916 VPB.n915 13.653
R730 VPB.n915 VPB.n914 13.653
R731 VPB.n923 VPB.n922 13.653
R732 VPB.n922 VPB.n921 13.653
R733 VPB.n928 VPB.n927 13.653
R734 VPB.n927 VPB.n926 13.653
R735 VPB.n933 VPB.n932 13.653
R736 VPB.n932 VPB.n931 13.653
R737 VPB.n107 VPB.n106 13.653
R738 VPB.n106 VPB.n105 13.653
R739 VPB.n110 VPB.n109 13.653
R740 VPB.n109 VPB.n108 13.653
R741 VPB.n115 VPB.n114 13.653
R742 VPB.n114 VPB.n113 13.653
R743 VPB.n118 VPB.n117 13.653
R744 VPB.n117 VPB.n116 13.653
R745 VPB.n122 VPB.n121 13.653
R746 VPB.n121 VPB.n120 13.653
R747 VPB.n126 VPB.n125 13.653
R748 VPB.n125 VPB.n124 13.653
R749 VPB.n130 VPB.n129 13.653
R750 VPB.n129 VPB.n128 13.653
R751 VPB.n135 VPB.n134 13.653
R752 VPB.n134 VPB.n133 13.653
R753 VPB.n139 VPB.n138 13.653
R754 VPB.n138 VPB.n137 13.653
R755 VPB.n144 VPB.n143 13.653
R756 VPB.n143 VPB.n142 13.653
R757 VPB.n949 VPB.n948 13.653
R758 VPB.n948 VPB.n947 13.653
R759 VPB.n953 VPB.n952 13.653
R760 VPB.n952 VPB.n951 13.653
R761 VPB.n957 VPB.n956 13.653
R762 VPB.n956 VPB.n955 13.653
R763 VPB.n961 VPB.n960 13.653
R764 VPB.n960 VPB.n959 13.653
R765 VPB.n988 VPB.n987 13.653
R766 VPB.n987 VPB.n986 13.653
R767 VPB.n992 VPB.n991 13.653
R768 VPB.n991 VPB.n990 13.653
R769 VPB.n997 VPB.n996 13.653
R770 VPB.n996 VPB.n995 13.653
R771 VPB.n1002 VPB.n1001 13.653
R772 VPB.n1001 VPB.n1000 13.653
R773 VPB.n1009 VPB.n1008 13.653
R774 VPB.n1008 VPB.n1007 13.653
R775 VPB.n1014 VPB.n1013 13.653
R776 VPB.n1013 VPB.n1012 13.653
R777 VPB.n1019 VPB.n1018 13.653
R778 VPB.n1018 VPB.n1017 13.653
R779 VPB.n1026 VPB.n1025 13.653
R780 VPB.n1025 VPB.n1024 13.653
R781 VPB.n1031 VPB.n1030 13.653
R782 VPB.n1030 VPB.n1029 13.653
R783 VPB.n1036 VPB.n1035 13.653
R784 VPB.n1035 VPB.n1034 13.653
R785 VPB.n1040 VPB.n1039 13.653
R786 VPB.n1039 VPB.n1038 13.653
R787 VPB.n1044 VPB.n1043 13.653
R788 VPB.n1043 VPB.n1042 13.653
R789 VPB.n1071 VPB.n1070 13.653
R790 VPB.n1070 VPB.n1069 13.653
R791 VPB.n1075 VPB.n1074 13.653
R792 VPB.n1074 VPB.n1073 13.653
R793 VPB.n1080 VPB.n1079 13.653
R794 VPB.n1079 VPB.n1078 13.653
R795 VPB.n1085 VPB.n1084 13.653
R796 VPB.n1084 VPB.n1083 13.653
R797 VPB.n1092 VPB.n1091 13.653
R798 VPB.n1091 VPB.n1090 13.653
R799 VPB.n1097 VPB.n1096 13.653
R800 VPB.n1096 VPB.n1095 13.653
R801 VPB.n1102 VPB.n1101 13.653
R802 VPB.n1101 VPB.n1100 13.653
R803 VPB.n1109 VPB.n1108 13.653
R804 VPB.n1108 VPB.n1107 13.653
R805 VPB.n1114 VPB.n1113 13.653
R806 VPB.n1113 VPB.n1112 13.653
R807 VPB.n1119 VPB.n1118 13.653
R808 VPB.n1118 VPB.n1117 13.653
R809 VPB.n1123 VPB.n1122 13.653
R810 VPB.n1122 VPB.n1121 13.653
R811 VPB.n1127 VPB.n1126 13.653
R812 VPB.n1126 VPB.n1125 13.653
R813 VPB.n1154 VPB.n1153 13.653
R814 VPB.n1153 VPB.n1152 13.653
R815 VPB.n1158 VPB.n1157 13.653
R816 VPB.n1157 VPB.n1156 13.653
R817 VPB.n1163 VPB.n1162 13.653
R818 VPB.n1162 VPB.n1161 13.653
R819 VPB.n1168 VPB.n1167 13.653
R820 VPB.n1167 VPB.n1166 13.653
R821 VPB.n1175 VPB.n1174 13.653
R822 VPB.n1174 VPB.n1173 13.653
R823 VPB.n1180 VPB.n1179 13.653
R824 VPB.n1179 VPB.n1178 13.653
R825 VPB.n1185 VPB.n1184 13.653
R826 VPB.n1184 VPB.n1183 13.653
R827 VPB.n1192 VPB.n1191 13.653
R828 VPB.n1191 VPB.n1190 13.653
R829 VPB.n1197 VPB.n1196 13.653
R830 VPB.n1196 VPB.n1195 13.653
R831 VPB.n1202 VPB.n1201 13.653
R832 VPB.n1201 VPB.n1200 13.653
R833 VPB.n1206 VPB.n1205 13.653
R834 VPB.n1205 VPB.n1204 13.653
R835 VPB.n1210 VPB.n1209 13.653
R836 VPB.n1209 VPB.n1208 13.653
R837 VPB.n1237 VPB.n1236 13.653
R838 VPB.n1236 VPB.n1235 13.653
R839 VPB.n1241 VPB.n1240 13.653
R840 VPB.n1240 VPB.n1239 13.653
R841 VPB.n1246 VPB.n1245 13.653
R842 VPB.n1245 VPB.n1244 13.653
R843 VPB.n1251 VPB.n1250 13.653
R844 VPB.n1250 VPB.n1249 13.653
R845 VPB.n1258 VPB.n1257 13.653
R846 VPB.n1257 VPB.n1256 13.653
R847 VPB.n1263 VPB.n1262 13.653
R848 VPB.n1262 VPB.n1261 13.653
R849 VPB.n1268 VPB.n1267 13.653
R850 VPB.n1267 VPB.n1266 13.653
R851 VPB.n1275 VPB.n1274 13.653
R852 VPB.n1274 VPB.n1273 13.653
R853 VPB.n1280 VPB.n1279 13.653
R854 VPB.n1279 VPB.n1278 13.653
R855 VPB.n1285 VPB.n1284 13.653
R856 VPB.n1284 VPB.n1283 13.653
R857 VPB.n1289 VPB.n1288 13.653
R858 VPB.n1288 VPB.n1287 13.653
R859 VPB.n1293 VPB.n1292 13.653
R860 VPB.n1292 VPB.n1291 13.653
R861 VPB.n1320 VPB.n1319 13.653
R862 VPB.n1319 VPB.n1318 13.653
R863 VPB.n1324 VPB.n1323 13.653
R864 VPB.n1323 VPB.n1322 13.653
R865 VPB.n1329 VPB.n1328 13.653
R866 VPB.n1328 VPB.n1327 13.653
R867 VPB.n1334 VPB.n1333 13.653
R868 VPB.n1333 VPB.n1332 13.653
R869 VPB.n1341 VPB.n1340 13.653
R870 VPB.n1340 VPB.n1339 13.653
R871 VPB.n1346 VPB.n1345 13.653
R872 VPB.n1345 VPB.n1344 13.653
R873 VPB.n1351 VPB.n1350 13.653
R874 VPB.n1350 VPB.n1349 13.653
R875 VPB.n1358 VPB.n1357 13.653
R876 VPB.n1357 VPB.n1356 13.653
R877 VPB.n1363 VPB.n1362 13.653
R878 VPB.n1362 VPB.n1361 13.653
R879 VPB.n1368 VPB.n1367 13.653
R880 VPB.n1367 VPB.n1366 13.653
R881 VPB.n1372 VPB.n1371 13.653
R882 VPB.n1371 VPB.n1370 13.653
R883 VPB.n1376 VPB.n1375 13.653
R884 VPB.n1375 VPB.n1374 13.653
R885 VPB.n1403 VPB.n1402 13.653
R886 VPB.n1402 VPB.n1401 13.653
R887 VPB.n1407 VPB.n1406 13.653
R888 VPB.n1406 VPB.n1405 13.653
R889 VPB.n1412 VPB.n1411 13.653
R890 VPB.n1411 VPB.n1410 13.653
R891 VPB.n1417 VPB.n1416 13.653
R892 VPB.n1416 VPB.n1415 13.653
R893 VPB.n1424 VPB.n1423 13.653
R894 VPB.n1423 VPB.n1422 13.653
R895 VPB.n1429 VPB.n1428 13.653
R896 VPB.n1428 VPB.n1427 13.653
R897 VPB.n1434 VPB.n1433 13.653
R898 VPB.n1433 VPB.n1432 13.653
R899 VPB.n1441 VPB.n1440 13.653
R900 VPB.n1440 VPB.n1439 13.653
R901 VPB.n1446 VPB.n1445 13.653
R902 VPB.n1445 VPB.n1444 13.653
R903 VPB.n1451 VPB.n1450 13.653
R904 VPB.n1450 VPB.n1449 13.653
R905 VPB.n1455 VPB.n1454 13.653
R906 VPB.n1454 VPB.n1453 13.653
R907 VPB.n1459 VPB.n1458 13.653
R908 VPB.n1458 VPB.n1457 13.653
R909 VPB.n1486 VPB.n1485 13.653
R910 VPB.n1485 VPB.n1484 13.653
R911 VPB.n1490 VPB.n1489 13.653
R912 VPB.n1489 VPB.n1488 13.653
R913 VPB.n1495 VPB.n1494 13.653
R914 VPB.n1494 VPB.n1493 13.653
R915 VPB.n1500 VPB.n1499 13.653
R916 VPB.n1499 VPB.n1498 13.653
R917 VPB.n1507 VPB.n1506 13.653
R918 VPB.n1506 VPB.n1505 13.653
R919 VPB.n1512 VPB.n1511 13.653
R920 VPB.n1511 VPB.n1510 13.653
R921 VPB.n1517 VPB.n1516 13.653
R922 VPB.n1516 VPB.n1515 13.653
R923 VPB.n1524 VPB.n1523 13.653
R924 VPB.n1523 VPB.n1522 13.653
R925 VPB.n1529 VPB.n1528 13.653
R926 VPB.n1528 VPB.n1527 13.653
R927 VPB.n1534 VPB.n1533 13.653
R928 VPB.n1533 VPB.n1532 13.653
R929 VPB.n1538 VPB.n1537 13.653
R930 VPB.n1537 VPB.n1536 13.653
R931 VPB.n1542 VPB.n1541 13.653
R932 VPB.n1541 VPB.n1540 13.653
R933 VPB.n1569 VPB.n1568 13.653
R934 VPB.n1568 VPB.n1567 13.653
R935 VPB.n1573 VPB.n1572 13.653
R936 VPB.n1572 VPB.n1571 13.653
R937 VPB.n1578 VPB.n1577 13.653
R938 VPB.n1577 VPB.n1576 13.653
R939 VPB.n1583 VPB.n1582 13.653
R940 VPB.n1582 VPB.n1581 13.653
R941 VPB.n1590 VPB.n1589 13.653
R942 VPB.n1589 VPB.n1588 13.653
R943 VPB.n1595 VPB.n1594 13.653
R944 VPB.n1594 VPB.n1593 13.653
R945 VPB.n1600 VPB.n1599 13.653
R946 VPB.n1599 VPB.n1598 13.653
R947 VPB.n1607 VPB.n1606 13.653
R948 VPB.n1606 VPB.n1605 13.653
R949 VPB.n1612 VPB.n1611 13.653
R950 VPB.n1611 VPB.n1610 13.653
R951 VPB.n1617 VPB.n1616 13.653
R952 VPB.n1616 VPB.n1615 13.653
R953 VPB.n1621 VPB.n1620 13.653
R954 VPB.n1620 VPB.n1619 13.653
R955 VPB.n1625 VPB.n1624 13.653
R956 VPB.n1624 VPB.n1623 13.653
R957 VPB.n1652 VPB.n1651 13.653
R958 VPB.n1651 VPB.n1650 13.653
R959 VPB.n1656 VPB.n1655 13.653
R960 VPB.n1655 VPB.n1654 13.653
R961 VPB.n1661 VPB.n1660 13.653
R962 VPB.n1660 VPB.n1659 13.653
R963 VPB.n1666 VPB.n1665 13.653
R964 VPB.n1665 VPB.n1664 13.653
R965 VPB.n1673 VPB.n1672 13.653
R966 VPB.n1672 VPB.n1671 13.653
R967 VPB.n1678 VPB.n1677 13.653
R968 VPB.n1677 VPB.n1676 13.653
R969 VPB.n1683 VPB.n1682 13.653
R970 VPB.n1682 VPB.n1681 13.653
R971 VPB.n1690 VPB.n1689 13.653
R972 VPB.n1689 VPB.n1688 13.653
R973 VPB.n1695 VPB.n1694 13.653
R974 VPB.n1694 VPB.n1693 13.653
R975 VPB.n1700 VPB.n1699 13.653
R976 VPB.n1699 VPB.n1698 13.653
R977 VPB.n1704 VPB.n1703 13.653
R978 VPB.n1703 VPB.n1702 13.653
R979 VPB.n1708 VPB.n1707 13.653
R980 VPB.n1707 VPB.n1706 13.653
R981 VPB.n41 VPB.n40 13.653
R982 VPB.n40 VPB.n39 13.653
R983 VPB.n44 VPB.n43 13.653
R984 VPB.n43 VPB.n42 13.653
R985 VPB.n48 VPB.n47 13.653
R986 VPB.n47 VPB.n46 13.653
R987 VPB.n52 VPB.n51 13.653
R988 VPB.n51 VPB.n50 13.653
R989 VPB.n56 VPB.n55 13.653
R990 VPB.n55 VPB.n54 13.653
R991 VPB.n61 VPB.n60 13.653
R992 VPB.n60 VPB.n59 13.653
R993 VPB.n65 VPB.n64 13.653
R994 VPB.n64 VPB.n63 13.653
R995 VPB.n70 VPB.n69 13.653
R996 VPB.n69 VPB.n68 13.653
R997 VPB.n74 VPB.n73 13.653
R998 VPB.n73 VPB.n72 13.653
R999 VPB.n77 VPB.n76 13.653
R1000 VPB.n76 VPB.n75 13.653
R1001 VPB.n81 VPB.n80 13.653
R1002 VPB.n80 VPB.n79 13.653
R1003 VPB.n1722 VPB.n0 13.653
R1004 VPB VPB.n0 13.653
R1005 VPB.n344 VPB.n343 13.35
R1006 VPB.n416 VPB.n415 13.35
R1007 VPB.n499 VPB.n498 13.35
R1008 VPB.n582 VPB.n581 13.35
R1009 VPB.n665 VPB.n664 13.35
R1010 VPB.n748 VPB.n747 13.35
R1011 VPB.n831 VPB.n830 13.35
R1012 VPB.n914 VPB.n913 13.35
R1013 VPB.n137 VPB.n136 13.35
R1014 VPB.n1017 VPB.n1016 13.35
R1015 VPB.n1100 VPB.n1099 13.35
R1016 VPB.n1183 VPB.n1182 13.35
R1017 VPB.n1266 VPB.n1265 13.35
R1018 VPB.n1349 VPB.n1348 13.35
R1019 VPB.n1432 VPB.n1431 13.35
R1020 VPB.n1515 VPB.n1514 13.35
R1021 VPB.n1598 VPB.n1597 13.35
R1022 VPB.n1681 VPB.n1680 13.35
R1023 VPB.n63 VPB.n62 13.35
R1024 VPB.n1726 VPB.n1725 13.276
R1025 VPB.n1725 VPB.n1723 13.276
R1026 VPB.n36 VPB.n18 13.276
R1027 VPB.n18 VPB.n16 13.276
R1028 VPB.n1647 VPB.n1629 13.276
R1029 VPB.n1629 VPB.n1627 13.276
R1030 VPB.n1564 VPB.n1546 13.276
R1031 VPB.n1546 VPB.n1544 13.276
R1032 VPB.n1481 VPB.n1463 13.276
R1033 VPB.n1463 VPB.n1461 13.276
R1034 VPB.n1398 VPB.n1380 13.276
R1035 VPB.n1380 VPB.n1378 13.276
R1036 VPB.n1315 VPB.n1297 13.276
R1037 VPB.n1297 VPB.n1295 13.276
R1038 VPB.n1232 VPB.n1214 13.276
R1039 VPB.n1214 VPB.n1212 13.276
R1040 VPB.n1149 VPB.n1131 13.276
R1041 VPB.n1131 VPB.n1129 13.276
R1042 VPB.n1066 VPB.n1048 13.276
R1043 VPB.n1048 VPB.n1046 13.276
R1044 VPB.n983 VPB.n965 13.276
R1045 VPB.n965 VPB.n963 13.276
R1046 VPB.n104 VPB.n86 13.276
R1047 VPB.n86 VPB.n84 13.276
R1048 VPB.n880 VPB.n862 13.276
R1049 VPB.n862 VPB.n860 13.276
R1050 VPB.n797 VPB.n779 13.276
R1051 VPB.n779 VPB.n777 13.276
R1052 VPB.n714 VPB.n696 13.276
R1053 VPB.n696 VPB.n694 13.276
R1054 VPB.n631 VPB.n613 13.276
R1055 VPB.n613 VPB.n611 13.276
R1056 VPB.n548 VPB.n530 13.276
R1057 VPB.n530 VPB.n528 13.276
R1058 VPB.n465 VPB.n447 13.276
R1059 VPB.n447 VPB.n445 13.276
R1060 VPB.n382 VPB.n364 13.276
R1061 VPB.n364 VPB.n362 13.276
R1062 VPB.n319 VPB.n301 13.276
R1063 VPB.n301 VPB.n299 13.276
R1064 VPB.n264 VPB.n246 13.276
R1065 VPB.n246 VPB.n244 13.276
R1066 VPB.n209 VPB.n191 13.276
R1067 VPB.n191 VPB.n189 13.276
R1068 VPB.n214 VPB.n210 13.276
R1069 VPB.n269 VPB.n265 13.276
R1070 VPB.n324 VPB.n320 13.276
R1071 VPB.n387 VPB.n383 13.276
R1072 VPB.n470 VPB.n466 13.276
R1073 VPB.n553 VPB.n549 13.276
R1074 VPB.n636 VPB.n632 13.276
R1075 VPB.n719 VPB.n715 13.276
R1076 VPB.n802 VPB.n798 13.276
R1077 VPB.n885 VPB.n881 13.276
R1078 VPB.n110 VPB.n107 13.276
R1079 VPB.n111 VPB.n110 13.276
R1080 VPB.n115 VPB.n111 13.276
R1081 VPB.n118 VPB.n115 13.276
R1082 VPB.n126 VPB.n122 13.276
R1083 VPB.n130 VPB.n126 13.276
R1084 VPB.n139 VPB.n135 13.276
R1085 VPB.n949 VPB.n144 13.276
R1086 VPB.n953 VPB.n949 13.276
R1087 VPB.n988 VPB.n984 13.276
R1088 VPB.n1071 VPB.n1067 13.276
R1089 VPB.n1154 VPB.n1150 13.276
R1090 VPB.n1237 VPB.n1233 13.276
R1091 VPB.n1320 VPB.n1316 13.276
R1092 VPB.n1403 VPB.n1399 13.276
R1093 VPB.n1486 VPB.n1482 13.276
R1094 VPB.n1569 VPB.n1565 13.276
R1095 VPB.n1652 VPB.n1648 13.276
R1096 VPB.n41 VPB.n37 13.276
R1097 VPB.n44 VPB.n41 13.276
R1098 VPB.n52 VPB.n48 13.276
R1099 VPB.n56 VPB.n52 13.276
R1100 VPB.n65 VPB.n61 13.276
R1101 VPB.n74 VPB.n70 13.276
R1102 VPB.n77 VPB.n74 13.276
R1103 VPB.n1722 VPB.n81 13.276
R1104 VPB.n165 VPB.n147 13.276
R1105 VPB.n147 VPB.n145 13.276
R1106 VPB.n152 VPB.n150 12.796
R1107 VPB.n152 VPB.n151 12.564
R1108 VPB.n81 VPB.n78 12.558
R1109 VPB.n119 VPB.n118 12.2
R1110 VPB.n45 VPB.n44 12.2
R1111 VPB.n161 VPB.n160 12.198
R1112 VPB.n158 VPB.n157 12.198
R1113 VPB.n158 VPB.n155 12.198
R1114 VPB.n135 VPB.n131 9.329
R1115 VPB.n61 VPB.n57 9.329
R1116 VPB.n140 VPB.n139 8.97
R1117 VPB.n66 VPB.n65 8.97
R1118 VPB.n165 VPB.n164 7.5
R1119 VPB.n150 VPB.n149 7.5
R1120 VPB.n157 VPB.n156 7.5
R1121 VPB.n155 VPB.n154 7.5
R1122 VPB.n147 VPB.n146 7.5
R1123 VPB.n162 VPB.n148 7.5
R1124 VPB.n191 VPB.n190 7.5
R1125 VPB.n204 VPB.n203 7.5
R1126 VPB.n198 VPB.n197 7.5
R1127 VPB.n200 VPB.n199 7.5
R1128 VPB.n193 VPB.n192 7.5
R1129 VPB.n209 VPB.n208 7.5
R1130 VPB.n246 VPB.n245 7.5
R1131 VPB.n259 VPB.n258 7.5
R1132 VPB.n253 VPB.n252 7.5
R1133 VPB.n255 VPB.n254 7.5
R1134 VPB.n248 VPB.n247 7.5
R1135 VPB.n264 VPB.n263 7.5
R1136 VPB.n301 VPB.n300 7.5
R1137 VPB.n314 VPB.n313 7.5
R1138 VPB.n308 VPB.n307 7.5
R1139 VPB.n310 VPB.n309 7.5
R1140 VPB.n303 VPB.n302 7.5
R1141 VPB.n319 VPB.n318 7.5
R1142 VPB.n364 VPB.n363 7.5
R1143 VPB.n377 VPB.n376 7.5
R1144 VPB.n371 VPB.n370 7.5
R1145 VPB.n373 VPB.n372 7.5
R1146 VPB.n366 VPB.n365 7.5
R1147 VPB.n382 VPB.n381 7.5
R1148 VPB.n447 VPB.n446 7.5
R1149 VPB.n460 VPB.n459 7.5
R1150 VPB.n454 VPB.n453 7.5
R1151 VPB.n456 VPB.n455 7.5
R1152 VPB.n449 VPB.n448 7.5
R1153 VPB.n465 VPB.n464 7.5
R1154 VPB.n530 VPB.n529 7.5
R1155 VPB.n543 VPB.n542 7.5
R1156 VPB.n537 VPB.n536 7.5
R1157 VPB.n539 VPB.n538 7.5
R1158 VPB.n532 VPB.n531 7.5
R1159 VPB.n548 VPB.n547 7.5
R1160 VPB.n613 VPB.n612 7.5
R1161 VPB.n626 VPB.n625 7.5
R1162 VPB.n620 VPB.n619 7.5
R1163 VPB.n622 VPB.n621 7.5
R1164 VPB.n615 VPB.n614 7.5
R1165 VPB.n631 VPB.n630 7.5
R1166 VPB.n696 VPB.n695 7.5
R1167 VPB.n709 VPB.n708 7.5
R1168 VPB.n703 VPB.n702 7.5
R1169 VPB.n705 VPB.n704 7.5
R1170 VPB.n698 VPB.n697 7.5
R1171 VPB.n714 VPB.n713 7.5
R1172 VPB.n779 VPB.n778 7.5
R1173 VPB.n792 VPB.n791 7.5
R1174 VPB.n786 VPB.n785 7.5
R1175 VPB.n788 VPB.n787 7.5
R1176 VPB.n781 VPB.n780 7.5
R1177 VPB.n797 VPB.n796 7.5
R1178 VPB.n862 VPB.n861 7.5
R1179 VPB.n875 VPB.n874 7.5
R1180 VPB.n869 VPB.n868 7.5
R1181 VPB.n871 VPB.n870 7.5
R1182 VPB.n864 VPB.n863 7.5
R1183 VPB.n880 VPB.n879 7.5
R1184 VPB.n86 VPB.n85 7.5
R1185 VPB.n99 VPB.n98 7.5
R1186 VPB.n93 VPB.n92 7.5
R1187 VPB.n95 VPB.n94 7.5
R1188 VPB.n88 VPB.n87 7.5
R1189 VPB.n104 VPB.n103 7.5
R1190 VPB.n965 VPB.n964 7.5
R1191 VPB.n978 VPB.n977 7.5
R1192 VPB.n972 VPB.n971 7.5
R1193 VPB.n974 VPB.n973 7.5
R1194 VPB.n967 VPB.n966 7.5
R1195 VPB.n983 VPB.n982 7.5
R1196 VPB.n1048 VPB.n1047 7.5
R1197 VPB.n1061 VPB.n1060 7.5
R1198 VPB.n1055 VPB.n1054 7.5
R1199 VPB.n1057 VPB.n1056 7.5
R1200 VPB.n1050 VPB.n1049 7.5
R1201 VPB.n1066 VPB.n1065 7.5
R1202 VPB.n1131 VPB.n1130 7.5
R1203 VPB.n1144 VPB.n1143 7.5
R1204 VPB.n1138 VPB.n1137 7.5
R1205 VPB.n1140 VPB.n1139 7.5
R1206 VPB.n1133 VPB.n1132 7.5
R1207 VPB.n1149 VPB.n1148 7.5
R1208 VPB.n1214 VPB.n1213 7.5
R1209 VPB.n1227 VPB.n1226 7.5
R1210 VPB.n1221 VPB.n1220 7.5
R1211 VPB.n1223 VPB.n1222 7.5
R1212 VPB.n1216 VPB.n1215 7.5
R1213 VPB.n1232 VPB.n1231 7.5
R1214 VPB.n1297 VPB.n1296 7.5
R1215 VPB.n1310 VPB.n1309 7.5
R1216 VPB.n1304 VPB.n1303 7.5
R1217 VPB.n1306 VPB.n1305 7.5
R1218 VPB.n1299 VPB.n1298 7.5
R1219 VPB.n1315 VPB.n1314 7.5
R1220 VPB.n1380 VPB.n1379 7.5
R1221 VPB.n1393 VPB.n1392 7.5
R1222 VPB.n1387 VPB.n1386 7.5
R1223 VPB.n1389 VPB.n1388 7.5
R1224 VPB.n1382 VPB.n1381 7.5
R1225 VPB.n1398 VPB.n1397 7.5
R1226 VPB.n1463 VPB.n1462 7.5
R1227 VPB.n1476 VPB.n1475 7.5
R1228 VPB.n1470 VPB.n1469 7.5
R1229 VPB.n1472 VPB.n1471 7.5
R1230 VPB.n1465 VPB.n1464 7.5
R1231 VPB.n1481 VPB.n1480 7.5
R1232 VPB.n1546 VPB.n1545 7.5
R1233 VPB.n1559 VPB.n1558 7.5
R1234 VPB.n1553 VPB.n1552 7.5
R1235 VPB.n1555 VPB.n1554 7.5
R1236 VPB.n1548 VPB.n1547 7.5
R1237 VPB.n1564 VPB.n1563 7.5
R1238 VPB.n1629 VPB.n1628 7.5
R1239 VPB.n1642 VPB.n1641 7.5
R1240 VPB.n1636 VPB.n1635 7.5
R1241 VPB.n1638 VPB.n1637 7.5
R1242 VPB.n1631 VPB.n1630 7.5
R1243 VPB.n1647 VPB.n1646 7.5
R1244 VPB.n18 VPB.n17 7.5
R1245 VPB.n31 VPB.n30 7.5
R1246 VPB.n25 VPB.n24 7.5
R1247 VPB.n27 VPB.n26 7.5
R1248 VPB.n20 VPB.n19 7.5
R1249 VPB.n36 VPB.n35 7.5
R1250 VPB.n1725 VPB.n1724 7.5
R1251 VPB.n12 VPB.n11 7.5
R1252 VPB.n6 VPB.n5 7.5
R1253 VPB.n8 VPB.n7 7.5
R1254 VPB.n2 VPB.n1 7.5
R1255 VPB.n1727 VPB.n1726 7.5
R1256 VPB.n37 VPB.n36 7.176
R1257 VPB.n1648 VPB.n1647 7.176
R1258 VPB.n1565 VPB.n1564 7.176
R1259 VPB.n1482 VPB.n1481 7.176
R1260 VPB.n1399 VPB.n1398 7.176
R1261 VPB.n1316 VPB.n1315 7.176
R1262 VPB.n1233 VPB.n1232 7.176
R1263 VPB.n1150 VPB.n1149 7.176
R1264 VPB.n1067 VPB.n1066 7.176
R1265 VPB.n984 VPB.n983 7.176
R1266 VPB.n111 VPB.n104 7.176
R1267 VPB.n881 VPB.n880 7.176
R1268 VPB.n798 VPB.n797 7.176
R1269 VPB.n715 VPB.n714 7.176
R1270 VPB.n632 VPB.n631 7.176
R1271 VPB.n549 VPB.n548 7.176
R1272 VPB.n466 VPB.n465 7.176
R1273 VPB.n383 VPB.n382 7.176
R1274 VPB.n320 VPB.n319 7.176
R1275 VPB.n265 VPB.n264 7.176
R1276 VPB.n210 VPB.n209 7.176
R1277 VPB.n205 VPB.n202 6.729
R1278 VPB.n201 VPB.n198 6.729
R1279 VPB.n196 VPB.n193 6.729
R1280 VPB.n260 VPB.n257 6.729
R1281 VPB.n256 VPB.n253 6.729
R1282 VPB.n251 VPB.n248 6.729
R1283 VPB.n315 VPB.n312 6.729
R1284 VPB.n311 VPB.n308 6.729
R1285 VPB.n306 VPB.n303 6.729
R1286 VPB.n378 VPB.n375 6.729
R1287 VPB.n374 VPB.n371 6.729
R1288 VPB.n369 VPB.n366 6.729
R1289 VPB.n461 VPB.n458 6.729
R1290 VPB.n457 VPB.n454 6.729
R1291 VPB.n452 VPB.n449 6.729
R1292 VPB.n544 VPB.n541 6.729
R1293 VPB.n540 VPB.n537 6.729
R1294 VPB.n535 VPB.n532 6.729
R1295 VPB.n627 VPB.n624 6.729
R1296 VPB.n623 VPB.n620 6.729
R1297 VPB.n618 VPB.n615 6.729
R1298 VPB.n710 VPB.n707 6.729
R1299 VPB.n706 VPB.n703 6.729
R1300 VPB.n701 VPB.n698 6.729
R1301 VPB.n793 VPB.n790 6.729
R1302 VPB.n789 VPB.n786 6.729
R1303 VPB.n784 VPB.n781 6.729
R1304 VPB.n876 VPB.n873 6.729
R1305 VPB.n872 VPB.n869 6.729
R1306 VPB.n867 VPB.n864 6.729
R1307 VPB.n100 VPB.n97 6.729
R1308 VPB.n96 VPB.n93 6.729
R1309 VPB.n91 VPB.n88 6.729
R1310 VPB.n979 VPB.n976 6.729
R1311 VPB.n975 VPB.n972 6.729
R1312 VPB.n970 VPB.n967 6.729
R1313 VPB.n1062 VPB.n1059 6.729
R1314 VPB.n1058 VPB.n1055 6.729
R1315 VPB.n1053 VPB.n1050 6.729
R1316 VPB.n1145 VPB.n1142 6.729
R1317 VPB.n1141 VPB.n1138 6.729
R1318 VPB.n1136 VPB.n1133 6.729
R1319 VPB.n1228 VPB.n1225 6.729
R1320 VPB.n1224 VPB.n1221 6.729
R1321 VPB.n1219 VPB.n1216 6.729
R1322 VPB.n1311 VPB.n1308 6.729
R1323 VPB.n1307 VPB.n1304 6.729
R1324 VPB.n1302 VPB.n1299 6.729
R1325 VPB.n1394 VPB.n1391 6.729
R1326 VPB.n1390 VPB.n1387 6.729
R1327 VPB.n1385 VPB.n1382 6.729
R1328 VPB.n1477 VPB.n1474 6.729
R1329 VPB.n1473 VPB.n1470 6.729
R1330 VPB.n1468 VPB.n1465 6.729
R1331 VPB.n1560 VPB.n1557 6.729
R1332 VPB.n1556 VPB.n1553 6.729
R1333 VPB.n1551 VPB.n1548 6.729
R1334 VPB.n1643 VPB.n1640 6.729
R1335 VPB.n1639 VPB.n1636 6.729
R1336 VPB.n1634 VPB.n1631 6.729
R1337 VPB.n32 VPB.n29 6.729
R1338 VPB.n28 VPB.n25 6.729
R1339 VPB.n23 VPB.n20 6.729
R1340 VPB.n13 VPB.n10 6.729
R1341 VPB.n9 VPB.n6 6.729
R1342 VPB.n4 VPB.n2 6.729
R1343 VPB.n196 VPB.n195 6.728
R1344 VPB.n201 VPB.n200 6.728
R1345 VPB.n205 VPB.n204 6.728
R1346 VPB.n208 VPB.n207 6.728
R1347 VPB.n251 VPB.n250 6.728
R1348 VPB.n256 VPB.n255 6.728
R1349 VPB.n260 VPB.n259 6.728
R1350 VPB.n263 VPB.n262 6.728
R1351 VPB.n306 VPB.n305 6.728
R1352 VPB.n311 VPB.n310 6.728
R1353 VPB.n315 VPB.n314 6.728
R1354 VPB.n318 VPB.n317 6.728
R1355 VPB.n369 VPB.n368 6.728
R1356 VPB.n374 VPB.n373 6.728
R1357 VPB.n378 VPB.n377 6.728
R1358 VPB.n381 VPB.n380 6.728
R1359 VPB.n452 VPB.n451 6.728
R1360 VPB.n457 VPB.n456 6.728
R1361 VPB.n461 VPB.n460 6.728
R1362 VPB.n464 VPB.n463 6.728
R1363 VPB.n535 VPB.n534 6.728
R1364 VPB.n540 VPB.n539 6.728
R1365 VPB.n544 VPB.n543 6.728
R1366 VPB.n547 VPB.n546 6.728
R1367 VPB.n618 VPB.n617 6.728
R1368 VPB.n623 VPB.n622 6.728
R1369 VPB.n627 VPB.n626 6.728
R1370 VPB.n630 VPB.n629 6.728
R1371 VPB.n701 VPB.n700 6.728
R1372 VPB.n706 VPB.n705 6.728
R1373 VPB.n710 VPB.n709 6.728
R1374 VPB.n713 VPB.n712 6.728
R1375 VPB.n784 VPB.n783 6.728
R1376 VPB.n789 VPB.n788 6.728
R1377 VPB.n793 VPB.n792 6.728
R1378 VPB.n796 VPB.n795 6.728
R1379 VPB.n867 VPB.n866 6.728
R1380 VPB.n872 VPB.n871 6.728
R1381 VPB.n876 VPB.n875 6.728
R1382 VPB.n879 VPB.n878 6.728
R1383 VPB.n91 VPB.n90 6.728
R1384 VPB.n96 VPB.n95 6.728
R1385 VPB.n100 VPB.n99 6.728
R1386 VPB.n103 VPB.n102 6.728
R1387 VPB.n970 VPB.n969 6.728
R1388 VPB.n975 VPB.n974 6.728
R1389 VPB.n979 VPB.n978 6.728
R1390 VPB.n982 VPB.n981 6.728
R1391 VPB.n1053 VPB.n1052 6.728
R1392 VPB.n1058 VPB.n1057 6.728
R1393 VPB.n1062 VPB.n1061 6.728
R1394 VPB.n1065 VPB.n1064 6.728
R1395 VPB.n1136 VPB.n1135 6.728
R1396 VPB.n1141 VPB.n1140 6.728
R1397 VPB.n1145 VPB.n1144 6.728
R1398 VPB.n1148 VPB.n1147 6.728
R1399 VPB.n1219 VPB.n1218 6.728
R1400 VPB.n1224 VPB.n1223 6.728
R1401 VPB.n1228 VPB.n1227 6.728
R1402 VPB.n1231 VPB.n1230 6.728
R1403 VPB.n1302 VPB.n1301 6.728
R1404 VPB.n1307 VPB.n1306 6.728
R1405 VPB.n1311 VPB.n1310 6.728
R1406 VPB.n1314 VPB.n1313 6.728
R1407 VPB.n1385 VPB.n1384 6.728
R1408 VPB.n1390 VPB.n1389 6.728
R1409 VPB.n1394 VPB.n1393 6.728
R1410 VPB.n1397 VPB.n1396 6.728
R1411 VPB.n1468 VPB.n1467 6.728
R1412 VPB.n1473 VPB.n1472 6.728
R1413 VPB.n1477 VPB.n1476 6.728
R1414 VPB.n1480 VPB.n1479 6.728
R1415 VPB.n1551 VPB.n1550 6.728
R1416 VPB.n1556 VPB.n1555 6.728
R1417 VPB.n1560 VPB.n1559 6.728
R1418 VPB.n1563 VPB.n1562 6.728
R1419 VPB.n1634 VPB.n1633 6.728
R1420 VPB.n1639 VPB.n1638 6.728
R1421 VPB.n1643 VPB.n1642 6.728
R1422 VPB.n1646 VPB.n1645 6.728
R1423 VPB.n23 VPB.n22 6.728
R1424 VPB.n28 VPB.n27 6.728
R1425 VPB.n32 VPB.n31 6.728
R1426 VPB.n35 VPB.n34 6.728
R1427 VPB.n4 VPB.n3 6.728
R1428 VPB.n9 VPB.n8 6.728
R1429 VPB.n13 VPB.n12 6.728
R1430 VPB.n1728 VPB.n1727 6.728
R1431 VPB.n341 VPB.n337 6.458
R1432 VPB.n164 VPB.n163 6.398
R1433 VPB.n425 VPB.n421 4.305
R1434 VPB.n508 VPB.n504 4.305
R1435 VPB.n591 VPB.n587 4.305
R1436 VPB.n674 VPB.n670 4.305
R1437 VPB.n757 VPB.n753 4.305
R1438 VPB.n840 VPB.n836 4.305
R1439 VPB.n923 VPB.n919 4.305
R1440 VPB.n144 VPB.n140 4.305
R1441 VPB.n1026 VPB.n1022 4.305
R1442 VPB.n1109 VPB.n1105 4.305
R1443 VPB.n1192 VPB.n1188 4.305
R1444 VPB.n1275 VPB.n1271 4.305
R1445 VPB.n1358 VPB.n1354 4.305
R1446 VPB.n1441 VPB.n1437 4.305
R1447 VPB.n1524 VPB.n1520 4.305
R1448 VPB.n1607 VPB.n1603 4.305
R1449 VPB.n1690 VPB.n1686 4.305
R1450 VPB.n70 VPB.n66 4.305
R1451 VPB.n408 VPB.n404 3.947
R1452 VPB.n491 VPB.n487 3.947
R1453 VPB.n574 VPB.n570 3.947
R1454 VPB.n657 VPB.n653 3.947
R1455 VPB.n740 VPB.n736 3.947
R1456 VPB.n823 VPB.n819 3.947
R1457 VPB.n906 VPB.n902 3.947
R1458 VPB.n131 VPB.n130 3.947
R1459 VPB.n1009 VPB.n1005 3.947
R1460 VPB.n1092 VPB.n1088 3.947
R1461 VPB.n1175 VPB.n1171 3.947
R1462 VPB.n1258 VPB.n1254 3.947
R1463 VPB.n1341 VPB.n1337 3.947
R1464 VPB.n1424 VPB.n1420 3.947
R1465 VPB.n1507 VPB.n1503 3.947
R1466 VPB.n1590 VPB.n1586 3.947
R1467 VPB.n1673 VPB.n1669 3.947
R1468 VPB.n57 VPB.n56 3.947
R1469 VPB.n173 VPB.n169 2.691
R1470 VPB.n183 VPB.n179 2.332
R1471 VPB.n356 VPB.n353 1.794
R1472 VPB.n329 VPB.n326 1.435
R1473 VPB.n162 VPB.n153 1.402
R1474 VPB.n162 VPB.n158 1.402
R1475 VPB.n162 VPB.n159 1.402
R1476 VPB.n162 VPB.n161 1.402
R1477 VPB.n396 VPB.n393 1.076
R1478 VPB.n479 VPB.n476 1.076
R1479 VPB.n562 VPB.n559 1.076
R1480 VPB.n645 VPB.n642 1.076
R1481 VPB.n728 VPB.n725 1.076
R1482 VPB.n811 VPB.n808 1.076
R1483 VPB.n894 VPB.n891 1.076
R1484 VPB.n122 VPB.n119 1.076
R1485 VPB.n997 VPB.n994 1.076
R1486 VPB.n1080 VPB.n1077 1.076
R1487 VPB.n1163 VPB.n1160 1.076
R1488 VPB.n1246 VPB.n1243 1.076
R1489 VPB.n1329 VPB.n1326 1.076
R1490 VPB.n1412 VPB.n1409 1.076
R1491 VPB.n1495 VPB.n1492 1.076
R1492 VPB.n1578 VPB.n1575 1.076
R1493 VPB.n1661 VPB.n1658 1.076
R1494 VPB.n48 VPB.n45 1.076
R1495 VPB.n163 VPB.n162 0.735
R1496 VPB.n162 VPB.n152 0.735
R1497 VPB.n435 VPB.n432 0.717
R1498 VPB.n518 VPB.n515 0.717
R1499 VPB.n601 VPB.n598 0.717
R1500 VPB.n684 VPB.n681 0.717
R1501 VPB.n767 VPB.n764 0.717
R1502 VPB.n850 VPB.n847 0.717
R1503 VPB.n933 VPB.n930 0.717
R1504 VPB.n953 VPB.n950 0.717
R1505 VPB.n1036 VPB.n1033 0.717
R1506 VPB.n1119 VPB.n1116 0.717
R1507 VPB.n1202 VPB.n1199 0.717
R1508 VPB.n1285 VPB.n1282 0.717
R1509 VPB.n1368 VPB.n1365 0.717
R1510 VPB.n1451 VPB.n1448 0.717
R1511 VPB.n1534 VPB.n1531 0.717
R1512 VPB.n1617 VPB.n1614 0.717
R1513 VPB.n1700 VPB.n1697 0.717
R1514 VPB.n78 VPB.n77 0.717
R1515 VPB.n206 VPB.n205 0.387
R1516 VPB.n206 VPB.n201 0.387
R1517 VPB.n206 VPB.n196 0.387
R1518 VPB.n207 VPB.n206 0.387
R1519 VPB.n261 VPB.n260 0.387
R1520 VPB.n261 VPB.n256 0.387
R1521 VPB.n261 VPB.n251 0.387
R1522 VPB.n262 VPB.n261 0.387
R1523 VPB.n316 VPB.n315 0.387
R1524 VPB.n316 VPB.n311 0.387
R1525 VPB.n316 VPB.n306 0.387
R1526 VPB.n317 VPB.n316 0.387
R1527 VPB.n379 VPB.n378 0.387
R1528 VPB.n379 VPB.n374 0.387
R1529 VPB.n379 VPB.n369 0.387
R1530 VPB.n380 VPB.n379 0.387
R1531 VPB.n462 VPB.n461 0.387
R1532 VPB.n462 VPB.n457 0.387
R1533 VPB.n462 VPB.n452 0.387
R1534 VPB.n463 VPB.n462 0.387
R1535 VPB.n545 VPB.n544 0.387
R1536 VPB.n545 VPB.n540 0.387
R1537 VPB.n545 VPB.n535 0.387
R1538 VPB.n546 VPB.n545 0.387
R1539 VPB.n628 VPB.n627 0.387
R1540 VPB.n628 VPB.n623 0.387
R1541 VPB.n628 VPB.n618 0.387
R1542 VPB.n629 VPB.n628 0.387
R1543 VPB.n711 VPB.n710 0.387
R1544 VPB.n711 VPB.n706 0.387
R1545 VPB.n711 VPB.n701 0.387
R1546 VPB.n712 VPB.n711 0.387
R1547 VPB.n794 VPB.n793 0.387
R1548 VPB.n794 VPB.n789 0.387
R1549 VPB.n794 VPB.n784 0.387
R1550 VPB.n795 VPB.n794 0.387
R1551 VPB.n877 VPB.n876 0.387
R1552 VPB.n877 VPB.n872 0.387
R1553 VPB.n877 VPB.n867 0.387
R1554 VPB.n878 VPB.n877 0.387
R1555 VPB.n101 VPB.n100 0.387
R1556 VPB.n101 VPB.n96 0.387
R1557 VPB.n101 VPB.n91 0.387
R1558 VPB.n102 VPB.n101 0.387
R1559 VPB.n980 VPB.n979 0.387
R1560 VPB.n980 VPB.n975 0.387
R1561 VPB.n980 VPB.n970 0.387
R1562 VPB.n981 VPB.n980 0.387
R1563 VPB.n1063 VPB.n1062 0.387
R1564 VPB.n1063 VPB.n1058 0.387
R1565 VPB.n1063 VPB.n1053 0.387
R1566 VPB.n1064 VPB.n1063 0.387
R1567 VPB.n1146 VPB.n1145 0.387
R1568 VPB.n1146 VPB.n1141 0.387
R1569 VPB.n1146 VPB.n1136 0.387
R1570 VPB.n1147 VPB.n1146 0.387
R1571 VPB.n1229 VPB.n1228 0.387
R1572 VPB.n1229 VPB.n1224 0.387
R1573 VPB.n1229 VPB.n1219 0.387
R1574 VPB.n1230 VPB.n1229 0.387
R1575 VPB.n1312 VPB.n1311 0.387
R1576 VPB.n1312 VPB.n1307 0.387
R1577 VPB.n1312 VPB.n1302 0.387
R1578 VPB.n1313 VPB.n1312 0.387
R1579 VPB.n1395 VPB.n1394 0.387
R1580 VPB.n1395 VPB.n1390 0.387
R1581 VPB.n1395 VPB.n1385 0.387
R1582 VPB.n1396 VPB.n1395 0.387
R1583 VPB.n1478 VPB.n1477 0.387
R1584 VPB.n1478 VPB.n1473 0.387
R1585 VPB.n1478 VPB.n1468 0.387
R1586 VPB.n1479 VPB.n1478 0.387
R1587 VPB.n1561 VPB.n1560 0.387
R1588 VPB.n1561 VPB.n1556 0.387
R1589 VPB.n1561 VPB.n1551 0.387
R1590 VPB.n1562 VPB.n1561 0.387
R1591 VPB.n1644 VPB.n1643 0.387
R1592 VPB.n1644 VPB.n1639 0.387
R1593 VPB.n1644 VPB.n1634 0.387
R1594 VPB.n1645 VPB.n1644 0.387
R1595 VPB.n33 VPB.n32 0.387
R1596 VPB.n33 VPB.n28 0.387
R1597 VPB.n33 VPB.n23 0.387
R1598 VPB.n34 VPB.n33 0.387
R1599 VPB.n1729 VPB.n13 0.387
R1600 VPB.n1729 VPB.n9 0.387
R1601 VPB.n1729 VPB.n4 0.387
R1602 VPB.n1729 VPB.n1728 0.387
R1603 VPB.n215 VPB.n188 0.272
R1604 VPB.n270 VPB.n243 0.272
R1605 VPB.n325 VPB.n298 0.272
R1606 VPB.n388 VPB.n361 0.272
R1607 VPB.n471 VPB.n444 0.272
R1608 VPB.n554 VPB.n527 0.272
R1609 VPB.n637 VPB.n610 0.272
R1610 VPB.n720 VPB.n693 0.272
R1611 VPB.n803 VPB.n776 0.272
R1612 VPB.n886 VPB.n859 0.272
R1613 VPB.n937 VPB.n936 0.272
R1614 VPB.n989 VPB.n962 0.272
R1615 VPB.n1072 VPB.n1045 0.272
R1616 VPB.n1155 VPB.n1128 0.272
R1617 VPB.n1238 VPB.n1211 0.272
R1618 VPB.n1321 VPB.n1294 0.272
R1619 VPB.n1404 VPB.n1377 0.272
R1620 VPB.n1487 VPB.n1460 0.272
R1621 VPB.n1570 VPB.n1543 0.272
R1622 VPB.n1653 VPB.n1626 0.272
R1623 VPB.n1710 VPB.n1709 0.272
R1624 VPB.n1721 VPB 0.198
R1625 VPB.n178 VPB.n174 0.136
R1626 VPB.n184 VPB.n178 0.136
R1627 VPB.n188 VPB.n184 0.136
R1628 VPB.n219 VPB.n215 0.136
R1629 VPB.n223 VPB.n219 0.136
R1630 VPB.n227 VPB.n223 0.136
R1631 VPB.n231 VPB.n227 0.136
R1632 VPB.n235 VPB.n231 0.136
R1633 VPB.n239 VPB.n235 0.136
R1634 VPB.n243 VPB.n239 0.136
R1635 VPB.n274 VPB.n270 0.136
R1636 VPB.n278 VPB.n274 0.136
R1637 VPB.n282 VPB.n278 0.136
R1638 VPB.n286 VPB.n282 0.136
R1639 VPB.n290 VPB.n286 0.136
R1640 VPB.n294 VPB.n290 0.136
R1641 VPB.n298 VPB.n294 0.136
R1642 VPB.n330 VPB.n325 0.136
R1643 VPB.n335 VPB.n330 0.136
R1644 VPB.n342 VPB.n335 0.136
R1645 VPB.n347 VPB.n342 0.136
R1646 VPB.n352 VPB.n347 0.136
R1647 VPB.n357 VPB.n352 0.136
R1648 VPB.n361 VPB.n357 0.136
R1649 VPB.n392 VPB.n388 0.136
R1650 VPB.n397 VPB.n392 0.136
R1651 VPB.n402 VPB.n397 0.136
R1652 VPB.n409 VPB.n402 0.136
R1653 VPB.n414 VPB.n409 0.136
R1654 VPB.n419 VPB.n414 0.136
R1655 VPB.n426 VPB.n419 0.136
R1656 VPB.n431 VPB.n426 0.136
R1657 VPB.n436 VPB.n431 0.136
R1658 VPB.n440 VPB.n436 0.136
R1659 VPB.n444 VPB.n440 0.136
R1660 VPB.n475 VPB.n471 0.136
R1661 VPB.n480 VPB.n475 0.136
R1662 VPB.n485 VPB.n480 0.136
R1663 VPB.n492 VPB.n485 0.136
R1664 VPB.n497 VPB.n492 0.136
R1665 VPB.n502 VPB.n497 0.136
R1666 VPB.n509 VPB.n502 0.136
R1667 VPB.n514 VPB.n509 0.136
R1668 VPB.n519 VPB.n514 0.136
R1669 VPB.n523 VPB.n519 0.136
R1670 VPB.n527 VPB.n523 0.136
R1671 VPB.n558 VPB.n554 0.136
R1672 VPB.n563 VPB.n558 0.136
R1673 VPB.n568 VPB.n563 0.136
R1674 VPB.n575 VPB.n568 0.136
R1675 VPB.n580 VPB.n575 0.136
R1676 VPB.n585 VPB.n580 0.136
R1677 VPB.n592 VPB.n585 0.136
R1678 VPB.n597 VPB.n592 0.136
R1679 VPB.n602 VPB.n597 0.136
R1680 VPB.n606 VPB.n602 0.136
R1681 VPB.n610 VPB.n606 0.136
R1682 VPB.n641 VPB.n637 0.136
R1683 VPB.n646 VPB.n641 0.136
R1684 VPB.n651 VPB.n646 0.136
R1685 VPB.n658 VPB.n651 0.136
R1686 VPB.n663 VPB.n658 0.136
R1687 VPB.n668 VPB.n663 0.136
R1688 VPB.n675 VPB.n668 0.136
R1689 VPB.n680 VPB.n675 0.136
R1690 VPB.n685 VPB.n680 0.136
R1691 VPB.n689 VPB.n685 0.136
R1692 VPB.n693 VPB.n689 0.136
R1693 VPB.n724 VPB.n720 0.136
R1694 VPB.n729 VPB.n724 0.136
R1695 VPB.n734 VPB.n729 0.136
R1696 VPB.n741 VPB.n734 0.136
R1697 VPB.n746 VPB.n741 0.136
R1698 VPB.n751 VPB.n746 0.136
R1699 VPB.n758 VPB.n751 0.136
R1700 VPB.n763 VPB.n758 0.136
R1701 VPB.n768 VPB.n763 0.136
R1702 VPB.n772 VPB.n768 0.136
R1703 VPB.n776 VPB.n772 0.136
R1704 VPB.n807 VPB.n803 0.136
R1705 VPB.n812 VPB.n807 0.136
R1706 VPB.n817 VPB.n812 0.136
R1707 VPB.n824 VPB.n817 0.136
R1708 VPB.n829 VPB.n824 0.136
R1709 VPB.n834 VPB.n829 0.136
R1710 VPB.n841 VPB.n834 0.136
R1711 VPB.n846 VPB.n841 0.136
R1712 VPB.n851 VPB.n846 0.136
R1713 VPB.n855 VPB.n851 0.136
R1714 VPB.n859 VPB.n855 0.136
R1715 VPB.n890 VPB.n886 0.136
R1716 VPB.n895 VPB.n890 0.136
R1717 VPB.n900 VPB.n895 0.136
R1718 VPB.n907 VPB.n900 0.136
R1719 VPB.n912 VPB.n907 0.136
R1720 VPB.n917 VPB.n912 0.136
R1721 VPB.n924 VPB.n917 0.136
R1722 VPB.n929 VPB.n924 0.136
R1723 VPB.n934 VPB.n929 0.136
R1724 VPB.n935 VPB.n934 0.136
R1725 VPB.n936 VPB.n935 0.136
R1726 VPB.n938 VPB.n937 0.136
R1727 VPB.n939 VPB.n938 0.136
R1728 VPB.n940 VPB.n939 0.136
R1729 VPB.n941 VPB.n940 0.136
R1730 VPB.n942 VPB.n941 0.136
R1731 VPB.n943 VPB.n942 0.136
R1732 VPB.n944 VPB.n943 0.136
R1733 VPB.n945 VPB.n944 0.136
R1734 VPB.n958 VPB.n954 0.136
R1735 VPB.n962 VPB.n958 0.136
R1736 VPB.n993 VPB.n989 0.136
R1737 VPB.n998 VPB.n993 0.136
R1738 VPB.n1003 VPB.n998 0.136
R1739 VPB.n1010 VPB.n1003 0.136
R1740 VPB.n1015 VPB.n1010 0.136
R1741 VPB.n1020 VPB.n1015 0.136
R1742 VPB.n1027 VPB.n1020 0.136
R1743 VPB.n1032 VPB.n1027 0.136
R1744 VPB.n1037 VPB.n1032 0.136
R1745 VPB.n1041 VPB.n1037 0.136
R1746 VPB.n1045 VPB.n1041 0.136
R1747 VPB.n1076 VPB.n1072 0.136
R1748 VPB.n1081 VPB.n1076 0.136
R1749 VPB.n1086 VPB.n1081 0.136
R1750 VPB.n1093 VPB.n1086 0.136
R1751 VPB.n1098 VPB.n1093 0.136
R1752 VPB.n1103 VPB.n1098 0.136
R1753 VPB.n1110 VPB.n1103 0.136
R1754 VPB.n1115 VPB.n1110 0.136
R1755 VPB.n1120 VPB.n1115 0.136
R1756 VPB.n1124 VPB.n1120 0.136
R1757 VPB.n1128 VPB.n1124 0.136
R1758 VPB.n1159 VPB.n1155 0.136
R1759 VPB.n1164 VPB.n1159 0.136
R1760 VPB.n1169 VPB.n1164 0.136
R1761 VPB.n1176 VPB.n1169 0.136
R1762 VPB.n1181 VPB.n1176 0.136
R1763 VPB.n1186 VPB.n1181 0.136
R1764 VPB.n1193 VPB.n1186 0.136
R1765 VPB.n1198 VPB.n1193 0.136
R1766 VPB.n1203 VPB.n1198 0.136
R1767 VPB.n1207 VPB.n1203 0.136
R1768 VPB.n1211 VPB.n1207 0.136
R1769 VPB.n1242 VPB.n1238 0.136
R1770 VPB.n1247 VPB.n1242 0.136
R1771 VPB.n1252 VPB.n1247 0.136
R1772 VPB.n1259 VPB.n1252 0.136
R1773 VPB.n1264 VPB.n1259 0.136
R1774 VPB.n1269 VPB.n1264 0.136
R1775 VPB.n1276 VPB.n1269 0.136
R1776 VPB.n1281 VPB.n1276 0.136
R1777 VPB.n1286 VPB.n1281 0.136
R1778 VPB.n1290 VPB.n1286 0.136
R1779 VPB.n1294 VPB.n1290 0.136
R1780 VPB.n1325 VPB.n1321 0.136
R1781 VPB.n1330 VPB.n1325 0.136
R1782 VPB.n1335 VPB.n1330 0.136
R1783 VPB.n1342 VPB.n1335 0.136
R1784 VPB.n1347 VPB.n1342 0.136
R1785 VPB.n1352 VPB.n1347 0.136
R1786 VPB.n1359 VPB.n1352 0.136
R1787 VPB.n1364 VPB.n1359 0.136
R1788 VPB.n1369 VPB.n1364 0.136
R1789 VPB.n1373 VPB.n1369 0.136
R1790 VPB.n1377 VPB.n1373 0.136
R1791 VPB.n1408 VPB.n1404 0.136
R1792 VPB.n1413 VPB.n1408 0.136
R1793 VPB.n1418 VPB.n1413 0.136
R1794 VPB.n1425 VPB.n1418 0.136
R1795 VPB.n1430 VPB.n1425 0.136
R1796 VPB.n1435 VPB.n1430 0.136
R1797 VPB.n1442 VPB.n1435 0.136
R1798 VPB.n1447 VPB.n1442 0.136
R1799 VPB.n1452 VPB.n1447 0.136
R1800 VPB.n1456 VPB.n1452 0.136
R1801 VPB.n1460 VPB.n1456 0.136
R1802 VPB.n1491 VPB.n1487 0.136
R1803 VPB.n1496 VPB.n1491 0.136
R1804 VPB.n1501 VPB.n1496 0.136
R1805 VPB.n1508 VPB.n1501 0.136
R1806 VPB.n1513 VPB.n1508 0.136
R1807 VPB.n1518 VPB.n1513 0.136
R1808 VPB.n1525 VPB.n1518 0.136
R1809 VPB.n1530 VPB.n1525 0.136
R1810 VPB.n1535 VPB.n1530 0.136
R1811 VPB.n1539 VPB.n1535 0.136
R1812 VPB.n1543 VPB.n1539 0.136
R1813 VPB.n1574 VPB.n1570 0.136
R1814 VPB.n1579 VPB.n1574 0.136
R1815 VPB.n1584 VPB.n1579 0.136
R1816 VPB.n1591 VPB.n1584 0.136
R1817 VPB.n1596 VPB.n1591 0.136
R1818 VPB.n1601 VPB.n1596 0.136
R1819 VPB.n1608 VPB.n1601 0.136
R1820 VPB.n1613 VPB.n1608 0.136
R1821 VPB.n1618 VPB.n1613 0.136
R1822 VPB.n1622 VPB.n1618 0.136
R1823 VPB.n1626 VPB.n1622 0.136
R1824 VPB.n1657 VPB.n1653 0.136
R1825 VPB.n1662 VPB.n1657 0.136
R1826 VPB.n1667 VPB.n1662 0.136
R1827 VPB.n1674 VPB.n1667 0.136
R1828 VPB.n1679 VPB.n1674 0.136
R1829 VPB.n1684 VPB.n1679 0.136
R1830 VPB.n1691 VPB.n1684 0.136
R1831 VPB.n1696 VPB.n1691 0.136
R1832 VPB.n1701 VPB.n1696 0.136
R1833 VPB.n1705 VPB.n1701 0.136
R1834 VPB.n1709 VPB.n1705 0.136
R1835 VPB.n1711 VPB.n1710 0.136
R1836 VPB.n1712 VPB.n1711 0.136
R1837 VPB.n1713 VPB.n1712 0.136
R1838 VPB.n1714 VPB.n1713 0.136
R1839 VPB.n1715 VPB.n1714 0.136
R1840 VPB.n1716 VPB.n1715 0.136
R1841 VPB.n1717 VPB.n1716 0.136
R1842 VPB.n1718 VPB.n1717 0.136
R1843 VPB.n1719 VPB.n1718 0.136
R1844 VPB.n1720 VPB.n1719 0.136
R1845 VPB.n1721 VPB.n1720 0.136
R1846 VPB.n945 VPB 0.068
R1847 VPB.n954 VPB 0.068
R1848 a_4447_943.n7 a_4447_943.t7 512.525
R1849 a_4447_943.n5 a_4447_943.t14 477.179
R1850 a_4447_943.n11 a_4447_943.t10 454.685
R1851 a_4447_943.n11 a_4447_943.t13 428.979
R1852 a_4447_943.n5 a_4447_943.t11 406.485
R1853 a_4447_943.n7 a_4447_943.t9 371.139
R1854 a_4447_943.n6 a_4447_943.t12 346.633
R1855 a_4447_943.n8 a_4447_943.t15 340.206
R1856 a_4447_943.n12 a_4447_943.t8 221.453
R1857 a_4447_943.n15 a_4447_943.n13 203.12
R1858 a_4447_943.n13 a_4447_943.n12 156.035
R1859 a_4447_943.n10 a_4447_943.n9 119.618
R1860 a_4447_943.n12 a_4447_943.n11 108.494
R1861 a_4447_943.n13 a_4447_943.n10 106.211
R1862 a_4447_943.n8 a_4447_943.n7 89.615
R1863 a_4447_943.n3 a_4447_943.n2 79.232
R1864 a_4447_943.n9 a_4447_943.n6 78.675
R1865 a_4447_943.n9 a_4447_943.n8 76
R1866 a_4447_943.n10 a_4447_943.n4 74.634
R1867 a_4447_943.n4 a_4447_943.n3 63.152
R1868 a_4447_943.n6 a_4447_943.n5 29.194
R1869 a_4447_943.n4 a_4447_943.n0 16.08
R1870 a_4447_943.n3 a_4447_943.n1 16.08
R1871 a_4447_943.n15 a_4447_943.n14 15.218
R1872 a_4447_943.n0 a_4447_943.t0 14.282
R1873 a_4447_943.n0 a_4447_943.t6 14.282
R1874 a_4447_943.n1 a_4447_943.t2 14.282
R1875 a_4447_943.n1 a_4447_943.t3 14.282
R1876 a_4447_943.n2 a_4447_943.t5 14.282
R1877 a_4447_943.n2 a_4447_943.t4 14.282
R1878 a_4447_943.n16 a_4447_943.n15 12.014
R1879 a_6371_943.n5 a_6371_943.t11 512.525
R1880 a_6371_943.n7 a_6371_943.t12 454.685
R1881 a_6371_943.n7 a_6371_943.t8 428.979
R1882 a_6371_943.n5 a_6371_943.t7 371.139
R1883 a_6371_943.n6 a_6371_943.t10 271.162
R1884 a_6371_943.n8 a_6371_943.t9 221.453
R1885 a_6371_943.n12 a_6371_943.n10 203.12
R1886 a_6371_943.n10 a_6371_943.n4 180.846
R1887 a_6371_943.n6 a_6371_943.n5 172.76
R1888 a_6371_943.n8 a_6371_943.n7 108.494
R1889 a_6371_943.n9 a_6371_943.n6 84.388
R1890 a_6371_943.n9 a_6371_943.n8 80.035
R1891 a_6371_943.n3 a_6371_943.n2 79.232
R1892 a_6371_943.n10 a_6371_943.n9 76
R1893 a_6371_943.n4 a_6371_943.n3 63.152
R1894 a_6371_943.n4 a_6371_943.n0 16.08
R1895 a_6371_943.n3 a_6371_943.n1 16.08
R1896 a_6371_943.n12 a_6371_943.n11 15.218
R1897 a_6371_943.n0 a_6371_943.t3 14.282
R1898 a_6371_943.n0 a_6371_943.t1 14.282
R1899 a_6371_943.n1 a_6371_943.t5 14.282
R1900 a_6371_943.n1 a_6371_943.t4 14.282
R1901 a_6371_943.n2 a_6371_943.t2 14.282
R1902 a_6371_943.n2 a_6371_943.t6 14.282
R1903 a_6371_943.n13 a_6371_943.n12 12.014
R1904 a_7333_943.n8 a_7333_943.t10 454.685
R1905 a_7333_943.n10 a_7333_943.t13 454.685
R1906 a_7333_943.n6 a_7333_943.t12 454.685
R1907 a_7333_943.n8 a_7333_943.t15 428.979
R1908 a_7333_943.n10 a_7333_943.t7 428.979
R1909 a_7333_943.n6 a_7333_943.t14 428.979
R1910 a_7333_943.n9 a_7333_943.t9 248.006
R1911 a_7333_943.n11 a_7333_943.t8 248.006
R1912 a_7333_943.n7 a_7333_943.t11 248.006
R1913 a_7333_943.n16 a_7333_943.n14 223.151
R1914 a_7333_943.n14 a_7333_943.n5 154.293
R1915 a_7333_943.n13 a_7333_943.n7 82.484
R1916 a_7333_943.n9 a_7333_943.n8 81.941
R1917 a_7333_943.n11 a_7333_943.n10 81.941
R1918 a_7333_943.n7 a_7333_943.n6 81.941
R1919 a_7333_943.n12 a_7333_943.n11 79.491
R1920 a_7333_943.n4 a_7333_943.n3 79.232
R1921 a_7333_943.n12 a_7333_943.n9 76
R1922 a_7333_943.n14 a_7333_943.n13 76
R1923 a_7333_943.n5 a_7333_943.n4 63.152
R1924 a_7333_943.n16 a_7333_943.n15 30
R1925 a_7333_943.n17 a_7333_943.n0 24.383
R1926 a_7333_943.n17 a_7333_943.n16 23.684
R1927 a_7333_943.n5 a_7333_943.n1 16.08
R1928 a_7333_943.n4 a_7333_943.n2 16.08
R1929 a_7333_943.n1 a_7333_943.t2 14.282
R1930 a_7333_943.n1 a_7333_943.t3 14.282
R1931 a_7333_943.n2 a_7333_943.t5 14.282
R1932 a_7333_943.n2 a_7333_943.t6 14.282
R1933 a_7333_943.n3 a_7333_943.t0 14.282
R1934 a_7333_943.n3 a_7333_943.t1 14.282
R1935 a_7333_943.n13 a_7333_943.n12 4.035
R1936 a_12143_943.n6 a_12143_943.t12 512.525
R1937 a_12143_943.n8 a_12143_943.t8 454.685
R1938 a_12143_943.n8 a_12143_943.t11 428.979
R1939 a_12143_943.n6 a_12143_943.t10 371.139
R1940 a_12143_943.n7 a_12143_943.t7 271.162
R1941 a_12143_943.n9 a_12143_943.t9 221.453
R1942 a_12143_943.n13 a_12143_943.n11 196.598
R1943 a_12143_943.n11 a_12143_943.n5 180.846
R1944 a_12143_943.n7 a_12143_943.n6 172.76
R1945 a_12143_943.n9 a_12143_943.n8 108.494
R1946 a_12143_943.n10 a_12143_943.n7 84.388
R1947 a_12143_943.n10 a_12143_943.n9 80.035
R1948 a_12143_943.n4 a_12143_943.n3 79.232
R1949 a_12143_943.n11 a_12143_943.n10 76
R1950 a_12143_943.n5 a_12143_943.n4 63.152
R1951 a_12143_943.n13 a_12143_943.n12 30
R1952 a_12143_943.n14 a_12143_943.n0 24.383
R1953 a_12143_943.n14 a_12143_943.n13 23.684
R1954 a_12143_943.n5 a_12143_943.n1 16.08
R1955 a_12143_943.n4 a_12143_943.n2 16.08
R1956 a_12143_943.n1 a_12143_943.t1 14.282
R1957 a_12143_943.n1 a_12143_943.t0 14.282
R1958 a_12143_943.n2 a_12143_943.t6 14.282
R1959 a_12143_943.n2 a_12143_943.t5 14.282
R1960 a_12143_943.n3 a_12143_943.t3 14.282
R1961 a_12143_943.n3 a_12143_943.t4 14.282
R1962 a_15483_75.t0 a_15483_75.n0 117.777
R1963 a_15483_75.n2 a_15483_75.n1 55.228
R1964 a_15483_75.n4 a_15483_75.n3 9.111
R1965 a_15483_75.n8 a_15483_75.n6 7.859
R1966 a_15483_75.t0 a_15483_75.n2 4.04
R1967 a_15483_75.t0 a_15483_75.n8 3.034
R1968 a_15483_75.n6 a_15483_75.n4 1.964
R1969 a_15483_75.n6 a_15483_75.n5 1.964
R1970 a_15483_75.n8 a_15483_75.n7 0.443
R1971 VNB VNB.n1505 300.778
R1972 VNB.n171 VNB.n170 199.897
R1973 VNB.n223 VNB.n222 199.897
R1974 VNB.n282 VNB.n281 199.897
R1975 VNB.n341 VNB.n340 199.897
R1976 VNB.n416 VNB.n415 199.897
R1977 VNB.n484 VNB.n483 199.897
R1978 VNB.n559 VNB.n558 199.897
R1979 VNB.n627 VNB.n626 199.897
R1980 VNB.n695 VNB.n694 199.897
R1981 VNB.n770 VNB.n769 199.897
R1982 VNB.n74 VNB.n73 199.897
R1983 VNB.n871 VNB.n870 199.897
R1984 VNB.n939 VNB.n938 199.897
R1985 VNB.n1007 VNB.n1006 199.897
R1986 VNB.n1075 VNB.n1074 199.897
R1987 VNB.n1150 VNB.n1149 199.897
R1988 VNB.n1218 VNB.n1217 199.897
R1989 VNB.n1286 VNB.n1285 199.897
R1990 VNB.n1354 VNB.n1353 199.897
R1991 VNB.n1422 VNB.n1421 199.897
R1992 VNB.n18 VNB.n17 199.897
R1993 VNB.n232 VNB.n230 154.509
R1994 VNB.n180 VNB.n178 154.509
R1995 VNB.n350 VNB.n348 154.509
R1996 VNB.n291 VNB.n289 154.509
R1997 VNB.n493 VNB.n491 154.509
R1998 VNB.n425 VNB.n423 154.509
R1999 VNB.n636 VNB.n634 154.509
R2000 VNB.n568 VNB.n566 154.509
R2001 VNB.n779 VNB.n777 154.509
R2002 VNB.n704 VNB.n702 154.509
R2003 VNB.n880 VNB.n878 154.509
R2004 VNB.n90 VNB.n88 154.509
R2005 VNB.n1016 VNB.n1014 154.509
R2006 VNB.n948 VNB.n946 154.509
R2007 VNB.n1159 VNB.n1157 154.509
R2008 VNB.n1084 VNB.n1082 154.509
R2009 VNB.n1295 VNB.n1293 154.509
R2010 VNB.n1227 VNB.n1225 154.509
R2011 VNB.n1431 VNB.n1429 154.509
R2012 VNB.n1363 VNB.n1361 154.509
R2013 VNB.n27 VNB.n25 154.509
R2014 VNB.n382 VNB.n381 147.75
R2015 VNB.n525 VNB.n524 147.75
R2016 VNB.n736 VNB.n735 147.75
R2017 VNB.n811 VNB.n810 147.75
R2018 VNB.n838 VNB.n837 147.75
R2019 VNB.n1116 VNB.n1115 147.75
R2020 VNB.n51 VNB.n50 147.75
R2021 VNB.n248 VNB.n247 121.366
R2022 VNB.n307 VNB.n306 121.366
R2023 VNB.n394 VNB.n391 121.366
R2024 VNB.n537 VNB.n534 121.366
R2025 VNB.n748 VNB.n745 121.366
R2026 VNB.n822 VNB.n820 121.366
R2027 VNB.n849 VNB.n846 121.366
R2028 VNB.n1128 VNB.n1125 121.366
R2029 VNB.n56 VNB.n54 121.366
R2030 VNB.n461 VNB.n460 85.559
R2031 VNB.n604 VNB.n603 85.559
R2032 VNB.n672 VNB.n671 85.559
R2033 VNB.n916 VNB.n915 85.559
R2034 VNB.n984 VNB.n983 85.559
R2035 VNB.n1052 VNB.n1051 85.559
R2036 VNB.n1195 VNB.n1194 85.559
R2037 VNB.n1263 VNB.n1262 85.559
R2038 VNB.n1331 VNB.n1330 85.559
R2039 VNB.n1399 VNB.n1398 85.559
R2040 VNB.n1467 VNB.n1466 85.559
R2041 VNB.n200 VNB.n199 84.842
R2042 VNB.n139 VNB.n130 76.136
R2043 VNB.n139 VNB.n138 76
R2044 VNB.n1492 VNB.n1491 76
R2045 VNB.n1479 VNB.n1478 76
R2046 VNB.n1475 VNB.n1474 76
R2047 VNB.n1471 VNB.n1470 76
R2048 VNB.n1465 VNB.n1464 76
R2049 VNB.n1461 VNB.n1460 76
R2050 VNB.n1457 VNB.n1456 76
R2051 VNB.n1453 VNB.n1452 76
R2052 VNB.n1449 VNB.n1448 76
R2053 VNB.n1445 VNB.n1444 76
R2054 VNB.n1441 VNB.n1440 76
R2055 VNB.n1437 VNB.n1436 76
R2056 VNB.n1433 VNB.n1432 76
R2057 VNB.n1411 VNB.n1410 76
R2058 VNB.n1407 VNB.n1406 76
R2059 VNB.n1403 VNB.n1402 76
R2060 VNB.n1397 VNB.n1396 76
R2061 VNB.n1393 VNB.n1392 76
R2062 VNB.n1389 VNB.n1388 76
R2063 VNB.n1385 VNB.n1384 76
R2064 VNB.n1381 VNB.n1380 76
R2065 VNB.n1377 VNB.n1376 76
R2066 VNB.n1373 VNB.n1372 76
R2067 VNB.n1369 VNB.n1368 76
R2068 VNB.n1365 VNB.n1364 76
R2069 VNB.n1343 VNB.n1342 76
R2070 VNB.n1339 VNB.n1338 76
R2071 VNB.n1335 VNB.n1334 76
R2072 VNB.n1329 VNB.n1328 76
R2073 VNB.n1325 VNB.n1324 76
R2074 VNB.n1321 VNB.n1320 76
R2075 VNB.n1317 VNB.n1316 76
R2076 VNB.n1313 VNB.n1312 76
R2077 VNB.n1309 VNB.n1308 76
R2078 VNB.n1305 VNB.n1304 76
R2079 VNB.n1301 VNB.n1300 76
R2080 VNB.n1297 VNB.n1296 76
R2081 VNB.n1275 VNB.n1274 76
R2082 VNB.n1271 VNB.n1270 76
R2083 VNB.n1267 VNB.n1266 76
R2084 VNB.n1261 VNB.n1260 76
R2085 VNB.n1257 VNB.n1256 76
R2086 VNB.n1253 VNB.n1252 76
R2087 VNB.n1249 VNB.n1248 76
R2088 VNB.n1245 VNB.n1244 76
R2089 VNB.n1241 VNB.n1240 76
R2090 VNB.n1237 VNB.n1236 76
R2091 VNB.n1233 VNB.n1232 76
R2092 VNB.n1229 VNB.n1228 76
R2093 VNB.n1207 VNB.n1206 76
R2094 VNB.n1203 VNB.n1202 76
R2095 VNB.n1199 VNB.n1198 76
R2096 VNB.n1193 VNB.n1192 76
R2097 VNB.n1189 VNB.n1188 76
R2098 VNB.n1185 VNB.n1184 76
R2099 VNB.n1181 VNB.n1180 76
R2100 VNB.n1177 VNB.n1176 76
R2101 VNB.n1173 VNB.n1172 76
R2102 VNB.n1169 VNB.n1168 76
R2103 VNB.n1165 VNB.n1164 76
R2104 VNB.n1161 VNB.n1160 76
R2105 VNB.n1139 VNB.n1138 76
R2106 VNB.n1135 VNB.n1134 76
R2107 VNB.n1131 VNB.n1130 76
R2108 VNB.n1119 VNB.n1118 76
R2109 VNB.n1114 VNB.n1113 76
R2110 VNB.n1110 VNB.n1109 76
R2111 VNB.n1106 VNB.n1105 76
R2112 VNB.n1102 VNB.n1101 76
R2113 VNB.n1098 VNB.n1097 76
R2114 VNB.n1094 VNB.n1093 76
R2115 VNB.n1090 VNB.n1089 76
R2116 VNB.n1086 VNB.n1085 76
R2117 VNB.n1064 VNB.n1063 76
R2118 VNB.n1060 VNB.n1059 76
R2119 VNB.n1056 VNB.n1055 76
R2120 VNB.n1050 VNB.n1049 76
R2121 VNB.n1046 VNB.n1045 76
R2122 VNB.n1042 VNB.n1041 76
R2123 VNB.n1038 VNB.n1037 76
R2124 VNB.n1034 VNB.n1033 76
R2125 VNB.n1030 VNB.n1029 76
R2126 VNB.n1026 VNB.n1025 76
R2127 VNB.n1022 VNB.n1021 76
R2128 VNB.n1018 VNB.n1017 76
R2129 VNB.n996 VNB.n995 76
R2130 VNB.n992 VNB.n991 76
R2131 VNB.n988 VNB.n987 76
R2132 VNB.n982 VNB.n981 76
R2133 VNB.n978 VNB.n977 76
R2134 VNB.n974 VNB.n973 76
R2135 VNB.n970 VNB.n969 76
R2136 VNB.n966 VNB.n965 76
R2137 VNB.n962 VNB.n961 76
R2138 VNB.n958 VNB.n957 76
R2139 VNB.n954 VNB.n953 76
R2140 VNB.n950 VNB.n949 76
R2141 VNB.n928 VNB.n927 76
R2142 VNB.n924 VNB.n923 76
R2143 VNB.n920 VNB.n919 76
R2144 VNB.n914 VNB.n913 76
R2145 VNB.n910 VNB.n909 76
R2146 VNB.n906 VNB.n905 76
R2147 VNB.n902 VNB.n901 76
R2148 VNB.n898 VNB.n897 76
R2149 VNB.n894 VNB.n893 76
R2150 VNB.n890 VNB.n889 76
R2151 VNB.n886 VNB.n885 76
R2152 VNB.n882 VNB.n881 76
R2153 VNB.n860 VNB.n859 76
R2154 VNB.n856 VNB.n855 76
R2155 VNB.n852 VNB.n851 76
R2156 VNB.n840 VNB.n836 76
R2157 VNB.n825 VNB.n824 76
R2158 VNB.n814 VNB.n813 76
R2159 VNB.n809 VNB.n808 76
R2160 VNB.n805 VNB.n804 76
R2161 VNB.n801 VNB.n800 76
R2162 VNB.n797 VNB.n796 76
R2163 VNB.n793 VNB.n792 76
R2164 VNB.n789 VNB.n788 76
R2165 VNB.n785 VNB.n784 76
R2166 VNB.n781 VNB.n780 76
R2167 VNB.n759 VNB.n758 76
R2168 VNB.n755 VNB.n754 76
R2169 VNB.n751 VNB.n750 76
R2170 VNB.n739 VNB.n738 76
R2171 VNB.n734 VNB.n733 76
R2172 VNB.n730 VNB.n729 76
R2173 VNB.n726 VNB.n725 76
R2174 VNB.n722 VNB.n721 76
R2175 VNB.n718 VNB.n717 76
R2176 VNB.n714 VNB.n713 76
R2177 VNB.n710 VNB.n709 76
R2178 VNB.n706 VNB.n705 76
R2179 VNB.n684 VNB.n683 76
R2180 VNB.n680 VNB.n679 76
R2181 VNB.n676 VNB.n675 76
R2182 VNB.n670 VNB.n669 76
R2183 VNB.n666 VNB.n665 76
R2184 VNB.n662 VNB.n661 76
R2185 VNB.n658 VNB.n657 76
R2186 VNB.n654 VNB.n653 76
R2187 VNB.n650 VNB.n649 76
R2188 VNB.n646 VNB.n645 76
R2189 VNB.n642 VNB.n641 76
R2190 VNB.n638 VNB.n637 76
R2191 VNB.n616 VNB.n615 76
R2192 VNB.n612 VNB.n611 76
R2193 VNB.n608 VNB.n607 76
R2194 VNB.n602 VNB.n601 76
R2195 VNB.n598 VNB.n597 76
R2196 VNB.n594 VNB.n593 76
R2197 VNB.n590 VNB.n589 76
R2198 VNB.n586 VNB.n585 76
R2199 VNB.n582 VNB.n581 76
R2200 VNB.n578 VNB.n577 76
R2201 VNB.n574 VNB.n573 76
R2202 VNB.n570 VNB.n569 76
R2203 VNB.n548 VNB.n547 76
R2204 VNB.n544 VNB.n543 76
R2205 VNB.n540 VNB.n539 76
R2206 VNB.n528 VNB.n527 76
R2207 VNB.n523 VNB.n522 76
R2208 VNB.n519 VNB.n518 76
R2209 VNB.n515 VNB.n514 76
R2210 VNB.n511 VNB.n510 76
R2211 VNB.n507 VNB.n506 76
R2212 VNB.n503 VNB.n502 76
R2213 VNB.n499 VNB.n498 76
R2214 VNB.n495 VNB.n494 76
R2215 VNB.n473 VNB.n472 76
R2216 VNB.n469 VNB.n468 76
R2217 VNB.n465 VNB.n464 76
R2218 VNB.n459 VNB.n458 76
R2219 VNB.n455 VNB.n454 76
R2220 VNB.n451 VNB.n450 76
R2221 VNB.n447 VNB.n446 76
R2222 VNB.n443 VNB.n442 76
R2223 VNB.n439 VNB.n438 76
R2224 VNB.n435 VNB.n434 76
R2225 VNB.n431 VNB.n430 76
R2226 VNB.n427 VNB.n426 76
R2227 VNB.n405 VNB.n404 76
R2228 VNB.n401 VNB.n400 76
R2229 VNB.n397 VNB.n396 76
R2230 VNB.n385 VNB.n384 76
R2231 VNB.n380 VNB.n379 76
R2232 VNB.n376 VNB.n375 76
R2233 VNB.n372 VNB.n371 76
R2234 VNB.n368 VNB.n367 76
R2235 VNB.n364 VNB.n363 76
R2236 VNB.n360 VNB.n359 76
R2237 VNB.n356 VNB.n355 76
R2238 VNB.n352 VNB.n351 76
R2239 VNB.n330 VNB.n329 76
R2240 VNB.n326 VNB.n325 76
R2241 VNB.n322 VNB.n321 76
R2242 VNB.n311 VNB.n310 76
R2243 VNB.n305 VNB.n304 76
R2244 VNB.n301 VNB.n300 76
R2245 VNB.n297 VNB.n296 76
R2246 VNB.n293 VNB.n292 76
R2247 VNB.n271 VNB.n270 76
R2248 VNB.n267 VNB.n266 76
R2249 VNB.n263 VNB.n262 76
R2250 VNB.n252 VNB.n251 76
R2251 VNB.n246 VNB.n245 76
R2252 VNB.n242 VNB.n241 76
R2253 VNB.n238 VNB.n237 76
R2254 VNB.n234 VNB.n233 76
R2255 VNB.n212 VNB.n211 76
R2256 VNB.n208 VNB.n207 76
R2257 VNB.n204 VNB.n203 76
R2258 VNB.n198 VNB.n197 76
R2259 VNB.n194 VNB.n193 76
R2260 VNB.n190 VNB.n189 76
R2261 VNB.n186 VNB.n185 76
R2262 VNB.n182 VNB.n181 76
R2263 VNB.n160 VNB.n159 76
R2264 VNB.n156 VNB.n155 76
R2265 VNB.n148 VNB.n147 76
R2266 VNB.n81 VNB.n80 73.875
R2267 VNB.n61 VNB.n60 73.875
R2268 VNB.n390 VNB.n389 64.552
R2269 VNB.n533 VNB.n532 64.552
R2270 VNB.n744 VNB.n743 64.552
R2271 VNB.n819 VNB.n818 64.552
R2272 VNB.n845 VNB.n844 64.552
R2273 VNB.n1124 VNB.n1123 64.552
R2274 VNB.n59 VNB.n7 64.552
R2275 VNB.n257 VNB.n256 63.835
R2276 VNB.n316 VNB.n315 63.835
R2277 VNB.n146 VNB.n145 49.896
R2278 VNB.n463 VNB.n462 41.971
R2279 VNB.n606 VNB.n605 41.971
R2280 VNB.n674 VNB.n673 41.971
R2281 VNB.n918 VNB.n917 41.971
R2282 VNB.n986 VNB.n985 41.971
R2283 VNB.n1054 VNB.n1053 41.971
R2284 VNB.n1197 VNB.n1196 41.971
R2285 VNB.n1265 VNB.n1264 41.971
R2286 VNB.n1333 VNB.n1332 41.971
R2287 VNB.n1401 VNB.n1400 41.971
R2288 VNB.n1469 VNB.n1468 41.971
R2289 VNB.n249 VNB.n248 36.937
R2290 VNB.n308 VNB.n307 36.937
R2291 VNB.n394 VNB.n393 36.937
R2292 VNB.n537 VNB.n536 36.937
R2293 VNB.n748 VNB.n747 36.937
R2294 VNB.n822 VNB.n821 36.937
R2295 VNB.n849 VNB.n848 36.937
R2296 VNB.n1128 VNB.n1127 36.937
R2297 VNB.n56 VNB.n55 36.937
R2298 VNB.n202 VNB.n201 36.678
R2299 VNB.n134 VNB.n133 35.01
R2300 VNB.n393 VNB.n392 29.844
R2301 VNB.n536 VNB.n535 29.844
R2302 VNB.n747 VNB.n746 29.844
R2303 VNB.n848 VNB.n847 29.844
R2304 VNB.n1127 VNB.n1126 29.844
R2305 VNB.n132 VNB.n131 29.127
R2306 VNB.n256 VNB.n255 28.421
R2307 VNB.n315 VNB.n314 28.421
R2308 VNB.n389 VNB.n388 28.421
R2309 VNB.n532 VNB.n531 28.421
R2310 VNB.n743 VNB.n742 28.421
R2311 VNB.n818 VNB.n817 28.421
R2312 VNB.n844 VNB.n843 28.421
R2313 VNB.n1123 VNB.n1122 28.421
R2314 VNB.n7 VNB.n6 28.421
R2315 VNB.n260 VNB.n259 27.855
R2316 VNB.n319 VNB.n318 27.855
R2317 VNB.n256 VNB.n254 25.263
R2318 VNB.n315 VNB.n313 25.263
R2319 VNB.n389 VNB.n387 25.263
R2320 VNB.n532 VNB.n530 25.263
R2321 VNB.n743 VNB.n741 25.263
R2322 VNB.n818 VNB.n816 25.263
R2323 VNB.n844 VNB.n842 25.263
R2324 VNB.n1123 VNB.n1121 25.263
R2325 VNB.n7 VNB.n5 25.263
R2326 VNB.n254 VNB.n253 24.383
R2327 VNB.n313 VNB.n312 24.383
R2328 VNB.n387 VNB.n386 24.383
R2329 VNB.n530 VNB.n529 24.383
R2330 VNB.n741 VNB.n740 24.383
R2331 VNB.n816 VNB.n815 24.383
R2332 VNB.n842 VNB.n841 24.383
R2333 VNB.n1121 VNB.n1120 24.383
R2334 VNB.n5 VNB.n4 24.383
R2335 VNB.n142 VNB.t19 20.794
R2336 VNB.n130 VNB.n127 20.452
R2337 VNB.n1493 VNB.n1492 20.452
R2338 VNB.n135 VNB.n134 20.094
R2339 VNB.n144 VNB.n143 20.094
R2340 VNB.n152 VNB.n151 20.094
R2341 VNB.n134 VNB.n132 19.017
R2342 VNB.n261 VNB.n260 16.721
R2343 VNB.n320 VNB.n319 16.721
R2344 VNB.n138 VNB.n137 13.653
R2345 VNB.n137 VNB.n136 13.653
R2346 VNB.n147 VNB.n146 13.653
R2347 VNB.n155 VNB.n154 13.653
R2348 VNB.n154 VNB.n153 13.653
R2349 VNB.n159 VNB.n158 13.653
R2350 VNB.n158 VNB.n157 13.653
R2351 VNB.n181 VNB.n180 13.653
R2352 VNB.n180 VNB.n179 13.653
R2353 VNB.n185 VNB.n184 13.653
R2354 VNB.n184 VNB.n183 13.653
R2355 VNB.n189 VNB.n188 13.653
R2356 VNB.n188 VNB.n187 13.653
R2357 VNB.n193 VNB.n192 13.653
R2358 VNB.n192 VNB.n191 13.653
R2359 VNB.n197 VNB.n196 13.653
R2360 VNB.n196 VNB.n195 13.653
R2361 VNB.n203 VNB.n202 13.653
R2362 VNB.n207 VNB.n206 13.653
R2363 VNB.n206 VNB.n205 13.653
R2364 VNB.n211 VNB.n210 13.653
R2365 VNB.n210 VNB.n209 13.653
R2366 VNB.n233 VNB.n232 13.653
R2367 VNB.n232 VNB.n231 13.653
R2368 VNB.n237 VNB.n236 13.653
R2369 VNB.n236 VNB.n235 13.653
R2370 VNB.n241 VNB.n240 13.653
R2371 VNB.n240 VNB.n239 13.653
R2372 VNB.n245 VNB.n244 13.653
R2373 VNB.n244 VNB.n243 13.653
R2374 VNB.n251 VNB.n250 13.653
R2375 VNB.n250 VNB.n249 13.653
R2376 VNB.n262 VNB.n261 13.653
R2377 VNB.n266 VNB.n265 13.653
R2378 VNB.n265 VNB.n264 13.653
R2379 VNB.n270 VNB.n269 13.653
R2380 VNB.n269 VNB.n268 13.653
R2381 VNB.n292 VNB.n291 13.653
R2382 VNB.n291 VNB.n290 13.653
R2383 VNB.n296 VNB.n295 13.653
R2384 VNB.n295 VNB.n294 13.653
R2385 VNB.n300 VNB.n299 13.653
R2386 VNB.n299 VNB.n298 13.653
R2387 VNB.n304 VNB.n303 13.653
R2388 VNB.n303 VNB.n302 13.653
R2389 VNB.n310 VNB.n309 13.653
R2390 VNB.n309 VNB.n308 13.653
R2391 VNB.n321 VNB.n320 13.653
R2392 VNB.n325 VNB.n324 13.653
R2393 VNB.n324 VNB.n323 13.653
R2394 VNB.n329 VNB.n328 13.653
R2395 VNB.n328 VNB.n327 13.653
R2396 VNB.n351 VNB.n350 13.653
R2397 VNB.n350 VNB.n349 13.653
R2398 VNB.n355 VNB.n354 13.653
R2399 VNB.n354 VNB.n353 13.653
R2400 VNB.n359 VNB.n358 13.653
R2401 VNB.n358 VNB.n357 13.653
R2402 VNB.n363 VNB.n362 13.653
R2403 VNB.n362 VNB.n361 13.653
R2404 VNB.n367 VNB.n366 13.653
R2405 VNB.n366 VNB.n365 13.653
R2406 VNB.n371 VNB.n370 13.653
R2407 VNB.n370 VNB.n369 13.653
R2408 VNB.n375 VNB.n374 13.653
R2409 VNB.n374 VNB.n373 13.653
R2410 VNB.n379 VNB.n378 13.653
R2411 VNB.n378 VNB.n377 13.653
R2412 VNB.n384 VNB.n383 13.653
R2413 VNB.n383 VNB.n382 13.653
R2414 VNB.n396 VNB.n395 13.653
R2415 VNB.n395 VNB.n394 13.653
R2416 VNB.n400 VNB.n399 13.653
R2417 VNB.n399 VNB.n398 13.653
R2418 VNB.n404 VNB.n403 13.653
R2419 VNB.n403 VNB.n402 13.653
R2420 VNB.n426 VNB.n425 13.653
R2421 VNB.n425 VNB.n424 13.653
R2422 VNB.n430 VNB.n429 13.653
R2423 VNB.n429 VNB.n428 13.653
R2424 VNB.n434 VNB.n433 13.653
R2425 VNB.n433 VNB.n432 13.653
R2426 VNB.n438 VNB.n437 13.653
R2427 VNB.n437 VNB.n436 13.653
R2428 VNB.n442 VNB.n441 13.653
R2429 VNB.n441 VNB.n440 13.653
R2430 VNB.n446 VNB.n445 13.653
R2431 VNB.n445 VNB.n444 13.653
R2432 VNB.n450 VNB.n449 13.653
R2433 VNB.n449 VNB.n448 13.653
R2434 VNB.n454 VNB.n453 13.653
R2435 VNB.n453 VNB.n452 13.653
R2436 VNB.n458 VNB.n457 13.653
R2437 VNB.n457 VNB.n456 13.653
R2438 VNB.n464 VNB.n463 13.653
R2439 VNB.n468 VNB.n467 13.653
R2440 VNB.n467 VNB.n466 13.653
R2441 VNB.n472 VNB.n471 13.653
R2442 VNB.n471 VNB.n470 13.653
R2443 VNB.n494 VNB.n493 13.653
R2444 VNB.n493 VNB.n492 13.653
R2445 VNB.n498 VNB.n497 13.653
R2446 VNB.n497 VNB.n496 13.653
R2447 VNB.n502 VNB.n501 13.653
R2448 VNB.n501 VNB.n500 13.653
R2449 VNB.n506 VNB.n505 13.653
R2450 VNB.n505 VNB.n504 13.653
R2451 VNB.n510 VNB.n509 13.653
R2452 VNB.n509 VNB.n508 13.653
R2453 VNB.n514 VNB.n513 13.653
R2454 VNB.n513 VNB.n512 13.653
R2455 VNB.n518 VNB.n517 13.653
R2456 VNB.n517 VNB.n516 13.653
R2457 VNB.n522 VNB.n521 13.653
R2458 VNB.n521 VNB.n520 13.653
R2459 VNB.n527 VNB.n526 13.653
R2460 VNB.n526 VNB.n525 13.653
R2461 VNB.n539 VNB.n538 13.653
R2462 VNB.n538 VNB.n537 13.653
R2463 VNB.n543 VNB.n542 13.653
R2464 VNB.n542 VNB.n541 13.653
R2465 VNB.n547 VNB.n546 13.653
R2466 VNB.n546 VNB.n545 13.653
R2467 VNB.n569 VNB.n568 13.653
R2468 VNB.n568 VNB.n567 13.653
R2469 VNB.n573 VNB.n572 13.653
R2470 VNB.n572 VNB.n571 13.653
R2471 VNB.n577 VNB.n576 13.653
R2472 VNB.n576 VNB.n575 13.653
R2473 VNB.n581 VNB.n580 13.653
R2474 VNB.n580 VNB.n579 13.653
R2475 VNB.n585 VNB.n584 13.653
R2476 VNB.n584 VNB.n583 13.653
R2477 VNB.n589 VNB.n588 13.653
R2478 VNB.n588 VNB.n587 13.653
R2479 VNB.n593 VNB.n592 13.653
R2480 VNB.n592 VNB.n591 13.653
R2481 VNB.n597 VNB.n596 13.653
R2482 VNB.n596 VNB.n595 13.653
R2483 VNB.n601 VNB.n600 13.653
R2484 VNB.n600 VNB.n599 13.653
R2485 VNB.n607 VNB.n606 13.653
R2486 VNB.n611 VNB.n610 13.653
R2487 VNB.n610 VNB.n609 13.653
R2488 VNB.n615 VNB.n614 13.653
R2489 VNB.n614 VNB.n613 13.653
R2490 VNB.n637 VNB.n636 13.653
R2491 VNB.n636 VNB.n635 13.653
R2492 VNB.n641 VNB.n640 13.653
R2493 VNB.n640 VNB.n639 13.653
R2494 VNB.n645 VNB.n644 13.653
R2495 VNB.n644 VNB.n643 13.653
R2496 VNB.n649 VNB.n648 13.653
R2497 VNB.n648 VNB.n647 13.653
R2498 VNB.n653 VNB.n652 13.653
R2499 VNB.n652 VNB.n651 13.653
R2500 VNB.n657 VNB.n656 13.653
R2501 VNB.n656 VNB.n655 13.653
R2502 VNB.n661 VNB.n660 13.653
R2503 VNB.n660 VNB.n659 13.653
R2504 VNB.n665 VNB.n664 13.653
R2505 VNB.n664 VNB.n663 13.653
R2506 VNB.n669 VNB.n668 13.653
R2507 VNB.n668 VNB.n667 13.653
R2508 VNB.n675 VNB.n674 13.653
R2509 VNB.n679 VNB.n678 13.653
R2510 VNB.n678 VNB.n677 13.653
R2511 VNB.n683 VNB.n682 13.653
R2512 VNB.n682 VNB.n681 13.653
R2513 VNB.n705 VNB.n704 13.653
R2514 VNB.n704 VNB.n703 13.653
R2515 VNB.n709 VNB.n708 13.653
R2516 VNB.n708 VNB.n707 13.653
R2517 VNB.n713 VNB.n712 13.653
R2518 VNB.n712 VNB.n711 13.653
R2519 VNB.n717 VNB.n716 13.653
R2520 VNB.n716 VNB.n715 13.653
R2521 VNB.n721 VNB.n720 13.653
R2522 VNB.n720 VNB.n719 13.653
R2523 VNB.n725 VNB.n724 13.653
R2524 VNB.n724 VNB.n723 13.653
R2525 VNB.n729 VNB.n728 13.653
R2526 VNB.n728 VNB.n727 13.653
R2527 VNB.n733 VNB.n732 13.653
R2528 VNB.n732 VNB.n731 13.653
R2529 VNB.n738 VNB.n737 13.653
R2530 VNB.n737 VNB.n736 13.653
R2531 VNB.n750 VNB.n749 13.653
R2532 VNB.n749 VNB.n748 13.653
R2533 VNB.n754 VNB.n753 13.653
R2534 VNB.n753 VNB.n752 13.653
R2535 VNB.n758 VNB.n757 13.653
R2536 VNB.n757 VNB.n756 13.653
R2537 VNB.n780 VNB.n779 13.653
R2538 VNB.n779 VNB.n778 13.653
R2539 VNB.n784 VNB.n783 13.653
R2540 VNB.n783 VNB.n782 13.653
R2541 VNB.n788 VNB.n787 13.653
R2542 VNB.n787 VNB.n786 13.653
R2543 VNB.n792 VNB.n791 13.653
R2544 VNB.n791 VNB.n790 13.653
R2545 VNB.n796 VNB.n795 13.653
R2546 VNB.n795 VNB.n794 13.653
R2547 VNB.n800 VNB.n799 13.653
R2548 VNB.n799 VNB.n798 13.653
R2549 VNB.n804 VNB.n803 13.653
R2550 VNB.n803 VNB.n802 13.653
R2551 VNB.n808 VNB.n807 13.653
R2552 VNB.n807 VNB.n806 13.653
R2553 VNB.n813 VNB.n812 13.653
R2554 VNB.n812 VNB.n811 13.653
R2555 VNB.n824 VNB.n823 13.653
R2556 VNB.n823 VNB.n822 13.653
R2557 VNB.n83 VNB.n82 13.653
R2558 VNB.n82 VNB.n81 13.653
R2559 VNB.n86 VNB.n85 13.653
R2560 VNB.n85 VNB.n84 13.653
R2561 VNB.n91 VNB.n90 13.653
R2562 VNB.n90 VNB.n89 13.653
R2563 VNB.n94 VNB.n93 13.653
R2564 VNB.n93 VNB.n92 13.653
R2565 VNB.n97 VNB.n96 13.653
R2566 VNB.n96 VNB.n95 13.653
R2567 VNB.n100 VNB.n99 13.653
R2568 VNB.n99 VNB.n98 13.653
R2569 VNB.n103 VNB.n102 13.653
R2570 VNB.n102 VNB.n101 13.653
R2571 VNB.n106 VNB.n105 13.653
R2572 VNB.n105 VNB.n104 13.653
R2573 VNB.n109 VNB.n108 13.653
R2574 VNB.n108 VNB.n107 13.653
R2575 VNB.n112 VNB.n111 13.653
R2576 VNB.n111 VNB.n110 13.653
R2577 VNB.n840 VNB.n839 13.653
R2578 VNB.n839 VNB.n838 13.653
R2579 VNB.n851 VNB.n850 13.653
R2580 VNB.n850 VNB.n849 13.653
R2581 VNB.n855 VNB.n854 13.653
R2582 VNB.n854 VNB.n853 13.653
R2583 VNB.n859 VNB.n858 13.653
R2584 VNB.n858 VNB.n857 13.653
R2585 VNB.n881 VNB.n880 13.653
R2586 VNB.n880 VNB.n879 13.653
R2587 VNB.n885 VNB.n884 13.653
R2588 VNB.n884 VNB.n883 13.653
R2589 VNB.n889 VNB.n888 13.653
R2590 VNB.n888 VNB.n887 13.653
R2591 VNB.n893 VNB.n892 13.653
R2592 VNB.n892 VNB.n891 13.653
R2593 VNB.n897 VNB.n896 13.653
R2594 VNB.n896 VNB.n895 13.653
R2595 VNB.n901 VNB.n900 13.653
R2596 VNB.n900 VNB.n899 13.653
R2597 VNB.n905 VNB.n904 13.653
R2598 VNB.n904 VNB.n903 13.653
R2599 VNB.n909 VNB.n908 13.653
R2600 VNB.n908 VNB.n907 13.653
R2601 VNB.n913 VNB.n912 13.653
R2602 VNB.n912 VNB.n911 13.653
R2603 VNB.n919 VNB.n918 13.653
R2604 VNB.n923 VNB.n922 13.653
R2605 VNB.n922 VNB.n921 13.653
R2606 VNB.n927 VNB.n926 13.653
R2607 VNB.n926 VNB.n925 13.653
R2608 VNB.n949 VNB.n948 13.653
R2609 VNB.n948 VNB.n947 13.653
R2610 VNB.n953 VNB.n952 13.653
R2611 VNB.n952 VNB.n951 13.653
R2612 VNB.n957 VNB.n956 13.653
R2613 VNB.n956 VNB.n955 13.653
R2614 VNB.n961 VNB.n960 13.653
R2615 VNB.n960 VNB.n959 13.653
R2616 VNB.n965 VNB.n964 13.653
R2617 VNB.n964 VNB.n963 13.653
R2618 VNB.n969 VNB.n968 13.653
R2619 VNB.n968 VNB.n967 13.653
R2620 VNB.n973 VNB.n972 13.653
R2621 VNB.n972 VNB.n971 13.653
R2622 VNB.n977 VNB.n976 13.653
R2623 VNB.n976 VNB.n975 13.653
R2624 VNB.n981 VNB.n980 13.653
R2625 VNB.n980 VNB.n979 13.653
R2626 VNB.n987 VNB.n986 13.653
R2627 VNB.n991 VNB.n990 13.653
R2628 VNB.n990 VNB.n989 13.653
R2629 VNB.n995 VNB.n994 13.653
R2630 VNB.n994 VNB.n993 13.653
R2631 VNB.n1017 VNB.n1016 13.653
R2632 VNB.n1016 VNB.n1015 13.653
R2633 VNB.n1021 VNB.n1020 13.653
R2634 VNB.n1020 VNB.n1019 13.653
R2635 VNB.n1025 VNB.n1024 13.653
R2636 VNB.n1024 VNB.n1023 13.653
R2637 VNB.n1029 VNB.n1028 13.653
R2638 VNB.n1028 VNB.n1027 13.653
R2639 VNB.n1033 VNB.n1032 13.653
R2640 VNB.n1032 VNB.n1031 13.653
R2641 VNB.n1037 VNB.n1036 13.653
R2642 VNB.n1036 VNB.n1035 13.653
R2643 VNB.n1041 VNB.n1040 13.653
R2644 VNB.n1040 VNB.n1039 13.653
R2645 VNB.n1045 VNB.n1044 13.653
R2646 VNB.n1044 VNB.n1043 13.653
R2647 VNB.n1049 VNB.n1048 13.653
R2648 VNB.n1048 VNB.n1047 13.653
R2649 VNB.n1055 VNB.n1054 13.653
R2650 VNB.n1059 VNB.n1058 13.653
R2651 VNB.n1058 VNB.n1057 13.653
R2652 VNB.n1063 VNB.n1062 13.653
R2653 VNB.n1062 VNB.n1061 13.653
R2654 VNB.n1085 VNB.n1084 13.653
R2655 VNB.n1084 VNB.n1083 13.653
R2656 VNB.n1089 VNB.n1088 13.653
R2657 VNB.n1088 VNB.n1087 13.653
R2658 VNB.n1093 VNB.n1092 13.653
R2659 VNB.n1092 VNB.n1091 13.653
R2660 VNB.n1097 VNB.n1096 13.653
R2661 VNB.n1096 VNB.n1095 13.653
R2662 VNB.n1101 VNB.n1100 13.653
R2663 VNB.n1100 VNB.n1099 13.653
R2664 VNB.n1105 VNB.n1104 13.653
R2665 VNB.n1104 VNB.n1103 13.653
R2666 VNB.n1109 VNB.n1108 13.653
R2667 VNB.n1108 VNB.n1107 13.653
R2668 VNB.n1113 VNB.n1112 13.653
R2669 VNB.n1112 VNB.n1111 13.653
R2670 VNB.n1118 VNB.n1117 13.653
R2671 VNB.n1117 VNB.n1116 13.653
R2672 VNB.n1130 VNB.n1129 13.653
R2673 VNB.n1129 VNB.n1128 13.653
R2674 VNB.n1134 VNB.n1133 13.653
R2675 VNB.n1133 VNB.n1132 13.653
R2676 VNB.n1138 VNB.n1137 13.653
R2677 VNB.n1137 VNB.n1136 13.653
R2678 VNB.n1160 VNB.n1159 13.653
R2679 VNB.n1159 VNB.n1158 13.653
R2680 VNB.n1164 VNB.n1163 13.653
R2681 VNB.n1163 VNB.n1162 13.653
R2682 VNB.n1168 VNB.n1167 13.653
R2683 VNB.n1167 VNB.n1166 13.653
R2684 VNB.n1172 VNB.n1171 13.653
R2685 VNB.n1171 VNB.n1170 13.653
R2686 VNB.n1176 VNB.n1175 13.653
R2687 VNB.n1175 VNB.n1174 13.653
R2688 VNB.n1180 VNB.n1179 13.653
R2689 VNB.n1179 VNB.n1178 13.653
R2690 VNB.n1184 VNB.n1183 13.653
R2691 VNB.n1183 VNB.n1182 13.653
R2692 VNB.n1188 VNB.n1187 13.653
R2693 VNB.n1187 VNB.n1186 13.653
R2694 VNB.n1192 VNB.n1191 13.653
R2695 VNB.n1191 VNB.n1190 13.653
R2696 VNB.n1198 VNB.n1197 13.653
R2697 VNB.n1202 VNB.n1201 13.653
R2698 VNB.n1201 VNB.n1200 13.653
R2699 VNB.n1206 VNB.n1205 13.653
R2700 VNB.n1205 VNB.n1204 13.653
R2701 VNB.n1228 VNB.n1227 13.653
R2702 VNB.n1227 VNB.n1226 13.653
R2703 VNB.n1232 VNB.n1231 13.653
R2704 VNB.n1231 VNB.n1230 13.653
R2705 VNB.n1236 VNB.n1235 13.653
R2706 VNB.n1235 VNB.n1234 13.653
R2707 VNB.n1240 VNB.n1239 13.653
R2708 VNB.n1239 VNB.n1238 13.653
R2709 VNB.n1244 VNB.n1243 13.653
R2710 VNB.n1243 VNB.n1242 13.653
R2711 VNB.n1248 VNB.n1247 13.653
R2712 VNB.n1247 VNB.n1246 13.653
R2713 VNB.n1252 VNB.n1251 13.653
R2714 VNB.n1251 VNB.n1250 13.653
R2715 VNB.n1256 VNB.n1255 13.653
R2716 VNB.n1255 VNB.n1254 13.653
R2717 VNB.n1260 VNB.n1259 13.653
R2718 VNB.n1259 VNB.n1258 13.653
R2719 VNB.n1266 VNB.n1265 13.653
R2720 VNB.n1270 VNB.n1269 13.653
R2721 VNB.n1269 VNB.n1268 13.653
R2722 VNB.n1274 VNB.n1273 13.653
R2723 VNB.n1273 VNB.n1272 13.653
R2724 VNB.n1296 VNB.n1295 13.653
R2725 VNB.n1295 VNB.n1294 13.653
R2726 VNB.n1300 VNB.n1299 13.653
R2727 VNB.n1299 VNB.n1298 13.653
R2728 VNB.n1304 VNB.n1303 13.653
R2729 VNB.n1303 VNB.n1302 13.653
R2730 VNB.n1308 VNB.n1307 13.653
R2731 VNB.n1307 VNB.n1306 13.653
R2732 VNB.n1312 VNB.n1311 13.653
R2733 VNB.n1311 VNB.n1310 13.653
R2734 VNB.n1316 VNB.n1315 13.653
R2735 VNB.n1315 VNB.n1314 13.653
R2736 VNB.n1320 VNB.n1319 13.653
R2737 VNB.n1319 VNB.n1318 13.653
R2738 VNB.n1324 VNB.n1323 13.653
R2739 VNB.n1323 VNB.n1322 13.653
R2740 VNB.n1328 VNB.n1327 13.653
R2741 VNB.n1327 VNB.n1326 13.653
R2742 VNB.n1334 VNB.n1333 13.653
R2743 VNB.n1338 VNB.n1337 13.653
R2744 VNB.n1337 VNB.n1336 13.653
R2745 VNB.n1342 VNB.n1341 13.653
R2746 VNB.n1341 VNB.n1340 13.653
R2747 VNB.n1364 VNB.n1363 13.653
R2748 VNB.n1363 VNB.n1362 13.653
R2749 VNB.n1368 VNB.n1367 13.653
R2750 VNB.n1367 VNB.n1366 13.653
R2751 VNB.n1372 VNB.n1371 13.653
R2752 VNB.n1371 VNB.n1370 13.653
R2753 VNB.n1376 VNB.n1375 13.653
R2754 VNB.n1375 VNB.n1374 13.653
R2755 VNB.n1380 VNB.n1379 13.653
R2756 VNB.n1379 VNB.n1378 13.653
R2757 VNB.n1384 VNB.n1383 13.653
R2758 VNB.n1383 VNB.n1382 13.653
R2759 VNB.n1388 VNB.n1387 13.653
R2760 VNB.n1387 VNB.n1386 13.653
R2761 VNB.n1392 VNB.n1391 13.653
R2762 VNB.n1391 VNB.n1390 13.653
R2763 VNB.n1396 VNB.n1395 13.653
R2764 VNB.n1395 VNB.n1394 13.653
R2765 VNB.n1402 VNB.n1401 13.653
R2766 VNB.n1406 VNB.n1405 13.653
R2767 VNB.n1405 VNB.n1404 13.653
R2768 VNB.n1410 VNB.n1409 13.653
R2769 VNB.n1409 VNB.n1408 13.653
R2770 VNB.n1432 VNB.n1431 13.653
R2771 VNB.n1431 VNB.n1430 13.653
R2772 VNB.n1436 VNB.n1435 13.653
R2773 VNB.n1435 VNB.n1434 13.653
R2774 VNB.n1440 VNB.n1439 13.653
R2775 VNB.n1439 VNB.n1438 13.653
R2776 VNB.n1444 VNB.n1443 13.653
R2777 VNB.n1443 VNB.n1442 13.653
R2778 VNB.n1448 VNB.n1447 13.653
R2779 VNB.n1447 VNB.n1446 13.653
R2780 VNB.n1452 VNB.n1451 13.653
R2781 VNB.n1451 VNB.n1450 13.653
R2782 VNB.n1456 VNB.n1455 13.653
R2783 VNB.n1455 VNB.n1454 13.653
R2784 VNB.n1460 VNB.n1459 13.653
R2785 VNB.n1459 VNB.n1458 13.653
R2786 VNB.n1464 VNB.n1463 13.653
R2787 VNB.n1463 VNB.n1462 13.653
R2788 VNB.n1470 VNB.n1469 13.653
R2789 VNB.n1474 VNB.n1473 13.653
R2790 VNB.n1473 VNB.n1472 13.653
R2791 VNB.n1478 VNB.n1477 13.653
R2792 VNB.n1477 VNB.n1476 13.653
R2793 VNB.n28 VNB.n27 13.653
R2794 VNB.n27 VNB.n26 13.653
R2795 VNB.n31 VNB.n30 13.653
R2796 VNB.n30 VNB.n29 13.653
R2797 VNB.n34 VNB.n33 13.653
R2798 VNB.n33 VNB.n32 13.653
R2799 VNB.n37 VNB.n36 13.653
R2800 VNB.n36 VNB.n35 13.653
R2801 VNB.n40 VNB.n39 13.653
R2802 VNB.n39 VNB.n38 13.653
R2803 VNB.n43 VNB.n42 13.653
R2804 VNB.n42 VNB.n41 13.653
R2805 VNB.n46 VNB.n45 13.653
R2806 VNB.n45 VNB.n44 13.653
R2807 VNB.n49 VNB.n48 13.653
R2808 VNB.n48 VNB.n47 13.653
R2809 VNB.n53 VNB.n52 13.653
R2810 VNB.n52 VNB.n51 13.653
R2811 VNB.n58 VNB.n57 13.653
R2812 VNB.n57 VNB.n56 13.653
R2813 VNB.n63 VNB.n62 13.653
R2814 VNB.n62 VNB.n61 13.653
R2815 VNB.n1492 VNB.n0 13.653
R2816 VNB VNB.n0 13.653
R2817 VNB.n130 VNB.n129 13.653
R2818 VNB.n129 VNB.n128 13.653
R2819 VNB.n1500 VNB.n1497 13.577
R2820 VNB.n115 VNB.n113 13.276
R2821 VNB.n127 VNB.n115 13.276
R2822 VNB.n163 VNB.n161 13.276
R2823 VNB.n176 VNB.n163 13.276
R2824 VNB.n215 VNB.n213 13.276
R2825 VNB.n228 VNB.n215 13.276
R2826 VNB.n274 VNB.n272 13.276
R2827 VNB.n287 VNB.n274 13.276
R2828 VNB.n333 VNB.n331 13.276
R2829 VNB.n346 VNB.n333 13.276
R2830 VNB.n408 VNB.n406 13.276
R2831 VNB.n421 VNB.n408 13.276
R2832 VNB.n476 VNB.n474 13.276
R2833 VNB.n489 VNB.n476 13.276
R2834 VNB.n551 VNB.n549 13.276
R2835 VNB.n564 VNB.n551 13.276
R2836 VNB.n619 VNB.n617 13.276
R2837 VNB.n632 VNB.n619 13.276
R2838 VNB.n687 VNB.n685 13.276
R2839 VNB.n700 VNB.n687 13.276
R2840 VNB.n762 VNB.n760 13.276
R2841 VNB.n775 VNB.n762 13.276
R2842 VNB.n66 VNB.n64 13.276
R2843 VNB.n79 VNB.n66 13.276
R2844 VNB.n863 VNB.n861 13.276
R2845 VNB.n876 VNB.n863 13.276
R2846 VNB.n931 VNB.n929 13.276
R2847 VNB.n944 VNB.n931 13.276
R2848 VNB.n999 VNB.n997 13.276
R2849 VNB.n1012 VNB.n999 13.276
R2850 VNB.n1067 VNB.n1065 13.276
R2851 VNB.n1080 VNB.n1067 13.276
R2852 VNB.n1142 VNB.n1140 13.276
R2853 VNB.n1155 VNB.n1142 13.276
R2854 VNB.n1210 VNB.n1208 13.276
R2855 VNB.n1223 VNB.n1210 13.276
R2856 VNB.n1278 VNB.n1276 13.276
R2857 VNB.n1291 VNB.n1278 13.276
R2858 VNB.n1346 VNB.n1344 13.276
R2859 VNB.n1359 VNB.n1346 13.276
R2860 VNB.n1414 VNB.n1412 13.276
R2861 VNB.n1427 VNB.n1414 13.276
R2862 VNB.n10 VNB.n8 13.276
R2863 VNB.n23 VNB.n10 13.276
R2864 VNB.n181 VNB.n177 13.276
R2865 VNB.n233 VNB.n229 13.276
R2866 VNB.n292 VNB.n288 13.276
R2867 VNB.n351 VNB.n347 13.276
R2868 VNB.n426 VNB.n422 13.276
R2869 VNB.n494 VNB.n490 13.276
R2870 VNB.n569 VNB.n565 13.276
R2871 VNB.n637 VNB.n633 13.276
R2872 VNB.n705 VNB.n701 13.276
R2873 VNB.n780 VNB.n776 13.276
R2874 VNB.n86 VNB.n83 13.276
R2875 VNB.n87 VNB.n86 13.276
R2876 VNB.n91 VNB.n87 13.276
R2877 VNB.n94 VNB.n91 13.276
R2878 VNB.n97 VNB.n94 13.276
R2879 VNB.n100 VNB.n97 13.276
R2880 VNB.n103 VNB.n100 13.276
R2881 VNB.n106 VNB.n103 13.276
R2882 VNB.n109 VNB.n106 13.276
R2883 VNB.n112 VNB.n109 13.276
R2884 VNB.n840 VNB.n112 13.276
R2885 VNB.n851 VNB.n840 13.276
R2886 VNB.n881 VNB.n877 13.276
R2887 VNB.n949 VNB.n945 13.276
R2888 VNB.n1017 VNB.n1013 13.276
R2889 VNB.n1085 VNB.n1081 13.276
R2890 VNB.n1160 VNB.n1156 13.276
R2891 VNB.n1228 VNB.n1224 13.276
R2892 VNB.n1296 VNB.n1292 13.276
R2893 VNB.n1364 VNB.n1360 13.276
R2894 VNB.n1432 VNB.n1428 13.276
R2895 VNB.n28 VNB.n24 13.276
R2896 VNB.n31 VNB.n28 13.276
R2897 VNB.n34 VNB.n31 13.276
R2898 VNB.n37 VNB.n34 13.276
R2899 VNB.n40 VNB.n37 13.276
R2900 VNB.n43 VNB.n40 13.276
R2901 VNB.n46 VNB.n43 13.276
R2902 VNB.n49 VNB.n46 13.276
R2903 VNB.n53 VNB.n49 13.276
R2904 VNB.n58 VNB.n53 13.276
R2905 VNB.n1492 VNB.n63 13.276
R2906 VNB.n3 VNB.n1 13.276
R2907 VNB.n1493 VNB.n3 13.276
R2908 VNB.n151 VNB.n150 12.837
R2909 VNB.n63 VNB.n59 12.02
R2910 VNB.n150 VNB.n149 7.566
R2911 VNB.n1502 VNB.n1501 7.5
R2912 VNB.n169 VNB.n168 7.5
R2913 VNB.n165 VNB.n164 7.5
R2914 VNB.n163 VNB.n162 7.5
R2915 VNB.n176 VNB.n175 7.5
R2916 VNB.n221 VNB.n220 7.5
R2917 VNB.n217 VNB.n216 7.5
R2918 VNB.n215 VNB.n214 7.5
R2919 VNB.n228 VNB.n227 7.5
R2920 VNB.n280 VNB.n279 7.5
R2921 VNB.n276 VNB.n275 7.5
R2922 VNB.n274 VNB.n273 7.5
R2923 VNB.n287 VNB.n286 7.5
R2924 VNB.n339 VNB.n338 7.5
R2925 VNB.n335 VNB.n334 7.5
R2926 VNB.n333 VNB.n332 7.5
R2927 VNB.n346 VNB.n345 7.5
R2928 VNB.n414 VNB.n413 7.5
R2929 VNB.n410 VNB.n409 7.5
R2930 VNB.n408 VNB.n407 7.5
R2931 VNB.n421 VNB.n420 7.5
R2932 VNB.n482 VNB.n481 7.5
R2933 VNB.n478 VNB.n477 7.5
R2934 VNB.n476 VNB.n475 7.5
R2935 VNB.n489 VNB.n488 7.5
R2936 VNB.n557 VNB.n556 7.5
R2937 VNB.n553 VNB.n552 7.5
R2938 VNB.n551 VNB.n550 7.5
R2939 VNB.n564 VNB.n563 7.5
R2940 VNB.n625 VNB.n624 7.5
R2941 VNB.n621 VNB.n620 7.5
R2942 VNB.n619 VNB.n618 7.5
R2943 VNB.n632 VNB.n631 7.5
R2944 VNB.n693 VNB.n692 7.5
R2945 VNB.n689 VNB.n688 7.5
R2946 VNB.n687 VNB.n686 7.5
R2947 VNB.n700 VNB.n699 7.5
R2948 VNB.n768 VNB.n767 7.5
R2949 VNB.n764 VNB.n763 7.5
R2950 VNB.n762 VNB.n761 7.5
R2951 VNB.n775 VNB.n774 7.5
R2952 VNB.n72 VNB.n71 7.5
R2953 VNB.n68 VNB.n67 7.5
R2954 VNB.n66 VNB.n65 7.5
R2955 VNB.n79 VNB.n78 7.5
R2956 VNB.n869 VNB.n868 7.5
R2957 VNB.n865 VNB.n864 7.5
R2958 VNB.n863 VNB.n862 7.5
R2959 VNB.n876 VNB.n875 7.5
R2960 VNB.n937 VNB.n936 7.5
R2961 VNB.n933 VNB.n932 7.5
R2962 VNB.n931 VNB.n930 7.5
R2963 VNB.n944 VNB.n943 7.5
R2964 VNB.n1005 VNB.n1004 7.5
R2965 VNB.n1001 VNB.n1000 7.5
R2966 VNB.n999 VNB.n998 7.5
R2967 VNB.n1012 VNB.n1011 7.5
R2968 VNB.n1073 VNB.n1072 7.5
R2969 VNB.n1069 VNB.n1068 7.5
R2970 VNB.n1067 VNB.n1066 7.5
R2971 VNB.n1080 VNB.n1079 7.5
R2972 VNB.n1148 VNB.n1147 7.5
R2973 VNB.n1144 VNB.n1143 7.5
R2974 VNB.n1142 VNB.n1141 7.5
R2975 VNB.n1155 VNB.n1154 7.5
R2976 VNB.n1216 VNB.n1215 7.5
R2977 VNB.n1212 VNB.n1211 7.5
R2978 VNB.n1210 VNB.n1209 7.5
R2979 VNB.n1223 VNB.n1222 7.5
R2980 VNB.n1284 VNB.n1283 7.5
R2981 VNB.n1280 VNB.n1279 7.5
R2982 VNB.n1278 VNB.n1277 7.5
R2983 VNB.n1291 VNB.n1290 7.5
R2984 VNB.n1352 VNB.n1351 7.5
R2985 VNB.n1348 VNB.n1347 7.5
R2986 VNB.n1346 VNB.n1345 7.5
R2987 VNB.n1359 VNB.n1358 7.5
R2988 VNB.n1420 VNB.n1419 7.5
R2989 VNB.n1416 VNB.n1415 7.5
R2990 VNB.n1414 VNB.n1413 7.5
R2991 VNB.n1427 VNB.n1426 7.5
R2992 VNB.n16 VNB.n15 7.5
R2993 VNB.n12 VNB.n11 7.5
R2994 VNB.n10 VNB.n9 7.5
R2995 VNB.n23 VNB.n22 7.5
R2996 VNB.n1494 VNB.n1493 7.5
R2997 VNB.n3 VNB.n2 7.5
R2998 VNB.n1499 VNB.n1498 7.5
R2999 VNB.n121 VNB.n120 7.5
R3000 VNB.n117 VNB.n116 7.5
R3001 VNB.n115 VNB.n114 7.5
R3002 VNB.n127 VNB.n126 7.5
R3003 VNB.n177 VNB.n176 7.176
R3004 VNB.n229 VNB.n228 7.176
R3005 VNB.n288 VNB.n287 7.176
R3006 VNB.n347 VNB.n346 7.176
R3007 VNB.n422 VNB.n421 7.176
R3008 VNB.n490 VNB.n489 7.176
R3009 VNB.n565 VNB.n564 7.176
R3010 VNB.n633 VNB.n632 7.176
R3011 VNB.n701 VNB.n700 7.176
R3012 VNB.n776 VNB.n775 7.176
R3013 VNB.n87 VNB.n79 7.176
R3014 VNB.n877 VNB.n876 7.176
R3015 VNB.n945 VNB.n944 7.176
R3016 VNB.n1013 VNB.n1012 7.176
R3017 VNB.n1081 VNB.n1080 7.176
R3018 VNB.n1156 VNB.n1155 7.176
R3019 VNB.n1224 VNB.n1223 7.176
R3020 VNB.n1292 VNB.n1291 7.176
R3021 VNB.n1360 VNB.n1359 7.176
R3022 VNB.n1428 VNB.n1427 7.176
R3023 VNB.n24 VNB.n23 7.176
R3024 VNB.n1504 VNB.n1502 7.011
R3025 VNB.n172 VNB.n169 7.011
R3026 VNB.n167 VNB.n165 7.011
R3027 VNB.n224 VNB.n221 7.011
R3028 VNB.n219 VNB.n217 7.011
R3029 VNB.n283 VNB.n280 7.011
R3030 VNB.n278 VNB.n276 7.011
R3031 VNB.n342 VNB.n339 7.011
R3032 VNB.n337 VNB.n335 7.011
R3033 VNB.n417 VNB.n414 7.011
R3034 VNB.n412 VNB.n410 7.011
R3035 VNB.n485 VNB.n482 7.011
R3036 VNB.n480 VNB.n478 7.011
R3037 VNB.n560 VNB.n557 7.011
R3038 VNB.n555 VNB.n553 7.011
R3039 VNB.n628 VNB.n625 7.011
R3040 VNB.n623 VNB.n621 7.011
R3041 VNB.n696 VNB.n693 7.011
R3042 VNB.n691 VNB.n689 7.011
R3043 VNB.n771 VNB.n768 7.011
R3044 VNB.n766 VNB.n764 7.011
R3045 VNB.n75 VNB.n72 7.011
R3046 VNB.n70 VNB.n68 7.011
R3047 VNB.n872 VNB.n869 7.011
R3048 VNB.n867 VNB.n865 7.011
R3049 VNB.n940 VNB.n937 7.011
R3050 VNB.n935 VNB.n933 7.011
R3051 VNB.n1008 VNB.n1005 7.011
R3052 VNB.n1003 VNB.n1001 7.011
R3053 VNB.n1076 VNB.n1073 7.011
R3054 VNB.n1071 VNB.n1069 7.011
R3055 VNB.n1151 VNB.n1148 7.011
R3056 VNB.n1146 VNB.n1144 7.011
R3057 VNB.n1219 VNB.n1216 7.011
R3058 VNB.n1214 VNB.n1212 7.011
R3059 VNB.n1287 VNB.n1284 7.011
R3060 VNB.n1282 VNB.n1280 7.011
R3061 VNB.n1355 VNB.n1352 7.011
R3062 VNB.n1350 VNB.n1348 7.011
R3063 VNB.n1423 VNB.n1420 7.011
R3064 VNB.n1418 VNB.n1416 7.011
R3065 VNB.n19 VNB.n16 7.011
R3066 VNB.n14 VNB.n12 7.011
R3067 VNB.n123 VNB.n121 7.011
R3068 VNB.n119 VNB.n117 7.011
R3069 VNB.n175 VNB.n174 7.01
R3070 VNB.n167 VNB.n166 7.01
R3071 VNB.n172 VNB.n171 7.01
R3072 VNB.n227 VNB.n226 7.01
R3073 VNB.n219 VNB.n218 7.01
R3074 VNB.n224 VNB.n223 7.01
R3075 VNB.n286 VNB.n285 7.01
R3076 VNB.n278 VNB.n277 7.01
R3077 VNB.n283 VNB.n282 7.01
R3078 VNB.n345 VNB.n344 7.01
R3079 VNB.n337 VNB.n336 7.01
R3080 VNB.n342 VNB.n341 7.01
R3081 VNB.n420 VNB.n419 7.01
R3082 VNB.n412 VNB.n411 7.01
R3083 VNB.n417 VNB.n416 7.01
R3084 VNB.n488 VNB.n487 7.01
R3085 VNB.n480 VNB.n479 7.01
R3086 VNB.n485 VNB.n484 7.01
R3087 VNB.n563 VNB.n562 7.01
R3088 VNB.n555 VNB.n554 7.01
R3089 VNB.n560 VNB.n559 7.01
R3090 VNB.n631 VNB.n630 7.01
R3091 VNB.n623 VNB.n622 7.01
R3092 VNB.n628 VNB.n627 7.01
R3093 VNB.n699 VNB.n698 7.01
R3094 VNB.n691 VNB.n690 7.01
R3095 VNB.n696 VNB.n695 7.01
R3096 VNB.n774 VNB.n773 7.01
R3097 VNB.n766 VNB.n765 7.01
R3098 VNB.n771 VNB.n770 7.01
R3099 VNB.n78 VNB.n77 7.01
R3100 VNB.n70 VNB.n69 7.01
R3101 VNB.n75 VNB.n74 7.01
R3102 VNB.n875 VNB.n874 7.01
R3103 VNB.n867 VNB.n866 7.01
R3104 VNB.n872 VNB.n871 7.01
R3105 VNB.n943 VNB.n942 7.01
R3106 VNB.n935 VNB.n934 7.01
R3107 VNB.n940 VNB.n939 7.01
R3108 VNB.n1011 VNB.n1010 7.01
R3109 VNB.n1003 VNB.n1002 7.01
R3110 VNB.n1008 VNB.n1007 7.01
R3111 VNB.n1079 VNB.n1078 7.01
R3112 VNB.n1071 VNB.n1070 7.01
R3113 VNB.n1076 VNB.n1075 7.01
R3114 VNB.n1154 VNB.n1153 7.01
R3115 VNB.n1146 VNB.n1145 7.01
R3116 VNB.n1151 VNB.n1150 7.01
R3117 VNB.n1222 VNB.n1221 7.01
R3118 VNB.n1214 VNB.n1213 7.01
R3119 VNB.n1219 VNB.n1218 7.01
R3120 VNB.n1290 VNB.n1289 7.01
R3121 VNB.n1282 VNB.n1281 7.01
R3122 VNB.n1287 VNB.n1286 7.01
R3123 VNB.n1358 VNB.n1357 7.01
R3124 VNB.n1350 VNB.n1349 7.01
R3125 VNB.n1355 VNB.n1354 7.01
R3126 VNB.n1426 VNB.n1425 7.01
R3127 VNB.n1418 VNB.n1417 7.01
R3128 VNB.n1423 VNB.n1422 7.01
R3129 VNB.n22 VNB.n21 7.01
R3130 VNB.n14 VNB.n13 7.01
R3131 VNB.n19 VNB.n18 7.01
R3132 VNB.n126 VNB.n125 7.01
R3133 VNB.n119 VNB.n118 7.01
R3134 VNB.n123 VNB.n122 7.01
R3135 VNB.n1504 VNB.n1503 7.01
R3136 VNB.n1500 VNB.n1499 6.788
R3137 VNB.n1495 VNB.n1494 6.788
R3138 VNB.n141 VNB.n140 4.551
R3139 VNB.n138 VNB.n135 4.305
R3140 VNB.n155 VNB.n152 3.947
R3141 VNB.n203 VNB.n200 2.511
R3142 VNB.n262 VNB.n257 2.511
R3143 VNB.n321 VNB.n316 2.511
R3144 VNB.t19 VNB.n141 2.238
R3145 VNB.n260 VNB.n258 1.99
R3146 VNB.n319 VNB.n317 1.99
R3147 VNB.n396 VNB.n390 1.255
R3148 VNB.n464 VNB.n461 1.255
R3149 VNB.n539 VNB.n533 1.255
R3150 VNB.n607 VNB.n604 1.255
R3151 VNB.n675 VNB.n672 1.255
R3152 VNB.n750 VNB.n744 1.255
R3153 VNB.n824 VNB.n819 1.255
R3154 VNB.n851 VNB.n845 1.255
R3155 VNB.n919 VNB.n916 1.255
R3156 VNB.n987 VNB.n984 1.255
R3157 VNB.n1055 VNB.n1052 1.255
R3158 VNB.n1130 VNB.n1124 1.255
R3159 VNB.n1198 VNB.n1195 1.255
R3160 VNB.n1266 VNB.n1263 1.255
R3161 VNB.n1334 VNB.n1331 1.255
R3162 VNB.n1402 VNB.n1399 1.255
R3163 VNB.n1470 VNB.n1467 1.255
R3164 VNB.n59 VNB.n58 1.255
R3165 VNB.n1505 VNB.n1496 0.921
R3166 VNB.n1505 VNB.n1500 0.476
R3167 VNB.n1505 VNB.n1495 0.475
R3168 VNB.n143 VNB.n142 0.358
R3169 VNB.n182 VNB.n160 0.272
R3170 VNB.n234 VNB.n212 0.272
R3171 VNB.n293 VNB.n271 0.272
R3172 VNB.n352 VNB.n330 0.272
R3173 VNB.n427 VNB.n405 0.272
R3174 VNB.n495 VNB.n473 0.272
R3175 VNB.n570 VNB.n548 0.272
R3176 VNB.n638 VNB.n616 0.272
R3177 VNB.n706 VNB.n684 0.272
R3178 VNB.n781 VNB.n759 0.272
R3179 VNB.n828 VNB.n827 0.272
R3180 VNB.n882 VNB.n860 0.272
R3181 VNB.n950 VNB.n928 0.272
R3182 VNB.n1018 VNB.n996 0.272
R3183 VNB.n1086 VNB.n1064 0.272
R3184 VNB.n1161 VNB.n1139 0.272
R3185 VNB.n1229 VNB.n1207 0.272
R3186 VNB.n1297 VNB.n1275 0.272
R3187 VNB.n1365 VNB.n1343 0.272
R3188 VNB.n1433 VNB.n1411 0.272
R3189 VNB.n1480 VNB.n1479 0.272
R3190 VNB.n173 VNB.n167 0.246
R3191 VNB.n174 VNB.n173 0.246
R3192 VNB.n173 VNB.n172 0.246
R3193 VNB.n225 VNB.n219 0.246
R3194 VNB.n226 VNB.n225 0.246
R3195 VNB.n225 VNB.n224 0.246
R3196 VNB.n284 VNB.n278 0.246
R3197 VNB.n285 VNB.n284 0.246
R3198 VNB.n284 VNB.n283 0.246
R3199 VNB.n343 VNB.n337 0.246
R3200 VNB.n344 VNB.n343 0.246
R3201 VNB.n343 VNB.n342 0.246
R3202 VNB.n418 VNB.n412 0.246
R3203 VNB.n419 VNB.n418 0.246
R3204 VNB.n418 VNB.n417 0.246
R3205 VNB.n486 VNB.n480 0.246
R3206 VNB.n487 VNB.n486 0.246
R3207 VNB.n486 VNB.n485 0.246
R3208 VNB.n561 VNB.n555 0.246
R3209 VNB.n562 VNB.n561 0.246
R3210 VNB.n561 VNB.n560 0.246
R3211 VNB.n629 VNB.n623 0.246
R3212 VNB.n630 VNB.n629 0.246
R3213 VNB.n629 VNB.n628 0.246
R3214 VNB.n697 VNB.n691 0.246
R3215 VNB.n698 VNB.n697 0.246
R3216 VNB.n697 VNB.n696 0.246
R3217 VNB.n772 VNB.n766 0.246
R3218 VNB.n773 VNB.n772 0.246
R3219 VNB.n772 VNB.n771 0.246
R3220 VNB.n76 VNB.n70 0.246
R3221 VNB.n77 VNB.n76 0.246
R3222 VNB.n76 VNB.n75 0.246
R3223 VNB.n873 VNB.n867 0.246
R3224 VNB.n874 VNB.n873 0.246
R3225 VNB.n873 VNB.n872 0.246
R3226 VNB.n941 VNB.n935 0.246
R3227 VNB.n942 VNB.n941 0.246
R3228 VNB.n941 VNB.n940 0.246
R3229 VNB.n1009 VNB.n1003 0.246
R3230 VNB.n1010 VNB.n1009 0.246
R3231 VNB.n1009 VNB.n1008 0.246
R3232 VNB.n1077 VNB.n1071 0.246
R3233 VNB.n1078 VNB.n1077 0.246
R3234 VNB.n1077 VNB.n1076 0.246
R3235 VNB.n1152 VNB.n1146 0.246
R3236 VNB.n1153 VNB.n1152 0.246
R3237 VNB.n1152 VNB.n1151 0.246
R3238 VNB.n1220 VNB.n1214 0.246
R3239 VNB.n1221 VNB.n1220 0.246
R3240 VNB.n1220 VNB.n1219 0.246
R3241 VNB.n1288 VNB.n1282 0.246
R3242 VNB.n1289 VNB.n1288 0.246
R3243 VNB.n1288 VNB.n1287 0.246
R3244 VNB.n1356 VNB.n1350 0.246
R3245 VNB.n1357 VNB.n1356 0.246
R3246 VNB.n1356 VNB.n1355 0.246
R3247 VNB.n1424 VNB.n1418 0.246
R3248 VNB.n1425 VNB.n1424 0.246
R3249 VNB.n1424 VNB.n1423 0.246
R3250 VNB.n20 VNB.n14 0.246
R3251 VNB.n21 VNB.n20 0.246
R3252 VNB.n20 VNB.n19 0.246
R3253 VNB.n124 VNB.n119 0.246
R3254 VNB.n125 VNB.n124 0.246
R3255 VNB.n124 VNB.n123 0.246
R3256 VNB.n1505 VNB.n1504 0.246
R3257 VNB.n1491 VNB 0.198
R3258 VNB.n147 VNB.n144 0.179
R3259 VNB.n148 VNB.n139 0.136
R3260 VNB.n156 VNB.n148 0.136
R3261 VNB.n160 VNB.n156 0.136
R3262 VNB.n186 VNB.n182 0.136
R3263 VNB.n190 VNB.n186 0.136
R3264 VNB.n194 VNB.n190 0.136
R3265 VNB.n198 VNB.n194 0.136
R3266 VNB.n204 VNB.n198 0.136
R3267 VNB.n208 VNB.n204 0.136
R3268 VNB.n212 VNB.n208 0.136
R3269 VNB.n238 VNB.n234 0.136
R3270 VNB.n242 VNB.n238 0.136
R3271 VNB.n246 VNB.n242 0.136
R3272 VNB.n252 VNB.n246 0.136
R3273 VNB.n263 VNB.n252 0.136
R3274 VNB.n267 VNB.n263 0.136
R3275 VNB.n271 VNB.n267 0.136
R3276 VNB.n297 VNB.n293 0.136
R3277 VNB.n301 VNB.n297 0.136
R3278 VNB.n305 VNB.n301 0.136
R3279 VNB.n311 VNB.n305 0.136
R3280 VNB.n322 VNB.n311 0.136
R3281 VNB.n326 VNB.n322 0.136
R3282 VNB.n330 VNB.n326 0.136
R3283 VNB.n356 VNB.n352 0.136
R3284 VNB.n360 VNB.n356 0.136
R3285 VNB.n364 VNB.n360 0.136
R3286 VNB.n368 VNB.n364 0.136
R3287 VNB.n372 VNB.n368 0.136
R3288 VNB.n376 VNB.n372 0.136
R3289 VNB.n380 VNB.n376 0.136
R3290 VNB.n385 VNB.n380 0.136
R3291 VNB.n397 VNB.n385 0.136
R3292 VNB.n401 VNB.n397 0.136
R3293 VNB.n405 VNB.n401 0.136
R3294 VNB.n431 VNB.n427 0.136
R3295 VNB.n435 VNB.n431 0.136
R3296 VNB.n439 VNB.n435 0.136
R3297 VNB.n443 VNB.n439 0.136
R3298 VNB.n447 VNB.n443 0.136
R3299 VNB.n451 VNB.n447 0.136
R3300 VNB.n455 VNB.n451 0.136
R3301 VNB.n459 VNB.n455 0.136
R3302 VNB.n465 VNB.n459 0.136
R3303 VNB.n469 VNB.n465 0.136
R3304 VNB.n473 VNB.n469 0.136
R3305 VNB.n499 VNB.n495 0.136
R3306 VNB.n503 VNB.n499 0.136
R3307 VNB.n507 VNB.n503 0.136
R3308 VNB.n511 VNB.n507 0.136
R3309 VNB.n515 VNB.n511 0.136
R3310 VNB.n519 VNB.n515 0.136
R3311 VNB.n523 VNB.n519 0.136
R3312 VNB.n528 VNB.n523 0.136
R3313 VNB.n540 VNB.n528 0.136
R3314 VNB.n544 VNB.n540 0.136
R3315 VNB.n548 VNB.n544 0.136
R3316 VNB.n574 VNB.n570 0.136
R3317 VNB.n578 VNB.n574 0.136
R3318 VNB.n582 VNB.n578 0.136
R3319 VNB.n586 VNB.n582 0.136
R3320 VNB.n590 VNB.n586 0.136
R3321 VNB.n594 VNB.n590 0.136
R3322 VNB.n598 VNB.n594 0.136
R3323 VNB.n602 VNB.n598 0.136
R3324 VNB.n608 VNB.n602 0.136
R3325 VNB.n612 VNB.n608 0.136
R3326 VNB.n616 VNB.n612 0.136
R3327 VNB.n642 VNB.n638 0.136
R3328 VNB.n646 VNB.n642 0.136
R3329 VNB.n650 VNB.n646 0.136
R3330 VNB.n654 VNB.n650 0.136
R3331 VNB.n658 VNB.n654 0.136
R3332 VNB.n662 VNB.n658 0.136
R3333 VNB.n666 VNB.n662 0.136
R3334 VNB.n670 VNB.n666 0.136
R3335 VNB.n676 VNB.n670 0.136
R3336 VNB.n680 VNB.n676 0.136
R3337 VNB.n684 VNB.n680 0.136
R3338 VNB.n710 VNB.n706 0.136
R3339 VNB.n714 VNB.n710 0.136
R3340 VNB.n718 VNB.n714 0.136
R3341 VNB.n722 VNB.n718 0.136
R3342 VNB.n726 VNB.n722 0.136
R3343 VNB.n730 VNB.n726 0.136
R3344 VNB.n734 VNB.n730 0.136
R3345 VNB.n739 VNB.n734 0.136
R3346 VNB.n751 VNB.n739 0.136
R3347 VNB.n755 VNB.n751 0.136
R3348 VNB.n759 VNB.n755 0.136
R3349 VNB.n785 VNB.n781 0.136
R3350 VNB.n789 VNB.n785 0.136
R3351 VNB.n793 VNB.n789 0.136
R3352 VNB.n797 VNB.n793 0.136
R3353 VNB.n801 VNB.n797 0.136
R3354 VNB.n805 VNB.n801 0.136
R3355 VNB.n809 VNB.n805 0.136
R3356 VNB.n814 VNB.n809 0.136
R3357 VNB.n825 VNB.n814 0.136
R3358 VNB.n826 VNB.n825 0.136
R3359 VNB.n827 VNB.n826 0.136
R3360 VNB.n829 VNB.n828 0.136
R3361 VNB.n830 VNB.n829 0.136
R3362 VNB.n831 VNB.n830 0.136
R3363 VNB.n832 VNB.n831 0.136
R3364 VNB.n833 VNB.n832 0.136
R3365 VNB.n834 VNB.n833 0.136
R3366 VNB.n835 VNB.n834 0.136
R3367 VNB.n836 VNB.n835 0.136
R3368 VNB.n856 VNB.n852 0.136
R3369 VNB.n860 VNB.n856 0.136
R3370 VNB.n886 VNB.n882 0.136
R3371 VNB.n890 VNB.n886 0.136
R3372 VNB.n894 VNB.n890 0.136
R3373 VNB.n898 VNB.n894 0.136
R3374 VNB.n902 VNB.n898 0.136
R3375 VNB.n906 VNB.n902 0.136
R3376 VNB.n910 VNB.n906 0.136
R3377 VNB.n914 VNB.n910 0.136
R3378 VNB.n920 VNB.n914 0.136
R3379 VNB.n924 VNB.n920 0.136
R3380 VNB.n928 VNB.n924 0.136
R3381 VNB.n954 VNB.n950 0.136
R3382 VNB.n958 VNB.n954 0.136
R3383 VNB.n962 VNB.n958 0.136
R3384 VNB.n966 VNB.n962 0.136
R3385 VNB.n970 VNB.n966 0.136
R3386 VNB.n974 VNB.n970 0.136
R3387 VNB.n978 VNB.n974 0.136
R3388 VNB.n982 VNB.n978 0.136
R3389 VNB.n988 VNB.n982 0.136
R3390 VNB.n992 VNB.n988 0.136
R3391 VNB.n996 VNB.n992 0.136
R3392 VNB.n1022 VNB.n1018 0.136
R3393 VNB.n1026 VNB.n1022 0.136
R3394 VNB.n1030 VNB.n1026 0.136
R3395 VNB.n1034 VNB.n1030 0.136
R3396 VNB.n1038 VNB.n1034 0.136
R3397 VNB.n1042 VNB.n1038 0.136
R3398 VNB.n1046 VNB.n1042 0.136
R3399 VNB.n1050 VNB.n1046 0.136
R3400 VNB.n1056 VNB.n1050 0.136
R3401 VNB.n1060 VNB.n1056 0.136
R3402 VNB.n1064 VNB.n1060 0.136
R3403 VNB.n1090 VNB.n1086 0.136
R3404 VNB.n1094 VNB.n1090 0.136
R3405 VNB.n1098 VNB.n1094 0.136
R3406 VNB.n1102 VNB.n1098 0.136
R3407 VNB.n1106 VNB.n1102 0.136
R3408 VNB.n1110 VNB.n1106 0.136
R3409 VNB.n1114 VNB.n1110 0.136
R3410 VNB.n1119 VNB.n1114 0.136
R3411 VNB.n1131 VNB.n1119 0.136
R3412 VNB.n1135 VNB.n1131 0.136
R3413 VNB.n1139 VNB.n1135 0.136
R3414 VNB.n1165 VNB.n1161 0.136
R3415 VNB.n1169 VNB.n1165 0.136
R3416 VNB.n1173 VNB.n1169 0.136
R3417 VNB.n1177 VNB.n1173 0.136
R3418 VNB.n1181 VNB.n1177 0.136
R3419 VNB.n1185 VNB.n1181 0.136
R3420 VNB.n1189 VNB.n1185 0.136
R3421 VNB.n1193 VNB.n1189 0.136
R3422 VNB.n1199 VNB.n1193 0.136
R3423 VNB.n1203 VNB.n1199 0.136
R3424 VNB.n1207 VNB.n1203 0.136
R3425 VNB.n1233 VNB.n1229 0.136
R3426 VNB.n1237 VNB.n1233 0.136
R3427 VNB.n1241 VNB.n1237 0.136
R3428 VNB.n1245 VNB.n1241 0.136
R3429 VNB.n1249 VNB.n1245 0.136
R3430 VNB.n1253 VNB.n1249 0.136
R3431 VNB.n1257 VNB.n1253 0.136
R3432 VNB.n1261 VNB.n1257 0.136
R3433 VNB.n1267 VNB.n1261 0.136
R3434 VNB.n1271 VNB.n1267 0.136
R3435 VNB.n1275 VNB.n1271 0.136
R3436 VNB.n1301 VNB.n1297 0.136
R3437 VNB.n1305 VNB.n1301 0.136
R3438 VNB.n1309 VNB.n1305 0.136
R3439 VNB.n1313 VNB.n1309 0.136
R3440 VNB.n1317 VNB.n1313 0.136
R3441 VNB.n1321 VNB.n1317 0.136
R3442 VNB.n1325 VNB.n1321 0.136
R3443 VNB.n1329 VNB.n1325 0.136
R3444 VNB.n1335 VNB.n1329 0.136
R3445 VNB.n1339 VNB.n1335 0.136
R3446 VNB.n1343 VNB.n1339 0.136
R3447 VNB.n1369 VNB.n1365 0.136
R3448 VNB.n1373 VNB.n1369 0.136
R3449 VNB.n1377 VNB.n1373 0.136
R3450 VNB.n1381 VNB.n1377 0.136
R3451 VNB.n1385 VNB.n1381 0.136
R3452 VNB.n1389 VNB.n1385 0.136
R3453 VNB.n1393 VNB.n1389 0.136
R3454 VNB.n1397 VNB.n1393 0.136
R3455 VNB.n1403 VNB.n1397 0.136
R3456 VNB.n1407 VNB.n1403 0.136
R3457 VNB.n1411 VNB.n1407 0.136
R3458 VNB.n1437 VNB.n1433 0.136
R3459 VNB.n1441 VNB.n1437 0.136
R3460 VNB.n1445 VNB.n1441 0.136
R3461 VNB.n1449 VNB.n1445 0.136
R3462 VNB.n1453 VNB.n1449 0.136
R3463 VNB.n1457 VNB.n1453 0.136
R3464 VNB.n1461 VNB.n1457 0.136
R3465 VNB.n1465 VNB.n1461 0.136
R3466 VNB.n1471 VNB.n1465 0.136
R3467 VNB.n1475 VNB.n1471 0.136
R3468 VNB.n1479 VNB.n1475 0.136
R3469 VNB.n1481 VNB.n1480 0.136
R3470 VNB.n1482 VNB.n1481 0.136
R3471 VNB.n1483 VNB.n1482 0.136
R3472 VNB.n1484 VNB.n1483 0.136
R3473 VNB.n1485 VNB.n1484 0.136
R3474 VNB.n1486 VNB.n1485 0.136
R3475 VNB.n1487 VNB.n1486 0.136
R3476 VNB.n1488 VNB.n1487 0.136
R3477 VNB.n1489 VNB.n1488 0.136
R3478 VNB.n1490 VNB.n1489 0.136
R3479 VNB.n1491 VNB.n1490 0.136
R3480 VNB.n836 VNB 0.068
R3481 VNB.n852 VNB 0.068
R3482 a_6049_1004.n8 a_6049_1004.t12 512.525
R3483 a_6049_1004.n6 a_6049_1004.t9 512.525
R3484 a_6049_1004.n8 a_6049_1004.t7 371.139
R3485 a_6049_1004.n6 a_6049_1004.t11 371.139
R3486 a_6049_1004.n11 a_6049_1004.n5 233.952
R3487 a_6049_1004.n9 a_6049_1004.n8 225.866
R3488 a_6049_1004.n7 a_6049_1004.n6 225.866
R3489 a_6049_1004.n9 a_6049_1004.t8 218.057
R3490 a_6049_1004.n7 a_6049_1004.t10 218.057
R3491 a_6049_1004.n13 a_6049_1004.n11 143.492
R3492 a_6049_1004.n10 a_6049_1004.n7 79.491
R3493 a_6049_1004.n4 a_6049_1004.n3 79.232
R3494 a_6049_1004.n11 a_6049_1004.n10 77.315
R3495 a_6049_1004.n10 a_6049_1004.n9 76
R3496 a_6049_1004.n5 a_6049_1004.n4 63.152
R3497 a_6049_1004.n13 a_6049_1004.n12 30
R3498 a_6049_1004.n14 a_6049_1004.n0 24.383
R3499 a_6049_1004.n14 a_6049_1004.n13 23.684
R3500 a_6049_1004.n5 a_6049_1004.n1 16.08
R3501 a_6049_1004.n4 a_6049_1004.n2 16.08
R3502 a_6049_1004.n1 a_6049_1004.t5 14.282
R3503 a_6049_1004.n1 a_6049_1004.t4 14.282
R3504 a_6049_1004.n2 a_6049_1004.t3 14.282
R3505 a_6049_1004.n2 a_6049_1004.t2 14.282
R3506 a_6049_1004.n3 a_6049_1004.t1 14.282
R3507 a_6049_1004.n3 a_6049_1004.t0 14.282
R3508 a_7973_1004.n6 a_7973_1004.t7 512.525
R3509 a_7973_1004.n6 a_7973_1004.t8 371.139
R3510 a_7973_1004.n8 a_7973_1004.n5 233.952
R3511 a_7973_1004.n7 a_7973_1004.n6 225.866
R3512 a_7973_1004.n7 a_7973_1004.t9 218.057
R3513 a_7973_1004.n8 a_7973_1004.n7 153.315
R3514 a_7973_1004.n10 a_7973_1004.n8 143.492
R3515 a_7973_1004.n4 a_7973_1004.n3 79.232
R3516 a_7973_1004.n5 a_7973_1004.n4 63.152
R3517 a_7973_1004.n10 a_7973_1004.n9 30
R3518 a_7973_1004.n11 a_7973_1004.n0 24.383
R3519 a_7973_1004.n11 a_7973_1004.n10 23.684
R3520 a_7973_1004.n5 a_7973_1004.n1 16.08
R3521 a_7973_1004.n4 a_7973_1004.n2 16.08
R3522 a_7973_1004.n1 a_7973_1004.t4 14.282
R3523 a_7973_1004.n1 a_7973_1004.t5 14.282
R3524 a_7973_1004.n2 a_7973_1004.t2 14.282
R3525 a_7973_1004.n2 a_7973_1004.t3 14.282
R3526 a_7973_1004.n3 a_7973_1004.t1 14.282
R3527 a_7973_1004.n3 a_7973_1004.t0 14.282
R3528 a_10219_943.n6 a_10219_943.t7 475.572
R3529 a_10219_943.n8 a_10219_943.t14 469.145
R3530 a_10219_943.n12 a_10219_943.t11 454.685
R3531 a_10219_943.n12 a_10219_943.t15 428.979
R3532 a_10219_943.n8 a_10219_943.t8 384.527
R3533 a_10219_943.n6 a_10219_943.t12 384.527
R3534 a_10219_943.n9 a_10219_943.t9 277.772
R3535 a_10219_943.n7 a_10219_943.t13 277.772
R3536 a_10219_943.n13 a_10219_943.t10 221.453
R3537 a_10219_943.n16 a_10219_943.n14 196.598
R3538 a_10219_943.n14 a_10219_943.n13 156.035
R3539 a_10219_943.n11 a_10219_943.n5 154.293
R3540 a_10219_943.n13 a_10219_943.n12 108.494
R3541 a_10219_943.n11 a_10219_943.n10 99.226
R3542 a_10219_943.n10 a_10219_943.n7 80.851
R3543 a_10219_943.n4 a_10219_943.n3 79.232
R3544 a_10219_943.n10 a_10219_943.n9 76
R3545 a_10219_943.n7 a_10219_943.n6 67.889
R3546 a_10219_943.n9 a_10219_943.n8 66.88
R3547 a_10219_943.n5 a_10219_943.n4 63.152
R3548 a_10219_943.n16 a_10219_943.n15 30
R3549 a_10219_943.n14 a_10219_943.n11 26.552
R3550 a_10219_943.n17 a_10219_943.n0 24.383
R3551 a_10219_943.n17 a_10219_943.n16 23.684
R3552 a_10219_943.n5 a_10219_943.n1 16.08
R3553 a_10219_943.n4 a_10219_943.n2 16.08
R3554 a_10219_943.n1 a_10219_943.t3 14.282
R3555 a_10219_943.n1 a_10219_943.t4 14.282
R3556 a_10219_943.n2 a_10219_943.t0 14.282
R3557 a_10219_943.n2 a_10219_943.t1 14.282
R3558 a_10219_943.n3 a_10219_943.t5 14.282
R3559 a_10219_943.n3 a_10219_943.t6 14.282
R3560 a_17708_181.n4 a_17708_181.t7 512.525
R3561 a_17708_181.n4 a_17708_181.t9 371.139
R3562 a_17708_181.n5 a_17708_181.t8 273.368
R3563 a_17708_181.n10 a_17708_181.n6 226.775
R3564 a_17708_181.n6 a_17708_181.n5 153.043
R3565 a_17708_181.n6 a_17708_181.n3 110.158
R3566 a_17708_181.n5 a_17708_181.n4 105.194
R3567 a_17708_181.n17 a_17708_181.n15 103.718
R3568 a_17708_181.n15 a_17708_181.n14 98.501
R3569 a_17708_181.n9 a_17708_181.n7 80.526
R3570 a_17708_181.n15 a_17708_181.n10 78.403
R3571 a_17708_181.n3 a_17708_181.n2 75.271
R3572 a_17708_181.n14 a_17708_181.n13 30
R3573 a_17708_181.n9 a_17708_181.n8 30
R3574 a_17708_181.n12 a_17708_181.n11 24.383
R3575 a_17708_181.n18 a_17708_181.n0 24.383
R3576 a_17708_181.n14 a_17708_181.n12 23.684
R3577 a_17708_181.n10 a_17708_181.n9 20.417
R3578 a_17708_181.n1 a_17708_181.t2 14.282
R3579 a_17708_181.n1 a_17708_181.t3 14.282
R3580 a_17708_181.n2 a_17708_181.t6 14.282
R3581 a_17708_181.n2 a_17708_181.t0 14.282
R3582 a_17708_181.n17 a_17708_181.n16 13.452
R3583 a_17708_181.n3 a_17708_181.n1 12.119
R3584 a_17708_181.n18 a_17708_181.n17 10.62
R3585 a_18197_1005.n4 a_18197_1005.n3 196.002
R3586 a_18197_1005.t3 a_18197_1005.n5 89.556
R3587 a_18197_1005.n3 a_18197_1005.n2 75.271
R3588 a_18197_1005.n5 a_18197_1005.n4 75.214
R3589 a_18197_1005.n3 a_18197_1005.n1 36.52
R3590 a_18197_1005.n4 a_18197_1005.t0 14.338
R3591 a_18197_1005.n1 a_18197_1005.t1 14.282
R3592 a_18197_1005.n1 a_18197_1005.t7 14.282
R3593 a_18197_1005.n2 a_18197_1005.t5 14.282
R3594 a_18197_1005.n2 a_18197_1005.t6 14.282
R3595 a_18197_1005.n0 a_18197_1005.t2 14.282
R3596 a_18197_1005.n0 a_18197_1005.t4 14.282
R3597 a_18197_1005.n5 a_18197_1005.n0 12.119
R3598 a_17533_1005.n4 a_17533_1005.n3 195.987
R3599 a_17533_1005.n2 a_17533_1005.t0 89.553
R3600 a_17533_1005.n4 a_17533_1005.n0 75.271
R3601 a_17533_1005.n3 a_17533_1005.n2 75.214
R3602 a_17533_1005.n5 a_17533_1005.n4 36.517
R3603 a_17533_1005.n3 a_17533_1005.t6 14.338
R3604 a_17533_1005.n1 a_17533_1005.t7 14.282
R3605 a_17533_1005.n1 a_17533_1005.t5 14.282
R3606 a_17533_1005.n0 a_17533_1005.t4 14.282
R3607 a_17533_1005.n0 a_17533_1005.t3 14.282
R3608 a_17533_1005.n5 a_17533_1005.t1 14.282
R3609 a_17533_1005.t2 a_17533_1005.n5 14.282
R3610 a_17533_1005.n2 a_17533_1005.n1 12.119
R3611 a_14521_75.n4 a_14521_75.n3 19.724
R3612 a_14521_75.t0 a_14521_75.n5 11.595
R3613 a_14521_75.t0 a_14521_75.n4 9.207
R3614 a_14521_75.n2 a_14521_75.n0 8.543
R3615 a_14521_75.t0 a_14521_75.n2 3.034
R3616 a_14521_75.n2 a_14521_75.n1 0.443
R3617 a_14802_182.n12 a_14802_182.n5 96.467
R3618 a_14802_182.t0 a_14802_182.n1 46.91
R3619 a_14802_182.n9 a_14802_182.n7 34.805
R3620 a_14802_182.n9 a_14802_182.n8 32.622
R3621 a_14802_182.t0 a_14802_182.n12 32.417
R3622 a_14802_182.n5 a_14802_182.n4 22.349
R3623 a_14802_182.n11 a_14802_182.n9 19.017
R3624 a_14802_182.n1 a_14802_182.n0 17.006
R3625 a_14802_182.n5 a_14802_182.n3 8.443
R3626 a_14802_182.t0 a_14802_182.n2 8.137
R3627 a_14802_182.n7 a_14802_182.n6 7.5
R3628 a_14802_182.n11 a_14802_182.n10 7.5
R3629 a_14802_182.n12 a_14802_182.n11 1.435
R3630 a_277_1004.n7 a_277_1004.t10 512.525
R3631 a_277_1004.n5 a_277_1004.t7 512.525
R3632 a_277_1004.n7 a_277_1004.t11 371.139
R3633 a_277_1004.n5 a_277_1004.t12 371.139
R3634 a_277_1004.n10 a_277_1004.n4 233.952
R3635 a_277_1004.n8 a_277_1004.n7 225.866
R3636 a_277_1004.n6 a_277_1004.n5 225.866
R3637 a_277_1004.n8 a_277_1004.t9 218.057
R3638 a_277_1004.n6 a_277_1004.t8 218.057
R3639 a_277_1004.n12 a_277_1004.n10 150.014
R3640 a_277_1004.n9 a_277_1004.n6 79.491
R3641 a_277_1004.n3 a_277_1004.n2 79.232
R3642 a_277_1004.n10 a_277_1004.n9 77.315
R3643 a_277_1004.n9 a_277_1004.n8 76
R3644 a_277_1004.n4 a_277_1004.n3 63.152
R3645 a_277_1004.n4 a_277_1004.n0 16.08
R3646 a_277_1004.n3 a_277_1004.n1 16.08
R3647 a_277_1004.n12 a_277_1004.n11 15.218
R3648 a_277_1004.n0 a_277_1004.t4 14.282
R3649 a_277_1004.n0 a_277_1004.t0 14.282
R3650 a_277_1004.n1 a_277_1004.t6 14.282
R3651 a_277_1004.n1 a_277_1004.t5 14.282
R3652 a_277_1004.n2 a_277_1004.t2 14.282
R3653 a_277_1004.n2 a_277_1004.t1 14.282
R3654 a_277_1004.n13 a_277_1004.n12 12.014
R3655 a_11821_1004.n8 a_11821_1004.t10 512.525
R3656 a_11821_1004.n6 a_11821_1004.t8 512.525
R3657 a_11821_1004.n8 a_11821_1004.t7 371.139
R3658 a_11821_1004.n6 a_11821_1004.t11 371.139
R3659 a_11821_1004.n11 a_11821_1004.n5 233.952
R3660 a_11821_1004.n9 a_11821_1004.n8 225.866
R3661 a_11821_1004.n7 a_11821_1004.n6 225.866
R3662 a_11821_1004.n9 a_11821_1004.t9 218.057
R3663 a_11821_1004.n7 a_11821_1004.t12 218.057
R3664 a_11821_1004.n13 a_11821_1004.n11 143.492
R3665 a_11821_1004.n10 a_11821_1004.n7 79.491
R3666 a_11821_1004.n4 a_11821_1004.n3 79.232
R3667 a_11821_1004.n11 a_11821_1004.n10 77.315
R3668 a_11821_1004.n10 a_11821_1004.n9 76
R3669 a_11821_1004.n5 a_11821_1004.n4 63.152
R3670 a_11821_1004.n13 a_11821_1004.n12 30
R3671 a_11821_1004.n14 a_11821_1004.n0 24.383
R3672 a_11821_1004.n14 a_11821_1004.n13 23.684
R3673 a_11821_1004.n5 a_11821_1004.n1 16.08
R3674 a_11821_1004.n4 a_11821_1004.n2 16.08
R3675 a_11821_1004.n1 a_11821_1004.t4 14.282
R3676 a_11821_1004.n1 a_11821_1004.t5 14.282
R3677 a_11821_1004.n2 a_11821_1004.t3 14.282
R3678 a_11821_1004.n2 a_11821_1004.t2 14.282
R3679 a_11821_1004.n3 a_11821_1004.t1 14.282
R3680 a_11821_1004.n3 a_11821_1004.t0 14.282
R3681 a_15991_943.n8 a_15991_943.t8 512.525
R3682 a_15991_943.n6 a_15991_943.t9 512.525
R3683 a_15991_943.n11 a_15991_943.t13 454.685
R3684 a_15991_943.n11 a_15991_943.t10 428.979
R3685 a_15991_943.n8 a_15991_943.t15 371.139
R3686 a_15991_943.n6 a_15991_943.t14 371.139
R3687 a_15991_943.n14 a_15991_943.n5 260.505
R3688 a_15991_943.n9 a_15991_943.n8 258.98
R3689 a_15991_943.n7 a_15991_943.n6 258.98
R3690 a_15991_943.n12 a_15991_943.n11 189.419
R3691 a_15991_943.n7 a_15991_943.t12 176.995
R3692 a_15991_943.n9 a_15991_943.t7 170.569
R3693 a_15991_943.n12 a_15991_943.t11 126.558
R3694 a_15991_943.n16 a_15991_943.n14 116.939
R3695 a_15991_943.n4 a_15991_943.n3 79.232
R3696 a_15991_943.n10 a_15991_943.n7 77.027
R3697 a_15991_943.n10 a_15991_943.n9 76
R3698 a_15991_943.n14 a_15991_943.n13 76
R3699 a_15991_943.n5 a_15991_943.n4 63.152
R3700 a_15991_943.n13 a_15991_943.n12 53.379
R3701 a_15991_943.n16 a_15991_943.n15 30
R3702 a_15991_943.n17 a_15991_943.n0 24.383
R3703 a_15991_943.n17 a_15991_943.n16 23.684
R3704 a_15991_943.n5 a_15991_943.n1 16.08
R3705 a_15991_943.n4 a_15991_943.n2 16.08
R3706 a_15991_943.n1 a_15991_943.t5 14.282
R3707 a_15991_943.n1 a_15991_943.t6 14.282
R3708 a_15991_943.n2 a_15991_943.t2 14.282
R3709 a_15991_943.n2 a_15991_943.t3 14.282
R3710 a_15991_943.n3 a_15991_943.t1 14.282
R3711 a_15991_943.n3 a_15991_943.t0 14.282
R3712 a_15991_943.n13 a_15991_943.n10 4.825
R3713 a_18094_73.n2 a_18094_73.n0 34.602
R3714 a_18094_73.n2 a_18094_73.n1 2.138
R3715 a_18094_73.t0 a_18094_73.n2 0.069
R3716 a_16445_75.n4 a_16445_75.n3 19.724
R3717 a_16445_75.t0 a_16445_75.n5 11.595
R3718 a_16445_75.t0 a_16445_75.n4 9.207
R3719 a_16445_75.n2 a_16445_75.n0 8.543
R3720 a_16445_75.t0 a_16445_75.n2 3.034
R3721 a_16445_75.n2 a_16445_75.n1 0.443
R3722 a_16726_182.n10 a_16726_182.n8 82.852
R3723 a_16726_182.n11 a_16726_182.n0 49.6
R3724 a_16726_182.n7 a_16726_182.n6 32.833
R3725 a_16726_182.n8 a_16726_182.t1 32.416
R3726 a_16726_182.n10 a_16726_182.n9 27.2
R3727 a_16726_182.n3 a_16726_182.n2 23.284
R3728 a_16726_182.n11 a_16726_182.n10 22.4
R3729 a_16726_182.n7 a_16726_182.n4 19.017
R3730 a_16726_182.n6 a_16726_182.n5 13.494
R3731 a_16726_182.t1 a_16726_182.n1 7.04
R3732 a_16726_182.t1 a_16726_182.n3 5.727
R3733 a_16726_182.n8 a_16726_182.n7 1.435
R3734 a_10673_75.n4 a_10673_75.n3 19.724
R3735 a_10673_75.t0 a_10673_75.n5 11.595
R3736 a_10673_75.t0 a_10673_75.n4 9.207
R3737 a_10673_75.n2 a_10673_75.n0 8.543
R3738 a_10673_75.t0 a_10673_75.n2 3.034
R3739 a_10673_75.n2 a_10673_75.n1 0.443
R3740 a_10954_182.n10 a_10954_182.n8 82.852
R3741 a_10954_182.n11 a_10954_182.n0 49.6
R3742 a_10954_182.n7 a_10954_182.n6 32.833
R3743 a_10954_182.n8 a_10954_182.t1 32.416
R3744 a_10954_182.n10 a_10954_182.n9 27.2
R3745 a_10954_182.n3 a_10954_182.n2 23.284
R3746 a_10954_182.n11 a_10954_182.n10 22.4
R3747 a_10954_182.n7 a_10954_182.n4 19.017
R3748 a_10954_182.n6 a_10954_182.n5 13.494
R3749 a_10954_182.t1 a_10954_182.n1 7.04
R3750 a_10954_182.t1 a_10954_182.n3 5.727
R3751 a_10954_182.n8 a_10954_182.n7 1.435
R3752 a_12597_75.n1 a_12597_75.n0 25.576
R3753 a_12597_75.n3 a_12597_75.n2 9.111
R3754 a_12597_75.n7 a_12597_75.n5 7.859
R3755 a_12597_75.t0 a_12597_75.n7 3.034
R3756 a_12597_75.n5 a_12597_75.n3 1.964
R3757 a_12597_75.n5 a_12597_75.n4 1.964
R3758 a_12597_75.t0 a_12597_75.n1 1.871
R3759 a_12597_75.n7 a_12597_75.n6 0.443
R3760 a_12878_182.n8 a_12878_182.n6 96.467
R3761 a_12878_182.n3 a_12878_182.n1 44.628
R3762 a_12878_182.t0 a_12878_182.n8 32.417
R3763 a_12878_182.n3 a_12878_182.n2 23.284
R3764 a_12878_182.n6 a_12878_182.n5 22.349
R3765 a_12878_182.t0 a_12878_182.n10 20.241
R3766 a_12878_182.n10 a_12878_182.n9 13.494
R3767 a_12878_182.n6 a_12878_182.n4 8.443
R3768 a_12878_182.t0 a_12878_182.n0 8.137
R3769 a_12878_182.t0 a_12878_182.n3 5.727
R3770 a_12878_182.n8 a_12878_182.n7 1.435
R3771 a_15669_1004.n6 a_15669_1004.t9 512.525
R3772 a_15669_1004.n6 a_15669_1004.t8 371.139
R3773 a_15669_1004.n8 a_15669_1004.n5 233.952
R3774 a_15669_1004.n7 a_15669_1004.n6 225.866
R3775 a_15669_1004.n7 a_15669_1004.t7 218.057
R3776 a_15669_1004.n8 a_15669_1004.n7 153.315
R3777 a_15669_1004.n10 a_15669_1004.n8 143.492
R3778 a_15669_1004.n4 a_15669_1004.n3 79.232
R3779 a_15669_1004.n5 a_15669_1004.n4 63.152
R3780 a_15669_1004.n10 a_15669_1004.n9 30
R3781 a_15669_1004.n11 a_15669_1004.n0 24.383
R3782 a_15669_1004.n11 a_15669_1004.n10 23.684
R3783 a_15669_1004.n5 a_15669_1004.n1 16.08
R3784 a_15669_1004.n4 a_15669_1004.n2 16.08
R3785 a_15669_1004.n1 a_15669_1004.t1 14.282
R3786 a_15669_1004.n1 a_15669_1004.t0 14.282
R3787 a_15669_1004.n2 a_15669_1004.t4 14.282
R3788 a_15669_1004.n2 a_15669_1004.t3 14.282
R3789 a_15669_1004.n3 a_15669_1004.t5 14.282
R3790 a_15669_1004.n3 a_15669_1004.t6 14.282
R3791 a_599_943.n5 a_599_943.t12 512.525
R3792 a_599_943.n7 a_599_943.t10 454.685
R3793 a_599_943.n7 a_599_943.t8 428.979
R3794 a_599_943.n5 a_599_943.t7 371.139
R3795 a_599_943.n6 a_599_943.t9 271.162
R3796 a_599_943.n8 a_599_943.t11 221.453
R3797 a_599_943.n12 a_599_943.n10 203.12
R3798 a_599_943.n10 a_599_943.n4 180.846
R3799 a_599_943.n6 a_599_943.n5 172.76
R3800 a_599_943.n8 a_599_943.n7 108.494
R3801 a_599_943.n9 a_599_943.n6 84.388
R3802 a_599_943.n9 a_599_943.n8 80.035
R3803 a_599_943.n3 a_599_943.n2 79.232
R3804 a_599_943.n10 a_599_943.n9 76
R3805 a_599_943.n4 a_599_943.n3 63.152
R3806 a_599_943.n4 a_599_943.n0 16.08
R3807 a_599_943.n3 a_599_943.n1 16.08
R3808 a_599_943.n12 a_599_943.n11 15.218
R3809 a_599_943.n0 a_599_943.t0 14.282
R3810 a_599_943.n0 a_599_943.t6 14.282
R3811 a_599_943.n1 a_599_943.t2 14.282
R3812 a_599_943.n1 a_599_943.t3 14.282
R3813 a_599_943.n2 a_599_943.t5 14.282
R3814 a_599_943.n2 a_599_943.t4 14.282
R3815 a_599_943.n13 a_599_943.n12 12.014
R3816 a_9897_1004.n6 a_9897_1004.t7 512.525
R3817 a_9897_1004.n6 a_9897_1004.t8 371.139
R3818 a_9897_1004.n8 a_9897_1004.n5 233.952
R3819 a_9897_1004.n7 a_9897_1004.n6 225.866
R3820 a_9897_1004.n7 a_9897_1004.t9 218.057
R3821 a_9897_1004.n8 a_9897_1004.n7 153.315
R3822 a_9897_1004.n10 a_9897_1004.n8 143.492
R3823 a_9897_1004.n4 a_9897_1004.n3 79.232
R3824 a_9897_1004.n5 a_9897_1004.n4 63.152
R3825 a_9897_1004.n10 a_9897_1004.n9 30
R3826 a_9897_1004.n11 a_9897_1004.n0 24.383
R3827 a_9897_1004.n11 a_9897_1004.n10 23.684
R3828 a_9897_1004.n5 a_9897_1004.n1 16.08
R3829 a_9897_1004.n4 a_9897_1004.n2 16.08
R3830 a_9897_1004.n1 a_9897_1004.t0 14.282
R3831 a_9897_1004.n1 a_9897_1004.t1 14.282
R3832 a_9897_1004.n2 a_9897_1004.t4 14.282
R3833 a_9897_1004.n2 a_9897_1004.t3 14.282
R3834 a_9897_1004.n3 a_9897_1004.t5 14.282
R3835 a_9897_1004.n3 a_9897_1004.t6 14.282
R3836 a_1561_943.n8 a_1561_943.t14 454.685
R3837 a_1561_943.n10 a_1561_943.t8 454.685
R3838 a_1561_943.n6 a_1561_943.t15 454.685
R3839 a_1561_943.n8 a_1561_943.t11 428.979
R3840 a_1561_943.n10 a_1561_943.t12 428.979
R3841 a_1561_943.n6 a_1561_943.t13 428.979
R3842 a_1561_943.n9 a_1561_943.t7 248.006
R3843 a_1561_943.n11 a_1561_943.t9 248.006
R3844 a_1561_943.n7 a_1561_943.t10 248.006
R3845 a_1561_943.n16 a_1561_943.n14 223.151
R3846 a_1561_943.n14 a_1561_943.n5 154.293
R3847 a_1561_943.n13 a_1561_943.n7 82.484
R3848 a_1561_943.n9 a_1561_943.n8 81.941
R3849 a_1561_943.n11 a_1561_943.n10 81.941
R3850 a_1561_943.n7 a_1561_943.n6 81.941
R3851 a_1561_943.n12 a_1561_943.n11 79.491
R3852 a_1561_943.n4 a_1561_943.n3 79.232
R3853 a_1561_943.n12 a_1561_943.n9 76
R3854 a_1561_943.n14 a_1561_943.n13 76
R3855 a_1561_943.n5 a_1561_943.n4 63.152
R3856 a_1561_943.n16 a_1561_943.n15 30
R3857 a_1561_943.n17 a_1561_943.n0 24.383
R3858 a_1561_943.n17 a_1561_943.n16 23.684
R3859 a_1561_943.n5 a_1561_943.n1 16.08
R3860 a_1561_943.n4 a_1561_943.n2 16.08
R3861 a_1561_943.n1 a_1561_943.t2 14.282
R3862 a_1561_943.n1 a_1561_943.t1 14.282
R3863 a_1561_943.n2 a_1561_943.t5 14.282
R3864 a_1561_943.n2 a_1561_943.t4 14.282
R3865 a_1561_943.n3 a_1561_943.t6 14.282
R3866 a_1561_943.n3 a_1561_943.t0 14.282
R3867 a_1561_943.n13 a_1561_943.n12 4.035
R3868 a_2296_182.n13 a_2296_182.n6 82.852
R3869 a_2296_182.t0 a_2296_182.n1 46.91
R3870 a_2296_182.n10 a_2296_182.n8 34.805
R3871 a_2296_182.n10 a_2296_182.n9 32.622
R3872 a_2296_182.t0 a_2296_182.n13 32.417
R3873 a_2296_182.n6 a_2296_182.n5 27.2
R3874 a_2296_182.n4 a_2296_182.n3 23.498
R3875 a_2296_182.n6 a_2296_182.n4 22.4
R3876 a_2296_182.n12 a_2296_182.n10 19.017
R3877 a_2296_182.n1 a_2296_182.n0 17.006
R3878 a_2296_182.t0 a_2296_182.n2 8.137
R3879 a_2296_182.n8 a_2296_182.n7 7.5
R3880 a_2296_182.n12 a_2296_182.n11 7.5
R3881 a_2296_182.n13 a_2296_182.n12 1.435
R3882 a_2201_1004.n5 a_2201_1004.t9 512.525
R3883 a_2201_1004.n5 a_2201_1004.t8 371.139
R3884 a_2201_1004.n7 a_2201_1004.n4 233.952
R3885 a_2201_1004.n6 a_2201_1004.n5 225.866
R3886 a_2201_1004.n6 a_2201_1004.t7 218.057
R3887 a_2201_1004.n7 a_2201_1004.n6 153.315
R3888 a_2201_1004.n9 a_2201_1004.n7 150.014
R3889 a_2201_1004.n3 a_2201_1004.n2 79.232
R3890 a_2201_1004.n4 a_2201_1004.n3 63.152
R3891 a_2201_1004.n4 a_2201_1004.n0 16.08
R3892 a_2201_1004.n3 a_2201_1004.n1 16.08
R3893 a_2201_1004.n9 a_2201_1004.n8 15.218
R3894 a_2201_1004.n0 a_2201_1004.t1 14.282
R3895 a_2201_1004.n0 a_2201_1004.t0 14.282
R3896 a_2201_1004.n1 a_2201_1004.t4 14.282
R3897 a_2201_1004.n1 a_2201_1004.t3 14.282
R3898 a_2201_1004.n2 a_2201_1004.t6 14.282
R3899 a_2201_1004.n2 a_2201_1004.t5 14.282
R3900 a_2201_1004.n10 a_2201_1004.n9 12.014
R3901 a_91_75.n4 a_91_75.n3 19.724
R3902 a_91_75.t0 a_91_75.n5 11.595
R3903 a_91_75.t0 a_91_75.n4 9.207
R3904 a_91_75.n2 a_91_75.n0 8.543
R3905 a_91_75.t0 a_91_75.n2 3.034
R3906 a_91_75.n2 a_91_75.n1 0.443
R3907 a_372_182.n10 a_372_182.n8 82.852
R3908 a_372_182.n11 a_372_182.n0 49.6
R3909 a_372_182.n7 a_372_182.n6 32.833
R3910 a_372_182.n8 a_372_182.t1 32.416
R3911 a_372_182.n10 a_372_182.n9 27.2
R3912 a_372_182.n3 a_372_182.n2 23.284
R3913 a_372_182.n11 a_372_182.n10 22.4
R3914 a_372_182.n7 a_372_182.n4 19.017
R3915 a_372_182.n6 a_372_182.n5 13.494
R3916 a_372_182.t1 a_372_182.n1 7.04
R3917 a_372_182.t1 a_372_182.n3 5.727
R3918 a_372_182.n8 a_372_182.n7 1.435
R3919 a_13105_943.n7 a_13105_943.t12 454.685
R3920 a_13105_943.n9 a_13105_943.t14 454.685
R3921 a_13105_943.n5 a_13105_943.t10 454.685
R3922 a_13105_943.n7 a_13105_943.t7 428.979
R3923 a_13105_943.n9 a_13105_943.t11 428.979
R3924 a_13105_943.n5 a_13105_943.t8 428.979
R3925 a_13105_943.n8 a_13105_943.t13 248.006
R3926 a_13105_943.n10 a_13105_943.t9 248.006
R3927 a_13105_943.n6 a_13105_943.t15 248.006
R3928 a_13105_943.n15 a_13105_943.n13 229.673
R3929 a_13105_943.n13 a_13105_943.n4 154.293
R3930 a_13105_943.n12 a_13105_943.n6 82.484
R3931 a_13105_943.n8 a_13105_943.n7 81.941
R3932 a_13105_943.n10 a_13105_943.n9 81.941
R3933 a_13105_943.n6 a_13105_943.n5 81.941
R3934 a_13105_943.n11 a_13105_943.n10 79.491
R3935 a_13105_943.n3 a_13105_943.n2 79.232
R3936 a_13105_943.n11 a_13105_943.n8 76
R3937 a_13105_943.n13 a_13105_943.n12 76
R3938 a_13105_943.n4 a_13105_943.n3 63.152
R3939 a_13105_943.n4 a_13105_943.n0 16.08
R3940 a_13105_943.n3 a_13105_943.n1 16.08
R3941 a_13105_943.n15 a_13105_943.n14 15.218
R3942 a_13105_943.n0 a_13105_943.t2 14.282
R3943 a_13105_943.n0 a_13105_943.t3 14.282
R3944 a_13105_943.n1 a_13105_943.t6 14.282
R3945 a_13105_943.n1 a_13105_943.t5 14.282
R3946 a_13105_943.n2 a_13105_943.t1 14.282
R3947 a_13105_943.n2 a_13105_943.t0 14.282
R3948 a_13105_943.n16 a_13105_943.n15 12.014
R3949 a_13105_943.n12 a_13105_943.n11 4.035
R3950 a_13745_1004.n6 a_13745_1004.t7 512.525
R3951 a_13745_1004.n6 a_13745_1004.t8 371.139
R3952 a_13745_1004.n8 a_13745_1004.n5 233.952
R3953 a_13745_1004.n7 a_13745_1004.n6 225.866
R3954 a_13745_1004.n7 a_13745_1004.t9 218.057
R3955 a_13745_1004.n8 a_13745_1004.n7 153.315
R3956 a_13745_1004.n10 a_13745_1004.n8 143.492
R3957 a_13745_1004.n4 a_13745_1004.n3 79.232
R3958 a_13745_1004.n5 a_13745_1004.n4 63.152
R3959 a_13745_1004.n10 a_13745_1004.n9 30
R3960 a_13745_1004.n11 a_13745_1004.n0 24.383
R3961 a_13745_1004.n11 a_13745_1004.n10 23.684
R3962 a_13745_1004.n5 a_13745_1004.n1 16.08
R3963 a_13745_1004.n4 a_13745_1004.n2 16.08
R3964 a_13745_1004.n1 a_13745_1004.t1 14.282
R3965 a_13745_1004.n1 a_13745_1004.t0 14.282
R3966 a_13745_1004.n2 a_13745_1004.t3 14.282
R3967 a_13745_1004.n2 a_13745_1004.t4 14.282
R3968 a_13745_1004.n3 a_13745_1004.t6 14.282
R3969 a_13745_1004.n3 a_13745_1004.t5 14.282
R3970 a_4220_182.n12 a_4220_182.n10 82.852
R3971 a_4220_182.t1 a_4220_182.n2 46.91
R3972 a_4220_182.n7 a_4220_182.n5 34.805
R3973 a_4220_182.n7 a_4220_182.n6 32.622
R3974 a_4220_182.n10 a_4220_182.t1 32.416
R3975 a_4220_182.n12 a_4220_182.n11 27.2
R3976 a_4220_182.n13 a_4220_182.n0 23.498
R3977 a_4220_182.n13 a_4220_182.n12 22.4
R3978 a_4220_182.n9 a_4220_182.n7 19.017
R3979 a_4220_182.n2 a_4220_182.n1 17.006
R3980 a_4220_182.n5 a_4220_182.n4 7.5
R3981 a_4220_182.n9 a_4220_182.n8 7.5
R3982 a_4220_182.t1 a_4220_182.n3 7.04
R3983 a_4220_182.n10 a_4220_182.n9 1.435
R3984 a_4125_1004.n5 a_4125_1004.t7 512.525
R3985 a_4125_1004.n5 a_4125_1004.t9 371.139
R3986 a_4125_1004.n7 a_4125_1004.n4 233.952
R3987 a_4125_1004.n6 a_4125_1004.n5 225.866
R3988 a_4125_1004.n6 a_4125_1004.t8 218.057
R3989 a_4125_1004.n7 a_4125_1004.n6 153.315
R3990 a_4125_1004.n9 a_4125_1004.n7 150.014
R3991 a_4125_1004.n3 a_4125_1004.n2 79.232
R3992 a_4125_1004.n4 a_4125_1004.n3 63.152
R3993 a_4125_1004.n4 a_4125_1004.n0 16.08
R3994 a_4125_1004.n3 a_4125_1004.n1 16.08
R3995 a_4125_1004.n9 a_4125_1004.n8 15.218
R3996 a_4125_1004.n0 a_4125_1004.t4 14.282
R3997 a_4125_1004.n0 a_4125_1004.t5 14.282
R3998 a_4125_1004.n1 a_4125_1004.t0 14.282
R3999 a_4125_1004.n1 a_4125_1004.t1 14.282
R4000 a_4125_1004.n2 a_4125_1004.t2 14.282
R4001 a_4125_1004.n2 a_4125_1004.t3 14.282
R4002 a_4125_1004.n10 a_4125_1004.n9 12.014
R4003 Q.n2 Q.n1 263.549
R4004 Q.n2 Q.n0 114.038
R4005 Q.n3 Q.n2 76
R4006 Q.n0 Q.t1 14.282
R4007 Q.n0 Q.t0 14.282
R4008 Q.n3 Q 0.046
R4009 a_13559_75.n1 a_13559_75.n0 25.576
R4010 a_13559_75.n3 a_13559_75.n2 9.111
R4011 a_13559_75.n7 a_13559_75.n5 7.859
R4012 a_13559_75.t0 a_13559_75.n7 3.034
R4013 a_13559_75.n5 a_13559_75.n3 1.964
R4014 a_13559_75.n5 a_13559_75.n4 1.964
R4015 a_13559_75.t0 a_13559_75.n1 1.871
R4016 a_13559_75.n7 a_13559_75.n6 0.443
R4017 a_13840_182.n8 a_13840_182.n6 96.467
R4018 a_13840_182.n3 a_13840_182.n1 44.628
R4019 a_13840_182.t0 a_13840_182.n8 32.417
R4020 a_13840_182.n3 a_13840_182.n2 23.284
R4021 a_13840_182.n6 a_13840_182.n5 22.349
R4022 a_13840_182.t0 a_13840_182.n10 20.241
R4023 a_13840_182.n10 a_13840_182.n9 13.494
R4024 a_13840_182.n6 a_13840_182.n4 8.443
R4025 a_13840_182.t0 a_13840_182.n0 8.137
R4026 a_13840_182.t0 a_13840_182.n3 5.727
R4027 a_13840_182.n8 a_13840_182.n7 1.435
R4028 a_15764_182.n8 a_15764_182.n6 96.467
R4029 a_15764_182.n3 a_15764_182.n1 44.628
R4030 a_15764_182.t0 a_15764_182.n8 32.417
R4031 a_15764_182.n3 a_15764_182.n2 23.284
R4032 a_15764_182.n6 a_15764_182.n5 22.349
R4033 a_15764_182.t0 a_15764_182.n10 20.241
R4034 a_15764_182.n10 a_15764_182.n9 13.494
R4035 a_15764_182.n6 a_15764_182.n4 8.443
R4036 a_15764_182.t0 a_15764_182.n0 8.137
R4037 a_15764_182.t0 a_15764_182.n3 5.727
R4038 a_15764_182.n8 a_15764_182.n7 1.435
R4039 a_7106_182.n10 a_7106_182.n8 82.852
R4040 a_7106_182.n7 a_7106_182.n6 32.833
R4041 a_7106_182.n8 a_7106_182.t1 32.416
R4042 a_7106_182.n10 a_7106_182.n9 27.2
R4043 a_7106_182.n11 a_7106_182.n0 23.498
R4044 a_7106_182.n3 a_7106_182.n2 23.284
R4045 a_7106_182.n11 a_7106_182.n10 22.4
R4046 a_7106_182.n7 a_7106_182.n4 19.017
R4047 a_7106_182.n6 a_7106_182.n5 13.494
R4048 a_7106_182.t1 a_7106_182.n1 7.04
R4049 a_7106_182.t1 a_7106_182.n3 5.727
R4050 a_7106_182.n8 a_7106_182.n7 1.435
R4051 a_2015_75.n1 a_2015_75.n0 25.576
R4052 a_2015_75.n3 a_2015_75.n2 9.111
R4053 a_2015_75.n7 a_2015_75.n6 2.455
R4054 a_2015_75.n5 a_2015_75.n3 1.964
R4055 a_2015_75.n5 a_2015_75.n4 1.964
R4056 a_2015_75.t0 a_2015_75.n1 1.871
R4057 a_2015_75.n7 a_2015_75.n5 0.636
R4058 a_2015_75.t0 a_2015_75.n7 0.246
R4059 a_1334_182.n9 a_1334_182.n7 82.852
R4060 a_1334_182.n3 a_1334_182.n1 44.628
R4061 a_1334_182.t0 a_1334_182.n9 32.417
R4062 a_1334_182.n7 a_1334_182.n6 27.2
R4063 a_1334_182.n5 a_1334_182.n4 23.498
R4064 a_1334_182.n3 a_1334_182.n2 23.284
R4065 a_1334_182.n7 a_1334_182.n5 22.4
R4066 a_1334_182.t0 a_1334_182.n11 20.241
R4067 a_1334_182.n11 a_1334_182.n10 13.494
R4068 a_1334_182.t0 a_1334_182.n0 8.137
R4069 a_1334_182.t0 a_1334_182.n3 5.727
R4070 a_1334_182.n9 a_1334_182.n8 1.435
R4071 a_3258_182.n9 a_3258_182.n7 82.852
R4072 a_3258_182.n3 a_3258_182.n1 44.628
R4073 a_3258_182.t0 a_3258_182.n9 32.417
R4074 a_3258_182.n7 a_3258_182.n6 27.2
R4075 a_3258_182.n5 a_3258_182.n4 23.498
R4076 a_3258_182.n3 a_3258_182.n2 23.284
R4077 a_3258_182.n7 a_3258_182.n5 22.4
R4078 a_3258_182.t0 a_3258_182.n11 20.241
R4079 a_3258_182.n11 a_3258_182.n10 13.494
R4080 a_3258_182.t0 a_3258_182.n0 8.137
R4081 a_3258_182.t0 a_3258_182.n3 5.727
R4082 a_3258_182.n9 a_3258_182.n8 1.435
R4083 a_5182_182.n9 a_5182_182.n7 82.852
R4084 a_5182_182.n3 a_5182_182.n1 44.628
R4085 a_5182_182.t0 a_5182_182.n9 32.417
R4086 a_5182_182.n7 a_5182_182.n6 27.2
R4087 a_5182_182.n5 a_5182_182.n4 23.498
R4088 a_5182_182.n3 a_5182_182.n2 23.284
R4089 a_5182_182.n7 a_5182_182.n5 22.4
R4090 a_5182_182.t0 a_5182_182.n11 20.241
R4091 a_5182_182.n11 a_5182_182.n10 13.494
R4092 a_5182_182.t0 a_5182_182.n0 8.137
R4093 a_5182_182.t0 a_5182_182.n3 5.727
R4094 a_5182_182.n9 a_5182_182.n8 1.435
R4095 a_11916_182.n10 a_11916_182.n8 82.852
R4096 a_11916_182.n7 a_11916_182.n6 32.833
R4097 a_11916_182.n8 a_11916_182.t1 32.416
R4098 a_11916_182.n10 a_11916_182.n9 27.2
R4099 a_11916_182.n11 a_11916_182.n0 23.498
R4100 a_11916_182.n3 a_11916_182.n2 23.284
R4101 a_11916_182.n11 a_11916_182.n10 22.4
R4102 a_11916_182.n7 a_11916_182.n4 19.017
R4103 a_11916_182.n6 a_11916_182.n5 13.494
R4104 a_11916_182.t1 a_11916_182.n1 7.04
R4105 a_11916_182.t1 a_11916_182.n3 5.727
R4106 a_11916_182.n8 a_11916_182.n7 1.435
R4107 a_17428_73.n1 a_17428_73.n0 32.249
R4108 a_17428_73.t0 a_17428_73.n5 7.911
R4109 a_17428_73.n4 a_17428_73.n2 4.032
R4110 a_17428_73.n4 a_17428_73.n3 3.644
R4111 a_17428_73.t0 a_17428_73.n1 2.534
R4112 a_17428_73.t0 a_17428_73.n4 1.099
R4113 a_9992_182.n9 a_9992_182.n7 82.852
R4114 a_9992_182.n3 a_9992_182.n1 44.628
R4115 a_9992_182.t0 a_9992_182.n9 32.417
R4116 a_9992_182.n7 a_9992_182.n6 27.2
R4117 a_9992_182.n5 a_9992_182.n4 23.498
R4118 a_9992_182.n3 a_9992_182.n2 23.284
R4119 a_9992_182.n7 a_9992_182.n5 22.4
R4120 a_9992_182.t0 a_9992_182.n11 20.241
R4121 a_9992_182.n11 a_9992_182.n10 13.494
R4122 a_9992_182.t0 a_9992_182.n0 8.137
R4123 a_9992_182.t0 a_9992_182.n3 5.727
R4124 a_9992_182.n9 a_9992_182.n8 1.435
R4125 a_6144_182.n10 a_6144_182.n8 82.852
R4126 a_6144_182.n7 a_6144_182.n6 32.833
R4127 a_6144_182.n8 a_6144_182.t1 32.416
R4128 a_6144_182.n10 a_6144_182.n9 27.2
R4129 a_6144_182.n11 a_6144_182.n0 23.498
R4130 a_6144_182.n3 a_6144_182.n2 23.284
R4131 a_6144_182.n11 a_6144_182.n10 22.4
R4132 a_6144_182.n7 a_6144_182.n4 19.017
R4133 a_6144_182.n6 a_6144_182.n5 13.494
R4134 a_6144_182.t1 a_6144_182.n1 7.04
R4135 a_6144_182.t1 a_6144_182.n3 5.727
R4136 a_6144_182.n8 a_6144_182.n7 1.435
R4137 a_8068_182.n10 a_8068_182.n8 82.852
R4138 a_8068_182.n7 a_8068_182.n6 32.833
R4139 a_8068_182.n8 a_8068_182.t1 32.416
R4140 a_8068_182.n10 a_8068_182.n9 27.2
R4141 a_8068_182.n11 a_8068_182.n0 23.498
R4142 a_8068_182.n3 a_8068_182.n2 23.284
R4143 a_8068_182.n11 a_8068_182.n10 22.4
R4144 a_8068_182.n7 a_8068_182.n4 19.017
R4145 a_8068_182.n6 a_8068_182.n5 13.494
R4146 a_8068_182.t1 a_8068_182.n1 7.04
R4147 a_8068_182.t1 a_8068_182.n3 5.727
R4148 a_8068_182.n8 a_8068_182.n7 1.435
R4149 a_2977_75.n1 a_2977_75.n0 25.576
R4150 a_2977_75.n3 a_2977_75.n2 9.111
R4151 a_2977_75.n7 a_2977_75.n6 2.455
R4152 a_2977_75.n5 a_2977_75.n3 1.964
R4153 a_2977_75.n5 a_2977_75.n4 1.964
R4154 a_2977_75.t0 a_2977_75.n1 1.871
R4155 a_2977_75.n7 a_2977_75.n5 0.636
R4156 a_2977_75.t0 a_2977_75.n7 0.246
R4157 a_1053_75.n1 a_1053_75.n0 25.576
R4158 a_1053_75.n3 a_1053_75.n2 9.111
R4159 a_1053_75.n7 a_1053_75.n6 2.455
R4160 a_1053_75.n5 a_1053_75.n3 1.964
R4161 a_1053_75.n5 a_1053_75.n4 1.964
R4162 a_1053_75.t0 a_1053_75.n1 1.871
R4163 a_1053_75.n7 a_1053_75.n5 0.636
R4164 a_1053_75.t0 a_1053_75.n7 0.246
R4165 a_3939_75.n1 a_3939_75.n0 25.576
R4166 a_3939_75.n3 a_3939_75.n2 9.111
R4167 a_3939_75.n7 a_3939_75.n6 2.455
R4168 a_3939_75.n5 a_3939_75.n3 1.964
R4169 a_3939_75.n5 a_3939_75.n4 1.964
R4170 a_3939_75.t0 a_3939_75.n1 1.871
R4171 a_3939_75.n7 a_3939_75.n5 0.636
R4172 a_3939_75.t0 a_3939_75.n7 0.246
R4173 a_9030_182.n9 a_9030_182.n7 82.852
R4174 a_9030_182.n3 a_9030_182.n1 44.628
R4175 a_9030_182.t0 a_9030_182.n9 32.417
R4176 a_9030_182.n7 a_9030_182.n6 27.2
R4177 a_9030_182.n5 a_9030_182.n4 23.498
R4178 a_9030_182.n3 a_9030_182.n2 23.284
R4179 a_9030_182.n7 a_9030_182.n5 22.4
R4180 a_9030_182.t0 a_9030_182.n11 20.241
R4181 a_9030_182.n11 a_9030_182.n10 13.494
R4182 a_9030_182.t0 a_9030_182.n0 8.137
R4183 a_9030_182.t0 a_9030_182.n3 5.727
R4184 a_9030_182.n9 a_9030_182.n8 1.435
R4185 a_4901_75.n1 a_4901_75.n0 25.576
R4186 a_4901_75.n3 a_4901_75.n2 9.111
R4187 a_4901_75.n7 a_4901_75.n6 2.455
R4188 a_4901_75.n5 a_4901_75.n3 1.964
R4189 a_4901_75.n5 a_4901_75.n4 1.964
R4190 a_4901_75.t0 a_4901_75.n1 1.871
R4191 a_4901_75.n7 a_4901_75.n5 0.636
R4192 a_4901_75.t0 a_4901_75.n7 0.246
R4193 a_6825_75.n5 a_6825_75.n4 19.724
R4194 a_6825_75.t0 a_6825_75.n3 11.595
R4195 a_6825_75.t0 a_6825_75.n5 9.207
R4196 a_6825_75.n2 a_6825_75.n1 2.455
R4197 a_6825_75.n2 a_6825_75.n0 1.32
R4198 a_6825_75.t0 a_6825_75.n2 0.246
R4199 a_18760_73.t0 a_18760_73.n1 34.62
R4200 a_18760_73.t0 a_18760_73.n0 8.137
R4201 a_18760_73.t0 a_18760_73.n2 4.69
R4202 a_11635_75.n5 a_11635_75.n4 19.724
R4203 a_11635_75.t0 a_11635_75.n3 11.595
R4204 a_11635_75.t0 a_11635_75.n5 9.207
R4205 a_11635_75.n2 a_11635_75.n1 2.455
R4206 a_11635_75.n2 a_11635_75.n0 1.32
R4207 a_11635_75.t0 a_11635_75.n2 0.246
R4208 a_5863_75.n5 a_5863_75.n4 19.724
R4209 a_5863_75.t0 a_5863_75.n3 11.595
R4210 a_5863_75.t0 a_5863_75.n5 9.207
R4211 a_5863_75.n2 a_5863_75.n1 2.455
R4212 a_5863_75.n2 a_5863_75.n0 1.32
R4213 a_5863_75.t0 a_5863_75.n2 0.246
R4214 a_7787_75.n5 a_7787_75.n4 19.724
R4215 a_7787_75.t0 a_7787_75.n3 11.595
R4216 a_7787_75.t0 a_7787_75.n5 9.207
R4217 a_7787_75.n2 a_7787_75.n1 2.455
R4218 a_7787_75.n2 a_7787_75.n0 1.32
R4219 a_7787_75.t0 a_7787_75.n2 0.246
R4220 a_9711_75.n1 a_9711_75.n0 25.576
R4221 a_9711_75.n3 a_9711_75.n2 9.111
R4222 a_9711_75.n7 a_9711_75.n6 2.455
R4223 a_9711_75.n5 a_9711_75.n3 1.964
R4224 a_9711_75.n5 a_9711_75.n4 1.964
R4225 a_9711_75.t0 a_9711_75.n1 1.871
R4226 a_9711_75.n7 a_9711_75.n5 0.636
R4227 a_9711_75.t0 a_9711_75.n7 0.246
R4228 a_8749_75.n1 a_8749_75.n0 25.576
R4229 a_8749_75.n3 a_8749_75.n2 9.111
R4230 a_8749_75.n7 a_8749_75.n6 2.455
R4231 a_8749_75.n5 a_8749_75.n3 1.964
R4232 a_8749_75.n5 a_8749_75.n4 1.964
R4233 a_8749_75.t0 a_8749_75.n1 1.871
R4234 a_8749_75.n7 a_8749_75.n5 0.636
R4235 a_8749_75.t0 a_8749_75.n7 0.246
C11 VPB VNB 72.65fF
C12 a_8749_75.n0 VNB 0.09fF
C13 a_8749_75.n1 VNB 0.10fF
C14 a_8749_75.n2 VNB 0.05fF
C15 a_8749_75.n3 VNB 0.03fF
C16 a_8749_75.n4 VNB 0.04fF
C17 a_8749_75.n5 VNB 0.03fF
C18 a_8749_75.n6 VNB 0.04fF
C19 a_9711_75.n0 VNB 0.09fF
C20 a_9711_75.n1 VNB 0.10fF
C21 a_9711_75.n2 VNB 0.05fF
C22 a_9711_75.n3 VNB 0.03fF
C23 a_9711_75.n4 VNB 0.04fF
C24 a_9711_75.n5 VNB 0.03fF
C25 a_9711_75.n6 VNB 0.04fF
C26 a_7787_75.n0 VNB 0.10fF
C27 a_7787_75.n1 VNB 0.04fF
C28 a_7787_75.n2 VNB 0.03fF
C29 a_7787_75.n3 VNB 0.07fF
C30 a_7787_75.n4 VNB 0.08fF
C31 a_7787_75.n5 VNB 0.06fF
C32 a_5863_75.n0 VNB 0.10fF
C33 a_5863_75.n1 VNB 0.04fF
C34 a_5863_75.n2 VNB 0.03fF
C35 a_5863_75.n3 VNB 0.07fF
C36 a_5863_75.n4 VNB 0.08fF
C37 a_5863_75.n5 VNB 0.06fF
C38 a_11635_75.n0 VNB 0.10fF
C39 a_11635_75.n1 VNB 0.04fF
C40 a_11635_75.n2 VNB 0.03fF
C41 a_11635_75.n3 VNB 0.07fF
C42 a_11635_75.n4 VNB 0.08fF
C43 a_11635_75.n5 VNB 0.06fF
C44 a_18760_73.n0 VNB 0.06fF
C45 a_18760_73.n1 VNB 0.13fF
C46 a_18760_73.n2 VNB 0.04fF
C47 a_6825_75.n0 VNB 0.10fF
C48 a_6825_75.n1 VNB 0.04fF
C49 a_6825_75.n2 VNB 0.03fF
C50 a_6825_75.n3 VNB 0.07fF
C51 a_6825_75.n4 VNB 0.08fF
C52 a_6825_75.n5 VNB 0.06fF
C53 a_4901_75.n0 VNB 0.09fF
C54 a_4901_75.n1 VNB 0.10fF
C55 a_4901_75.n2 VNB 0.05fF
C56 a_4901_75.n3 VNB 0.03fF
C57 a_4901_75.n4 VNB 0.04fF
C58 a_4901_75.n5 VNB 0.03fF
C59 a_4901_75.n6 VNB 0.04fF
C60 a_9030_182.n0 VNB 0.07fF
C61 a_9030_182.n1 VNB 0.09fF
C62 a_9030_182.n2 VNB 0.13fF
C63 a_9030_182.n3 VNB 0.11fF
C64 a_9030_182.n4 VNB 0.02fF
C65 a_9030_182.n5 VNB 0.03fF
C66 a_9030_182.n6 VNB 0.02fF
C67 a_9030_182.n7 VNB 0.05fF
C68 a_9030_182.n8 VNB 0.03fF
C69 a_9030_182.n9 VNB 0.11fF
C70 a_9030_182.n10 VNB 0.06fF
C71 a_9030_182.n11 VNB 0.01fF
C72 a_9030_182.t0 VNB 0.33fF
C73 a_3939_75.n0 VNB 0.09fF
C74 a_3939_75.n1 VNB 0.10fF
C75 a_3939_75.n2 VNB 0.05fF
C76 a_3939_75.n3 VNB 0.03fF
C77 a_3939_75.n4 VNB 0.04fF
C78 a_3939_75.n5 VNB 0.03fF
C79 a_3939_75.n6 VNB 0.04fF
C80 a_1053_75.n0 VNB 0.09fF
C81 a_1053_75.n1 VNB 0.10fF
C82 a_1053_75.n2 VNB 0.05fF
C83 a_1053_75.n3 VNB 0.03fF
C84 a_1053_75.n4 VNB 0.04fF
C85 a_1053_75.n5 VNB 0.03fF
C86 a_1053_75.n6 VNB 0.04fF
C87 a_2977_75.n0 VNB 0.09fF
C88 a_2977_75.n1 VNB 0.10fF
C89 a_2977_75.n2 VNB 0.05fF
C90 a_2977_75.n3 VNB 0.03fF
C91 a_2977_75.n4 VNB 0.04fF
C92 a_2977_75.n5 VNB 0.03fF
C93 a_2977_75.n6 VNB 0.04fF
C94 a_8068_182.n0 VNB 0.02fF
C95 a_8068_182.n1 VNB 0.09fF
C96 a_8068_182.n2 VNB 0.13fF
C97 a_8068_182.n3 VNB 0.11fF
C98 a_8068_182.t1 VNB 0.30fF
C99 a_8068_182.n4 VNB 0.09fF
C100 a_8068_182.n5 VNB 0.06fF
C101 a_8068_182.n6 VNB 0.01fF
C102 a_8068_182.n7 VNB 0.03fF
C103 a_8068_182.n8 VNB 0.11fF
C104 a_8068_182.n9 VNB 0.02fF
C105 a_8068_182.n10 VNB 0.05fF
C106 a_8068_182.n11 VNB 0.03fF
C107 a_6144_182.n0 VNB 0.02fF
C108 a_6144_182.n1 VNB 0.09fF
C109 a_6144_182.n2 VNB 0.13fF
C110 a_6144_182.n3 VNB 0.11fF
C111 a_6144_182.t1 VNB 0.30fF
C112 a_6144_182.n4 VNB 0.09fF
C113 a_6144_182.n5 VNB 0.06fF
C114 a_6144_182.n6 VNB 0.01fF
C115 a_6144_182.n7 VNB 0.03fF
C116 a_6144_182.n8 VNB 0.11fF
C117 a_6144_182.n9 VNB 0.02fF
C118 a_6144_182.n10 VNB 0.05fF
C119 a_6144_182.n11 VNB 0.03fF
C120 a_9992_182.n0 VNB 0.07fF
C121 a_9992_182.n1 VNB 0.09fF
C122 a_9992_182.n2 VNB 0.13fF
C123 a_9992_182.n3 VNB 0.11fF
C124 a_9992_182.n4 VNB 0.02fF
C125 a_9992_182.n5 VNB 0.03fF
C126 a_9992_182.n6 VNB 0.02fF
C127 a_9992_182.n7 VNB 0.05fF
C128 a_9992_182.n8 VNB 0.03fF
C129 a_9992_182.n9 VNB 0.11fF
C130 a_9992_182.n10 VNB 0.06fF
C131 a_9992_182.n11 VNB 0.01fF
C132 a_9992_182.t0 VNB 0.33fF
C133 a_17428_73.n0 VNB 0.11fF
C134 a_17428_73.n1 VNB 0.09fF
C135 a_17428_73.n2 VNB 0.08fF
C136 a_17428_73.n3 VNB 0.02fF
C137 a_17428_73.n4 VNB 0.01fF
C138 a_17428_73.n5 VNB 0.06fF
C139 a_11916_182.n0 VNB 0.02fF
C140 a_11916_182.n1 VNB 0.09fF
C141 a_11916_182.n2 VNB 0.13fF
C142 a_11916_182.n3 VNB 0.11fF
C143 a_11916_182.t1 VNB 0.30fF
C144 a_11916_182.n4 VNB 0.09fF
C145 a_11916_182.n5 VNB 0.06fF
C146 a_11916_182.n6 VNB 0.01fF
C147 a_11916_182.n7 VNB 0.03fF
C148 a_11916_182.n8 VNB 0.11fF
C149 a_11916_182.n9 VNB 0.02fF
C150 a_11916_182.n10 VNB 0.05fF
C151 a_11916_182.n11 VNB 0.03fF
C152 a_5182_182.n0 VNB 0.07fF
C153 a_5182_182.n1 VNB 0.09fF
C154 a_5182_182.n2 VNB 0.13fF
C155 a_5182_182.n3 VNB 0.11fF
C156 a_5182_182.n4 VNB 0.02fF
C157 a_5182_182.n5 VNB 0.03fF
C158 a_5182_182.n6 VNB 0.02fF
C159 a_5182_182.n7 VNB 0.05fF
C160 a_5182_182.n8 VNB 0.03fF
C161 a_5182_182.n9 VNB 0.11fF
C162 a_5182_182.n10 VNB 0.06fF
C163 a_5182_182.n11 VNB 0.01fF
C164 a_5182_182.t0 VNB 0.33fF
C165 a_3258_182.n0 VNB 0.07fF
C166 a_3258_182.n1 VNB 0.09fF
C167 a_3258_182.n2 VNB 0.13fF
C168 a_3258_182.n3 VNB 0.11fF
C169 a_3258_182.n4 VNB 0.02fF
C170 a_3258_182.n5 VNB 0.03fF
C171 a_3258_182.n6 VNB 0.02fF
C172 a_3258_182.n7 VNB 0.05fF
C173 a_3258_182.n8 VNB 0.03fF
C174 a_3258_182.n9 VNB 0.11fF
C175 a_3258_182.n10 VNB 0.06fF
C176 a_3258_182.n11 VNB 0.01fF
C177 a_3258_182.t0 VNB 0.33fF
C178 a_1334_182.n0 VNB 0.07fF
C179 a_1334_182.n1 VNB 0.09fF
C180 a_1334_182.n2 VNB 0.13fF
C181 a_1334_182.n3 VNB 0.11fF
C182 a_1334_182.n4 VNB 0.02fF
C183 a_1334_182.n5 VNB 0.03fF
C184 a_1334_182.n6 VNB 0.02fF
C185 a_1334_182.n7 VNB 0.05fF
C186 a_1334_182.n8 VNB 0.03fF
C187 a_1334_182.n9 VNB 0.11fF
C188 a_1334_182.n10 VNB 0.06fF
C189 a_1334_182.n11 VNB 0.01fF
C190 a_1334_182.t0 VNB 0.33fF
C191 a_2015_75.n0 VNB 0.09fF
C192 a_2015_75.n1 VNB 0.10fF
C193 a_2015_75.n2 VNB 0.05fF
C194 a_2015_75.n3 VNB 0.03fF
C195 a_2015_75.n4 VNB 0.04fF
C196 a_2015_75.n5 VNB 0.03fF
C197 a_2015_75.n6 VNB 0.04fF
C198 a_7106_182.n0 VNB 0.02fF
C199 a_7106_182.n1 VNB 0.09fF
C200 a_7106_182.n2 VNB 0.13fF
C201 a_7106_182.n3 VNB 0.11fF
C202 a_7106_182.t1 VNB 0.30fF
C203 a_7106_182.n4 VNB 0.09fF
C204 a_7106_182.n5 VNB 0.06fF
C205 a_7106_182.n6 VNB 0.01fF
C206 a_7106_182.n7 VNB 0.03fF
C207 a_7106_182.n8 VNB 0.11fF
C208 a_7106_182.n9 VNB 0.02fF
C209 a_7106_182.n10 VNB 0.05fF
C210 a_7106_182.n11 VNB 0.03fF
C211 a_15764_182.n0 VNB 0.07fF
C212 a_15764_182.n1 VNB 0.09fF
C213 a_15764_182.n2 VNB 0.13fF
C214 a_15764_182.n3 VNB 0.11fF
C215 a_15764_182.n4 VNB 0.02fF
C216 a_15764_182.n5 VNB 0.03fF
C217 a_15764_182.n6 VNB 0.06fF
C218 a_15764_182.n7 VNB 0.03fF
C219 a_15764_182.n8 VNB 0.12fF
C220 a_15764_182.n9 VNB 0.06fF
C221 a_15764_182.n10 VNB 0.01fF
C222 a_15764_182.t0 VNB 0.33fF
C223 a_13840_182.n0 VNB 0.07fF
C224 a_13840_182.n1 VNB 0.09fF
C225 a_13840_182.n2 VNB 0.13fF
C226 a_13840_182.n3 VNB 0.11fF
C227 a_13840_182.n4 VNB 0.02fF
C228 a_13840_182.n5 VNB 0.03fF
C229 a_13840_182.n6 VNB 0.06fF
C230 a_13840_182.n7 VNB 0.03fF
C231 a_13840_182.n8 VNB 0.12fF
C232 a_13840_182.n9 VNB 0.06fF
C233 a_13840_182.n10 VNB 0.01fF
C234 a_13840_182.t0 VNB 0.33fF
C235 a_13559_75.n0 VNB 0.09fF
C236 a_13559_75.n1 VNB 0.10fF
C237 a_13559_75.n2 VNB 0.05fF
C238 a_13559_75.n3 VNB 0.03fF
C239 a_13559_75.n4 VNB 0.04fF
C240 a_13559_75.n5 VNB 0.11fF
C241 a_13559_75.n6 VNB 0.04fF
C242 Q.n0 VNB 0.73fF
C243 Q.n1 VNB 0.47fF
C244 Q.n2 VNB 0.50fF
C245 Q.n3 VNB 0.01fF
C246 a_4125_1004.n0 VNB 0.54fF
C247 a_4125_1004.n1 VNB 0.54fF
C248 a_4125_1004.n2 VNB 0.64fF
C249 a_4125_1004.n3 VNB 0.20fF
C250 a_4125_1004.n4 VNB 0.38fF
C251 a_4125_1004.n5 VNB 0.41fF
C252 a_4125_1004.n6 VNB 0.64fF
C253 a_4125_1004.n7 VNB 0.64fF
C254 a_4125_1004.n8 VNB 0.08fF
C255 a_4125_1004.n9 VNB 0.21fF
C256 a_4125_1004.n10 VNB 0.05fF
C257 a_4220_182.n0 VNB 0.02fF
C258 a_4220_182.n1 VNB 0.07fF
C259 a_4220_182.n2 VNB 0.13fF
C260 a_4220_182.n3 VNB 0.09fF
C261 a_4220_182.t1 VNB 0.25fF
C262 a_4220_182.n4 VNB 0.05fF
C263 a_4220_182.n5 VNB 0.06fF
C264 a_4220_182.n6 VNB 0.07fF
C265 a_4220_182.n7 VNB 0.07fF
C266 a_4220_182.n8 VNB 0.03fF
C267 a_4220_182.n9 VNB 0.01fF
C268 a_4220_182.n10 VNB 0.11fF
C269 a_4220_182.n11 VNB 0.02fF
C270 a_4220_182.n12 VNB 0.05fF
C271 a_4220_182.n13 VNB 0.03fF
C272 a_13745_1004.n0 VNB 0.04fF
C273 a_13745_1004.n1 VNB 0.55fF
C274 a_13745_1004.n2 VNB 0.55fF
C275 a_13745_1004.n3 VNB 0.65fF
C276 a_13745_1004.n4 VNB 0.20fF
C277 a_13745_1004.n5 VNB 0.39fF
C278 a_13745_1004.n6 VNB 0.42fF
C279 a_13745_1004.n7 VNB 0.65fF
C280 a_13745_1004.n8 VNB 0.64fF
C281 a_13745_1004.n9 VNB 0.04fF
C282 a_13745_1004.n10 VNB 0.22fF
C283 a_13745_1004.n11 VNB 0.06fF
C284 a_13105_943.n0 VNB 0.91fF
C285 a_13105_943.n1 VNB 0.91fF
C286 a_13105_943.n2 VNB 1.07fF
C287 a_13105_943.n3 VNB 0.34fF
C288 a_13105_943.n4 VNB 0.49fF
C289 a_13105_943.n5 VNB 0.61fF
C290 a_13105_943.t15 VNB 0.93fF
C291 a_13105_943.n6 VNB 0.72fF
C292 a_13105_943.n7 VNB 0.61fF
C293 a_13105_943.t13 VNB 0.93fF
C294 a_13105_943.n8 VNB 0.62fF
C295 a_13105_943.n9 VNB 0.61fF
C296 a_13105_943.t9 VNB 0.93fF
C297 a_13105_943.n10 VNB 0.65fF
C298 a_13105_943.n11 VNB 2.14fF
C299 a_13105_943.n12 VNB 3.20fF
C300 a_13105_943.n13 VNB 0.77fF
C301 a_13105_943.n14 VNB 0.14fF
C302 a_13105_943.n15 VNB 0.52fF
C303 a_13105_943.n16 VNB 0.08fF
C304 a_372_182.n0 VNB 0.02fF
C305 a_372_182.n1 VNB 0.09fF
C306 a_372_182.n2 VNB 0.13fF
C307 a_372_182.n3 VNB 0.11fF
C308 a_372_182.t1 VNB 0.30fF
C309 a_372_182.n4 VNB 0.09fF
C310 a_372_182.n5 VNB 0.06fF
C311 a_372_182.n6 VNB 0.01fF
C312 a_372_182.n7 VNB 0.03fF
C313 a_372_182.n8 VNB 0.11fF
C314 a_372_182.n9 VNB 0.02fF
C315 a_372_182.n10 VNB 0.05fF
C316 a_372_182.n11 VNB 0.02fF
C317 a_91_75.n0 VNB 0.19fF
C318 a_91_75.n1 VNB 0.04fF
C319 a_91_75.n2 VNB 0.01fF
C320 a_91_75.n3 VNB 0.08fF
C321 a_91_75.n4 VNB 0.06fF
C322 a_91_75.n5 VNB 0.06fF
C323 a_2201_1004.n0 VNB 0.54fF
C324 a_2201_1004.n1 VNB 0.54fF
C325 a_2201_1004.n2 VNB 0.64fF
C326 a_2201_1004.n3 VNB 0.20fF
C327 a_2201_1004.n4 VNB 0.38fF
C328 a_2201_1004.n5 VNB 0.41fF
C329 a_2201_1004.n6 VNB 0.64fF
C330 a_2201_1004.n7 VNB 0.64fF
C331 a_2201_1004.n8 VNB 0.08fF
C332 a_2201_1004.n9 VNB 0.21fF
C333 a_2201_1004.n10 VNB 0.05fF
C334 a_2296_182.n0 VNB 0.07fF
C335 a_2296_182.n1 VNB 0.13fF
C336 a_2296_182.n2 VNB 0.07fF
C337 a_2296_182.n3 VNB 0.02fF
C338 a_2296_182.n4 VNB 0.03fF
C339 a_2296_182.n5 VNB 0.02fF
C340 a_2296_182.n6 VNB 0.05fF
C341 a_2296_182.n7 VNB 0.05fF
C342 a_2296_182.n8 VNB 0.06fF
C343 a_2296_182.n9 VNB 0.07fF
C344 a_2296_182.n10 VNB 0.07fF
C345 a_2296_182.n11 VNB 0.03fF
C346 a_2296_182.n12 VNB 0.01fF
C347 a_2296_182.n13 VNB 0.11fF
C348 a_2296_182.t0 VNB 0.28fF
C349 a_1561_943.n0 VNB 0.07fF
C350 a_1561_943.n1 VNB 0.93fF
C351 a_1561_943.n2 VNB 0.93fF
C352 a_1561_943.n3 VNB 1.10fF
C353 a_1561_943.n4 VNB 0.35fF
C354 a_1561_943.n5 VNB 0.50fF
C355 a_1561_943.n6 VNB 0.62fF
C356 a_1561_943.t10 VNB 0.95fF
C357 a_1561_943.n7 VNB 0.73fF
C358 a_1561_943.n8 VNB 0.62fF
C359 a_1561_943.t7 VNB 0.95fF
C360 a_1561_943.n9 VNB 0.63fF
C361 a_1561_943.n10 VNB 0.62fF
C362 a_1561_943.t9 VNB 0.95fF
C363 a_1561_943.n11 VNB 0.66fF
C364 a_1561_943.n12 VNB 2.19fF
C365 a_1561_943.n13 VNB 3.27fF
C366 a_1561_943.n14 VNB 0.77fF
C367 a_1561_943.n15 VNB 0.06fF
C368 a_1561_943.n16 VNB 0.54fF
C369 a_1561_943.n17 VNB 0.09fF
C370 a_9897_1004.n0 VNB 0.04fF
C371 a_9897_1004.n1 VNB 0.55fF
C372 a_9897_1004.n2 VNB 0.55fF
C373 a_9897_1004.n3 VNB 0.65fF
C374 a_9897_1004.n4 VNB 0.20fF
C375 a_9897_1004.n5 VNB 0.39fF
C376 a_9897_1004.n6 VNB 0.42fF
C377 a_9897_1004.n7 VNB 0.65fF
C378 a_9897_1004.n8 VNB 0.64fF
C379 a_9897_1004.n9 VNB 0.04fF
C380 a_9897_1004.n10 VNB 0.22fF
C381 a_9897_1004.n11 VNB 0.06fF
C382 a_599_943.n0 VNB 0.83fF
C383 a_599_943.n1 VNB 0.83fF
C384 a_599_943.n2 VNB 0.98fF
C385 a_599_943.n3 VNB 0.31fF
C386 a_599_943.n4 VNB 0.49fF
C387 a_599_943.n5 VNB 0.54fF
C388 a_599_943.n6 VNB 0.87fF
C389 a_599_943.n7 VNB 0.60fF
C390 a_599_943.t11 VNB 0.80fF
C391 a_599_943.n8 VNB 0.59fF
C392 a_599_943.n9 VNB 4.22fF
C393 a_599_943.n10 VNB 0.70fF
C394 a_599_943.n11 VNB 0.13fF
C395 a_599_943.n12 VNB 0.42fF
C396 a_599_943.n13 VNB 0.07fF
C397 a_15669_1004.n0 VNB 0.04fF
C398 a_15669_1004.n1 VNB 0.52fF
C399 a_15669_1004.n2 VNB 0.52fF
C400 a_15669_1004.n3 VNB 0.61fF
C401 a_15669_1004.n4 VNB 0.19fF
C402 a_15669_1004.n5 VNB 0.37fF
C403 a_15669_1004.n6 VNB 0.40fF
C404 a_15669_1004.n7 VNB 0.61fF
C405 a_15669_1004.n8 VNB 0.61fF
C406 a_15669_1004.n9 VNB 0.03fF
C407 a_15669_1004.n10 VNB 0.21fF
C408 a_15669_1004.n11 VNB 0.05fF
C409 a_12878_182.n0 VNB 0.07fF
C410 a_12878_182.n1 VNB 0.09fF
C411 a_12878_182.n2 VNB 0.13fF
C412 a_12878_182.n3 VNB 0.11fF
C413 a_12878_182.n4 VNB 0.02fF
C414 a_12878_182.n5 VNB 0.03fF
C415 a_12878_182.n6 VNB 0.06fF
C416 a_12878_182.n7 VNB 0.03fF
C417 a_12878_182.n8 VNB 0.12fF
C418 a_12878_182.n9 VNB 0.06fF
C419 a_12878_182.n10 VNB 0.01fF
C420 a_12878_182.t0 VNB 0.33fF
C421 a_12597_75.n0 VNB 0.09fF
C422 a_12597_75.n1 VNB 0.10fF
C423 a_12597_75.n2 VNB 0.05fF
C424 a_12597_75.n3 VNB 0.03fF
C425 a_12597_75.n4 VNB 0.04fF
C426 a_12597_75.n5 VNB 0.11fF
C427 a_12597_75.n6 VNB 0.04fF
C428 a_10954_182.n0 VNB 0.02fF
C429 a_10954_182.n1 VNB 0.09fF
C430 a_10954_182.n2 VNB 0.13fF
C431 a_10954_182.n3 VNB 0.11fF
C432 a_10954_182.t1 VNB 0.30fF
C433 a_10954_182.n4 VNB 0.09fF
C434 a_10954_182.n5 VNB 0.06fF
C435 a_10954_182.n6 VNB 0.01fF
C436 a_10954_182.n7 VNB 0.03fF
C437 a_10954_182.n8 VNB 0.11fF
C438 a_10954_182.n9 VNB 0.02fF
C439 a_10954_182.n10 VNB 0.05fF
C440 a_10954_182.n11 VNB 0.02fF
C441 a_10673_75.n0 VNB 0.20fF
C442 a_10673_75.n1 VNB 0.04fF
C443 a_10673_75.n2 VNB 0.01fF
C444 a_10673_75.n3 VNB 0.08fF
C445 a_10673_75.n4 VNB 0.06fF
C446 a_10673_75.n5 VNB 0.07fF
C447 a_16726_182.n0 VNB 0.02fF
C448 a_16726_182.n1 VNB 0.09fF
C449 a_16726_182.n2 VNB 0.13fF
C450 a_16726_182.n3 VNB 0.11fF
C451 a_16726_182.t1 VNB 0.30fF
C452 a_16726_182.n4 VNB 0.09fF
C453 a_16726_182.n5 VNB 0.06fF
C454 a_16726_182.n6 VNB 0.01fF
C455 a_16726_182.n7 VNB 0.03fF
C456 a_16726_182.n8 VNB 0.11fF
C457 a_16726_182.n9 VNB 0.02fF
C458 a_16726_182.n10 VNB 0.05fF
C459 a_16726_182.n11 VNB 0.02fF
C460 a_16445_75.n0 VNB 0.20fF
C461 a_16445_75.n1 VNB 0.04fF
C462 a_16445_75.n2 VNB 0.01fF
C463 a_16445_75.n3 VNB 0.08fF
C464 a_16445_75.n4 VNB 0.06fF
C465 a_16445_75.n5 VNB 0.07fF
C466 a_18094_73.n0 VNB 0.13fF
C467 a_18094_73.n1 VNB 0.13fF
C468 a_18094_73.n2 VNB 0.14fF
C469 a_15991_943.n0 VNB 0.04fF
C470 a_15991_943.n1 VNB 0.48fF
C471 a_15991_943.n2 VNB 0.48fF
C472 a_15991_943.n3 VNB 0.56fF
C473 a_15991_943.n4 VNB 0.18fF
C474 a_15991_943.n5 VNB 0.36fF
C475 a_15991_943.n6 VNB 0.41fF
C476 a_15991_943.n7 VNB 0.38fF
C477 a_15991_943.n8 VNB 0.41fF
C478 a_15991_943.t7 VNB 0.39fF
C479 a_15991_943.n9 VNB 0.38fF
C480 a_15991_943.n10 VNB 0.75fF
C481 a_15991_943.n11 VNB 0.43fF
C482 a_15991_943.t11 VNB 0.39fF
C483 a_15991_943.n12 VNB 0.34fF
C484 a_15991_943.n13 VNB 1.29fF
C485 a_15991_943.n14 VNB 0.40fF
C486 a_15991_943.n15 VNB 0.03fF
C487 a_15991_943.n16 VNB 0.16fF
C488 a_15991_943.n17 VNB 0.05fF
C489 a_11821_1004.n0 VNB 0.05fF
C490 a_11821_1004.n1 VNB 0.68fF
C491 a_11821_1004.n2 VNB 0.68fF
C492 a_11821_1004.n3 VNB 0.80fF
C493 a_11821_1004.n4 VNB 0.25fF
C494 a_11821_1004.n5 VNB 0.48fF
C495 a_11821_1004.n6 VNB 0.52fF
C496 a_11821_1004.n7 VNB 0.60fF
C497 a_11821_1004.n8 VNB 0.52fF
C498 a_11821_1004.n9 VNB 0.58fF
C499 a_11821_1004.n10 VNB 1.44fF
C500 a_11821_1004.n11 VNB 0.57fF
C501 a_11821_1004.n12 VNB 0.04fF
C502 a_11821_1004.n13 VNB 0.28fF
C503 a_11821_1004.n14 VNB 0.07fF
C504 a_277_1004.n0 VNB 0.55fF
C505 a_277_1004.n1 VNB 0.55fF
C506 a_277_1004.n2 VNB 0.65fF
C507 a_277_1004.n3 VNB 0.20fF
C508 a_277_1004.n4 VNB 0.39fF
C509 a_277_1004.n5 VNB 0.42fF
C510 a_277_1004.n6 VNB 0.49fF
C511 a_277_1004.n7 VNB 0.42fF
C512 a_277_1004.n8 VNB 0.47fF
C513 a_277_1004.n9 VNB 1.16fF
C514 a_277_1004.n10 VNB 0.47fF
C515 a_277_1004.n11 VNB 0.09fF
C516 a_277_1004.n12 VNB 0.21fF
C517 a_277_1004.n13 VNB 0.05fF
C518 a_14802_182.n0 VNB 0.07fF
C519 a_14802_182.n1 VNB 0.13fF
C520 a_14802_182.n2 VNB 0.07fF
C521 a_14802_182.n3 VNB 0.02fF
C522 a_14802_182.n4 VNB 0.03fF
C523 a_14802_182.n5 VNB 0.06fF
C524 a_14802_182.n6 VNB 0.05fF
C525 a_14802_182.n7 VNB 0.06fF
C526 a_14802_182.n8 VNB 0.07fF
C527 a_14802_182.n9 VNB 0.07fF
C528 a_14802_182.n10 VNB 0.03fF
C529 a_14802_182.n11 VNB 0.01fF
C530 a_14802_182.n12 VNB 0.12fF
C531 a_14802_182.t0 VNB 0.28fF
C532 a_14521_75.n0 VNB 0.20fF
C533 a_14521_75.n1 VNB 0.04fF
C534 a_14521_75.n2 VNB 0.01fF
C535 a_14521_75.n3 VNB 0.08fF
C536 a_14521_75.n4 VNB 0.06fF
C537 a_14521_75.n5 VNB 0.07fF
C538 a_17533_1005.n0 VNB 0.40fF
C539 a_17533_1005.n1 VNB 0.32fF
C540 a_17533_1005.n2 VNB 0.23fF
C541 a_17533_1005.n3 VNB 0.62fF
C542 a_17533_1005.n4 VNB 0.28fF
C543 a_17533_1005.n5 VNB 0.36fF
C544 a_18197_1005.n0 VNB 0.29fF
C545 a_18197_1005.n1 VNB 0.28fF
C546 a_18197_1005.n2 VNB 0.36fF
C547 a_18197_1005.n3 VNB 0.25fF
C548 a_18197_1005.n4 VNB 0.57fF
C549 a_18197_1005.n5 VNB 0.20fF
C550 a_17708_181.n0 VNB 0.03fF
C551 a_17708_181.n1 VNB 0.39fF
C552 a_17708_181.n2 VNB 0.47fF
C553 a_17708_181.n3 VNB 0.22fF
C554 a_17708_181.n4 VNB 0.25fF
C555 a_17708_181.n5 VNB 0.50fF
C556 a_17708_181.n6 VNB 0.46fF
C557 a_17708_181.n7 VNB 0.05fF
C558 a_17708_181.n8 VNB 0.03fF
C559 a_17708_181.n9 VNB 0.08fF
C560 a_17708_181.n10 VNB 0.27fF
C561 a_17708_181.n11 VNB 0.03fF
C562 a_17708_181.n12 VNB 0.05fF
C563 a_17708_181.n13 VNB 0.03fF
C564 a_17708_181.n14 VNB 0.09fF
C565 a_17708_181.n15 VNB 1.00fF
C566 a_17708_181.n16 VNB 0.02fF
C567 a_17708_181.n17 VNB 0.08fF
C568 a_17708_181.n18 VNB 0.05fF
C569 a_10219_943.n0 VNB 0.08fF
C570 a_10219_943.n1 VNB 1.09fF
C571 a_10219_943.n2 VNB 1.09fF
C572 a_10219_943.n3 VNB 1.28fF
C573 a_10219_943.n4 VNB 0.40fF
C574 a_10219_943.n5 VNB 0.59fF
C575 a_10219_943.n6 VNB 0.66fF
C576 a_10219_943.t13 VNB 1.16fF
C577 a_10219_943.n7 VNB 0.87fF
C578 a_10219_943.n8 VNB 0.59fF
C579 a_10219_943.t9 VNB 1.17fF
C580 a_10219_943.n9 VNB 0.76fF
C581 a_10219_943.n10 VNB 11.60fF
C582 a_10219_943.n11 VNB 1.68fF
C583 a_10219_943.n12 VNB 0.79fF
C584 a_10219_943.t10 VNB 1.05fF
C585 a_10219_943.n13 VNB 1.71fF
C586 a_10219_943.n14 VNB 1.51fF
C587 a_10219_943.n15 VNB 0.07fF
C588 a_10219_943.n16 VNB 0.57fF
C589 a_10219_943.n17 VNB 0.11fF
C590 a_7973_1004.n0 VNB 0.04fF
C591 a_7973_1004.n1 VNB 0.55fF
C592 a_7973_1004.n2 VNB 0.55fF
C593 a_7973_1004.n3 VNB 0.65fF
C594 a_7973_1004.n4 VNB 0.20fF
C595 a_7973_1004.n5 VNB 0.39fF
C596 a_7973_1004.n6 VNB 0.42fF
C597 a_7973_1004.n7 VNB 0.65fF
C598 a_7973_1004.n8 VNB 0.64fF
C599 a_7973_1004.n9 VNB 0.04fF
C600 a_7973_1004.n10 VNB 0.22fF
C601 a_7973_1004.n11 VNB 0.06fF
C602 a_6049_1004.n0 VNB 0.05fF
C603 a_6049_1004.n1 VNB 0.68fF
C604 a_6049_1004.n2 VNB 0.68fF
C605 a_6049_1004.n3 VNB 0.80fF
C606 a_6049_1004.n4 VNB 0.25fF
C607 a_6049_1004.n5 VNB 0.48fF
C608 a_6049_1004.n6 VNB 0.52fF
C609 a_6049_1004.n7 VNB 0.60fF
C610 a_6049_1004.n8 VNB 0.52fF
C611 a_6049_1004.n9 VNB 0.58fF
C612 a_6049_1004.n10 VNB 1.44fF
C613 a_6049_1004.n11 VNB 0.57fF
C614 a_6049_1004.n12 VNB 0.04fF
C615 a_6049_1004.n13 VNB 0.28fF
C616 a_6049_1004.n14 VNB 0.07fF
C617 a_15483_75.n0 VNB 0.03fF
C618 a_15483_75.n1 VNB 0.10fF
C619 a_15483_75.n2 VNB 0.10fF
C620 a_15483_75.n3 VNB 0.05fF
C621 a_15483_75.n4 VNB 0.03fF
C622 a_15483_75.n5 VNB 0.04fF
C623 a_15483_75.n6 VNB 0.11fF
C624 a_15483_75.n7 VNB 0.04fF
C625 a_12143_943.n0 VNB 0.08fF
C626 a_12143_943.n1 VNB 1.01fF
C627 a_12143_943.n2 VNB 1.01fF
C628 a_12143_943.n3 VNB 1.19fF
C629 a_12143_943.n4 VNB 0.37fF
C630 a_12143_943.n5 VNB 0.60fF
C631 a_12143_943.n6 VNB 0.66fF
C632 a_12143_943.n7 VNB 1.06fF
C633 a_12143_943.n8 VNB 0.73fF
C634 a_12143_943.t9 VNB 0.97fF
C635 a_12143_943.n9 VNB 0.72fF
C636 a_12143_943.n10 VNB 5.12fF
C637 a_12143_943.n11 VNB 0.83fF
C638 a_12143_943.n12 VNB 0.06fF
C639 a_12143_943.n13 VNB 0.53fF
C640 a_12143_943.n14 VNB 0.10fF
C641 a_7333_943.n0 VNB 0.08fF
C642 a_7333_943.n1 VNB 1.00fF
C643 a_7333_943.n2 VNB 1.00fF
C644 a_7333_943.n3 VNB 1.17fF
C645 a_7333_943.n4 VNB 0.37fF
C646 a_7333_943.n5 VNB 0.54fF
C647 a_7333_943.n6 VNB 0.66fF
C648 a_7333_943.t11 VNB 1.01fF
C649 a_7333_943.n7 VNB 0.78fF
C650 a_7333_943.n8 VNB 0.66fF
C651 a_7333_943.t9 VNB 1.01fF
C652 a_7333_943.n9 VNB 0.67fF
C653 a_7333_943.n10 VNB 0.66fF
C654 a_7333_943.t8 VNB 1.01fF
C655 a_7333_943.n11 VNB 0.71fF
C656 a_7333_943.n12 VNB 2.35fF
C657 a_7333_943.n13 VNB 3.51fF
C658 a_7333_943.n14 VNB 0.83fF
C659 a_7333_943.n15 VNB 0.06fF
C660 a_7333_943.n16 VNB 0.58fF
C661 a_7333_943.n17 VNB 0.10fF
C662 a_6371_943.n0 VNB 0.99fF
C663 a_6371_943.n1 VNB 0.99fF
C664 a_6371_943.n2 VNB 1.16fF
C665 a_6371_943.n3 VNB 0.37fF
C666 a_6371_943.n4 VNB 0.59fF
C667 a_6371_943.n5 VNB 0.64fF
C668 a_6371_943.n6 VNB 1.04fF
C669 a_6371_943.n7 VNB 0.71fF
C670 a_6371_943.t9 VNB 0.95fF
C671 a_6371_943.n8 VNB 0.71fF
C672 a_6371_943.n9 VNB 5.02fF
C673 a_6371_943.n10 VNB 0.83fF
C674 a_6371_943.n11 VNB 0.15fF
C675 a_6371_943.n12 VNB 0.50fF
C676 a_6371_943.n13 VNB 0.08fF
C677 a_4447_943.n0 VNB 1.10fF
C678 a_4447_943.n1 VNB 1.10fF
C679 a_4447_943.n2 VNB 1.29fF
C680 a_4447_943.n3 VNB 0.41fF
C681 a_4447_943.n4 VNB 0.39fF
C682 a_4447_943.n5 VNB 0.59fF
C683 a_4447_943.n6 VNB 0.84fF
C684 a_4447_943.n7 VNB 0.53fF
C685 a_4447_943.n8 VNB 0.97fF
C686 a_4447_943.n9 VNB 17.57fF
C687 a_4447_943.n10 VNB 4.08fF
C688 a_4447_943.n11 VNB 0.79fF
C689 a_4447_943.t8 VNB 1.06fF
C690 a_4447_943.n12 VNB 1.71fF
C691 a_4447_943.n13 VNB 1.72fF
C692 a_4447_943.n14 VNB 0.17fF
C693 a_4447_943.n15 VNB 0.56fF
C694 a_4447_943.n16 VNB 0.09fF
C695 VPB.n0 VNB 0.03fF
C696 VPB.n1 VNB 0.04fF
C697 VPB.n2 VNB 0.02fF
C698 VPB.n3 VNB 0.19fF
C699 VPB.n5 VNB 0.02fF
C700 VPB.n6 VNB 0.02fF
C701 VPB.n7 VNB 0.02fF
C702 VPB.n8 VNB 0.02fF
C703 VPB.n10 VNB 0.02fF
C704 VPB.n11 VNB 0.02fF
C705 VPB.n12 VNB 0.02fF
C706 VPB.n14 VNB 0.10fF
C707 VPB.n15 VNB 0.10fF
C708 VPB.n16 VNB 0.02fF
C709 VPB.n17 VNB 0.02fF
C710 VPB.n18 VNB 0.02fF
C711 VPB.n19 VNB 0.04fF
C712 VPB.n20 VNB 0.02fF
C713 VPB.n21 VNB 0.29fF
C714 VPB.n22 VNB 0.04fF
C715 VPB.n24 VNB 0.02fF
C716 VPB.n25 VNB 0.02fF
C717 VPB.n26 VNB 0.02fF
C718 VPB.n27 VNB 0.02fF
C719 VPB.n29 VNB 0.02fF
C720 VPB.n30 VNB 0.02fF
C721 VPB.n31 VNB 0.02fF
C722 VPB.n33 VNB 0.28fF
C723 VPB.n35 VNB 0.03fF
C724 VPB.n36 VNB 0.02fF
C725 VPB.n37 VNB 0.03fF
C726 VPB.n38 VNB 0.03fF
C727 VPB.n39 VNB 0.28fF
C728 VPB.n40 VNB 0.01fF
C729 VPB.n41 VNB 0.02fF
C730 VPB.n42 VNB 0.28fF
C731 VPB.n43 VNB 0.02fF
C732 VPB.n44 VNB 0.02fF
C733 VPB.n45 VNB 0.05fF
C734 VPB.n46 VNB 0.21fF
C735 VPB.n47 VNB 0.02fF
C736 VPB.n48 VNB 0.01fF
C737 VPB.n49 VNB 0.14fF
C738 VPB.n50 VNB 0.16fF
C739 VPB.n51 VNB 0.02fF
C740 VPB.n52 VNB 0.02fF
C741 VPB.n53 VNB 0.14fF
C742 VPB.n54 VNB 0.16fF
C743 VPB.n55 VNB 0.02fF
C744 VPB.n56 VNB 0.02fF
C745 VPB.n57 VNB 0.02fF
C746 VPB.n58 VNB 0.14fF
C747 VPB.n59 VNB 0.15fF
C748 VPB.n60 VNB 0.02fF
C749 VPB.n61 VNB 0.02fF
C750 VPB.n62 VNB 0.14fF
C751 VPB.n63 VNB 0.15fF
C752 VPB.n64 VNB 0.02fF
C753 VPB.n65 VNB 0.02fF
C754 VPB.n66 VNB 0.02fF
C755 VPB.n67 VNB 0.14fF
C756 VPB.n68 VNB 0.16fF
C757 VPB.n69 VNB 0.02fF
C758 VPB.n70 VNB 0.02fF
C759 VPB.n71 VNB 0.14fF
C760 VPB.n72 VNB 0.16fF
C761 VPB.n73 VNB 0.02fF
C762 VPB.n74 VNB 0.02fF
C763 VPB.n75 VNB 0.21fF
C764 VPB.n76 VNB 0.02fF
C765 VPB.n77 VNB 0.01fF
C766 VPB.n78 VNB 0.06fF
C767 VPB.n79 VNB 0.28fF
C768 VPB.n80 VNB 0.02fF
C769 VPB.n81 VNB 0.02fF
C770 VPB.n82 VNB 0.10fF
C771 VPB.n83 VNB 0.10fF
C772 VPB.n84 VNB 0.02fF
C773 VPB.n85 VNB 0.02fF
C774 VPB.n86 VNB 0.02fF
C775 VPB.n87 VNB 0.04fF
C776 VPB.n88 VNB 0.02fF
C777 VPB.n89 VNB 0.29fF
C778 VPB.n90 VNB 0.04fF
C779 VPB.n92 VNB 0.02fF
C780 VPB.n93 VNB 0.02fF
C781 VPB.n94 VNB 0.02fF
C782 VPB.n95 VNB 0.02fF
C783 VPB.n97 VNB 0.02fF
C784 VPB.n98 VNB 0.02fF
C785 VPB.n99 VNB 0.02fF
C786 VPB.n101 VNB 0.28fF
C787 VPB.n103 VNB 0.03fF
C788 VPB.n104 VNB 0.02fF
C789 VPB.n105 VNB 0.28fF
C790 VPB.n106 VNB 0.02fF
C791 VPB.n107 VNB 0.02fF
C792 VPB.n108 VNB 0.28fF
C793 VPB.n109 VNB 0.01fF
C794 VPB.n110 VNB 0.02fF
C795 VPB.n111 VNB 0.03fF
C796 VPB.n112 VNB 0.03fF
C797 VPB.n113 VNB 0.28fF
C798 VPB.n114 VNB 0.01fF
C799 VPB.n115 VNB 0.02fF
C800 VPB.n116 VNB 0.28fF
C801 VPB.n117 VNB 0.02fF
C802 VPB.n118 VNB 0.02fF
C803 VPB.n119 VNB 0.05fF
C804 VPB.n120 VNB 0.21fF
C805 VPB.n121 VNB 0.02fF
C806 VPB.n122 VNB 0.01fF
C807 VPB.n123 VNB 0.14fF
C808 VPB.n124 VNB 0.16fF
C809 VPB.n125 VNB 0.02fF
C810 VPB.n126 VNB 0.02fF
C811 VPB.n127 VNB 0.14fF
C812 VPB.n128 VNB 0.16fF
C813 VPB.n129 VNB 0.02fF
C814 VPB.n130 VNB 0.02fF
C815 VPB.n131 VNB 0.02fF
C816 VPB.n132 VNB 0.14fF
C817 VPB.n133 VNB 0.15fF
C818 VPB.n134 VNB 0.02fF
C819 VPB.n135 VNB 0.02fF
C820 VPB.n136 VNB 0.14fF
C821 VPB.n137 VNB 0.15fF
C822 VPB.n138 VNB 0.02fF
C823 VPB.n139 VNB 0.02fF
C824 VPB.n140 VNB 0.02fF
C825 VPB.n141 VNB 0.14fF
C826 VPB.n142 VNB 0.16fF
C827 VPB.n143 VNB 0.02fF
C828 VPB.n144 VNB 0.02fF
C829 VPB.n145 VNB 0.02fF
C830 VPB.n146 VNB 0.02fF
C831 VPB.n147 VNB 0.02fF
C832 VPB.n148 VNB 0.11fF
C833 VPB.n149 VNB 0.03fF
C834 VPB.n150 VNB 0.02fF
C835 VPB.n151 VNB 0.05fF
C836 VPB.n152 VNB 0.01fF
C837 VPB.n154 VNB 0.02fF
C838 VPB.n155 VNB 0.02fF
C839 VPB.n156 VNB 0.02fF
C840 VPB.n157 VNB 0.02fF
C841 VPB.n160 VNB 0.02fF
C842 VPB.n162 VNB 0.46fF
C843 VPB.n164 VNB 0.04fF
C844 VPB.n165 VNB 0.04fF
C845 VPB.n166 VNB 0.28fF
C846 VPB.n167 VNB 0.03fF
C847 VPB.n168 VNB 0.03fF
C848 VPB.n169 VNB 0.06fF
C849 VPB.n170 VNB 0.14fF
C850 VPB.n171 VNB 0.19fF
C851 VPB.n172 VNB 0.02fF
C852 VPB.n173 VNB 0.01fF
C853 VPB.n174 VNB 0.07fF
C854 VPB.n175 VNB 0.16fF
C855 VPB.n176 VNB 0.02fF
C856 VPB.n177 VNB 0.02fF
C857 VPB.n178 VNB 0.02fF
C858 VPB.n179 VNB 0.06fF
C859 VPB.n180 VNB 0.14fF
C860 VPB.n181 VNB 0.20fF
C861 VPB.n182 VNB 0.02fF
C862 VPB.n183 VNB 0.01fF
C863 VPB.n184 VNB 0.02fF
C864 VPB.n185 VNB 0.28fF
C865 VPB.n186 VNB 0.01fF
C866 VPB.n187 VNB 0.02fF
C867 VPB.n188 VNB 0.04fF
C868 VPB.n189 VNB 0.02fF
C869 VPB.n190 VNB 0.02fF
C870 VPB.n191 VNB 0.02fF
C871 VPB.n192 VNB 0.04fF
C872 VPB.n193 VNB 0.02fF
C873 VPB.n194 VNB 0.17fF
C874 VPB.n195 VNB 0.04fF
C875 VPB.n197 VNB 0.02fF
C876 VPB.n198 VNB 0.02fF
C877 VPB.n199 VNB 0.02fF
C878 VPB.n200 VNB 0.02fF
C879 VPB.n202 VNB 0.02fF
C880 VPB.n203 VNB 0.02fF
C881 VPB.n204 VNB 0.02fF
C882 VPB.n206 VNB 0.28fF
C883 VPB.n208 VNB 0.03fF
C884 VPB.n209 VNB 0.02fF
C885 VPB.n210 VNB 0.03fF
C886 VPB.n211 VNB 0.03fF
C887 VPB.n212 VNB 0.28fF
C888 VPB.n213 VNB 0.01fF
C889 VPB.n214 VNB 0.02fF
C890 VPB.n215 VNB 0.04fF
C891 VPB.n216 VNB 0.28fF
C892 VPB.n217 VNB 0.02fF
C893 VPB.n218 VNB 0.02fF
C894 VPB.n219 VNB 0.02fF
C895 VPB.n220 VNB 0.28fF
C896 VPB.n221 VNB 0.02fF
C897 VPB.n222 VNB 0.02fF
C898 VPB.n223 VNB 0.02fF
C899 VPB.n224 VNB 0.28fF
C900 VPB.n225 VNB 0.02fF
C901 VPB.n226 VNB 0.02fF
C902 VPB.n227 VNB 0.02fF
C903 VPB.n228 VNB 0.28fF
C904 VPB.n229 VNB 0.02fF
C905 VPB.n230 VNB 0.02fF
C906 VPB.n231 VNB 0.02fF
C907 VPB.n232 VNB 0.28fF
C908 VPB.n233 VNB 0.02fF
C909 VPB.n234 VNB 0.02fF
C910 VPB.n235 VNB 0.02fF
C911 VPB.n236 VNB 0.28fF
C912 VPB.n237 VNB 0.02fF
C913 VPB.n238 VNB 0.02fF
C914 VPB.n239 VNB 0.02fF
C915 VPB.n240 VNB 0.28fF
C916 VPB.n241 VNB 0.01fF
C917 VPB.n242 VNB 0.02fF
C918 VPB.n243 VNB 0.04fF
C919 VPB.n244 VNB 0.02fF
C920 VPB.n245 VNB 0.02fF
C921 VPB.n246 VNB 0.02fF
C922 VPB.n247 VNB 0.04fF
C923 VPB.n248 VNB 0.02fF
C924 VPB.n249 VNB 0.20fF
C925 VPB.n250 VNB 0.04fF
C926 VPB.n252 VNB 0.02fF
C927 VPB.n253 VNB 0.02fF
C928 VPB.n254 VNB 0.02fF
C929 VPB.n255 VNB 0.02fF
C930 VPB.n257 VNB 0.02fF
C931 VPB.n258 VNB 0.02fF
C932 VPB.n259 VNB 0.02fF
C933 VPB.n261 VNB 0.28fF
C934 VPB.n263 VNB 0.03fF
C935 VPB.n264 VNB 0.02fF
C936 VPB.n265 VNB 0.03fF
C937 VPB.n266 VNB 0.03fF
C938 VPB.n267 VNB 0.28fF
C939 VPB.n268 VNB 0.01fF
C940 VPB.n269 VNB 0.02fF
C941 VPB.n270 VNB 0.04fF
C942 VPB.n271 VNB 0.28fF
C943 VPB.n272 VNB 0.02fF
C944 VPB.n273 VNB 0.02fF
C945 VPB.n274 VNB 0.02fF
C946 VPB.n275 VNB 0.28fF
C947 VPB.n276 VNB 0.02fF
C948 VPB.n277 VNB 0.02fF
C949 VPB.n278 VNB 0.02fF
C950 VPB.n279 VNB 0.28fF
C951 VPB.n280 VNB 0.02fF
C952 VPB.n281 VNB 0.02fF
C953 VPB.n282 VNB 0.02fF
C954 VPB.n283 VNB 0.28fF
C955 VPB.n284 VNB 0.02fF
C956 VPB.n285 VNB 0.02fF
C957 VPB.n286 VNB 0.02fF
C958 VPB.n287 VNB 0.28fF
C959 VPB.n288 VNB 0.02fF
C960 VPB.n289 VNB 0.02fF
C961 VPB.n290 VNB 0.02fF
C962 VPB.n291 VNB 0.28fF
C963 VPB.n292 VNB 0.02fF
C964 VPB.n293 VNB 0.02fF
C965 VPB.n294 VNB 0.02fF
C966 VPB.n295 VNB 0.28fF
C967 VPB.n296 VNB 0.01fF
C968 VPB.n297 VNB 0.02fF
C969 VPB.n298 VNB 0.04fF
C970 VPB.n299 VNB 0.02fF
C971 VPB.n300 VNB 0.02fF
C972 VPB.n301 VNB 0.02fF
C973 VPB.n302 VNB 0.04fF
C974 VPB.n303 VNB 0.02fF
C975 VPB.n304 VNB 0.20fF
C976 VPB.n305 VNB 0.04fF
C977 VPB.n307 VNB 0.02fF
C978 VPB.n308 VNB 0.02fF
C979 VPB.n309 VNB 0.02fF
C980 VPB.n310 VNB 0.02fF
C981 VPB.n312 VNB 0.02fF
C982 VPB.n313 VNB 0.02fF
C983 VPB.n314 VNB 0.02fF
C984 VPB.n316 VNB 0.28fF
C985 VPB.n318 VNB 0.03fF
C986 VPB.n319 VNB 0.02fF
C987 VPB.n320 VNB 0.03fF
C988 VPB.n321 VNB 0.03fF
C989 VPB.n322 VNB 0.28fF
C990 VPB.n323 VNB 0.01fF
C991 VPB.n324 VNB 0.02fF
C992 VPB.n325 VNB 0.04fF
C993 VPB.n326 VNB 0.06fF
C994 VPB.n327 VNB 0.24fF
C995 VPB.n328 VNB 0.02fF
C996 VPB.n329 VNB 0.01fF
C997 VPB.n330 VNB 0.02fF
C998 VPB.n331 VNB 0.14fF
C999 VPB.n332 VNB 0.16fF
C1000 VPB.n333 VNB 0.02fF
C1001 VPB.n334 VNB 0.02fF
C1002 VPB.n335 VNB 0.02fF
C1003 VPB.n336 VNB 0.10fF
C1004 VPB.n337 VNB 0.02fF
C1005 VPB.n338 VNB 0.14fF
C1006 VPB.n339 VNB 0.15fF
C1007 VPB.n340 VNB 0.02fF
C1008 VPB.n341 VNB 0.02fF
C1009 VPB.n342 VNB 0.02fF
C1010 VPB.n343 VNB 0.14fF
C1011 VPB.n344 VNB 0.15fF
C1012 VPB.n345 VNB 0.02fF
C1013 VPB.n346 VNB 0.02fF
C1014 VPB.n347 VNB 0.02fF
C1015 VPB.n348 VNB 0.14fF
C1016 VPB.n349 VNB 0.16fF
C1017 VPB.n350 VNB 0.02fF
C1018 VPB.n351 VNB 0.02fF
C1019 VPB.n352 VNB 0.02fF
C1020 VPB.n353 VNB 0.06fF
C1021 VPB.n354 VNB 0.24fF
C1022 VPB.n355 VNB 0.02fF
C1023 VPB.n356 VNB 0.01fF
C1024 VPB.n357 VNB 0.02fF
C1025 VPB.n358 VNB 0.28fF
C1026 VPB.n359 VNB 0.01fF
C1027 VPB.n360 VNB 0.02fF
C1028 VPB.n361 VNB 0.04fF
C1029 VPB.n362 VNB 0.02fF
C1030 VPB.n363 VNB 0.02fF
C1031 VPB.n364 VNB 0.02fF
C1032 VPB.n365 VNB 0.04fF
C1033 VPB.n366 VNB 0.02fF
C1034 VPB.n367 VNB 0.24fF
C1035 VPB.n368 VNB 0.04fF
C1036 VPB.n370 VNB 0.02fF
C1037 VPB.n371 VNB 0.02fF
C1038 VPB.n372 VNB 0.02fF
C1039 VPB.n373 VNB 0.02fF
C1040 VPB.n375 VNB 0.02fF
C1041 VPB.n376 VNB 0.02fF
C1042 VPB.n377 VNB 0.02fF
C1043 VPB.n379 VNB 0.28fF
C1044 VPB.n381 VNB 0.03fF
C1045 VPB.n382 VNB 0.02fF
C1046 VPB.n383 VNB 0.03fF
C1047 VPB.n384 VNB 0.03fF
C1048 VPB.n385 VNB 0.28fF
C1049 VPB.n386 VNB 0.01fF
C1050 VPB.n387 VNB 0.02fF
C1051 VPB.n388 VNB 0.04fF
C1052 VPB.n389 VNB 0.28fF
C1053 VPB.n390 VNB 0.02fF
C1054 VPB.n391 VNB 0.02fF
C1055 VPB.n392 VNB 0.02fF
C1056 VPB.n393 VNB 0.05fF
C1057 VPB.n394 VNB 0.21fF
C1058 VPB.n395 VNB 0.02fF
C1059 VPB.n396 VNB 0.01fF
C1060 VPB.n397 VNB 0.02fF
C1061 VPB.n398 VNB 0.14fF
C1062 VPB.n399 VNB 0.16fF
C1063 VPB.n400 VNB 0.02fF
C1064 VPB.n401 VNB 0.02fF
C1065 VPB.n402 VNB 0.02fF
C1066 VPB.n403 VNB 0.10fF
C1067 VPB.n404 VNB 0.02fF
C1068 VPB.n405 VNB 0.14fF
C1069 VPB.n406 VNB 0.16fF
C1070 VPB.n407 VNB 0.02fF
C1071 VPB.n408 VNB 0.02fF
C1072 VPB.n409 VNB 0.02fF
C1073 VPB.n410 VNB 0.14fF
C1074 VPB.n411 VNB 0.15fF
C1075 VPB.n412 VNB 0.02fF
C1076 VPB.n413 VNB 0.02fF
C1077 VPB.n414 VNB 0.02fF
C1078 VPB.n415 VNB 0.14fF
C1079 VPB.n416 VNB 0.15fF
C1080 VPB.n417 VNB 0.02fF
C1081 VPB.n418 VNB 0.02fF
C1082 VPB.n419 VNB 0.02fF
C1083 VPB.n420 VNB 0.10fF
C1084 VPB.n421 VNB 0.02fF
C1085 VPB.n422 VNB 0.14fF
C1086 VPB.n423 VNB 0.16fF
C1087 VPB.n424 VNB 0.02fF
C1088 VPB.n425 VNB 0.02fF
C1089 VPB.n426 VNB 0.02fF
C1090 VPB.n427 VNB 0.14fF
C1091 VPB.n428 VNB 0.16fF
C1092 VPB.n429 VNB 0.02fF
C1093 VPB.n430 VNB 0.02fF
C1094 VPB.n431 VNB 0.02fF
C1095 VPB.n432 VNB 0.06fF
C1096 VPB.n433 VNB 0.21fF
C1097 VPB.n434 VNB 0.02fF
C1098 VPB.n435 VNB 0.01fF
C1099 VPB.n436 VNB 0.02fF
C1100 VPB.n437 VNB 0.28fF
C1101 VPB.n438 VNB 0.02fF
C1102 VPB.n439 VNB 0.02fF
C1103 VPB.n440 VNB 0.02fF
C1104 VPB.n441 VNB 0.28fF
C1105 VPB.n442 VNB 0.01fF
C1106 VPB.n443 VNB 0.02fF
C1107 VPB.n444 VNB 0.04fF
C1108 VPB.n445 VNB 0.02fF
C1109 VPB.n446 VNB 0.02fF
C1110 VPB.n447 VNB 0.02fF
C1111 VPB.n448 VNB 0.04fF
C1112 VPB.n449 VNB 0.02fF
C1113 VPB.n450 VNB 0.29fF
C1114 VPB.n451 VNB 0.04fF
C1115 VPB.n453 VNB 0.02fF
C1116 VPB.n454 VNB 0.02fF
C1117 VPB.n455 VNB 0.02fF
C1118 VPB.n456 VNB 0.02fF
C1119 VPB.n458 VNB 0.02fF
C1120 VPB.n459 VNB 0.02fF
C1121 VPB.n460 VNB 0.02fF
C1122 VPB.n462 VNB 0.28fF
C1123 VPB.n464 VNB 0.03fF
C1124 VPB.n465 VNB 0.02fF
C1125 VPB.n466 VNB 0.03fF
C1126 VPB.n467 VNB 0.03fF
C1127 VPB.n468 VNB 0.28fF
C1128 VPB.n469 VNB 0.01fF
C1129 VPB.n470 VNB 0.02fF
C1130 VPB.n471 VNB 0.04fF
C1131 VPB.n472 VNB 0.28fF
C1132 VPB.n473 VNB 0.02fF
C1133 VPB.n474 VNB 0.02fF
C1134 VPB.n475 VNB 0.02fF
C1135 VPB.n476 VNB 0.05fF
C1136 VPB.n477 VNB 0.21fF
C1137 VPB.n478 VNB 0.02fF
C1138 VPB.n479 VNB 0.01fF
C1139 VPB.n480 VNB 0.02fF
C1140 VPB.n481 VNB 0.14fF
C1141 VPB.n482 VNB 0.16fF
C1142 VPB.n483 VNB 0.02fF
C1143 VPB.n484 VNB 0.02fF
C1144 VPB.n485 VNB 0.02fF
C1145 VPB.n486 VNB 0.10fF
C1146 VPB.n487 VNB 0.02fF
C1147 VPB.n488 VNB 0.14fF
C1148 VPB.n489 VNB 0.16fF
C1149 VPB.n490 VNB 0.02fF
C1150 VPB.n491 VNB 0.02fF
C1151 VPB.n492 VNB 0.02fF
C1152 VPB.n493 VNB 0.14fF
C1153 VPB.n494 VNB 0.15fF
C1154 VPB.n495 VNB 0.02fF
C1155 VPB.n496 VNB 0.02fF
C1156 VPB.n497 VNB 0.02fF
C1157 VPB.n498 VNB 0.14fF
C1158 VPB.n499 VNB 0.15fF
C1159 VPB.n500 VNB 0.02fF
C1160 VPB.n501 VNB 0.02fF
C1161 VPB.n502 VNB 0.02fF
C1162 VPB.n503 VNB 0.10fF
C1163 VPB.n504 VNB 0.02fF
C1164 VPB.n505 VNB 0.14fF
C1165 VPB.n506 VNB 0.16fF
C1166 VPB.n507 VNB 0.02fF
C1167 VPB.n508 VNB 0.02fF
C1168 VPB.n509 VNB 0.02fF
C1169 VPB.n510 VNB 0.14fF
C1170 VPB.n511 VNB 0.16fF
C1171 VPB.n512 VNB 0.02fF
C1172 VPB.n513 VNB 0.02fF
C1173 VPB.n514 VNB 0.02fF
C1174 VPB.n515 VNB 0.06fF
C1175 VPB.n516 VNB 0.21fF
C1176 VPB.n517 VNB 0.02fF
C1177 VPB.n518 VNB 0.01fF
C1178 VPB.n519 VNB 0.02fF
C1179 VPB.n520 VNB 0.28fF
C1180 VPB.n521 VNB 0.02fF
C1181 VPB.n522 VNB 0.02fF
C1182 VPB.n523 VNB 0.02fF
C1183 VPB.n524 VNB 0.28fF
C1184 VPB.n525 VNB 0.01fF
C1185 VPB.n526 VNB 0.02fF
C1186 VPB.n527 VNB 0.04fF
C1187 VPB.n528 VNB 0.02fF
C1188 VPB.n529 VNB 0.02fF
C1189 VPB.n530 VNB 0.02fF
C1190 VPB.n531 VNB 0.04fF
C1191 VPB.n532 VNB 0.02fF
C1192 VPB.n533 VNB 0.29fF
C1193 VPB.n534 VNB 0.04fF
C1194 VPB.n536 VNB 0.02fF
C1195 VPB.n537 VNB 0.02fF
C1196 VPB.n538 VNB 0.02fF
C1197 VPB.n539 VNB 0.02fF
C1198 VPB.n541 VNB 0.02fF
C1199 VPB.n542 VNB 0.02fF
C1200 VPB.n543 VNB 0.02fF
C1201 VPB.n545 VNB 0.28fF
C1202 VPB.n547 VNB 0.03fF
C1203 VPB.n548 VNB 0.02fF
C1204 VPB.n549 VNB 0.03fF
C1205 VPB.n550 VNB 0.03fF
C1206 VPB.n551 VNB 0.28fF
C1207 VPB.n552 VNB 0.01fF
C1208 VPB.n553 VNB 0.02fF
C1209 VPB.n554 VNB 0.04fF
C1210 VPB.n555 VNB 0.28fF
C1211 VPB.n556 VNB 0.02fF
C1212 VPB.n557 VNB 0.02fF
C1213 VPB.n558 VNB 0.02fF
C1214 VPB.n559 VNB 0.05fF
C1215 VPB.n560 VNB 0.21fF
C1216 VPB.n561 VNB 0.02fF
C1217 VPB.n562 VNB 0.01fF
C1218 VPB.n563 VNB 0.02fF
C1219 VPB.n564 VNB 0.14fF
C1220 VPB.n565 VNB 0.16fF
C1221 VPB.n566 VNB 0.02fF
C1222 VPB.n567 VNB 0.02fF
C1223 VPB.n568 VNB 0.02fF
C1224 VPB.n569 VNB 0.10fF
C1225 VPB.n570 VNB 0.02fF
C1226 VPB.n571 VNB 0.14fF
C1227 VPB.n572 VNB 0.16fF
C1228 VPB.n573 VNB 0.02fF
C1229 VPB.n574 VNB 0.02fF
C1230 VPB.n575 VNB 0.02fF
C1231 VPB.n576 VNB 0.14fF
C1232 VPB.n577 VNB 0.15fF
C1233 VPB.n578 VNB 0.02fF
C1234 VPB.n579 VNB 0.02fF
C1235 VPB.n580 VNB 0.02fF
C1236 VPB.n581 VNB 0.14fF
C1237 VPB.n582 VNB 0.15fF
C1238 VPB.n583 VNB 0.02fF
C1239 VPB.n584 VNB 0.02fF
C1240 VPB.n585 VNB 0.02fF
C1241 VPB.n586 VNB 0.10fF
C1242 VPB.n587 VNB 0.02fF
C1243 VPB.n588 VNB 0.14fF
C1244 VPB.n589 VNB 0.16fF
C1245 VPB.n590 VNB 0.02fF
C1246 VPB.n591 VNB 0.02fF
C1247 VPB.n592 VNB 0.02fF
C1248 VPB.n593 VNB 0.14fF
C1249 VPB.n594 VNB 0.16fF
C1250 VPB.n595 VNB 0.02fF
C1251 VPB.n596 VNB 0.02fF
C1252 VPB.n597 VNB 0.02fF
C1253 VPB.n598 VNB 0.06fF
C1254 VPB.n599 VNB 0.21fF
C1255 VPB.n600 VNB 0.02fF
C1256 VPB.n601 VNB 0.01fF
C1257 VPB.n602 VNB 0.02fF
C1258 VPB.n603 VNB 0.28fF
C1259 VPB.n604 VNB 0.02fF
C1260 VPB.n605 VNB 0.02fF
C1261 VPB.n606 VNB 0.02fF
C1262 VPB.n607 VNB 0.28fF
C1263 VPB.n608 VNB 0.01fF
C1264 VPB.n609 VNB 0.02fF
C1265 VPB.n610 VNB 0.04fF
C1266 VPB.n611 VNB 0.02fF
C1267 VPB.n612 VNB 0.02fF
C1268 VPB.n613 VNB 0.02fF
C1269 VPB.n614 VNB 0.04fF
C1270 VPB.n615 VNB 0.02fF
C1271 VPB.n616 VNB 0.29fF
C1272 VPB.n617 VNB 0.04fF
C1273 VPB.n619 VNB 0.02fF
C1274 VPB.n620 VNB 0.02fF
C1275 VPB.n621 VNB 0.02fF
C1276 VPB.n622 VNB 0.02fF
C1277 VPB.n624 VNB 0.02fF
C1278 VPB.n625 VNB 0.02fF
C1279 VPB.n626 VNB 0.02fF
C1280 VPB.n628 VNB 0.28fF
C1281 VPB.n630 VNB 0.03fF
C1282 VPB.n631 VNB 0.02fF
C1283 VPB.n632 VNB 0.03fF
C1284 VPB.n633 VNB 0.03fF
C1285 VPB.n634 VNB 0.28fF
C1286 VPB.n635 VNB 0.01fF
C1287 VPB.n636 VNB 0.02fF
C1288 VPB.n637 VNB 0.04fF
C1289 VPB.n638 VNB 0.28fF
C1290 VPB.n639 VNB 0.02fF
C1291 VPB.n640 VNB 0.02fF
C1292 VPB.n641 VNB 0.02fF
C1293 VPB.n642 VNB 0.05fF
C1294 VPB.n643 VNB 0.21fF
C1295 VPB.n644 VNB 0.02fF
C1296 VPB.n645 VNB 0.01fF
C1297 VPB.n646 VNB 0.02fF
C1298 VPB.n647 VNB 0.14fF
C1299 VPB.n648 VNB 0.16fF
C1300 VPB.n649 VNB 0.02fF
C1301 VPB.n650 VNB 0.02fF
C1302 VPB.n651 VNB 0.02fF
C1303 VPB.n652 VNB 0.10fF
C1304 VPB.n653 VNB 0.02fF
C1305 VPB.n654 VNB 0.14fF
C1306 VPB.n655 VNB 0.16fF
C1307 VPB.n656 VNB 0.02fF
C1308 VPB.n657 VNB 0.02fF
C1309 VPB.n658 VNB 0.02fF
C1310 VPB.n659 VNB 0.14fF
C1311 VPB.n660 VNB 0.15fF
C1312 VPB.n661 VNB 0.02fF
C1313 VPB.n662 VNB 0.02fF
C1314 VPB.n663 VNB 0.02fF
C1315 VPB.n664 VNB 0.14fF
C1316 VPB.n665 VNB 0.15fF
C1317 VPB.n666 VNB 0.02fF
C1318 VPB.n667 VNB 0.02fF
C1319 VPB.n668 VNB 0.02fF
C1320 VPB.n669 VNB 0.10fF
C1321 VPB.n670 VNB 0.02fF
C1322 VPB.n671 VNB 0.14fF
C1323 VPB.n672 VNB 0.16fF
C1324 VPB.n673 VNB 0.02fF
C1325 VPB.n674 VNB 0.02fF
C1326 VPB.n675 VNB 0.02fF
C1327 VPB.n676 VNB 0.14fF
C1328 VPB.n677 VNB 0.16fF
C1329 VPB.n678 VNB 0.02fF
C1330 VPB.n679 VNB 0.02fF
C1331 VPB.n680 VNB 0.02fF
C1332 VPB.n681 VNB 0.06fF
C1333 VPB.n682 VNB 0.21fF
C1334 VPB.n683 VNB 0.02fF
C1335 VPB.n684 VNB 0.01fF
C1336 VPB.n685 VNB 0.02fF
C1337 VPB.n686 VNB 0.28fF
C1338 VPB.n687 VNB 0.02fF
C1339 VPB.n688 VNB 0.02fF
C1340 VPB.n689 VNB 0.02fF
C1341 VPB.n690 VNB 0.28fF
C1342 VPB.n691 VNB 0.01fF
C1343 VPB.n692 VNB 0.02fF
C1344 VPB.n693 VNB 0.04fF
C1345 VPB.n694 VNB 0.02fF
C1346 VPB.n695 VNB 0.02fF
C1347 VPB.n696 VNB 0.02fF
C1348 VPB.n697 VNB 0.04fF
C1349 VPB.n698 VNB 0.02fF
C1350 VPB.n699 VNB 0.29fF
C1351 VPB.n700 VNB 0.04fF
C1352 VPB.n702 VNB 0.02fF
C1353 VPB.n703 VNB 0.02fF
C1354 VPB.n704 VNB 0.02fF
C1355 VPB.n705 VNB 0.02fF
C1356 VPB.n707 VNB 0.02fF
C1357 VPB.n708 VNB 0.02fF
C1358 VPB.n709 VNB 0.02fF
C1359 VPB.n711 VNB 0.28fF
C1360 VPB.n713 VNB 0.03fF
C1361 VPB.n714 VNB 0.02fF
C1362 VPB.n715 VNB 0.03fF
C1363 VPB.n716 VNB 0.03fF
C1364 VPB.n717 VNB 0.28fF
C1365 VPB.n718 VNB 0.01fF
C1366 VPB.n719 VNB 0.02fF
C1367 VPB.n720 VNB 0.04fF
C1368 VPB.n721 VNB 0.28fF
C1369 VPB.n722 VNB 0.02fF
C1370 VPB.n723 VNB 0.02fF
C1371 VPB.n724 VNB 0.02fF
C1372 VPB.n725 VNB 0.05fF
C1373 VPB.n726 VNB 0.21fF
C1374 VPB.n727 VNB 0.02fF
C1375 VPB.n728 VNB 0.01fF
C1376 VPB.n729 VNB 0.02fF
C1377 VPB.n730 VNB 0.14fF
C1378 VPB.n731 VNB 0.16fF
C1379 VPB.n732 VNB 0.02fF
C1380 VPB.n733 VNB 0.02fF
C1381 VPB.n734 VNB 0.02fF
C1382 VPB.n735 VNB 0.10fF
C1383 VPB.n736 VNB 0.02fF
C1384 VPB.n737 VNB 0.14fF
C1385 VPB.n738 VNB 0.16fF
C1386 VPB.n739 VNB 0.02fF
C1387 VPB.n740 VNB 0.02fF
C1388 VPB.n741 VNB 0.02fF
C1389 VPB.n742 VNB 0.14fF
C1390 VPB.n743 VNB 0.15fF
C1391 VPB.n744 VNB 0.02fF
C1392 VPB.n745 VNB 0.02fF
C1393 VPB.n746 VNB 0.02fF
C1394 VPB.n747 VNB 0.14fF
C1395 VPB.n748 VNB 0.15fF
C1396 VPB.n749 VNB 0.02fF
C1397 VPB.n750 VNB 0.02fF
C1398 VPB.n751 VNB 0.02fF
C1399 VPB.n752 VNB 0.10fF
C1400 VPB.n753 VNB 0.02fF
C1401 VPB.n754 VNB 0.14fF
C1402 VPB.n755 VNB 0.16fF
C1403 VPB.n756 VNB 0.02fF
C1404 VPB.n757 VNB 0.02fF
C1405 VPB.n758 VNB 0.02fF
C1406 VPB.n759 VNB 0.14fF
C1407 VPB.n760 VNB 0.16fF
C1408 VPB.n761 VNB 0.02fF
C1409 VPB.n762 VNB 0.02fF
C1410 VPB.n763 VNB 0.02fF
C1411 VPB.n764 VNB 0.06fF
C1412 VPB.n765 VNB 0.21fF
C1413 VPB.n766 VNB 0.02fF
C1414 VPB.n767 VNB 0.01fF
C1415 VPB.n768 VNB 0.02fF
C1416 VPB.n769 VNB 0.28fF
C1417 VPB.n770 VNB 0.02fF
C1418 VPB.n771 VNB 0.02fF
C1419 VPB.n772 VNB 0.02fF
C1420 VPB.n773 VNB 0.28fF
C1421 VPB.n774 VNB 0.01fF
C1422 VPB.n775 VNB 0.02fF
C1423 VPB.n776 VNB 0.04fF
C1424 VPB.n777 VNB 0.02fF
C1425 VPB.n778 VNB 0.02fF
C1426 VPB.n779 VNB 0.02fF
C1427 VPB.n780 VNB 0.04fF
C1428 VPB.n781 VNB 0.02fF
C1429 VPB.n782 VNB 0.29fF
C1430 VPB.n783 VNB 0.04fF
C1431 VPB.n785 VNB 0.02fF
C1432 VPB.n786 VNB 0.02fF
C1433 VPB.n787 VNB 0.02fF
C1434 VPB.n788 VNB 0.02fF
C1435 VPB.n790 VNB 0.02fF
C1436 VPB.n791 VNB 0.02fF
C1437 VPB.n792 VNB 0.02fF
C1438 VPB.n794 VNB 0.28fF
C1439 VPB.n796 VNB 0.03fF
C1440 VPB.n797 VNB 0.02fF
C1441 VPB.n798 VNB 0.03fF
C1442 VPB.n799 VNB 0.03fF
C1443 VPB.n800 VNB 0.28fF
C1444 VPB.n801 VNB 0.01fF
C1445 VPB.n802 VNB 0.02fF
C1446 VPB.n803 VNB 0.04fF
C1447 VPB.n804 VNB 0.28fF
C1448 VPB.n805 VNB 0.02fF
C1449 VPB.n806 VNB 0.02fF
C1450 VPB.n807 VNB 0.02fF
C1451 VPB.n808 VNB 0.05fF
C1452 VPB.n809 VNB 0.21fF
C1453 VPB.n810 VNB 0.02fF
C1454 VPB.n811 VNB 0.01fF
C1455 VPB.n812 VNB 0.02fF
C1456 VPB.n813 VNB 0.14fF
C1457 VPB.n814 VNB 0.16fF
C1458 VPB.n815 VNB 0.02fF
C1459 VPB.n816 VNB 0.02fF
C1460 VPB.n817 VNB 0.02fF
C1461 VPB.n818 VNB 0.10fF
C1462 VPB.n819 VNB 0.02fF
C1463 VPB.n820 VNB 0.14fF
C1464 VPB.n821 VNB 0.16fF
C1465 VPB.n822 VNB 0.02fF
C1466 VPB.n823 VNB 0.02fF
C1467 VPB.n824 VNB 0.02fF
C1468 VPB.n825 VNB 0.14fF
C1469 VPB.n826 VNB 0.15fF
C1470 VPB.n827 VNB 0.02fF
C1471 VPB.n828 VNB 0.02fF
C1472 VPB.n829 VNB 0.02fF
C1473 VPB.n830 VNB 0.14fF
C1474 VPB.n831 VNB 0.15fF
C1475 VPB.n832 VNB 0.02fF
C1476 VPB.n833 VNB 0.02fF
C1477 VPB.n834 VNB 0.02fF
C1478 VPB.n835 VNB 0.10fF
C1479 VPB.n836 VNB 0.02fF
C1480 VPB.n837 VNB 0.14fF
C1481 VPB.n838 VNB 0.16fF
C1482 VPB.n839 VNB 0.02fF
C1483 VPB.n840 VNB 0.02fF
C1484 VPB.n841 VNB 0.02fF
C1485 VPB.n842 VNB 0.14fF
C1486 VPB.n843 VNB 0.16fF
C1487 VPB.n844 VNB 0.02fF
C1488 VPB.n845 VNB 0.02fF
C1489 VPB.n846 VNB 0.02fF
C1490 VPB.n847 VNB 0.06fF
C1491 VPB.n848 VNB 0.21fF
C1492 VPB.n849 VNB 0.02fF
C1493 VPB.n850 VNB 0.01fF
C1494 VPB.n851 VNB 0.02fF
C1495 VPB.n852 VNB 0.28fF
C1496 VPB.n853 VNB 0.02fF
C1497 VPB.n854 VNB 0.02fF
C1498 VPB.n855 VNB 0.02fF
C1499 VPB.n856 VNB 0.28fF
C1500 VPB.n857 VNB 0.01fF
C1501 VPB.n858 VNB 0.02fF
C1502 VPB.n859 VNB 0.04fF
C1503 VPB.n860 VNB 0.02fF
C1504 VPB.n861 VNB 0.02fF
C1505 VPB.n862 VNB 0.02fF
C1506 VPB.n863 VNB 0.04fF
C1507 VPB.n864 VNB 0.02fF
C1508 VPB.n865 VNB 0.29fF
C1509 VPB.n866 VNB 0.04fF
C1510 VPB.n868 VNB 0.02fF
C1511 VPB.n869 VNB 0.02fF
C1512 VPB.n870 VNB 0.02fF
C1513 VPB.n871 VNB 0.02fF
C1514 VPB.n873 VNB 0.02fF
C1515 VPB.n874 VNB 0.02fF
C1516 VPB.n875 VNB 0.02fF
C1517 VPB.n877 VNB 0.28fF
C1518 VPB.n879 VNB 0.03fF
C1519 VPB.n880 VNB 0.02fF
C1520 VPB.n881 VNB 0.03fF
C1521 VPB.n882 VNB 0.03fF
C1522 VPB.n883 VNB 0.28fF
C1523 VPB.n884 VNB 0.01fF
C1524 VPB.n885 VNB 0.02fF
C1525 VPB.n886 VNB 0.04fF
C1526 VPB.n887 VNB 0.28fF
C1527 VPB.n888 VNB 0.02fF
C1528 VPB.n889 VNB 0.02fF
C1529 VPB.n890 VNB 0.02fF
C1530 VPB.n891 VNB 0.05fF
C1531 VPB.n892 VNB 0.21fF
C1532 VPB.n893 VNB 0.02fF
C1533 VPB.n894 VNB 0.01fF
C1534 VPB.n895 VNB 0.02fF
C1535 VPB.n896 VNB 0.14fF
C1536 VPB.n897 VNB 0.16fF
C1537 VPB.n898 VNB 0.02fF
C1538 VPB.n899 VNB 0.02fF
C1539 VPB.n900 VNB 0.02fF
C1540 VPB.n901 VNB 0.10fF
C1541 VPB.n902 VNB 0.02fF
C1542 VPB.n903 VNB 0.14fF
C1543 VPB.n904 VNB 0.16fF
C1544 VPB.n905 VNB 0.02fF
C1545 VPB.n906 VNB 0.02fF
C1546 VPB.n907 VNB 0.02fF
C1547 VPB.n908 VNB 0.14fF
C1548 VPB.n909 VNB 0.15fF
C1549 VPB.n910 VNB 0.02fF
C1550 VPB.n911 VNB 0.02fF
C1551 VPB.n912 VNB 0.02fF
C1552 VPB.n913 VNB 0.14fF
C1553 VPB.n914 VNB 0.15fF
C1554 VPB.n915 VNB 0.02fF
C1555 VPB.n916 VNB 0.02fF
C1556 VPB.n917 VNB 0.02fF
C1557 VPB.n918 VNB 0.10fF
C1558 VPB.n919 VNB 0.02fF
C1559 VPB.n920 VNB 0.14fF
C1560 VPB.n921 VNB 0.16fF
C1561 VPB.n922 VNB 0.02fF
C1562 VPB.n923 VNB 0.02fF
C1563 VPB.n924 VNB 0.02fF
C1564 VPB.n925 VNB 0.14fF
C1565 VPB.n926 VNB 0.16fF
C1566 VPB.n927 VNB 0.02fF
C1567 VPB.n928 VNB 0.02fF
C1568 VPB.n929 VNB 0.02fF
C1569 VPB.n930 VNB 0.06fF
C1570 VPB.n931 VNB 0.21fF
C1571 VPB.n932 VNB 0.02fF
C1572 VPB.n933 VNB 0.01fF
C1573 VPB.n934 VNB 0.02fF
C1574 VPB.n935 VNB 0.02fF
C1575 VPB.n936 VNB 0.04fF
C1576 VPB.n937 VNB 0.04fF
C1577 VPB.n938 VNB 0.02fF
C1578 VPB.n939 VNB 0.02fF
C1579 VPB.n940 VNB 0.02fF
C1580 VPB.n941 VNB 0.02fF
C1581 VPB.n942 VNB 0.02fF
C1582 VPB.n943 VNB 0.02fF
C1583 VPB.n944 VNB 0.02fF
C1584 VPB.n945 VNB 0.02fF
C1585 VPB.n946 VNB 0.14fF
C1586 VPB.n947 VNB 0.16fF
C1587 VPB.n948 VNB 0.02fF
C1588 VPB.n949 VNB 0.02fF
C1589 VPB.n950 VNB 0.06fF
C1590 VPB.n951 VNB 0.21fF
C1591 VPB.n952 VNB 0.02fF
C1592 VPB.n953 VNB 0.01fF
C1593 VPB.n954 VNB 0.02fF
C1594 VPB.n955 VNB 0.28fF
C1595 VPB.n956 VNB 0.02fF
C1596 VPB.n957 VNB 0.02fF
C1597 VPB.n958 VNB 0.02fF
C1598 VPB.n959 VNB 0.28fF
C1599 VPB.n960 VNB 0.01fF
C1600 VPB.n961 VNB 0.02fF
C1601 VPB.n962 VNB 0.04fF
C1602 VPB.n963 VNB 0.02fF
C1603 VPB.n964 VNB 0.02fF
C1604 VPB.n965 VNB 0.02fF
C1605 VPB.n966 VNB 0.04fF
C1606 VPB.n967 VNB 0.02fF
C1607 VPB.n968 VNB 0.29fF
C1608 VPB.n969 VNB 0.04fF
C1609 VPB.n971 VNB 0.02fF
C1610 VPB.n972 VNB 0.02fF
C1611 VPB.n973 VNB 0.02fF
C1612 VPB.n974 VNB 0.02fF
C1613 VPB.n976 VNB 0.02fF
C1614 VPB.n977 VNB 0.02fF
C1615 VPB.n978 VNB 0.02fF
C1616 VPB.n980 VNB 0.28fF
C1617 VPB.n982 VNB 0.03fF
C1618 VPB.n983 VNB 0.02fF
C1619 VPB.n984 VNB 0.03fF
C1620 VPB.n985 VNB 0.03fF
C1621 VPB.n986 VNB 0.28fF
C1622 VPB.n987 VNB 0.01fF
C1623 VPB.n988 VNB 0.02fF
C1624 VPB.n989 VNB 0.04fF
C1625 VPB.n990 VNB 0.28fF
C1626 VPB.n991 VNB 0.02fF
C1627 VPB.n992 VNB 0.02fF
C1628 VPB.n993 VNB 0.02fF
C1629 VPB.n994 VNB 0.05fF
C1630 VPB.n995 VNB 0.21fF
C1631 VPB.n996 VNB 0.02fF
C1632 VPB.n997 VNB 0.01fF
C1633 VPB.n998 VNB 0.02fF
C1634 VPB.n999 VNB 0.14fF
C1635 VPB.n1000 VNB 0.16fF
C1636 VPB.n1001 VNB 0.02fF
C1637 VPB.n1002 VNB 0.02fF
C1638 VPB.n1003 VNB 0.02fF
C1639 VPB.n1004 VNB 0.10fF
C1640 VPB.n1005 VNB 0.02fF
C1641 VPB.n1006 VNB 0.14fF
C1642 VPB.n1007 VNB 0.16fF
C1643 VPB.n1008 VNB 0.02fF
C1644 VPB.n1009 VNB 0.02fF
C1645 VPB.n1010 VNB 0.02fF
C1646 VPB.n1011 VNB 0.14fF
C1647 VPB.n1012 VNB 0.15fF
C1648 VPB.n1013 VNB 0.02fF
C1649 VPB.n1014 VNB 0.02fF
C1650 VPB.n1015 VNB 0.02fF
C1651 VPB.n1016 VNB 0.14fF
C1652 VPB.n1017 VNB 0.15fF
C1653 VPB.n1018 VNB 0.02fF
C1654 VPB.n1019 VNB 0.02fF
C1655 VPB.n1020 VNB 0.02fF
C1656 VPB.n1021 VNB 0.10fF
C1657 VPB.n1022 VNB 0.02fF
C1658 VPB.n1023 VNB 0.14fF
C1659 VPB.n1024 VNB 0.16fF
C1660 VPB.n1025 VNB 0.02fF
C1661 VPB.n1026 VNB 0.02fF
C1662 VPB.n1027 VNB 0.02fF
C1663 VPB.n1028 VNB 0.14fF
C1664 VPB.n1029 VNB 0.16fF
C1665 VPB.n1030 VNB 0.02fF
C1666 VPB.n1031 VNB 0.02fF
C1667 VPB.n1032 VNB 0.02fF
C1668 VPB.n1033 VNB 0.06fF
C1669 VPB.n1034 VNB 0.21fF
C1670 VPB.n1035 VNB 0.02fF
C1671 VPB.n1036 VNB 0.01fF
C1672 VPB.n1037 VNB 0.02fF
C1673 VPB.n1038 VNB 0.28fF
C1674 VPB.n1039 VNB 0.02fF
C1675 VPB.n1040 VNB 0.02fF
C1676 VPB.n1041 VNB 0.02fF
C1677 VPB.n1042 VNB 0.28fF
C1678 VPB.n1043 VNB 0.01fF
C1679 VPB.n1044 VNB 0.02fF
C1680 VPB.n1045 VNB 0.04fF
C1681 VPB.n1046 VNB 0.02fF
C1682 VPB.n1047 VNB 0.02fF
C1683 VPB.n1048 VNB 0.02fF
C1684 VPB.n1049 VNB 0.04fF
C1685 VPB.n1050 VNB 0.02fF
C1686 VPB.n1051 VNB 0.29fF
C1687 VPB.n1052 VNB 0.04fF
C1688 VPB.n1054 VNB 0.02fF
C1689 VPB.n1055 VNB 0.02fF
C1690 VPB.n1056 VNB 0.02fF
C1691 VPB.n1057 VNB 0.02fF
C1692 VPB.n1059 VNB 0.02fF
C1693 VPB.n1060 VNB 0.02fF
C1694 VPB.n1061 VNB 0.02fF
C1695 VPB.n1063 VNB 0.28fF
C1696 VPB.n1065 VNB 0.03fF
C1697 VPB.n1066 VNB 0.02fF
C1698 VPB.n1067 VNB 0.03fF
C1699 VPB.n1068 VNB 0.03fF
C1700 VPB.n1069 VNB 0.28fF
C1701 VPB.n1070 VNB 0.01fF
C1702 VPB.n1071 VNB 0.02fF
C1703 VPB.n1072 VNB 0.04fF
C1704 VPB.n1073 VNB 0.28fF
C1705 VPB.n1074 VNB 0.02fF
C1706 VPB.n1075 VNB 0.02fF
C1707 VPB.n1076 VNB 0.02fF
C1708 VPB.n1077 VNB 0.05fF
C1709 VPB.n1078 VNB 0.21fF
C1710 VPB.n1079 VNB 0.02fF
C1711 VPB.n1080 VNB 0.01fF
C1712 VPB.n1081 VNB 0.02fF
C1713 VPB.n1082 VNB 0.14fF
C1714 VPB.n1083 VNB 0.16fF
C1715 VPB.n1084 VNB 0.02fF
C1716 VPB.n1085 VNB 0.02fF
C1717 VPB.n1086 VNB 0.02fF
C1718 VPB.n1087 VNB 0.10fF
C1719 VPB.n1088 VNB 0.02fF
C1720 VPB.n1089 VNB 0.14fF
C1721 VPB.n1090 VNB 0.16fF
C1722 VPB.n1091 VNB 0.02fF
C1723 VPB.n1092 VNB 0.02fF
C1724 VPB.n1093 VNB 0.02fF
C1725 VPB.n1094 VNB 0.14fF
C1726 VPB.n1095 VNB 0.15fF
C1727 VPB.n1096 VNB 0.02fF
C1728 VPB.n1097 VNB 0.02fF
C1729 VPB.n1098 VNB 0.02fF
C1730 VPB.n1099 VNB 0.14fF
C1731 VPB.n1100 VNB 0.15fF
C1732 VPB.n1101 VNB 0.02fF
C1733 VPB.n1102 VNB 0.02fF
C1734 VPB.n1103 VNB 0.02fF
C1735 VPB.n1104 VNB 0.10fF
C1736 VPB.n1105 VNB 0.02fF
C1737 VPB.n1106 VNB 0.14fF
C1738 VPB.n1107 VNB 0.16fF
C1739 VPB.n1108 VNB 0.02fF
C1740 VPB.n1109 VNB 0.02fF
C1741 VPB.n1110 VNB 0.02fF
C1742 VPB.n1111 VNB 0.14fF
C1743 VPB.n1112 VNB 0.16fF
C1744 VPB.n1113 VNB 0.02fF
C1745 VPB.n1114 VNB 0.02fF
C1746 VPB.n1115 VNB 0.02fF
C1747 VPB.n1116 VNB 0.06fF
C1748 VPB.n1117 VNB 0.21fF
C1749 VPB.n1118 VNB 0.02fF
C1750 VPB.n1119 VNB 0.01fF
C1751 VPB.n1120 VNB 0.02fF
C1752 VPB.n1121 VNB 0.28fF
C1753 VPB.n1122 VNB 0.02fF
C1754 VPB.n1123 VNB 0.02fF
C1755 VPB.n1124 VNB 0.02fF
C1756 VPB.n1125 VNB 0.28fF
C1757 VPB.n1126 VNB 0.01fF
C1758 VPB.n1127 VNB 0.02fF
C1759 VPB.n1128 VNB 0.04fF
C1760 VPB.n1129 VNB 0.02fF
C1761 VPB.n1130 VNB 0.02fF
C1762 VPB.n1131 VNB 0.02fF
C1763 VPB.n1132 VNB 0.04fF
C1764 VPB.n1133 VNB 0.02fF
C1765 VPB.n1134 VNB 0.29fF
C1766 VPB.n1135 VNB 0.04fF
C1767 VPB.n1137 VNB 0.02fF
C1768 VPB.n1138 VNB 0.02fF
C1769 VPB.n1139 VNB 0.02fF
C1770 VPB.n1140 VNB 0.02fF
C1771 VPB.n1142 VNB 0.02fF
C1772 VPB.n1143 VNB 0.02fF
C1773 VPB.n1144 VNB 0.02fF
C1774 VPB.n1146 VNB 0.28fF
C1775 VPB.n1148 VNB 0.03fF
C1776 VPB.n1149 VNB 0.02fF
C1777 VPB.n1150 VNB 0.03fF
C1778 VPB.n1151 VNB 0.03fF
C1779 VPB.n1152 VNB 0.28fF
C1780 VPB.n1153 VNB 0.01fF
C1781 VPB.n1154 VNB 0.02fF
C1782 VPB.n1155 VNB 0.04fF
C1783 VPB.n1156 VNB 0.28fF
C1784 VPB.n1157 VNB 0.02fF
C1785 VPB.n1158 VNB 0.02fF
C1786 VPB.n1159 VNB 0.02fF
C1787 VPB.n1160 VNB 0.05fF
C1788 VPB.n1161 VNB 0.21fF
C1789 VPB.n1162 VNB 0.02fF
C1790 VPB.n1163 VNB 0.01fF
C1791 VPB.n1164 VNB 0.02fF
C1792 VPB.n1165 VNB 0.14fF
C1793 VPB.n1166 VNB 0.16fF
C1794 VPB.n1167 VNB 0.02fF
C1795 VPB.n1168 VNB 0.02fF
C1796 VPB.n1169 VNB 0.02fF
C1797 VPB.n1170 VNB 0.10fF
C1798 VPB.n1171 VNB 0.02fF
C1799 VPB.n1172 VNB 0.14fF
C1800 VPB.n1173 VNB 0.16fF
C1801 VPB.n1174 VNB 0.02fF
C1802 VPB.n1175 VNB 0.02fF
C1803 VPB.n1176 VNB 0.02fF
C1804 VPB.n1177 VNB 0.14fF
C1805 VPB.n1178 VNB 0.15fF
C1806 VPB.n1179 VNB 0.02fF
C1807 VPB.n1180 VNB 0.02fF
C1808 VPB.n1181 VNB 0.02fF
C1809 VPB.n1182 VNB 0.14fF
C1810 VPB.n1183 VNB 0.15fF
C1811 VPB.n1184 VNB 0.02fF
C1812 VPB.n1185 VNB 0.02fF
C1813 VPB.n1186 VNB 0.02fF
C1814 VPB.n1187 VNB 0.10fF
C1815 VPB.n1188 VNB 0.02fF
C1816 VPB.n1189 VNB 0.14fF
C1817 VPB.n1190 VNB 0.16fF
C1818 VPB.n1191 VNB 0.02fF
C1819 VPB.n1192 VNB 0.02fF
C1820 VPB.n1193 VNB 0.02fF
C1821 VPB.n1194 VNB 0.14fF
C1822 VPB.n1195 VNB 0.16fF
C1823 VPB.n1196 VNB 0.02fF
C1824 VPB.n1197 VNB 0.02fF
C1825 VPB.n1198 VNB 0.02fF
C1826 VPB.n1199 VNB 0.06fF
C1827 VPB.n1200 VNB 0.21fF
C1828 VPB.n1201 VNB 0.02fF
C1829 VPB.n1202 VNB 0.01fF
C1830 VPB.n1203 VNB 0.02fF
C1831 VPB.n1204 VNB 0.28fF
C1832 VPB.n1205 VNB 0.02fF
C1833 VPB.n1206 VNB 0.02fF
C1834 VPB.n1207 VNB 0.02fF
C1835 VPB.n1208 VNB 0.28fF
C1836 VPB.n1209 VNB 0.01fF
C1837 VPB.n1210 VNB 0.02fF
C1838 VPB.n1211 VNB 0.04fF
C1839 VPB.n1212 VNB 0.02fF
C1840 VPB.n1213 VNB 0.02fF
C1841 VPB.n1214 VNB 0.02fF
C1842 VPB.n1215 VNB 0.04fF
C1843 VPB.n1216 VNB 0.02fF
C1844 VPB.n1217 VNB 0.29fF
C1845 VPB.n1218 VNB 0.04fF
C1846 VPB.n1220 VNB 0.02fF
C1847 VPB.n1221 VNB 0.02fF
C1848 VPB.n1222 VNB 0.02fF
C1849 VPB.n1223 VNB 0.02fF
C1850 VPB.n1225 VNB 0.02fF
C1851 VPB.n1226 VNB 0.02fF
C1852 VPB.n1227 VNB 0.02fF
C1853 VPB.n1229 VNB 0.28fF
C1854 VPB.n1231 VNB 0.03fF
C1855 VPB.n1232 VNB 0.02fF
C1856 VPB.n1233 VNB 0.03fF
C1857 VPB.n1234 VNB 0.03fF
C1858 VPB.n1235 VNB 0.28fF
C1859 VPB.n1236 VNB 0.01fF
C1860 VPB.n1237 VNB 0.02fF
C1861 VPB.n1238 VNB 0.04fF
C1862 VPB.n1239 VNB 0.28fF
C1863 VPB.n1240 VNB 0.02fF
C1864 VPB.n1241 VNB 0.02fF
C1865 VPB.n1242 VNB 0.02fF
C1866 VPB.n1243 VNB 0.05fF
C1867 VPB.n1244 VNB 0.21fF
C1868 VPB.n1245 VNB 0.02fF
C1869 VPB.n1246 VNB 0.01fF
C1870 VPB.n1247 VNB 0.02fF
C1871 VPB.n1248 VNB 0.14fF
C1872 VPB.n1249 VNB 0.16fF
C1873 VPB.n1250 VNB 0.02fF
C1874 VPB.n1251 VNB 0.02fF
C1875 VPB.n1252 VNB 0.02fF
C1876 VPB.n1253 VNB 0.10fF
C1877 VPB.n1254 VNB 0.02fF
C1878 VPB.n1255 VNB 0.14fF
C1879 VPB.n1256 VNB 0.16fF
C1880 VPB.n1257 VNB 0.02fF
C1881 VPB.n1258 VNB 0.02fF
C1882 VPB.n1259 VNB 0.02fF
C1883 VPB.n1260 VNB 0.14fF
C1884 VPB.n1261 VNB 0.15fF
C1885 VPB.n1262 VNB 0.02fF
C1886 VPB.n1263 VNB 0.02fF
C1887 VPB.n1264 VNB 0.02fF
C1888 VPB.n1265 VNB 0.14fF
C1889 VPB.n1266 VNB 0.15fF
C1890 VPB.n1267 VNB 0.02fF
C1891 VPB.n1268 VNB 0.02fF
C1892 VPB.n1269 VNB 0.02fF
C1893 VPB.n1270 VNB 0.10fF
C1894 VPB.n1271 VNB 0.02fF
C1895 VPB.n1272 VNB 0.14fF
C1896 VPB.n1273 VNB 0.16fF
C1897 VPB.n1274 VNB 0.02fF
C1898 VPB.n1275 VNB 0.02fF
C1899 VPB.n1276 VNB 0.02fF
C1900 VPB.n1277 VNB 0.14fF
C1901 VPB.n1278 VNB 0.16fF
C1902 VPB.n1279 VNB 0.02fF
C1903 VPB.n1280 VNB 0.02fF
C1904 VPB.n1281 VNB 0.02fF
C1905 VPB.n1282 VNB 0.06fF
C1906 VPB.n1283 VNB 0.21fF
C1907 VPB.n1284 VNB 0.02fF
C1908 VPB.n1285 VNB 0.01fF
C1909 VPB.n1286 VNB 0.02fF
C1910 VPB.n1287 VNB 0.28fF
C1911 VPB.n1288 VNB 0.02fF
C1912 VPB.n1289 VNB 0.02fF
C1913 VPB.n1290 VNB 0.02fF
C1914 VPB.n1291 VNB 0.28fF
C1915 VPB.n1292 VNB 0.01fF
C1916 VPB.n1293 VNB 0.02fF
C1917 VPB.n1294 VNB 0.04fF
C1918 VPB.n1295 VNB 0.02fF
C1919 VPB.n1296 VNB 0.02fF
C1920 VPB.n1297 VNB 0.02fF
C1921 VPB.n1298 VNB 0.04fF
C1922 VPB.n1299 VNB 0.02fF
C1923 VPB.n1300 VNB 0.29fF
C1924 VPB.n1301 VNB 0.04fF
C1925 VPB.n1303 VNB 0.02fF
C1926 VPB.n1304 VNB 0.02fF
C1927 VPB.n1305 VNB 0.02fF
C1928 VPB.n1306 VNB 0.02fF
C1929 VPB.n1308 VNB 0.02fF
C1930 VPB.n1309 VNB 0.02fF
C1931 VPB.n1310 VNB 0.02fF
C1932 VPB.n1312 VNB 0.28fF
C1933 VPB.n1314 VNB 0.03fF
C1934 VPB.n1315 VNB 0.02fF
C1935 VPB.n1316 VNB 0.03fF
C1936 VPB.n1317 VNB 0.03fF
C1937 VPB.n1318 VNB 0.28fF
C1938 VPB.n1319 VNB 0.01fF
C1939 VPB.n1320 VNB 0.02fF
C1940 VPB.n1321 VNB 0.04fF
C1941 VPB.n1322 VNB 0.28fF
C1942 VPB.n1323 VNB 0.02fF
C1943 VPB.n1324 VNB 0.02fF
C1944 VPB.n1325 VNB 0.02fF
C1945 VPB.n1326 VNB 0.05fF
C1946 VPB.n1327 VNB 0.21fF
C1947 VPB.n1328 VNB 0.02fF
C1948 VPB.n1329 VNB 0.01fF
C1949 VPB.n1330 VNB 0.02fF
C1950 VPB.n1331 VNB 0.14fF
C1951 VPB.n1332 VNB 0.16fF
C1952 VPB.n1333 VNB 0.02fF
C1953 VPB.n1334 VNB 0.02fF
C1954 VPB.n1335 VNB 0.02fF
C1955 VPB.n1336 VNB 0.10fF
C1956 VPB.n1337 VNB 0.02fF
C1957 VPB.n1338 VNB 0.14fF
C1958 VPB.n1339 VNB 0.16fF
C1959 VPB.n1340 VNB 0.02fF
C1960 VPB.n1341 VNB 0.02fF
C1961 VPB.n1342 VNB 0.02fF
C1962 VPB.n1343 VNB 0.14fF
C1963 VPB.n1344 VNB 0.15fF
C1964 VPB.n1345 VNB 0.02fF
C1965 VPB.n1346 VNB 0.02fF
C1966 VPB.n1347 VNB 0.02fF
C1967 VPB.n1348 VNB 0.14fF
C1968 VPB.n1349 VNB 0.15fF
C1969 VPB.n1350 VNB 0.02fF
C1970 VPB.n1351 VNB 0.02fF
C1971 VPB.n1352 VNB 0.02fF
C1972 VPB.n1353 VNB 0.10fF
C1973 VPB.n1354 VNB 0.02fF
C1974 VPB.n1355 VNB 0.14fF
C1975 VPB.n1356 VNB 0.16fF
C1976 VPB.n1357 VNB 0.02fF
C1977 VPB.n1358 VNB 0.02fF
C1978 VPB.n1359 VNB 0.02fF
C1979 VPB.n1360 VNB 0.14fF
C1980 VPB.n1361 VNB 0.16fF
C1981 VPB.n1362 VNB 0.02fF
C1982 VPB.n1363 VNB 0.02fF
C1983 VPB.n1364 VNB 0.02fF
C1984 VPB.n1365 VNB 0.06fF
C1985 VPB.n1366 VNB 0.21fF
C1986 VPB.n1367 VNB 0.02fF
C1987 VPB.n1368 VNB 0.01fF
C1988 VPB.n1369 VNB 0.02fF
C1989 VPB.n1370 VNB 0.28fF
C1990 VPB.n1371 VNB 0.02fF
C1991 VPB.n1372 VNB 0.02fF
C1992 VPB.n1373 VNB 0.02fF
C1993 VPB.n1374 VNB 0.28fF
C1994 VPB.n1375 VNB 0.01fF
C1995 VPB.n1376 VNB 0.02fF
C1996 VPB.n1377 VNB 0.04fF
C1997 VPB.n1378 VNB 0.02fF
C1998 VPB.n1379 VNB 0.02fF
C1999 VPB.n1380 VNB 0.02fF
C2000 VPB.n1381 VNB 0.04fF
C2001 VPB.n1382 VNB 0.02fF
C2002 VPB.n1383 VNB 0.29fF
C2003 VPB.n1384 VNB 0.04fF
C2004 VPB.n1386 VNB 0.02fF
C2005 VPB.n1387 VNB 0.02fF
C2006 VPB.n1388 VNB 0.02fF
C2007 VPB.n1389 VNB 0.02fF
C2008 VPB.n1391 VNB 0.02fF
C2009 VPB.n1392 VNB 0.02fF
C2010 VPB.n1393 VNB 0.02fF
C2011 VPB.n1395 VNB 0.28fF
C2012 VPB.n1397 VNB 0.03fF
C2013 VPB.n1398 VNB 0.02fF
C2014 VPB.n1399 VNB 0.03fF
C2015 VPB.n1400 VNB 0.03fF
C2016 VPB.n1401 VNB 0.28fF
C2017 VPB.n1402 VNB 0.01fF
C2018 VPB.n1403 VNB 0.02fF
C2019 VPB.n1404 VNB 0.04fF
C2020 VPB.n1405 VNB 0.28fF
C2021 VPB.n1406 VNB 0.02fF
C2022 VPB.n1407 VNB 0.02fF
C2023 VPB.n1408 VNB 0.02fF
C2024 VPB.n1409 VNB 0.05fF
C2025 VPB.n1410 VNB 0.21fF
C2026 VPB.n1411 VNB 0.02fF
C2027 VPB.n1412 VNB 0.01fF
C2028 VPB.n1413 VNB 0.02fF
C2029 VPB.n1414 VNB 0.14fF
C2030 VPB.n1415 VNB 0.16fF
C2031 VPB.n1416 VNB 0.02fF
C2032 VPB.n1417 VNB 0.02fF
C2033 VPB.n1418 VNB 0.02fF
C2034 VPB.n1419 VNB 0.10fF
C2035 VPB.n1420 VNB 0.02fF
C2036 VPB.n1421 VNB 0.14fF
C2037 VPB.n1422 VNB 0.16fF
C2038 VPB.n1423 VNB 0.02fF
C2039 VPB.n1424 VNB 0.02fF
C2040 VPB.n1425 VNB 0.02fF
C2041 VPB.n1426 VNB 0.14fF
C2042 VPB.n1427 VNB 0.15fF
C2043 VPB.n1428 VNB 0.02fF
C2044 VPB.n1429 VNB 0.02fF
C2045 VPB.n1430 VNB 0.02fF
C2046 VPB.n1431 VNB 0.14fF
C2047 VPB.n1432 VNB 0.15fF
C2048 VPB.n1433 VNB 0.02fF
C2049 VPB.n1434 VNB 0.02fF
C2050 VPB.n1435 VNB 0.02fF
C2051 VPB.n1436 VNB 0.10fF
C2052 VPB.n1437 VNB 0.02fF
C2053 VPB.n1438 VNB 0.14fF
C2054 VPB.n1439 VNB 0.16fF
C2055 VPB.n1440 VNB 0.02fF
C2056 VPB.n1441 VNB 0.02fF
C2057 VPB.n1442 VNB 0.02fF
C2058 VPB.n1443 VNB 0.14fF
C2059 VPB.n1444 VNB 0.16fF
C2060 VPB.n1445 VNB 0.02fF
C2061 VPB.n1446 VNB 0.02fF
C2062 VPB.n1447 VNB 0.02fF
C2063 VPB.n1448 VNB 0.06fF
C2064 VPB.n1449 VNB 0.21fF
C2065 VPB.n1450 VNB 0.02fF
C2066 VPB.n1451 VNB 0.01fF
C2067 VPB.n1452 VNB 0.02fF
C2068 VPB.n1453 VNB 0.28fF
C2069 VPB.n1454 VNB 0.02fF
C2070 VPB.n1455 VNB 0.02fF
C2071 VPB.n1456 VNB 0.02fF
C2072 VPB.n1457 VNB 0.28fF
C2073 VPB.n1458 VNB 0.01fF
C2074 VPB.n1459 VNB 0.02fF
C2075 VPB.n1460 VNB 0.04fF
C2076 VPB.n1461 VNB 0.02fF
C2077 VPB.n1462 VNB 0.02fF
C2078 VPB.n1463 VNB 0.02fF
C2079 VPB.n1464 VNB 0.04fF
C2080 VPB.n1465 VNB 0.02fF
C2081 VPB.n1466 VNB 0.29fF
C2082 VPB.n1467 VNB 0.04fF
C2083 VPB.n1469 VNB 0.02fF
C2084 VPB.n1470 VNB 0.02fF
C2085 VPB.n1471 VNB 0.02fF
C2086 VPB.n1472 VNB 0.02fF
C2087 VPB.n1474 VNB 0.02fF
C2088 VPB.n1475 VNB 0.02fF
C2089 VPB.n1476 VNB 0.02fF
C2090 VPB.n1478 VNB 0.28fF
C2091 VPB.n1480 VNB 0.03fF
C2092 VPB.n1481 VNB 0.02fF
C2093 VPB.n1482 VNB 0.03fF
C2094 VPB.n1483 VNB 0.03fF
C2095 VPB.n1484 VNB 0.28fF
C2096 VPB.n1485 VNB 0.01fF
C2097 VPB.n1486 VNB 0.02fF
C2098 VPB.n1487 VNB 0.04fF
C2099 VPB.n1488 VNB 0.28fF
C2100 VPB.n1489 VNB 0.02fF
C2101 VPB.n1490 VNB 0.02fF
C2102 VPB.n1491 VNB 0.02fF
C2103 VPB.n1492 VNB 0.05fF
C2104 VPB.n1493 VNB 0.21fF
C2105 VPB.n1494 VNB 0.02fF
C2106 VPB.n1495 VNB 0.01fF
C2107 VPB.n1496 VNB 0.02fF
C2108 VPB.n1497 VNB 0.14fF
C2109 VPB.n1498 VNB 0.16fF
C2110 VPB.n1499 VNB 0.02fF
C2111 VPB.n1500 VNB 0.02fF
C2112 VPB.n1501 VNB 0.02fF
C2113 VPB.n1502 VNB 0.10fF
C2114 VPB.n1503 VNB 0.02fF
C2115 VPB.n1504 VNB 0.14fF
C2116 VPB.n1505 VNB 0.16fF
C2117 VPB.n1506 VNB 0.02fF
C2118 VPB.n1507 VNB 0.02fF
C2119 VPB.n1508 VNB 0.02fF
C2120 VPB.n1509 VNB 0.14fF
C2121 VPB.n1510 VNB 0.15fF
C2122 VPB.n1511 VNB 0.02fF
C2123 VPB.n1512 VNB 0.02fF
C2124 VPB.n1513 VNB 0.02fF
C2125 VPB.n1514 VNB 0.14fF
C2126 VPB.n1515 VNB 0.15fF
C2127 VPB.n1516 VNB 0.02fF
C2128 VPB.n1517 VNB 0.02fF
C2129 VPB.n1518 VNB 0.02fF
C2130 VPB.n1519 VNB 0.10fF
C2131 VPB.n1520 VNB 0.02fF
C2132 VPB.n1521 VNB 0.14fF
C2133 VPB.n1522 VNB 0.16fF
C2134 VPB.n1523 VNB 0.02fF
C2135 VPB.n1524 VNB 0.02fF
C2136 VPB.n1525 VNB 0.02fF
C2137 VPB.n1526 VNB 0.14fF
C2138 VPB.n1527 VNB 0.16fF
C2139 VPB.n1528 VNB 0.02fF
C2140 VPB.n1529 VNB 0.02fF
C2141 VPB.n1530 VNB 0.02fF
C2142 VPB.n1531 VNB 0.06fF
C2143 VPB.n1532 VNB 0.21fF
C2144 VPB.n1533 VNB 0.02fF
C2145 VPB.n1534 VNB 0.01fF
C2146 VPB.n1535 VNB 0.02fF
C2147 VPB.n1536 VNB 0.28fF
C2148 VPB.n1537 VNB 0.02fF
C2149 VPB.n1538 VNB 0.02fF
C2150 VPB.n1539 VNB 0.02fF
C2151 VPB.n1540 VNB 0.28fF
C2152 VPB.n1541 VNB 0.01fF
C2153 VPB.n1542 VNB 0.02fF
C2154 VPB.n1543 VNB 0.04fF
C2155 VPB.n1544 VNB 0.02fF
C2156 VPB.n1545 VNB 0.02fF
C2157 VPB.n1546 VNB 0.02fF
C2158 VPB.n1547 VNB 0.04fF
C2159 VPB.n1548 VNB 0.02fF
C2160 VPB.n1549 VNB 0.29fF
C2161 VPB.n1550 VNB 0.04fF
C2162 VPB.n1552 VNB 0.02fF
C2163 VPB.n1553 VNB 0.02fF
C2164 VPB.n1554 VNB 0.02fF
C2165 VPB.n1555 VNB 0.02fF
C2166 VPB.n1557 VNB 0.02fF
C2167 VPB.n1558 VNB 0.02fF
C2168 VPB.n1559 VNB 0.02fF
C2169 VPB.n1561 VNB 0.28fF
C2170 VPB.n1563 VNB 0.03fF
C2171 VPB.n1564 VNB 0.02fF
C2172 VPB.n1565 VNB 0.03fF
C2173 VPB.n1566 VNB 0.03fF
C2174 VPB.n1567 VNB 0.28fF
C2175 VPB.n1568 VNB 0.01fF
C2176 VPB.n1569 VNB 0.02fF
C2177 VPB.n1570 VNB 0.04fF
C2178 VPB.n1571 VNB 0.28fF
C2179 VPB.n1572 VNB 0.02fF
C2180 VPB.n1573 VNB 0.02fF
C2181 VPB.n1574 VNB 0.02fF
C2182 VPB.n1575 VNB 0.05fF
C2183 VPB.n1576 VNB 0.21fF
C2184 VPB.n1577 VNB 0.02fF
C2185 VPB.n1578 VNB 0.01fF
C2186 VPB.n1579 VNB 0.02fF
C2187 VPB.n1580 VNB 0.14fF
C2188 VPB.n1581 VNB 0.16fF
C2189 VPB.n1582 VNB 0.02fF
C2190 VPB.n1583 VNB 0.02fF
C2191 VPB.n1584 VNB 0.02fF
C2192 VPB.n1585 VNB 0.10fF
C2193 VPB.n1586 VNB 0.02fF
C2194 VPB.n1587 VNB 0.14fF
C2195 VPB.n1588 VNB 0.16fF
C2196 VPB.n1589 VNB 0.02fF
C2197 VPB.n1590 VNB 0.02fF
C2198 VPB.n1591 VNB 0.02fF
C2199 VPB.n1592 VNB 0.14fF
C2200 VPB.n1593 VNB 0.15fF
C2201 VPB.n1594 VNB 0.02fF
C2202 VPB.n1595 VNB 0.02fF
C2203 VPB.n1596 VNB 0.02fF
C2204 VPB.n1597 VNB 0.14fF
C2205 VPB.n1598 VNB 0.15fF
C2206 VPB.n1599 VNB 0.02fF
C2207 VPB.n1600 VNB 0.02fF
C2208 VPB.n1601 VNB 0.02fF
C2209 VPB.n1602 VNB 0.10fF
C2210 VPB.n1603 VNB 0.02fF
C2211 VPB.n1604 VNB 0.14fF
C2212 VPB.n1605 VNB 0.16fF
C2213 VPB.n1606 VNB 0.02fF
C2214 VPB.n1607 VNB 0.02fF
C2215 VPB.n1608 VNB 0.02fF
C2216 VPB.n1609 VNB 0.14fF
C2217 VPB.n1610 VNB 0.16fF
C2218 VPB.n1611 VNB 0.02fF
C2219 VPB.n1612 VNB 0.02fF
C2220 VPB.n1613 VNB 0.02fF
C2221 VPB.n1614 VNB 0.06fF
C2222 VPB.n1615 VNB 0.21fF
C2223 VPB.n1616 VNB 0.02fF
C2224 VPB.n1617 VNB 0.01fF
C2225 VPB.n1618 VNB 0.02fF
C2226 VPB.n1619 VNB 0.28fF
C2227 VPB.n1620 VNB 0.02fF
C2228 VPB.n1621 VNB 0.02fF
C2229 VPB.n1622 VNB 0.02fF
C2230 VPB.n1623 VNB 0.28fF
C2231 VPB.n1624 VNB 0.01fF
C2232 VPB.n1625 VNB 0.02fF
C2233 VPB.n1626 VNB 0.04fF
C2234 VPB.n1627 VNB 0.02fF
C2235 VPB.n1628 VNB 0.02fF
C2236 VPB.n1629 VNB 0.02fF
C2237 VPB.n1630 VNB 0.04fF
C2238 VPB.n1631 VNB 0.02fF
C2239 VPB.n1632 VNB 0.29fF
C2240 VPB.n1633 VNB 0.04fF
C2241 VPB.n1635 VNB 0.02fF
C2242 VPB.n1636 VNB 0.02fF
C2243 VPB.n1637 VNB 0.02fF
C2244 VPB.n1638 VNB 0.02fF
C2245 VPB.n1640 VNB 0.02fF
C2246 VPB.n1641 VNB 0.02fF
C2247 VPB.n1642 VNB 0.02fF
C2248 VPB.n1644 VNB 0.28fF
C2249 VPB.n1646 VNB 0.03fF
C2250 VPB.n1647 VNB 0.02fF
C2251 VPB.n1648 VNB 0.03fF
C2252 VPB.n1649 VNB 0.03fF
C2253 VPB.n1650 VNB 0.28fF
C2254 VPB.n1651 VNB 0.01fF
C2255 VPB.n1652 VNB 0.02fF
C2256 VPB.n1653 VNB 0.04fF
C2257 VPB.n1654 VNB 0.28fF
C2258 VPB.n1655 VNB 0.02fF
C2259 VPB.n1656 VNB 0.02fF
C2260 VPB.n1657 VNB 0.02fF
C2261 VPB.n1658 VNB 0.05fF
C2262 VPB.n1659 VNB 0.21fF
C2263 VPB.n1660 VNB 0.02fF
C2264 VPB.n1661 VNB 0.01fF
C2265 VPB.n1662 VNB 0.02fF
C2266 VPB.n1663 VNB 0.14fF
C2267 VPB.n1664 VNB 0.16fF
C2268 VPB.n1665 VNB 0.02fF
C2269 VPB.n1666 VNB 0.02fF
C2270 VPB.n1667 VNB 0.02fF
C2271 VPB.n1668 VNB 0.10fF
C2272 VPB.n1669 VNB 0.02fF
C2273 VPB.n1670 VNB 0.14fF
C2274 VPB.n1671 VNB 0.16fF
C2275 VPB.n1672 VNB 0.02fF
C2276 VPB.n1673 VNB 0.02fF
C2277 VPB.n1674 VNB 0.02fF
C2278 VPB.n1675 VNB 0.14fF
C2279 VPB.n1676 VNB 0.15fF
C2280 VPB.n1677 VNB 0.02fF
C2281 VPB.n1678 VNB 0.02fF
C2282 VPB.n1679 VNB 0.02fF
C2283 VPB.n1680 VNB 0.14fF
C2284 VPB.n1681 VNB 0.15fF
C2285 VPB.n1682 VNB 0.02fF
C2286 VPB.n1683 VNB 0.02fF
C2287 VPB.n1684 VNB 0.02fF
C2288 VPB.n1685 VNB 0.10fF
C2289 VPB.n1686 VNB 0.02fF
C2290 VPB.n1687 VNB 0.14fF
C2291 VPB.n1688 VNB 0.16fF
C2292 VPB.n1689 VNB 0.02fF
C2293 VPB.n1690 VNB 0.02fF
C2294 VPB.n1691 VNB 0.02fF
C2295 VPB.n1692 VNB 0.14fF
C2296 VPB.n1693 VNB 0.16fF
C2297 VPB.n1694 VNB 0.02fF
C2298 VPB.n1695 VNB 0.02fF
C2299 VPB.n1696 VNB 0.02fF
C2300 VPB.n1697 VNB 0.06fF
C2301 VPB.n1698 VNB 0.21fF
C2302 VPB.n1699 VNB 0.02fF
C2303 VPB.n1700 VNB 0.01fF
C2304 VPB.n1701 VNB 0.02fF
C2305 VPB.n1702 VNB 0.28fF
C2306 VPB.n1703 VNB 0.02fF
C2307 VPB.n1704 VNB 0.02fF
C2308 VPB.n1705 VNB 0.02fF
C2309 VPB.n1706 VNB 0.28fF
C2310 VPB.n1707 VNB 0.01fF
C2311 VPB.n1708 VNB 0.02fF
C2312 VPB.n1709 VNB 0.04fF
C2313 VPB.n1710 VNB 0.04fF
C2314 VPB.n1711 VNB 0.02fF
C2315 VPB.n1712 VNB 0.02fF
C2316 VPB.n1713 VNB 0.02fF
C2317 VPB.n1714 VNB 0.02fF
C2318 VPB.n1715 VNB 0.02fF
C2319 VPB.n1716 VNB 0.02fF
C2320 VPB.n1717 VNB 0.02fF
C2321 VPB.n1718 VNB 0.02fF
C2322 VPB.n1719 VNB 0.02fF
C2323 VPB.n1720 VNB 0.02fF
C2324 VPB.n1721 VNB 0.03fF
C2325 VPB.n1722 VNB 0.04fF
C2326 VPB.n1723 VNB 0.02fF
C2327 VPB.n1724 VNB 0.02fF
C2328 VPB.n1725 VNB 0.02fF
C2329 VPB.n1726 VNB 0.04fF
C2330 VPB.n1727 VNB 0.04fF
C2331 VPB.n1729 VNB 0.43fF
.ends
