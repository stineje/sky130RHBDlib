VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFQX1
  CLASS CORE ;
  FOREIGN DFFQX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.460 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 19.275 5.285 19.445 7.020 ;
        RECT 20.155 5.285 20.325 7.020 ;
        RECT 19.275 5.115 20.805 5.285 ;
        RECT 16.595 4.710 16.765 4.865 ;
        RECT 16.565 4.535 16.765 4.710 ;
        RECT 16.565 1.915 16.735 4.535 ;
        RECT 20.635 1.740 20.805 5.115 ;
        RECT 20.195 1.570 20.805 1.740 ;
        RECT 20.195 0.835 20.365 1.570 ;
      LAYER mcon ;
        RECT 16.565 3.615 16.735 3.785 ;
        RECT 20.635 3.615 20.805 3.785 ;
      LAYER met1 ;
        RECT 16.535 3.785 16.765 3.815 ;
        RECT 20.605 3.785 20.835 3.815 ;
        RECT 16.505 3.615 20.865 3.785 ;
        RECT 16.535 3.585 16.765 3.615 ;
        RECT 20.605 3.585 20.835 3.615 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 6.605 4.710 6.775 4.865 ;
        RECT 6.575 4.535 6.775 4.710 ;
        RECT 6.575 1.915 6.745 4.535 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 13.265 4.710 13.435 4.865 ;
        RECT 13.235 4.535 13.435 4.710 ;
        RECT 13.235 1.915 13.405 4.535 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 13.235 4.355 13.405 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 13.205 4.525 13.435 4.555 ;
        RECT 2.075 4.355 13.465 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 13.205 4.325 13.435 4.355 ;
    END
  END CLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 21.895 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 21.630 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.515 5.135 5.685 7.230 ;
        RECT 6.395 5.555 6.565 7.230 ;
        RECT 7.275 5.555 7.445 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 8.845 5.135 9.015 7.230 ;
        RECT 9.725 5.555 9.895 7.230 ;
        RECT 10.605 5.555 10.775 7.230 ;
        RECT 11.300 4.110 11.640 7.230 ;
        RECT 12.175 5.135 12.345 7.230 ;
        RECT 13.055 5.555 13.225 7.230 ;
        RECT 13.935 5.555 14.105 7.230 ;
        RECT 14.630 4.110 14.970 7.230 ;
        RECT 15.505 5.135 15.675 7.230 ;
        RECT 16.385 5.555 16.555 7.230 ;
        RECT 17.265 5.555 17.435 7.230 ;
        RECT 17.960 4.110 18.300 7.230 ;
        RECT 18.835 5.135 19.005 7.230 ;
        RECT 19.715 5.555 19.885 7.230 ;
        RECT 20.595 5.555 20.765 7.230 ;
        RECT 21.290 4.110 21.630 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 21.630 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 21.630 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.905 0.170 6.075 1.120 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.235 0.170 9.405 1.120 ;
        RECT 11.300 0.170 11.640 2.720 ;
        RECT 12.565 0.170 12.735 1.120 ;
        RECT 14.630 0.170 14.970 2.720 ;
        RECT 15.895 0.170 16.065 1.120 ;
        RECT 17.960 0.170 18.300 2.720 ;
        RECT 19.225 0.170 19.395 1.120 ;
        RECT 21.290 0.170 21.630 2.720 ;
        RECT -0.170 -0.170 21.630 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 21.630 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 5.955 5.285 6.125 7.020 ;
        RECT 6.835 5.285 7.005 7.020 ;
        RECT 9.285 5.285 9.455 7.020 ;
        RECT 10.165 5.285 10.335 7.020 ;
        RECT 12.615 5.285 12.785 7.020 ;
        RECT 13.495 5.285 13.665 7.020 ;
        RECT 15.945 5.285 16.115 7.020 ;
        RECT 16.825 5.285 16.995 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 5.955 5.115 7.485 5.285 ;
        RECT 9.285 5.115 10.815 5.285 ;
        RECT 12.615 5.115 14.145 5.285 ;
        RECT 15.945 5.115 17.475 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.420 1.665 5.590 1.745 ;
        RECT 6.390 1.665 6.560 1.745 ;
        RECT 7.315 1.740 7.485 5.115 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 9.935 4.710 10.105 4.865 ;
        RECT 9.905 4.535 10.105 4.710 ;
        RECT 9.905 1.915 10.075 4.535 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.420 1.495 6.560 1.665 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.420 0.365 5.590 1.495 ;
        RECT 6.390 0.615 6.560 1.495 ;
        RECT 6.875 1.570 7.485 1.740 ;
        RECT 8.750 1.665 8.920 1.745 ;
        RECT 9.720 1.665 9.890 1.745 ;
        RECT 10.645 1.740 10.815 5.115 ;
        RECT 12.495 1.915 12.665 4.865 ;
        RECT 6.875 0.835 7.045 1.570 ;
        RECT 8.750 1.495 9.890 1.665 ;
        RECT 7.360 0.615 7.530 1.385 ;
        RECT 6.390 0.445 7.530 0.615 ;
        RECT 6.390 0.365 6.560 0.445 ;
        RECT 7.360 0.365 7.530 0.445 ;
        RECT 8.750 0.365 8.920 1.495 ;
        RECT 9.720 0.615 9.890 1.495 ;
        RECT 10.205 1.570 10.815 1.740 ;
        RECT 12.080 1.665 12.250 1.745 ;
        RECT 13.050 1.665 13.220 1.745 ;
        RECT 13.975 1.740 14.145 5.115 ;
        RECT 15.825 1.915 15.995 4.865 ;
        RECT 10.205 0.835 10.375 1.570 ;
        RECT 12.080 1.495 13.220 1.665 ;
        RECT 10.690 0.615 10.860 1.385 ;
        RECT 9.720 0.445 10.860 0.615 ;
        RECT 9.720 0.365 9.890 0.445 ;
        RECT 10.690 0.365 10.860 0.445 ;
        RECT 12.080 0.365 12.250 1.495 ;
        RECT 13.050 0.615 13.220 1.495 ;
        RECT 13.535 1.570 14.145 1.740 ;
        RECT 15.410 1.665 15.580 1.745 ;
        RECT 16.380 1.665 16.550 1.745 ;
        RECT 17.305 1.740 17.475 5.115 ;
        RECT 19.155 1.915 19.325 4.865 ;
        RECT 19.925 4.710 20.095 4.865 ;
        RECT 19.895 4.535 20.095 4.710 ;
        RECT 19.895 1.915 20.065 4.535 ;
        RECT 13.535 0.835 13.705 1.570 ;
        RECT 15.410 1.495 16.550 1.665 ;
        RECT 14.020 0.615 14.190 1.385 ;
        RECT 13.050 0.445 14.190 0.615 ;
        RECT 13.050 0.365 13.220 0.445 ;
        RECT 14.020 0.365 14.190 0.445 ;
        RECT 15.410 0.365 15.580 1.495 ;
        RECT 16.380 0.615 16.550 1.495 ;
        RECT 16.865 1.570 17.475 1.740 ;
        RECT 18.740 1.665 18.910 1.745 ;
        RECT 19.710 1.665 19.880 1.745 ;
        RECT 16.865 0.835 17.035 1.570 ;
        RECT 18.740 1.495 19.880 1.665 ;
        RECT 17.350 0.615 17.520 1.385 ;
        RECT 16.380 0.445 17.520 0.615 ;
        RECT 16.380 0.365 16.550 0.445 ;
        RECT 17.350 0.365 17.520 0.445 ;
        RECT 18.740 0.365 18.910 1.495 ;
        RECT 19.710 0.615 19.880 1.495 ;
        RECT 20.680 0.615 20.850 1.385 ;
        RECT 19.710 0.445 20.850 0.615 ;
        RECT 19.710 0.365 19.880 0.445 ;
        RECT 20.680 0.365 20.850 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 7.315 3.245 7.485 3.415 ;
        RECT 9.165 3.245 9.335 3.415 ;
        RECT 9.905 3.985 10.075 4.155 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 12.495 3.245 12.665 3.415 ;
        RECT 13.975 3.985 14.145 4.155 ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 17.305 3.245 17.475 3.415 ;
        RECT 19.155 3.245 19.325 3.415 ;
        RECT 19.895 3.985 20.065 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 9.875 4.155 10.105 4.185 ;
        RECT 13.945 4.155 14.175 4.185 ;
        RECT 19.865 4.155 20.095 4.185 ;
        RECT 0.965 3.985 20.125 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 9.875 3.955 10.105 3.985 ;
        RECT 13.945 3.955 14.175 3.985 ;
        RECT 19.865 3.955 20.095 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 3.925 3.615 16.055 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 7.285 3.415 7.515 3.445 ;
        RECT 9.135 3.415 9.365 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.465 3.415 12.695 3.445 ;
        RECT 17.275 3.415 17.505 3.445 ;
        RECT 19.125 3.415 19.355 3.445 ;
        RECT 3.185 3.245 9.395 3.415 ;
        RECT 10.585 3.245 12.725 3.415 ;
        RECT 17.245 3.245 19.385 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 7.285 3.215 7.515 3.245 ;
        RECT 9.135 3.215 9.365 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.465 3.215 12.695 3.245 ;
        RECT 17.275 3.215 17.505 3.245 ;
        RECT 19.125 3.215 19.355 3.245 ;
  END
END DFFQX1
END LIBRARY

