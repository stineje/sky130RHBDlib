VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO TMRDFFQNX1
  CLASS CORE ;
  FOREIGN TMRDFFQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 74.370 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.734950 ;
    PORT
      LAYER li1 ;
        RECT 72.185 5.295 72.355 6.565 ;
        RECT 73.065 5.295 73.235 6.565 ;
        RECT 72.185 5.125 73.715 5.295 ;
        RECT 73.545 1.730 73.715 5.125 ;
        RECT 73.105 1.560 73.715 1.730 ;
        RECT 66.445 1.170 66.615 1.345 ;
        RECT 66.440 1.015 66.615 1.170 ;
        RECT 66.440 0.835 66.610 1.015 ;
        RECT 69.775 0.835 69.945 1.345 ;
        RECT 73.105 0.835 73.275 1.560 ;
      LAYER mcon ;
        RECT 66.445 1.095 66.615 1.265 ;
        RECT 69.775 1.095 69.945 1.265 ;
        RECT 73.105 1.095 73.275 1.265 ;
      LAYER met1 ;
        RECT 66.415 1.265 66.645 1.295 ;
        RECT 69.745 1.265 69.975 1.295 ;
        RECT 73.075 1.265 73.305 1.295 ;
        RECT 66.385 1.095 73.335 1.265 ;
        RECT 66.415 1.065 66.645 1.095 ;
        RECT 69.745 1.065 69.975 1.095 ;
        RECT 73.075 1.065 73.305 1.095 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.081750 ;
    PORT
      LAYER li1 ;
        RECT 6.605 4.710 6.775 4.865 ;
        RECT 28.065 4.710 28.235 4.865 ;
        RECT 49.525 4.710 49.695 4.865 ;
        RECT 6.575 4.535 6.775 4.710 ;
        RECT 28.035 4.535 28.235 4.710 ;
        RECT 49.495 4.535 49.695 4.710 ;
        RECT 6.575 1.915 6.745 4.535 ;
        RECT 28.035 1.915 28.205 4.535 ;
        RECT 49.495 1.915 49.665 4.535 ;
      LAYER mcon ;
        RECT 6.575 2.505 6.745 2.675 ;
        RECT 28.035 2.505 28.205 2.675 ;
        RECT 49.495 2.505 49.665 2.675 ;
      LAYER met1 ;
        RECT 6.545 2.675 6.775 2.705 ;
        RECT 28.005 2.675 28.235 2.705 ;
        RECT 49.465 2.675 49.695 2.705 ;
        RECT 6.515 2.505 49.725 2.675 ;
        RECT 6.545 2.475 6.775 2.505 ;
        RECT 28.005 2.475 28.235 2.505 ;
        RECT 49.465 2.475 49.695 2.505 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.126300 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 13.265 4.710 13.435 4.865 ;
        RECT 13.235 4.535 13.435 4.710 ;
        RECT 13.235 1.915 13.405 4.535 ;
        RECT 23.595 1.915 23.765 4.865 ;
        RECT 34.725 4.710 34.895 4.865 ;
        RECT 34.695 4.535 34.895 4.710 ;
        RECT 34.695 1.915 34.865 4.535 ;
        RECT 45.055 1.915 45.225 4.865 ;
        RECT 56.185 4.710 56.355 4.865 ;
        RECT 56.155 4.535 56.355 4.710 ;
        RECT 56.155 1.915 56.325 4.535 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 13.235 4.355 13.405 4.525 ;
        RECT 23.595 4.355 23.765 4.525 ;
        RECT 34.695 4.355 34.865 4.525 ;
        RECT 45.055 4.355 45.225 4.525 ;
        RECT 56.155 4.355 56.325 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 13.205 4.525 13.435 4.555 ;
        RECT 23.565 4.525 23.795 4.555 ;
        RECT 34.665 4.525 34.895 4.555 ;
        RECT 45.025 4.525 45.255 4.555 ;
        RECT 56.125 4.525 56.355 4.555 ;
        RECT 2.075 4.520 13.465 4.525 ;
        RECT 16.745 4.520 56.385 4.525 ;
        RECT 2.075 4.365 56.385 4.520 ;
        RECT 2.075 4.355 13.465 4.365 ;
        RECT 16.745 4.355 56.385 4.365 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 13.205 4.325 13.435 4.355 ;
        RECT 23.565 4.325 23.795 4.355 ;
        RECT 34.665 4.325 34.895 4.355 ;
        RECT 45.025 4.325 45.255 4.355 ;
        RECT 56.125 4.325 56.355 4.355 ;
    END
  END CLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 74.805 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 74.540 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.515 5.135 5.685 7.230 ;
        RECT 6.395 5.555 6.565 7.230 ;
        RECT 7.275 5.555 7.445 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 8.845 5.135 9.015 7.230 ;
        RECT 9.725 5.555 9.895 7.230 ;
        RECT 10.605 5.555 10.775 7.230 ;
        RECT 11.300 4.110 11.640 7.230 ;
        RECT 12.175 5.135 12.345 7.230 ;
        RECT 13.055 5.555 13.225 7.230 ;
        RECT 13.935 5.555 14.105 7.230 ;
        RECT 14.630 4.110 14.970 7.230 ;
        RECT 15.505 5.135 15.675 7.230 ;
        RECT 16.385 5.555 16.555 7.230 ;
        RECT 17.265 5.555 17.435 7.230 ;
        RECT 17.960 4.110 18.300 7.230 ;
        RECT 18.835 5.135 19.005 7.230 ;
        RECT 19.715 5.555 19.885 7.230 ;
        RECT 20.595 5.555 20.765 7.230 ;
        RECT 21.290 4.110 21.630 7.230 ;
        RECT 22.465 5.215 22.635 7.230 ;
        RECT 23.345 5.555 23.515 7.230 ;
        RECT 24.225 5.555 24.395 7.230 ;
        RECT 25.105 5.555 25.275 7.230 ;
        RECT 26.100 4.110 26.440 7.230 ;
        RECT 26.975 5.135 27.145 7.230 ;
        RECT 27.855 5.555 28.025 7.230 ;
        RECT 28.735 5.555 28.905 7.230 ;
        RECT 29.430 4.110 29.770 7.230 ;
        RECT 30.305 5.135 30.475 7.230 ;
        RECT 31.185 5.555 31.355 7.230 ;
        RECT 32.065 5.555 32.235 7.230 ;
        RECT 32.760 4.110 33.100 7.230 ;
        RECT 33.635 5.135 33.805 7.230 ;
        RECT 34.515 5.555 34.685 7.230 ;
        RECT 35.395 5.555 35.565 7.230 ;
        RECT 36.090 4.110 36.430 7.230 ;
        RECT 36.965 5.135 37.135 7.230 ;
        RECT 37.845 5.555 38.015 7.230 ;
        RECT 38.725 5.555 38.895 7.230 ;
        RECT 39.420 4.110 39.760 7.230 ;
        RECT 40.295 5.135 40.465 7.230 ;
        RECT 41.175 5.555 41.345 7.230 ;
        RECT 42.055 5.555 42.225 7.230 ;
        RECT 42.750 4.110 43.090 7.230 ;
        RECT 43.925 5.215 44.095 7.230 ;
        RECT 44.805 5.555 44.975 7.230 ;
        RECT 45.685 5.555 45.855 7.230 ;
        RECT 46.565 5.555 46.735 7.230 ;
        RECT 47.560 4.110 47.900 7.230 ;
        RECT 48.435 5.135 48.605 7.230 ;
        RECT 49.315 5.555 49.485 7.230 ;
        RECT 50.195 5.555 50.365 7.230 ;
        RECT 50.890 4.110 51.230 7.230 ;
        RECT 51.765 5.135 51.935 7.230 ;
        RECT 52.645 5.555 52.815 7.230 ;
        RECT 53.525 5.555 53.695 7.230 ;
        RECT 54.220 4.110 54.560 7.230 ;
        RECT 55.095 5.135 55.265 7.230 ;
        RECT 55.975 5.555 56.145 7.230 ;
        RECT 56.855 5.555 57.025 7.230 ;
        RECT 57.550 4.110 57.890 7.230 ;
        RECT 58.425 5.135 58.595 7.230 ;
        RECT 59.305 5.555 59.475 7.230 ;
        RECT 60.185 5.555 60.355 7.230 ;
        RECT 60.880 4.110 61.220 7.230 ;
        RECT 61.755 5.135 61.925 7.230 ;
        RECT 62.635 5.555 62.805 7.230 ;
        RECT 63.515 5.555 63.685 7.230 ;
        RECT 64.210 4.110 64.550 7.230 ;
        RECT 65.085 5.125 65.255 7.230 ;
        RECT 65.965 5.555 66.135 7.230 ;
        RECT 66.845 5.125 67.015 7.230 ;
        RECT 67.540 4.110 67.880 7.230 ;
        RECT 70.870 4.110 71.210 7.230 ;
        RECT 74.200 4.110 74.540 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.625 7.315 30.795 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.435 7.315 35.605 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
        RECT 38.765 7.315 38.935 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.615 7.315 40.785 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 43.205 7.315 43.375 7.485 ;
        RECT 43.575 7.315 43.745 7.485 ;
        RECT 43.945 7.315 44.115 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 48.015 7.315 48.185 7.485 ;
        RECT 48.385 7.315 48.555 7.485 ;
        RECT 48.755 7.315 48.925 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 51.715 7.315 51.885 7.485 ;
        RECT 52.085 7.315 52.255 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 52.825 7.315 52.995 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.525 7.315 56.695 7.485 ;
        RECT 56.895 7.315 57.065 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 61.335 7.315 61.505 7.485 ;
        RECT 61.705 7.315 61.875 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.445 7.315 62.615 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.665 7.315 64.835 7.485 ;
        RECT 65.035 7.315 65.205 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.255 7.315 67.425 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.365 7.315 68.535 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.475 7.315 69.645 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.065 7.315 72.235 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.175 7.315 73.345 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 74.540 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 74.540 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.905 0.170 6.075 1.120 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.235 0.170 9.405 1.120 ;
        RECT 11.300 0.170 11.640 2.720 ;
        RECT 12.565 0.170 12.735 1.120 ;
        RECT 14.630 0.170 14.970 2.720 ;
        RECT 15.895 0.170 16.065 1.120 ;
        RECT 17.960 0.170 18.300 2.720 ;
        RECT 19.225 0.170 19.395 1.120 ;
        RECT 21.290 0.170 21.630 2.720 ;
        RECT 22.450 0.170 22.620 1.130 ;
        RECT 26.100 0.170 26.440 2.720 ;
        RECT 27.365 0.170 27.535 1.120 ;
        RECT 29.430 0.170 29.770 2.720 ;
        RECT 30.695 0.170 30.865 1.120 ;
        RECT 32.760 0.170 33.100 2.720 ;
        RECT 34.025 0.170 34.195 1.120 ;
        RECT 36.090 0.170 36.430 2.720 ;
        RECT 37.355 0.170 37.525 1.120 ;
        RECT 39.420 0.170 39.760 2.720 ;
        RECT 40.685 0.170 40.855 1.120 ;
        RECT 42.750 0.170 43.090 2.720 ;
        RECT 43.910 0.170 44.080 1.130 ;
        RECT 47.560 0.170 47.900 2.720 ;
        RECT 48.825 0.170 48.995 1.120 ;
        RECT 50.890 0.170 51.230 2.720 ;
        RECT 52.155 0.170 52.325 1.120 ;
        RECT 54.220 0.170 54.560 2.720 ;
        RECT 55.485 0.170 55.655 1.120 ;
        RECT 57.550 0.170 57.890 2.720 ;
        RECT 58.815 0.170 58.985 1.120 ;
        RECT 60.880 0.170 61.220 2.720 ;
        RECT 62.145 0.170 62.315 1.120 ;
        RECT 64.210 0.170 64.550 2.720 ;
        RECT 65.475 0.170 65.645 1.120 ;
        RECT 67.540 0.170 67.880 2.720 ;
        RECT 68.805 0.170 68.975 1.120 ;
        RECT 70.870 0.170 71.210 2.720 ;
        RECT 72.135 0.170 72.305 1.120 ;
        RECT 74.200 0.170 74.540 2.720 ;
        RECT -0.170 -0.170 74.540 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.625 -0.085 30.795 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.435 -0.085 35.605 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
        RECT 38.765 -0.085 38.935 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.615 -0.085 40.785 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 43.205 -0.085 43.375 0.085 ;
        RECT 43.575 -0.085 43.745 0.085 ;
        RECT 43.945 -0.085 44.115 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 48.015 -0.085 48.185 0.085 ;
        RECT 48.385 -0.085 48.555 0.085 ;
        RECT 48.755 -0.085 48.925 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 51.715 -0.085 51.885 0.085 ;
        RECT 52.085 -0.085 52.255 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 52.825 -0.085 52.995 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.525 -0.085 56.695 0.085 ;
        RECT 56.895 -0.085 57.065 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 61.335 -0.085 61.505 0.085 ;
        RECT 61.705 -0.085 61.875 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.445 -0.085 62.615 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.665 -0.085 64.835 0.085 ;
        RECT 65.035 -0.085 65.205 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.255 -0.085 67.425 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.365 -0.085 68.535 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.475 -0.085 69.645 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.065 -0.085 72.235 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.175 -0.085 73.345 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 74.540 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 5.955 5.285 6.125 7.020 ;
        RECT 6.835 5.285 7.005 7.020 ;
        RECT 9.285 5.285 9.455 7.020 ;
        RECT 10.165 5.285 10.335 7.020 ;
        RECT 12.615 5.285 12.785 7.020 ;
        RECT 13.495 5.285 13.665 7.020 ;
        RECT 15.945 5.285 16.115 7.020 ;
        RECT 16.825 5.285 16.995 7.020 ;
        RECT 19.275 5.285 19.445 7.020 ;
        RECT 20.155 5.285 20.325 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 5.955 5.115 7.485 5.285 ;
        RECT 9.285 5.115 10.815 5.285 ;
        RECT 12.615 5.115 14.145 5.285 ;
        RECT 15.945 5.115 17.475 5.285 ;
        RECT 19.275 5.115 20.805 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.420 1.665 5.590 1.745 ;
        RECT 6.390 1.665 6.560 1.745 ;
        RECT 7.315 1.740 7.485 5.115 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 9.935 4.710 10.105 4.865 ;
        RECT 9.905 4.535 10.105 4.710 ;
        RECT 9.905 1.915 10.075 4.535 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.420 1.495 6.560 1.665 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.420 0.365 5.590 1.495 ;
        RECT 6.390 0.615 6.560 1.495 ;
        RECT 6.875 1.570 7.485 1.740 ;
        RECT 8.750 1.665 8.920 1.745 ;
        RECT 9.720 1.665 9.890 1.745 ;
        RECT 10.645 1.740 10.815 5.115 ;
        RECT 12.495 1.915 12.665 4.865 ;
        RECT 6.875 0.835 7.045 1.570 ;
        RECT 8.750 1.495 9.890 1.665 ;
        RECT 7.360 0.615 7.530 1.385 ;
        RECT 6.390 0.445 7.530 0.615 ;
        RECT 6.390 0.365 6.560 0.445 ;
        RECT 7.360 0.365 7.530 0.445 ;
        RECT 8.750 0.365 8.920 1.495 ;
        RECT 9.720 0.615 9.890 1.495 ;
        RECT 10.205 1.570 10.815 1.740 ;
        RECT 12.080 1.665 12.250 1.745 ;
        RECT 13.050 1.665 13.220 1.745 ;
        RECT 13.975 1.740 14.145 5.115 ;
        RECT 15.825 1.915 15.995 4.865 ;
        RECT 16.595 4.710 16.765 4.865 ;
        RECT 16.565 4.535 16.765 4.710 ;
        RECT 16.565 1.915 16.735 4.535 ;
        RECT 10.205 0.835 10.375 1.570 ;
        RECT 12.080 1.495 13.220 1.665 ;
        RECT 10.690 0.615 10.860 1.385 ;
        RECT 9.720 0.445 10.860 0.615 ;
        RECT 9.720 0.365 9.890 0.445 ;
        RECT 10.690 0.365 10.860 0.445 ;
        RECT 12.080 0.365 12.250 1.495 ;
        RECT 13.050 0.615 13.220 1.495 ;
        RECT 13.535 1.570 14.145 1.740 ;
        RECT 15.410 1.665 15.580 1.745 ;
        RECT 16.380 1.665 16.550 1.745 ;
        RECT 17.305 1.740 17.475 5.115 ;
        RECT 19.155 1.915 19.325 4.865 ;
        RECT 19.925 4.710 20.095 4.865 ;
        RECT 19.895 4.535 20.095 4.710 ;
        RECT 19.895 1.915 20.065 4.535 ;
        RECT 13.535 0.835 13.705 1.570 ;
        RECT 15.410 1.495 16.550 1.665 ;
        RECT 14.020 0.615 14.190 1.385 ;
        RECT 13.050 0.445 14.190 0.615 ;
        RECT 13.050 0.365 13.220 0.445 ;
        RECT 14.020 0.365 14.190 0.445 ;
        RECT 15.410 0.365 15.580 1.495 ;
        RECT 16.380 0.615 16.550 1.495 ;
        RECT 16.865 1.570 17.475 1.740 ;
        RECT 18.740 1.665 18.910 1.745 ;
        RECT 19.710 1.665 19.880 1.745 ;
        RECT 20.635 1.740 20.805 5.115 ;
        RECT 22.905 5.240 23.075 7.020 ;
        RECT 23.785 5.240 23.955 7.020 ;
        RECT 24.665 5.240 24.835 7.020 ;
        RECT 27.415 5.285 27.585 7.020 ;
        RECT 28.295 5.285 28.465 7.020 ;
        RECT 30.745 5.285 30.915 7.020 ;
        RECT 31.625 5.285 31.795 7.020 ;
        RECT 34.075 5.285 34.245 7.020 ;
        RECT 34.955 5.285 35.125 7.020 ;
        RECT 37.405 5.285 37.575 7.020 ;
        RECT 38.285 5.285 38.455 7.020 ;
        RECT 40.735 5.285 40.905 7.020 ;
        RECT 41.615 5.285 41.785 7.020 ;
        RECT 22.905 5.070 25.615 5.240 ;
        RECT 27.415 5.115 28.945 5.285 ;
        RECT 30.745 5.115 32.275 5.285 ;
        RECT 34.075 5.115 35.605 5.285 ;
        RECT 37.405 5.115 38.935 5.285 ;
        RECT 40.735 5.115 42.265 5.285 ;
        RECT 22.485 1.915 22.655 4.865 ;
        RECT 24.705 1.915 24.875 4.865 ;
        RECT 16.865 0.835 17.035 1.570 ;
        RECT 18.740 1.495 19.880 1.665 ;
        RECT 17.350 0.615 17.520 1.385 ;
        RECT 16.380 0.445 17.520 0.615 ;
        RECT 16.380 0.365 16.550 0.445 ;
        RECT 17.350 0.365 17.520 0.445 ;
        RECT 18.740 0.365 18.910 1.495 ;
        RECT 19.710 0.615 19.880 1.495 ;
        RECT 20.195 1.570 20.805 1.740 ;
        RECT 21.965 1.675 22.135 1.755 ;
        RECT 22.935 1.675 23.105 1.755 ;
        RECT 23.905 1.675 24.075 1.755 ;
        RECT 20.195 0.835 20.365 1.570 ;
        RECT 21.965 1.505 24.075 1.675 ;
        RECT 20.680 0.615 20.850 1.385 ;
        RECT 19.710 0.445 20.850 0.615 ;
        RECT 19.710 0.365 19.880 0.445 ;
        RECT 20.680 0.365 20.850 0.445 ;
        RECT 21.965 0.375 22.135 1.505 ;
        RECT 22.935 0.625 23.105 1.505 ;
        RECT 23.905 1.425 24.075 1.505 ;
        RECT 23.425 1.080 23.595 1.160 ;
        RECT 24.475 1.080 24.645 1.755 ;
        RECT 25.445 1.750 25.615 5.070 ;
        RECT 27.295 1.915 27.465 4.865 ;
        RECT 23.425 0.910 24.645 1.080 ;
        RECT 23.425 0.830 23.595 0.910 ;
        RECT 23.905 0.625 24.075 0.705 ;
        RECT 22.935 0.455 24.075 0.625 ;
        RECT 22.935 0.375 23.105 0.455 ;
        RECT 23.905 0.375 24.075 0.455 ;
        RECT 24.475 0.625 24.645 0.910 ;
        RECT 24.960 1.580 25.615 1.750 ;
        RECT 26.880 1.665 27.050 1.745 ;
        RECT 27.850 1.665 28.020 1.745 ;
        RECT 28.775 1.740 28.945 5.115 ;
        RECT 30.625 1.915 30.795 4.865 ;
        RECT 31.395 4.710 31.565 4.865 ;
        RECT 31.365 4.535 31.565 4.710 ;
        RECT 31.365 1.915 31.535 4.535 ;
        RECT 24.960 0.845 25.130 1.580 ;
        RECT 26.880 1.495 28.020 1.665 ;
        RECT 25.445 0.625 25.615 1.395 ;
        RECT 24.475 0.455 25.615 0.625 ;
        RECT 24.475 0.375 24.645 0.455 ;
        RECT 25.445 0.375 25.615 0.455 ;
        RECT 26.880 0.365 27.050 1.495 ;
        RECT 27.850 0.615 28.020 1.495 ;
        RECT 28.335 1.570 28.945 1.740 ;
        RECT 30.210 1.665 30.380 1.745 ;
        RECT 31.180 1.665 31.350 1.745 ;
        RECT 32.105 1.740 32.275 5.115 ;
        RECT 33.955 1.915 34.125 4.865 ;
        RECT 28.335 0.835 28.505 1.570 ;
        RECT 30.210 1.495 31.350 1.665 ;
        RECT 28.820 0.615 28.990 1.385 ;
        RECT 27.850 0.445 28.990 0.615 ;
        RECT 27.850 0.365 28.020 0.445 ;
        RECT 28.820 0.365 28.990 0.445 ;
        RECT 30.210 0.365 30.380 1.495 ;
        RECT 31.180 0.615 31.350 1.495 ;
        RECT 31.665 1.570 32.275 1.740 ;
        RECT 33.540 1.665 33.710 1.745 ;
        RECT 34.510 1.665 34.680 1.745 ;
        RECT 35.435 1.740 35.605 5.115 ;
        RECT 37.285 1.915 37.455 4.865 ;
        RECT 38.055 4.710 38.225 4.865 ;
        RECT 38.025 4.535 38.225 4.710 ;
        RECT 38.025 1.915 38.195 4.535 ;
        RECT 31.665 0.835 31.835 1.570 ;
        RECT 33.540 1.495 34.680 1.665 ;
        RECT 32.150 0.615 32.320 1.385 ;
        RECT 31.180 0.445 32.320 0.615 ;
        RECT 31.180 0.365 31.350 0.445 ;
        RECT 32.150 0.365 32.320 0.445 ;
        RECT 33.540 0.365 33.710 1.495 ;
        RECT 34.510 0.615 34.680 1.495 ;
        RECT 34.995 1.570 35.605 1.740 ;
        RECT 36.870 1.665 37.040 1.745 ;
        RECT 37.840 1.665 38.010 1.745 ;
        RECT 38.765 1.740 38.935 5.115 ;
        RECT 40.615 1.915 40.785 4.865 ;
        RECT 41.385 4.710 41.555 4.865 ;
        RECT 41.355 4.535 41.555 4.710 ;
        RECT 41.355 1.915 41.525 4.535 ;
        RECT 34.995 0.835 35.165 1.570 ;
        RECT 36.870 1.495 38.010 1.665 ;
        RECT 35.480 0.615 35.650 1.385 ;
        RECT 34.510 0.445 35.650 0.615 ;
        RECT 34.510 0.365 34.680 0.445 ;
        RECT 35.480 0.365 35.650 0.445 ;
        RECT 36.870 0.365 37.040 1.495 ;
        RECT 37.840 0.615 38.010 1.495 ;
        RECT 38.325 1.570 38.935 1.740 ;
        RECT 40.200 1.665 40.370 1.745 ;
        RECT 41.170 1.665 41.340 1.745 ;
        RECT 42.095 1.740 42.265 5.115 ;
        RECT 44.365 5.240 44.535 7.020 ;
        RECT 45.245 5.240 45.415 7.020 ;
        RECT 46.125 5.240 46.295 7.020 ;
        RECT 48.875 5.285 49.045 7.020 ;
        RECT 49.755 5.285 49.925 7.020 ;
        RECT 52.205 5.285 52.375 7.020 ;
        RECT 53.085 5.285 53.255 7.020 ;
        RECT 55.535 5.285 55.705 7.020 ;
        RECT 56.415 5.285 56.585 7.020 ;
        RECT 58.865 5.285 59.035 7.020 ;
        RECT 59.745 5.285 59.915 7.020 ;
        RECT 62.195 5.285 62.365 7.020 ;
        RECT 63.075 5.285 63.245 7.020 ;
        RECT 65.525 6.825 65.705 6.995 ;
        RECT 65.525 5.295 65.695 6.825 ;
        RECT 66.405 5.295 66.575 6.995 ;
        RECT 44.365 5.070 47.075 5.240 ;
        RECT 48.875 5.115 50.405 5.285 ;
        RECT 52.205 5.115 53.735 5.285 ;
        RECT 55.535 5.115 57.065 5.285 ;
        RECT 58.865 5.115 60.395 5.285 ;
        RECT 62.195 5.115 63.725 5.285 ;
        RECT 65.525 5.125 66.575 5.295 ;
        RECT 43.945 1.915 44.115 4.865 ;
        RECT 46.165 1.915 46.335 4.865 ;
        RECT 38.325 0.835 38.495 1.570 ;
        RECT 40.200 1.495 41.340 1.665 ;
        RECT 38.810 0.615 38.980 1.385 ;
        RECT 37.840 0.445 38.980 0.615 ;
        RECT 37.840 0.365 38.010 0.445 ;
        RECT 38.810 0.365 38.980 0.445 ;
        RECT 40.200 0.365 40.370 1.495 ;
        RECT 41.170 0.615 41.340 1.495 ;
        RECT 41.655 1.570 42.265 1.740 ;
        RECT 43.425 1.675 43.595 1.755 ;
        RECT 44.395 1.675 44.565 1.755 ;
        RECT 45.365 1.675 45.535 1.755 ;
        RECT 41.655 0.835 41.825 1.570 ;
        RECT 43.425 1.505 45.535 1.675 ;
        RECT 42.140 0.615 42.310 1.385 ;
        RECT 41.170 0.445 42.310 0.615 ;
        RECT 41.170 0.365 41.340 0.445 ;
        RECT 42.140 0.365 42.310 0.445 ;
        RECT 43.425 0.375 43.595 1.505 ;
        RECT 44.395 0.625 44.565 1.505 ;
        RECT 45.365 1.425 45.535 1.505 ;
        RECT 44.885 1.080 45.055 1.160 ;
        RECT 45.935 1.080 46.105 1.755 ;
        RECT 46.905 1.750 47.075 5.070 ;
        RECT 48.755 1.915 48.925 4.865 ;
        RECT 44.885 0.910 46.105 1.080 ;
        RECT 44.885 0.830 45.055 0.910 ;
        RECT 45.365 0.625 45.535 0.705 ;
        RECT 44.395 0.455 45.535 0.625 ;
        RECT 44.395 0.375 44.565 0.455 ;
        RECT 45.365 0.375 45.535 0.455 ;
        RECT 45.935 0.625 46.105 0.910 ;
        RECT 46.420 1.580 47.075 1.750 ;
        RECT 48.340 1.665 48.510 1.745 ;
        RECT 49.310 1.665 49.480 1.745 ;
        RECT 50.235 1.740 50.405 5.115 ;
        RECT 52.085 1.915 52.255 4.865 ;
        RECT 52.855 4.710 53.025 4.865 ;
        RECT 52.825 4.535 53.025 4.710 ;
        RECT 52.825 1.915 52.995 4.535 ;
        RECT 46.420 0.845 46.590 1.580 ;
        RECT 48.340 1.495 49.480 1.665 ;
        RECT 46.905 0.625 47.075 1.395 ;
        RECT 45.935 0.455 47.075 0.625 ;
        RECT 45.935 0.375 46.105 0.455 ;
        RECT 46.905 0.375 47.075 0.455 ;
        RECT 48.340 0.365 48.510 1.495 ;
        RECT 49.310 0.615 49.480 1.495 ;
        RECT 49.795 1.570 50.405 1.740 ;
        RECT 51.670 1.665 51.840 1.745 ;
        RECT 52.640 1.665 52.810 1.745 ;
        RECT 53.565 1.740 53.735 5.115 ;
        RECT 55.415 1.915 55.585 4.865 ;
        RECT 49.795 0.835 49.965 1.570 ;
        RECT 51.670 1.495 52.810 1.665 ;
        RECT 50.280 0.615 50.450 1.385 ;
        RECT 49.310 0.445 50.450 0.615 ;
        RECT 49.310 0.365 49.480 0.445 ;
        RECT 50.280 0.365 50.450 0.445 ;
        RECT 51.670 0.365 51.840 1.495 ;
        RECT 52.640 0.615 52.810 1.495 ;
        RECT 53.125 1.570 53.735 1.740 ;
        RECT 55.000 1.665 55.170 1.745 ;
        RECT 55.970 1.665 56.140 1.745 ;
        RECT 56.895 1.740 57.065 5.115 ;
        RECT 58.745 1.915 58.915 4.865 ;
        RECT 59.515 4.710 59.685 4.865 ;
        RECT 59.485 4.535 59.685 4.710 ;
        RECT 59.485 1.915 59.655 4.535 ;
        RECT 53.125 0.835 53.295 1.570 ;
        RECT 55.000 1.495 56.140 1.665 ;
        RECT 53.610 0.615 53.780 1.385 ;
        RECT 52.640 0.445 53.780 0.615 ;
        RECT 52.640 0.365 52.810 0.445 ;
        RECT 53.610 0.365 53.780 0.445 ;
        RECT 55.000 0.365 55.170 1.495 ;
        RECT 55.970 0.615 56.140 1.495 ;
        RECT 56.455 1.570 57.065 1.740 ;
        RECT 58.330 1.665 58.500 1.745 ;
        RECT 59.300 1.665 59.470 1.745 ;
        RECT 60.225 1.740 60.395 5.115 ;
        RECT 62.075 1.915 62.245 4.865 ;
        RECT 62.845 4.710 63.015 4.865 ;
        RECT 62.815 4.535 63.015 4.710 ;
        RECT 62.815 1.915 62.985 4.535 ;
        RECT 56.455 0.835 56.625 1.570 ;
        RECT 58.330 1.495 59.470 1.665 ;
        RECT 56.940 0.615 57.110 1.385 ;
        RECT 55.970 0.445 57.110 0.615 ;
        RECT 55.970 0.365 56.140 0.445 ;
        RECT 56.940 0.365 57.110 0.445 ;
        RECT 58.330 0.365 58.500 1.495 ;
        RECT 59.300 0.615 59.470 1.495 ;
        RECT 59.785 1.570 60.395 1.740 ;
        RECT 61.660 1.665 61.830 1.745 ;
        RECT 62.630 1.665 62.800 1.745 ;
        RECT 63.555 1.740 63.725 5.115 ;
        RECT 66.405 5.045 66.575 5.125 ;
        RECT 68.405 6.825 70.335 6.995 ;
        RECT 68.405 5.045 68.575 6.825 ;
        RECT 68.845 5.295 69.015 6.565 ;
        RECT 69.285 5.555 69.455 6.825 ;
        RECT 69.725 5.295 69.895 6.565 ;
        RECT 70.165 5.375 70.335 6.825 ;
        RECT 71.745 6.825 73.675 6.995 ;
        RECT 68.845 5.125 69.895 5.295 ;
        RECT 69.725 5.045 69.895 5.125 ;
        RECT 71.745 5.045 71.915 6.825 ;
        RECT 72.625 5.555 72.795 6.825 ;
        RECT 73.505 5.555 73.675 6.825 ;
        RECT 65.035 1.915 65.205 4.870 ;
        RECT 66.185 4.710 66.355 4.870 ;
        RECT 66.145 4.540 66.355 4.710 ;
        RECT 66.145 1.915 66.315 4.540 ;
        RECT 68.735 1.915 68.905 4.870 ;
        RECT 70.215 1.915 70.385 4.870 ;
        RECT 71.695 1.915 71.865 4.870 ;
        RECT 72.805 4.540 72.995 4.870 ;
        RECT 72.805 1.915 72.975 4.540 ;
        RECT 59.785 0.835 59.955 1.570 ;
        RECT 61.660 1.495 62.800 1.665 ;
        RECT 60.270 0.615 60.440 1.385 ;
        RECT 59.300 0.445 60.440 0.615 ;
        RECT 59.300 0.365 59.470 0.445 ;
        RECT 60.270 0.365 60.440 0.445 ;
        RECT 61.660 0.365 61.830 1.495 ;
        RECT 62.630 0.615 62.800 1.495 ;
        RECT 63.115 1.570 63.725 1.740 ;
        RECT 64.990 1.665 65.160 1.745 ;
        RECT 65.960 1.665 66.130 1.745 ;
        RECT 63.115 0.835 63.285 1.570 ;
        RECT 64.990 1.495 66.130 1.665 ;
        RECT 63.600 0.615 63.770 1.385 ;
        RECT 62.630 0.445 63.770 0.615 ;
        RECT 62.630 0.365 62.800 0.445 ;
        RECT 63.600 0.365 63.770 0.445 ;
        RECT 64.990 0.365 65.160 1.495 ;
        RECT 65.960 0.615 66.130 1.495 ;
        RECT 66.930 0.615 67.100 1.745 ;
        RECT 65.960 0.445 67.100 0.615 ;
        RECT 65.960 0.365 66.130 0.445 ;
        RECT 66.930 0.365 67.100 0.445 ;
        RECT 68.320 1.665 68.490 1.745 ;
        RECT 69.290 1.665 69.460 1.745 ;
        RECT 68.320 1.495 69.460 1.665 ;
        RECT 68.320 0.365 68.490 1.495 ;
        RECT 69.290 0.615 69.460 1.495 ;
        RECT 70.260 0.615 70.430 1.745 ;
        RECT 69.290 0.445 70.430 0.615 ;
        RECT 69.290 0.365 69.460 0.445 ;
        RECT 70.260 0.365 70.430 0.445 ;
        RECT 71.650 1.665 71.820 1.745 ;
        RECT 72.620 1.665 72.790 1.745 ;
        RECT 71.650 1.495 72.790 1.665 ;
        RECT 71.650 0.365 71.820 1.495 ;
        RECT 72.620 0.615 72.790 1.495 ;
        RECT 73.590 0.615 73.760 1.390 ;
        RECT 72.620 0.445 73.760 0.615 ;
        RECT 72.620 0.365 72.790 0.445 ;
        RECT 73.590 0.365 73.760 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 7.315 3.245 7.485 3.415 ;
        RECT 9.165 3.245 9.335 3.415 ;
        RECT 9.905 3.985 10.075 4.155 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 12.495 3.245 12.665 3.415 ;
        RECT 13.975 3.985 14.145 4.155 ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 16.565 2.875 16.735 3.045 ;
        RECT 17.305 3.615 17.475 3.785 ;
        RECT 19.155 3.615 19.325 3.785 ;
        RECT 19.895 3.985 20.065 4.155 ;
        RECT 20.635 2.875 20.805 3.045 ;
        RECT 22.485 3.985 22.655 4.155 ;
        RECT 24.705 3.245 24.875 3.415 ;
        RECT 25.445 3.615 25.615 3.785 ;
        RECT 27.295 3.615 27.465 3.785 ;
        RECT 28.775 3.245 28.945 3.415 ;
        RECT 30.625 3.245 30.795 3.415 ;
        RECT 31.365 3.985 31.535 4.155 ;
        RECT 32.105 3.245 32.275 3.415 ;
        RECT 33.955 3.245 34.125 3.415 ;
        RECT 35.435 3.985 35.605 4.155 ;
        RECT 37.285 3.615 37.455 3.785 ;
        RECT 38.025 2.135 38.195 2.305 ;
        RECT 38.765 3.615 38.935 3.785 ;
        RECT 40.615 3.615 40.785 3.785 ;
        RECT 41.355 3.985 41.525 4.155 ;
        RECT 66.405 5.125 66.575 5.295 ;
        RECT 42.095 2.135 42.265 2.305 ;
        RECT 43.945 3.985 44.115 4.155 ;
        RECT 46.165 3.245 46.335 3.415 ;
        RECT 46.905 3.615 47.075 3.785 ;
        RECT 48.755 3.615 48.925 3.785 ;
        RECT 50.235 3.245 50.405 3.415 ;
        RECT 52.085 3.245 52.255 3.415 ;
        RECT 52.825 3.985 52.995 4.155 ;
        RECT 53.565 3.245 53.735 3.415 ;
        RECT 55.415 3.245 55.585 3.415 ;
        RECT 56.895 3.985 57.065 4.155 ;
        RECT 58.745 3.615 58.915 3.785 ;
        RECT 59.485 3.615 59.655 3.785 ;
        RECT 60.225 4.355 60.395 4.525 ;
        RECT 62.075 4.355 62.245 4.525 ;
        RECT 62.815 3.985 62.985 4.155 ;
        RECT 68.405 5.125 68.575 5.295 ;
        RECT 69.725 5.125 69.895 5.295 ;
        RECT 71.745 5.125 71.915 5.295 ;
        RECT 63.555 3.615 63.725 3.785 ;
        RECT 65.035 4.355 65.205 4.525 ;
        RECT 65.035 3.615 65.205 3.785 ;
        RECT 66.145 3.985 66.315 4.155 ;
        RECT 66.145 2.135 66.315 2.305 ;
        RECT 68.735 4.355 68.905 4.525 ;
        RECT 70.215 2.875 70.385 3.045 ;
        RECT 70.215 1.995 70.385 2.165 ;
        RECT 71.695 1.995 71.865 2.165 ;
        RECT 72.805 3.985 72.975 4.155 ;
      LAYER met1 ;
        RECT 66.375 5.295 66.605 5.325 ;
        RECT 68.375 5.295 68.605 5.325 ;
        RECT 69.695 5.295 69.925 5.325 ;
        RECT 71.715 5.295 71.945 5.325 ;
        RECT 66.345 5.125 68.635 5.295 ;
        RECT 69.665 5.125 71.975 5.295 ;
        RECT 66.375 5.095 66.605 5.125 ;
        RECT 68.375 5.095 68.605 5.125 ;
        RECT 69.695 5.095 69.925 5.125 ;
        RECT 71.715 5.095 71.945 5.125 ;
        RECT 60.195 4.525 60.425 4.555 ;
        RECT 62.045 4.525 62.275 4.555 ;
        RECT 65.005 4.525 65.235 4.555 ;
        RECT 68.705 4.525 68.935 4.555 ;
        RECT 60.165 4.355 62.305 4.525 ;
        RECT 64.975 4.355 68.965 4.525 ;
        RECT 60.195 4.325 60.425 4.355 ;
        RECT 62.045 4.325 62.275 4.355 ;
        RECT 65.005 4.325 65.235 4.355 ;
        RECT 68.705 4.325 68.935 4.355 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 9.875 4.155 10.105 4.185 ;
        RECT 13.945 4.155 14.175 4.185 ;
        RECT 19.865 4.155 20.095 4.185 ;
        RECT 22.455 4.155 22.685 4.185 ;
        RECT 31.335 4.155 31.565 4.185 ;
        RECT 35.405 4.155 35.635 4.185 ;
        RECT 41.325 4.155 41.555 4.185 ;
        RECT 43.915 4.155 44.145 4.185 ;
        RECT 52.795 4.155 53.025 4.185 ;
        RECT 56.865 4.155 57.095 4.185 ;
        RECT 62.785 4.155 63.015 4.185 ;
        RECT 66.115 4.155 66.345 4.185 ;
        RECT 72.775 4.155 73.005 4.185 ;
        RECT 0.965 3.985 20.125 4.155 ;
        RECT 22.425 3.985 41.585 4.155 ;
        RECT 43.885 3.985 63.045 4.155 ;
        RECT 66.085 3.985 73.035 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 9.875 3.955 10.105 3.985 ;
        RECT 13.945 3.955 14.175 3.985 ;
        RECT 19.865 3.955 20.095 3.985 ;
        RECT 22.455 3.955 22.685 3.985 ;
        RECT 31.335 3.955 31.565 3.985 ;
        RECT 35.405 3.955 35.635 3.985 ;
        RECT 41.325 3.955 41.555 3.985 ;
        RECT 43.915 3.955 44.145 3.985 ;
        RECT 52.795 3.955 53.025 3.985 ;
        RECT 56.865 3.955 57.095 3.985 ;
        RECT 62.785 3.955 63.015 3.985 ;
        RECT 66.115 3.955 66.345 3.985 ;
        RECT 72.775 3.955 73.005 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 17.275 3.785 17.505 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 25.415 3.785 25.645 3.815 ;
        RECT 27.265 3.785 27.495 3.815 ;
        RECT 37.255 3.785 37.485 3.815 ;
        RECT 38.735 3.785 38.965 3.815 ;
        RECT 40.585 3.785 40.815 3.815 ;
        RECT 46.875 3.785 47.105 3.815 ;
        RECT 48.725 3.785 48.955 3.815 ;
        RECT 58.715 3.785 58.945 3.815 ;
        RECT 59.455 3.785 59.685 3.815 ;
        RECT 63.525 3.785 63.755 3.815 ;
        RECT 65.005 3.785 65.235 3.815 ;
        RECT 3.925 3.615 16.055 3.785 ;
        RECT 17.245 3.615 19.385 3.785 ;
        RECT 25.385 3.615 37.515 3.785 ;
        RECT 38.705 3.615 40.845 3.785 ;
        RECT 46.845 3.615 58.975 3.785 ;
        RECT 59.425 3.615 65.265 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 17.275 3.585 17.505 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
        RECT 25.415 3.585 25.645 3.615 ;
        RECT 27.265 3.585 27.495 3.615 ;
        RECT 37.255 3.585 37.485 3.615 ;
        RECT 38.735 3.585 38.965 3.615 ;
        RECT 40.585 3.585 40.815 3.615 ;
        RECT 46.875 3.585 47.105 3.615 ;
        RECT 48.725 3.585 48.955 3.615 ;
        RECT 58.715 3.585 58.945 3.615 ;
        RECT 59.455 3.585 59.685 3.615 ;
        RECT 63.525 3.585 63.755 3.615 ;
        RECT 65.005 3.585 65.235 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 7.285 3.415 7.515 3.445 ;
        RECT 9.135 3.415 9.365 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.465 3.415 12.695 3.445 ;
        RECT 24.675 3.415 24.905 3.445 ;
        RECT 28.745 3.415 28.975 3.445 ;
        RECT 30.595 3.415 30.825 3.445 ;
        RECT 32.075 3.415 32.305 3.445 ;
        RECT 33.925 3.415 34.155 3.445 ;
        RECT 46.135 3.415 46.365 3.445 ;
        RECT 50.205 3.415 50.435 3.445 ;
        RECT 52.055 3.415 52.285 3.445 ;
        RECT 53.535 3.415 53.765 3.445 ;
        RECT 55.385 3.415 55.615 3.445 ;
        RECT 3.185 3.245 9.395 3.415 ;
        RECT 10.585 3.245 12.725 3.415 ;
        RECT 24.645 3.245 30.855 3.415 ;
        RECT 32.045 3.245 34.185 3.415 ;
        RECT 46.105 3.245 52.315 3.415 ;
        RECT 53.505 3.245 55.645 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 7.285 3.215 7.515 3.245 ;
        RECT 9.135 3.215 9.365 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.465 3.215 12.695 3.245 ;
        RECT 24.675 3.215 24.905 3.245 ;
        RECT 28.745 3.215 28.975 3.245 ;
        RECT 30.595 3.215 30.825 3.245 ;
        RECT 32.075 3.215 32.305 3.245 ;
        RECT 33.925 3.215 34.155 3.245 ;
        RECT 46.135 3.215 46.365 3.245 ;
        RECT 50.205 3.215 50.435 3.245 ;
        RECT 52.055 3.215 52.285 3.245 ;
        RECT 53.535 3.215 53.765 3.245 ;
        RECT 55.385 3.215 55.615 3.245 ;
        RECT 16.535 3.045 16.765 3.075 ;
        RECT 20.605 3.045 20.835 3.075 ;
        RECT 70.185 3.045 70.415 3.075 ;
        RECT 16.505 2.875 70.445 3.045 ;
        RECT 16.535 2.845 16.765 2.875 ;
        RECT 20.605 2.845 20.835 2.875 ;
        RECT 70.185 2.845 70.415 2.875 ;
        RECT 37.995 2.305 38.225 2.335 ;
        RECT 42.065 2.305 42.295 2.335 ;
        RECT 66.115 2.305 66.345 2.335 ;
        RECT 37.965 2.135 66.375 2.305 ;
        RECT 70.185 2.165 70.415 2.195 ;
        RECT 71.665 2.165 71.895 2.195 ;
        RECT 37.995 2.105 38.225 2.135 ;
        RECT 42.065 2.105 42.295 2.135 ;
        RECT 66.115 2.105 66.345 2.135 ;
        RECT 70.155 1.995 71.925 2.165 ;
        RECT 70.185 1.965 70.415 1.995 ;
        RECT 71.665 1.965 71.895 1.995 ;
  END
END TMRDFFQNX1
END LIBRARY

