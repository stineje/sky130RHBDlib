* SPICE3 file created from HA.ext - technology: sky130A

.subckt HA SUM COUT A B VDD GND
M1000 a_2351_1051.t1 a_1295_209.t3 SUM.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_1685_1051.t3 A.t0 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t7 B.t0 a_2351_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 GND A.t3 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=3.9597p pd=29.01u as=0p ps=0u
M1004 VDD.t13 A.t1 a_217_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 COUT.t2 a_217_1050.t6 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 SUM a_1295_209.t4 a_2332_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.14u as=0p ps=0u
M1007 a_1295_209.t1 A.t2 VDD.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t6 B.t2 a_217_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 GND A.t4 a_1666_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1010 SUM.t1 a_1295_209.t5 a_2351_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VDD.t5 B.t3 a_1917_990.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1685_1051.t1 a_1917_990.t4 SUM.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_217_1050.t1 A.t6 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 SUM.t4 a_1917_990.t5 a_1685_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_217_1050.t0 B.t5 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VDD.t2 a_217_1050.t7 COUT.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VDD.t11 A.t7 a_1685_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 SUM B.t8 a_1666_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 VDD.t9 A.t8 a_1295_209.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 COUT a_217_1050.t5 GND.t3 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1021 GND a_1917_990.t3 a_2332_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_2351_1051.t2 B.t6 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1917_990.t0 B.t7 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 SUM B 0.89fF
C1 SUM A 0.08fF
C2 B COUT 0.07fF
C3 A COUT 0.12fF
C4 B A 1.08fF
C5 SUM VDD 0.53fF
C6 COUT VDD 0.82fF
C7 B VDD 0.99fF
C8 A VDD 1.13fF
R0 a_217_1050.n3 a_217_1050.t7 512.525
R1 a_217_1050.n3 a_217_1050.t6 371.139
R2 a_217_1050.n4 a_217_1050.t5 210.434
R3 a_217_1050.n7 a_217_1050.n5 190.561
R4 a_217_1050.n5 a_217_1050.n2 179.052
R5 a_217_1050.n4 a_217_1050.n3 173.2
R6 a_217_1050.n5 a_217_1050.n4 153.043
R7 a_217_1050.n2 a_217_1050.n1 76.002
R8 a_217_1050.n7 a_217_1050.n6 15.218
R9 a_217_1050.n0 a_217_1050.t2 14.282
R10 a_217_1050.n0 a_217_1050.t0 14.282
R11 a_217_1050.n1 a_217_1050.t4 14.282
R12 a_217_1050.n1 a_217_1050.t1 14.282
R13 a_217_1050.n2 a_217_1050.n0 12.85
R14 a_217_1050.n8 a_217_1050.n7 12.014
R15 GND.n29 GND.n27 219.745
R16 GND.n113 GND.n112 219.745
R17 GND.n148 GND.n146 219.745
R18 GND.n183 GND.n181 219.745
R19 GND.n59 GND.n58 219.745
R20 GND.n29 GND.n28 85.529
R21 GND.n113 GND.n111 85.529
R22 GND.n148 GND.n147 85.529
R23 GND.n183 GND.n182 85.529
R24 GND.n59 GND.n57 85.529
R25 GND.n47 GND.n46 84.842
R26 GND.n77 GND.n76 84.842
R27 GND.n91 GND.n90 84.842
R28 GND.n8 GND.n1 76.145
R29 GND.n86 GND.n85 76
R30 GND.n8 GND.n7 76
R31 GND.n16 GND.n15 76
R32 GND.n23 GND.n22 76
R33 GND.n26 GND.n25 76
R34 GND.n33 GND.n32 76
R35 GND.n36 GND.n35 76
R36 GND.n39 GND.n38 76
R37 GND.n42 GND.n41 76
R38 GND.n45 GND.n44 76
R39 GND.n50 GND.n49 76
R40 GND.n53 GND.n52 76
R41 GND.n56 GND.n55 76
R42 GND.n63 GND.n62 76
R43 GND.n66 GND.n65 76
R44 GND.n69 GND.n68 76
R45 GND.n72 GND.n71 76
R46 GND.n75 GND.n74 76
R47 GND.n80 GND.n79 76
R48 GND.n83 GND.n82 76
R49 GND.n186 GND.n185 76
R50 GND.n179 GND.n178 76
R51 GND.n176 GND.n175 76
R52 GND.n168 GND.n167 76
R53 GND.n160 GND.n159 76
R54 GND.n151 GND.n150 76
R55 GND.n144 GND.n143 76
R56 GND.n141 GND.n140 76
R57 GND.n133 GND.n132 76
R58 GND.n125 GND.n124 76
R59 GND.n116 GND.n115 76
R60 GND.n109 GND.n108 76
R61 GND.n106 GND.n105 76
R62 GND.n103 GND.n102 76
R63 GND.n100 GND.n99 76
R64 GND.n97 GND.n96 76
R65 GND.n94 GND.n93 76
R66 GND.n89 GND.n88 76
R67 GND.n3 GND.t5 39.413
R68 GND.n156 GND.t1 39.412
R69 GND.n121 GND.t3 39.412
R70 GND.n172 GND.n171 35.01
R71 GND.n137 GND.n136 35.01
R72 GND.n5 GND.n4 19.735
R73 GND.n14 GND.n13 19.735
R74 GND.n21 GND.n20 19.735
R75 GND.n173 GND.n172 19.735
R76 GND.n165 GND.n164 19.735
R77 GND.n158 GND.n157 19.735
R78 GND.n138 GND.n137 19.735
R79 GND.n130 GND.n129 19.735
R80 GND.n123 GND.n122 19.735
R81 GND.n172 GND.n170 19.017
R82 GND.n137 GND.n135 19.017
R83 GND.n19 GND.n18 18.345
R84 GND.n156 GND.n155 17.185
R85 GND.n121 GND.n120 17.185
R86 GND.n3 GND.n2 17.185
R87 GND.n32 GND.n30 14.167
R88 GND.n62 GND.n60 14.167
R89 GND.n185 GND.n184 14.167
R90 GND.n150 GND.n149 14.167
R91 GND.n115 GND.n114 14.167
R92 GND.n88 GND.n87 13.653
R93 GND.n93 GND.n92 13.653
R94 GND.n96 GND.n95 13.653
R95 GND.n99 GND.n98 13.653
R96 GND.n102 GND.n101 13.653
R97 GND.n105 GND.n104 13.653
R98 GND.n108 GND.n107 13.653
R99 GND.n115 GND.n110 13.653
R100 GND.n124 GND.n117 13.653
R101 GND.n132 GND.n131 13.653
R102 GND.n140 GND.n139 13.653
R103 GND.n143 GND.n142 13.653
R104 GND.n150 GND.n145 13.653
R105 GND.n159 GND.n152 13.653
R106 GND.n167 GND.n166 13.653
R107 GND.n175 GND.n174 13.653
R108 GND.n178 GND.n177 13.653
R109 GND.n185 GND.n180 13.653
R110 GND.n82 GND.n81 13.653
R111 GND.n79 GND.n78 13.653
R112 GND.n74 GND.n73 13.653
R113 GND.n71 GND.n70 13.653
R114 GND.n68 GND.n67 13.653
R115 GND.n65 GND.n64 13.653
R116 GND.n62 GND.n61 13.653
R117 GND.n55 GND.n54 13.653
R118 GND.n52 GND.n51 13.653
R119 GND.n49 GND.n48 13.653
R120 GND.n44 GND.n43 13.653
R121 GND.n41 GND.n40 13.653
R122 GND.n38 GND.n37 13.653
R123 GND.n35 GND.n34 13.653
R124 GND.n32 GND.n31 13.653
R125 GND.n25 GND.n24 13.653
R126 GND.n22 GND.n17 13.653
R127 GND.n15 GND.n9 13.653
R128 GND.n7 GND.n6 13.653
R129 GND.n12 GND.n11 7.5
R130 GND.n170 GND.n169 7.5
R131 GND.n163 GND.n162 7.5
R132 GND.n135 GND.n134 7.5
R133 GND.n128 GND.n127 7.5
R134 GND.n30 GND.n29 7.312
R135 GND.n114 GND.n113 7.312
R136 GND.n149 GND.n148 7.312
R137 GND.n184 GND.n183 7.312
R138 GND.n60 GND.n59 7.312
R139 GND.n20 GND.n19 6.358
R140 GND.n4 GND.n3 6.139
R141 GND.n157 GND.n156 6.139
R142 GND.n122 GND.n121 6.139
R143 GND.n154 GND.n153 4.551
R144 GND.n119 GND.n118 4.551
R145 GND.n22 GND.n21 3.935
R146 GND.n49 GND.n47 3.935
R147 GND.n79 GND.n77 3.935
R148 GND.n175 GND.n173 3.935
R149 GND.n140 GND.n138 3.935
R150 GND.n93 GND.n91 3.935
R151 GND.n7 GND.n5 3.541
R152 GND.n159 GND.n158 3.541
R153 GND.n124 GND.n123 3.541
R154 GND.t1 GND.n154 2.238
R155 GND.t3 GND.n119 2.238
R156 GND.n11 GND.n10 1.935
R157 GND.n162 GND.n161 1.935
R158 GND.n127 GND.n126 1.935
R159 GND.n1 GND.n0 0.596
R160 GND.n85 GND.n84 0.596
R161 GND.n13 GND.n12 0.358
R162 GND.n164 GND.n163 0.358
R163 GND.n129 GND.n128 0.358
R164 GND.n33 GND.n26 0.29
R165 GND.n63 GND.n56 0.29
R166 GND.n186 GND.n179 0.29
R167 GND.n151 GND.n144 0.29
R168 GND.n116 GND.n109 0.29
R169 GND.n86 GND 0.207
R170 GND.n15 GND.n14 0.196
R171 GND.n167 GND.n165 0.196
R172 GND.n132 GND.n130 0.196
R173 GND.n45 GND.n42 0.181
R174 GND.n75 GND.n72 0.181
R175 GND.n100 GND.n97 0.181
R176 GND.n16 GND.n8 0.157
R177 GND.n23 GND.n16 0.157
R178 GND.n176 GND.n168 0.157
R179 GND.n168 GND.n160 0.157
R180 GND.n141 GND.n133 0.157
R181 GND.n133 GND.n125 0.157
R182 GND.n26 GND.n23 0.145
R183 GND.n36 GND.n33 0.145
R184 GND.n39 GND.n36 0.145
R185 GND.n42 GND.n39 0.145
R186 GND.n50 GND.n45 0.145
R187 GND.n53 GND.n50 0.145
R188 GND.n56 GND.n53 0.145
R189 GND.n66 GND.n63 0.145
R190 GND.n69 GND.n66 0.145
R191 GND.n72 GND.n69 0.145
R192 GND.n80 GND.n75 0.145
R193 GND.n83 GND.n80 0.145
R194 GND.n179 GND.n176 0.145
R195 GND.n160 GND.n151 0.145
R196 GND.n144 GND.n141 0.145
R197 GND.n125 GND.n116 0.145
R198 GND.n109 GND.n106 0.145
R199 GND.n106 GND.n103 0.145
R200 GND.n103 GND.n100 0.145
R201 GND.n97 GND.n94 0.145
R202 GND.n94 GND.n89 0.145
R203 GND.n89 GND.n86 0.145
R204 GND GND.n186 0.078
R205 GND GND.n83 0.066
R206 COUT.n2 COUT.n0 210.56
R207 COUT.n2 COUT.n1 174.201
R208 COUT.n3 COUT.n2 76
R209 COUT.n0 COUT.t0 14.282
R210 COUT.n0 COUT.t2 14.282
R211 COUT.n3 COUT 0.046
R212 a_1295_209.n1 a_1295_209.t5 477.179
R213 a_1295_209.n1 a_1295_209.t3 406.485
R214 a_1295_209.n2 a_1295_209.t4 269.148
R215 a_1295_209.n5 a_1295_209.n3 185.537
R216 a_1295_209.n3 a_1295_209.n0 184.007
R217 a_1295_209.n3 a_1295_209.n2 156.579
R218 a_1295_209.n2 a_1295_209.n1 125.359
R219 a_1295_209.n5 a_1295_209.n4 15.218
R220 a_1295_209.n0 a_1295_209.t2 14.282
R221 a_1295_209.n0 a_1295_209.t1 14.282
R222 a_1295_209.n6 a_1295_209.n5 12.014
R223 SUM.n8 SUM.n7 232.332
R224 SUM.n5 SUM.n4 210.593
R225 SUM.n5 SUM.n0 165.336
R226 SUM.n8 SUM.n6 165.336
R227 SUM SUM.n8 78.357
R228 SUM.n9 SUM.n5 76
R229 SUM.n4 SUM.n3 30
R230 SUM.n2 SUM.n1 24.383
R231 SUM.n4 SUM.n2 23.684
R232 SUM.n0 SUM.t2 14.282
R233 SUM.n0 SUM.t1 14.282
R234 SUM.n6 SUM.t0 14.282
R235 SUM.n6 SUM.t4 14.282
R236 SUM.n9 SUM 0.046
R237 a_2351_1051.t1 a_2351_1051.n0 101.663
R238 a_2351_1051.n0 a_2351_1051.t3 101.661
R239 a_2351_1051.n0 a_2351_1051.t0 14.294
R240 a_2351_1051.n0 a_2351_1051.t2 14.282
R241 a_1917_990.n2 a_1917_990.t5 477.179
R242 a_1917_990.n2 a_1917_990.t4 406.485
R243 a_1917_990.n4 a_1917_990.t3 384.505
R244 a_1917_990.n3 a_1917_990.n2 228.016
R245 a_1917_990.n6 a_1917_990.n4 152.462
R246 a_1917_990.n3 a_1917_990.n1 130.901
R247 a_1917_990.n4 a_1917_990.n3 79.658
R248 a_1917_990.n7 a_1917_990.n0 55.263
R249 a_1917_990.n6 a_1917_990.n5 30
R250 a_1917_990.n7 a_1917_990.n6 23.684
R251 a_1917_990.n1 a_1917_990.t1 14.282
R252 a_1917_990.n1 a_1917_990.t0 14.282
R253 a_2332_101.t0 a_2332_101.n1 34.62
R254 a_2332_101.t0 a_2332_101.n0 8.137
R255 a_2332_101.t0 a_2332_101.n2 4.69
R256 A.n2 A.t8 512.525
R257 A.n5 A.t1 480.392
R258 A.n0 A.t0 480.392
R259 A.n5 A.t6 403.272
R260 A.n0 A.t7 403.272
R261 A.n2 A.t2 371.139
R262 A.n6 A.t3 336.586
R263 A.n1 A.t4 336.586
R264 A.n3 A.t5 290.093
R265 A.n3 A.n2 93.541
R266 A.n4 A.n1 77.859
R267 A.n4 A.n3 76
R268 A.n7 A.n6 76
R269 A.n1 A.n0 45.7
R270 A.n6 A.n5 45.341
R271 A.n7 A.n4 3.763
R272 A.n7 A 0.046
R273 VDD.n239 VDD.n237 144.705
R274 VDD.n264 VDD.n262 144.705
R275 VDD.n126 VDD.n124 144.705
R276 VDD.n331 VDD.n329 144.705
R277 VDD.n68 VDD.n66 144.705
R278 VDD.n26 VDD.n25 77.792
R279 VDD.n35 VDD.n34 77.792
R280 VDD.n300 VDD.n299 77.792
R281 VDD.n290 VDD.n289 77.792
R282 VDD.n254 VDD.n253 77.792
R283 VDD.n243 VDD.n242 77.792
R284 VDD.n29 VDD.n23 76.145
R285 VDD.n29 VDD.n28 76
R286 VDD.n33 VDD.n32 76
R287 VDD.n39 VDD.n38 76
R288 VDD.n43 VDD.n42 76
R289 VDD.n70 VDD.n69 76
R290 VDD.n74 VDD.n73 76
R291 VDD.n78 VDD.n77 76
R292 VDD.n82 VDD.n81 76
R293 VDD.n87 VDD.n86 76
R294 VDD.n94 VDD.n93 76
R295 VDD.n98 VDD.n97 76
R296 VDD.n102 VDD.n101 76
R297 VDD.n128 VDD.n127 76
R298 VDD.n132 VDD.n131 76
R299 VDD.n136 VDD.n135 76
R300 VDD.n140 VDD.n139 76
R301 VDD.n145 VDD.n144 76
R302 VDD.n152 VDD.n151 76
R303 VDD.n156 VDD.n155 76
R304 VDD.n333 VDD.n332 76
R305 VDD.n307 VDD.n306 76
R306 VDD.n303 VDD.n302 76
R307 VDD.n297 VDD.n296 76
R308 VDD.n293 VDD.n292 76
R309 VDD.n287 VDD.n286 76
R310 VDD.n261 VDD.n260 76
R311 VDD.n257 VDD.n256 76
R312 VDD.n251 VDD.n250 76
R313 VDD.n247 VDD.n246 76
R314 VDD.n241 VDD.n240 76
R315 VDD.n214 VDD.n213 76
R316 VDD.n210 VDD.n209 76
R317 VDD.n205 VDD.n204 76
R318 VDD.n200 VDD.n199 76
R319 VDD.n194 VDD.n193 76
R320 VDD.n189 VDD.n188 76
R321 VDD.n184 VDD.n183 76
R322 VDD.n179 VDD.n178 76
R323 VDD.n147 VDD.n146 65.585
R324 VDD.n89 VDD.n88 65.585
R325 VDD.n180 VDD.t12 55.106
R326 VDD.n245 VDD.t3 55.106
R327 VDD.n252 VDD.t2 55.106
R328 VDD.n288 VDD.t10 55.106
R329 VDD.n298 VDD.t9 55.106
R330 VDD.n37 VDD.t4 55.106
R331 VDD.n24 VDD.t5 55.106
R332 VDD.n206 VDD.t6 55.106
R333 VDD.n196 VDD.n195 40.824
R334 VDD.n269 VDD.n268 36.774
R335 VDD.n312 VDD.n311 36.774
R336 VDD.n107 VDD.n106 36.774
R337 VDD.n48 VDD.n47 36.774
R338 VDD.n230 VDD.n229 36.774
R339 VDD.n202 VDD.n201 36.608
R340 VDD.n91 VDD.n90 32.032
R341 VDD.n149 VDD.n148 32.032
R342 VDD.n186 VDD.n185 32.032
R343 VDD.n178 VDD.n175 21.841
R344 VDD.n23 VDD.n20 21.841
R345 VDD.n195 VDD.t0 14.282
R346 VDD.n195 VDD.t13 14.282
R347 VDD.n146 VDD.t8 14.282
R348 VDD.n146 VDD.t11 14.282
R349 VDD.n88 VDD.t1 14.282
R350 VDD.n88 VDD.t7 14.282
R351 VDD.n175 VDD.n158 14.167
R352 VDD.n158 VDD.n157 14.167
R353 VDD.n284 VDD.n266 14.167
R354 VDD.n266 VDD.n265 14.167
R355 VDD.n327 VDD.n309 14.167
R356 VDD.n309 VDD.n308 14.167
R357 VDD.n122 VDD.n104 14.167
R358 VDD.n104 VDD.n103 14.167
R359 VDD.n64 VDD.n45 14.167
R360 VDD.n45 VDD.n44 14.167
R361 VDD.n235 VDD.n216 14.167
R362 VDD.n216 VDD.n215 14.167
R363 VDD.n20 VDD.n19 14.167
R364 VDD.n19 VDD.n17 14.167
R365 VDD.n69 VDD.n65 14.167
R366 VDD.n127 VDD.n123 14.167
R367 VDD.n332 VDD.n328 14.167
R368 VDD.n286 VDD.n285 14.167
R369 VDD.n240 VDD.n236 14.167
R370 VDD.n23 VDD.n22 13.653
R371 VDD.n22 VDD.n21 13.653
R372 VDD.n28 VDD.n27 13.653
R373 VDD.n27 VDD.n26 13.653
R374 VDD.n32 VDD.n31 13.653
R375 VDD.n31 VDD.n30 13.653
R376 VDD.n38 VDD.n36 13.653
R377 VDD.n36 VDD.n35 13.653
R378 VDD.n42 VDD.n41 13.653
R379 VDD.n41 VDD.n40 13.653
R380 VDD.n69 VDD.n68 13.653
R381 VDD.n68 VDD.n67 13.653
R382 VDD.n73 VDD.n72 13.653
R383 VDD.n72 VDD.n71 13.653
R384 VDD.n77 VDD.n76 13.653
R385 VDD.n76 VDD.n75 13.653
R386 VDD.n81 VDD.n80 13.653
R387 VDD.n80 VDD.n79 13.653
R388 VDD.n86 VDD.n85 13.653
R389 VDD.n85 VDD.n84 13.653
R390 VDD.n93 VDD.n92 13.653
R391 VDD.n92 VDD.n91 13.653
R392 VDD.n97 VDD.n96 13.653
R393 VDD.n96 VDD.n95 13.653
R394 VDD.n101 VDD.n100 13.653
R395 VDD.n100 VDD.n99 13.653
R396 VDD.n127 VDD.n126 13.653
R397 VDD.n126 VDD.n125 13.653
R398 VDD.n131 VDD.n130 13.653
R399 VDD.n130 VDD.n129 13.653
R400 VDD.n135 VDD.n134 13.653
R401 VDD.n134 VDD.n133 13.653
R402 VDD.n139 VDD.n138 13.653
R403 VDD.n138 VDD.n137 13.653
R404 VDD.n144 VDD.n143 13.653
R405 VDD.n143 VDD.n142 13.653
R406 VDD.n151 VDD.n150 13.653
R407 VDD.n150 VDD.n149 13.653
R408 VDD.n155 VDD.n154 13.653
R409 VDD.n154 VDD.n153 13.653
R410 VDD.n332 VDD.n331 13.653
R411 VDD.n331 VDD.n330 13.653
R412 VDD.n306 VDD.n305 13.653
R413 VDD.n305 VDD.n304 13.653
R414 VDD.n302 VDD.n301 13.653
R415 VDD.n301 VDD.n300 13.653
R416 VDD.n296 VDD.n295 13.653
R417 VDD.n295 VDD.n294 13.653
R418 VDD.n292 VDD.n291 13.653
R419 VDD.n291 VDD.n290 13.653
R420 VDD.n286 VDD.n264 13.653
R421 VDD.n264 VDD.n263 13.653
R422 VDD.n260 VDD.n259 13.653
R423 VDD.n259 VDD.n258 13.653
R424 VDD.n256 VDD.n255 13.653
R425 VDD.n255 VDD.n254 13.653
R426 VDD.n250 VDD.n249 13.653
R427 VDD.n249 VDD.n248 13.653
R428 VDD.n246 VDD.n244 13.653
R429 VDD.n244 VDD.n243 13.653
R430 VDD.n240 VDD.n239 13.653
R431 VDD.n239 VDD.n238 13.653
R432 VDD.n213 VDD.n212 13.653
R433 VDD.n212 VDD.n211 13.653
R434 VDD.n209 VDD.n208 13.653
R435 VDD.n208 VDD.n207 13.653
R436 VDD.n204 VDD.n203 13.653
R437 VDD.n203 VDD.n202 13.653
R438 VDD.n199 VDD.n198 13.653
R439 VDD.n198 VDD.n197 13.653
R440 VDD.n193 VDD.n192 13.653
R441 VDD.n192 VDD.n191 13.653
R442 VDD.n188 VDD.n187 13.653
R443 VDD.n187 VDD.n186 13.653
R444 VDD.n183 VDD.n182 13.653
R445 VDD.n182 VDD.n181 13.653
R446 VDD.n178 VDD.n177 13.653
R447 VDD.n177 VDD.n176 13.653
R448 VDD.n4 VDD.n2 12.915
R449 VDD.n4 VDD.n3 12.66
R450 VDD.n13 VDD.n12 12.343
R451 VDD.n11 VDD.n10 12.343
R452 VDD.n7 VDD.n6 12.343
R453 VDD.n199 VDD.n196 8.658
R454 VDD.n285 VDD.n284 7.674
R455 VDD.n328 VDD.n327 7.674
R456 VDD.n123 VDD.n122 7.674
R457 VDD.n65 VDD.n64 7.674
R458 VDD.n236 VDD.n235 7.674
R459 VDD.n59 VDD.n58 7.5
R460 VDD.n53 VDD.n52 7.5
R461 VDD.n55 VDD.n54 7.5
R462 VDD.n50 VDD.n49 7.5
R463 VDD.n64 VDD.n63 7.5
R464 VDD.n117 VDD.n116 7.5
R465 VDD.n111 VDD.n110 7.5
R466 VDD.n113 VDD.n112 7.5
R467 VDD.n119 VDD.n109 7.5
R468 VDD.n119 VDD.n107 7.5
R469 VDD.n122 VDD.n121 7.5
R470 VDD.n322 VDD.n321 7.5
R471 VDD.n316 VDD.n315 7.5
R472 VDD.n318 VDD.n317 7.5
R473 VDD.n324 VDD.n314 7.5
R474 VDD.n324 VDD.n312 7.5
R475 VDD.n327 VDD.n326 7.5
R476 VDD.n279 VDD.n278 7.5
R477 VDD.n273 VDD.n272 7.5
R478 VDD.n275 VDD.n274 7.5
R479 VDD.n281 VDD.n271 7.5
R480 VDD.n281 VDD.n269 7.5
R481 VDD.n284 VDD.n283 7.5
R482 VDD.n220 VDD.n219 7.5
R483 VDD.n223 VDD.n222 7.5
R484 VDD.n225 VDD.n224 7.5
R485 VDD.n228 VDD.n227 7.5
R486 VDD.n235 VDD.n234 7.5
R487 VDD.n170 VDD.n169 7.5
R488 VDD.n164 VDD.n163 7.5
R489 VDD.n166 VDD.n165 7.5
R490 VDD.n172 VDD.n162 7.5
R491 VDD.n172 VDD.n160 7.5
R492 VDD.n175 VDD.n174 7.5
R493 VDD.n20 VDD.n16 7.5
R494 VDD.n2 VDD.n1 7.5
R495 VDD.n6 VDD.n5 7.5
R496 VDD.n10 VDD.n9 7.5
R497 VDD.n19 VDD.n18 7.5
R498 VDD.n14 VDD.n0 7.5
R499 VDD.n51 VDD.n48 6.772
R500 VDD.n62 VDD.n46 6.772
R501 VDD.n60 VDD.n57 6.772
R502 VDD.n56 VDD.n53 6.772
R503 VDD.n120 VDD.n105 6.772
R504 VDD.n118 VDD.n115 6.772
R505 VDD.n114 VDD.n111 6.772
R506 VDD.n325 VDD.n310 6.772
R507 VDD.n323 VDD.n320 6.772
R508 VDD.n319 VDD.n316 6.772
R509 VDD.n282 VDD.n267 6.772
R510 VDD.n280 VDD.n277 6.772
R511 VDD.n276 VDD.n273 6.772
R512 VDD.n173 VDD.n159 6.772
R513 VDD.n171 VDD.n168 6.772
R514 VDD.n167 VDD.n164 6.772
R515 VDD.n51 VDD.n50 6.772
R516 VDD.n56 VDD.n55 6.772
R517 VDD.n60 VDD.n59 6.772
R518 VDD.n63 VDD.n62 6.772
R519 VDD.n114 VDD.n113 6.772
R520 VDD.n118 VDD.n117 6.772
R521 VDD.n121 VDD.n120 6.772
R522 VDD.n319 VDD.n318 6.772
R523 VDD.n323 VDD.n322 6.772
R524 VDD.n326 VDD.n325 6.772
R525 VDD.n276 VDD.n275 6.772
R526 VDD.n280 VDD.n279 6.772
R527 VDD.n283 VDD.n282 6.772
R528 VDD.n167 VDD.n166 6.772
R529 VDD.n171 VDD.n170 6.772
R530 VDD.n174 VDD.n173 6.772
R531 VDD.n234 VDD.n233 6.772
R532 VDD.n221 VDD.n218 6.772
R533 VDD.n226 VDD.n223 6.772
R534 VDD.n231 VDD.n228 6.772
R535 VDD.n231 VDD.n230 6.772
R536 VDD.n226 VDD.n225 6.772
R537 VDD.n221 VDD.n220 6.772
R538 VDD.n233 VDD.n217 6.772
R539 VDD.n16 VDD.n15 6.458
R540 VDD.n109 VDD.n108 6.202
R541 VDD.n314 VDD.n313 6.202
R542 VDD.n271 VDD.n270 6.202
R543 VDD.n162 VDD.n161 6.202
R544 VDD.n93 VDD.n89 5.903
R545 VDD.n151 VDD.n147 5.903
R546 VDD.n84 VDD.n83 4.576
R547 VDD.n142 VDD.n141 4.576
R548 VDD.n191 VDD.n190 4.576
R549 VDD.n183 VDD.n180 2.754
R550 VDD.n209 VDD.n206 2.361
R551 VDD.n28 VDD.n24 1.967
R552 VDD.n38 VDD.n37 1.967
R553 VDD.n302 VDD.n298 1.967
R554 VDD.n292 VDD.n288 1.967
R555 VDD.n256 VDD.n252 1.967
R556 VDD.n246 VDD.n245 1.967
R557 VDD.n14 VDD.n7 1.329
R558 VDD.n14 VDD.n8 1.329
R559 VDD.n14 VDD.n11 1.329
R560 VDD.n14 VDD.n13 1.329
R561 VDD.n15 VDD.n14 0.696
R562 VDD.n14 VDD.n4 0.696
R563 VDD.n61 VDD.n60 0.365
R564 VDD.n61 VDD.n56 0.365
R565 VDD.n61 VDD.n51 0.365
R566 VDD.n62 VDD.n61 0.365
R567 VDD.n119 VDD.n118 0.365
R568 VDD.n119 VDD.n114 0.365
R569 VDD.n120 VDD.n119 0.365
R570 VDD.n324 VDD.n323 0.365
R571 VDD.n324 VDD.n319 0.365
R572 VDD.n325 VDD.n324 0.365
R573 VDD.n281 VDD.n280 0.365
R574 VDD.n281 VDD.n276 0.365
R575 VDD.n282 VDD.n281 0.365
R576 VDD.n172 VDD.n171 0.365
R577 VDD.n172 VDD.n167 0.365
R578 VDD.n173 VDD.n172 0.365
R579 VDD.n232 VDD.n231 0.365
R580 VDD.n232 VDD.n226 0.365
R581 VDD.n232 VDD.n221 0.365
R582 VDD.n233 VDD.n232 0.365
R583 VDD.n70 VDD.n43 0.29
R584 VDD.n128 VDD.n102 0.29
R585 VDD.n333 VDD.n307 0.29
R586 VDD.n287 VDD.n261 0.29
R587 VDD.n241 VDD.n214 0.29
R588 VDD.n179 VDD 0.207
R589 VDD.n87 VDD.n82 0.181
R590 VDD.n145 VDD.n140 0.181
R591 VDD.n200 VDD.n194 0.181
R592 VDD.n33 VDD.n29 0.157
R593 VDD.n39 VDD.n33 0.157
R594 VDD.n303 VDD.n297 0.157
R595 VDD.n297 VDD.n293 0.157
R596 VDD.n257 VDD.n251 0.157
R597 VDD.n251 VDD.n247 0.157
R598 VDD.n43 VDD.n39 0.145
R599 VDD.n74 VDD.n70 0.145
R600 VDD.n78 VDD.n74 0.145
R601 VDD.n82 VDD.n78 0.145
R602 VDD.n94 VDD.n87 0.145
R603 VDD.n98 VDD.n94 0.145
R604 VDD.n102 VDD.n98 0.145
R605 VDD.n132 VDD.n128 0.145
R606 VDD.n136 VDD.n132 0.145
R607 VDD.n140 VDD.n136 0.145
R608 VDD.n152 VDD.n145 0.145
R609 VDD.n156 VDD.n152 0.145
R610 VDD.n307 VDD.n303 0.145
R611 VDD.n293 VDD.n287 0.145
R612 VDD.n261 VDD.n257 0.145
R613 VDD.n247 VDD.n241 0.145
R614 VDD.n214 VDD.n210 0.145
R615 VDD.n210 VDD.n205 0.145
R616 VDD.n205 VDD.n200 0.145
R617 VDD.n194 VDD.n189 0.145
R618 VDD.n189 VDD.n184 0.145
R619 VDD.n184 VDD.n179 0.145
R620 VDD VDD.n333 0.078
R621 VDD VDD.n156 0.066
R622 a_1685_1051.t1 a_1685_1051.n0 101.663
R623 a_1685_1051.n0 a_1685_1051.t2 101.661
R624 a_1685_1051.n0 a_1685_1051.t0 14.294
R625 a_1685_1051.n0 a_1685_1051.t3 14.282
R626 B.n0 B.t7 512.525
R627 B.n3 B.t6 480.392
R628 B.n5 B.t2 472.359
R629 B.n3 B.t0 403.272
R630 B.n5 B.t5 384.527
R631 B.n1 B.t8 372.349
R632 B.n0 B.t3 371.139
R633 B.n6 B.t4 241.172
R634 B.n7 B.n4 212.632
R635 B.n1 B.t1 157.328
R636 B.n2 B.n1 132.764
R637 B.n4 B.n3 121.7
R638 B.n6 B.n5 110.06
R639 B.n2 B.n0 93.541
R640 B.n4 B.n2 78.675
R641 B.n7 B.n6 76
R642 B.n7 B 0.046
R643 a_112_101.t0 a_112_101.n1 34.62
R644 a_112_101.t0 a_112_101.n0 8.137
R645 a_112_101.t0 a_112_101.n2 4.69
R646 a_1666_101.t0 a_1666_101.n1 34.62
R647 a_1666_101.t0 a_1666_101.n0 8.137
R648 a_1666_101.t0 a_1666_101.n2 4.69
C9 VDD GND 13.28fF
C10 a_1666_101.n0 GND 0.05fF
C11 a_1666_101.n1 GND 0.12fF
C12 a_1666_101.n2 GND 0.04fF
C13 a_112_101.n0 GND 0.05fF
C14 a_112_101.n1 GND 0.12fF
C15 a_112_101.n2 GND 0.04fF
C16 a_1685_1051.n0 GND 0.52fF
C17 VDD.n0 GND 0.12fF
C18 VDD.n1 GND 0.03fF
C19 VDD.n2 GND 0.02fF
C20 VDD.n3 GND 0.05fF
C21 VDD.n4 GND 0.01fF
C22 VDD.n5 GND 0.02fF
C23 VDD.n6 GND 0.02fF
C24 VDD.n9 GND 0.02fF
C25 VDD.n10 GND 0.02fF
C26 VDD.n12 GND 0.02fF
C27 VDD.n14 GND 0.46fF
C28 VDD.n16 GND 0.03fF
C29 VDD.n17 GND 0.02fF
C30 VDD.n18 GND 0.02fF
C31 VDD.n19 GND 0.02fF
C32 VDD.n20 GND 0.04fF
C33 VDD.n21 GND 0.27fF
C34 VDD.n22 GND 0.02fF
C35 VDD.n23 GND 0.03fF
C36 VDD.n24 GND 0.06fF
C37 VDD.n25 GND 0.15fF
C38 VDD.n26 GND 0.20fF
C39 VDD.n27 GND 0.01fF
C40 VDD.n28 GND 0.01fF
C41 VDD.n29 GND 0.07fF
C42 VDD.n30 GND 0.17fF
C43 VDD.n31 GND 0.01fF
C44 VDD.n32 GND 0.02fF
C45 VDD.n33 GND 0.02fF
C46 VDD.n34 GND 0.15fF
C47 VDD.n35 GND 0.20fF
C48 VDD.n36 GND 0.01fF
C49 VDD.n37 GND 0.06fF
C50 VDD.n38 GND 0.01fF
C51 VDD.n39 GND 0.02fF
C52 VDD.n40 GND 0.27fF
C53 VDD.n41 GND 0.01fF
C54 VDD.n42 GND 0.02fF
C55 VDD.n43 GND 0.03fF
C56 VDD.n44 GND 0.02fF
C57 VDD.n45 GND 0.02fF
C58 VDD.n46 GND 0.02fF
C59 VDD.n47 GND 0.18fF
C60 VDD.n48 GND 0.04fF
C61 VDD.n49 GND 0.04fF
C62 VDD.n50 GND 0.02fF
C63 VDD.n52 GND 0.02fF
C64 VDD.n53 GND 0.02fF
C65 VDD.n54 GND 0.02fF
C66 VDD.n55 GND 0.02fF
C67 VDD.n57 GND 0.02fF
C68 VDD.n58 GND 0.02fF
C69 VDD.n59 GND 0.02fF
C70 VDD.n61 GND 0.27fF
C71 VDD.n63 GND 0.02fF
C72 VDD.n64 GND 0.02fF
C73 VDD.n65 GND 0.03fF
C74 VDD.n66 GND 0.02fF
C75 VDD.n67 GND 0.27fF
C76 VDD.n68 GND 0.01fF
C77 VDD.n69 GND 0.02fF
C78 VDD.n70 GND 0.03fF
C79 VDD.n71 GND 0.27fF
C80 VDD.n72 GND 0.01fF
C81 VDD.n73 GND 0.02fF
C82 VDD.n74 GND 0.02fF
C83 VDD.n75 GND 0.27fF
C84 VDD.n76 GND 0.01fF
C85 VDD.n77 GND 0.02fF
C86 VDD.n78 GND 0.02fF
C87 VDD.n79 GND 0.30fF
C88 VDD.n80 GND 0.01fF
C89 VDD.n81 GND 0.03fF
C90 VDD.n82 GND 0.03fF
C91 VDD.n83 GND 0.17fF
C92 VDD.n84 GND 0.14fF
C93 VDD.n85 GND 0.01fF
C94 VDD.n86 GND 0.02fF
C95 VDD.n87 GND 0.03fF
C96 VDD.n88 GND 0.10fF
C97 VDD.n89 GND 0.03fF
C98 VDD.n90 GND 0.14fF
C99 VDD.n91 GND 0.16fF
C100 VDD.n92 GND 0.01fF
C101 VDD.n93 GND 0.02fF
C102 VDD.n94 GND 0.02fF
C103 VDD.n95 GND 0.25fF
C104 VDD.n96 GND 0.01fF
C105 VDD.n97 GND 0.02fF
C106 VDD.n98 GND 0.02fF
C107 VDD.n99 GND 0.27fF
C108 VDD.n100 GND 0.01fF
C109 VDD.n101 GND 0.02fF
C110 VDD.n102 GND 0.03fF
C111 VDD.n103 GND 0.02fF
C112 VDD.n104 GND 0.02fF
C113 VDD.n105 GND 0.02fF
C114 VDD.n106 GND 0.21fF
C115 VDD.n107 GND 0.04fF
C116 VDD.n108 GND 0.03fF
C117 VDD.n109 GND 0.02fF
C118 VDD.n110 GND 0.02fF
C119 VDD.n111 GND 0.02fF
C120 VDD.n112 GND 0.03fF
C121 VDD.n113 GND 0.02fF
C122 VDD.n115 GND 0.02fF
C123 VDD.n116 GND 0.02fF
C124 VDD.n117 GND 0.02fF
C125 VDD.n119 GND 0.27fF
C126 VDD.n121 GND 0.02fF
C127 VDD.n122 GND 0.02fF
C128 VDD.n123 GND 0.03fF
C129 VDD.n124 GND 0.02fF
C130 VDD.n125 GND 0.27fF
C131 VDD.n126 GND 0.01fF
C132 VDD.n127 GND 0.02fF
C133 VDD.n128 GND 0.03fF
C134 VDD.n129 GND 0.27fF
C135 VDD.n130 GND 0.01fF
C136 VDD.n131 GND 0.02fF
C137 VDD.n132 GND 0.02fF
C138 VDD.n133 GND 0.27fF
C139 VDD.n134 GND 0.01fF
C140 VDD.n135 GND 0.02fF
C141 VDD.n136 GND 0.02fF
C142 VDD.n137 GND 0.30fF
C143 VDD.n138 GND 0.01fF
C144 VDD.n139 GND 0.03fF
C145 VDD.n140 GND 0.03fF
C146 VDD.n141 GND 0.17fF
C147 VDD.n142 GND 0.14fF
C148 VDD.n143 GND 0.01fF
C149 VDD.n144 GND 0.02fF
C150 VDD.n145 GND 0.03fF
C151 VDD.n146 GND 0.10fF
C152 VDD.n147 GND 0.03fF
C153 VDD.n148 GND 0.14fF
C154 VDD.n149 GND 0.16fF
C155 VDD.n150 GND 0.01fF
C156 VDD.n151 GND 0.02fF
C157 VDD.n152 GND 0.02fF
C158 VDD.n153 GND 0.25fF
C159 VDD.n154 GND 0.01fF
C160 VDD.n155 GND 0.02fF
C161 VDD.n156 GND 0.02fF
C162 VDD.n157 GND 0.02fF
C163 VDD.n158 GND 0.02fF
C164 VDD.n159 GND 0.02fF
C165 VDD.n160 GND 0.15fF
C166 VDD.n161 GND 0.03fF
C167 VDD.n162 GND 0.02fF
C168 VDD.n163 GND 0.02fF
C169 VDD.n164 GND 0.02fF
C170 VDD.n165 GND 0.03fF
C171 VDD.n166 GND 0.02fF
C172 VDD.n168 GND 0.02fF
C173 VDD.n169 GND 0.02fF
C174 VDD.n170 GND 0.02fF
C175 VDD.n172 GND 0.46fF
C176 VDD.n174 GND 0.03fF
C177 VDD.n175 GND 0.04fF
C178 VDD.n176 GND 0.27fF
C179 VDD.n177 GND 0.02fF
C180 VDD.n178 GND 0.03fF
C181 VDD.n179 GND 0.03fF
C182 VDD.n180 GND 0.06fF
C183 VDD.n181 GND 0.25fF
C184 VDD.n182 GND 0.01fF
C185 VDD.n183 GND 0.01fF
C186 VDD.n184 GND 0.02fF
C187 VDD.n185 GND 0.14fF
C188 VDD.n186 GND 0.16fF
C189 VDD.n187 GND 0.01fF
C190 VDD.n188 GND 0.02fF
C191 VDD.n189 GND 0.02fF
C192 VDD.n190 GND 0.17fF
C193 VDD.n191 GND 0.14fF
C194 VDD.n192 GND 0.01fF
C195 VDD.n193 GND 0.02fF
C196 VDD.n194 GND 0.03fF
C197 VDD.n195 GND 0.11fF
C198 VDD.n196 GND 0.03fF
C199 VDD.n197 GND 0.30fF
C200 VDD.n198 GND 0.01fF
C201 VDD.n199 GND 0.02fF
C202 VDD.n200 GND 0.03fF
C203 VDD.n201 GND 0.14fF
C204 VDD.n202 GND 0.17fF
C205 VDD.n203 GND 0.01fF
C206 VDD.n204 GND 0.02fF
C207 VDD.n205 GND 0.02fF
C208 VDD.n206 GND 0.06fF
C209 VDD.n207 GND 0.24fF
C210 VDD.n208 GND 0.01fF
C211 VDD.n209 GND 0.01fF
C212 VDD.n210 GND 0.02fF
C213 VDD.n211 GND 0.27fF
C214 VDD.n212 GND 0.01fF
C215 VDD.n213 GND 0.02fF
C216 VDD.n214 GND 0.03fF
C217 VDD.n215 GND 0.02fF
C218 VDD.n216 GND 0.02fF
C219 VDD.n217 GND 0.02fF
C220 VDD.n218 GND 0.02fF
C221 VDD.n219 GND 0.02fF
C222 VDD.n220 GND 0.02fF
C223 VDD.n222 GND 0.02fF
C224 VDD.n223 GND 0.02fF
C225 VDD.n224 GND 0.02fF
C226 VDD.n225 GND 0.02fF
C227 VDD.n227 GND 0.04fF
C228 VDD.n228 GND 0.02fF
C229 VDD.n229 GND 0.18fF
C230 VDD.n230 GND 0.04fF
C231 VDD.n232 GND 0.27fF
C232 VDD.n234 GND 0.02fF
C233 VDD.n235 GND 0.02fF
C234 VDD.n236 GND 0.03fF
C235 VDD.n237 GND 0.02fF
C236 VDD.n238 GND 0.27fF
C237 VDD.n239 GND 0.01fF
C238 VDD.n240 GND 0.02fF
C239 VDD.n241 GND 0.03fF
C240 VDD.n242 GND 0.15fF
C241 VDD.n243 GND 0.20fF
C242 VDD.n244 GND 0.01fF
C243 VDD.n245 GND 0.06fF
C244 VDD.n246 GND 0.01fF
C245 VDD.n247 GND 0.02fF
C246 VDD.n248 GND 0.17fF
C247 VDD.n249 GND 0.01fF
C248 VDD.n250 GND 0.02fF
C249 VDD.n251 GND 0.02fF
C250 VDD.n252 GND 0.06fF
C251 VDD.n253 GND 0.15fF
C252 VDD.n254 GND 0.20fF
C253 VDD.n255 GND 0.01fF
C254 VDD.n256 GND 0.01fF
C255 VDD.n257 GND 0.02fF
C256 VDD.n258 GND 0.27fF
C257 VDD.n259 GND 0.01fF
C258 VDD.n260 GND 0.02fF
C259 VDD.n261 GND 0.03fF
C260 VDD.n262 GND 0.02fF
C261 VDD.n263 GND 0.27fF
C262 VDD.n264 GND 0.01fF
C263 VDD.n265 GND 0.02fF
C264 VDD.n266 GND 0.02fF
C265 VDD.n267 GND 0.02fF
C266 VDD.n268 GND 0.14fF
C267 VDD.n269 GND 0.04fF
C268 VDD.n270 GND 0.03fF
C269 VDD.n271 GND 0.02fF
C270 VDD.n272 GND 0.02fF
C271 VDD.n273 GND 0.02fF
C272 VDD.n274 GND 0.03fF
C273 VDD.n275 GND 0.02fF
C274 VDD.n277 GND 0.02fF
C275 VDD.n278 GND 0.02fF
C276 VDD.n279 GND 0.02fF
C277 VDD.n281 GND 0.27fF
C278 VDD.n283 GND 0.02fF
C279 VDD.n284 GND 0.02fF
C280 VDD.n285 GND 0.03fF
C281 VDD.n286 GND 0.02fF
C282 VDD.n287 GND 0.03fF
C283 VDD.n288 GND 0.06fF
C284 VDD.n289 GND 0.15fF
C285 VDD.n290 GND 0.20fF
C286 VDD.n291 GND 0.01fF
C287 VDD.n292 GND 0.01fF
C288 VDD.n293 GND 0.02fF
C289 VDD.n294 GND 0.17fF
C290 VDD.n295 GND 0.01fF
C291 VDD.n296 GND 0.02fF
C292 VDD.n297 GND 0.02fF
C293 VDD.n298 GND 0.06fF
C294 VDD.n299 GND 0.15fF
C295 VDD.n300 GND 0.20fF
C296 VDD.n301 GND 0.01fF
C297 VDD.n302 GND 0.01fF
C298 VDD.n303 GND 0.02fF
C299 VDD.n304 GND 0.27fF
C300 VDD.n305 GND 0.01fF
C301 VDD.n306 GND 0.02fF
C302 VDD.n307 GND 0.03fF
C303 VDD.n308 GND 0.02fF
C304 VDD.n309 GND 0.02fF
C305 VDD.n310 GND 0.02fF
C306 VDD.n311 GND 0.18fF
C307 VDD.n312 GND 0.04fF
C308 VDD.n313 GND 0.03fF
C309 VDD.n314 GND 0.02fF
C310 VDD.n315 GND 0.02fF
C311 VDD.n316 GND 0.02fF
C312 VDD.n317 GND 0.03fF
C313 VDD.n318 GND 0.02fF
C314 VDD.n320 GND 0.02fF
C315 VDD.n321 GND 0.02fF
C316 VDD.n322 GND 0.02fF
C317 VDD.n324 GND 0.27fF
C318 VDD.n326 GND 0.02fF
C319 VDD.n327 GND 0.02fF
C320 VDD.n328 GND 0.03fF
C321 VDD.n329 GND 0.02fF
C322 VDD.n330 GND 0.27fF
C323 VDD.n331 GND 0.01fF
C324 VDD.n332 GND 0.02fF
C325 VDD.n333 GND 0.03fF
C326 a_2332_101.n0 GND 0.05fF
C327 a_2332_101.n1 GND 0.12fF
C328 a_2332_101.n2 GND 0.04fF
C329 a_1917_990.n0 GND 0.07fF
C330 a_1917_990.n1 GND 1.16fF
C331 a_1917_990.n2 GND 1.22fF
C332 a_1917_990.n3 GND 1.48fF
C333 a_1917_990.n4 GND 1.43fF
C334 a_1917_990.n5 GND 0.07fF
C335 a_1917_990.n6 GND 0.38fF
C336 a_1917_990.n7 GND 0.08fF
C337 a_2351_1051.n0 GND 0.52fF
C338 SUM.n0 GND 1.15fF
C339 SUM.n1 GND 0.07fF
C340 SUM.n2 GND 0.09fF
C341 SUM.n3 GND 0.06fF
C342 SUM.n4 GND 0.51fF
C343 SUM.n5 GND 0.76fF
C344 SUM.n6 GND 1.15fF
C345 SUM.n7 GND 0.68fF
C346 SUM.n8 GND 0.83fF
C347 SUM.n9 GND 0.05fF
C348 a_1295_209.n0 GND 1.13fF
C349 a_1295_209.n1 GND 0.61fF
C350 a_1295_209.n2 GND 1.41fF
C351 a_1295_209.n3 GND 1.48fF
C352 a_1295_209.n4 GND 0.12fF
C353 a_1295_209.n5 GND 0.37fF
C354 a_1295_209.n6 GND 0.07fF
C355 a_217_1050.n0 GND 0.48fF
C356 a_217_1050.n1 GND 0.57fF
C357 a_217_1050.n2 GND 0.31fF
C358 a_217_1050.n3 GND 0.34fF
C359 a_217_1050.n4 GND 0.53fF
C360 a_217_1050.n5 GND 0.53fF
C361 a_217_1050.n6 GND 0.08fF
C362 a_217_1050.n7 GND 0.23fF
C363 a_217_1050.n8 GND 0.04fF
.ends
