// File: nmos_side_right.spi.NMOS_SIDE_RIGHT.pxi
// Created: Tue Oct 15 15:58:31 2024
// 
simulator lang=spectre
cc_1 ( noxref_1 noxref_2 ) capacitor c=0.0464957f //x=0.435 //y=0.535 //x2=0 \
 //y2=0
cc_2 ( noxref_1 noxref_3 ) capacitor c=0.0254606f //x=0.435 //y=0.535 \
 //x2=0.622 //y2=0.925
cc_3 ( noxref_2 noxref_3 ) capacitor c=0.096254f //x=0 //y=0 //x2=0.622 \
 //y2=0.925
