// File: MUX2X1.spi.pex
// Created: Tue Oct 15 15:49:38 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_MUX2X1\%GND ( 1 23 35 39 42 47 53 59 65 73 81 94 97 108 111 113 115 \
 116 117 118 )
c165 ( 118 0 ) capacitor c=0.0207871f //x=9.87 //y=0.865
c166 ( 117 0 ) capacitor c=0.0207873f //x=6.54 //y=0.865
c167 ( 116 0 ) capacitor c=0.0207871f //x=3.21 //y=0.865
c168 ( 115 0 ) capacitor c=0.0583152f //x=0.495 //y=0.37
c169 ( 114 0 ) capacitor c=0.00440095f //x=10.06 //y=0
c170 ( 113 0 ) capacitor c=0.106543f //x=8.88 //y=0
c171 ( 112 0 ) capacitor c=0.00440095f //x=6.73 //y=0
c172 ( 111 0 ) capacitor c=0.106543f //x=5.55 //y=0
c173 ( 110 0 ) capacitor c=0.00440095f //x=3.33 //y=0
c174 ( 108 0 ) capacitor c=0.102231f //x=2.22 //y=0
c175 ( 97 0 ) capacitor c=0.192978f //x=0.63 //y=0
c176 ( 94 0 ) capacitor c=0.259331f //x=11.47 //y=0
c177 ( 81 0 ) capacitor c=0.0389171f //x=9.975 //y=0
c178 ( 73 0 ) capacitor c=0.0718766f //x=8.71 //y=0
c179 ( 65 0 ) capacitor c=0.0389171f //x=6.645 //y=0
c180 ( 59 0 ) capacitor c=0.0720496f //x=5.38 //y=0
c181 ( 53 0 ) capacitor c=0.0389171f //x=3.315 //y=0
c182 ( 48 0 ) capacitor c=0.036088f //x=1.685 //y=0
c183 ( 47 0 ) capacitor c=0.0160123f //x=2.05 //y=0
c184 ( 42 0 ) capacitor c=0.00583665f //x=1.6 //y=0.45
c185 ( 39 0 ) capacitor c=0.00531808f //x=1.515 //y=0.535
c186 ( 38 0 ) capacitor c=0.00479856f //x=1.115 //y=0.45
c187 ( 35 0 ) capacitor c=0.00644318f //x=1.03 //y=0.535
c188 ( 30 0 ) capacitor c=0.00592191f //x=0.63 //y=0.45
c189 ( 23 0 ) capacitor c=0.424473f //x=11.47 //y=0
r190 (  100 101 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.115 //y=0 //x2=1.6 //y2=0
r191 (  99 100 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.115 //y2=0
r192 (  97 99 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=0.63 //y=0 //x2=0.74 //y2=0
r193 (  92 94 ) resistor r=26.5322 //w=0.357 //l=0.74 //layer=li \
 //thickness=0.1 //x=10.73 //y=0 //x2=11.47 //y2=0
r194 (  90 114 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.145 //y=0 //x2=10.06 //y2=0
r195 (  90 92 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=10.145 //y=0 //x2=10.73 //y2=0
r196 (  85 114 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.06 //y=0.17 //x2=10.06 //y2=0
r197 (  85 118 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=10.06 //y=0.17 //x2=10.06 //y2=0.955
r198 (  82 113 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.05 //y=0 //x2=8.88 //y2=0
r199 (  82 84 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.05 //y=0 //x2=9.62 //y2=0
r200 (  81 114 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.975 //y=0 //x2=10.06 //y2=0
r201 (  81 84 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=9.975 //y=0 //x2=9.62 //y2=0
r202 (  76 78 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.03 //y=0 //x2=8.14 //y2=0
r203 (  74 112 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.815 //y=0 //x2=6.73 //y2=0
r204 (  74 76 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=6.815 //y=0 //x2=7.03 //y2=0
r205 (  73 113 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.71 //y=0 //x2=8.88 //y2=0
r206 (  73 78 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.71 //y=0 //x2=8.14 //y2=0
r207 (  69 112 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.73 //y=0.17 //x2=6.73 //y2=0
r208 (  69 117 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=6.73 //y=0.17 //x2=6.73 //y2=0.955
r209 (  66 111 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.55 //y2=0
r210 (  66 68 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.92 //y2=0
r211 (  65 112 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.645 //y=0 //x2=6.73 //y2=0
r212 (  65 68 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=6.645 //y=0 //x2=5.92 //y2=0
r213 (  60 110 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.485 //y=0 //x2=3.4 //y2=0
r214 (  60 62 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=3.485 //y=0 //x2=4.44 //y2=0
r215 (  59 111 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=5.55 //y2=0
r216 (  59 62 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=4.44 //y2=0
r217 (  55 110 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.4 //y=0.17 //x2=3.4 //y2=0
r218 (  55 116 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=3.4 //y=0.17 //x2=3.4 //y2=0.955
r219 (  54 108 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.39 //y=0 //x2=2.22 //y2=0
r220 (  53 110 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.315 //y=0 //x2=3.4 //y2=0
r221 (  53 54 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=3.315 //y=0 //x2=2.39 //y2=0
r222 (  48 101 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.6 //y2=0
r223 (  48 50 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.85 //y2=0
r224 (  47 108 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=2.22 //y2=0
r225 (  47 50 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=1.85 //y2=0
r226 (  43 115 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=0.535
r227 (  43 115 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=1.225
r228 (  42 115 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.45 //x2=1.6 //y2=0.535
r229 (  41 101 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0
r230 (  41 42 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0.45
r231 (  40 115 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.2 //y=0.535 //x2=1.115 //y2=0.535
r232 (  39 115 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.6 //y2=0.535
r233 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.2 //y2=0.535
r234 (  38 115 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.45 //x2=1.115 //y2=0.535
r235 (  37 100 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0
r236 (  37 38 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0.45
r237 (  36 115 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.715 //y=0.535 //x2=0.63 //y2=0.535
r238 (  35 115 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=1.115 //y2=0.535
r239 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=0.715 //y2=0.535
r240 (  31 115 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=0.535
r241 (  31 115 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=1.225
r242 (  30 115 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.45 //x2=0.63 //y2=0.535
r243 (  29 97 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0
r244 (  29 30 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0.45
r245 (  23 94 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r246 (  21 92 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=0 //x2=10.73 //y2=0
r247 (  21 23 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=0 //x2=11.47 //y2=0
r248 (  19 84 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=0 //x2=9.62 //y2=0
r249 (  19 21 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.62 //y=0 //x2=10.73 //y2=0
r250 (  17 78 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=0 //x2=8.14 //y2=0
r251 (  17 19 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=0 //x2=9.62 //y2=0
r252 (  15 76 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=0 //x2=7.03 //y2=0
r253 (  15 17 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=0 //x2=8.14 //y2=0
r254 (  12 68 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=0 //x2=5.92 //y2=0
r255 (  10 62 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r256 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.92 //y2=0
r257 (  8 110 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=0 //x2=3.33 //y2=0
r258 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=0 //x2=4.44 //y2=0
r259 (  6 50 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r260 (  6 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=3.33 //y2=0
r261 (  3 99 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r262 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r263 (  1 15 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=6.105 //y=0 //x2=7.03 //y2=0
r264 (  1 12 ) resistor r=0.0768272 //w=0.301 //l=0.185 //layer=m1 \
 //thickness=0.36 //x=6.105 //y=0 //x2=5.92 //y2=0
ends PM_MUX2X1\%GND

subckt PM_MUX2X1\%VDD ( 1 23 35 57 67 91 101 121 129 144 146 150 155 160 161 \
 162 163 164 165 166 167 168 169 170 171 )
c163 ( 171 0 ) capacitor c=0.0383753f //x=11.285 //y=5.02
c164 ( 170 0 ) capacitor c=0.0241901f //x=10.405 //y=5.02
c165 ( 169 0 ) capacitor c=0.0499723f //x=9.535 //y=5.02
c166 ( 168 0 ) capacitor c=0.0382536f //x=7.955 //y=5.02
c167 ( 167 0 ) capacitor c=0.024222f //x=7.075 //y=5.02
c168 ( 166 0 ) capacitor c=0.0499723f //x=6.205 //y=5.02
c169 ( 165 0 ) capacitor c=0.0382565f //x=4.625 //y=5.02
c170 ( 164 0 ) capacitor c=0.0241904f //x=3.745 //y=5.02
c171 ( 163 0 ) capacitor c=0.0500634f //x=2.875 //y=5.02
c172 ( 162 0 ) capacitor c=0.0436617f //x=1.41 //y=5.02
c173 ( 161 0 ) capacitor c=0.0423206f //x=0.54 //y=5.02
c174 ( 160 0 ) capacitor c=0.243792f //x=11.47 //y=7.4
c175 ( 158 0 ) capacitor c=0.00591168f //x=10.55 //y=7.4
c176 ( 157 0 ) capacitor c=0.00591168f //x=9.62 //y=7.4
c177 ( 155 0 ) capacitor c=0.119448f //x=8.88 //y=7.4
c178 ( 154 0 ) capacitor c=0.00591168f //x=8.14 //y=7.4
c179 ( 152 0 ) capacitor c=0.00591168f //x=7.22 //y=7.4
c180 ( 151 0 ) capacitor c=0.00591168f //x=6.34 //y=7.4
c181 ( 150 0 ) capacitor c=0.119448f //x=5.55 //y=7.4
c182 ( 149 0 ) capacitor c=0.00591168f //x=4.77 //y=7.4
c183 ( 148 0 ) capacitor c=0.00591168f //x=3.89 //y=7.4
c184 ( 147 0 ) capacitor c=0.00591168f //x=3.01 //y=7.4
c185 ( 146 0 ) capacitor c=0.116993f //x=2.22 //y=7.4
c186 ( 145 0 ) capacitor c=0.00591168f //x=1.555 //y=7.4
c187 ( 144 0 ) capacitor c=0.233263f //x=0.74 //y=7.4
c188 ( 129 0 ) capacitor c=0.0285035f //x=11.345 //y=7.4
c189 ( 121 0 ) capacitor c=0.0286367f //x=10.465 //y=7.4
c190 ( 113 0 ) capacitor c=0.0281468f //x=9.585 //y=7.4
c191 ( 109 0 ) capacitor c=0.0275781f //x=8.71 //y=7.4
c192 ( 101 0 ) capacitor c=0.0285035f //x=8.015 //y=7.4
c193 ( 91 0 ) capacitor c=0.0286367f //x=7.135 //y=7.4
c194 ( 81 0 ) capacitor c=0.0281468f //x=6.255 //y=7.4
c195 ( 77 0 ) capacitor c=0.0275781f //x=5.38 //y=7.4
c196 ( 67 0 ) capacitor c=0.0285035f //x=4.685 //y=7.4
c197 ( 57 0 ) capacitor c=0.0286367f //x=3.805 //y=7.4
c198 ( 49 0 ) capacitor c=0.0281468f //x=2.925 //y=7.4
c199 ( 43 0 ) capacitor c=0.0210379f //x=2.05 //y=7.4
c200 ( 35 0 ) capacitor c=0.0287207f //x=1.47 //y=7.4
c201 ( 23 0 ) capacitor c=0.450693f //x=11.47 //y=7.4
r202 (  133 160 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.43 //y=7.23 //x2=11.43 //y2=7.4
r203 (  133 171 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.43 //y=7.23 //x2=11.43 //y2=6.745
r204 (  130 158 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.635 //y=7.4 //x2=10.55 //y2=7.4
r205 (  130 132 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=10.635 //y=7.4 //x2=10.73 //y2=7.4
r206 (  129 160 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.345 //y=7.4 //x2=11.43 //y2=7.4
r207 (  129 132 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=11.345 //y=7.4 //x2=10.73 //y2=7.4
r208 (  123 158 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.55 //y=7.23 //x2=10.55 //y2=7.4
r209 (  123 170 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.55 //y=7.23 //x2=10.55 //y2=6.745
r210 (  122 157 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.755 //y=7.4 //x2=9.67 //y2=7.4
r211 (  121 158 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.465 //y=7.4 //x2=10.55 //y2=7.4
r212 (  121 122 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.465 //y=7.4 //x2=9.755 //y2=7.4
r213 (  115 157 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.67 //y=7.23 //x2=9.67 //y2=7.4
r214 (  115 169 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=9.67 //y=7.23 //x2=9.67 //y2=6.405
r215 (  114 155 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.05 //y=7.4 //x2=8.88 //y2=7.4
r216 (  113 157 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.585 //y=7.4 //x2=9.67 //y2=7.4
r217 (  113 114 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=9.585 //y=7.4 //x2=9.05 //y2=7.4
r218 (  110 154 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.185 //y=7.4 //x2=8.1 //y2=7.4
r219 (  109 155 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.71 //y=7.4 //x2=8.88 //y2=7.4
r220 (  109 110 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=8.71 //y=7.4 //x2=8.185 //y2=7.4
r221 (  103 154 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.1 //y=7.23 //x2=8.1 //y2=7.4
r222 (  103 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.1 //y=7.23 //x2=8.1 //y2=6.745
r223 (  102 152 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.305 //y=7.4 //x2=7.22 //y2=7.4
r224 (  101 154 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.015 //y=7.4 //x2=8.1 //y2=7.4
r225 (  101 102 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.015 //y=7.4 //x2=7.305 //y2=7.4
r226 (  95 152 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.22 //y=7.23 //x2=7.22 //y2=7.4
r227 (  95 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.22 //y=7.23 //x2=7.22 //y2=6.745
r228 (  92 151 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.425 //y=7.4 //x2=6.34 //y2=7.4
r229 (  92 94 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=6.425 //y=7.4 //x2=7.03 //y2=7.4
r230 (  91 152 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.135 //y=7.4 //x2=7.22 //y2=7.4
r231 (  91 94 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=7.135 //y=7.4 //x2=7.03 //y2=7.4
r232 (  85 151 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.34 //y=7.23 //x2=6.34 //y2=7.4
r233 (  85 166 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=6.34 //y=7.23 //x2=6.34 //y2=6.405
r234 (  82 150 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.55 //y2=7.4
r235 (  82 84 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.92 //y2=7.4
r236 (  81 151 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.255 //y=7.4 //x2=6.34 //y2=7.4
r237 (  81 84 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=6.255 //y=7.4 //x2=5.92 //y2=7.4
r238 (  78 149 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.855 //y=7.4 //x2=4.77 //y2=7.4
r239 (  77 150 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=5.55 //y2=7.4
r240 (  77 78 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=4.855 //y2=7.4
r241 (  71 149 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.77 //y=7.23 //x2=4.77 //y2=7.4
r242 (  71 165 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.77 //y=7.23 //x2=4.77 //y2=6.745
r243 (  68 148 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.975 //y=7.4 //x2=3.89 //y2=7.4
r244 (  68 70 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=3.975 //y=7.4 //x2=4.44 //y2=7.4
r245 (  67 149 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.685 //y=7.4 //x2=4.77 //y2=7.4
r246 (  67 70 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=4.685 //y=7.4 //x2=4.44 //y2=7.4
r247 (  61 148 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.89 //y=7.23 //x2=3.89 //y2=7.4
r248 (  61 164 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.89 //y=7.23 //x2=3.89 //y2=6.745
r249 (  58 147 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.095 //y=7.4 //x2=3.01 //y2=7.4
r250 (  58 60 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=3.095 //y=7.4 //x2=3.33 //y2=7.4
r251 (  57 148 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.805 //y=7.4 //x2=3.89 //y2=7.4
r252 (  57 60 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=3.805 //y=7.4 //x2=3.33 //y2=7.4
r253 (  51 147 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.01 //y=7.23 //x2=3.01 //y2=7.4
r254 (  51 163 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=3.01 //y=7.23 //x2=3.01 //y2=6.405
r255 (  50 146 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.39 //y=7.4 //x2=2.22 //y2=7.4
r256 (  49 147 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.925 //y=7.4 //x2=3.01 //y2=7.4
r257 (  49 50 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=2.925 //y=7.4 //x2=2.39 //y2=7.4
r258 (  44 145 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.555 //y2=7.4
r259 (  44 46 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.85 //y2=7.4
r260 (  43 146 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.05 //y=7.4 //x2=2.22 //y2=7.4
r261 (  43 46 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=7.4 //x2=1.85 //y2=7.4
r262 (  37 145 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=7.4
r263 (  37 162 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=6.405
r264 (  36 144 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.76 //y=7.4 //x2=0.675 //y2=7.4
r265 (  35 145 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=1.555 //y2=7.4
r266 (  35 36 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=0.76 //y2=7.4
r267 (  29 144 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=7.4
r268 (  29 161 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=6.405
r269 (  23 160 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r270 (  21 132 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=7.4 //x2=10.73 //y2=7.4
r271 (  21 23 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=7.4 //x2=11.47 //y2=7.4
r272 (  19 157 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=7.4 //x2=9.62 //y2=7.4
r273 (  19 21 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.62 //y=7.4 //x2=10.73 //y2=7.4
r274 (  17 154 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=7.4 //x2=8.14 //y2=7.4
r275 (  17 19 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=7.4 //x2=9.62 //y2=7.4
r276 (  15 94 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=7.4 //x2=7.03 //y2=7.4
r277 (  15 17 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=7.4 //x2=8.14 //y2=7.4
r278 (  12 84 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=7.4 //x2=5.92 //y2=7.4
r279 (  10 70 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r280 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.92 //y2=7.4
r281 (  8 60 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=7.4 //x2=3.33 //y2=7.4
r282 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=7.4 //x2=4.44 //y2=7.4
r283 (  6 46 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r284 (  6 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=3.33 //y2=7.4
r285 (  3 144 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r286 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r287 (  1 15 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=6.105 //y=7.4 //x2=7.03 //y2=7.4
r288 (  1 12 ) resistor r=0.0768272 //w=0.301 //l=0.185 //layer=m1 \
 //thickness=0.36 //x=6.105 //y=7.4 //x2=5.92 //y2=7.4
ends PM_MUX2X1\%VDD

subckt PM_MUX2X1\%S ( 1 2 7 8 9 10 11 12 13 14 15 16 17 18 19 21 35 47 48 49 \
 50 51 52 53 54 55 56 60 61 62 64 70 71 72 73 74 75 79 81 84 85 90 104 )
c127 ( 104 0 ) capacitor c=0.0667949f //x=3.33 //y=4.7
c128 ( 90 0 ) capacitor c=0.051138f //x=0.74 //y=2.085
c129 ( 85 0 ) capacitor c=0.0318948f //x=3.665 //y=1.21
c130 ( 84 0 ) capacitor c=0.0187384f //x=3.665 //y=0.865
c131 ( 81 0 ) capacitor c=0.0141798f //x=3.51 //y=1.365
c132 ( 79 0 ) capacitor c=0.0149844f //x=3.51 //y=0.71
c133 ( 75 0 ) capacitor c=0.0819722f //x=3.135 //y=1.915
c134 ( 74 0 ) capacitor c=0.0229722f //x=3.135 //y=1.52
c135 ( 73 0 ) capacitor c=0.0234352f //x=3.135 //y=1.21
c136 ( 72 0 ) capacitor c=0.0199343f //x=3.135 //y=0.865
c137 ( 71 0 ) capacitor c=0.0435629f //x=1.38 //y=1.255
c138 ( 70 0 ) capacitor c=0.0200386f //x=1.38 //y=0.91
c139 ( 64 0 ) capacitor c=0.0152946f //x=1.225 //y=1.41
c140 ( 62 0 ) capacitor c=0.0157804f //x=1.225 //y=0.755
c141 ( 61 0 ) capacitor c=0.0524167f //x=0.97 //y=4.79
c142 ( 60 0 ) capacitor c=0.0322983f //x=1.26 //y=4.79
c143 ( 56 0 ) capacitor c=0.0290017f //x=0.85 //y=1.92
c144 ( 55 0 ) capacitor c=0.0250027f //x=0.85 //y=1.565
c145 ( 54 0 ) capacitor c=0.0234316f //x=0.85 //y=1.255
c146 ( 53 0 ) capacitor c=0.0200596f //x=0.85 //y=0.91
c147 ( 52 0 ) capacitor c=0.110275f //x=3.67 //y=6.02
c148 ( 51 0 ) capacitor c=0.154305f //x=3.23 //y=6.02
c149 ( 50 0 ) capacitor c=0.154218f //x=1.335 //y=6.02
c150 ( 49 0 ) capacitor c=0.154243f //x=0.895 //y=6.02
c151 ( 35 0 ) capacitor c=0.0971096f //x=3.33 //y=2.08
c152 ( 21 0 ) capacitor c=0.110891f //x=0.74 //y=2.085
c153 ( 2 0 ) capacitor c=0.0133976f //x=0.855 //y=2.96
c154 ( 1 0 ) capacitor c=0.0813108f //x=3.215 //y=2.96
r155 (  102 104 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=3.23 //y=4.7 //x2=3.33 //y2=4.7
r156 (  90 91 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=0.74 //y=2.085 //x2=0.85 //y2=2.085
r157 (  86 104 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=3.67 //y=4.865 //x2=3.33 //y2=4.7
r158 (  85 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.665 //y=1.21 //x2=3.625 //y2=1.365
r159 (  84 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.665 //y=0.865 //x2=3.625 //y2=0.71
r160 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.665 //y=0.865 //x2=3.665 //y2=1.21
r161 (  82 101 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.29 //y=1.365 //x2=3.175 //y2=1.365
r162 (  81 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.51 //y=1.365 //x2=3.625 //y2=1.365
r163 (  80 100 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.29 //y=0.71 //x2=3.175 //y2=0.71
r164 (  79 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.51 //y=0.71 //x2=3.625 //y2=0.71
r165 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.51 //y=0.71 //x2=3.29 //y2=0.71
r166 (  76 102 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.23 //y=4.865 //x2=3.23 //y2=4.7
r167 (  75 99 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.915 //x2=3.33 //y2=2.08
r168 (  74 101 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.52 //x2=3.175 //y2=1.365
r169 (  74 75 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.52 //x2=3.135 //y2=1.915
r170 (  73 101 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.21 //x2=3.175 //y2=1.365
r171 (  72 100 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=0.865 //x2=3.175 //y2=0.71
r172 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.135 //y=0.865 //x2=3.135 //y2=1.21
r173 (  71 97 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=1.255 //x2=1.34 //y2=1.41
r174 (  70 96 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.34 //y2=0.755
r175 (  70 71 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.38 //y2=1.255
r176 (  65 95 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=1.41 //x2=0.89 //y2=1.41
r177 (  64 97 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=1.41 //x2=1.34 //y2=1.41
r178 (  63 94 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=0.755 //x2=0.89 //y2=0.755
r179 (  62 96 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.34 //y2=0.755
r180 (  62 63 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.005 //y2=0.755
r181 (  60 67 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=1.335 //y2=4.865
r182 (  60 61 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=0.97 //y2=4.79
r183 (  57 61 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.97 //y2=4.79
r184 (  57 93 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.74 //y2=4.7
r185 (  56 91 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.92 //x2=0.85 //y2=2.085
r186 (  55 95 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.89 //y2=1.41
r187 (  55 56 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.85 //y2=1.92
r188 (  54 95 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.255 //x2=0.89 //y2=1.41
r189 (  53 94 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.89 //y2=0.755
r190 (  53 54 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.85 //y2=1.255
r191 (  52 86 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.67 //y=6.02 //x2=3.67 //y2=4.865
r192 (  51 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.23 //y=6.02 //x2=3.23 //y2=4.865
r193 (  50 67 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.335 //y=6.02 //x2=1.335 //y2=4.865
r194 (  49 57 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.895 //y=6.02 //x2=0.895 //y2=4.865
r195 (  48 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.4 //y=1.365 //x2=3.51 //y2=1.365
r196 (  48 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.4 //y=1.365 //x2=3.29 //y2=1.365
r197 (  47 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.225 //y2=1.41
r198 (  47 65 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.005 //y2=1.41
r199 (  45 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r200 (  35 99 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r201 (  32 93 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.7 //x2=0.74 //y2=4.7
r202 (  21 90 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=2.085
r203 (  19 45 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=3.33 //y=4.44 //x2=3.33 //y2=4.7
r204 (  18 19 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=4.07 //x2=3.33 //y2=4.44
r205 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.7 //x2=3.33 //y2=4.07
r206 (  16 17 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.96 //x2=3.33 //y2=3.7
r207 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.59 //x2=3.33 //y2=2.96
r208 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.22 //x2=3.33 //y2=2.59
r209 (  14 35 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.22 //x2=3.33 //y2=2.08
r210 (  13 32 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=0.74 //y=4.44 //x2=0.74 //y2=4.7
r211 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=4.07 //x2=0.74 //y2=4.44
r212 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=3.7 //x2=0.74 //y2=4.07
r213 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=3.33 //x2=0.74 //y2=3.7
r214 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=2.96 //x2=0.74 //y2=3.33
r215 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.59 //x2=0.74 //y2=2.96
r216 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.22 //x2=0.74 //y2=2.59
r217 (  7 21 ) resistor r=9.24064 //w=0.187 //l=0.135 //layer=li \
 //thickness=0.1 //x=0.74 //y=2.22 //x2=0.74 //y2=2.085
r218 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=2.96 //x2=3.33 //y2=2.96
r219 (  4 9 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=0.74 \
 //y=2.96 //x2=0.74 //y2=2.96
r220 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=0.855 //y=2.96 //x2=0.74 //y2=2.96
r221 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.215 //y=2.96 //x2=3.33 //y2=2.96
r222 (  1 2 ) resistor r=2.25191 //w=0.131 //l=2.36 //layer=m1 \
 //thickness=0.36 //x=3.215 //y=2.96 //x2=0.855 //y2=2.96
ends PM_MUX2X1\%S

subckt PM_MUX2X1\%noxref_4 ( 1 2 17 18 19 20 24 26 33 34 35 36 37 38 39 43 45 \
 48 49 59 62 64 )
c139 ( 64 0 ) capacitor c=0.0288745f //x=0.97 //y=5.02
c140 ( 62 0 ) capacitor c=0.0173218f //x=0.925 //y=0.91
c141 ( 59 0 ) capacitor c=0.0667949f //x=6.66 //y=4.7
c142 ( 49 0 ) capacitor c=0.0318948f //x=6.995 //y=1.21
c143 ( 48 0 ) capacitor c=0.0187384f //x=6.995 //y=0.865
c144 ( 45 0 ) capacitor c=0.0141798f //x=6.84 //y=1.365
c145 ( 43 0 ) capacitor c=0.0149844f //x=6.84 //y=0.71
c146 ( 39 0 ) capacitor c=0.0819799f //x=6.465 //y=1.915
c147 ( 38 0 ) capacitor c=0.0229722f //x=6.465 //y=1.52
c148 ( 37 0 ) capacitor c=0.0234352f //x=6.465 //y=1.21
c149 ( 36 0 ) capacitor c=0.0199343f //x=6.465 //y=0.865
c150 ( 35 0 ) capacitor c=0.110275f //x=7 //y=6.02
c151 ( 34 0 ) capacitor c=0.154305f //x=6.56 //y=6.02
c152 ( 26 0 ) capacitor c=0.0969029f //x=6.66 //y=2.08
c153 ( 24 0 ) capacitor c=0.0857489f //x=1.48 //y=3.33
c154 ( 20 0 ) capacitor c=0.00560375f //x=1.2 //y=4.58
c155 ( 19 0 ) capacitor c=0.0134399f //x=1.395 //y=4.58
c156 ( 18 0 ) capacitor c=0.00549299f //x=1.195 //y=2.08
c157 ( 17 0 ) capacitor c=0.013178f //x=1.395 //y=2.08
c158 ( 2 0 ) capacitor c=0.0158256f //x=1.595 //y=3.33
c159 ( 1 0 ) capacitor c=0.183474f //x=6.545 //y=3.33
r160 (  57 59 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=6.56 //y=4.7 //x2=6.66 //y2=4.7
r161 (  50 59 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=7 //y=4.865 //x2=6.66 //y2=4.7
r162 (  49 61 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.995 //y=1.21 //x2=6.955 //y2=1.365
r163 (  48 60 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.995 //y=0.865 //x2=6.955 //y2=0.71
r164 (  48 49 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.995 //y=0.865 //x2=6.995 //y2=1.21
r165 (  46 56 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.62 //y=1.365 //x2=6.505 //y2=1.365
r166 (  45 61 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.84 //y=1.365 //x2=6.955 //y2=1.365
r167 (  44 55 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.62 //y=0.71 //x2=6.505 //y2=0.71
r168 (  43 60 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.84 //y=0.71 //x2=6.955 //y2=0.71
r169 (  43 44 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.84 //y=0.71 //x2=6.62 //y2=0.71
r170 (  40 57 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.56 //y=4.865 //x2=6.56 //y2=4.7
r171 (  39 54 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.915 //x2=6.66 //y2=2.08
r172 (  38 56 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.52 //x2=6.505 //y2=1.365
r173 (  38 39 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.52 //x2=6.465 //y2=1.915
r174 (  37 56 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.21 //x2=6.505 //y2=1.365
r175 (  36 55 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.465 //y=0.865 //x2=6.505 //y2=0.71
r176 (  36 37 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.465 //y=0.865 //x2=6.465 //y2=1.21
r177 (  35 50 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7 //y=6.02 //x2=7 //y2=4.865
r178 (  34 40 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.56 //y=6.02 //x2=6.56 //y2=4.865
r179 (  33 45 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.73 //y=1.365 //x2=6.84 //y2=1.365
r180 (  33 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.73 //y=1.365 //x2=6.62 //y2=1.365
r181 (  31 59 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=4.7 //x2=6.66 //y2=4.7
r182 (  29 31 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=6.66 //y=3.33 //x2=6.66 //y2=4.7
r183 (  26 54 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.08 //x2=6.66 //y2=2.08
r184 (  26 29 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.08 //x2=6.66 //y2=3.33
r185 (  22 24 ) resistor r=79.7433 //w=0.187 //l=1.165 //layer=li \
 //thickness=0.1 //x=1.48 //y=4.495 //x2=1.48 //y2=3.33
r186 (  21 24 ) resistor r=79.7433 //w=0.187 //l=1.165 //layer=li \
 //thickness=0.1 //x=1.48 //y=2.165 //x2=1.48 //y2=3.33
r187 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.48 //y2=4.495
r188 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.2 //y2=4.58
r189 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.48 //y2=2.165
r190 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.195 //y2=2.08
r191 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.2 //y2=4.58
r192 (  11 64 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.115 //y2=5.725
r193 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.195 //y2=2.08
r194 (  7 62 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.11 //y2=1.005
r195 (  6 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=3.33 //x2=6.66 //y2=3.33
r196 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.48 //y=3.33 //x2=1.48 //y2=3.33
r197 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.595 //y=3.33 //x2=1.48 //y2=3.33
r198 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.545 //y=3.33 //x2=6.66 //y2=3.33
r199 (  1 2 ) resistor r=4.72328 //w=0.131 //l=4.95 //layer=m1 \
 //thickness=0.36 //x=6.545 //y=3.33 //x2=1.595 //y2=3.33
ends PM_MUX2X1\%noxref_4

subckt PM_MUX2X1\%noxref_5 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 \
 52 54 57 58 68 71 73 74 )
c168 ( 74 0 ) capacitor c=0.0220291f //x=4.185 //y=5.02
c169 ( 73 0 ) capacitor c=0.0217503f //x=3.305 //y=5.02
c170 ( 71 0 ) capacitor c=0.00866655f //x=4.18 //y=0.905
c171 ( 68 0 ) capacitor c=0.0667949f //x=9.99 //y=4.7
c172 ( 58 0 ) capacitor c=0.0318948f //x=10.325 //y=1.21
c173 ( 57 0 ) capacitor c=0.0187384f //x=10.325 //y=0.865
c174 ( 54 0 ) capacitor c=0.0141798f //x=10.17 //y=1.365
c175 ( 52 0 ) capacitor c=0.0149844f //x=10.17 //y=0.71
c176 ( 48 0 ) capacitor c=0.0819722f //x=9.795 //y=1.915
c177 ( 47 0 ) capacitor c=0.0229722f //x=9.795 //y=1.52
c178 ( 46 0 ) capacitor c=0.0234352f //x=9.795 //y=1.21
c179 ( 45 0 ) capacitor c=0.0199343f //x=9.795 //y=0.865
c180 ( 44 0 ) capacitor c=0.110275f //x=10.33 //y=6.02
c181 ( 43 0 ) capacitor c=0.154305f //x=9.89 //y=6.02
c182 ( 41 0 ) capacitor c=0.00264586f //x=4.33 //y=5.2
c183 ( 34 0 ) capacitor c=0.09625f //x=9.99 //y=2.08
c184 ( 32 0 ) capacitor c=0.113528f //x=4.81 //y=2.96
c185 ( 28 0 ) capacitor c=0.00498573f //x=4.455 //y=1.655
c186 ( 27 0 ) capacitor c=0.0135368f //x=4.725 //y=1.655
c187 ( 25 0 ) capacitor c=0.0145797f //x=4.725 //y=5.2
c188 ( 14 0 ) capacitor c=0.00290084f //x=3.535 //y=5.2
c189 ( 13 0 ) capacitor c=0.0161139f //x=4.245 //y=5.2
c190 ( 2 0 ) capacitor c=0.00976349f //x=4.925 //y=2.96
c191 ( 1 0 ) capacitor c=0.168301f //x=9.875 //y=2.96
r192 (  66 68 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=9.89 //y=4.7 //x2=9.99 //y2=4.7
r193 (  59 68 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=10.33 //y=4.865 //x2=9.99 //y2=4.7
r194 (  58 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.325 //y=1.21 //x2=10.285 //y2=1.365
r195 (  57 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.325 //y=0.865 //x2=10.285 //y2=0.71
r196 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.325 //y=0.865 //x2=10.325 //y2=1.21
r197 (  55 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.95 //y=1.365 //x2=9.835 //y2=1.365
r198 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.17 //y=1.365 //x2=10.285 //y2=1.365
r199 (  53 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.95 //y=0.71 //x2=9.835 //y2=0.71
r200 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.17 //y=0.71 //x2=10.285 //y2=0.71
r201 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.17 //y=0.71 //x2=9.95 //y2=0.71
r202 (  49 66 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=9.89 //y=4.865 //x2=9.89 //y2=4.7
r203 (  48 63 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=9.795 //y=1.915 //x2=9.99 //y2=2.08
r204 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.795 //y=1.52 //x2=9.835 //y2=1.365
r205 (  47 48 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=9.795 //y=1.52 //x2=9.795 //y2=1.915
r206 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.795 //y=1.21 //x2=9.835 //y2=1.365
r207 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.795 //y=0.865 //x2=9.835 //y2=0.71
r208 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.795 //y=0.865 //x2=9.795 //y2=1.21
r209 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.33 //y=6.02 //x2=10.33 //y2=4.865
r210 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.89 //y=6.02 //x2=9.89 //y2=4.865
r211 (  42 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.06 //y=1.365 //x2=10.17 //y2=1.365
r212 (  42 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.06 //y=1.365 //x2=9.95 //y2=1.365
r213 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.99 //y=4.7 //x2=9.99 //y2=4.7
r214 (  37 39 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=9.99 //y=2.96 //x2=9.99 //y2=4.7
r215 (  34 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.99 //y=2.08 //x2=9.99 //y2=2.08
r216 (  34 37 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=9.99 //y=2.08 //x2=9.99 //y2=2.96
r217 (  30 32 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=4.81 //y=5.115 //x2=4.81 //y2=2.96
r218 (  29 32 ) resistor r=83.508 //w=0.187 //l=1.22 //layer=li \
 //thickness=0.1 //x=4.81 //y=1.74 //x2=4.81 //y2=2.96
r219 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=1.655 //x2=4.81 //y2=1.74
r220 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=4.725 //y=1.655 //x2=4.455 //y2=1.655
r221 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.415 //y=5.2 //x2=4.33 //y2=5.2
r222 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=5.2 //x2=4.81 //y2=5.115
r223 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=4.725 //y=5.2 //x2=4.415 //y2=5.2
r224 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.37 //y=1.57 //x2=4.455 //y2=1.655
r225 (  21 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.37 //y=1.57 //x2=4.37 //y2=1
r226 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.33 //y=5.285 //x2=4.33 //y2=5.2
r227 (  15 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=4.33 //y=5.285 //x2=4.33 //y2=5.725
r228 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.245 //y=5.2 //x2=4.33 //y2=5.2
r229 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=4.245 //y=5.2 //x2=3.535 //y2=5.2
r230 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.45 //y=5.285 //x2=3.535 //y2=5.2
r231 (  7 73 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=3.45 //y=5.285 //x2=3.45 //y2=5.725
r232 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.99 //y=2.96 //x2=9.99 //y2=2.96
r233 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.81 //y=2.96 //x2=4.81 //y2=2.96
r234 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.925 //y=2.96 //x2=4.81 //y2=2.96
r235 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.875 //y=2.96 //x2=9.99 //y2=2.96
r236 (  1 2 ) resistor r=4.72328 //w=0.131 //l=4.95 //layer=m1 \
 //thickness=0.36 //x=9.875 //y=2.96 //x2=4.925 //y2=2.96
ends PM_MUX2X1\%noxref_5

subckt PM_MUX2X1\%noxref_6 ( 1 2 13 14 25 27 28 32 33 35 39 42 43 44 45 46 47 \
 52 54 56 62 63 65 66 69 77 79 80 )
c155 ( 80 0 ) capacitor c=0.0220291f //x=7.515 //y=5.02
c156 ( 79 0 ) capacitor c=0.0217503f //x=6.635 //y=5.02
c157 ( 77 0 ) capacitor c=0.00866655f //x=7.51 //y=0.905
c158 ( 69 0 ) capacitor c=0.034715f //x=10.76 //y=4.7
c159 ( 66 0 ) capacitor c=0.0279499f //x=10.73 //y=1.915
c160 ( 65 0 ) capacitor c=0.0428694f //x=10.73 //y=2.08
c161 ( 63 0 ) capacitor c=0.0429696f //x=11.295 //y=1.25
c162 ( 62 0 ) capacitor c=0.0192208f //x=11.295 //y=0.905
c163 ( 56 0 ) capacitor c=0.0158629f //x=11.14 //y=1.405
c164 ( 54 0 ) capacitor c=0.0157803f //x=11.14 //y=0.75
c165 ( 52 0 ) capacitor c=0.0366192f //x=11.135 //y=4.79
c166 ( 47 0 ) capacitor c=0.0205163f //x=10.765 //y=1.56
c167 ( 46 0 ) capacitor c=0.0168481f //x=10.765 //y=1.25
c168 ( 45 0 ) capacitor c=0.0174783f //x=10.765 //y=0.905
c169 ( 44 0 ) capacitor c=0.15358f //x=11.21 //y=6.02
c170 ( 43 0 ) capacitor c=0.110281f //x=10.77 //y=6.02
c171 ( 39 0 ) capacitor c=0.00279371f //x=7.66 //y=5.2
c172 ( 35 0 ) capacitor c=0.0787765f //x=10.73 //y=2.08
c173 ( 33 0 ) capacitor c=0.00453889f //x=10.73 //y=4.535
c174 ( 32 0 ) capacitor c=0.113733f //x=8.14 //y=3.33
c175 ( 28 0 ) capacitor c=0.00468667f //x=7.785 //y=1.655
c176 ( 27 0 ) capacitor c=0.0131863f //x=8.055 //y=1.655
c177 ( 25 0 ) capacitor c=0.0147208f //x=8.055 //y=5.2
c178 ( 14 0 ) capacitor c=0.0029559f //x=6.865 //y=5.2
c179 ( 13 0 ) capacitor c=0.0166338f //x=7.575 //y=5.2
c180 ( 2 0 ) capacitor c=0.00897649f //x=8.255 //y=3.33
c181 ( 1 0 ) capacitor c=0.100712f //x=10.615 //y=3.33
r182 (  71 72 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=10.76 //y=4.79 //x2=10.76 //y2=4.865
r183 (  69 71 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=10.76 //y=4.7 //x2=10.76 //y2=4.79
r184 (  65 66 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=10.73 //y=2.08 //x2=10.73 //y2=1.915
r185 (  63 76 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.295 //y=1.25 //x2=11.255 //y2=1.405
r186 (  62 75 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.295 //y=0.905 //x2=11.255 //y2=0.75
r187 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.295 //y=0.905 //x2=11.295 //y2=1.25
r188 (  57 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.92 //y=1.405 //x2=10.805 //y2=1.405
r189 (  56 76 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.14 //y=1.405 //x2=11.255 //y2=1.405
r190 (  55 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.92 //y=0.75 //x2=10.805 //y2=0.75
r191 (  54 75 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.14 //y=0.75 //x2=11.255 //y2=0.75
r192 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=11.14 //y=0.75 //x2=10.92 //y2=0.75
r193 (  53 71 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=10.895 //y=4.79 //x2=10.76 //y2=4.79
r194 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.135 //y=4.79 //x2=11.21 //y2=4.865
r195 (  52 53 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=11.135 //y=4.79 //x2=10.895 //y2=4.79
r196 (  47 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.765 //y=1.56 //x2=10.805 //y2=1.405
r197 (  47 66 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=10.765 //y=1.56 //x2=10.765 //y2=1.915
r198 (  46 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.765 //y=1.25 //x2=10.805 //y2=1.405
r199 (  45 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.765 //y=0.905 //x2=10.805 //y2=0.75
r200 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.765 //y=0.905 //x2=10.765 //y2=1.25
r201 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.21 //y=6.02 //x2=11.21 //y2=4.865
r202 (  43 72 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.77 //y=6.02 //x2=10.77 //y2=4.865
r203 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.03 //y=1.405 //x2=11.14 //y2=1.405
r204 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.03 //y=1.405 //x2=10.92 //y2=1.405
r205 (  41 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.76 //y=4.7 //x2=10.76 //y2=4.7
r206 (  35 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=2.08 //x2=10.73 //y2=2.08
r207 (  35 38 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.08 //x2=10.73 //y2=3.33
r208 (  33 41 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=10.73 //y=4.535 //x2=10.745 //y2=4.7
r209 (  33 38 ) resistor r=82.4813 //w=0.187 //l=1.205 //layer=li \
 //thickness=0.1 //x=10.73 //y=4.535 //x2=10.73 //y2=3.33
r210 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=8.14 //y=5.115 //x2=8.14 //y2=3.33
r211 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=8.14 //y=1.74 //x2=8.14 //y2=3.33
r212 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.055 //y=1.655 //x2=8.14 //y2=1.74
r213 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=8.055 //y=1.655 //x2=7.785 //y2=1.655
r214 (  26 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.745 //y=5.2 //x2=7.66 //y2=5.2
r215 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.055 //y=5.2 //x2=8.14 //y2=5.115
r216 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=8.055 //y=5.2 //x2=7.745 //y2=5.2
r217 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.7 //y=1.57 //x2=7.785 //y2=1.655
r218 (  21 77 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=7.7 //y=1.57 //x2=7.7 //y2=1
r219 (  15 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.66 //y=5.285 //x2=7.66 //y2=5.2
r220 (  15 80 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=7.66 //y=5.285 //x2=7.66 //y2=5.725
r221 (  13 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.575 //y=5.2 //x2=7.66 //y2=5.2
r222 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.575 //y=5.2 //x2=6.865 //y2=5.2
r223 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.78 //y=5.285 //x2=6.865 //y2=5.2
r224 (  7 79 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.78 //y=5.285 //x2=6.78 //y2=5.725
r225 (  6 38 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=3.33 //x2=10.73 //y2=3.33
r226 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.14 //y=3.33 //x2=8.14 //y2=3.33
r227 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.255 //y=3.33 //x2=8.14 //y2=3.33
r228 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=3.33 //x2=10.73 //y2=3.33
r229 (  1 2 ) resistor r=2.25191 //w=0.131 //l=2.36 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=3.33 //x2=8.255 //y2=3.33
ends PM_MUX2X1\%noxref_6

subckt PM_MUX2X1\%A0 ( 1 2 3 4 5 6 7 9 19 20 21 22 23 24 29 31 33 39 40 42 43 \
 46 )
c68 ( 46 0 ) capacitor c=0.034715f //x=4.1 //y=4.7
c69 ( 43 0 ) capacitor c=0.0279499f //x=4.07 //y=1.915
c70 ( 42 0 ) capacitor c=0.0437302f //x=4.07 //y=2.08
c71 ( 40 0 ) capacitor c=0.0429696f //x=4.635 //y=1.25
c72 ( 39 0 ) capacitor c=0.0192208f //x=4.635 //y=0.905
c73 ( 33 0 ) capacitor c=0.0158629f //x=4.48 //y=1.405
c74 ( 31 0 ) capacitor c=0.0157803f //x=4.48 //y=0.75
c75 ( 29 0 ) capacitor c=0.0366192f //x=4.475 //y=4.79
c76 ( 24 0 ) capacitor c=0.0205163f //x=4.105 //y=1.56
c77 ( 23 0 ) capacitor c=0.0168481f //x=4.105 //y=1.25
c78 ( 22 0 ) capacitor c=0.0174783f //x=4.105 //y=0.905
c79 ( 21 0 ) capacitor c=0.15358f //x=4.55 //y=6.02
c80 ( 20 0 ) capacitor c=0.110281f //x=4.11 //y=6.02
c81 ( 9 0 ) capacitor c=0.0784233f //x=4.07 //y=2.08
c82 ( 7 0 ) capacitor c=0.00453889f //x=4.07 //y=4.535
r83 (  48 49 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=4.1 //y=4.79 //x2=4.1 //y2=4.865
r84 (  46 48 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=4.1 //y=4.7 //x2=4.1 //y2=4.79
r85 (  42 43 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=4.07 //y=2.08 //x2=4.07 //y2=1.915
r86 (  40 53 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.635 //y=1.25 //x2=4.595 //y2=1.405
r87 (  39 52 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.635 //y=0.905 //x2=4.595 //y2=0.75
r88 (  39 40 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.635 //y=0.905 //x2=4.635 //y2=1.25
r89 (  34 51 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.26 //y=1.405 //x2=4.145 //y2=1.405
r90 (  33 53 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.48 //y=1.405 //x2=4.595 //y2=1.405
r91 (  32 50 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.26 //y=0.75 //x2=4.145 //y2=0.75
r92 (  31 52 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.48 //y=0.75 //x2=4.595 //y2=0.75
r93 (  31 32 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.48 //y=0.75 //x2=4.26 //y2=0.75
r94 (  30 48 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=4.235 //y=4.79 //x2=4.1 //y2=4.79
r95 (  29 36 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.475 //y=4.79 //x2=4.55 //y2=4.865
r96 (  29 30 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=4.475 //y=4.79 //x2=4.235 //y2=4.79
r97 (  24 51 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.56 //x2=4.145 //y2=1.405
r98 (  24 43 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.56 //x2=4.105 //y2=1.915
r99 (  23 51 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.25 //x2=4.145 //y2=1.405
r100 (  22 50 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=0.905 //x2=4.145 //y2=0.75
r101 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.105 //y=0.905 //x2=4.105 //y2=1.25
r102 (  21 36 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.55 //y=6.02 //x2=4.55 //y2=4.865
r103 (  20 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.11 //y=6.02 //x2=4.11 //y2=4.865
r104 (  19 33 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.37 //y=1.405 //x2=4.48 //y2=1.405
r105 (  19 34 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.37 //y=1.405 //x2=4.26 //y2=1.405
r106 (  18 46 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.1 //y=4.7 //x2=4.1 //y2=4.7
r107 (  9 42 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=2.08 //x2=4.07 //y2=2.08
r108 (  7 18 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=4.07 //y=4.535 //x2=4.085 //y2=4.7
r109 (  6 7 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=4.07 //y=4.44 //x2=4.07 //y2=4.535
r110 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.07 //y=4.07 //x2=4.07 //y2=4.44
r111 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.07 //y=3.7 //x2=4.07 //y2=4.07
r112 (  3 4 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li //thickness=0.1 \
 //x=4.07 //y=2.96 //x2=4.07 //y2=3.7
r113 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.07 //y=2.59 //x2=4.07 //y2=2.96
r114 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.07 //y=2.22 //x2=4.07 //y2=2.59
r115 (  1 9 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li //thickness=0.1 \
 //x=4.07 //y=2.22 //x2=4.07 //y2=2.08
ends PM_MUX2X1\%A0

subckt PM_MUX2X1\%noxref_8 ( 1 5 9 10 13 17 29 )
c57 ( 29 0 ) capacitor c=0.0632369f //x=2.78 //y=0.365
c58 ( 17 0 ) capacitor c=0.00722223f //x=4.855 //y=0.615
c59 ( 13 0 ) capacitor c=0.0148778f //x=4.77 //y=0.53
c60 ( 10 0 ) capacitor c=0.00664066f //x=3.885 //y=1.495
c61 ( 9 0 ) capacitor c=0.006761f //x=3.885 //y=0.615
c62 ( 5 0 ) capacitor c=0.0194491f //x=3.8 //y=1.58
c63 ( 1 0 ) capacitor c=0.00798521f //x=2.915 //y=1.495
r64 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.855 //y=0.615 //x2=4.855 //y2=0.49
r65 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.855 //y=0.615 //x2=4.855 //y2=0.88
r66 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.97 //y=0.53 //x2=3.885 //y2=0.49
r67 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.97 //y=0.53 //x2=4.37 //y2=0.53
r68 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.77 //y=0.53 //x2=4.855 //y2=0.49
r69 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.77 //y=0.53 //x2=4.37 //y2=0.53
r70 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=3.885 //y=1.495 //x2=3.885 //y2=1.62
r71 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=3.885 //y=1.495 //x2=3.885 //y2=0.88
r72 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.885 //y=0.615 //x2=3.885 //y2=0.49
r73 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.885 //y=0.615 //x2=3.885 //y2=0.88
r74 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3 //y=1.58 //x2=2.915 //y2=1.62
r75 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3 //y=1.58 //x2=3.4 //y2=1.58
r76 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.8 //y=1.58 //x2=3.885 //y2=1.62
r77 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.8 //y=1.58 //x2=3.4 //y2=1.58
r78 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=2.915 //y=1.495 //x2=2.915 //y2=1.62
r79 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.915 //y=1.495 //x2=2.915 //y2=0.88
ends PM_MUX2X1\%noxref_8

subckt PM_MUX2X1\%A1 ( 1 2 3 4 5 6 7 9 19 20 21 22 23 24 29 31 33 39 40 42 43 \
 46 )
c69 ( 46 0 ) capacitor c=0.034715f //x=7.43 //y=4.7
c70 ( 43 0 ) capacitor c=0.0279499f //x=7.4 //y=1.915
c71 ( 42 0 ) capacitor c=0.0422587f //x=7.4 //y=2.08
c72 ( 40 0 ) capacitor c=0.0429696f //x=7.965 //y=1.25
c73 ( 39 0 ) capacitor c=0.0192208f //x=7.965 //y=0.905
c74 ( 33 0 ) capacitor c=0.0158629f //x=7.81 //y=1.405
c75 ( 31 0 ) capacitor c=0.0157803f //x=7.81 //y=0.75
c76 ( 29 0 ) capacitor c=0.0366192f //x=7.805 //y=4.79
c77 ( 24 0 ) capacitor c=0.0205163f //x=7.435 //y=1.56
c78 ( 23 0 ) capacitor c=0.0168481f //x=7.435 //y=1.25
c79 ( 22 0 ) capacitor c=0.0174783f //x=7.435 //y=0.905
c80 ( 21 0 ) capacitor c=0.15358f //x=7.88 //y=6.02
c81 ( 20 0 ) capacitor c=0.110281f //x=7.44 //y=6.02
c82 ( 9 0 ) capacitor c=0.0784233f //x=7.4 //y=2.08
c83 ( 7 0 ) capacitor c=0.00453889f //x=7.4 //y=4.535
r84 (  48 49 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=7.43 //y=4.79 //x2=7.43 //y2=4.865
r85 (  46 48 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=7.43 //y=4.7 //x2=7.43 //y2=4.79
r86 (  42 43 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=7.4 //y=2.08 //x2=7.4 //y2=1.915
r87 (  40 53 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.965 //y=1.25 //x2=7.925 //y2=1.405
r88 (  39 52 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.965 //y=0.905 //x2=7.925 //y2=0.75
r89 (  39 40 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.965 //y=0.905 //x2=7.965 //y2=1.25
r90 (  34 51 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.59 //y=1.405 //x2=7.475 //y2=1.405
r91 (  33 53 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.81 //y=1.405 //x2=7.925 //y2=1.405
r92 (  32 50 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.59 //y=0.75 //x2=7.475 //y2=0.75
r93 (  31 52 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.81 //y=0.75 //x2=7.925 //y2=0.75
r94 (  31 32 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.81 //y=0.75 //x2=7.59 //y2=0.75
r95 (  30 48 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=7.565 //y=4.79 //x2=7.43 //y2=4.79
r96 (  29 36 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.805 //y=4.79 //x2=7.88 //y2=4.865
r97 (  29 30 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=7.805 //y=4.79 //x2=7.565 //y2=4.79
r98 (  24 51 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.56 //x2=7.475 //y2=1.405
r99 (  24 43 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.56 //x2=7.435 //y2=1.915
r100 (  23 51 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.25 //x2=7.475 //y2=1.405
r101 (  22 50 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.435 //y=0.905 //x2=7.475 //y2=0.75
r102 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.435 //y=0.905 //x2=7.435 //y2=1.25
r103 (  21 36 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.88 //y=6.02 //x2=7.88 //y2=4.865
r104 (  20 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.44 //y=6.02 //x2=7.44 //y2=4.865
r105 (  19 33 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.7 //y=1.405 //x2=7.81 //y2=1.405
r106 (  19 34 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.7 //y=1.405 //x2=7.59 //y2=1.405
r107 (  18 46 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.43 //y=4.7 //x2=7.43 //y2=4.7
r108 (  9 42 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.4 //y=2.08 //x2=7.4 //y2=2.08
r109 (  7 18 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=7.4 //y=4.535 //x2=7.415 //y2=4.7
r110 (  6 7 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=7.4 //y=4.44 //x2=7.4 //y2=4.535
r111 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=7.4 //y=4.07 //x2=7.4 //y2=4.44
r112 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=7.4 //y=3.7 //x2=7.4 //y2=4.07
r113 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=7.4 //y=3.33 //x2=7.4 //y2=3.7
r114 (  2 3 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li //thickness=0.1 \
 //x=7.4 //y=2.59 //x2=7.4 //y2=3.33
r115 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=7.4 //y=2.22 //x2=7.4 //y2=2.59
r116 (  1 9 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li //thickness=0.1 \
 //x=7.4 //y=2.22 //x2=7.4 //y2=2.08
ends PM_MUX2X1\%A1

subckt PM_MUX2X1\%noxref_10 ( 1 5 9 10 13 17 29 )
c55 ( 29 0 ) capacitor c=0.0635478f //x=6.11 //y=0.365
c56 ( 17 0 ) capacitor c=0.00722223f //x=8.185 //y=0.615
c57 ( 13 0 ) capacitor c=0.0147854f //x=8.1 //y=0.53
c58 ( 10 0 ) capacitor c=0.00638095f //x=7.215 //y=1.495
c59 ( 9 0 ) capacitor c=0.006761f //x=7.215 //y=0.615
c60 ( 5 0 ) capacitor c=0.0189075f //x=7.13 //y=1.58
c61 ( 1 0 ) capacitor c=0.00798521f //x=6.245 //y=1.495
r62 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.185 //y=0.615 //x2=8.185 //y2=0.49
r63 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=8.185 //y=0.615 //x2=8.185 //y2=0.88
r64 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.3 //y=0.53 //x2=7.215 //y2=0.49
r65 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.3 //y=0.53 //x2=7.7 //y2=0.53
r66 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.1 //y=0.53 //x2=8.185 //y2=0.49
r67 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.1 //y=0.53 //x2=7.7 //y2=0.53
r68 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.215 //y=1.495 //x2=7.215 //y2=1.62
r69 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=7.215 //y=1.495 //x2=7.215 //y2=0.88
r70 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.215 //y=0.615 //x2=7.215 //y2=0.49
r71 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=7.215 //y=0.615 //x2=7.215 //y2=0.88
r72 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.33 //y=1.58 //x2=6.245 //y2=1.62
r73 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.33 //y=1.58 //x2=6.73 //y2=1.58
r74 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.13 //y=1.58 //x2=7.215 //y2=1.62
r75 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.13 //y=1.58 //x2=6.73 //y2=1.58
r76 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.245 //y=1.495 //x2=6.245 //y2=1.62
r77 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.245 //y=1.495 //x2=6.245 //y2=0.88
ends PM_MUX2X1\%noxref_10

subckt PM_MUX2X1\%Y ( 1 2 3 4 5 6 7 8 15 16 27 29 30 41 42 44 45 )
c65 ( 45 0 ) capacitor c=0.0220291f //x=10.845 //y=5.02
c66 ( 44 0 ) capacitor c=0.0217503f //x=9.965 //y=5.02
c67 ( 42 0 ) capacitor c=0.0084702f //x=10.84 //y=0.905
c68 ( 41 0 ) capacitor c=0.00427536f //x=10.99 //y=5.2
c69 ( 30 0 ) capacitor c=0.00781917f //x=11.115 //y=1.655
c70 ( 29 0 ) capacitor c=0.0167625f //x=11.385 //y=1.655
c71 ( 27 0 ) capacitor c=0.0162757f //x=11.385 //y=5.2
c72 ( 16 0 ) capacitor c=0.00289676f //x=10.195 //y=5.2
c73 ( 15 0 ) capacitor c=0.0167385f //x=10.905 //y=5.2
c74 ( 1 0 ) capacitor c=0.132268f //x=11.47 //y=2.22
r75 (  29 31 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.385 //y=1.655 //x2=11.47 //y2=1.74
r76 (  29 30 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=11.385 //y=1.655 //x2=11.115 //y2=1.655
r77 (  28 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.075 //y=5.2 //x2=10.99 //y2=5.2
r78 (  27 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.385 //y=5.2 //x2=11.47 //y2=5.115
r79 (  27 28 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=11.385 //y=5.2 //x2=11.075 //y2=5.2
r80 (  23 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.03 //y=1.57 //x2=11.115 //y2=1.655
r81 (  23 42 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=11.03 //y=1.57 //x2=11.03 //y2=1
r82 (  17 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.99 //y=5.285 //x2=10.99 //y2=5.2
r83 (  17 45 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=10.99 //y=5.285 //x2=10.99 //y2=5.725
r84 (  15 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=10.905 //y=5.2 //x2=10.99 //y2=5.2
r85 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.905 //y=5.2 //x2=10.195 //y2=5.2
r86 (  9 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.11 //y=5.285 //x2=10.195 //y2=5.2
r87 (  9 44 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li //thickness=0.1 \
 //x=10.11 //y=5.285 //x2=10.11 //y2=5.725
r88 (  8 32 ) resistor r=20.877 //w=0.187 //l=0.305 //layer=li //thickness=0.1 \
 //x=11.47 //y=4.81 //x2=11.47 //y2=5.115
r89 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=11.47 //y=4.44 //x2=11.47 //y2=4.81
r90 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=11.47 //y=4.07 //x2=11.47 //y2=4.44
r91 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=11.47 //y=3.7 //x2=11.47 //y2=4.07
r92 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=11.47 //y=3.33 //x2=11.47 //y2=3.7
r93 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=11.47 //y=2.96 //x2=11.47 //y2=3.33
r94 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=11.47 //y=2.59 //x2=11.47 //y2=2.96
r95 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=11.47 //y=2.22 //x2=11.47 //y2=2.59
r96 (  1 31 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li //thickness=0.1 \
 //x=11.47 //y=2.22 //x2=11.47 //y2=1.74
ends PM_MUX2X1\%Y

subckt PM_MUX2X1\%noxref_12 ( 1 5 9 10 13 17 29 )
c49 ( 29 0 ) capacitor c=0.0644508f //x=9.44 //y=0.365
c50 ( 17 0 ) capacitor c=0.00722223f //x=11.515 //y=0.615
c51 ( 13 0 ) capacitor c=0.0152085f //x=11.43 //y=0.53
c52 ( 10 0 ) capacitor c=0.00664f //x=10.545 //y=1.495
c53 ( 9 0 ) capacitor c=0.006761f //x=10.545 //y=0.615
c54 ( 5 0 ) capacitor c=0.0194491f //x=10.46 //y=1.58
c55 ( 1 0 ) capacitor c=0.00798521f //x=9.575 //y=1.495
r56 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=11.515 //y=0.615 //x2=11.515 //y2=0.49
r57 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=11.515 //y=0.615 //x2=11.515 //y2=0.88
r58 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.63 //y=0.53 //x2=10.545 //y2=0.49
r59 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.63 //y=0.53 //x2=11.03 //y2=0.53
r60 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.43 //y=0.53 //x2=11.515 //y2=0.49
r61 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.43 //y=0.53 //x2=11.03 //y2=0.53
r62 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=10.545 //y=1.495 //x2=10.545 //y2=1.62
r63 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.545 //y=1.495 //x2=10.545 //y2=0.88
r64 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=10.545 //y=0.615 //x2=10.545 //y2=0.49
r65 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=10.545 //y=0.615 //x2=10.545 //y2=0.88
r66 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.66 //y=1.58 //x2=9.575 //y2=1.62
r67 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.66 //y=1.58 //x2=10.06 //y2=1.58
r68 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.46 //y=1.58 //x2=10.545 //y2=1.62
r69 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.46 //y=1.58 //x2=10.06 //y2=1.58
r70 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.575 //y=1.495 //x2=9.575 //y2=1.62
r71 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.575 //y=1.495 //x2=9.575 //y2=0.88
ends PM_MUX2X1\%noxref_12

