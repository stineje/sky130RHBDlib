magic
tech sky130A
magscale 1 2
timestamp 1652323563
<< nwell >>
rect 87 786 579 1550
<< pwell >>
rect 34 -34 632 544
<< pdiffc >>
rect 141 1331 175 1365
rect 229 1331 263 1365
rect 317 1331 351 1365
rect 493 1331 527 1365
rect 141 1059 175 1093
rect 317 1059 351 1093
rect 405 1059 439 1093
<< psubdiff >>
rect 34 482 632 544
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 632 17
rect 34 -34 632 -17
<< nsubdiff >>
rect 34 1497 632 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 632 1497
rect 34 822 632 884
<< psubdiffcont >>
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
<< poly >>
rect 168 375 198 413
rect 362 382 392 383
<< locali >>
rect 34 1497 632 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 632 1497
rect 34 1446 632 1463
rect 141 1365 175 1405
rect 141 1313 175 1331
rect 229 1365 263 1446
rect 229 1313 263 1331
rect 317 1365 527 1399
rect 317 1313 351 1331
rect 493 1313 527 1331
rect 141 1093 175 1111
rect 317 1093 351 1111
rect 141 1025 351 1059
rect 405 1093 439 1111
rect 405 1025 535 1059
rect 205 433 239 942
rect 353 908 361 942
rect 353 441 387 908
rect 353 433 357 441
rect 501 348 535 1025
rect 219 314 535 348
rect 219 233 253 314
rect 413 233 447 314
rect 122 34 156 73
rect 219 34 253 89
rect 316 34 350 73
rect 413 34 447 89
rect 510 34 544 73
rect 34 17 632 34
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 632 17
rect 34 -34 632 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
<< metal1 >>
rect 34 1497 632 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 632 1497
rect 34 1446 632 1463
rect 34 17 632 34
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 632 17
rect 34 -34 632 -17
use pmos2_1  pmos2_1_0
timestamp 1647326732
transform 1 0 43 0 1 1404
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 192 -1 0 942
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 223 -1 0 417
box -32 -28 34 26
use nmos_top_trim1  nmos_top_trim1_1
timestamp 1651256895
transform -1 0 360 0 1 73
box 0 0 248 309
use pmos2_1  pmos2_1_1
timestamp 1647326732
transform 1 0 219 0 1 1404
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 378 -1 0 942
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 -1 369 1 0 415
box -32 -28 34 26
use nmos_top_trim2  nmos_top_trim2_0
timestamp 1651256905
transform -1 0 554 0 1 73
box 0 0 248 309
use diff_ring_side  diff_ring_side_1
timestamp 1652319726
transform 1 0 0 0 1 0
box -87 -34 87 1550
use diff_ring_side  diff_ring_side_0
timestamp 1652319726
transform 1 0 666 0 1 0
box -87 -34 87 1550
<< end >>
