// File: DFFSNQX1.spi.pex
// Created: Tue Oct 15 15:47:07 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_DFFSNQX1\%GND ( 1 43 47 50 55 63 69 79 85 95 101 107 115 123 138 142 \
 145 148 151 153 155 156 157 158 159 160 )
c286 ( 160 0 ) capacitor c=0.0226075f //x=20.495 //y=0.875
c287 ( 159 0 ) capacitor c=0.0207407f //x=17.27 //y=0.865
c288 ( 158 0 ) capacitor c=0.0207407f //x=13.94 //y=0.865
c289 ( 157 0 ) capacitor c=0.0226205f //x=9.025 //y=0.875
c290 ( 156 0 ) capacitor c=0.0226323f //x=4.215 //y=0.875
c291 ( 155 0 ) capacitor c=0.0208404f //x=0.99 //y=0.865
c292 ( 154 0 ) capacitor c=0.00440144f //x=20.685 //y=0
c293 ( 153 0 ) capacitor c=0.104091f //x=19.61 //y=0
c294 ( 152 0 ) capacitor c=0.00440095f //x=17.46 //y=0
c295 ( 151 0 ) capacitor c=0.106174f //x=16.28 //y=0
c296 ( 150 0 ) capacitor c=0.00440095f //x=14.06 //y=0
c297 ( 148 0 ) capacitor c=0.108248f //x=12.95 //y=0
c298 ( 147 0 ) capacitor c=0.00440144f //x=9.25 //y=0
c299 ( 145 0 ) capacitor c=0.108235f //x=8.14 //y=0
c300 ( 144 0 ) capacitor c=0.00440144f //x=4.44 //y=0
c301 ( 142 0 ) capacitor c=0.105313f //x=3.33 //y=0
c302 ( 141 0 ) capacitor c=0.00440095f //x=1.18 //y=0
c303 ( 138 0 ) capacitor c=0.324351f //x=23.68 //y=0
c304 ( 123 0 ) capacitor c=0.0339325f //x=20.6 //y=0
c305 ( 115 0 ) capacitor c=0.0718026f //x=19.44 //y=0
c306 ( 107 0 ) capacitor c=0.0388888f //x=17.375 //y=0
c307 ( 101 0 ) capacitor c=0.0718026f //x=16.11 //y=0
c308 ( 95 0 ) capacitor c=0.0388888f //x=14.045 //y=0
c309 ( 85 0 ) capacitor c=0.133402f //x=12.78 //y=0
c310 ( 79 0 ) capacitor c=0.0339482f //x=9.13 //y=0
c311 ( 69 0 ) capacitor c=0.133515f //x=7.97 //y=0
c312 ( 63 0 ) capacitor c=0.0339482f //x=4.32 //y=0
c313 ( 55 0 ) capacitor c=0.0720582f //x=3.16 //y=0
c314 ( 50 0 ) capacitor c=0.179262f //x=0.74 //y=0
c315 ( 47 0 ) capacitor c=0.0426751f //x=1.095 //y=0
c316 ( 43 0 ) capacitor c=0.775533f //x=23.68 //y=0
r317 (  136 138 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=22.57 //y=0 //x2=23.68 //y2=0
r318 (  134 136 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.46 //y=0 //x2=22.57 //y2=0
r319 (  132 154 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.77 //y=0 //x2=20.685 //y2=0
r320 (  132 134 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=20.77 //y=0 //x2=21.46 //y2=0
r321 (  127 154 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.685 //y=0.17 //x2=20.685 //y2=0
r322 (  127 160 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=20.685 //y=0.17 //x2=20.685 //y2=0.965
r323 (  124 153 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.78 //y=0 //x2=19.61 //y2=0
r324 (  124 126 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.78 //y=0 //x2=20.35 //y2=0
r325 (  123 154 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.6 //y=0 //x2=20.685 //y2=0
r326 (  123 126 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=20.6 //y=0 //x2=20.35 //y2=0
r327 (  118 120 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.76 //y=0 //x2=18.87 //y2=0
r328 (  116 152 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.545 //y=0 //x2=17.46 //y2=0
r329 (  116 118 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=17.545 //y=0 //x2=17.76 //y2=0
r330 (  115 153 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.44 //y=0 //x2=19.61 //y2=0
r331 (  115 120 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.44 //y=0 //x2=18.87 //y2=0
r332 (  111 152 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.46 //y=0.17 //x2=17.46 //y2=0
r333 (  111 159 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=17.46 //y=0.17 //x2=17.46 //y2=0.955
r334 (  108 151 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.45 //y=0 //x2=16.28 //y2=0
r335 (  108 110 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=16.45 //y=0 //x2=16.65 //y2=0
r336 (  107 152 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.375 //y=0 //x2=17.46 //y2=0
r337 (  107 110 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=17.375 //y=0 //x2=16.65 //y2=0
r338 (  102 150 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.215 //y=0 //x2=14.13 //y2=0
r339 (  102 104 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=14.215 //y=0 //x2=15.17 //y2=0
r340 (  101 151 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.11 //y=0 //x2=16.28 //y2=0
r341 (  101 104 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=16.11 //y=0 //x2=15.17 //y2=0
r342 (  97 150 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.13 //y=0.17 //x2=14.13 //y2=0
r343 (  97 158 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=14.13 //y=0.17 //x2=14.13 //y2=0.955
r344 (  96 148 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=0 //x2=12.95 //y2=0
r345 (  95 150 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.045 //y=0 //x2=14.13 //y2=0
r346 (  95 96 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=14.045 //y=0 //x2=13.12 //y2=0
r347 (  90 92 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r348 (  88 90 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=10.36 //y=0 //x2=11.47 //y2=0
r349 (  86 147 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.3 //y=0 //x2=9.215 //y2=0
r350 (  86 88 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=9.3 //y=0 //x2=10.36 //y2=0
r351 (  85 148 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.95 //y2=0
r352 (  85 92 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.58 //y2=0
r353 (  81 147 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.215 //y=0.17 //x2=9.215 //y2=0
r354 (  81 157 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=9.215 //y=0.17 //x2=9.215 //y2=0.965
r355 (  80 145 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=0 //x2=8.14 //y2=0
r356 (  79 147 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.13 //y=0 //x2=9.215 //y2=0
r357 (  79 80 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=9.13 //y=0 //x2=8.31 //y2=0
r358 (  74 76 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r359 (  72 74 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=5.55 //y=0 //x2=6.66 //y2=0
r360 (  70 144 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.49 //y=0 //x2=4.405 //y2=0
r361 (  70 72 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=4.49 //y=0 //x2=5.55 //y2=0
r362 (  69 145 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=8.14 //y2=0
r363 (  69 76 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=7.77 //y2=0
r364 (  65 144 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.405 //y=0.17 //x2=4.405 //y2=0
r365 (  65 156 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=4.405 //y=0.17 //x2=4.405 //y2=0.965
r366 (  64 142 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=0 //x2=3.33 //y2=0
r367 (  63 144 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.32 //y=0 //x2=4.405 //y2=0
r368 (  63 64 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=4.32 //y=0 //x2=3.5 //y2=0
r369 (  58 60 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r370 (  56 141 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.18 //y2=0
r371 (  56 58 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.85 //y2=0
r372 (  55 142 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=3.33 //y2=0
r373 (  55 60 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r374 (  51 141 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r375 (  51 155 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.955
r376 (  47 141 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=1.18 //y2=0
r377 (  47 50 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=0.74 //y2=0
r378 (  43 138 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=0 //x2=23.68 //y2=0
r379 (  41 136 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=0 //x2=22.57 //y2=0
r380 (  41 43 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=0 //x2=23.68 //y2=0
r381 (  39 134 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.46 //y=0 //x2=21.46 //y2=0
r382 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.46 //y=0 //x2=22.57 //y2=0
r383 (  37 126 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=0 //x2=20.35 //y2=0
r384 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=0 //x2=21.46 //y2=0
r385 (  35 120 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=0 //x2=18.87 //y2=0
r386 (  35 37 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=0 //x2=20.35 //y2=0
r387 (  33 118 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=0 //x2=17.76 //y2=0
r388 (  33 35 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=0 //x2=18.87 //y2=0
r389 (  31 110 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=0 //x2=16.65 //y2=0
r390 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=0 //x2=17.76 //y2=0
r391 (  29 104 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r392 (  29 31 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.65 //y2=0
r393 (  27 150 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=0 //x2=14.06 //y2=0
r394 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=0 //x2=15.17 //y2=0
r395 (  25 92 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r396 (  25 27 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=0 //x2=14.06 //y2=0
r397 (  22 90 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r398 (  20 88 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r399 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r400 (  18 147 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=0 //x2=9.25 //y2=0
r401 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=0 //x2=10.36 //y2=0
r402 (  16 76 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r403 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=9.25 //y2=0
r404 (  14 74 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r405 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r406 (  12 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r407 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r408 (  10 144 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r409 (  10 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.55 //y2=0
r410 (  8 60 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r411 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r412 (  6 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r413 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r414 (  3 50 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r415 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r416 (  1 25 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=0 //x2=12.58 //y2=0
r417 (  1 22 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=0 //x2=11.47 //y2=0
ends PM_DFFSNQX1\%GND

subckt PM_DFFSNQX1\%VDD ( 1 43 55 63 73 79 87 95 105 115 121 129 137 147 157 \
 163 171 181 191 195 205 215 237 247 255 268 272 275 281 287 291 296 301 302 \
 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 )
c304 ( 321 0 ) capacitor c=0.0454188f //x=23.195 //y=5.02
c305 ( 320 0 ) capacitor c=0.0243052f //x=22.315 //y=5.02
c306 ( 319 0 ) capacitor c=0.0243052f //x=21.435 //y=5.02
c307 ( 318 0 ) capacitor c=0.0532751f //x=20.565 //y=5.02
c308 ( 317 0 ) capacitor c=0.0382117f //x=18.685 //y=5.02
c309 ( 316 0 ) capacitor c=0.024147f //x=17.805 //y=5.02
c310 ( 315 0 ) capacitor c=0.0493657f //x=16.935 //y=5.02
c311 ( 314 0 ) capacitor c=0.0381505f //x=15.355 //y=5.02
c312 ( 313 0 ) capacitor c=0.0240074f //x=14.475 //y=5.02
c313 ( 312 0 ) capacitor c=0.049209f //x=13.605 //y=5.02
c314 ( 311 0 ) capacitor c=0.0452179f //x=11.725 //y=5.02
c315 ( 310 0 ) capacitor c=0.024152f //x=10.845 //y=5.02
c316 ( 309 0 ) capacitor c=0.024152f //x=9.965 //y=5.02
c317 ( 308 0 ) capacitor c=0.053132f //x=9.095 //y=5.02
c318 ( 307 0 ) capacitor c=0.0452179f //x=6.915 //y=5.02
c319 ( 306 0 ) capacitor c=0.024152f //x=6.035 //y=5.02
c320 ( 305 0 ) capacitor c=0.02424f //x=5.155 //y=5.02
c321 ( 304 0 ) capacitor c=0.0532367f //x=4.285 //y=5.02
c322 ( 303 0 ) capacitor c=0.0381505f //x=2.405 //y=5.02
c323 ( 302 0 ) capacitor c=0.024246f //x=1.525 //y=5.02
c324 ( 301 0 ) capacitor c=0.053196f //x=0.655 //y=5.02
c325 ( 300 0 ) capacitor c=0.00591168f //x=23.34 //y=7.4
c326 ( 299 0 ) capacitor c=0.00591168f //x=22.46 //y=7.4
c327 ( 298 0 ) capacitor c=0.00591168f //x=21.58 //y=7.4
c328 ( 297 0 ) capacitor c=0.00591168f //x=20.7 //y=7.4
c329 ( 296 0 ) capacitor c=0.139422f //x=19.61 //y=7.4
c330 ( 295 0 ) capacitor c=0.00591168f //x=18.87 //y=7.4
c331 ( 293 0 ) capacitor c=0.00591168f //x=17.95 //y=7.4
c332 ( 292 0 ) capacitor c=0.00591168f //x=17.07 //y=7.4
c333 ( 291 0 ) capacitor c=0.116163f //x=16.28 //y=7.4
c334 ( 290 0 ) capacitor c=0.00591168f //x=15.5 //y=7.4
c335 ( 289 0 ) capacitor c=0.00591168f //x=14.62 //y=7.4
c336 ( 288 0 ) capacitor c=0.00591168f //x=13.74 //y=7.4
c337 ( 287 0 ) capacitor c=0.13452f //x=12.95 //y=7.4
c338 ( 286 0 ) capacitor c=0.00591168f //x=11.87 //y=7.4
c339 ( 285 0 ) capacitor c=0.00591168f //x=10.99 //y=7.4
c340 ( 284 0 ) capacitor c=0.00591168f //x=10.11 //y=7.4
c341 ( 283 0 ) capacitor c=0.00591168f //x=9.25 //y=7.4
c342 ( 281 0 ) capacitor c=0.155082f //x=8.14 //y=7.4
c343 ( 280 0 ) capacitor c=0.00591168f //x=7.06 //y=7.4
c344 ( 279 0 ) capacitor c=0.00591168f //x=6.18 //y=7.4
c345 ( 278 0 ) capacitor c=0.00591168f //x=5.3 //y=7.4
c346 ( 277 0 ) capacitor c=0.00591168f //x=4.44 //y=7.4
c347 ( 275 0 ) capacitor c=0.137403f //x=3.33 //y=7.4
c348 ( 274 0 ) capacitor c=0.00591168f //x=2.55 //y=7.4
c349 ( 273 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c350 ( 272 0 ) capacitor c=0.248311f //x=0.74 //y=7.4
c351 ( 268 0 ) capacitor c=0.272255f //x=23.68 //y=7.4
c352 ( 255 0 ) capacitor c=0.028513f //x=23.255 //y=7.4
c353 ( 247 0 ) capacitor c=0.0287069f //x=22.375 //y=7.4
c354 ( 237 0 ) capacitor c=0.0292055f //x=21.495 //y=7.4
c355 ( 227 0 ) capacitor c=0.0452081f //x=20.615 //y=7.4
c356 ( 223 0 ) capacitor c=0.0275781f //x=19.44 //y=7.4
c357 ( 215 0 ) capacitor c=0.0285035f //x=18.745 //y=7.4
c358 ( 205 0 ) capacitor c=0.0291038f //x=17.865 //y=7.4
c359 ( 195 0 ) capacitor c=0.0240981f //x=16.985 //y=7.4
c360 ( 191 0 ) capacitor c=0.0236224f //x=16.11 //y=7.4
c361 ( 181 0 ) capacitor c=0.0288598f //x=15.415 //y=7.4
c362 ( 171 0 ) capacitor c=0.0288369f //x=14.535 //y=7.4
c363 ( 163 0 ) capacitor c=0.0240981f //x=13.655 //y=7.4
c364 ( 157 0 ) capacitor c=0.0394667f //x=12.78 //y=7.4
c365 ( 147 0 ) capacitor c=0.0288488f //x=11.785 //y=7.4
c366 ( 137 0 ) capacitor c=0.0287514f //x=10.905 //y=7.4
c367 ( 129 0 ) capacitor c=0.0284966f //x=10.025 //y=7.4
c368 ( 121 0 ) capacitor c=0.0383672f //x=9.145 //y=7.4
c369 ( 115 0 ) capacitor c=0.0394667f //x=7.97 //y=7.4
c370 ( 105 0 ) capacitor c=0.0288488f //x=6.975 //y=7.4
c371 ( 95 0 ) capacitor c=0.0287505f //x=6.095 //y=7.4
c372 ( 87 0 ) capacitor c=0.028511f //x=5.215 //y=7.4
c373 ( 79 0 ) capacitor c=0.0383672f //x=4.335 //y=7.4
c374 ( 73 0 ) capacitor c=0.0236224f //x=3.16 //y=7.4
c375 ( 63 0 ) capacitor c=0.0288637f //x=2.465 //y=7.4
c376 ( 55 0 ) capacitor c=0.0286367f //x=1.585 //y=7.4
c377 ( 43 0 ) capacitor c=0.851956f //x=23.68 //y=7.4
r378 (  266 300 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.425 //y=7.4 //x2=23.34 //y2=7.4
r379 (  266 268 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=23.425 //y=7.4 //x2=23.68 //y2=7.4
r380 (  259 300 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.34 //y=7.23 //x2=23.34 //y2=7.4
r381 (  259 321 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=23.34 //y=7.23 //x2=23.34 //y2=6.745
r382 (  256 299 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.545 //y=7.4 //x2=22.46 //y2=7.4
r383 (  256 258 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=22.545 //y=7.4 //x2=22.57 //y2=7.4
r384 (  255 300 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.255 //y=7.4 //x2=23.34 //y2=7.4
r385 (  255 258 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=23.255 //y=7.4 //x2=22.57 //y2=7.4
r386 (  249 299 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.46 //y=7.23 //x2=22.46 //y2=7.4
r387 (  249 320 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.46 //y=7.23 //x2=22.46 //y2=6.745
r388 (  248 298 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.665 //y=7.4 //x2=21.58 //y2=7.4
r389 (  247 299 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.375 //y=7.4 //x2=22.46 //y2=7.4
r390 (  247 248 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.375 //y=7.4 //x2=21.665 //y2=7.4
r391 (  241 298 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.58 //y=7.23 //x2=21.58 //y2=7.4
r392 (  241 319 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.58 //y=7.23 //x2=21.58 //y2=6.745
r393 (  238 297 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.785 //y=7.4 //x2=20.7 //y2=7.4
r394 (  238 240 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=20.785 //y=7.4 //x2=21.46 //y2=7.4
r395 (  237 298 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.495 //y=7.4 //x2=21.58 //y2=7.4
r396 (  237 240 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=21.495 //y=7.4 //x2=21.46 //y2=7.4
r397 (  231 297 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.7 //y=7.23 //x2=20.7 //y2=7.4
r398 (  231 318 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=20.7 //y=7.23 //x2=20.7 //y2=6.405
r399 (  228 296 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.78 //y=7.4 //x2=19.61 //y2=7.4
r400 (  228 230 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.78 //y=7.4 //x2=20.35 //y2=7.4
r401 (  227 297 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.615 //y=7.4 //x2=20.7 //y2=7.4
r402 (  227 230 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.615 //y=7.4 //x2=20.35 //y2=7.4
r403 (  224 295 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.915 //y=7.4 //x2=18.83 //y2=7.4
r404 (  223 296 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.44 //y=7.4 //x2=19.61 //y2=7.4
r405 (  223 224 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=19.44 //y=7.4 //x2=18.915 //y2=7.4
r406 (  217 295 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.83 //y=7.23 //x2=18.83 //y2=7.4
r407 (  217 317 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=18.83 //y=7.23 //x2=18.83 //y2=6.745
r408 (  216 293 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.035 //y=7.4 //x2=17.95 //y2=7.4
r409 (  215 295 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.745 //y=7.4 //x2=18.83 //y2=7.4
r410 (  215 216 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=18.745 //y=7.4 //x2=18.035 //y2=7.4
r411 (  209 293 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.95 //y=7.23 //x2=17.95 //y2=7.4
r412 (  209 316 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.95 //y=7.23 //x2=17.95 //y2=6.745
r413 (  206 292 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.155 //y=7.4 //x2=17.07 //y2=7.4
r414 (  206 208 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=17.155 //y=7.4 //x2=17.76 //y2=7.4
r415 (  205 293 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.865 //y=7.4 //x2=17.95 //y2=7.4
r416 (  205 208 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=17.865 //y=7.4 //x2=17.76 //y2=7.4
r417 (  199 292 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.07 //y=7.23 //x2=17.07 //y2=7.4
r418 (  199 315 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=17.07 //y=7.23 //x2=17.07 //y2=6.405
r419 (  196 291 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.45 //y=7.4 //x2=16.28 //y2=7.4
r420 (  196 198 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=16.45 //y=7.4 //x2=16.65 //y2=7.4
r421 (  195 292 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.985 //y=7.4 //x2=17.07 //y2=7.4
r422 (  195 198 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=16.985 //y=7.4 //x2=16.65 //y2=7.4
r423 (  192 290 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.585 //y=7.4 //x2=15.5 //y2=7.4
r424 (  191 291 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.11 //y=7.4 //x2=16.28 //y2=7.4
r425 (  191 192 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=16.11 //y=7.4 //x2=15.585 //y2=7.4
r426 (  185 290 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.5 //y=7.23 //x2=15.5 //y2=7.4
r427 (  185 314 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.5 //y=7.23 //x2=15.5 //y2=6.745
r428 (  182 289 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.705 //y=7.4 //x2=14.62 //y2=7.4
r429 (  182 184 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=14.705 //y=7.4 //x2=15.17 //y2=7.4
r430 (  181 290 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.415 //y=7.4 //x2=15.5 //y2=7.4
r431 (  181 184 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=15.415 //y=7.4 //x2=15.17 //y2=7.4
r432 (  175 289 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.62 //y=7.23 //x2=14.62 //y2=7.4
r433 (  175 313 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.62 //y=7.23 //x2=14.62 //y2=6.745
r434 (  172 288 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.825 //y=7.4 //x2=13.74 //y2=7.4
r435 (  172 174 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=13.825 //y=7.4 //x2=14.06 //y2=7.4
r436 (  171 289 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.535 //y=7.4 //x2=14.62 //y2=7.4
r437 (  171 174 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=14.535 //y=7.4 //x2=14.06 //y2=7.4
r438 (  165 288 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.74 //y=7.23 //x2=13.74 //y2=7.4
r439 (  165 312 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=13.74 //y=7.23 //x2=13.74 //y2=6.405
r440 (  164 287 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=7.4 //x2=12.95 //y2=7.4
r441 (  163 288 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.655 //y=7.4 //x2=13.74 //y2=7.4
r442 (  163 164 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=13.655 //y=7.4 //x2=13.12 //y2=7.4
r443 (  158 286 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.955 //y=7.4 //x2=11.87 //y2=7.4
r444 (  158 160 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=11.955 //y=7.4 //x2=12.58 //y2=7.4
r445 (  157 287 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.95 //y2=7.4
r446 (  157 160 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.58 //y2=7.4
r447 (  151 286 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.87 //y=7.23 //x2=11.87 //y2=7.4
r448 (  151 311 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.87 //y=7.23 //x2=11.87 //y2=6.745
r449 (  148 285 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.075 //y=7.4 //x2=10.99 //y2=7.4
r450 (  148 150 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=11.075 //y=7.4 //x2=11.47 //y2=7.4
r451 (  147 286 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.785 //y=7.4 //x2=11.87 //y2=7.4
r452 (  147 150 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=11.785 //y=7.4 //x2=11.47 //y2=7.4
r453 (  141 285 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.99 //y=7.23 //x2=10.99 //y2=7.4
r454 (  141 310 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.99 //y=7.23 //x2=10.99 //y2=6.745
r455 (  138 284 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.195 //y=7.4 //x2=10.11 //y2=7.4
r456 (  138 140 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=10.195 //y=7.4 //x2=10.36 //y2=7.4
r457 (  137 285 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.905 //y=7.4 //x2=10.99 //y2=7.4
r458 (  137 140 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=10.905 //y=7.4 //x2=10.36 //y2=7.4
r459 (  131 284 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.11 //y=7.23 //x2=10.11 //y2=7.4
r460 (  131 309 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.11 //y=7.23 //x2=10.11 //y2=6.745
r461 (  130 283 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.315 //y=7.4 //x2=9.23 //y2=7.4
r462 (  129 284 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.025 //y=7.4 //x2=10.11 //y2=7.4
r463 (  129 130 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.025 //y=7.4 //x2=9.315 //y2=7.4
r464 (  123 283 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.23 //y=7.23 //x2=9.23 //y2=7.4
r465 (  123 308 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=9.23 //y=7.23 //x2=9.23 //y2=6.405
r466 (  122 281 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=7.4 //x2=8.14 //y2=7.4
r467 (  121 283 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.145 //y=7.4 //x2=9.23 //y2=7.4
r468 (  121 122 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=9.145 //y=7.4 //x2=8.31 //y2=7.4
r469 (  116 280 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.145 //y=7.4 //x2=7.06 //y2=7.4
r470 (  116 118 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=7.145 //y=7.4 //x2=7.77 //y2=7.4
r471 (  115 281 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=8.14 //y2=7.4
r472 (  115 118 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=7.77 //y2=7.4
r473 (  109 280 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.06 //y=7.23 //x2=7.06 //y2=7.4
r474 (  109 307 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.06 //y=7.23 //x2=7.06 //y2=6.745
r475 (  106 279 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.265 //y=7.4 //x2=6.18 //y2=7.4
r476 (  106 108 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=6.265 //y=7.4 //x2=6.66 //y2=7.4
r477 (  105 280 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.975 //y=7.4 //x2=7.06 //y2=7.4
r478 (  105 108 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=6.975 //y=7.4 //x2=6.66 //y2=7.4
r479 (  99 279 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.18 //y=7.23 //x2=6.18 //y2=7.4
r480 (  99 306 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.18 //y=7.23 //x2=6.18 //y2=6.745
r481 (  96 278 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.385 //y=7.4 //x2=5.3 //y2=7.4
r482 (  96 98 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=5.385 //y=7.4 //x2=5.55 //y2=7.4
r483 (  95 279 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.095 //y=7.4 //x2=6.18 //y2=7.4
r484 (  95 98 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=6.095 //y=7.4 //x2=5.55 //y2=7.4
r485 (  89 278 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.3 //y=7.23 //x2=5.3 //y2=7.4
r486 (  89 305 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=5.3 //y=7.23 //x2=5.3 //y2=6.745
r487 (  88 277 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.505 //y=7.4 //x2=4.42 //y2=7.4
r488 (  87 278 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.215 //y=7.4 //x2=5.3 //y2=7.4
r489 (  87 88 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.215 //y=7.4 //x2=4.505 //y2=7.4
r490 (  81 277 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.42 //y=7.23 //x2=4.42 //y2=7.4
r491 (  81 304 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.42 //y=7.23 //x2=4.42 //y2=6.405
r492 (  80 275 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r493 (  79 277 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.335 //y=7.4 //x2=4.42 //y2=7.4
r494 (  79 80 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=4.335 //y=7.4 //x2=3.5 //y2=7.4
r495 (  74 274 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.55 //y2=7.4
r496 (  74 76 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.96 //y2=7.4
r497 (  73 275 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r498 (  73 76 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r499 (  67 274 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r500 (  67 303 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.745
r501 (  64 273 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r502 (  64 66 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r503 (  63 274 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r504 (  63 66 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r505 (  57 273 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r506 (  57 302 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.745
r507 (  56 272 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r508 (  55 273 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r509 (  55 56 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r510 (  49 272 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r511 (  49 301 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.405
r512 (  43 268 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=7.4 //x2=23.68 //y2=7.4
r513 (  41 258 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=7.4 //x2=22.57 //y2=7.4
r514 (  41 43 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=7.4 //x2=23.68 //y2=7.4
r515 (  39 240 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.46 //y=7.4 //x2=21.46 //y2=7.4
r516 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.46 //y=7.4 //x2=22.57 //y2=7.4
r517 (  37 230 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=7.4 //x2=20.35 //y2=7.4
r518 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=7.4 //x2=21.46 //y2=7.4
r519 (  35 295 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=7.4 //x2=18.87 //y2=7.4
r520 (  35 37 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=7.4 //x2=20.35 //y2=7.4
r521 (  33 208 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=7.4 //x2=17.76 //y2=7.4
r522 (  33 35 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=7.4 //x2=18.87 //y2=7.4
r523 (  31 198 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=7.4 //x2=16.65 //y2=7.4
r524 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=7.4 //x2=17.76 //y2=7.4
r525 (  29 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r526 (  29 31 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.65 //y2=7.4
r527 (  27 174 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=7.4 //x2=14.06 //y2=7.4
r528 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=7.4 //x2=15.17 //y2=7.4
r529 (  25 160 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r530 (  25 27 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.4 //x2=14.06 //y2=7.4
r531 (  22 150 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r532 (  20 140 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r533 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r534 (  18 283 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=7.4 //x2=9.25 //y2=7.4
r535 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=7.4 //x2=10.36 //y2=7.4
r536 (  16 118 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r537 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=9.25 //y2=7.4
r538 (  14 108 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r539 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r540 (  12 98 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r541 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r542 (  10 277 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r543 (  10 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.55 //y2=7.4
r544 (  8 76 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r545 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r546 (  6 66 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r547 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r548 (  3 272 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r549 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r550 (  1 25 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=7.4 //x2=12.58 //y2=7.4
r551 (  1 22 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=7.4 //x2=11.47 //y2=7.4
ends PM_DFFSNQX1\%VDD

subckt PM_DFFSNQX1\%noxref_3 ( 1 2 3 4 17 18 29 31 32 36 38 46 53 54 55 56 57 \
 58 59 60 61 62 63 64 66 72 73 74 75 79 80 81 82 83 85 91 92 93 94 114 116 117 )
c240 ( 117 0 ) capacitor c=0.0220291f //x=1.965 //y=5.02
c241 ( 116 0 ) capacitor c=0.0217503f //x=1.085 //y=5.02
c242 ( 114 0 ) capacitor c=0.0084702f //x=1.96 //y=0.905
c243 ( 94 0 ) capacitor c=0.0556143f //x=9.525 //y=4.79
c244 ( 93 0 ) capacitor c=0.0293157f //x=9.815 //y=4.79
c245 ( 92 0 ) capacitor c=0.0347816f //x=9.48 //y=1.22
c246 ( 91 0 ) capacitor c=0.0187487f //x=9.48 //y=0.875
c247 ( 85 0 ) capacitor c=0.0137055f //x=9.325 //y=1.375
c248 ( 83 0 ) capacitor c=0.0149861f //x=9.325 //y=0.72
c249 ( 82 0 ) capacitor c=0.0965257f //x=8.95 //y=1.915
c250 ( 81 0 ) capacitor c=0.0229444f //x=8.95 //y=1.53
c251 ( 80 0 ) capacitor c=0.0234352f //x=8.95 //y=1.22
c252 ( 79 0 ) capacitor c=0.0198724f //x=8.95 //y=0.875
c253 ( 75 0 ) capacitor c=0.055995f //x=4.715 //y=4.79
c254 ( 74 0 ) capacitor c=0.0298189f //x=5.005 //y=4.79
c255 ( 73 0 ) capacitor c=0.0347816f //x=4.67 //y=1.22
c256 ( 72 0 ) capacitor c=0.0187487f //x=4.67 //y=0.875
c257 ( 66 0 ) capacitor c=0.0137055f //x=4.515 //y=1.375
c258 ( 64 0 ) capacitor c=0.0149861f //x=4.515 //y=0.72
c259 ( 63 0 ) capacitor c=0.0965245f //x=4.14 //y=1.915
c260 ( 62 0 ) capacitor c=0.0229444f //x=4.14 //y=1.53
c261 ( 61 0 ) capacitor c=0.0234352f //x=4.14 //y=1.22
c262 ( 60 0 ) capacitor c=0.0198724f //x=4.14 //y=0.875
c263 ( 59 0 ) capacitor c=0.110114f //x=9.89 //y=6.02
c264 ( 58 0 ) capacitor c=0.158956f //x=9.45 //y=6.02
c265 ( 57 0 ) capacitor c=0.110114f //x=5.08 //y=6.02
c266 ( 56 0 ) capacitor c=0.158956f //x=4.64 //y=6.02
c267 ( 53 0 ) capacitor c=0.0023043f //x=2.11 //y=5.2
c268 ( 46 0 ) capacitor c=0.10363f //x=9.25 //y=2.08
c269 ( 38 0 ) capacitor c=0.108245f //x=4.44 //y=2.08
c270 ( 36 0 ) capacitor c=0.114138f //x=2.59 //y=2.59
c271 ( 32 0 ) capacitor c=0.00550359f //x=2.235 //y=1.655
c272 ( 31 0 ) capacitor c=0.0140493f //x=2.505 //y=1.655
c273 ( 29 0 ) capacitor c=0.0140934f //x=2.505 //y=5.2
c274 ( 18 0 ) capacitor c=0.00387264f //x=1.315 //y=5.2
c275 ( 17 0 ) capacitor c=0.019002f //x=2.025 //y=5.2
c276 ( 4 0 ) capacitor c=0.012652f //x=4.705 //y=2.59
c277 ( 3 0 ) capacitor c=0.143287f //x=9.135 //y=2.59
c278 ( 2 0 ) capacitor c=0.0148669f //x=2.705 //y=2.59
c279 ( 1 0 ) capacitor c=0.0543359f //x=4.295 //y=2.59
r280 (  93 95 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.815 //y=4.79 //x2=9.89 //y2=4.865
r281 (  93 94 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=9.815 //y=4.79 //x2=9.525 //y2=4.79
r282 (  92 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.48 //y=1.22 //x2=9.44 //y2=1.375
r283 (  91 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.48 //y=0.875 //x2=9.44 //y2=0.72
r284 (  91 92 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.48 //y=0.875 //x2=9.48 //y2=1.22
r285 (  88 94 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.45 //y=4.865 //x2=9.525 //y2=4.79
r286 (  88 111 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=9.45 //y=4.865 //x2=9.25 //y2=4.7
r287 (  86 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.105 //y=1.375 //x2=8.99 //y2=1.375
r288 (  85 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.325 //y=1.375 //x2=9.44 //y2=1.375
r289 (  84 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.105 //y=0.72 //x2=8.99 //y2=0.72
r290 (  83 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.325 //y=0.72 //x2=9.44 //y2=0.72
r291 (  83 84 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=9.325 //y=0.72 //x2=9.105 //y2=0.72
r292 (  82 109 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.915 //x2=9.25 //y2=2.08
r293 (  81 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.53 //x2=8.99 //y2=1.375
r294 (  81 82 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.53 //x2=8.95 //y2=1.915
r295 (  80 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.22 //x2=8.99 //y2=1.375
r296 (  79 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=0.875 //x2=8.99 //y2=0.72
r297 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.95 //y=0.875 //x2=8.95 //y2=1.22
r298 (  74 76 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.005 //y=4.79 //x2=5.08 //y2=4.865
r299 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=5.005 //y=4.79 //x2=4.715 //y2=4.79
r300 (  73 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.67 //y=1.22 //x2=4.63 //y2=1.375
r301 (  72 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.67 //y=0.875 //x2=4.63 //y2=0.72
r302 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.67 //y=0.875 //x2=4.67 //y2=1.22
r303 (  69 75 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.64 //y=4.865 //x2=4.715 //y2=4.79
r304 (  69 103 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=4.64 //y=4.865 //x2=4.44 //y2=4.7
r305 (  67 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.295 //y=1.375 //x2=4.18 //y2=1.375
r306 (  66 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.515 //y=1.375 //x2=4.63 //y2=1.375
r307 (  65 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.295 //y=0.72 //x2=4.18 //y2=0.72
r308 (  64 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.515 //y=0.72 //x2=4.63 //y2=0.72
r309 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.515 //y=0.72 //x2=4.295 //y2=0.72
r310 (  63 101 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.915 //x2=4.44 //y2=2.08
r311 (  62 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.53 //x2=4.18 //y2=1.375
r312 (  62 63 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.53 //x2=4.14 //y2=1.915
r313 (  61 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.22 //x2=4.18 //y2=1.375
r314 (  60 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=0.875 //x2=4.18 //y2=0.72
r315 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.14 //y=0.875 //x2=4.14 //y2=1.22
r316 (  59 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.89 //y=6.02 //x2=9.89 //y2=4.865
r317 (  58 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.45 //y=6.02 //x2=9.45 //y2=4.865
r318 (  57 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.08 //y=6.02 //x2=5.08 //y2=4.865
r319 (  56 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.64 //y=6.02 //x2=4.64 //y2=4.865
r320 (  55 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.375 //x2=9.325 //y2=1.375
r321 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.375 //x2=9.105 //y2=1.375
r322 (  54 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.405 //y=1.375 //x2=4.515 //y2=1.375
r323 (  54 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.405 //y=1.375 //x2=4.295 //y2=1.375
r324 (  51 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=4.7 //x2=9.25 //y2=4.7
r325 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.59 //x2=9.25 //y2=4.7
r326 (  46 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=2.08 //x2=9.25 //y2=2.08
r327 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.08 //x2=9.25 //y2=2.59
r328 (  43 103 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=4.7 //x2=4.44 //y2=4.7
r329 (  41 43 ) resistor r=144.77 //w=0.187 //l=2.115 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.585 //x2=4.44 //y2=4.7
r330 (  38 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=2.08 //x2=4.44 //y2=2.08
r331 (  38 41 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.08 //x2=4.44 //y2=2.585
r332 (  34 36 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.115 //x2=2.59 //y2=2.59
r333 (  33 36 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=2.59
r334 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r335 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r336 (  30 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.195 //y=5.2 //x2=2.11 //y2=5.2
r337 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.59 //y2=5.115
r338 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.195 //y2=5.2
r339 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.235 //y2=1.655
r340 (  25 114 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r341 (  19 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.2
r342 (  19 117 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.725
r343 (  17 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=2.11 //y2=5.2
r344 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=1.315 //y2=5.2
r345 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.315 //y2=5.2
r346 (  11 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.23 //y2=5.725
r347 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.25 //y=2.59 //x2=9.25 //y2=2.59
r348 (  8 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=2.585 //x2=4.44 //y2=2.585
r349 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=2.59 //x2=2.59 //y2=2.59
r350 (  4 8 ) resistor r=0.164988 //w=0.206 //l=0.267488 //layer=m1 \
 //thickness=0.36 //x=4.705 //y=2.59 //x2=4.44 //y2=2.585
r351 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.135 //y=2.59 //x2=9.25 //y2=2.59
r352 (  3 4 ) resistor r=4.2271 //w=0.131 //l=4.43 //layer=m1 //thickness=0.36 \
 //x=9.135 //y=2.59 //x2=4.705 //y2=2.59
r353 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=2.59 //x2=2.59 //y2=2.59
r354 (  1 8 ) resistor r=0.0921728 //w=0.206 //l=0.147479 //layer=m1 \
 //thickness=0.36 //x=4.295 //y=2.59 //x2=4.44 //y2=2.585
r355 (  1 2 ) resistor r=1.51718 //w=0.131 //l=1.59 //layer=m1 \
 //thickness=0.36 //x=4.295 //y=2.59 //x2=2.705 //y2=2.59
ends PM_DFFSNQX1\%noxref_3

subckt PM_DFFSNQX1\%noxref_4 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 54 \
 55 56 57 61 63 66 67 77 80 82 83 84 )
c160 ( 84 0 ) capacitor c=0.023087f //x=11.285 //y=5.02
c161 ( 83 0 ) capacitor c=0.023519f //x=10.405 //y=5.02
c162 ( 82 0 ) capacitor c=0.0224735f //x=9.525 //y=5.02
c163 ( 80 0 ) capacitor c=0.00872971f //x=11.535 //y=0.915
c164 ( 77 0 ) capacitor c=0.0588816f //x=14.06 //y=4.7
c165 ( 67 0 ) capacitor c=0.0318948f //x=14.395 //y=1.21
c166 ( 66 0 ) capacitor c=0.0187384f //x=14.395 //y=0.865
c167 ( 63 0 ) capacitor c=0.0141798f //x=14.24 //y=1.365
c168 ( 61 0 ) capacitor c=0.0149844f //x=14.24 //y=0.71
c169 ( 57 0 ) capacitor c=0.0813322f //x=13.865 //y=1.915
c170 ( 56 0 ) capacitor c=0.0229267f //x=13.865 //y=1.52
c171 ( 55 0 ) capacitor c=0.0234352f //x=13.865 //y=1.21
c172 ( 54 0 ) capacitor c=0.0199343f //x=13.865 //y=0.865
c173 ( 53 0 ) capacitor c=0.110275f //x=14.4 //y=6.02
c174 ( 52 0 ) capacitor c=0.154305f //x=13.96 //y=6.02
c175 ( 50 0 ) capacitor c=0.00106608f //x=11.43 //y=5.155
c176 ( 49 0 ) capacitor c=0.00207319f //x=10.55 //y=5.155
c177 ( 42 0 ) capacitor c=0.0900192f //x=14.06 //y=2.08
c178 ( 40 0 ) capacitor c=0.110109f //x=12.21 //y=2.59
c179 ( 36 0 ) capacitor c=0.00398962f //x=11.81 //y=1.665
c180 ( 35 0 ) capacitor c=0.0137288f //x=12.125 //y=1.665
c181 ( 29 0 ) capacitor c=0.0284988f //x=12.125 //y=5.155
c182 ( 21 0 ) capacitor c=0.0176454f //x=11.345 //y=5.155
c183 ( 14 0 ) capacitor c=0.00332903f //x=9.755 //y=5.155
c184 ( 13 0 ) capacitor c=0.0148427f //x=10.465 //y=5.155
c185 ( 2 0 ) capacitor c=0.00879187f //x=12.325 //y=2.59
c186 ( 1 0 ) capacitor c=0.0476269f //x=13.945 //y=2.59
r187 (  75 77 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=13.96 //y=4.7 //x2=14.06 //y2=4.7
r188 (  68 77 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=14.4 //y=4.865 //x2=14.06 //y2=4.7
r189 (  67 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.395 //y=1.21 //x2=14.355 //y2=1.365
r190 (  66 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.395 //y=0.865 //x2=14.355 //y2=0.71
r191 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.395 //y=0.865 //x2=14.395 //y2=1.21
r192 (  64 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.02 //y=1.365 //x2=13.905 //y2=1.365
r193 (  63 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.24 //y=1.365 //x2=14.355 //y2=1.365
r194 (  62 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.02 //y=0.71 //x2=13.905 //y2=0.71
r195 (  61 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.24 //y=0.71 //x2=14.355 //y2=0.71
r196 (  61 62 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=14.24 //y=0.71 //x2=14.02 //y2=0.71
r197 (  58 75 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=13.96 //y=4.865 //x2=13.96 //y2=4.7
r198 (  57 72 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.915 //x2=14.06 //y2=2.08
r199 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.52 //x2=13.905 //y2=1.365
r200 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.52 //x2=13.865 //y2=1.915
r201 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.21 //x2=13.905 //y2=1.365
r202 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=0.865 //x2=13.905 //y2=0.71
r203 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.865 //y=0.865 //x2=13.865 //y2=1.21
r204 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.4 //y=6.02 //x2=14.4 //y2=4.865
r205 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.96 //y=6.02 //x2=13.96 //y2=4.865
r206 (  51 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.13 //y=1.365 //x2=14.24 //y2=1.365
r207 (  51 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.13 //y=1.365 //x2=14.02 //y2=1.365
r208 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=4.7 //x2=14.06 //y2=4.7
r209 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.59 //x2=14.06 //y2=4.7
r210 (  42 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=2.08 //x2=14.06 //y2=2.08
r211 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.08 //x2=14.06 //y2=2.59
r212 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=12.21 //y=5.07 //x2=12.21 //y2=2.59
r213 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.75 //x2=12.21 //y2=2.59
r214 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.665 //x2=12.21 //y2=1.75
r215 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.665 //x2=11.81 //y2=1.665
r216 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.725 //y=1.58 //x2=11.81 //y2=1.665
r217 (  31 80 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=11.725 //y=1.58 //x2=11.725 //y2=1.01
r218 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.515 //y=5.155 //x2=11.43 //y2=5.155
r219 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.155 //x2=12.21 //y2=5.07
r220 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.155 //x2=11.515 //y2=5.155
r221 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.43 //y=5.24 //x2=11.43 //y2=5.155
r222 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.43 //y=5.24 //x2=11.43 //y2=5.725
r223 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.635 //y=5.155 //x2=10.55 //y2=5.155
r224 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.345 //y=5.155 //x2=11.43 //y2=5.155
r225 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.345 //y=5.155 //x2=10.635 //y2=5.155
r226 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.55 //y=5.24 //x2=10.55 //y2=5.155
r227 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.55 //y=5.24 //x2=10.55 //y2=5.725
r228 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.465 //y=5.155 //x2=10.55 //y2=5.155
r229 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.465 //y=5.155 //x2=9.755 //y2=5.155
r230 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.67 //y=5.24 //x2=9.755 //y2=5.155
r231 (  7 82 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.67 //y=5.24 //x2=9.67 //y2=5.725
r232 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=2.59 //x2=14.06 //y2=2.59
r233 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.21 //y=2.59 //x2=12.21 //y2=2.59
r234 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.325 //y=2.59 //x2=12.21 //y2=2.59
r235 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=2.59 //x2=14.06 //y2=2.59
r236 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=13.945 //y=2.59 //x2=12.325 //y2=2.59
ends PM_DFFSNQX1\%noxref_4

subckt PM_DFFSNQX1\%CLK ( 1 2 7 8 9 10 11 12 13 14 16 26 28 37 38 39 40 41 42 \
 43 44 45 47 53 54 55 56 57 62 63 64 69 71 73 79 80 84 93 94 97 )
c198 ( 97 0 ) capacitor c=0.0331838f //x=14.83 //y=4.7
c199 ( 94 0 ) capacitor c=0.0279499f //x=14.8 //y=1.915
c200 ( 93 0 ) capacitor c=0.0425269f //x=14.8 //y=2.08
c201 ( 84 0 ) capacitor c=0.0334842f //x=5.55 //y=4.7
c202 ( 80 0 ) capacitor c=0.0429696f //x=15.365 //y=1.25
c203 ( 79 0 ) capacitor c=0.0192208f //x=15.365 //y=0.905
c204 ( 73 0 ) capacitor c=0.0148884f //x=15.21 //y=1.405
c205 ( 71 0 ) capacitor c=0.0157803f //x=15.21 //y=0.75
c206 ( 69 0 ) capacitor c=0.0299681f //x=15.205 //y=4.79
c207 ( 64 0 ) capacitor c=0.0205163f //x=14.835 //y=1.56
c208 ( 63 0 ) capacitor c=0.0168481f //x=14.835 //y=1.25
c209 ( 62 0 ) capacitor c=0.0174783f //x=14.835 //y=0.905
c210 ( 57 0 ) capacitor c=0.0245352f //x=5.885 //y=4.79
c211 ( 56 0 ) capacitor c=0.0826403f //x=5.64 //y=1.915
c212 ( 55 0 ) capacitor c=0.0170266f //x=5.64 //y=1.45
c213 ( 54 0 ) capacitor c=0.018609f //x=5.64 //y=1.22
c214 ( 53 0 ) capacitor c=0.0187309f //x=5.64 //y=0.91
c215 ( 47 0 ) capacitor c=0.014725f //x=5.485 //y=1.375
c216 ( 45 0 ) capacitor c=0.0146567f //x=5.485 //y=0.755
c217 ( 44 0 ) capacitor c=0.0335408f //x=5.115 //y=1.22
c218 ( 43 0 ) capacitor c=0.0173761f //x=5.115 //y=0.91
c219 ( 42 0 ) capacitor c=0.15358f //x=15.28 //y=6.02
c220 ( 41 0 ) capacitor c=0.110281f //x=14.84 //y=6.02
c221 ( 40 0 ) capacitor c=0.110114f //x=5.96 //y=6.02
c222 ( 39 0 ) capacitor c=0.11012f //x=5.52 //y=6.02
c223 ( 28 0 ) capacitor c=0.0726007f //x=14.8 //y=2.08
c224 ( 26 0 ) capacitor c=0.00369614f //x=14.8 //y=4.535
c225 ( 16 0 ) capacitor c=0.0979973f //x=5.55 //y=2.08
c226 ( 2 0 ) capacitor c=0.0154455f //x=5.665 //y=4.44
c227 ( 1 0 ) capacitor c=0.21665f //x=14.685 //y=4.44
r228 (  99 100 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=14.83 //y=4.79 //x2=14.83 //y2=4.865
r229 (  97 99 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=14.83 //y=4.7 //x2=14.83 //y2=4.79
r230 (  93 94 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=14.8 //y=2.08 //x2=14.8 //y2=1.915
r231 (  86 87 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=5.55 //y=4.79 //x2=5.55 //y2=4.865
r232 (  84 86 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=5.55 //y=4.7 //x2=5.55 //y2=4.79
r233 (  80 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.365 //y=1.25 //x2=15.325 //y2=1.405
r234 (  79 103 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.365 //y=0.905 //x2=15.325 //y2=0.75
r235 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.365 //y=0.905 //x2=15.365 //y2=1.25
r236 (  74 102 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.99 //y=1.405 //x2=14.875 //y2=1.405
r237 (  73 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.21 //y=1.405 //x2=15.325 //y2=1.405
r238 (  72 101 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.99 //y=0.75 //x2=14.875 //y2=0.75
r239 (  71 103 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.21 //y=0.75 //x2=15.325 //y2=0.75
r240 (  71 72 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.21 //y=0.75 //x2=14.99 //y2=0.75
r241 (  70 99 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=14.965 //y=4.79 //x2=14.83 //y2=4.79
r242 (  69 76 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.79 //x2=15.28 //y2=4.865
r243 (  69 70 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.79 //x2=14.965 //y2=4.79
r244 (  64 102 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.56 //x2=14.875 //y2=1.405
r245 (  64 94 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.56 //x2=14.835 //y2=1.915
r246 (  63 102 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.25 //x2=14.875 //y2=1.405
r247 (  62 101 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=0.905 //x2=14.875 //y2=0.75
r248 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.835 //y=0.905 //x2=14.835 //y2=1.25
r249 (  58 86 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=5.685 //y=4.79 //x2=5.55 //y2=4.79
r250 (  57 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.885 //y=4.79 //x2=5.96 //y2=4.865
r251 (  57 58 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=5.885 //y=4.79 //x2=5.685 //y2=4.79
r252 (  56 91 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.915 //x2=5.565 //y2=2.08
r253 (  55 89 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.45 //x2=5.6 //y2=1.375
r254 (  55 56 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.45 //x2=5.64 //y2=1.915
r255 (  54 89 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.22 //x2=5.6 //y2=1.375
r256 (  53 88 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.64 //y=0.91 //x2=5.6 //y2=0.755
r257 (  53 54 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=5.64 //y=0.91 //x2=5.64 //y2=1.22
r258 (  48 82 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.27 //y=1.375 //x2=5.155 //y2=1.375
r259 (  47 89 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.485 //y=1.375 //x2=5.6 //y2=1.375
r260 (  46 81 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.27 //y=0.755 //x2=5.155 //y2=0.755
r261 (  45 88 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.485 //y=0.755 //x2=5.6 //y2=0.755
r262 (  45 46 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=5.485 //y=0.755 //x2=5.27 //y2=0.755
r263 (  44 82 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.115 //y=1.22 //x2=5.155 //y2=1.375
r264 (  43 81 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.115 //y=0.91 //x2=5.155 //y2=0.755
r265 (  43 44 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=5.115 //y=0.91 //x2=5.115 //y2=1.22
r266 (  42 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.28 //y=6.02 //x2=15.28 //y2=4.865
r267 (  41 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.84 //y=6.02 //x2=14.84 //y2=4.865
r268 (  40 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.96 //y=6.02 //x2=5.96 //y2=4.865
r269 (  39 87 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.52 //y=6.02 //x2=5.52 //y2=4.865
r270 (  38 73 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.1 //y=1.405 //x2=15.21 //y2=1.405
r271 (  38 74 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.1 //y=1.405 //x2=14.99 //y2=1.405
r272 (  37 47 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=5.377 //y=1.375 //x2=5.485 //y2=1.375
r273 (  37 48 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=5.377 //y=1.375 //x2=5.27 //y2=1.375
r274 (  36 97 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.83 //y=4.7 //x2=14.83 //y2=4.7
r275 (  28 93 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.8 //y=2.08 //x2=14.8 //y2=2.08
r276 (  26 36 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=14.8 //y=4.535 //x2=14.815 //y2=4.7
r277 (  24 84 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=4.7 //x2=5.55 //y2=4.7
r278 (  16 91 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=2.08 //x2=5.55 //y2=2.08
r279 (  14 26 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=14.8 //y=4.44 //x2=14.8 //y2=4.535
r280 (  13 14 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=14.8 //y=3.33 //x2=14.8 //y2=4.44
r281 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=14.8 //y=2.96 //x2=14.8 //y2=3.33
r282 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=14.8 //y=2.59 //x2=14.8 //y2=2.96
r283 (  11 28 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=14.8 //y=2.59 //x2=14.8 //y2=2.08
r284 (  10 24 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=5.55 //y=4.44 //x2=5.55 //y2=4.7
r285 (  9 10 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=5.55 //y=3.7 //x2=5.55 //y2=4.44
r286 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=5.55 //y=3.33 //x2=5.55 //y2=3.7
r287 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=5.55 //y=2.96 //x2=5.55 //y2=3.33
r288 (  7 16 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=5.55 //y=2.96 //x2=5.55 //y2=2.08
r289 (  6 14 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.8 //y=4.44 //x2=14.8 //y2=4.44
r290 (  4 10 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.55 //y=4.44 //x2=5.55 //y2=4.44
r291 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.665 //y=4.44 //x2=5.55 //y2=4.44
r292 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.685 //y=4.44 //x2=14.8 //y2=4.44
r293 (  1 2 ) resistor r=8.60687 //w=0.131 //l=9.02 //layer=m1 \
 //thickness=0.36 //x=14.685 //y=4.44 //x2=5.665 //y2=4.44
ends PM_DFFSNQX1\%CLK

subckt PM_DFFSNQX1\%noxref_6 ( 1 2 3 4 11 13 23 24 31 39 45 46 50 52 61 62 64 \
 65 67 68 69 70 71 72 73 74 75 80 82 84 90 91 92 93 94 95 99 101 104 105 110 \
 111 114 128 131 133 134 135 )
c286 ( 135 0 ) capacitor c=0.023087f //x=6.475 //y=5.02
c287 ( 134 0 ) capacitor c=0.023519f //x=5.595 //y=5.02
c288 ( 133 0 ) capacitor c=0.0224735f //x=4.715 //y=5.02
c289 ( 131 0 ) capacitor c=0.00853354f //x=6.725 //y=0.915
c290 ( 128 0 ) capacitor c=0.0597793f //x=17.39 //y=4.7
c291 ( 114 0 ) capacitor c=0.0331534f //x=1.88 //y=4.7
c292 ( 111 0 ) capacitor c=0.0279499f //x=1.85 //y=1.915
c293 ( 110 0 ) capacitor c=0.0437302f //x=1.85 //y=2.08
c294 ( 105 0 ) capacitor c=0.0318948f //x=17.725 //y=1.21
c295 ( 104 0 ) capacitor c=0.0187384f //x=17.725 //y=0.865
c296 ( 101 0 ) capacitor c=0.0141798f //x=17.57 //y=1.365
c297 ( 99 0 ) capacitor c=0.0149844f //x=17.57 //y=0.71
c298 ( 95 0 ) capacitor c=0.0813322f //x=17.195 //y=1.915
c299 ( 94 0 ) capacitor c=0.0229267f //x=17.195 //y=1.52
c300 ( 93 0 ) capacitor c=0.0234352f //x=17.195 //y=1.21
c301 ( 92 0 ) capacitor c=0.0199343f //x=17.195 //y=0.865
c302 ( 91 0 ) capacitor c=0.0429696f //x=2.415 //y=1.25
c303 ( 90 0 ) capacitor c=0.0192208f //x=2.415 //y=0.905
c304 ( 84 0 ) capacitor c=0.0158629f //x=2.26 //y=1.405
c305 ( 82 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c306 ( 80 0 ) capacitor c=0.0299681f //x=2.255 //y=4.79
c307 ( 75 0 ) capacitor c=0.0205163f //x=1.885 //y=1.56
c308 ( 74 0 ) capacitor c=0.0168481f //x=1.885 //y=1.25
c309 ( 73 0 ) capacitor c=0.0174783f //x=1.885 //y=0.905
c310 ( 72 0 ) capacitor c=0.110275f //x=17.73 //y=6.02
c311 ( 71 0 ) capacitor c=0.154305f //x=17.29 //y=6.02
c312 ( 70 0 ) capacitor c=0.15358f //x=2.33 //y=6.02
c313 ( 69 0 ) capacitor c=0.110281f //x=1.89 //y=6.02
c314 ( 65 0 ) capacitor c=0.0786338f //x=7.397 //y=3.905
c315 ( 64 0 ) capacitor c=0.0101843f //x=7.395 //y=4.07
c316 ( 62 0 ) capacitor c=0.00106608f //x=6.62 //y=5.155
c317 ( 61 0 ) capacitor c=0.00207162f //x=5.74 //y=5.155
c318 ( 52 0 ) capacitor c=0.0929759f //x=17.39 //y=2.08
c319 ( 50 0 ) capacitor c=0.0236247f //x=7.4 //y=5.07
c320 ( 46 0 ) capacitor c=0.00431225f //x=7 //y=1.665
c321 ( 45 0 ) capacitor c=0.0141453f //x=7.315 //y=1.665
c322 ( 39 0 ) capacitor c=0.0281378f //x=7.315 //y=5.155
c323 ( 31 0 ) capacitor c=0.0176454f //x=6.535 //y=5.155
c324 ( 24 0 ) capacitor c=0.00351598f //x=4.945 //y=5.155
c325 ( 23 0 ) capacitor c=0.0154196f //x=5.655 //y=5.155
c326 ( 13 0 ) capacitor c=0.0787953f //x=1.85 //y=2.08
c327 ( 11 0 ) capacitor c=0.00453889f //x=1.85 //y=4.535
c328 ( 4 0 ) capacitor c=0.00551102f //x=7.51 //y=4.07
c329 ( 3 0 ) capacitor c=0.180782f //x=17.275 //y=4.07
c330 ( 2 0 ) capacitor c=0.0180257f //x=1.965 //y=4.07
c331 ( 1 0 ) capacitor c=0.159166f //x=7.28 //y=4.07
r332 (  126 128 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=17.29 //y=4.7 //x2=17.39 //y2=4.7
r333 (  116 117 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.79 //x2=1.88 //y2=4.865
r334 (  114 116 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.7 //x2=1.88 //y2=4.79
r335 (  110 111 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r336 (  106 128 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=17.73 //y=4.865 //x2=17.39 //y2=4.7
r337 (  105 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.725 //y=1.21 //x2=17.685 //y2=1.365
r338 (  104 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.725 //y=0.865 //x2=17.685 //y2=0.71
r339 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.725 //y=0.865 //x2=17.725 //y2=1.21
r340 (  102 125 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.35 //y=1.365 //x2=17.235 //y2=1.365
r341 (  101 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.57 //y=1.365 //x2=17.685 //y2=1.365
r342 (  100 124 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.35 //y=0.71 //x2=17.235 //y2=0.71
r343 (  99 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.57 //y=0.71 //x2=17.685 //y2=0.71
r344 (  99 100 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.57 //y=0.71 //x2=17.35 //y2=0.71
r345 (  96 126 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.29 //y=4.865 //x2=17.29 //y2=4.7
r346 (  95 123 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.915 //x2=17.39 //y2=2.08
r347 (  94 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.52 //x2=17.235 //y2=1.365
r348 (  94 95 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.52 //x2=17.195 //y2=1.915
r349 (  93 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.21 //x2=17.235 //y2=1.365
r350 (  92 124 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=0.865 //x2=17.235 //y2=0.71
r351 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.195 //y=0.865 //x2=17.195 //y2=1.21
r352 (  91 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r353 (  90 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r354 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r355 (  85 119 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r356 (  84 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r357 (  83 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r358 (  82 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r359 (  82 83 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r360 (  81 116 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.015 //y=4.79 //x2=1.88 //y2=4.79
r361 (  80 87 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.33 //y2=4.865
r362 (  80 81 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.015 //y2=4.79
r363 (  75 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r364 (  75 111 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r365 (  74 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r366 (  73 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r367 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r368 (  72 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.73 //y=6.02 //x2=17.73 //y2=4.865
r369 (  71 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.29 //y=6.02 //x2=17.29 //y2=4.865
r370 (  70 87 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.02 //x2=2.33 //y2=4.865
r371 (  69 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.02 //x2=1.89 //y2=4.865
r372 (  68 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.46 //y=1.365 //x2=17.57 //y2=1.365
r373 (  68 102 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.46 //y=1.365 //x2=17.35 //y2=1.365
r374 (  67 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r375 (  67 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r376 (  64 66 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=7.397 //y=4.07 //x2=7.397 //y2=4.235
r377 (  64 65 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=7.397 //y=4.07 //x2=7.397 //y2=3.905
r378 (  60 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.88 //y=4.7 //x2=1.88 //y2=4.7
r379 (  57 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.39 //y=4.7 //x2=17.39 //y2=4.7
r380 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=17.39 //y=4.07 //x2=17.39 //y2=4.7
r381 (  52 123 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.39 //y=2.08 //x2=17.39 //y2=2.08
r382 (  52 55 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=17.39 //y=2.08 //x2=17.39 //y2=4.07
r383 (  50 66 ) resistor r=57.1551 //w=0.187 //l=0.835 //layer=li \
 //thickness=0.1 //x=7.4 //y=5.07 //x2=7.4 //y2=4.235
r384 (  47 65 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=7.4 //y=1.75 //x2=7.4 //y2=3.905
r385 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.665 //x2=7.4 //y2=1.75
r386 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.665 //x2=7 //y2=1.665
r387 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.915 //y=1.58 //x2=7 //y2=1.665
r388 (  41 131 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=6.915 //y=1.58 //x2=6.915 //y2=1.01
r389 (  40 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.705 //y=5.155 //x2=6.62 //y2=5.155
r390 (  39 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.155 //x2=7.4 //y2=5.07
r391 (  39 40 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.155 //x2=6.705 //y2=5.155
r392 (  33 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.62 //y=5.24 //x2=6.62 //y2=5.155
r393 (  33 135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.62 //y=5.24 //x2=6.62 //y2=5.725
r394 (  32 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.825 //y=5.155 //x2=5.74 //y2=5.155
r395 (  31 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.535 //y=5.155 //x2=6.62 //y2=5.155
r396 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.535 //y=5.155 //x2=5.825 //y2=5.155
r397 (  25 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.74 //y=5.24 //x2=5.74 //y2=5.155
r398 (  25 134 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=5.74 //y=5.24 //x2=5.74 //y2=5.725
r399 (  23 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.655 //y=5.155 //x2=5.74 //y2=5.155
r400 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.655 //y=5.155 //x2=4.945 //y2=5.155
r401 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.86 //y=5.24 //x2=4.945 //y2=5.155
r402 (  17 133 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.86 //y=5.24 //x2=4.86 //y2=5.725
r403 (  13 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r404 (  13 16 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.08 //x2=1.85 //y2=4.07
r405 (  11 60 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.865 //y2=4.7
r406 (  11 16 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.85 //y2=4.07
r407 (  10 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.39 //y=4.07 //x2=17.39 //y2=4.07
r408 (  8 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.395 //y=4.07 //x2=7.395 //y2=4.07
r409 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.85 //y=4.07 //x2=1.85 //y2=4.07
r410 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.51 //y=4.07 //x2=7.395 //y2=4.07
r411 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.275 //y=4.07 //x2=17.39 //y2=4.07
r412 (  3 4 ) resistor r=9.31775 //w=0.131 //l=9.765 //layer=m1 \
 //thickness=0.36 //x=17.275 //y=4.07 //x2=7.51 //y2=4.07
r413 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.965 //y=4.07 //x2=1.85 //y2=4.07
r414 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.28 //y=4.07 //x2=7.395 //y2=4.07
r415 (  1 2 ) resistor r=5.07156 //w=0.131 //l=5.315 //layer=m1 \
 //thickness=0.36 //x=7.28 //y=4.07 //x2=1.965 //y2=4.07
ends PM_DFFSNQX1\%noxref_6

subckt PM_DFFSNQX1\%noxref_7 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 \
 48 49 51 57 58 59 60 72 74 75 )
c145 ( 75 0 ) capacitor c=0.0220291f //x=18.245 //y=5.02
c146 ( 74 0 ) capacitor c=0.0217503f //x=17.365 //y=5.02
c147 ( 72 0 ) capacitor c=0.0084702f //x=18.24 //y=0.905
c148 ( 60 0 ) capacitor c=0.0562318f //x=20.995 //y=4.79
c149 ( 59 0 ) capacitor c=0.0305765f //x=21.285 //y=4.79
c150 ( 58 0 ) capacitor c=0.0347816f //x=20.95 //y=1.22
c151 ( 57 0 ) capacitor c=0.0187487f //x=20.95 //y=0.875
c152 ( 51 0 ) capacitor c=0.0137055f //x=20.795 //y=1.375
c153 ( 49 0 ) capacitor c=0.0149861f //x=20.795 //y=0.72
c154 ( 48 0 ) capacitor c=0.096037f //x=20.42 //y=1.915
c155 ( 47 0 ) capacitor c=0.0228993f //x=20.42 //y=1.53
c156 ( 46 0 ) capacitor c=0.0234352f //x=20.42 //y=1.22
c157 ( 45 0 ) capacitor c=0.0198724f //x=20.42 //y=0.875
c158 ( 44 0 ) capacitor c=0.110114f //x=21.36 //y=6.02
c159 ( 43 0 ) capacitor c=0.158956f //x=20.92 //y=6.02
c160 ( 41 0 ) capacitor c=0.0024826f //x=18.39 //y=5.2
c161 ( 34 0 ) capacitor c=0.101911f //x=20.72 //y=2.08
c162 ( 32 0 ) capacitor c=0.108434f //x=18.87 //y=2.96
c163 ( 28 0 ) capacitor c=0.00404073f //x=18.515 //y=1.655
c164 ( 27 0 ) capacitor c=0.0122201f //x=18.785 //y=1.655
c165 ( 25 0 ) capacitor c=0.0143719f //x=18.785 //y=5.2
c166 ( 14 0 ) capacitor c=0.00272496f //x=17.595 //y=5.2
c167 ( 13 0 ) capacitor c=0.0155386f //x=18.305 //y=5.2
c168 ( 2 0 ) capacitor c=0.0123518f //x=18.985 //y=2.96
c169 ( 1 0 ) capacitor c=0.0446552f //x=20.605 //y=2.96
r170 (  59 61 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.285 //y=4.79 //x2=21.36 //y2=4.865
r171 (  59 60 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=21.285 //y=4.79 //x2=20.995 //y2=4.79
r172 (  58 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.95 //y=1.22 //x2=20.91 //y2=1.375
r173 (  57 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.95 //y=0.875 //x2=20.91 //y2=0.72
r174 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.95 //y=0.875 //x2=20.95 //y2=1.22
r175 (  54 60 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.92 //y=4.865 //x2=20.995 //y2=4.79
r176 (  54 69 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=20.92 //y=4.865 //x2=20.72 //y2=4.7
r177 (  52 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.575 //y=1.375 //x2=20.46 //y2=1.375
r178 (  51 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.795 //y=1.375 //x2=20.91 //y2=1.375
r179 (  50 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.575 //y=0.72 //x2=20.46 //y2=0.72
r180 (  49 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.795 //y=0.72 //x2=20.91 //y2=0.72
r181 (  49 50 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.795 //y=0.72 //x2=20.575 //y2=0.72
r182 (  48 67 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.915 //x2=20.72 //y2=2.08
r183 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.53 //x2=20.46 //y2=1.375
r184 (  47 48 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.53 //x2=20.42 //y2=1.915
r185 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.22 //x2=20.46 //y2=1.375
r186 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=0.875 //x2=20.46 //y2=0.72
r187 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.42 //y=0.875 //x2=20.42 //y2=1.22
r188 (  44 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.36 //y=6.02 //x2=21.36 //y2=4.865
r189 (  43 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.92 //y=6.02 //x2=20.92 //y2=4.865
r190 (  42 51 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.685 //y=1.375 //x2=20.795 //y2=1.375
r191 (  42 52 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.685 //y=1.375 //x2=20.575 //y2=1.375
r192 (  39 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.72 //y=4.7 //x2=20.72 //y2=4.7
r193 (  37 39 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.96 //x2=20.72 //y2=4.7
r194 (  34 67 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.72 //y=2.08 //x2=20.72 //y2=2.08
r195 (  34 37 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.08 //x2=20.72 //y2=2.96
r196 (  30 32 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=18.87 //y=5.115 //x2=18.87 //y2=2.96
r197 (  29 32 ) resistor r=83.508 //w=0.187 //l=1.22 //layer=li \
 //thickness=0.1 //x=18.87 //y=1.74 //x2=18.87 //y2=2.96
r198 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.785 //y=1.655 //x2=18.87 //y2=1.74
r199 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=18.785 //y=1.655 //x2=18.515 //y2=1.655
r200 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.475 //y=5.2 //x2=18.39 //y2=5.2
r201 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.785 //y=5.2 //x2=18.87 //y2=5.115
r202 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=18.785 //y=5.2 //x2=18.475 //y2=5.2
r203 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.43 //y=1.57 //x2=18.515 //y2=1.655
r204 (  21 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=18.43 //y=1.57 //x2=18.43 //y2=1
r205 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.39 //y=5.285 //x2=18.39 //y2=5.2
r206 (  15 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=18.39 //y=5.285 //x2=18.39 //y2=5.725
r207 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.305 //y=5.2 //x2=18.39 //y2=5.2
r208 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=18.305 //y=5.2 //x2=17.595 //y2=5.2
r209 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.51 //y=5.285 //x2=17.595 //y2=5.2
r210 (  7 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=17.51 //y=5.285 //x2=17.51 //y2=5.725
r211 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.72 //y=2.96 //x2=20.72 //y2=2.96
r212 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.87 //y=2.96 //x2=18.87 //y2=2.96
r213 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.985 //y=2.96 //x2=18.87 //y2=2.96
r214 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=2.96 //x2=20.72 //y2=2.96
r215 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=20.605 //y=2.96 //x2=18.985 //y2=2.96
ends PM_DFFSNQX1\%noxref_7

subckt PM_DFFSNQX1\%SN ( 1 2 7 8 9 10 11 12 13 14 15 17 28 39 40 41 42 43 44 \
 45 46 47 49 55 56 57 58 59 64 65 66 68 74 75 76 77 78 86 97 )
c226 ( 97 0 ) capacitor c=0.0337728f //x=21.83 //y=4.7
c227 ( 86 0 ) capacitor c=0.0335551f //x=10.36 //y=4.7
c228 ( 78 0 ) capacitor c=0.025532f //x=22.165 //y=4.79
c229 ( 77 0 ) capacitor c=0.0831166f //x=21.92 //y=1.915
c230 ( 76 0 ) capacitor c=0.0170266f //x=21.92 //y=1.45
c231 ( 75 0 ) capacitor c=0.018609f //x=21.92 //y=1.22
c232 ( 74 0 ) capacitor c=0.0187309f //x=21.92 //y=0.91
c233 ( 68 0 ) capacitor c=0.014725f //x=21.765 //y=1.375
c234 ( 66 0 ) capacitor c=0.0146567f //x=21.765 //y=0.755
c235 ( 65 0 ) capacitor c=0.0335408f //x=21.395 //y=1.22
c236 ( 64 0 ) capacitor c=0.0173761f //x=21.395 //y=0.91
c237 ( 59 0 ) capacitor c=0.0245352f //x=10.695 //y=4.79
c238 ( 58 0 ) capacitor c=0.0826756f //x=10.45 //y=1.915
c239 ( 57 0 ) capacitor c=0.0170266f //x=10.45 //y=1.45
c240 ( 56 0 ) capacitor c=0.018609f //x=10.45 //y=1.22
c241 ( 55 0 ) capacitor c=0.0187309f //x=10.45 //y=0.91
c242 ( 49 0 ) capacitor c=0.014725f //x=10.295 //y=1.375
c243 ( 47 0 ) capacitor c=0.0146567f //x=10.295 //y=0.755
c244 ( 46 0 ) capacitor c=0.0335408f //x=9.925 //y=1.22
c245 ( 45 0 ) capacitor c=0.0173761f //x=9.925 //y=0.91
c246 ( 44 0 ) capacitor c=0.110114f //x=22.24 //y=6.02
c247 ( 43 0 ) capacitor c=0.11012f //x=21.8 //y=6.02
c248 ( 42 0 ) capacitor c=0.110114f //x=10.77 //y=6.02
c249 ( 41 0 ) capacitor c=0.11012f //x=10.33 //y=6.02
c250 ( 28 0 ) capacitor c=0.0978105f //x=21.83 //y=2.08
c251 ( 17 0 ) capacitor c=0.094794f //x=10.36 //y=2.08
c252 ( 2 0 ) capacitor c=0.0160685f //x=10.475 //y=2.22
c253 ( 1 0 ) capacitor c=0.295394f //x=21.715 //y=2.22
r254 (  99 100 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=21.83 //y=4.79 //x2=21.83 //y2=4.865
r255 (  97 99 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=21.83 //y=4.7 //x2=21.83 //y2=4.79
r256 (  88 89 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=10.36 //y=4.79 //x2=10.36 //y2=4.865
r257 (  86 88 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=10.36 //y=4.7 //x2=10.36 //y2=4.79
r258 (  79 99 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=21.965 //y=4.79 //x2=21.83 //y2=4.79
r259 (  78 80 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=22.165 //y=4.79 //x2=22.24 //y2=4.865
r260 (  78 79 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=22.165 //y=4.79 //x2=21.965 //y2=4.79
r261 (  77 104 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.915 //x2=21.845 //y2=2.08
r262 (  76 102 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.45 //x2=21.88 //y2=1.375
r263 (  76 77 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.45 //x2=21.92 //y2=1.915
r264 (  75 102 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.22 //x2=21.88 //y2=1.375
r265 (  74 101 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.92 //y=0.91 //x2=21.88 //y2=0.755
r266 (  74 75 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.92 //y=0.91 //x2=21.92 //y2=1.22
r267 (  69 95 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.375 //x2=21.435 //y2=1.375
r268 (  68 102 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.765 //y=1.375 //x2=21.88 //y2=1.375
r269 (  67 94 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.755 //x2=21.435 //y2=0.755
r270 (  66 101 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.765 //y=0.755 //x2=21.88 //y2=0.755
r271 (  66 67 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=21.765 //y=0.755 //x2=21.55 //y2=0.755
r272 (  65 95 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.395 //y=1.22 //x2=21.435 //y2=1.375
r273 (  64 94 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.91 //x2=21.435 //y2=0.755
r274 (  64 65 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.91 //x2=21.395 //y2=1.22
r275 (  60 88 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=10.495 //y=4.79 //x2=10.36 //y2=4.79
r276 (  59 61 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.695 //y=4.79 //x2=10.77 //y2=4.865
r277 (  59 60 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=10.695 //y=4.79 //x2=10.495 //y2=4.79
r278 (  58 93 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.915 //x2=10.375 //y2=2.08
r279 (  57 91 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.45 //x2=10.41 //y2=1.375
r280 (  57 58 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.45 //x2=10.45 //y2=1.915
r281 (  56 91 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.22 //x2=10.41 //y2=1.375
r282 (  55 90 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.45 //y=0.91 //x2=10.41 //y2=0.755
r283 (  55 56 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=10.45 //y=0.91 //x2=10.45 //y2=1.22
r284 (  50 84 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.08 //y=1.375 //x2=9.965 //y2=1.375
r285 (  49 91 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.295 //y=1.375 //x2=10.41 //y2=1.375
r286 (  48 83 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.08 //y=0.755 //x2=9.965 //y2=0.755
r287 (  47 90 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.295 //y=0.755 //x2=10.41 //y2=0.755
r288 (  47 48 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=10.295 //y=0.755 //x2=10.08 //y2=0.755
r289 (  46 84 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.925 //y=1.22 //x2=9.965 //y2=1.375
r290 (  45 83 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.925 //y=0.91 //x2=9.965 //y2=0.755
r291 (  45 46 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=9.925 //y=0.91 //x2=9.925 //y2=1.22
r292 (  44 80 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.24 //y=6.02 //x2=22.24 //y2=4.865
r293 (  43 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.8 //y=6.02 //x2=21.8 //y2=4.865
r294 (  42 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.77 //y=6.02 //x2=10.77 //y2=4.865
r295 (  41 89 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.33 //y=6.02 //x2=10.33 //y2=4.865
r296 (  40 68 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=21.657 //y=1.375 //x2=21.765 //y2=1.375
r297 (  40 69 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=21.657 //y=1.375 //x2=21.55 //y2=1.375
r298 (  39 49 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=10.187 //y=1.375 //x2=10.295 //y2=1.375
r299 (  39 50 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=10.187 //y=1.375 //x2=10.08 //y2=1.375
r300 (  37 97 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.83 //y=4.7 //x2=21.83 //y2=4.7
r301 (  28 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.83 //y=2.08 //x2=21.83 //y2=2.08
r302 (  25 86 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=4.7 //x2=10.36 //y2=4.7
r303 (  17 93 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=2.08 //x2=10.36 //y2=2.08
r304 (  15 37 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=21.83 //y=4.44 //x2=21.83 //y2=4.7
r305 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.83 //y=4.07 //x2=21.83 //y2=4.44
r306 (  13 14 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.96 //x2=21.83 //y2=4.07
r307 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.59 //x2=21.83 //y2=2.96
r308 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.22 //x2=21.83 //y2=2.59
r309 (  11 28 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.22 //x2=21.83 //y2=2.08
r310 (  10 25 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=10.36 //y=3.33 //x2=10.36 //y2=4.7
r311 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.96 //x2=10.36 //y2=3.33
r312 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=10.36 //y=2.59 //x2=10.36 //y2=2.96
r313 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=10.36 //y=2.22 //x2=10.36 //y2=2.59
r314 (  7 17 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.22 //x2=10.36 //y2=2.08
r315 (  6 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.83 //y=2.22 //x2=21.83 //y2=2.22
r316 (  4 7 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=2.22 //x2=10.36 //y2=2.22
r317 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.475 //y=2.22 //x2=10.36 //y2=2.22
r318 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=2.22 //x2=21.83 //y2=2.22
r319 (  1 2 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=2.22 //x2=10.475 //y2=2.22
ends PM_DFFSNQX1\%SN

subckt PM_DFFSNQX1\%noxref_9 ( 1 2 3 4 5 6 16 24 37 38 49 51 52 56 58 65 66 67 \
 68 69 70 71 72 73 74 78 79 80 85 87 90 91 95 96 97 102 104 107 108 112 113 \
 114 119 121 124 125 127 128 133 137 138 143 147 148 153 156 158 159 )
c324 ( 159 0 ) capacitor c=0.0220291f //x=14.915 //y=5.02
c325 ( 158 0 ) capacitor c=0.0217503f //x=14.035 //y=5.02
c326 ( 156 0 ) capacitor c=0.00866655f //x=14.91 //y=0.905
c327 ( 153 0 ) capacitor c=0.0617593f //x=22.94 //y=4.7
c328 ( 148 0 ) capacitor c=0.0273931f //x=22.94 //y=1.915
c329 ( 147 0 ) capacitor c=0.0471168f //x=22.94 //y=2.08
c330 ( 143 0 ) capacitor c=0.0587755f //x=11.47 //y=4.7
c331 ( 138 0 ) capacitor c=0.0273931f //x=11.47 //y=1.915
c332 ( 137 0 ) capacitor c=0.0462455f //x=11.47 //y=2.08
c333 ( 133 0 ) capacitor c=0.058931f //x=6.66 //y=4.7
c334 ( 128 0 ) capacitor c=0.0267105f //x=6.66 //y=1.915
c335 ( 127 0 ) capacitor c=0.0457054f //x=6.66 //y=2.08
c336 ( 125 0 ) capacitor c=0.0432517f //x=23.46 //y=1.26
c337 ( 124 0 ) capacitor c=0.0200379f //x=23.46 //y=0.915
c338 ( 121 0 ) capacitor c=0.0158629f //x=23.305 //y=1.415
c339 ( 119 0 ) capacitor c=0.0157803f //x=23.305 //y=0.76
c340 ( 114 0 ) capacitor c=0.0218028f //x=22.93 //y=1.57
c341 ( 113 0 ) capacitor c=0.0207459f //x=22.93 //y=1.26
c342 ( 112 0 ) capacitor c=0.0194308f //x=22.93 //y=0.915
c343 ( 108 0 ) capacitor c=0.0432517f //x=11.99 //y=1.26
c344 ( 107 0 ) capacitor c=0.0200379f //x=11.99 //y=0.915
c345 ( 104 0 ) capacitor c=0.0148873f //x=11.835 //y=1.415
c346 ( 102 0 ) capacitor c=0.0157803f //x=11.835 //y=0.76
c347 ( 97 0 ) capacitor c=0.0218028f //x=11.46 //y=1.57
c348 ( 96 0 ) capacitor c=0.0207459f //x=11.46 //y=1.26
c349 ( 95 0 ) capacitor c=0.0194308f //x=11.46 //y=0.915
c350 ( 91 0 ) capacitor c=0.0432517f //x=7.18 //y=1.26
c351 ( 90 0 ) capacitor c=0.0200379f //x=7.18 //y=0.915
c352 ( 87 0 ) capacitor c=0.0158629f //x=7.025 //y=1.415
c353 ( 85 0 ) capacitor c=0.0157803f //x=7.025 //y=0.76
c354 ( 80 0 ) capacitor c=0.0218028f //x=6.65 //y=1.57
c355 ( 79 0 ) capacitor c=0.0207459f //x=6.65 //y=1.26
c356 ( 78 0 ) capacitor c=0.0194308f //x=6.65 //y=0.915
c357 ( 74 0 ) capacitor c=0.158794f //x=23.12 //y=6.02
c358 ( 73 0 ) capacitor c=0.110114f //x=22.68 //y=6.02
c359 ( 72 0 ) capacitor c=0.158794f //x=11.65 //y=6.02
c360 ( 71 0 ) capacitor c=0.110114f //x=11.21 //y=6.02
c361 ( 70 0 ) capacitor c=0.158048f //x=6.84 //y=6.02
c362 ( 69 0 ) capacitor c=0.110114f //x=6.4 //y=6.02
c363 ( 65 0 ) capacitor c=0.0023043f //x=15.06 //y=5.2
c364 ( 58 0 ) capacitor c=0.0908639f //x=22.94 //y=2.08
c365 ( 56 0 ) capacitor c=0.110723f //x=15.54 //y=3.7
c366 ( 52 0 ) capacitor c=0.00404073f //x=15.185 //y=1.655
c367 ( 51 0 ) capacitor c=0.0122201f //x=15.455 //y=1.655
c368 ( 49 0 ) capacitor c=0.0140462f //x=15.455 //y=5.2
c369 ( 38 0 ) capacitor c=0.00251635f //x=14.265 //y=5.2
c370 ( 37 0 ) capacitor c=0.0143111f //x=14.975 //y=5.2
c371 ( 24 0 ) capacitor c=0.0857928f //x=11.47 //y=2.08
c372 ( 16 0 ) capacitor c=0.0865938f //x=6.66 //y=2.08
c373 ( 6 0 ) capacitor c=0.00472158f //x=15.655 //y=3.7
c374 ( 5 0 ) capacitor c=0.215022f //x=22.825 //y=3.7
c375 ( 4 0 ) capacitor c=0.00493991f //x=11.585 //y=3.7
c376 ( 3 0 ) capacitor c=0.0805272f //x=15.425 //y=3.7
c377 ( 2 0 ) capacitor c=0.0147097f //x=6.775 //y=3.7
c378 ( 1 0 ) capacitor c=0.105064f //x=11.355 //y=3.7
r379 (  147 148 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=22.94 //y=2.08 //x2=22.94 //y2=1.915
r380 (  137 138 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11.47 //y=2.08 //x2=11.47 //y2=1.915
r381 (  127 128 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.66 //y=2.08 //x2=6.66 //y2=1.915
r382 (  125 155 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.46 //y=1.26 //x2=23.42 //y2=1.415
r383 (  124 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.46 //y=0.915 //x2=23.42 //y2=0.76
r384 (  124 125 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.46 //y=0.915 //x2=23.46 //y2=1.26
r385 (  122 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.085 //y=1.415 //x2=22.97 //y2=1.415
r386 (  121 155 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.305 //y=1.415 //x2=23.42 //y2=1.415
r387 (  120 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.085 //y=0.76 //x2=22.97 //y2=0.76
r388 (  119 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.305 //y=0.76 //x2=23.42 //y2=0.76
r389 (  119 120 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=23.305 //y=0.76 //x2=23.085 //y2=0.76
r390 (  116 153 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=23.12 //y=4.865 //x2=22.94 //y2=4.7
r391 (  114 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.57 //x2=22.97 //y2=1.415
r392 (  114 148 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.57 //x2=22.93 //y2=1.915
r393 (  113 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.26 //x2=22.97 //y2=1.415
r394 (  112 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=0.915 //x2=22.97 //y2=0.76
r395 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.93 //y=0.915 //x2=22.93 //y2=1.26
r396 (  109 153 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=22.68 //y=4.865 //x2=22.94 //y2=4.7
r397 (  108 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.99 //y=1.26 //x2=11.95 //y2=1.415
r398 (  107 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.99 //y=0.915 //x2=11.95 //y2=0.76
r399 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.99 //y=0.915 //x2=11.99 //y2=1.26
r400 (  105 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.615 //y=1.415 //x2=11.5 //y2=1.415
r401 (  104 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.835 //y=1.415 //x2=11.95 //y2=1.415
r402 (  103 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.615 //y=0.76 //x2=11.5 //y2=0.76
r403 (  102 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.835 //y=0.76 //x2=11.95 //y2=0.76
r404 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=11.835 //y=0.76 //x2=11.615 //y2=0.76
r405 (  99 143 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=11.65 //y=4.865 //x2=11.47 //y2=4.7
r406 (  97 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.57 //x2=11.5 //y2=1.415
r407 (  97 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.57 //x2=11.46 //y2=1.915
r408 (  96 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.26 //x2=11.5 //y2=1.415
r409 (  95 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=0.915 //x2=11.5 //y2=0.76
r410 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.46 //y=0.915 //x2=11.46 //y2=1.26
r411 (  92 143 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=11.21 //y=4.865 //x2=11.47 //y2=4.7
r412 (  91 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.18 //y=1.26 //x2=7.14 //y2=1.415
r413 (  90 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.18 //y=0.915 //x2=7.14 //y2=0.76
r414 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.18 //y=0.915 //x2=7.18 //y2=1.26
r415 (  88 131 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.805 //y=1.415 //x2=6.69 //y2=1.415
r416 (  87 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.025 //y=1.415 //x2=7.14 //y2=1.415
r417 (  86 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.805 //y=0.76 //x2=6.69 //y2=0.76
r418 (  85 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.025 //y=0.76 //x2=7.14 //y2=0.76
r419 (  85 86 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.025 //y=0.76 //x2=6.805 //y2=0.76
r420 (  82 133 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=6.84 //y=4.865 //x2=6.66 //y2=4.7
r421 (  80 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.57 //x2=6.69 //y2=1.415
r422 (  80 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.57 //x2=6.65 //y2=1.915
r423 (  79 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.26 //x2=6.69 //y2=1.415
r424 (  78 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=0.915 //x2=6.69 //y2=0.76
r425 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.65 //y=0.915 //x2=6.65 //y2=1.26
r426 (  75 133 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=6.4 //y=4.865 //x2=6.66 //y2=4.7
r427 (  74 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.12 //y=6.02 //x2=23.12 //y2=4.865
r428 (  73 109 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.68 //y=6.02 //x2=22.68 //y2=4.865
r429 (  72 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.65 //y=6.02 //x2=11.65 //y2=4.865
r430 (  71 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.21 //y=6.02 //x2=11.21 //y2=4.865
r431 (  70 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.84 //y=6.02 //x2=6.84 //y2=4.865
r432 (  69 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.4 //y=6.02 //x2=6.4 //y2=4.865
r433 (  68 121 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.195 //y=1.415 //x2=23.305 //y2=1.415
r434 (  68 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.195 //y=1.415 //x2=23.085 //y2=1.415
r435 (  67 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.725 //y=1.415 //x2=11.835 //y2=1.415
r436 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.725 //y=1.415 //x2=11.615 //y2=1.415
r437 (  66 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.915 //y=1.415 //x2=7.025 //y2=1.415
r438 (  66 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.915 //y=1.415 //x2=6.805 //y2=1.415
r439 (  63 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.94 //y=4.7 //x2=22.94 //y2=4.7
r440 (  61 63 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=22.94 //y=3.7 //x2=22.94 //y2=4.7
r441 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.94 //y=2.08 //x2=22.94 //y2=2.08
r442 (  58 61 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=22.94 //y=2.08 //x2=22.94 //y2=3.7
r443 (  54 56 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=15.54 //y=5.115 //x2=15.54 //y2=3.7
r444 (  53 56 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=15.54 //y=1.74 //x2=15.54 //y2=3.7
r445 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.455 //y=1.655 //x2=15.54 //y2=1.74
r446 (  51 52 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=15.455 //y=1.655 //x2=15.185 //y2=1.655
r447 (  50 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.145 //y=5.2 //x2=15.06 //y2=5.2
r448 (  49 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.455 //y=5.2 //x2=15.54 //y2=5.115
r449 (  49 50 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=15.455 //y=5.2 //x2=15.145 //y2=5.2
r450 (  45 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.1 //y=1.57 //x2=15.185 //y2=1.655
r451 (  45 156 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=15.1 //y=1.57 //x2=15.1 //y2=1
r452 (  39 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.06 //y=5.285 //x2=15.06 //y2=5.2
r453 (  39 159 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=15.06 //y=5.285 //x2=15.06 //y2=5.725
r454 (  37 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.975 //y=5.2 //x2=15.06 //y2=5.2
r455 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=14.975 //y=5.2 //x2=14.265 //y2=5.2
r456 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.18 //y=5.285 //x2=14.265 //y2=5.2
r457 (  31 158 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=14.18 //y=5.285 //x2=14.18 //y2=5.725
r458 (  29 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=4.7 //x2=11.47 //y2=4.7
r459 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=11.47 //y=3.7 //x2=11.47 //y2=4.7
r460 (  24 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=2.08 //x2=11.47 //y2=2.08
r461 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=11.47 //y=2.08 //x2=11.47 //y2=3.7
r462 (  21 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=4.7 //x2=6.66 //y2=4.7
r463 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=6.66 //y=3.7 //x2=6.66 //y2=4.7
r464 (  16 127 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.08 //x2=6.66 //y2=2.08
r465 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.08 //x2=6.66 //y2=3.7
r466 (  14 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=22.94 //y=3.7 //x2=22.94 //y2=3.7
r467 (  12 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=3.7 //x2=15.54 //y2=3.7
r468 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.47 //y=3.7 //x2=11.47 //y2=3.7
r469 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=3.7 //x2=6.66 //y2=3.7
r470 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.655 //y=3.7 //x2=15.54 //y2=3.7
r471 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=22.825 //y=3.7 //x2=22.94 //y2=3.7
r472 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=22.825 //y=3.7 //x2=15.655 //y2=3.7
r473 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.585 //y=3.7 //x2=11.47 //y2=3.7
r474 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=3.7 //x2=15.54 //y2=3.7
r475 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=3.7 //x2=11.585 //y2=3.7
r476 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.775 //y=3.7 //x2=6.66 //y2=3.7
r477 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=3.7 //x2=11.47 //y2=3.7
r478 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=3.7 //x2=6.775 //y2=3.7
ends PM_DFFSNQX1\%noxref_9

subckt PM_DFFSNQX1\%Q ( 1 2 7 8 9 10 11 12 13 14 15 16 17 18 19 20 22 36 37 44 \
 52 58 59 73 74 75 76 77 78 79 80 85 87 89 95 96 98 99 102 110 112 113 114 )
c170 ( 114 0 ) capacitor c=0.023087f //x=22.755 //y=5.02
c171 ( 113 0 ) capacitor c=0.023519f //x=21.875 //y=5.02
c172 ( 112 0 ) capacitor c=0.0224735f //x=20.995 //y=5.02
c173 ( 110 0 ) capacitor c=0.00853354f //x=23.005 //y=0.915
c174 ( 102 0 ) capacitor c=0.0332623f //x=18.16 //y=4.7
c175 ( 99 0 ) capacitor c=0.0279499f //x=18.13 //y=1.915
c176 ( 98 0 ) capacitor c=0.0422904f //x=18.13 //y=2.08
c177 ( 96 0 ) capacitor c=0.0429696f //x=18.695 //y=1.25
c178 ( 95 0 ) capacitor c=0.0192208f //x=18.695 //y=0.905
c179 ( 89 0 ) capacitor c=0.0148884f //x=18.54 //y=1.405
c180 ( 87 0 ) capacitor c=0.0157803f //x=18.54 //y=0.75
c181 ( 85 0 ) capacitor c=0.0306375f //x=18.535 //y=4.79
c182 ( 80 0 ) capacitor c=0.0205163f //x=18.165 //y=1.56
c183 ( 79 0 ) capacitor c=0.0168481f //x=18.165 //y=1.25
c184 ( 78 0 ) capacitor c=0.0174783f //x=18.165 //y=0.905
c185 ( 77 0 ) capacitor c=0.15358f //x=18.61 //y=6.02
c186 ( 76 0 ) capacitor c=0.110281f //x=18.17 //y=6.02
c187 ( 74 0 ) capacitor c=0.00125237f //x=22.9 //y=5.155
c188 ( 73 0 ) capacitor c=0.00243871f //x=22.02 //y=5.155
c189 ( 59 0 ) capacitor c=0.00493499f //x=23.28 //y=1.665
c190 ( 58 0 ) capacitor c=0.0154014f //x=23.595 //y=1.665
c191 ( 52 0 ) capacitor c=0.0304842f //x=23.595 //y=5.155
c192 ( 44 0 ) capacitor c=0.0191592f //x=22.815 //y=5.155
c193 ( 37 0 ) capacitor c=0.00369455f //x=21.225 //y=5.155
c194 ( 36 0 ) capacitor c=0.0161734f //x=21.935 //y=5.155
c195 ( 22 0 ) capacitor c=0.0737377f //x=18.13 //y=2.08
c196 ( 20 0 ) capacitor c=0.00453889f //x=18.13 //y=4.535
c197 ( 12 0 ) capacitor c=0.130008f //x=23.68 //y=2.22
c198 ( 2 0 ) capacitor c=0.0143991f //x=18.245 //y=3.33
c199 ( 1 0 ) capacitor c=0.130302f //x=23.565 //y=3.33
r200 (  104 105 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=18.16 //y=4.79 //x2=18.16 //y2=4.865
r201 (  102 104 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=18.16 //y=4.7 //x2=18.16 //y2=4.79
r202 (  98 99 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=18.13 //y=2.08 //x2=18.13 //y2=1.915
r203 (  96 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.695 //y=1.25 //x2=18.655 //y2=1.405
r204 (  95 108 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.695 //y=0.905 //x2=18.655 //y2=0.75
r205 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.695 //y=0.905 //x2=18.695 //y2=1.25
r206 (  90 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.32 //y=1.405 //x2=18.205 //y2=1.405
r207 (  89 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.54 //y=1.405 //x2=18.655 //y2=1.405
r208 (  88 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.32 //y=0.75 //x2=18.205 //y2=0.75
r209 (  87 108 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.54 //y=0.75 //x2=18.655 //y2=0.75
r210 (  87 88 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.54 //y=0.75 //x2=18.32 //y2=0.75
r211 (  86 104 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=18.295 //y=4.79 //x2=18.16 //y2=4.79
r212 (  85 92 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.79 //x2=18.61 //y2=4.865
r213 (  85 86 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.79 //x2=18.295 //y2=4.79
r214 (  80 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.56 //x2=18.205 //y2=1.405
r215 (  80 99 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.56 //x2=18.165 //y2=1.915
r216 (  79 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.25 //x2=18.205 //y2=1.405
r217 (  78 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=0.905 //x2=18.205 //y2=0.75
r218 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.165 //y=0.905 //x2=18.165 //y2=1.25
r219 (  77 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.61 //y=6.02 //x2=18.61 //y2=4.865
r220 (  76 105 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.17 //y=6.02 //x2=18.17 //y2=4.865
r221 (  75 89 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.43 //y=1.405 //x2=18.54 //y2=1.405
r222 (  75 90 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.43 //y=1.405 //x2=18.32 //y2=1.405
r223 (  72 102 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.16 //y=4.7 //x2=18.16 //y2=4.7
r224 (  58 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.595 //y=1.665 //x2=23.68 //y2=1.75
r225 (  58 59 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=23.595 //y=1.665 //x2=23.28 //y2=1.665
r226 (  54 59 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.195 //y=1.58 //x2=23.28 //y2=1.665
r227 (  54 110 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.195 //y=1.58 //x2=23.195 //y2=1.01
r228 (  53 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.985 //y=5.155 //x2=22.9 //y2=5.155
r229 (  52 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.595 //y=5.155 //x2=23.68 //y2=5.07
r230 (  52 53 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=23.595 //y=5.155 //x2=22.985 //y2=5.155
r231 (  46 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.9 //y=5.24 //x2=22.9 //y2=5.155
r232 (  46 114 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.9 //y=5.24 //x2=22.9 //y2=5.725
r233 (  45 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.105 //y=5.155 //x2=22.02 //y2=5.155
r234 (  44 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.815 //y=5.155 //x2=22.9 //y2=5.155
r235 (  44 45 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.815 //y=5.155 //x2=22.105 //y2=5.155
r236 (  38 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.02 //y=5.24 //x2=22.02 //y2=5.155
r237 (  38 113 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.02 //y=5.24 //x2=22.02 //y2=5.725
r238 (  36 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.935 //y=5.155 //x2=22.02 //y2=5.155
r239 (  36 37 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=21.935 //y=5.155 //x2=21.225 //y2=5.155
r240 (  30 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.14 //y=5.24 //x2=21.225 //y2=5.155
r241 (  30 112 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.14 //y=5.24 //x2=21.14 //y2=5.725
r242 (  22 98 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.13 //y=2.08 //x2=18.13 //y2=2.08
r243 (  20 72 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.535 //x2=18.145 //y2=4.7
r244 (  19 61 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=23.68 //y=4.81 //x2=23.68 //y2=5.07
r245 (  18 19 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=4.44 //x2=23.68 //y2=4.81
r246 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=4.07 //x2=23.68 //y2=4.44
r247 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=3.7 //x2=23.68 //y2=4.07
r248 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=3.33 //x2=23.68 //y2=3.7
r249 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=2.96 //x2=23.68 //y2=3.33
r250 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=2.59 //x2=23.68 //y2=2.96
r251 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=2.22 //x2=23.68 //y2=2.59
r252 (  12 60 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=23.68 //y=2.22 //x2=23.68 //y2=1.75
r253 (  11 20 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.44 //x2=18.13 //y2=4.535
r254 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.07 //x2=18.13 //y2=4.44
r255 (  9 10 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=18.13 //y=3.33 //x2=18.13 //y2=4.07
r256 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=18.13 //y=2.96 //x2=18.13 //y2=3.33
r257 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=18.13 //y=2.59 //x2=18.13 //y2=2.96
r258 (  7 22 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=18.13 //y=2.59 //x2=18.13 //y2=2.08
r259 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.68 //y=3.33 //x2=23.68 //y2=3.33
r260 (  4 9 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.13 //y=3.33 //x2=18.13 //y2=3.33
r261 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.245 //y=3.33 //x2=18.13 //y2=3.33
r262 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.565 //y=3.33 //x2=23.68 //y2=3.33
r263 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=23.565 //y=3.33 //x2=18.245 //y2=3.33
ends PM_DFFSNQX1\%Q

subckt PM_DFFSNQX1\%D ( 1 2 3 4 5 6 8 19 20 21 22 23 24 25 29 31 34 35 45 )
c57 ( 45 0 ) capacitor c=0.0667949f //x=1.11 //y=4.7
c58 ( 35 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c59 ( 34 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c60 ( 31 0 ) capacitor c=0.0141798f //x=1.29 //y=1.365
c61 ( 29 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c62 ( 25 0 ) capacitor c=0.0860049f //x=0.915 //y=1.915
c63 ( 24 0 ) capacitor c=0.0229722f //x=0.915 //y=1.52
c64 ( 23 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c65 ( 22 0 ) capacitor c=0.0199343f //x=0.915 //y=0.865
c66 ( 21 0 ) capacitor c=0.110275f //x=1.45 //y=6.02
c67 ( 20 0 ) capacitor c=0.154305f //x=1.01 //y=6.02
c68 ( 8 0 ) capacitor c=0.115639f //x=1.11 //y=2.08
r69 (  43 45 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.7 //x2=1.11 //y2=4.7
r70 (  36 45 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=1.45 //y=4.865 //x2=1.11 //y2=4.7
r71 (  35 47 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r72 (  34 46 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r73 (  34 35 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r74 (  32 42 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r75 (  31 47 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r76 (  30 41 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r77 (  29 46 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r78 (  29 30 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r79 (  26 43 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.865 //x2=1.01 //y2=4.7
r80 (  25 40 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r81 (  24 42 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r82 (  24 25 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r83 (  23 42 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r84 (  22 41 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r85 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r86 (  21 36 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.02 //x2=1.45 //y2=4.865
r87 (  20 26 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.02 //x2=1.01 //y2=4.865
r88 (  19 31 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r89 (  19 32 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r90 (  17 45 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r91 (  8 40 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r92 (  6 17 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.44 //x2=1.11 //y2=4.7
r93 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r94 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r95 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r96 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r97 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r98 (  1 8 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.59 //x2=1.11 //y2=2.08
ends PM_DFFSNQX1\%D

subckt PM_DFFSNQX1\%noxref_12 ( 1 5 9 10 13 17 29 )
c48 ( 29 0 ) capacitor c=0.0632971f //x=0.56 //y=0.365
c49 ( 17 0 ) capacitor c=0.0072343f //x=2.635 //y=0.615
c50 ( 13 0 ) capacitor c=0.015427f //x=2.55 //y=0.53
c51 ( 10 0 ) capacitor c=0.00896024f //x=1.665 //y=1.495
c52 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c53 ( 5 0 ) capacitor c=0.0255599f //x=1.58 //y=1.58
c54 ( 1 0 ) capacitor c=0.0113547f //x=0.695 //y=1.495
r55 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r56 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r57 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r58 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=2.15 //y2=0.53
r59 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r60 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.15 //y2=0.53
r61 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r62 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r63 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r64 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r65 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r66 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r67 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r68 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r69 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r70 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_DFFSNQX1\%noxref_12

subckt PM_DFFSNQX1\%noxref_13 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0680128f //x=3.785 //y=0.375
c53 ( 17 0 ) capacitor c=0.018806f //x=5.775 //y=1.59
c54 ( 13 0 ) capacitor c=0.0155484f //x=5.775 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=4.89 //y=0.625
c56 ( 5 0 ) capacitor c=0.017077f //x=4.805 //y=1.59
c57 ( 1 0 ) capacitor c=0.00729042f //x=3.92 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.975 //y=1.59 //x2=4.89 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.975 //y=1.59 //x2=5.375 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.775 //y=1.59 //x2=5.86 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.775 //y=1.59 //x2=5.375 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.975 //y=0.54 //x2=4.89 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.975 //y=0.54 //x2=5.375 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.775 //y=0.54 //x2=5.86 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.775 //y=0.54 //x2=5.375 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.89 //y=1.505 //x2=4.89 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=4.89 //y=1.505 //x2=4.89 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=4.89 //y=0.625 //x2=4.89 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=4.89 //y=0.625 //x2=4.89 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.005 //y=1.59 //x2=3.92 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.005 //y=1.59 //x2=4.405 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.805 //y=1.59 //x2=4.89 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.805 //y=1.59 //x2=4.405 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.92 //y=1.505 //x2=3.92 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=3.92 //y=1.505 //x2=3.92 //y2=0.89
ends PM_DFFSNQX1\%noxref_13

subckt PM_DFFSNQX1\%noxref_14 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.041888f //x=6.295 //y=0.375
c54 ( 28 0 ) capacitor c=0.00460056f //x=5.19 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=6.43 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=7.4 //y=0.625
c57 ( 11 0 ) capacitor c=0.0145763f //x=7.315 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=6.43 //y=0.625
c59 ( 1 0 ) capacitor c=0.022894f //x=6.345 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.4 //y=0.625 //x2=7.4 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=7.4 //y=0.625 //x2=7.4 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.515 //y=0.54 //x2=6.43 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.515 //y=0.54 //x2=6.915 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.315 //y=0.54 //x2=7.4 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.315 //y=0.54 //x2=6.915 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.43 //y=1.08 //x2=6.43 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=6.43 //y=1.08 //x2=6.43 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.91 //x2=6.43 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.91 //x2=6.43 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.625 //x2=6.43 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.625 //x2=6.43 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.465 //y=0.995 //x2=5.38 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.345 //y=0.995 //x2=6.43 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=6.345 //y=0.995 //x2=5.465 //y2=0.995
ends PM_DFFSNQX1\%noxref_14

subckt PM_DFFSNQX1\%noxref_15 ( 1 5 9 13 17 35 )
c54 ( 35 0 ) capacitor c=0.0685332f //x=8.595 //y=0.375
c55 ( 17 0 ) capacitor c=0.0207646f //x=10.585 //y=1.59
c56 ( 13 0 ) capacitor c=0.0155144f //x=10.585 //y=0.54
c57 ( 9 0 ) capacitor c=0.00678203f //x=9.7 //y=0.625
c58 ( 5 0 ) capacitor c=0.0181938f //x=9.615 //y=1.59
c59 ( 1 0 ) capacitor c=0.00729042f //x=8.73 //y=1.505
r60 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.785 //y=1.59 //x2=9.7 //y2=1.63
r61 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.785 //y=1.59 //x2=10.185 //y2=1.59
r62 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.585 //y=1.59 //x2=10.67 //y2=1.59
r63 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.585 //y=1.59 //x2=10.185 //y2=1.59
r64 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.785 //y=0.54 //x2=9.7 //y2=0.5
r65 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.785 //y=0.54 //x2=10.185 //y2=0.54
r66 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.585 //y=0.54 //x2=10.67 //y2=0.54
r67 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.585 //y=0.54 //x2=10.185 //y2=0.54
r68 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.7 //y=1.505 //x2=9.7 //y2=1.63
r69 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.7 //y=1.505 //x2=9.7 //y2=0.89
r70 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.7 //y=0.625 //x2=9.7 //y2=0.5
r71 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=9.7 //y=0.625 //x2=9.7 //y2=0.89
r72 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.815 //y=1.59 //x2=8.73 //y2=1.63
r73 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.815 //y=1.59 //x2=9.215 //y2=1.59
r74 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.615 //y=1.59 //x2=9.7 //y2=1.63
r75 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.615 //y=1.59 //x2=9.215 //y2=1.59
r76 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.73 //y=1.505 //x2=8.73 //y2=1.63
r77 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.73 //y=1.505 //x2=8.73 //y2=0.89
ends PM_DFFSNQX1\%noxref_15

subckt PM_DFFSNQX1\%noxref_16 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0414744f //x=11.105 //y=0.375
c54 ( 28 0 ) capacitor c=0.00461914f //x=10 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=11.24 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=12.21 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144274f //x=12.125 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=11.24 //y=0.625
c59 ( 1 0 ) capacitor c=0.0220663f //x=11.155 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=12.21 //y=0.625 //x2=12.21 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=12.21 //y=0.625 //x2=12.21 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.325 //y=0.54 //x2=11.24 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.325 //y=0.54 //x2=11.725 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.125 //y=0.54 //x2=12.21 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.125 //y=0.54 //x2=11.725 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.24 //y=1.08 //x2=11.24 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=11.24 //y=1.08 //x2=11.24 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.91 //x2=11.24 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.91 //x2=11.24 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.625 //x2=11.24 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.625 //x2=11.24 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.275 //y=0.995 //x2=10.19 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.155 //y=0.995 //x2=11.24 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=11.155 //y=0.995 //x2=10.275 //y2=0.995
ends PM_DFFSNQX1\%noxref_16

subckt PM_DFFSNQX1\%noxref_17 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632682f //x=13.51 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=15.585 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=15.5 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=14.615 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=14.615 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=14.53 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=13.645 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=15.585 //y=0.615 //x2=15.585 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.585 //y=0.615 //x2=15.585 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.7 //y=0.53 //x2=14.615 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.7 //y=0.53 //x2=15.1 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.5 //y=0.53 //x2=15.585 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.5 //y=0.53 //x2=15.1 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.615 //y=1.495 //x2=14.615 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=14.615 //y=1.495 //x2=14.615 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=14.615 //y=0.615 //x2=14.615 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=14.615 //y=0.615 //x2=14.615 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.73 //y=1.58 //x2=13.645 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.73 //y=1.58 //x2=14.13 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.53 //y=1.58 //x2=14.615 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.53 //y=1.58 //x2=14.13 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=13.645 //y=1.495 //x2=13.645 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.645 //y=1.495 //x2=13.645 //y2=0.88
ends PM_DFFSNQX1\%noxref_17

subckt PM_DFFSNQX1\%noxref_18 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632684f //x=16.84 //y=0.365
c53 ( 17 0 ) capacitor c=0.0072343f //x=18.915 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=18.83 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=17.945 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=17.945 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=17.86 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=16.975 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=18.915 //y=0.615 //x2=18.915 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.915 //y=0.615 //x2=18.915 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.03 //y=0.53 //x2=17.945 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.03 //y=0.53 //x2=18.43 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.83 //y=0.53 //x2=18.915 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.83 //y=0.53 //x2=18.43 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=17.945 //y=1.495 //x2=17.945 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=17.945 //y=1.495 //x2=17.945 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=17.945 //y=0.615 //x2=17.945 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=17.945 //y=0.615 //x2=17.945 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.06 //y=1.58 //x2=16.975 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.06 //y=1.58 //x2=17.46 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.86 //y=1.58 //x2=17.945 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.86 //y=1.58 //x2=17.46 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=16.975 //y=1.495 //x2=16.975 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=16.975 //y=1.495 //x2=16.975 //y2=0.88
ends PM_DFFSNQX1\%noxref_18

subckt PM_DFFSNQX1\%noxref_19 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0683476f //x=20.065 //y=0.375
c51 ( 17 0 ) capacitor c=0.018143f //x=22.055 //y=1.59
c52 ( 13 0 ) capacitor c=0.0155396f //x=22.055 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=21.17 //y=0.625
c54 ( 5 0 ) capacitor c=0.0164013f //x=21.085 //y=1.59
c55 ( 1 0 ) capacitor c=0.00696517f //x=20.2 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.255 //y=1.59 //x2=21.17 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.255 //y=1.59 //x2=21.655 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.055 //y=1.59 //x2=22.14 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.055 //y=1.59 //x2=21.655 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.255 //y=0.54 //x2=21.17 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.255 //y=0.54 //x2=21.655 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.055 //y=0.54 //x2=22.14 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.055 //y=0.54 //x2=21.655 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=21.17 //y=1.505 //x2=21.17 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=21.17 //y=1.505 //x2=21.17 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=21.17 //y=0.625 //x2=21.17 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=21.17 //y=0.625 //x2=21.17 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.285 //y=1.59 //x2=20.2 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.285 //y=1.59 //x2=20.685 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.085 //y=1.59 //x2=21.17 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.085 //y=1.59 //x2=20.685 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.2 //y=1.505 //x2=20.2 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=20.2 //y=1.505 //x2=20.2 //y2=0.89
ends PM_DFFSNQX1\%noxref_19

subckt PM_DFFSNQX1\%noxref_20 ( 1 3 11 15 25 28 29 )
c50 ( 29 0 ) capacitor c=0.0425456f //x=22.575 //y=0.375
c51 ( 28 0 ) capacitor c=0.00457437f //x=21.47 //y=0.91
c52 ( 25 0 ) capacitor c=0.00156479f //x=22.71 //y=0.995
c53 ( 15 0 ) capacitor c=0.00737666f //x=23.68 //y=0.625
c54 ( 11 0 ) capacitor c=0.0147903f //x=23.595 //y=0.54
c55 ( 3 0 ) capacitor c=0.00718386f //x=22.71 //y=0.625
c56 ( 1 0 ) capacitor c=0.0240499f //x=22.625 //y=0.995
r57 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.68 //y=0.625 //x2=23.68 //y2=0.5
r58 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=23.68 //y=0.625 //x2=23.68 //y2=0.89
r59 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.795 //y=0.54 //x2=22.71 //y2=0.5
r60 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.795 //y=0.54 //x2=23.195 //y2=0.54
r61 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.595 //y=0.54 //x2=23.68 //y2=0.5
r62 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.595 //y=0.54 //x2=23.195 //y2=0.54
r63 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.71 //y=1.08 //x2=22.71 //y2=0.995
r64 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=22.71 //y=1.08 //x2=22.71 //y2=1.23
r65 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.91 //x2=22.71 //y2=0.995
r66 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.91 //x2=22.71 //y2=0.89
r67 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.625 //x2=22.71 //y2=0.5
r68 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.625 //x2=22.71 //y2=0.89
r69 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.745 //y=0.995 //x2=21.66 //y2=0.995
r70 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.625 //y=0.995 //x2=22.71 //y2=0.995
r71 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=22.625 //y=0.995 //x2=21.745 //y2=0.995
ends PM_DFFSNQX1\%noxref_20

