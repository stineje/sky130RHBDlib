magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 145 157 415 203
rect 48 21 415 157
rect 48 17 63 21
rect 29 -17 63 17
<< locali >>
rect 331 370 443 493
rect 20 145 65 265
rect 192 213 265 265
rect 407 179 443 370
rect 247 145 443 179
rect 247 51 313 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 83 336 135 381
rect 175 371 241 527
rect 83 302 341 336
rect 99 109 135 302
rect 307 249 341 302
rect 307 215 373 249
rect 66 74 135 109
rect 171 17 213 179
rect 347 17 424 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 20 145 65 265 6 A
port 1 nsew signal input
rlabel locali s 192 213 265 265 6 SLEEP
port 2 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 48 17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 48 21 415 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 145 157 415 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 247 51 313 145 6 X
port 7 nsew signal output
rlabel locali s 247 145 443 179 6 X
port 7 nsew signal output
rlabel locali s 407 179 443 370 6 X
port 7 nsew signal output
rlabel locali s 331 370 443 493 6 X
port 7 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 460 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2370900
string GDS_START 2366634
<< end >>
