// File: dffsnrnx1_pcell.spi.DFFSNRNX1_PCELL.pxi
// Created: Tue Oct 15 15:56:04 2024
// 
simulator lang=spectre
x_PM_DFFSNRNX1_PCELL\%noxref_1 ( N_noxref_1_c_71_p N_noxref_1_c_106_p \
 N_noxref_1_c_1_p N_noxref_1_c_72_p N_noxref_1_c_16_p N_noxref_1_c_23_p \
 N_noxref_1_c_26_p N_noxref_1_c_33_p N_noxref_1_c_42_p N_noxref_1_c_49_p \
 N_noxref_1_c_60_p N_noxref_1_c_67_p N_noxref_1_c_93_p N_noxref_1_c_2_p \
 N_noxref_1_c_3_p N_noxref_1_c_4_p N_noxref_1_c_5_p N_noxref_1_c_6_p \
 N_noxref_1_c_7_p N_noxref_1_M0_noxref_d N_noxref_1_M3_noxref_d \
 N_noxref_1_M6_noxref_d N_noxref_1_M9_noxref_d N_noxref_1_M12_noxref_d \
 N_noxref_1_M15_noxref_d )  PM_DFFSNRNX1_PCELL\%noxref_1
x_PM_DFFSNRNX1_PCELL\%noxref_2 ( N_noxref_2_c_320_p N_noxref_2_c_313_n \
 N_noxref_2_c_321_p N_noxref_2_c_322_p N_noxref_2_c_328_p N_noxref_2_c_332_p \
 N_noxref_2_c_341_p N_noxref_2_c_423_p N_noxref_2_c_444_p N_noxref_2_c_408_p \
 N_noxref_2_c_409_p N_noxref_2_c_345_p N_noxref_2_c_370_p N_noxref_2_c_376_p \
 N_noxref_2_c_380_p N_noxref_2_c_412_p N_noxref_2_c_386_p N_noxref_2_c_427_p \
 N_noxref_2_c_488_p N_noxref_2_c_531_p N_noxref_2_c_458_p N_noxref_2_c_492_p \
 N_noxref_2_c_572_p N_noxref_2_c_588_p N_noxref_2_c_609_p N_noxref_2_c_504_p \
 N_noxref_2_c_543_p N_noxref_2_c_314_n N_noxref_2_c_315_n N_noxref_2_c_316_n \
 N_noxref_2_c_317_n N_noxref_2_c_318_n N_noxref_2_c_319_n \
 N_noxref_2_M18_noxref_s N_noxref_2_M19_noxref_d N_noxref_2_M21_noxref_d \
 N_noxref_2_M23_noxref_d N_noxref_2_M24_noxref_s N_noxref_2_M25_noxref_d \
 N_noxref_2_M27_noxref_d N_noxref_2_M29_noxref_d N_noxref_2_M30_noxref_s \
 N_noxref_2_M31_noxref_d N_noxref_2_M33_noxref_d N_noxref_2_M35_noxref_d \
 N_noxref_2_M36_noxref_s N_noxref_2_M37_noxref_d N_noxref_2_M39_noxref_d \
 N_noxref_2_M41_noxref_d N_noxref_2_M42_noxref_s N_noxref_2_M43_noxref_d \
 N_noxref_2_M45_noxref_d N_noxref_2_M47_noxref_d N_noxref_2_M48_noxref_s \
 N_noxref_2_M49_noxref_d N_noxref_2_M51_noxref_d N_noxref_2_M53_noxref_d )  \
 PM_DFFSNRNX1_PCELL\%noxref_2
x_PM_DFFSNRNX1_PCELL\%noxref_3 ( N_noxref_3_c_644_n N_noxref_3_c_645_n \
 N_noxref_3_c_646_n N_noxref_3_c_647_n N_noxref_3_c_673_n N_noxref_3_c_677_n \
 N_noxref_3_c_679_n N_noxref_3_c_683_n N_noxref_3_c_648_n N_noxref_3_c_803_p \
 N_noxref_3_c_649_n N_noxref_3_c_650_n N_noxref_3_c_651_n N_noxref_3_c_807_p \
 N_noxref_3_c_764_p N_noxref_3_M3_noxref_g N_noxref_3_M6_noxref_g \
 N_noxref_3_M24_noxref_g N_noxref_3_M25_noxref_g N_noxref_3_M30_noxref_g \
 N_noxref_3_M31_noxref_g N_noxref_3_c_652_n N_noxref_3_c_654_n \
 N_noxref_3_c_655_n N_noxref_3_c_656_n N_noxref_3_c_657_n N_noxref_3_c_658_n \
 N_noxref_3_c_659_n N_noxref_3_c_661_n N_noxref_3_c_736_p N_noxref_3_c_702_n \
 N_noxref_3_c_662_n N_noxref_3_c_664_n N_noxref_3_c_665_n N_noxref_3_c_666_n \
 N_noxref_3_c_667_n N_noxref_3_c_668_n N_noxref_3_c_669_n N_noxref_3_c_671_n \
 N_noxref_3_c_724_p N_noxref_3_c_704_n N_noxref_3_M2_noxref_d \
 N_noxref_3_M18_noxref_d N_noxref_3_M20_noxref_d N_noxref_3_M22_noxref_d )  \
 PM_DFFSNRNX1_PCELL\%noxref_3
x_PM_DFFSNRNX1_PCELL\%noxref_4 ( N_noxref_4_c_881_n N_noxref_4_c_882_n \
 N_noxref_4_c_897_n N_noxref_4_c_901_n N_noxref_4_c_903_n N_noxref_4_c_907_n \
 N_noxref_4_c_883_n N_noxref_4_c_976_p N_noxref_4_c_884_n N_noxref_4_c_885_n \
 N_noxref_4_c_991_p N_noxref_4_c_999_p N_noxref_4_M9_noxref_g \
 N_noxref_4_M36_noxref_g N_noxref_4_M37_noxref_g N_noxref_4_c_886_n \
 N_noxref_4_c_888_n N_noxref_4_c_889_n N_noxref_4_c_890_n N_noxref_4_c_891_n \
 N_noxref_4_c_892_n N_noxref_4_c_893_n N_noxref_4_c_895_n N_noxref_4_c_951_p \
 N_noxref_4_c_919_n N_noxref_4_M8_noxref_d N_noxref_4_M30_noxref_d \
 N_noxref_4_M32_noxref_d N_noxref_4_M34_noxref_d )  PM_DFFSNRNX1_PCELL\%noxref_4
x_PM_DFFSNRNX1_PCELL\%noxref_5 ( N_noxref_5_c_1045_n N_noxref_5_c_1056_n \
 N_noxref_5_c_1043_n N_noxref_5_c_1044_n N_noxref_5_M4_noxref_g \
 N_noxref_5_M10_noxref_g N_noxref_5_M26_noxref_g N_noxref_5_M27_noxref_g \
 N_noxref_5_M38_noxref_g N_noxref_5_M39_noxref_g N_noxref_5_c_1084_n \
 N_noxref_5_c_1087_n N_noxref_5_c_1215_p N_noxref_5_c_1222_p \
 N_noxref_5_c_1089_n N_noxref_5_c_1090_n N_noxref_5_c_1091_n \
 N_noxref_5_c_1092_n N_noxref_5_c_1140_p N_noxref_5_c_1112_n \
 N_noxref_5_c_1115_n N_noxref_5_c_1235_p N_noxref_5_c_1242_p \
 N_noxref_5_c_1117_n N_noxref_5_c_1118_n N_noxref_5_c_1119_n \
 N_noxref_5_c_1120_n N_noxref_5_c_1163_p N_noxref_5_c_1094_n \
 N_noxref_5_c_1122_n )  PM_DFFSNRNX1_PCELL\%noxref_5
x_PM_DFFSNRNX1_PCELL\%noxref_6 ( N_noxref_6_c_1247_n N_noxref_6_c_1266_n \
 N_noxref_6_c_1248_n N_noxref_6_c_1324_n N_noxref_6_c_1249_n \
 N_noxref_6_c_1268_n N_noxref_6_c_1272_n N_noxref_6_c_1274_n \
 N_noxref_6_c_1278_n N_noxref_6_c_1250_n N_noxref_6_c_1384_p \
 N_noxref_6_c_1282_n N_noxref_6_c_1251_n N_noxref_6_c_1375_n \
 N_noxref_6_c_1454_p N_noxref_6_M2_noxref_g N_noxref_6_M12_noxref_g \
 N_noxref_6_M22_noxref_g N_noxref_6_M23_noxref_g N_noxref_6_M42_noxref_g \
 N_noxref_6_M43_noxref_g N_noxref_6_c_1340_n N_noxref_6_c_1341_n \
 N_noxref_6_c_1342_n N_noxref_6_c_1343_n N_noxref_6_c_1344_n \
 N_noxref_6_c_1346_n N_noxref_6_c_1347_n N_noxref_6_c_1252_n \
 N_noxref_6_c_1254_n N_noxref_6_c_1255_n N_noxref_6_c_1256_n \
 N_noxref_6_c_1257_n N_noxref_6_c_1258_n N_noxref_6_c_1259_n \
 N_noxref_6_c_1261_n N_noxref_6_c_1403_p N_noxref_6_c_1294_n \
 N_noxref_6_c_1349_n N_noxref_6_c_1350_n N_noxref_6_c_1352_n \
 N_noxref_6_M5_noxref_d N_noxref_6_M24_noxref_d N_noxref_6_M26_noxref_d \
 N_noxref_6_M28_noxref_d )  PM_DFFSNRNX1_PCELL\%noxref_6
x_PM_DFFSNRNX1_PCELL\%noxref_7 ( N_noxref_7_c_1511_n N_noxref_7_c_1522_n \
 N_noxref_7_c_1523_n N_noxref_7_c_1527_n N_noxref_7_c_1528_n \
 N_noxref_7_c_1529_n N_noxref_7_c_1530_n N_noxref_7_M1_noxref_g \
 N_noxref_7_M11_noxref_g N_noxref_7_M13_noxref_g N_noxref_7_M20_noxref_g \
 N_noxref_7_M21_noxref_g N_noxref_7_M40_noxref_g N_noxref_7_M41_noxref_g \
 N_noxref_7_M44_noxref_g N_noxref_7_M45_noxref_g N_noxref_7_c_1706_p \
 N_noxref_7_c_1708_p N_noxref_7_c_1733_p N_noxref_7_c_1741_p \
 N_noxref_7_c_1629_n N_noxref_7_c_1630_n N_noxref_7_c_1631_n \
 N_noxref_7_c_1632_n N_noxref_7_c_1566_n N_noxref_7_c_1588_n \
 N_noxref_7_c_1589_n N_noxref_7_c_1590_n N_noxref_7_c_1692_p \
 N_noxref_7_c_1673_p N_noxref_7_c_1694_p N_noxref_7_c_1674_p \
 N_noxref_7_c_1636_n N_noxref_7_c_1639_n N_noxref_7_c_1815_p \
 N_noxref_7_c_1822_p N_noxref_7_c_1641_n N_noxref_7_c_1642_n \
 N_noxref_7_c_1643_n N_noxref_7_c_1644_n N_noxref_7_c_1665_p \
 N_noxref_7_c_1567_n N_noxref_7_c_1591_n N_noxref_7_c_1593_n \
 N_noxref_7_c_1594_n N_noxref_7_c_1648_n )  PM_DFFSNRNX1_PCELL\%noxref_7
x_PM_DFFSNRNX1_PCELL\%noxref_8 ( N_noxref_8_c_1827_n N_noxref_8_c_1847_n \
 N_noxref_8_c_1833_n N_noxref_8_c_1834_n N_noxref_8_M7_noxref_g \
 N_noxref_8_M16_noxref_g N_noxref_8_M32_noxref_g N_noxref_8_M33_noxref_g \
 N_noxref_8_M50_noxref_g N_noxref_8_M51_noxref_g N_noxref_8_c_1856_n \
 N_noxref_8_c_1859_n N_noxref_8_c_1952_p N_noxref_8_c_1959_p \
 N_noxref_8_c_1861_n N_noxref_8_c_1862_n N_noxref_8_c_1863_n \
 N_noxref_8_c_1864_n N_noxref_8_c_1879_n N_noxref_8_c_1981_p \
 N_noxref_8_c_1983_p N_noxref_8_c_2016_p N_noxref_8_c_2023_p \
 N_noxref_8_c_1929_p N_noxref_8_c_1930_p N_noxref_8_c_1931_p \
 N_noxref_8_c_1918_p N_noxref_8_c_1907_p N_noxref_8_c_1866_n \
 N_noxref_8_c_1908_p )  PM_DFFSNRNX1_PCELL\%noxref_8
x_PM_DFFSNRNX1_PCELL\%noxref_9 ( N_noxref_9_c_2034_n N_noxref_9_c_2090_n \
 N_noxref_9_c_2035_n N_noxref_9_c_2097_n N_noxref_9_c_2028_n \
 N_noxref_9_c_2042_n N_noxref_9_c_2029_n N_noxref_9_c_2030_n \
 N_noxref_9_c_2045_n N_noxref_9_c_2049_n N_noxref_9_c_2051_n \
 N_noxref_9_c_2055_n N_noxref_9_c_2031_n N_noxref_9_c_2218_n \
 N_noxref_9_c_2059_n N_noxref_9_c_2032_n N_noxref_9_c_2146_n \
 N_noxref_9_c_2226_n N_noxref_9_M5_noxref_g N_noxref_9_M8_noxref_g \
 N_noxref_9_M17_noxref_g N_noxref_9_M28_noxref_g N_noxref_9_M29_noxref_g \
 N_noxref_9_M34_noxref_g N_noxref_9_M35_noxref_g N_noxref_9_M52_noxref_g \
 N_noxref_9_M53_noxref_g N_noxref_9_c_2151_n N_noxref_9_c_2152_n \
 N_noxref_9_c_2153_n N_noxref_9_c_2191_n N_noxref_9_c_2192_n \
 N_noxref_9_c_2194_n N_noxref_9_c_2195_n N_noxref_9_c_2110_n \
 N_noxref_9_c_2111_n N_noxref_9_c_2112_n N_noxref_9_c_2113_n \
 N_noxref_9_c_2114_n N_noxref_9_c_2116_n N_noxref_9_c_2117_n \
 N_noxref_9_c_2272_n N_noxref_9_c_2273_n N_noxref_9_c_2274_n \
 N_noxref_9_c_2345_p N_noxref_9_c_2332_p N_noxref_9_c_2347_p \
 N_noxref_9_c_2333_p N_noxref_9_c_2154_n N_noxref_9_c_2156_n \
 N_noxref_9_c_2157_n N_noxref_9_c_2119_n N_noxref_9_c_2120_n \
 N_noxref_9_c_2122_n N_noxref_9_c_2281_n N_noxref_9_c_2283_n \
 N_noxref_9_c_2284_n N_noxref_9_M11_noxref_d N_noxref_9_M36_noxref_d \
 N_noxref_9_M38_noxref_d N_noxref_9_M40_noxref_d )  PM_DFFSNRNX1_PCELL\%noxref_9
x_PM_DFFSNRNX1_PCELL\%noxref_10 ( N_noxref_10_c_2364_n N_noxref_10_M0_noxref_g \
 N_noxref_10_M18_noxref_g N_noxref_10_M19_noxref_g N_noxref_10_c_2365_n \
 N_noxref_10_c_2367_n N_noxref_10_c_2368_n N_noxref_10_c_2369_n \
 N_noxref_10_c_2370_n N_noxref_10_c_2371_n N_noxref_10_c_2372_n \
 N_noxref_10_c_2374_n N_noxref_10_c_2387_n N_noxref_10_c_2382_n )  \
 PM_DFFSNRNX1_PCELL\%noxref_10
x_PM_DFFSNRNX1_PCELL\%noxref_11 ( N_noxref_11_c_2449_n N_noxref_11_c_2421_n \
 N_noxref_11_c_2425_n N_noxref_11_c_2428_n N_noxref_11_c_2440_n \
 N_noxref_11_M0_noxref_s )  PM_DFFSNRNX1_PCELL\%noxref_11
x_PM_DFFSNRNX1_PCELL\%noxref_12 ( N_noxref_12_c_2467_n N_noxref_12_c_2470_n \
 N_noxref_12_c_2473_n N_noxref_12_c_2476_n N_noxref_12_c_2484_n \
 N_noxref_12_M1_noxref_d N_noxref_12_M2_noxref_s )  \
 PM_DFFSNRNX1_PCELL\%noxref_12
x_PM_DFFSNRNX1_PCELL\%noxref_13 ( N_noxref_13_c_2537_n N_noxref_13_c_2521_n \
 N_noxref_13_c_2525_n N_noxref_13_c_2528_n N_noxref_13_c_2551_n \
 N_noxref_13_M3_noxref_s )  PM_DFFSNRNX1_PCELL\%noxref_13
x_PM_DFFSNRNX1_PCELL\%noxref_14 ( N_noxref_14_c_2571_n N_noxref_14_c_2574_n \
 N_noxref_14_c_2577_n N_noxref_14_c_2580_n N_noxref_14_c_2600_n \
 N_noxref_14_M4_noxref_d N_noxref_14_M5_noxref_s )  \
 PM_DFFSNRNX1_PCELL\%noxref_14
x_PM_DFFSNRNX1_PCELL\%noxref_15 ( N_noxref_15_c_2641_n N_noxref_15_c_2625_n \
 N_noxref_15_c_2629_n N_noxref_15_c_2632_n N_noxref_15_c_2656_n \
 N_noxref_15_M6_noxref_s )  PM_DFFSNRNX1_PCELL\%noxref_15
x_PM_DFFSNRNX1_PCELL\%noxref_16 ( N_noxref_16_c_2675_n N_noxref_16_c_2678_n \
 N_noxref_16_c_2681_n N_noxref_16_c_2684_n N_noxref_16_c_2692_n \
 N_noxref_16_M7_noxref_d N_noxref_16_M8_noxref_s )  \
 PM_DFFSNRNX1_PCELL\%noxref_16
x_PM_DFFSNRNX1_PCELL\%noxref_17 ( N_noxref_17_c_2745_n N_noxref_17_c_2729_n \
 N_noxref_17_c_2733_n N_noxref_17_c_2736_n N_noxref_17_c_2759_n \
 N_noxref_17_M9_noxref_s )  PM_DFFSNRNX1_PCELL\%noxref_17
x_PM_DFFSNRNX1_PCELL\%noxref_18 ( N_noxref_18_c_2779_n N_noxref_18_c_2782_n \
 N_noxref_18_c_2785_n N_noxref_18_c_2788_n N_noxref_18_c_2813_n \
 N_noxref_18_M10_noxref_d N_noxref_18_M11_noxref_s )  \
 PM_DFFSNRNX1_PCELL\%noxref_18
x_PM_DFFSNRNX1_PCELL\%noxref_19 ( N_noxref_19_c_2850_n N_noxref_19_c_2834_n \
 N_noxref_19_c_2838_n N_noxref_19_c_2841_n N_noxref_19_c_2864_n \
 N_noxref_19_M12_noxref_s )  PM_DFFSNRNX1_PCELL\%noxref_19
x_PM_DFFSNRNX1_PCELL\%noxref_20 ( N_noxref_20_c_2886_n \
 N_noxref_20_M14_noxref_g N_noxref_20_M46_noxref_g N_noxref_20_M47_noxref_g \
 N_noxref_20_c_2900_n N_noxref_20_c_2901_n N_noxref_20_c_2902_n \
 N_noxref_20_c_2928_p N_noxref_20_c_2917_p N_noxref_20_c_2930_p \
 N_noxref_20_c_2918_p N_noxref_20_c_2903_n N_noxref_20_c_2906_n \
 N_noxref_20_c_2907_n )  PM_DFFSNRNX1_PCELL\%noxref_20
x_PM_DFFSNRNX1_PCELL\%noxref_21 ( N_noxref_21_c_2947_n N_noxref_21_c_2951_n \
 N_noxref_21_c_2953_n N_noxref_21_c_2957_n N_noxref_21_c_2945_n \
 N_noxref_21_c_2989_n N_noxref_21_c_2961_n N_noxref_21_c_2986_n \
 N_noxref_21_c_3007_n N_noxref_21_M14_noxref_d N_noxref_21_M42_noxref_d \
 N_noxref_21_M44_noxref_d N_noxref_21_M46_noxref_d )  \
 PM_DFFSNRNX1_PCELL\%noxref_21
x_PM_DFFSNRNX1_PCELL\%noxref_22 ( N_noxref_22_c_3029_n N_noxref_22_c_3032_n \
 N_noxref_22_c_3035_n N_noxref_22_c_3038_n N_noxref_22_c_3071_n \
 N_noxref_22_M13_noxref_d N_noxref_22_M14_noxref_s )  \
 PM_DFFSNRNX1_PCELL\%noxref_22
x_PM_DFFSNRNX1_PCELL\%noxref_23 ( N_noxref_23_c_3083_n \
 N_noxref_23_M15_noxref_g N_noxref_23_M48_noxref_g N_noxref_23_M49_noxref_g \
 N_noxref_23_c_3084_n N_noxref_23_c_3086_n N_noxref_23_c_3087_n \
 N_noxref_23_c_3088_n N_noxref_23_c_3089_n N_noxref_23_c_3090_n \
 N_noxref_23_c_3091_n N_noxref_23_c_3093_n N_noxref_23_c_3121_n \
 N_noxref_23_c_3101_n )  PM_DFFSNRNX1_PCELL\%noxref_23
x_PM_DFFSNRNX1_PCELL\%noxref_24 ( N_noxref_24_c_3158_n N_noxref_24_c_3144_n \
 N_noxref_24_c_3148_n N_noxref_24_c_3151_n N_noxref_24_c_3162_n \
 N_noxref_24_M15_noxref_s )  PM_DFFSNRNX1_PCELL\%noxref_24
x_PM_DFFSNRNX1_PCELL\%noxref_25 ( N_noxref_25_c_3196_n N_noxref_25_c_3200_n \
 N_noxref_25_c_3202_n N_noxref_25_c_3206_n N_noxref_25_c_3194_n \
 N_noxref_25_c_3267_p N_noxref_25_c_3210_n N_noxref_25_c_3230_n \
 N_noxref_25_c_3246_n N_noxref_25_M17_noxref_d N_noxref_25_M48_noxref_d \
 N_noxref_25_M50_noxref_d N_noxref_25_M52_noxref_d )  \
 PM_DFFSNRNX1_PCELL\%noxref_25
x_PM_DFFSNRNX1_PCELL\%noxref_26 ( N_noxref_26_c_3271_n N_noxref_26_c_3273_n \
 N_noxref_26_c_3276_n N_noxref_26_c_3278_n N_noxref_26_c_3301_n \
 N_noxref_26_M16_noxref_d N_noxref_26_M17_noxref_s )  \
 PM_DFFSNRNX1_PCELL\%noxref_26
cc_1 ( N_noxref_1_c_1_p N_noxref_2_c_313_n ) capacitor c=0.00989031f //x=0.74 \
 //y=0 //x2=0.74 //y2=7.4
cc_2 ( N_noxref_1_c_2_p N_noxref_2_c_314_n ) capacitor c=0.00989031f //x=28.12 \
 //y=0 //x2=28.12 //y2=7.4
cc_3 ( N_noxref_1_c_3_p N_noxref_2_c_315_n ) capacitor c=0.00927471f //x=4.81 \
 //y=0 //x2=4.81 //y2=7.4
cc_4 ( N_noxref_1_c_4_p N_noxref_2_c_316_n ) capacitor c=0.00989031f //x=9.62 \
 //y=0 //x2=9.62 //y2=7.4
cc_5 ( N_noxref_1_c_5_p N_noxref_2_c_317_n ) capacitor c=0.00989031f //x=14.43 \
 //y=0 //x2=14.43 //y2=7.4
cc_6 ( N_noxref_1_c_6_p N_noxref_2_c_318_n ) capacitor c=0.00802221f //x=19.24 \
 //y=0 //x2=19.24 //y2=7.4
cc_7 ( N_noxref_1_c_7_p N_noxref_2_c_319_n ) capacitor c=0.00802221f //x=24.05 \
 //y=0 //x2=24.05 //y2=7.4
cc_8 ( N_noxref_1_c_3_p N_noxref_3_c_644_n ) capacitor c=0.0238274f //x=4.81 \
 //y=0 //x2=5.805 //y2=2.59
cc_9 ( N_noxref_1_c_3_p N_noxref_3_c_645_n ) capacitor c=0.00102529f //x=4.81 \
 //y=0 //x2=4.185 //y2=2.59
cc_10 ( N_noxref_1_c_4_p N_noxref_3_c_646_n ) capacitor c=0.0253329f //x=9.62 \
 //y=0 //x2=10.615 //y2=2.59
cc_11 ( N_noxref_1_c_3_p N_noxref_3_c_647_n ) capacitor c=7.16565e-19 //x=4.81 \
 //y=0 //x2=6.035 //y2=2.59
cc_12 ( N_noxref_1_c_3_p N_noxref_3_c_648_n ) capacitor c=0.04008f //x=4.81 \
 //y=0 //x2=3.985 //y2=1.665
cc_13 ( N_noxref_1_c_3_p N_noxref_3_c_649_n ) capacitor c=5.56859e-19 //x=4.81 \
 //y=0 //x2=4.07 //y2=2.59
cc_14 ( N_noxref_1_c_3_p N_noxref_3_c_650_n ) capacitor c=0.0128021f //x=4.81 \
 //y=0 //x2=5.92 //y2=2.08
cc_15 ( N_noxref_1_c_4_p N_noxref_3_c_651_n ) capacitor c=0.0126655f //x=9.62 \
 //y=0 //x2=10.73 //y2=2.08
cc_16 ( N_noxref_1_c_16_p N_noxref_3_c_652_n ) capacitor c=0.00132755f //x=5.8 \
 //y=0 //x2=5.62 //y2=0.875
cc_17 ( N_noxref_1_M3_noxref_d N_noxref_3_c_652_n ) capacitor c=0.00211996f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=0.875
cc_18 ( N_noxref_1_M3_noxref_d N_noxref_3_c_654_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=1.22
cc_19 ( N_noxref_1_c_3_p N_noxref_3_c_655_n ) capacitor c=0.00204716f //x=4.81 \
 //y=0 //x2=5.62 //y2=1.53
cc_20 ( N_noxref_1_c_3_p N_noxref_3_c_656_n ) capacitor c=0.0110952f //x=4.81 \
 //y=0 //x2=5.62 //y2=1.915
cc_21 ( N_noxref_1_M3_noxref_d N_noxref_3_c_657_n ) capacitor c=0.0131341f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=0.72
cc_22 ( N_noxref_1_M3_noxref_d N_noxref_3_c_658_n ) capacitor c=0.00193146f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=1.375
cc_23 ( N_noxref_1_c_23_p N_noxref_3_c_659_n ) capacitor c=0.00129018f \
 //x=9.45 //y=0 //x2=6.15 //y2=0.875
cc_24 ( N_noxref_1_M3_noxref_d N_noxref_3_c_659_n ) capacitor c=0.00257848f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=0.875
cc_25 ( N_noxref_1_M3_noxref_d N_noxref_3_c_661_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=1.22
cc_26 ( N_noxref_1_c_26_p N_noxref_3_c_662_n ) capacitor c=0.00132755f \
 //x=10.61 //y=0 //x2=10.43 //y2=0.875
cc_27 ( N_noxref_1_M6_noxref_d N_noxref_3_c_662_n ) capacitor c=0.00211996f \
 //x=10.505 //y=0.875 //x2=10.43 //y2=0.875
cc_28 ( N_noxref_1_M6_noxref_d N_noxref_3_c_664_n ) capacitor c=0.00255985f \
 //x=10.505 //y=0.875 //x2=10.43 //y2=1.22
cc_29 ( N_noxref_1_c_4_p N_noxref_3_c_665_n ) capacitor c=0.00204716f //x=9.62 \
 //y=0 //x2=10.43 //y2=1.53
cc_30 ( N_noxref_1_c_4_p N_noxref_3_c_666_n ) capacitor c=0.0112696f //x=9.62 \
 //y=0 //x2=10.43 //y2=1.915
cc_31 ( N_noxref_1_M6_noxref_d N_noxref_3_c_667_n ) capacitor c=0.0131341f \
 //x=10.505 //y=0.875 //x2=10.805 //y2=0.72
cc_32 ( N_noxref_1_M6_noxref_d N_noxref_3_c_668_n ) capacitor c=0.00193146f \
 //x=10.505 //y=0.875 //x2=10.805 //y2=1.375
cc_33 ( N_noxref_1_c_33_p N_noxref_3_c_669_n ) capacitor c=0.00129018f \
 //x=14.26 //y=0 //x2=10.96 //y2=0.875
cc_34 ( N_noxref_1_M6_noxref_d N_noxref_3_c_669_n ) capacitor c=0.00257848f \
 //x=10.505 //y=0.875 //x2=10.96 //y2=0.875
cc_35 ( N_noxref_1_M6_noxref_d N_noxref_3_c_671_n ) capacitor c=0.00255985f \
 //x=10.505 //y=0.875 //x2=10.96 //y2=1.22
cc_36 ( N_noxref_1_c_3_p N_noxref_3_M2_noxref_d ) capacitor c=0.00591582f \
 //x=4.81 //y=0 //x2=3.395 //y2=0.915
cc_37 ( N_noxref_1_c_5_p N_noxref_4_c_881_n ) capacitor c=0.0222748f //x=14.43 \
 //y=0 //x2=15.425 //y2=2.59
cc_38 ( N_noxref_1_c_5_p N_noxref_4_c_882_n ) capacitor c=0.00102529f \
 //x=14.43 //y=0 //x2=13.805 //y2=2.59
cc_39 ( N_noxref_1_c_5_p N_noxref_4_c_883_n ) capacitor c=0.0401826f //x=14.43 \
 //y=0 //x2=13.605 //y2=1.665
cc_40 ( N_noxref_1_c_5_p N_noxref_4_c_884_n ) capacitor c=5.56859e-19 \
 //x=14.43 //y=0 //x2=13.69 //y2=2.59
cc_41 ( N_noxref_1_c_5_p N_noxref_4_c_885_n ) capacitor c=0.0127664f //x=14.43 \
 //y=0 //x2=15.54 //y2=2.08
cc_42 ( N_noxref_1_c_42_p N_noxref_4_c_886_n ) capacitor c=0.00132755f \
 //x=15.42 //y=0 //x2=15.24 //y2=0.875
cc_43 ( N_noxref_1_M9_noxref_d N_noxref_4_c_886_n ) capacitor c=0.00211996f \
 //x=15.315 //y=0.875 //x2=15.24 //y2=0.875
cc_44 ( N_noxref_1_M9_noxref_d N_noxref_4_c_888_n ) capacitor c=0.00255985f \
 //x=15.315 //y=0.875 //x2=15.24 //y2=1.22
cc_45 ( N_noxref_1_c_5_p N_noxref_4_c_889_n ) capacitor c=0.00204716f \
 //x=14.43 //y=0 //x2=15.24 //y2=1.53
cc_46 ( N_noxref_1_c_5_p N_noxref_4_c_890_n ) capacitor c=0.0110952f //x=14.43 \
 //y=0 //x2=15.24 //y2=1.915
cc_47 ( N_noxref_1_M9_noxref_d N_noxref_4_c_891_n ) capacitor c=0.0131341f \
 //x=15.315 //y=0.875 //x2=15.615 //y2=0.72
cc_48 ( N_noxref_1_M9_noxref_d N_noxref_4_c_892_n ) capacitor c=0.00193146f \
 //x=15.315 //y=0.875 //x2=15.615 //y2=1.375
cc_49 ( N_noxref_1_c_49_p N_noxref_4_c_893_n ) capacitor c=0.00129018f \
 //x=19.07 //y=0 //x2=15.77 //y2=0.875
cc_50 ( N_noxref_1_M9_noxref_d N_noxref_4_c_893_n ) capacitor c=0.00257848f \
 //x=15.315 //y=0.875 //x2=15.77 //y2=0.875
cc_51 ( N_noxref_1_M9_noxref_d N_noxref_4_c_895_n ) capacitor c=0.00255985f \
 //x=15.315 //y=0.875 //x2=15.77 //y2=1.22
cc_52 ( N_noxref_1_c_5_p N_noxref_4_M8_noxref_d ) capacitor c=0.00591582f \
 //x=14.43 //y=0 //x2=13.015 //y2=0.915
cc_53 ( N_noxref_1_c_3_p N_noxref_5_c_1043_n ) capacitor c=5.58077e-19 \
 //x=4.81 //y=0 //x2=7.03 //y2=2.08
cc_54 ( N_noxref_1_c_5_p N_noxref_5_c_1044_n ) capacitor c=7.67786e-19 \
 //x=14.43 //y=0 //x2=16.65 //y2=2.08
cc_55 ( N_noxref_1_c_3_p N_noxref_6_c_1247_n ) capacitor c=0.00505527f \
 //x=4.81 //y=0 //x2=8.765 //y2=3.33
cc_56 ( N_noxref_1_c_4_p N_noxref_6_c_1248_n ) capacitor c=0.00505527f \
 //x=9.62 //y=0 //x2=20.235 //y2=3.33
cc_57 ( N_noxref_1_c_3_p N_noxref_6_c_1249_n ) capacitor c=0.00101012f \
 //x=4.81 //y=0 //x2=3.33 //y2=2.08
cc_58 ( N_noxref_1_c_4_p N_noxref_6_c_1250_n ) capacitor c=0.0405987f //x=9.62 \
 //y=0 //x2=8.795 //y2=1.665
cc_59 ( N_noxref_1_c_6_p N_noxref_6_c_1251_n ) capacitor c=0.0155796f \
 //x=19.24 //y=0 //x2=20.35 //y2=2.08
cc_60 ( N_noxref_1_c_60_p N_noxref_6_c_1252_n ) capacitor c=0.00132755f \
 //x=20.23 //y=0 //x2=20.05 //y2=0.875
cc_61 ( N_noxref_1_M12_noxref_d N_noxref_6_c_1252_n ) capacitor c=0.00211996f \
 //x=20.125 //y=0.875 //x2=20.05 //y2=0.875
cc_62 ( N_noxref_1_M12_noxref_d N_noxref_6_c_1254_n ) capacitor c=0.00255985f \
 //x=20.125 //y=0.875 //x2=20.05 //y2=1.22
cc_63 ( N_noxref_1_c_6_p N_noxref_6_c_1255_n ) capacitor c=0.00204716f \
 //x=19.24 //y=0 //x2=20.05 //y2=1.53
cc_64 ( N_noxref_1_c_6_p N_noxref_6_c_1256_n ) capacitor c=0.0110952f \
 //x=19.24 //y=0 //x2=20.05 //y2=1.915
cc_65 ( N_noxref_1_M12_noxref_d N_noxref_6_c_1257_n ) capacitor c=0.0131341f \
 //x=20.125 //y=0.875 //x2=20.425 //y2=0.72
cc_66 ( N_noxref_1_M12_noxref_d N_noxref_6_c_1258_n ) capacitor c=0.00193146f \
 //x=20.125 //y=0.875 //x2=20.425 //y2=1.375
cc_67 ( N_noxref_1_c_67_p N_noxref_6_c_1259_n ) capacitor c=0.00129018f \
 //x=23.88 //y=0 //x2=20.58 //y2=0.875
cc_68 ( N_noxref_1_M12_noxref_d N_noxref_6_c_1259_n ) capacitor c=0.00257848f \
 //x=20.125 //y=0.875 //x2=20.58 //y2=0.875
cc_69 ( N_noxref_1_M12_noxref_d N_noxref_6_c_1261_n ) capacitor c=0.00255985f \
 //x=20.125 //y=0.875 //x2=20.58 //y2=1.22
cc_70 ( N_noxref_1_c_4_p N_noxref_6_M5_noxref_d ) capacitor c=0.00591582f \
 //x=9.62 //y=0 //x2=8.205 //y2=0.915
cc_71 ( N_noxref_1_c_71_p N_noxref_7_c_1511_n ) capacitor c=0.145588f \
 //x=28.12 //y=0 //x2=17.645 //y2=2.22
cc_72 ( N_noxref_1_c_72_p N_noxref_7_c_1511_n ) capacitor c=0.00447829f \
 //x=4.64 //y=0 //x2=17.645 //y2=2.22
cc_73 ( N_noxref_1_c_16_p N_noxref_7_c_1511_n ) capacitor c=0.00274252f \
 //x=5.8 //y=0 //x2=17.645 //y2=2.22
cc_74 ( N_noxref_1_c_23_p N_noxref_7_c_1511_n ) capacitor c=0.00450506f \
 //x=9.45 //y=0 //x2=17.645 //y2=2.22
cc_75 ( N_noxref_1_c_26_p N_noxref_7_c_1511_n ) capacitor c=0.00274252f \
 //x=10.61 //y=0 //x2=17.645 //y2=2.22
cc_76 ( N_noxref_1_c_33_p N_noxref_7_c_1511_n ) capacitor c=0.00450506f \
 //x=14.26 //y=0 //x2=17.645 //y2=2.22
cc_77 ( N_noxref_1_c_42_p N_noxref_7_c_1511_n ) capacitor c=0.00274252f \
 //x=15.42 //y=0 //x2=17.645 //y2=2.22
cc_78 ( N_noxref_1_c_49_p N_noxref_7_c_1511_n ) capacitor c=0.00111309f \
 //x=19.07 //y=0 //x2=17.645 //y2=2.22
cc_79 ( N_noxref_1_c_3_p N_noxref_7_c_1511_n ) capacitor c=0.0379964f //x=4.81 \
 //y=0 //x2=17.645 //y2=2.22
cc_80 ( N_noxref_1_c_4_p N_noxref_7_c_1511_n ) capacitor c=0.0379964f //x=9.62 \
 //y=0 //x2=17.645 //y2=2.22
cc_81 ( N_noxref_1_c_5_p N_noxref_7_c_1511_n ) capacitor c=0.0379964f \
 //x=14.43 //y=0 //x2=17.645 //y2=2.22
cc_82 ( N_noxref_1_c_71_p N_noxref_7_c_1522_n ) capacitor c=0.0019104f \
 //x=28.12 //y=0 //x2=2.335 //y2=2.22
cc_83 ( N_noxref_1_c_71_p N_noxref_7_c_1523_n ) capacitor c=0.0355717f \
 //x=28.12 //y=0 //x2=21.345 //y2=2.22
cc_84 ( N_noxref_1_c_49_p N_noxref_7_c_1523_n ) capacitor c=0.00318526f \
 //x=19.07 //y=0 //x2=21.345 //y2=2.22
cc_85 ( N_noxref_1_c_60_p N_noxref_7_c_1523_n ) capacitor c=0.00274252f \
 //x=20.23 //y=0 //x2=21.345 //y2=2.22
cc_86 ( N_noxref_1_c_6_p N_noxref_7_c_1523_n ) capacitor c=0.0401775f \
 //x=19.24 //y=0 //x2=21.345 //y2=2.22
cc_87 ( N_noxref_1_c_71_p N_noxref_7_c_1527_n ) capacitor c=0.00195247f \
 //x=28.12 //y=0 //x2=17.875 //y2=2.22
cc_88 ( N_noxref_1_c_1_p N_noxref_7_c_1528_n ) capacitor c=8.20622e-19 \
 //x=0.74 //y=0 //x2=2.22 //y2=2.08
cc_89 ( N_noxref_1_c_6_p N_noxref_7_c_1529_n ) capacitor c=8.37259e-19 \
 //x=19.24 //y=0 //x2=17.76 //y2=2.08
cc_90 ( N_noxref_1_c_6_p N_noxref_7_c_1530_n ) capacitor c=5.94159e-19 \
 //x=19.24 //y=0 //x2=21.46 //y2=2.08
cc_91 ( N_noxref_1_c_71_p N_noxref_8_c_1827_n ) capacitor c=0.0528755f \
 //x=28.12 //y=0 //x2=26.155 //y2=2.96
cc_92 ( N_noxref_1_c_67_p N_noxref_8_c_1827_n ) capacitor c=0.00282695f \
 //x=23.88 //y=0 //x2=26.155 //y2=2.96
cc_93 ( N_noxref_1_c_93_p N_noxref_8_c_1827_n ) capacitor c=0.00184476f \
 //x=25.04 //y=0 //x2=26.155 //y2=2.96
cc_94 ( N_noxref_1_c_5_p N_noxref_8_c_1827_n ) capacitor c=0.00750857f \
 //x=14.43 //y=0 //x2=26.155 //y2=2.96
cc_95 ( N_noxref_1_c_6_p N_noxref_8_c_1827_n ) capacitor c=0.00949826f \
 //x=19.24 //y=0 //x2=26.155 //y2=2.96
cc_96 ( N_noxref_1_c_7_p N_noxref_8_c_1827_n ) capacitor c=0.0144849f \
 //x=24.05 //y=0 //x2=26.155 //y2=2.96
cc_97 ( N_noxref_1_c_4_p N_noxref_8_c_1833_n ) capacitor c=7.37634e-19 \
 //x=9.62 //y=0 //x2=11.84 //y2=2.08
cc_98 ( N_noxref_1_c_7_p N_noxref_8_c_1834_n ) capacitor c=7.64246e-19 \
 //x=24.05 //y=0 //x2=26.27 //y2=2.08
cc_99 ( N_noxref_1_c_71_p N_noxref_9_c_2028_n ) capacitor c=0.0159588f \
 //x=28.12 //y=0 //x2=27.265 //y2=3.7
cc_100 ( N_noxref_1_c_4_p N_noxref_9_c_2029_n ) capacitor c=6.0472e-19 \
 //x=9.62 //y=0 //x2=8.14 //y2=2.08
cc_101 ( N_noxref_1_c_5_p N_noxref_9_c_2030_n ) capacitor c=9.24123e-19 \
 //x=14.43 //y=0 //x2=12.95 //y2=2.08
cc_102 ( N_noxref_1_c_6_p N_noxref_9_c_2031_n ) capacitor c=0.0430857f \
 //x=19.24 //y=0 //x2=18.415 //y2=1.665
cc_103 ( N_noxref_1_c_2_p N_noxref_9_c_2032_n ) capacitor c=9.53263e-19 \
 //x=28.12 //y=0 //x2=27.38 //y2=2.08
cc_104 ( N_noxref_1_c_6_p N_noxref_9_M11_noxref_d ) capacitor c=0.00591582f \
 //x=19.24 //y=0 //x2=17.825 //y2=0.915
cc_105 ( N_noxref_1_c_1_p N_noxref_10_c_2364_n ) capacitor c=0.0178706f \
 //x=0.74 //y=0 //x2=1.11 //y2=2.08
cc_106 ( N_noxref_1_c_106_p N_noxref_10_c_2365_n ) capacitor c=0.00132755f \
 //x=0.99 //y=0 //x2=0.81 //y2=0.875
cc_107 ( N_noxref_1_M0_noxref_d N_noxref_10_c_2365_n ) capacitor c=0.00211996f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=0.875
cc_108 ( N_noxref_1_M0_noxref_d N_noxref_10_c_2367_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=1.22
cc_109 ( N_noxref_1_c_1_p N_noxref_10_c_2368_n ) capacitor c=0.00295461f \
 //x=0.74 //y=0 //x2=0.81 //y2=1.53
cc_110 ( N_noxref_1_c_1_p N_noxref_10_c_2369_n ) capacitor c=0.0126075f \
 //x=0.74 //y=0 //x2=0.81 //y2=1.915
cc_111 ( N_noxref_1_M0_noxref_d N_noxref_10_c_2370_n ) capacitor c=0.0131341f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=0.72
cc_112 ( N_noxref_1_M0_noxref_d N_noxref_10_c_2371_n ) capacitor c=0.00193146f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=1.375
cc_113 ( N_noxref_1_c_72_p N_noxref_10_c_2372_n ) capacitor c=0.00129018f \
 //x=4.64 //y=0 //x2=1.34 //y2=0.875
cc_114 ( N_noxref_1_M0_noxref_d N_noxref_10_c_2372_n ) capacitor c=0.00257848f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=0.875
cc_115 ( N_noxref_1_M0_noxref_d N_noxref_10_c_2374_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=1.22
cc_116 ( N_noxref_1_c_71_p N_noxref_11_c_2421_n ) capacitor c=0.00710541f \
 //x=28.12 //y=0 //x2=1.475 //y2=1.59
cc_117 ( N_noxref_1_c_106_p N_noxref_11_c_2421_n ) capacitor c=0.00110021f \
 //x=0.99 //y=0 //x2=1.475 //y2=1.59
cc_118 ( N_noxref_1_c_72_p N_noxref_11_c_2421_n ) capacitor c=0.00179185f \
 //x=4.64 //y=0 //x2=1.475 //y2=1.59
cc_119 ( N_noxref_1_M0_noxref_d N_noxref_11_c_2421_n ) capacitor c=0.00900091f \
 //x=0.885 //y=0.875 //x2=1.475 //y2=1.59
cc_120 ( N_noxref_1_c_71_p N_noxref_11_c_2425_n ) capacitor c=0.00709506f \
 //x=28.12 //y=0 //x2=1.56 //y2=0.625
cc_121 ( N_noxref_1_c_72_p N_noxref_11_c_2425_n ) capacitor c=0.0140218f \
 //x=4.64 //y=0 //x2=1.56 //y2=0.625
cc_122 ( N_noxref_1_M0_noxref_d N_noxref_11_c_2425_n ) capacitor c=0.033954f \
 //x=0.885 //y=0.875 //x2=1.56 //y2=0.625
cc_123 ( N_noxref_1_c_71_p N_noxref_11_c_2428_n ) capacitor c=0.0151387f \
 //x=28.12 //y=0 //x2=2.445 //y2=0.54
cc_124 ( N_noxref_1_c_72_p N_noxref_11_c_2428_n ) capacitor c=0.0358309f \
 //x=4.64 //y=0 //x2=2.445 //y2=0.54
cc_125 ( N_noxref_1_c_2_p N_noxref_11_c_2428_n ) capacitor c=0.00265129f \
 //x=28.12 //y=0 //x2=2.445 //y2=0.54
cc_126 ( N_noxref_1_c_71_p N_noxref_11_M0_noxref_s ) capacitor c=0.00962687f \
 //x=28.12 //y=0 //x2=0.455 //y2=0.375
cc_127 ( N_noxref_1_c_106_p N_noxref_11_M0_noxref_s ) capacitor c=0.0140218f \
 //x=0.99 //y=0 //x2=0.455 //y2=0.375
cc_128 ( N_noxref_1_c_1_p N_noxref_11_M0_noxref_s ) capacitor c=0.0712607f \
 //x=0.74 //y=0 //x2=0.455 //y2=0.375
cc_129 ( N_noxref_1_c_72_p N_noxref_11_M0_noxref_s ) capacitor c=0.0131437f \
 //x=4.64 //y=0 //x2=0.455 //y2=0.375
cc_130 ( N_noxref_1_c_3_p N_noxref_11_M0_noxref_s ) capacitor c=3.31601e-19 \
 //x=4.81 //y=0 //x2=0.455 //y2=0.375
cc_131 ( N_noxref_1_M0_noxref_d N_noxref_11_M0_noxref_s ) capacitor \
 c=0.033718f //x=0.885 //y=0.875 //x2=0.455 //y2=0.375
cc_132 ( N_noxref_1_c_71_p N_noxref_12_c_2467_n ) capacitor c=0.00352952f \
 //x=28.12 //y=0 //x2=3.015 //y2=0.995
cc_133 ( N_noxref_1_c_72_p N_noxref_12_c_2467_n ) capacitor c=0.00934524f \
 //x=4.64 //y=0 //x2=3.015 //y2=0.995
cc_134 ( N_noxref_1_c_2_p N_noxref_12_c_2467_n ) capacitor c=3.54249e-19 \
 //x=28.12 //y=0 //x2=3.015 //y2=0.995
cc_135 ( N_noxref_1_c_71_p N_noxref_12_c_2470_n ) capacitor c=0.00254475f \
 //x=28.12 //y=0 //x2=3.1 //y2=0.625
cc_136 ( N_noxref_1_c_72_p N_noxref_12_c_2470_n ) capacitor c=0.0140928f \
 //x=4.64 //y=0 //x2=3.1 //y2=0.625
cc_137 ( N_noxref_1_M0_noxref_d N_noxref_12_c_2470_n ) capacitor c=6.21394e-19 \
 //x=0.885 //y=0.875 //x2=3.1 //y2=0.625
cc_138 ( N_noxref_1_c_71_p N_noxref_12_c_2473_n ) capacitor c=0.0105317f \
 //x=28.12 //y=0 //x2=3.985 //y2=0.54
cc_139 ( N_noxref_1_c_72_p N_noxref_12_c_2473_n ) capacitor c=0.0363691f \
 //x=4.64 //y=0 //x2=3.985 //y2=0.54
cc_140 ( N_noxref_1_c_2_p N_noxref_12_c_2473_n ) capacitor c=0.00283214f \
 //x=28.12 //y=0 //x2=3.985 //y2=0.54
cc_141 ( N_noxref_1_c_71_p N_noxref_12_c_2476_n ) capacitor c=0.00254232f \
 //x=28.12 //y=0 //x2=4.07 //y2=0.625
cc_142 ( N_noxref_1_c_72_p N_noxref_12_c_2476_n ) capacitor c=0.0140304f \
 //x=4.64 //y=0 //x2=4.07 //y2=0.625
cc_143 ( N_noxref_1_c_3_p N_noxref_12_c_2476_n ) capacitor c=0.0404137f \
 //x=4.81 //y=0 //x2=4.07 //y2=0.625
cc_144 ( N_noxref_1_M0_noxref_d N_noxref_12_M1_noxref_d ) capacitor \
 c=0.00162435f //x=0.885 //y=0.875 //x2=1.86 //y2=0.91
cc_145 ( N_noxref_1_c_1_p N_noxref_12_M2_noxref_s ) capacitor c=8.16352e-19 \
 //x=0.74 //y=0 //x2=2.965 //y2=0.375
cc_146 ( N_noxref_1_c_3_p N_noxref_12_M2_noxref_s ) capacitor c=0.00183204f \
 //x=4.81 //y=0 //x2=2.965 //y2=0.375
cc_147 ( N_noxref_1_c_71_p N_noxref_13_c_2521_n ) capacitor c=0.00517576f \
 //x=28.12 //y=0 //x2=6.285 //y2=1.59
cc_148 ( N_noxref_1_c_16_p N_noxref_13_c_2521_n ) capacitor c=0.00111448f \
 //x=5.8 //y=0 //x2=6.285 //y2=1.59
cc_149 ( N_noxref_1_c_23_p N_noxref_13_c_2521_n ) capacitor c=0.00180612f \
 //x=9.45 //y=0 //x2=6.285 //y2=1.59
cc_150 ( N_noxref_1_M3_noxref_d N_noxref_13_c_2521_n ) capacitor c=0.00853078f \
 //x=5.695 //y=0.875 //x2=6.285 //y2=1.59
cc_151 ( N_noxref_1_c_71_p N_noxref_13_c_2525_n ) capacitor c=0.00254475f \
 //x=28.12 //y=0 //x2=6.37 //y2=0.625
cc_152 ( N_noxref_1_c_23_p N_noxref_13_c_2525_n ) capacitor c=0.0140928f \
 //x=9.45 //y=0 //x2=6.37 //y2=0.625
cc_153 ( N_noxref_1_M3_noxref_d N_noxref_13_c_2525_n ) capacitor c=0.033954f \
 //x=5.695 //y=0.875 //x2=6.37 //y2=0.625
cc_154 ( N_noxref_1_c_71_p N_noxref_13_c_2528_n ) capacitor c=0.0104506f \
 //x=28.12 //y=0 //x2=7.255 //y2=0.54
cc_155 ( N_noxref_1_c_23_p N_noxref_13_c_2528_n ) capacitor c=0.0360726f \
 //x=9.45 //y=0 //x2=7.255 //y2=0.54
cc_156 ( N_noxref_1_c_2_p N_noxref_13_c_2528_n ) capacitor c=0.00265129f \
 //x=28.12 //y=0 //x2=7.255 //y2=0.54
cc_157 ( N_noxref_1_c_71_p N_noxref_13_M3_noxref_s ) capacitor c=0.00507657f \
 //x=28.12 //y=0 //x2=5.265 //y2=0.375
cc_158 ( N_noxref_1_c_16_p N_noxref_13_M3_noxref_s ) capacitor c=0.0140928f \
 //x=5.8 //y=0 //x2=5.265 //y2=0.375
cc_159 ( N_noxref_1_c_23_p N_noxref_13_M3_noxref_s ) capacitor c=0.0136651f \
 //x=9.45 //y=0 //x2=5.265 //y2=0.375
cc_160 ( N_noxref_1_c_3_p N_noxref_13_M3_noxref_s ) capacitor c=0.0696963f \
 //x=4.81 //y=0 //x2=5.265 //y2=0.375
cc_161 ( N_noxref_1_c_4_p N_noxref_13_M3_noxref_s ) capacitor c=3.31601e-19 \
 //x=9.62 //y=0 //x2=5.265 //y2=0.375
cc_162 ( N_noxref_1_M3_noxref_d N_noxref_13_M3_noxref_s ) capacitor \
 c=0.033718f //x=5.695 //y=0.875 //x2=5.265 //y2=0.375
cc_163 ( N_noxref_1_c_71_p N_noxref_14_c_2571_n ) capacitor c=0.00352952f \
 //x=28.12 //y=0 //x2=7.825 //y2=0.995
cc_164 ( N_noxref_1_c_23_p N_noxref_14_c_2571_n ) capacitor c=0.00934524f \
 //x=9.45 //y=0 //x2=7.825 //y2=0.995
cc_165 ( N_noxref_1_c_2_p N_noxref_14_c_2571_n ) capacitor c=3.54249e-19 \
 //x=28.12 //y=0 //x2=7.825 //y2=0.995
cc_166 ( N_noxref_1_c_71_p N_noxref_14_c_2574_n ) capacitor c=0.00254475f \
 //x=28.12 //y=0 //x2=7.91 //y2=0.625
cc_167 ( N_noxref_1_c_23_p N_noxref_14_c_2574_n ) capacitor c=0.0140928f \
 //x=9.45 //y=0 //x2=7.91 //y2=0.625
cc_168 ( N_noxref_1_M3_noxref_d N_noxref_14_c_2574_n ) capacitor c=6.21394e-19 \
 //x=5.695 //y=0.875 //x2=7.91 //y2=0.625
cc_169 ( N_noxref_1_c_71_p N_noxref_14_c_2577_n ) capacitor c=0.0105317f \
 //x=28.12 //y=0 //x2=8.795 //y2=0.54
cc_170 ( N_noxref_1_c_23_p N_noxref_14_c_2577_n ) capacitor c=0.0364215f \
 //x=9.45 //y=0 //x2=8.795 //y2=0.54
cc_171 ( N_noxref_1_c_2_p N_noxref_14_c_2577_n ) capacitor c=0.00283214f \
 //x=28.12 //y=0 //x2=8.795 //y2=0.54
cc_172 ( N_noxref_1_c_71_p N_noxref_14_c_2580_n ) capacitor c=0.00254232f \
 //x=28.12 //y=0 //x2=8.88 //y2=0.625
cc_173 ( N_noxref_1_c_23_p N_noxref_14_c_2580_n ) capacitor c=0.0140304f \
 //x=9.45 //y=0 //x2=8.88 //y2=0.625
cc_174 ( N_noxref_1_c_4_p N_noxref_14_c_2580_n ) capacitor c=0.0404137f \
 //x=9.62 //y=0 //x2=8.88 //y2=0.625
cc_175 ( N_noxref_1_M3_noxref_d N_noxref_14_M4_noxref_d ) capacitor \
 c=0.00162435f //x=5.695 //y=0.875 //x2=6.67 //y2=0.91
cc_176 ( N_noxref_1_c_3_p N_noxref_14_M5_noxref_s ) capacitor c=8.16352e-19 \
 //x=4.81 //y=0 //x2=7.775 //y2=0.375
cc_177 ( N_noxref_1_c_4_p N_noxref_14_M5_noxref_s ) capacitor c=0.00183204f \
 //x=9.62 //y=0 //x2=7.775 //y2=0.375
cc_178 ( N_noxref_1_c_71_p N_noxref_15_c_2625_n ) capacitor c=0.00517576f \
 //x=28.12 //y=0 //x2=11.095 //y2=1.59
cc_179 ( N_noxref_1_c_26_p N_noxref_15_c_2625_n ) capacitor c=0.00111448f \
 //x=10.61 //y=0 //x2=11.095 //y2=1.59
cc_180 ( N_noxref_1_c_33_p N_noxref_15_c_2625_n ) capacitor c=0.00180612f \
 //x=14.26 //y=0 //x2=11.095 //y2=1.59
cc_181 ( N_noxref_1_M6_noxref_d N_noxref_15_c_2625_n ) capacitor c=0.00853078f \
 //x=10.505 //y=0.875 //x2=11.095 //y2=1.59
cc_182 ( N_noxref_1_c_71_p N_noxref_15_c_2629_n ) capacitor c=0.00254475f \
 //x=28.12 //y=0 //x2=11.18 //y2=0.625
cc_183 ( N_noxref_1_c_33_p N_noxref_15_c_2629_n ) capacitor c=0.0140928f \
 //x=14.26 //y=0 //x2=11.18 //y2=0.625
cc_184 ( N_noxref_1_M6_noxref_d N_noxref_15_c_2629_n ) capacitor c=0.033954f \
 //x=10.505 //y=0.875 //x2=11.18 //y2=0.625
cc_185 ( N_noxref_1_c_71_p N_noxref_15_c_2632_n ) capacitor c=0.0104506f \
 //x=28.12 //y=0 //x2=12.065 //y2=0.54
cc_186 ( N_noxref_1_c_33_p N_noxref_15_c_2632_n ) capacitor c=0.0360726f \
 //x=14.26 //y=0 //x2=12.065 //y2=0.54
cc_187 ( N_noxref_1_c_2_p N_noxref_15_c_2632_n ) capacitor c=0.00265129f \
 //x=28.12 //y=0 //x2=12.065 //y2=0.54
cc_188 ( N_noxref_1_c_71_p N_noxref_15_M6_noxref_s ) capacitor c=0.00507657f \
 //x=28.12 //y=0 //x2=10.075 //y2=0.375
cc_189 ( N_noxref_1_c_26_p N_noxref_15_M6_noxref_s ) capacitor c=0.0140928f \
 //x=10.61 //y=0 //x2=10.075 //y2=0.375
cc_190 ( N_noxref_1_c_33_p N_noxref_15_M6_noxref_s ) capacitor c=0.0131437f \
 //x=14.26 //y=0 //x2=10.075 //y2=0.375
cc_191 ( N_noxref_1_c_4_p N_noxref_15_M6_noxref_s ) capacitor c=0.0696963f \
 //x=9.62 //y=0 //x2=10.075 //y2=0.375
cc_192 ( N_noxref_1_c_5_p N_noxref_15_M6_noxref_s ) capacitor c=3.31601e-19 \
 //x=14.43 //y=0 //x2=10.075 //y2=0.375
cc_193 ( N_noxref_1_M6_noxref_d N_noxref_15_M6_noxref_s ) capacitor \
 c=0.033718f //x=10.505 //y=0.875 //x2=10.075 //y2=0.375
cc_194 ( N_noxref_1_c_71_p N_noxref_16_c_2675_n ) capacitor c=0.00352952f \
 //x=28.12 //y=0 //x2=12.635 //y2=0.995
cc_195 ( N_noxref_1_c_33_p N_noxref_16_c_2675_n ) capacitor c=0.00934524f \
 //x=14.26 //y=0 //x2=12.635 //y2=0.995
cc_196 ( N_noxref_1_c_2_p N_noxref_16_c_2675_n ) capacitor c=3.54249e-19 \
 //x=28.12 //y=0 //x2=12.635 //y2=0.995
cc_197 ( N_noxref_1_c_71_p N_noxref_16_c_2678_n ) capacitor c=0.00254475f \
 //x=28.12 //y=0 //x2=12.72 //y2=0.625
cc_198 ( N_noxref_1_c_33_p N_noxref_16_c_2678_n ) capacitor c=0.0140928f \
 //x=14.26 //y=0 //x2=12.72 //y2=0.625
cc_199 ( N_noxref_1_M6_noxref_d N_noxref_16_c_2678_n ) capacitor c=6.21394e-19 \
 //x=10.505 //y=0.875 //x2=12.72 //y2=0.625
cc_200 ( N_noxref_1_c_71_p N_noxref_16_c_2681_n ) capacitor c=0.0105317f \
 //x=28.12 //y=0 //x2=13.605 //y2=0.54
cc_201 ( N_noxref_1_c_33_p N_noxref_16_c_2681_n ) capacitor c=0.0364215f \
 //x=14.26 //y=0 //x2=13.605 //y2=0.54
cc_202 ( N_noxref_1_c_2_p N_noxref_16_c_2681_n ) capacitor c=0.00283214f \
 //x=28.12 //y=0 //x2=13.605 //y2=0.54
cc_203 ( N_noxref_1_c_71_p N_noxref_16_c_2684_n ) capacitor c=0.00254232f \
 //x=28.12 //y=0 //x2=13.69 //y2=0.625
cc_204 ( N_noxref_1_c_33_p N_noxref_16_c_2684_n ) capacitor c=0.0140304f \
 //x=14.26 //y=0 //x2=13.69 //y2=0.625
cc_205 ( N_noxref_1_c_5_p N_noxref_16_c_2684_n ) capacitor c=0.0404137f \
 //x=14.43 //y=0 //x2=13.69 //y2=0.625
cc_206 ( N_noxref_1_M6_noxref_d N_noxref_16_M7_noxref_d ) capacitor \
 c=0.00162435f //x=10.505 //y=0.875 //x2=11.48 //y2=0.91
cc_207 ( N_noxref_1_c_4_p N_noxref_16_M8_noxref_s ) capacitor c=8.16352e-19 \
 //x=9.62 //y=0 //x2=12.585 //y2=0.375
cc_208 ( N_noxref_1_c_5_p N_noxref_16_M8_noxref_s ) capacitor c=0.00183204f \
 //x=14.43 //y=0 //x2=12.585 //y2=0.375
cc_209 ( N_noxref_1_c_71_p N_noxref_17_c_2729_n ) capacitor c=0.00517576f \
 //x=28.12 //y=0 //x2=15.905 //y2=1.59
cc_210 ( N_noxref_1_c_42_p N_noxref_17_c_2729_n ) capacitor c=0.00111448f \
 //x=15.42 //y=0 //x2=15.905 //y2=1.59
cc_211 ( N_noxref_1_c_49_p N_noxref_17_c_2729_n ) capacitor c=0.00180612f \
 //x=19.07 //y=0 //x2=15.905 //y2=1.59
cc_212 ( N_noxref_1_M9_noxref_d N_noxref_17_c_2729_n ) capacitor c=0.00853078f \
 //x=15.315 //y=0.875 //x2=15.905 //y2=1.59
cc_213 ( N_noxref_1_c_71_p N_noxref_17_c_2733_n ) capacitor c=0.00254475f \
 //x=28.12 //y=0 //x2=15.99 //y2=0.625
cc_214 ( N_noxref_1_c_49_p N_noxref_17_c_2733_n ) capacitor c=0.0140928f \
 //x=19.07 //y=0 //x2=15.99 //y2=0.625
cc_215 ( N_noxref_1_M9_noxref_d N_noxref_17_c_2733_n ) capacitor c=0.033954f \
 //x=15.315 //y=0.875 //x2=15.99 //y2=0.625
cc_216 ( N_noxref_1_c_71_p N_noxref_17_c_2736_n ) capacitor c=0.0104506f \
 //x=28.12 //y=0 //x2=16.875 //y2=0.54
cc_217 ( N_noxref_1_c_49_p N_noxref_17_c_2736_n ) capacitor c=0.0360726f \
 //x=19.07 //y=0 //x2=16.875 //y2=0.54
cc_218 ( N_noxref_1_c_2_p N_noxref_17_c_2736_n ) capacitor c=0.00265129f \
 //x=28.12 //y=0 //x2=16.875 //y2=0.54
cc_219 ( N_noxref_1_c_71_p N_noxref_17_M9_noxref_s ) capacitor c=0.00507657f \
 //x=28.12 //y=0 //x2=14.885 //y2=0.375
cc_220 ( N_noxref_1_c_42_p N_noxref_17_M9_noxref_s ) capacitor c=0.0140928f \
 //x=15.42 //y=0 //x2=14.885 //y2=0.375
cc_221 ( N_noxref_1_c_49_p N_noxref_17_M9_noxref_s ) capacitor c=0.0131437f \
 //x=19.07 //y=0 //x2=14.885 //y2=0.375
cc_222 ( N_noxref_1_c_5_p N_noxref_17_M9_noxref_s ) capacitor c=0.0696963f \
 //x=14.43 //y=0 //x2=14.885 //y2=0.375
cc_223 ( N_noxref_1_c_6_p N_noxref_17_M9_noxref_s ) capacitor c=3.31601e-19 \
 //x=19.24 //y=0 //x2=14.885 //y2=0.375
cc_224 ( N_noxref_1_M9_noxref_d N_noxref_17_M9_noxref_s ) capacitor \
 c=0.033718f //x=15.315 //y=0.875 //x2=14.885 //y2=0.375
cc_225 ( N_noxref_1_c_71_p N_noxref_18_c_2779_n ) capacitor c=0.00352952f \
 //x=28.12 //y=0 //x2=17.445 //y2=0.995
cc_226 ( N_noxref_1_c_49_p N_noxref_18_c_2779_n ) capacitor c=0.00934524f \
 //x=19.07 //y=0 //x2=17.445 //y2=0.995
cc_227 ( N_noxref_1_c_2_p N_noxref_18_c_2779_n ) capacitor c=3.54249e-19 \
 //x=28.12 //y=0 //x2=17.445 //y2=0.995
cc_228 ( N_noxref_1_c_71_p N_noxref_18_c_2782_n ) capacitor c=0.00254475f \
 //x=28.12 //y=0 //x2=17.53 //y2=0.625
cc_229 ( N_noxref_1_c_49_p N_noxref_18_c_2782_n ) capacitor c=0.0140928f \
 //x=19.07 //y=0 //x2=17.53 //y2=0.625
cc_230 ( N_noxref_1_M9_noxref_d N_noxref_18_c_2782_n ) capacitor c=6.21394e-19 \
 //x=15.315 //y=0.875 //x2=17.53 //y2=0.625
cc_231 ( N_noxref_1_c_71_p N_noxref_18_c_2785_n ) capacitor c=0.0105197f \
 //x=28.12 //y=0 //x2=18.415 //y2=0.54
cc_232 ( N_noxref_1_c_49_p N_noxref_18_c_2785_n ) capacitor c=0.0364139f \
 //x=19.07 //y=0 //x2=18.415 //y2=0.54
cc_233 ( N_noxref_1_c_2_p N_noxref_18_c_2785_n ) capacitor c=0.00283214f \
 //x=28.12 //y=0 //x2=18.415 //y2=0.54
cc_234 ( N_noxref_1_c_71_p N_noxref_18_c_2788_n ) capacitor c=0.00254232f \
 //x=28.12 //y=0 //x2=18.5 //y2=0.625
cc_235 ( N_noxref_1_c_49_p N_noxref_18_c_2788_n ) capacitor c=0.0140304f \
 //x=19.07 //y=0 //x2=18.5 //y2=0.625
cc_236 ( N_noxref_1_c_6_p N_noxref_18_c_2788_n ) capacitor c=0.0404137f \
 //x=19.24 //y=0 //x2=18.5 //y2=0.625
cc_237 ( N_noxref_1_M9_noxref_d N_noxref_18_M10_noxref_d ) capacitor \
 c=0.00162435f //x=15.315 //y=0.875 //x2=16.29 //y2=0.91
cc_238 ( N_noxref_1_c_5_p N_noxref_18_M11_noxref_s ) capacitor c=8.16352e-19 \
 //x=14.43 //y=0 //x2=17.395 //y2=0.375
cc_239 ( N_noxref_1_c_6_p N_noxref_18_M11_noxref_s ) capacitor c=0.00183204f \
 //x=19.24 //y=0 //x2=17.395 //y2=0.375
cc_240 ( N_noxref_1_c_71_p N_noxref_19_c_2834_n ) capacitor c=0.00517576f \
 //x=28.12 //y=0 //x2=20.715 //y2=1.59
cc_241 ( N_noxref_1_c_60_p N_noxref_19_c_2834_n ) capacitor c=0.00111448f \
 //x=20.23 //y=0 //x2=20.715 //y2=1.59
cc_242 ( N_noxref_1_c_67_p N_noxref_19_c_2834_n ) capacitor c=0.00180612f \
 //x=23.88 //y=0 //x2=20.715 //y2=1.59
cc_243 ( N_noxref_1_M12_noxref_d N_noxref_19_c_2834_n ) capacitor \
 c=0.00853078f //x=20.125 //y=0.875 //x2=20.715 //y2=1.59
cc_244 ( N_noxref_1_c_71_p N_noxref_19_c_2838_n ) capacitor c=0.00254475f \
 //x=28.12 //y=0 //x2=20.8 //y2=0.625
cc_245 ( N_noxref_1_c_67_p N_noxref_19_c_2838_n ) capacitor c=0.0140928f \
 //x=23.88 //y=0 //x2=20.8 //y2=0.625
cc_246 ( N_noxref_1_M12_noxref_d N_noxref_19_c_2838_n ) capacitor c=0.033954f \
 //x=20.125 //y=0.875 //x2=20.8 //y2=0.625
cc_247 ( N_noxref_1_c_71_p N_noxref_19_c_2841_n ) capacitor c=0.0105304f \
 //x=28.12 //y=0 //x2=21.685 //y2=0.54
cc_248 ( N_noxref_1_c_67_p N_noxref_19_c_2841_n ) capacitor c=0.0361183f \
 //x=23.88 //y=0 //x2=21.685 //y2=0.54
cc_249 ( N_noxref_1_c_2_p N_noxref_19_c_2841_n ) capacitor c=0.00265129f \
 //x=28.12 //y=0 //x2=21.685 //y2=0.54
cc_250 ( N_noxref_1_c_71_p N_noxref_19_M12_noxref_s ) capacitor c=0.00531539f \
 //x=28.12 //y=0 //x2=19.695 //y2=0.375
cc_251 ( N_noxref_1_c_60_p N_noxref_19_M12_noxref_s ) capacitor c=0.0140928f \
 //x=20.23 //y=0 //x2=19.695 //y2=0.375
cc_252 ( N_noxref_1_c_67_p N_noxref_19_M12_noxref_s ) capacitor c=0.0133155f \
 //x=23.88 //y=0 //x2=19.695 //y2=0.375
cc_253 ( N_noxref_1_c_6_p N_noxref_19_M12_noxref_s ) capacitor c=0.0696963f \
 //x=19.24 //y=0 //x2=19.695 //y2=0.375
cc_254 ( N_noxref_1_c_7_p N_noxref_19_M12_noxref_s ) capacitor c=3.31601e-19 \
 //x=24.05 //y=0 //x2=19.695 //y2=0.375
cc_255 ( N_noxref_1_M12_noxref_d N_noxref_19_M12_noxref_s ) capacitor \
 c=0.033718f //x=20.125 //y=0.875 //x2=19.695 //y2=0.375
cc_256 ( N_noxref_1_c_7_p N_noxref_20_c_2886_n ) capacitor c=0.00128267f \
 //x=24.05 //y=0 //x2=22.57 //y2=2.08
cc_257 ( N_noxref_1_c_7_p N_noxref_21_c_2945_n ) capacitor c=0.045554f \
 //x=24.05 //y=0 //x2=23.225 //y2=1.665
cc_258 ( N_noxref_1_c_7_p N_noxref_21_M14_noxref_d ) capacitor c=0.00591582f \
 //x=24.05 //y=0 //x2=22.635 //y2=0.915
cc_259 ( N_noxref_1_c_71_p N_noxref_22_c_3029_n ) capacitor c=0.00375441f \
 //x=28.12 //y=0 //x2=22.255 //y2=0.995
cc_260 ( N_noxref_1_c_67_p N_noxref_22_c_3029_n ) capacitor c=0.00944862f \
 //x=23.88 //y=0 //x2=22.255 //y2=0.995
cc_261 ( N_noxref_1_c_2_p N_noxref_22_c_3029_n ) capacitor c=3.54249e-19 \
 //x=28.12 //y=0 //x2=22.255 //y2=0.995
cc_262 ( N_noxref_1_c_71_p N_noxref_22_c_3032_n ) capacitor c=0.00277579f \
 //x=28.12 //y=0 //x2=22.34 //y2=0.625
cc_263 ( N_noxref_1_c_67_p N_noxref_22_c_3032_n ) capacitor c=0.0142586f \
 //x=23.88 //y=0 //x2=22.34 //y2=0.625
cc_264 ( N_noxref_1_M12_noxref_d N_noxref_22_c_3032_n ) capacitor \
 c=6.21394e-19 //x=20.125 //y=0.875 //x2=22.34 //y2=0.625
cc_265 ( N_noxref_1_c_71_p N_noxref_22_c_3035_n ) capacitor c=0.011473f \
 //x=28.12 //y=0 //x2=23.225 //y2=0.54
cc_266 ( N_noxref_1_c_67_p N_noxref_22_c_3035_n ) capacitor c=0.0365589f \
 //x=23.88 //y=0 //x2=23.225 //y2=0.54
cc_267 ( N_noxref_1_c_2_p N_noxref_22_c_3035_n ) capacitor c=0.00283214f \
 //x=28.12 //y=0 //x2=23.225 //y2=0.54
cc_268 ( N_noxref_1_c_71_p N_noxref_22_c_3038_n ) capacitor c=0.00277442f \
 //x=28.12 //y=0 //x2=23.31 //y2=0.625
cc_269 ( N_noxref_1_c_67_p N_noxref_22_c_3038_n ) capacitor c=0.014197f \
 //x=23.88 //y=0 //x2=23.31 //y2=0.625
cc_270 ( N_noxref_1_c_7_p N_noxref_22_c_3038_n ) capacitor c=0.0404137f \
 //x=24.05 //y=0 //x2=23.31 //y2=0.625
cc_271 ( N_noxref_1_M12_noxref_d N_noxref_22_M13_noxref_d ) capacitor \
 c=0.00162435f //x=20.125 //y=0.875 //x2=21.1 //y2=0.91
cc_272 ( N_noxref_1_c_6_p N_noxref_22_M14_noxref_s ) capacitor c=8.16352e-19 \
 //x=19.24 //y=0 //x2=22.205 //y2=0.375
cc_273 ( N_noxref_1_c_7_p N_noxref_22_M14_noxref_s ) capacitor c=0.00183204f \
 //x=24.05 //y=0 //x2=22.205 //y2=0.375
cc_274 ( N_noxref_1_c_7_p N_noxref_23_c_3083_n ) capacitor c=0.0179249f \
 //x=24.05 //y=0 //x2=25.16 //y2=2.08
cc_275 ( N_noxref_1_c_93_p N_noxref_23_c_3084_n ) capacitor c=0.00132755f \
 //x=25.04 //y=0 //x2=24.86 //y2=0.875
cc_276 ( N_noxref_1_M15_noxref_d N_noxref_23_c_3084_n ) capacitor \
 c=0.00211996f //x=24.935 //y=0.875 //x2=24.86 //y2=0.875
cc_277 ( N_noxref_1_M15_noxref_d N_noxref_23_c_3086_n ) capacitor \
 c=0.00255985f //x=24.935 //y=0.875 //x2=24.86 //y2=1.22
cc_278 ( N_noxref_1_c_7_p N_noxref_23_c_3087_n ) capacitor c=0.00204716f \
 //x=24.05 //y=0 //x2=24.86 //y2=1.53
cc_279 ( N_noxref_1_c_7_p N_noxref_23_c_3088_n ) capacitor c=0.0118433f \
 //x=24.05 //y=0 //x2=24.86 //y2=1.915
cc_280 ( N_noxref_1_M15_noxref_d N_noxref_23_c_3089_n ) capacitor c=0.0131341f \
 //x=24.935 //y=0.875 //x2=25.235 //y2=0.72
cc_281 ( N_noxref_1_M15_noxref_d N_noxref_23_c_3090_n ) capacitor \
 c=0.00193146f //x=24.935 //y=0.875 //x2=25.235 //y2=1.375
cc_282 ( N_noxref_1_c_2_p N_noxref_23_c_3091_n ) capacitor c=0.00129018f \
 //x=28.12 //y=0 //x2=25.39 //y2=0.875
cc_283 ( N_noxref_1_M15_noxref_d N_noxref_23_c_3091_n ) capacitor \
 c=0.00257848f //x=24.935 //y=0.875 //x2=25.39 //y2=0.875
cc_284 ( N_noxref_1_M15_noxref_d N_noxref_23_c_3093_n ) capacitor \
 c=0.00255985f //x=24.935 //y=0.875 //x2=25.39 //y2=1.22
cc_285 ( N_noxref_1_c_71_p N_noxref_24_c_3144_n ) capacitor c=0.00540905f \
 //x=28.12 //y=0 //x2=25.525 //y2=1.59
cc_286 ( N_noxref_1_c_93_p N_noxref_24_c_3144_n ) capacitor c=0.00111539f \
 //x=25.04 //y=0 //x2=25.525 //y2=1.59
cc_287 ( N_noxref_1_c_2_p N_noxref_24_c_3144_n ) capacitor c=0.00180702f \
 //x=28.12 //y=0 //x2=25.525 //y2=1.59
cc_288 ( N_noxref_1_M15_noxref_d N_noxref_24_c_3144_n ) capacitor \
 c=0.00880514f //x=24.935 //y=0.875 //x2=25.525 //y2=1.59
cc_289 ( N_noxref_1_c_71_p N_noxref_24_c_3148_n ) capacitor c=0.00277579f \
 //x=28.12 //y=0 //x2=25.61 //y2=0.625
cc_290 ( N_noxref_1_c_2_p N_noxref_24_c_3148_n ) capacitor c=0.0142586f \
 //x=28.12 //y=0 //x2=25.61 //y2=0.625
cc_291 ( N_noxref_1_M15_noxref_d N_noxref_24_c_3148_n ) capacitor c=0.033954f \
 //x=24.935 //y=0.875 //x2=25.61 //y2=0.625
cc_292 ( N_noxref_1_c_71_p N_noxref_24_c_3151_n ) capacitor c=0.011436f \
 //x=28.12 //y=0 //x2=26.495 //y2=0.54
cc_293 ( N_noxref_1_c_2_p N_noxref_24_c_3151_n ) capacitor c=0.0385503f \
 //x=28.12 //y=0 //x2=26.495 //y2=0.54
cc_294 ( N_noxref_1_c_71_p N_noxref_24_M15_noxref_s ) capacitor c=0.00574679f \
 //x=28.12 //y=0 //x2=24.505 //y2=0.375
cc_295 ( N_noxref_1_c_93_p N_noxref_24_M15_noxref_s ) capacitor c=0.0142586f \
 //x=25.04 //y=0 //x2=24.505 //y2=0.375
cc_296 ( N_noxref_1_c_2_p N_noxref_24_M15_noxref_s ) capacitor c=0.0129524f \
 //x=28.12 //y=0 //x2=24.505 //y2=0.375
cc_297 ( N_noxref_1_c_7_p N_noxref_24_M15_noxref_s ) capacitor c=0.0696963f \
 //x=24.05 //y=0 //x2=24.505 //y2=0.375
cc_298 ( N_noxref_1_M15_noxref_d N_noxref_24_M15_noxref_s ) capacitor \
 c=0.033718f //x=24.935 //y=0.875 //x2=24.505 //y2=0.375
cc_299 ( N_noxref_1_c_2_p N_noxref_25_c_3194_n ) capacitor c=0.0465819f \
 //x=28.12 //y=0 //x2=28.035 //y2=1.665
cc_300 ( N_noxref_1_c_2_p N_noxref_25_M17_noxref_d ) capacitor c=0.00593061f \
 //x=28.12 //y=0 //x2=27.445 //y2=0.915
cc_301 ( N_noxref_1_c_71_p N_noxref_26_c_3271_n ) capacitor c=0.00394306f \
 //x=28.12 //y=0 //x2=27.065 //y2=0.995
cc_302 ( N_noxref_1_c_2_p N_noxref_26_c_3271_n ) capacitor c=0.00865404f \
 //x=28.12 //y=0 //x2=27.065 //y2=0.995
cc_303 ( N_noxref_1_c_71_p N_noxref_26_c_3273_n ) capacitor c=0.00296961f \
 //x=28.12 //y=0 //x2=27.15 //y2=0.625
cc_304 ( N_noxref_1_c_2_p N_noxref_26_c_3273_n ) capacitor c=0.0140218f \
 //x=28.12 //y=0 //x2=27.15 //y2=0.625
cc_305 ( N_noxref_1_M15_noxref_d N_noxref_26_c_3273_n ) capacitor \
 c=6.21394e-19 //x=24.935 //y=0.875 //x2=27.15 //y2=0.625
cc_306 ( N_noxref_1_c_71_p N_noxref_26_c_3276_n ) capacitor c=0.0167017f \
 //x=28.12 //y=0 //x2=28.035 //y2=0.54
cc_307 ( N_noxref_1_c_2_p N_noxref_26_c_3276_n ) capacitor c=0.0388692f \
 //x=28.12 //y=0 //x2=28.035 //y2=0.54
cc_308 ( N_noxref_1_c_71_p N_noxref_26_c_3278_n ) capacitor c=0.00705484f \
 //x=28.12 //y=0 //x2=28.12 //y2=0.625
cc_309 ( N_noxref_1_c_2_p N_noxref_26_c_3278_n ) capacitor c=0.0549101f \
 //x=28.12 //y=0 //x2=28.12 //y2=0.625
cc_310 ( N_noxref_1_M15_noxref_d N_noxref_26_M16_noxref_d ) capacitor \
 c=0.00162435f //x=24.935 //y=0.875 //x2=25.91 //y2=0.91
cc_311 ( N_noxref_1_c_2_p N_noxref_26_M17_noxref_s ) capacitor c=0.00183576f \
 //x=28.12 //y=0 //x2=27.015 //y2=0.375
cc_312 ( N_noxref_1_c_7_p N_noxref_26_M17_noxref_s ) capacitor c=8.16352e-19 \
 //x=24.05 //y=0 //x2=27.015 //y2=0.375
cc_313 ( N_noxref_2_c_320_p N_noxref_3_c_673_n ) capacitor c=0.0058961f \
 //x=28.12 //y=7.4 //x2=2.325 //y2=5.155
cc_314 ( N_noxref_2_c_321_p N_noxref_3_c_673_n ) capacitor c=4.18223e-19 \
 //x=1.885 //y=7.4 //x2=2.325 //y2=5.155
cc_315 ( N_noxref_2_c_322_p N_noxref_3_c_673_n ) capacitor c=4.18223e-19 \
 //x=2.765 //y=7.4 //x2=2.325 //y2=5.155
cc_316 ( N_noxref_2_M19_noxref_d N_noxref_3_c_673_n ) capacitor c=0.0119114f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_317 ( N_noxref_2_c_313_n N_noxref_3_c_677_n ) capacitor c=0.00880189f \
 //x=0.74 //y=7.4 //x2=1.615 //y2=5.155
cc_318 ( N_noxref_2_M18_noxref_s N_noxref_3_c_677_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_319 ( N_noxref_2_c_320_p N_noxref_3_c_679_n ) capacitor c=0.00539117f \
 //x=28.12 //y=7.4 //x2=3.205 //y2=5.155
cc_320 ( N_noxref_2_c_322_p N_noxref_3_c_679_n ) capacitor c=4.18223e-19 \
 //x=2.765 //y=7.4 //x2=3.205 //y2=5.155
cc_321 ( N_noxref_2_c_328_p N_noxref_3_c_679_n ) capacitor c=4.18223e-19 \
 //x=3.645 //y=7.4 //x2=3.205 //y2=5.155
cc_322 ( N_noxref_2_M21_noxref_d N_noxref_3_c_679_n ) capacitor c=0.0118689f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_323 ( N_noxref_2_c_320_p N_noxref_3_c_683_n ) capacitor c=0.00456797f \
 //x=28.12 //y=7.4 //x2=3.985 //y2=5.155
cc_324 ( N_noxref_2_c_328_p N_noxref_3_c_683_n ) capacitor c=6.98646e-19 \
 //x=3.645 //y=7.4 //x2=3.985 //y2=5.155
cc_325 ( N_noxref_2_c_332_p N_noxref_3_c_683_n ) capacitor c=0.00179956f \
 //x=4.64 //y=7.4 //x2=3.985 //y2=5.155
cc_326 ( N_noxref_2_M23_noxref_d N_noxref_3_c_683_n ) capacitor c=0.0117481f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_327 ( N_noxref_2_c_315_n N_noxref_3_c_649_n ) capacitor c=0.0457553f \
 //x=4.81 //y=7.4 //x2=4.07 //y2=2.59
cc_328 ( N_noxref_2_c_320_p N_noxref_3_c_650_n ) capacitor c=9.47191e-19 \
 //x=28.12 //y=7.4 //x2=5.92 //y2=2.08
cc_329 ( N_noxref_2_c_315_n N_noxref_3_c_650_n ) capacitor c=0.0164579f \
 //x=4.81 //y=7.4 //x2=5.92 //y2=2.08
cc_330 ( N_noxref_2_M24_noxref_s N_noxref_3_c_650_n ) capacitor c=0.0126291f \
 //x=5.765 //y=5.02 //x2=5.92 //y2=2.08
cc_331 ( N_noxref_2_c_320_p N_noxref_3_c_651_n ) capacitor c=9.10347e-19 \
 //x=28.12 //y=7.4 //x2=10.73 //y2=2.08
cc_332 ( N_noxref_2_c_316_n N_noxref_3_c_651_n ) capacitor c=0.0141571f \
 //x=9.62 //y=7.4 //x2=10.73 //y2=2.08
cc_333 ( N_noxref_2_M30_noxref_s N_noxref_3_c_651_n ) capacitor c=0.0125322f \
 //x=10.575 //y=5.02 //x2=10.73 //y2=2.08
cc_334 ( N_noxref_2_c_341_p N_noxref_3_M24_noxref_g ) capacitor c=0.00749687f \
 //x=6.695 //y=7.4 //x2=6.12 //y2=6.02
cc_335 ( N_noxref_2_M24_noxref_s N_noxref_3_M24_noxref_g ) capacitor \
 c=0.0477201f //x=5.765 //y=5.02 //x2=6.12 //y2=6.02
cc_336 ( N_noxref_2_c_341_p N_noxref_3_M25_noxref_g ) capacitor c=0.00675175f \
 //x=6.695 //y=7.4 //x2=6.56 //y2=6.02
cc_337 ( N_noxref_2_M25_noxref_d N_noxref_3_M25_noxref_g ) capacitor \
 c=0.015318f //x=6.635 //y=5.02 //x2=6.56 //y2=6.02
cc_338 ( N_noxref_2_c_345_p N_noxref_3_M30_noxref_g ) capacitor c=0.00749687f \
 //x=11.505 //y=7.4 //x2=10.93 //y2=6.02
cc_339 ( N_noxref_2_M30_noxref_s N_noxref_3_M30_noxref_g ) capacitor \
 c=0.0477201f //x=10.575 //y=5.02 //x2=10.93 //y2=6.02
cc_340 ( N_noxref_2_c_345_p N_noxref_3_M31_noxref_g ) capacitor c=0.00675175f \
 //x=11.505 //y=7.4 //x2=11.37 //y2=6.02
cc_341 ( N_noxref_2_M31_noxref_d N_noxref_3_M31_noxref_g ) capacitor \
 c=0.015318f //x=11.445 //y=5.02 //x2=11.37 //y2=6.02
cc_342 ( N_noxref_2_c_315_n N_noxref_3_c_702_n ) capacitor c=0.00757682f \
 //x=4.81 //y=7.4 //x2=6.195 //y2=4.79
cc_343 ( N_noxref_2_M24_noxref_s N_noxref_3_c_702_n ) capacitor c=0.00446175f \
 //x=5.765 //y=5.02 //x2=6.195 //y2=4.79
cc_344 ( N_noxref_2_c_316_n N_noxref_3_c_704_n ) capacitor c=0.00757682f \
 //x=9.62 //y=7.4 //x2=11.005 //y2=4.79
cc_345 ( N_noxref_2_M30_noxref_s N_noxref_3_c_704_n ) capacitor c=0.00444914f \
 //x=10.575 //y=5.02 //x2=11.005 //y2=4.79
cc_346 ( N_noxref_2_c_320_p N_noxref_3_M18_noxref_d ) capacitor c=0.00706456f \
 //x=28.12 //y=7.4 //x2=1.385 //y2=5.02
cc_347 ( N_noxref_2_c_321_p N_noxref_3_M18_noxref_d ) capacitor c=0.0138437f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_348 ( N_noxref_2_M19_noxref_d N_noxref_3_M18_noxref_d ) capacitor \
 c=0.0664752f //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_349 ( N_noxref_2_c_320_p N_noxref_3_M20_noxref_d ) capacitor c=0.00706456f \
 //x=28.12 //y=7.4 //x2=2.265 //y2=5.02
cc_350 ( N_noxref_2_c_322_p N_noxref_3_M20_noxref_d ) capacitor c=0.0138437f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_351 ( N_noxref_2_c_315_n N_noxref_3_M20_noxref_d ) capacitor c=4.9285e-19 \
 //x=4.81 //y=7.4 //x2=2.265 //y2=5.02
cc_352 ( N_noxref_2_M18_noxref_s N_noxref_3_M20_noxref_d ) capacitor \
 c=0.00130656f //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_353 ( N_noxref_2_M19_noxref_d N_noxref_3_M20_noxref_d ) capacitor \
 c=0.0664752f //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_354 ( N_noxref_2_M21_noxref_d N_noxref_3_M20_noxref_d ) capacitor \
 c=0.0664752f //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_355 ( N_noxref_2_c_320_p N_noxref_3_M22_noxref_d ) capacitor c=0.00574237f \
 //x=28.12 //y=7.4 //x2=3.145 //y2=5.02
cc_356 ( N_noxref_2_c_328_p N_noxref_3_M22_noxref_d ) capacitor c=0.0137718f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_357 ( N_noxref_2_c_315_n N_noxref_3_M22_noxref_d ) capacitor c=0.00939849f \
 //x=4.81 //y=7.4 //x2=3.145 //y2=5.02
cc_358 ( N_noxref_2_M21_noxref_d N_noxref_3_M22_noxref_d ) capacitor \
 c=0.0664752f //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_359 ( N_noxref_2_M23_noxref_d N_noxref_3_M22_noxref_d ) capacitor \
 c=0.0664752f //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_360 ( N_noxref_2_M24_noxref_s N_noxref_3_M22_noxref_d ) capacitor \
 c=3.57641e-19 //x=5.765 //y=5.02 //x2=3.145 //y2=5.02
cc_361 ( N_noxref_2_c_320_p N_noxref_4_c_897_n ) capacitor c=0.00444892f \
 //x=28.12 //y=7.4 //x2=11.945 //y2=5.155
cc_362 ( N_noxref_2_c_345_p N_noxref_4_c_897_n ) capacitor c=4.31931e-19 \
 //x=11.505 //y=7.4 //x2=11.945 //y2=5.155
cc_363 ( N_noxref_2_c_370_p N_noxref_4_c_897_n ) capacitor c=4.31931e-19 \
 //x=12.385 //y=7.4 //x2=11.945 //y2=5.155
cc_364 ( N_noxref_2_M31_noxref_d N_noxref_4_c_897_n ) capacitor c=0.0112985f \
 //x=11.445 //y=5.02 //x2=11.945 //y2=5.155
cc_365 ( N_noxref_2_c_316_n N_noxref_4_c_901_n ) capacitor c=0.00863585f \
 //x=9.62 //y=7.4 //x2=11.235 //y2=5.155
cc_366 ( N_noxref_2_M30_noxref_s N_noxref_4_c_901_n ) capacitor c=0.0831083f \
 //x=10.575 //y=5.02 //x2=11.235 //y2=5.155
cc_367 ( N_noxref_2_c_320_p N_noxref_4_c_903_n ) capacitor c=0.0044221f \
 //x=28.12 //y=7.4 //x2=12.825 //y2=5.155
cc_368 ( N_noxref_2_c_370_p N_noxref_4_c_903_n ) capacitor c=4.31931e-19 \
 //x=12.385 //y=7.4 //x2=12.825 //y2=5.155
cc_369 ( N_noxref_2_c_376_p N_noxref_4_c_903_n ) capacitor c=4.31931e-19 \
 //x=13.265 //y=7.4 //x2=12.825 //y2=5.155
cc_370 ( N_noxref_2_M33_noxref_d N_noxref_4_c_903_n ) capacitor c=0.0112985f \
 //x=12.325 //y=5.02 //x2=12.825 //y2=5.155
cc_371 ( N_noxref_2_c_320_p N_noxref_4_c_907_n ) capacitor c=0.00434174f \
 //x=28.12 //y=7.4 //x2=13.605 //y2=5.155
cc_372 ( N_noxref_2_c_376_p N_noxref_4_c_907_n ) capacitor c=7.46626e-19 \
 //x=13.265 //y=7.4 //x2=13.605 //y2=5.155
cc_373 ( N_noxref_2_c_380_p N_noxref_4_c_907_n ) capacitor c=0.00198565f \
 //x=14.26 //y=7.4 //x2=13.605 //y2=5.155
cc_374 ( N_noxref_2_M35_noxref_d N_noxref_4_c_907_n ) capacitor c=0.0112985f \
 //x=13.205 //y=5.02 //x2=13.605 //y2=5.155
cc_375 ( N_noxref_2_c_317_n N_noxref_4_c_884_n ) capacitor c=0.0434114f \
 //x=14.43 //y=7.4 //x2=13.69 //y2=2.59
cc_376 ( N_noxref_2_c_320_p N_noxref_4_c_885_n ) capacitor c=9.10347e-19 \
 //x=28.12 //y=7.4 //x2=15.54 //y2=2.08
cc_377 ( N_noxref_2_c_317_n N_noxref_4_c_885_n ) capacitor c=0.0140972f \
 //x=14.43 //y=7.4 //x2=15.54 //y2=2.08
cc_378 ( N_noxref_2_M36_noxref_s N_noxref_4_c_885_n ) capacitor c=0.0125322f \
 //x=15.385 //y=5.02 //x2=15.54 //y2=2.08
cc_379 ( N_noxref_2_c_386_p N_noxref_4_M36_noxref_g ) capacitor c=0.00749687f \
 //x=16.315 //y=7.4 //x2=15.74 //y2=6.02
cc_380 ( N_noxref_2_M36_noxref_s N_noxref_4_M36_noxref_g ) capacitor \
 c=0.0477201f //x=15.385 //y=5.02 //x2=15.74 //y2=6.02
cc_381 ( N_noxref_2_c_386_p N_noxref_4_M37_noxref_g ) capacitor c=0.00675175f \
 //x=16.315 //y=7.4 //x2=16.18 //y2=6.02
cc_382 ( N_noxref_2_M37_noxref_d N_noxref_4_M37_noxref_g ) capacitor \
 c=0.015318f //x=16.255 //y=5.02 //x2=16.18 //y2=6.02
cc_383 ( N_noxref_2_c_317_n N_noxref_4_c_919_n ) capacitor c=0.00757682f \
 //x=14.43 //y=7.4 //x2=15.815 //y2=4.79
cc_384 ( N_noxref_2_M36_noxref_s N_noxref_4_c_919_n ) capacitor c=0.00444914f \
 //x=15.385 //y=5.02 //x2=15.815 //y2=4.79
cc_385 ( N_noxref_2_c_320_p N_noxref_4_M30_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=11.005 //y2=5.02
cc_386 ( N_noxref_2_c_345_p N_noxref_4_M30_noxref_d ) capacitor c=0.014035f \
 //x=11.505 //y=7.4 //x2=11.005 //y2=5.02
cc_387 ( N_noxref_2_M31_noxref_d N_noxref_4_M30_noxref_d ) capacitor \
 c=0.0664752f //x=11.445 //y=5.02 //x2=11.005 //y2=5.02
cc_388 ( N_noxref_2_c_320_p N_noxref_4_M32_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=11.885 //y2=5.02
cc_389 ( N_noxref_2_c_370_p N_noxref_4_M32_noxref_d ) capacitor c=0.014035f \
 //x=12.385 //y=7.4 //x2=11.885 //y2=5.02
cc_390 ( N_noxref_2_c_317_n N_noxref_4_M32_noxref_d ) capacitor c=4.9285e-19 \
 //x=14.43 //y=7.4 //x2=11.885 //y2=5.02
cc_391 ( N_noxref_2_M30_noxref_s N_noxref_4_M32_noxref_d ) capacitor \
 c=0.00130656f //x=10.575 //y=5.02 //x2=11.885 //y2=5.02
cc_392 ( N_noxref_2_M31_noxref_d N_noxref_4_M32_noxref_d ) capacitor \
 c=0.0664752f //x=11.445 //y=5.02 //x2=11.885 //y2=5.02
cc_393 ( N_noxref_2_M33_noxref_d N_noxref_4_M32_noxref_d ) capacitor \
 c=0.0664752f //x=12.325 //y=5.02 //x2=11.885 //y2=5.02
cc_394 ( N_noxref_2_c_320_p N_noxref_4_M34_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=12.765 //y2=5.02
cc_395 ( N_noxref_2_c_376_p N_noxref_4_M34_noxref_d ) capacitor c=0.0137384f \
 //x=13.265 //y=7.4 //x2=12.765 //y2=5.02
cc_396 ( N_noxref_2_c_317_n N_noxref_4_M34_noxref_d ) capacitor c=0.00939849f \
 //x=14.43 //y=7.4 //x2=12.765 //y2=5.02
cc_397 ( N_noxref_2_M33_noxref_d N_noxref_4_M34_noxref_d ) capacitor \
 c=0.0664752f //x=12.325 //y=5.02 //x2=12.765 //y2=5.02
cc_398 ( N_noxref_2_M35_noxref_d N_noxref_4_M34_noxref_d ) capacitor \
 c=0.0664752f //x=13.205 //y=5.02 //x2=12.765 //y2=5.02
cc_399 ( N_noxref_2_M36_noxref_s N_noxref_4_M34_noxref_d ) capacitor \
 c=3.57641e-19 //x=15.385 //y=5.02 //x2=12.765 //y2=5.02
cc_400 ( N_noxref_2_c_320_p N_noxref_5_c_1045_n ) capacitor c=0.0725458f \
 //x=28.12 //y=7.4 //x2=16.535 //y2=4.44
cc_401 ( N_noxref_2_c_408_p N_noxref_5_c_1045_n ) capacitor c=0.00258496f \
 //x=9.45 //y=7.4 //x2=16.535 //y2=4.44
cc_402 ( N_noxref_2_c_409_p N_noxref_5_c_1045_n ) capacitor c=0.00328994f \
 //x=10.625 //y=7.4 //x2=16.535 //y2=4.44
cc_403 ( N_noxref_2_c_345_p N_noxref_5_c_1045_n ) capacitor c=0.00135925f \
 //x=11.505 //y=7.4 //x2=16.535 //y2=4.44
cc_404 ( N_noxref_2_c_380_p N_noxref_5_c_1045_n ) capacitor c=0.00258496f \
 //x=14.26 //y=7.4 //x2=16.535 //y2=4.44
cc_405 ( N_noxref_2_c_412_p N_noxref_5_c_1045_n ) capacitor c=0.00328994f \
 //x=15.435 //y=7.4 //x2=16.535 //y2=4.44
cc_406 ( N_noxref_2_c_386_p N_noxref_5_c_1045_n ) capacitor c=0.00135925f \
 //x=16.315 //y=7.4 //x2=16.535 //y2=4.44
cc_407 ( N_noxref_2_c_316_n N_noxref_5_c_1045_n ) capacitor c=0.0375613f \
 //x=9.62 //y=7.4 //x2=16.535 //y2=4.44
cc_408 ( N_noxref_2_c_317_n N_noxref_5_c_1045_n ) capacitor c=0.0375613f \
 //x=14.43 //y=7.4 //x2=16.535 //y2=4.44
cc_409 ( N_noxref_2_M30_noxref_s N_noxref_5_c_1045_n ) capacitor c=0.00179496f \
 //x=10.575 //y=5.02 //x2=16.535 //y2=4.44
cc_410 ( N_noxref_2_M36_noxref_s N_noxref_5_c_1045_n ) capacitor c=0.00179496f \
 //x=15.385 //y=5.02 //x2=16.535 //y2=4.44
cc_411 ( N_noxref_2_c_320_p N_noxref_5_c_1056_n ) capacitor c=0.00146064f \
 //x=28.12 //y=7.4 //x2=7.145 //y2=4.44
cc_412 ( N_noxref_2_c_320_p N_noxref_5_c_1043_n ) capacitor c=2.03287e-19 \
 //x=28.12 //y=7.4 //x2=7.03 //y2=2.08
cc_413 ( N_noxref_2_c_315_n N_noxref_5_c_1043_n ) capacitor c=8.7832e-19 \
 //x=4.81 //y=7.4 //x2=7.03 //y2=2.08
cc_414 ( N_noxref_2_c_320_p N_noxref_5_c_1044_n ) capacitor c=2.03287e-19 \
 //x=28.12 //y=7.4 //x2=16.65 //y2=2.08
cc_415 ( N_noxref_2_c_317_n N_noxref_5_c_1044_n ) capacitor c=6.46361e-19 \
 //x=14.43 //y=7.4 //x2=16.65 //y2=2.08
cc_416 ( N_noxref_2_c_423_p N_noxref_5_M26_noxref_g ) capacitor c=0.00676195f \
 //x=7.575 //y=7.4 //x2=7 //y2=6.02
cc_417 ( N_noxref_2_M25_noxref_d N_noxref_5_M26_noxref_g ) capacitor \
 c=0.015318f //x=6.635 //y=5.02 //x2=7 //y2=6.02
cc_418 ( N_noxref_2_c_423_p N_noxref_5_M27_noxref_g ) capacitor c=0.00675175f \
 //x=7.575 //y=7.4 //x2=7.44 //y2=6.02
cc_419 ( N_noxref_2_M27_noxref_d N_noxref_5_M27_noxref_g ) capacitor \
 c=0.015318f //x=7.515 //y=5.02 //x2=7.44 //y2=6.02
cc_420 ( N_noxref_2_c_427_p N_noxref_5_M38_noxref_g ) capacitor c=0.00676195f \
 //x=17.195 //y=7.4 //x2=16.62 //y2=6.02
cc_421 ( N_noxref_2_M37_noxref_d N_noxref_5_M38_noxref_g ) capacitor \
 c=0.015318f //x=16.255 //y=5.02 //x2=16.62 //y2=6.02
cc_422 ( N_noxref_2_c_427_p N_noxref_5_M39_noxref_g ) capacitor c=0.00675175f \
 //x=17.195 //y=7.4 //x2=17.06 //y2=6.02
cc_423 ( N_noxref_2_M39_noxref_d N_noxref_5_M39_noxref_g ) capacitor \
 c=0.015318f //x=17.135 //y=5.02 //x2=17.06 //y2=6.02
cc_424 ( N_noxref_2_c_320_p N_noxref_6_c_1247_n ) capacitor c=0.0217405f \
 //x=28.12 //y=7.4 //x2=8.765 //y2=3.33
cc_425 ( N_noxref_2_c_315_n N_noxref_6_c_1247_n ) capacitor c=0.0069465f \
 //x=4.81 //y=7.4 //x2=8.765 //y2=3.33
cc_426 ( N_noxref_2_M24_noxref_s N_noxref_6_c_1247_n ) capacitor c=7.16349e-19 \
 //x=5.765 //y=5.02 //x2=8.765 //y2=3.33
cc_427 ( N_noxref_2_c_320_p N_noxref_6_c_1266_n ) capacitor c=0.00148944f \
 //x=28.12 //y=7.4 //x2=3.445 //y2=3.33
cc_428 ( N_noxref_2_c_315_n N_noxref_6_c_1249_n ) capacitor c=8.81482e-19 \
 //x=4.81 //y=7.4 //x2=3.33 //y2=2.08
cc_429 ( N_noxref_2_c_320_p N_noxref_6_c_1268_n ) capacitor c=0.00456856f \
 //x=28.12 //y=7.4 //x2=7.135 //y2=5.155
cc_430 ( N_noxref_2_c_341_p N_noxref_6_c_1268_n ) capacitor c=4.18223e-19 \
 //x=6.695 //y=7.4 //x2=7.135 //y2=5.155
cc_431 ( N_noxref_2_c_423_p N_noxref_6_c_1268_n ) capacitor c=4.31906e-19 \
 //x=7.575 //y=7.4 //x2=7.135 //y2=5.155
cc_432 ( N_noxref_2_M25_noxref_d N_noxref_6_c_1268_n ) capacitor c=0.0117481f \
 //x=6.635 //y=5.02 //x2=7.135 //y2=5.155
cc_433 ( N_noxref_2_c_315_n N_noxref_6_c_1272_n ) capacitor c=0.00863585f \
 //x=4.81 //y=7.4 //x2=6.425 //y2=5.155
cc_434 ( N_noxref_2_M24_noxref_s N_noxref_6_c_1272_n ) capacitor c=0.0831083f \
 //x=5.765 //y=5.02 //x2=6.425 //y2=5.155
cc_435 ( N_noxref_2_c_320_p N_noxref_6_c_1274_n ) capacitor c=0.0044221f \
 //x=28.12 //y=7.4 //x2=8.015 //y2=5.155
cc_436 ( N_noxref_2_c_423_p N_noxref_6_c_1274_n ) capacitor c=4.31931e-19 \
 //x=7.575 //y=7.4 //x2=8.015 //y2=5.155
cc_437 ( N_noxref_2_c_444_p N_noxref_6_c_1274_n ) capacitor c=4.31931e-19 \
 //x=8.455 //y=7.4 //x2=8.015 //y2=5.155
cc_438 ( N_noxref_2_M27_noxref_d N_noxref_6_c_1274_n ) capacitor c=0.0112985f \
 //x=7.515 //y=5.02 //x2=8.015 //y2=5.155
cc_439 ( N_noxref_2_c_320_p N_noxref_6_c_1278_n ) capacitor c=0.00434174f \
 //x=28.12 //y=7.4 //x2=8.795 //y2=5.155
cc_440 ( N_noxref_2_c_444_p N_noxref_6_c_1278_n ) capacitor c=7.46626e-19 \
 //x=8.455 //y=7.4 //x2=8.795 //y2=5.155
cc_441 ( N_noxref_2_c_408_p N_noxref_6_c_1278_n ) capacitor c=0.00198565f \
 //x=9.45 //y=7.4 //x2=8.795 //y2=5.155
cc_442 ( N_noxref_2_M29_noxref_d N_noxref_6_c_1278_n ) capacitor c=0.0112985f \
 //x=8.395 //y=5.02 //x2=8.795 //y2=5.155
cc_443 ( N_noxref_2_c_316_n N_noxref_6_c_1282_n ) capacitor c=0.043403f \
 //x=9.62 //y=7.4 //x2=8.88 //y2=3.33
cc_444 ( N_noxref_2_c_320_p N_noxref_6_c_1251_n ) capacitor c=9.35768e-19 \
 //x=28.12 //y=7.4 //x2=20.35 //y2=2.08
cc_445 ( N_noxref_2_c_318_n N_noxref_6_c_1251_n ) capacitor c=0.0167484f \
 //x=19.24 //y=7.4 //x2=20.35 //y2=2.08
cc_446 ( N_noxref_2_M42_noxref_s N_noxref_6_c_1251_n ) capacitor c=0.0125045f \
 //x=20.195 //y=5.02 //x2=20.35 //y2=2.08
cc_447 ( N_noxref_2_c_328_p N_noxref_6_M22_noxref_g ) capacitor c=0.00675175f \
 //x=3.645 //y=7.4 //x2=3.07 //y2=6.02
cc_448 ( N_noxref_2_M21_noxref_d N_noxref_6_M22_noxref_g ) capacitor \
 c=0.015318f //x=2.705 //y=5.02 //x2=3.07 //y2=6.02
cc_449 ( N_noxref_2_c_328_p N_noxref_6_M23_noxref_g ) capacitor c=0.00675379f \
 //x=3.645 //y=7.4 //x2=3.51 //y2=6.02
cc_450 ( N_noxref_2_M23_noxref_d N_noxref_6_M23_noxref_g ) capacitor \
 c=0.0394719f //x=3.585 //y=5.02 //x2=3.51 //y2=6.02
cc_451 ( N_noxref_2_c_458_p N_noxref_6_M42_noxref_g ) capacitor c=0.00749687f \
 //x=21.125 //y=7.4 //x2=20.55 //y2=6.02
cc_452 ( N_noxref_2_M42_noxref_s N_noxref_6_M42_noxref_g ) capacitor \
 c=0.0477201f //x=20.195 //y=5.02 //x2=20.55 //y2=6.02
cc_453 ( N_noxref_2_c_458_p N_noxref_6_M43_noxref_g ) capacitor c=0.00675175f \
 //x=21.125 //y=7.4 //x2=20.99 //y2=6.02
cc_454 ( N_noxref_2_M43_noxref_d N_noxref_6_M43_noxref_g ) capacitor \
 c=0.015318f //x=21.065 //y=5.02 //x2=20.99 //y2=6.02
cc_455 ( N_noxref_2_c_318_n N_noxref_6_c_1294_n ) capacitor c=0.00757682f \
 //x=19.24 //y=7.4 //x2=20.625 //y2=4.79
cc_456 ( N_noxref_2_M42_noxref_s N_noxref_6_c_1294_n ) capacitor c=0.00446175f \
 //x=20.195 //y=5.02 //x2=20.625 //y2=4.79
cc_457 ( N_noxref_2_c_320_p N_noxref_6_M24_noxref_d ) capacitor c=0.00574869f \
 //x=28.12 //y=7.4 //x2=6.195 //y2=5.02
cc_458 ( N_noxref_2_c_341_p N_noxref_6_M24_noxref_d ) capacitor c=0.0138437f \
 //x=6.695 //y=7.4 //x2=6.195 //y2=5.02
cc_459 ( N_noxref_2_M25_noxref_d N_noxref_6_M24_noxref_d ) capacitor \
 c=0.0664752f //x=6.635 //y=5.02 //x2=6.195 //y2=5.02
cc_460 ( N_noxref_2_c_320_p N_noxref_6_M26_noxref_d ) capacitor c=0.00275186f \
 //x=28.12 //y=7.4 //x2=7.075 //y2=5.02
cc_461 ( N_noxref_2_c_423_p N_noxref_6_M26_noxref_d ) capacitor c=0.0140346f \
 //x=7.575 //y=7.4 //x2=7.075 //y2=5.02
cc_462 ( N_noxref_2_c_316_n N_noxref_6_M26_noxref_d ) capacitor c=4.9285e-19 \
 //x=9.62 //y=7.4 //x2=7.075 //y2=5.02
cc_463 ( N_noxref_2_M24_noxref_s N_noxref_6_M26_noxref_d ) capacitor \
 c=0.00130656f //x=5.765 //y=5.02 //x2=7.075 //y2=5.02
cc_464 ( N_noxref_2_M25_noxref_d N_noxref_6_M26_noxref_d ) capacitor \
 c=0.0664752f //x=6.635 //y=5.02 //x2=7.075 //y2=5.02
cc_465 ( N_noxref_2_M27_noxref_d N_noxref_6_M26_noxref_d ) capacitor \
 c=0.0664752f //x=7.515 //y=5.02 //x2=7.075 //y2=5.02
cc_466 ( N_noxref_2_c_320_p N_noxref_6_M28_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=7.955 //y2=5.02
cc_467 ( N_noxref_2_c_444_p N_noxref_6_M28_noxref_d ) capacitor c=0.0137384f \
 //x=8.455 //y=7.4 //x2=7.955 //y2=5.02
cc_468 ( N_noxref_2_c_316_n N_noxref_6_M28_noxref_d ) capacitor c=0.00939849f \
 //x=9.62 //y=7.4 //x2=7.955 //y2=5.02
cc_469 ( N_noxref_2_M27_noxref_d N_noxref_6_M28_noxref_d ) capacitor \
 c=0.0664752f //x=7.515 //y=5.02 //x2=7.955 //y2=5.02
cc_470 ( N_noxref_2_M29_noxref_d N_noxref_6_M28_noxref_d ) capacitor \
 c=0.0664752f //x=8.395 //y=5.02 //x2=7.955 //y2=5.02
cc_471 ( N_noxref_2_M30_noxref_s N_noxref_6_M28_noxref_d ) capacitor \
 c=3.57641e-19 //x=10.575 //y=5.02 //x2=7.955 //y2=5.02
cc_472 ( N_noxref_2_c_320_p N_noxref_7_c_1528_n ) capacitor c=2.41299e-19 \
 //x=28.12 //y=7.4 //x2=2.22 //y2=2.08
cc_473 ( N_noxref_2_c_313_n N_noxref_7_c_1528_n ) capacitor c=7.34553e-19 \
 //x=0.74 //y=7.4 //x2=2.22 //y2=2.08
cc_474 ( N_noxref_2_c_318_n N_noxref_7_c_1529_n ) capacitor c=0.00121089f \
 //x=19.24 //y=7.4 //x2=17.76 //y2=2.08
cc_475 ( N_noxref_2_c_320_p N_noxref_7_c_1530_n ) capacitor c=2.07998e-19 \
 //x=28.12 //y=7.4 //x2=21.46 //y2=2.08
cc_476 ( N_noxref_2_c_318_n N_noxref_7_c_1530_n ) capacitor c=7.34553e-19 \
 //x=19.24 //y=7.4 //x2=21.46 //y2=2.08
cc_477 ( N_noxref_2_c_322_p N_noxref_7_M20_noxref_g ) capacitor c=0.00676195f \
 //x=2.765 //y=7.4 //x2=2.19 //y2=6.02
cc_478 ( N_noxref_2_M19_noxref_d N_noxref_7_M20_noxref_g ) capacitor \
 c=0.015318f //x=1.825 //y=5.02 //x2=2.19 //y2=6.02
cc_479 ( N_noxref_2_c_322_p N_noxref_7_M21_noxref_g ) capacitor c=0.00675175f \
 //x=2.765 //y=7.4 //x2=2.63 //y2=6.02
cc_480 ( N_noxref_2_M21_noxref_d N_noxref_7_M21_noxref_g ) capacitor \
 c=0.015318f //x=2.705 //y=5.02 //x2=2.63 //y2=6.02
cc_481 ( N_noxref_2_c_488_p N_noxref_7_M40_noxref_g ) capacitor c=0.00675175f \
 //x=18.075 //y=7.4 //x2=17.5 //y2=6.02
cc_482 ( N_noxref_2_M39_noxref_d N_noxref_7_M40_noxref_g ) capacitor \
 c=0.015318f //x=17.135 //y=5.02 //x2=17.5 //y2=6.02
cc_483 ( N_noxref_2_c_488_p N_noxref_7_M41_noxref_g ) capacitor c=0.00675379f \
 //x=18.075 //y=7.4 //x2=17.94 //y2=6.02
cc_484 ( N_noxref_2_M41_noxref_d N_noxref_7_M41_noxref_g ) capacitor \
 c=0.0394719f //x=18.015 //y=5.02 //x2=17.94 //y2=6.02
cc_485 ( N_noxref_2_c_492_p N_noxref_7_M44_noxref_g ) capacitor c=0.00676195f \
 //x=22.005 //y=7.4 //x2=21.43 //y2=6.02
cc_486 ( N_noxref_2_M43_noxref_d N_noxref_7_M44_noxref_g ) capacitor \
 c=0.015318f //x=21.065 //y=5.02 //x2=21.43 //y2=6.02
cc_487 ( N_noxref_2_c_492_p N_noxref_7_M45_noxref_g ) capacitor c=0.00675175f \
 //x=22.005 //y=7.4 //x2=21.87 //y2=6.02
cc_488 ( N_noxref_2_M45_noxref_d N_noxref_7_M45_noxref_g ) capacitor \
 c=0.015318f //x=21.945 //y=5.02 //x2=21.87 //y2=6.02
cc_489 ( N_noxref_2_c_320_p N_noxref_8_c_1833_n ) capacitor c=2.03486e-19 \
 //x=28.12 //y=7.4 //x2=11.84 //y2=2.08
cc_490 ( N_noxref_2_c_316_n N_noxref_8_c_1833_n ) capacitor c=6.19557e-19 \
 //x=9.62 //y=7.4 //x2=11.84 //y2=2.08
cc_491 ( N_noxref_2_c_320_p N_noxref_8_c_1834_n ) capacitor c=2.07998e-19 \
 //x=28.12 //y=7.4 //x2=26.27 //y2=2.08
cc_492 ( N_noxref_2_c_319_n N_noxref_8_c_1834_n ) capacitor c=7.34553e-19 \
 //x=24.05 //y=7.4 //x2=26.27 //y2=2.08
cc_493 ( N_noxref_2_c_370_p N_noxref_8_M32_noxref_g ) capacitor c=0.00676195f \
 //x=12.385 //y=7.4 //x2=11.81 //y2=6.02
cc_494 ( N_noxref_2_M31_noxref_d N_noxref_8_M32_noxref_g ) capacitor \
 c=0.015318f //x=11.445 //y=5.02 //x2=11.81 //y2=6.02
cc_495 ( N_noxref_2_c_370_p N_noxref_8_M33_noxref_g ) capacitor c=0.00675175f \
 //x=12.385 //y=7.4 //x2=12.25 //y2=6.02
cc_496 ( N_noxref_2_M33_noxref_d N_noxref_8_M33_noxref_g ) capacitor \
 c=0.015318f //x=12.325 //y=5.02 //x2=12.25 //y2=6.02
cc_497 ( N_noxref_2_c_504_p N_noxref_8_M50_noxref_g ) capacitor c=0.00676195f \
 //x=26.815 //y=7.4 //x2=26.24 //y2=6.02
cc_498 ( N_noxref_2_M49_noxref_d N_noxref_8_M50_noxref_g ) capacitor \
 c=0.015318f //x=25.875 //y=5.02 //x2=26.24 //y2=6.02
cc_499 ( N_noxref_2_c_504_p N_noxref_8_M51_noxref_g ) capacitor c=0.00675175f \
 //x=26.815 //y=7.4 //x2=26.68 //y2=6.02
cc_500 ( N_noxref_2_M51_noxref_d N_noxref_8_M51_noxref_g ) capacitor \
 c=0.015318f //x=26.755 //y=5.02 //x2=26.68 //y2=6.02
cc_501 ( N_noxref_2_c_316_n N_noxref_9_c_2034_n ) capacitor c=0.00686843f \
 //x=9.62 //y=7.4 //x2=12.835 //y2=3.7
cc_502 ( N_noxref_2_c_320_p N_noxref_9_c_2035_n ) capacitor c=0.0159925f \
 //x=28.12 //y=7.4 //x2=18.385 //y2=3.7
cc_503 ( N_noxref_2_c_317_n N_noxref_9_c_2035_n ) capacitor c=0.00686843f \
 //x=14.43 //y=7.4 //x2=18.385 //y2=3.7
cc_504 ( N_noxref_2_c_320_p N_noxref_9_c_2028_n ) capacitor c=0.0562032f \
 //x=28.12 //y=7.4 //x2=27.265 //y2=3.7
cc_505 ( N_noxref_2_c_318_n N_noxref_9_c_2028_n ) capacitor c=0.0109524f \
 //x=19.24 //y=7.4 //x2=27.265 //y2=3.7
cc_506 ( N_noxref_2_c_319_n N_noxref_9_c_2028_n ) capacitor c=0.0109524f \
 //x=24.05 //y=7.4 //x2=27.265 //y2=3.7
cc_507 ( N_noxref_2_M42_noxref_s N_noxref_9_c_2028_n ) capacitor c=9.16752e-19 \
 //x=20.195 //y=5.02 //x2=27.265 //y2=3.7
cc_508 ( N_noxref_2_M48_noxref_s N_noxref_9_c_2028_n ) capacitor c=9.16752e-19 \
 //x=25.005 //y=5.02 //x2=27.265 //y2=3.7
cc_509 ( N_noxref_2_c_320_p N_noxref_9_c_2042_n ) capacitor c=0.00155789f \
 //x=28.12 //y=7.4 //x2=18.615 //y2=3.7
cc_510 ( N_noxref_2_c_316_n N_noxref_9_c_2029_n ) capacitor c=7.23426e-19 \
 //x=9.62 //y=7.4 //x2=8.14 //y2=2.08
cc_511 ( N_noxref_2_c_317_n N_noxref_9_c_2030_n ) capacitor c=6.37426e-19 \
 //x=14.43 //y=7.4 //x2=12.95 //y2=2.08
cc_512 ( N_noxref_2_c_320_p N_noxref_9_c_2045_n ) capacitor c=0.00444751f \
 //x=28.12 //y=7.4 //x2=16.755 //y2=5.155
cc_513 ( N_noxref_2_c_386_p N_noxref_9_c_2045_n ) capacitor c=4.31931e-19 \
 //x=16.315 //y=7.4 //x2=16.755 //y2=5.155
cc_514 ( N_noxref_2_c_427_p N_noxref_9_c_2045_n ) capacitor c=4.31906e-19 \
 //x=17.195 //y=7.4 //x2=16.755 //y2=5.155
cc_515 ( N_noxref_2_M37_noxref_d N_noxref_9_c_2045_n ) capacitor c=0.0112985f \
 //x=16.255 //y=5.02 //x2=16.755 //y2=5.155
cc_516 ( N_noxref_2_c_317_n N_noxref_9_c_2049_n ) capacitor c=0.00863585f \
 //x=14.43 //y=7.4 //x2=16.045 //y2=5.155
cc_517 ( N_noxref_2_M36_noxref_s N_noxref_9_c_2049_n ) capacitor c=0.0831083f \
 //x=15.385 //y=5.02 //x2=16.045 //y2=5.155
cc_518 ( N_noxref_2_c_320_p N_noxref_9_c_2051_n ) capacitor c=0.00454915f \
 //x=28.12 //y=7.4 //x2=17.635 //y2=5.155
cc_519 ( N_noxref_2_c_427_p N_noxref_9_c_2051_n ) capacitor c=4.18223e-19 \
 //x=17.195 //y=7.4 //x2=17.635 //y2=5.155
cc_520 ( N_noxref_2_c_488_p N_noxref_9_c_2051_n ) capacitor c=4.18223e-19 \
 //x=18.075 //y=7.4 //x2=17.635 //y2=5.155
cc_521 ( N_noxref_2_M39_noxref_d N_noxref_9_c_2051_n ) capacitor c=0.0116565f \
 //x=17.135 //y=5.02 //x2=17.635 //y2=5.155
cc_522 ( N_noxref_2_c_320_p N_noxref_9_c_2055_n ) capacitor c=0.00449936f \
 //x=28.12 //y=7.4 //x2=18.415 //y2=5.155
cc_523 ( N_noxref_2_c_488_p N_noxref_9_c_2055_n ) capacitor c=6.98646e-19 \
 //x=18.075 //y=7.4 //x2=18.415 //y2=5.155
cc_524 ( N_noxref_2_c_531_p N_noxref_9_c_2055_n ) capacitor c=0.00179956f \
 //x=19.07 //y=7.4 //x2=18.415 //y2=5.155
cc_525 ( N_noxref_2_M41_noxref_d N_noxref_9_c_2055_n ) capacitor c=0.0116565f \
 //x=18.015 //y=5.02 //x2=18.415 //y2=5.155
cc_526 ( N_noxref_2_c_318_n N_noxref_9_c_2059_n ) capacitor c=0.0457225f \
 //x=19.24 //y=7.4 //x2=18.5 //y2=3.7
cc_527 ( N_noxref_2_c_314_n N_noxref_9_c_2032_n ) capacitor c=8.81482e-19 \
 //x=28.12 //y=7.4 //x2=27.38 //y2=2.08
cc_528 ( N_noxref_2_c_444_p N_noxref_9_M28_noxref_g ) capacitor c=0.00675175f \
 //x=8.455 //y=7.4 //x2=7.88 //y2=6.02
cc_529 ( N_noxref_2_M27_noxref_d N_noxref_9_M28_noxref_g ) capacitor \
 c=0.015318f //x=7.515 //y=5.02 //x2=7.88 //y2=6.02
cc_530 ( N_noxref_2_c_444_p N_noxref_9_M29_noxref_g ) capacitor c=0.00675379f \
 //x=8.455 //y=7.4 //x2=8.32 //y2=6.02
cc_531 ( N_noxref_2_M29_noxref_d N_noxref_9_M29_noxref_g ) capacitor \
 c=0.0394719f //x=8.395 //y=5.02 //x2=8.32 //y2=6.02
cc_532 ( N_noxref_2_c_376_p N_noxref_9_M34_noxref_g ) capacitor c=0.00675175f \
 //x=13.265 //y=7.4 //x2=12.69 //y2=6.02
cc_533 ( N_noxref_2_M33_noxref_d N_noxref_9_M34_noxref_g ) capacitor \
 c=0.015318f //x=12.325 //y=5.02 //x2=12.69 //y2=6.02
cc_534 ( N_noxref_2_c_376_p N_noxref_9_M35_noxref_g ) capacitor c=0.00675379f \
 //x=13.265 //y=7.4 //x2=13.13 //y2=6.02
cc_535 ( N_noxref_2_M35_noxref_d N_noxref_9_M35_noxref_g ) capacitor \
 c=0.0394719f //x=13.205 //y=5.02 //x2=13.13 //y2=6.02
cc_536 ( N_noxref_2_c_543_p N_noxref_9_M52_noxref_g ) capacitor c=0.00675175f \
 //x=27.695 //y=7.4 //x2=27.12 //y2=6.02
cc_537 ( N_noxref_2_M51_noxref_d N_noxref_9_M52_noxref_g ) capacitor \
 c=0.015318f //x=26.755 //y=5.02 //x2=27.12 //y2=6.02
cc_538 ( N_noxref_2_c_543_p N_noxref_9_M53_noxref_g ) capacitor c=0.00675379f \
 //x=27.695 //y=7.4 //x2=27.56 //y2=6.02
cc_539 ( N_noxref_2_M53_noxref_d N_noxref_9_M53_noxref_g ) capacitor \
 c=0.0394719f //x=27.635 //y=5.02 //x2=27.56 //y2=6.02
cc_540 ( N_noxref_2_c_320_p N_noxref_9_M36_noxref_d ) capacitor c=0.00275235f \
 //x=28.12 //y=7.4 //x2=15.815 //y2=5.02
cc_541 ( N_noxref_2_c_386_p N_noxref_9_M36_noxref_d ) capacitor c=0.014035f \
 //x=16.315 //y=7.4 //x2=15.815 //y2=5.02
cc_542 ( N_noxref_2_M37_noxref_d N_noxref_9_M36_noxref_d ) capacitor \
 c=0.0664752f //x=16.255 //y=5.02 //x2=15.815 //y2=5.02
cc_543 ( N_noxref_2_c_320_p N_noxref_9_M38_noxref_d ) capacitor c=0.00289706f \
 //x=28.12 //y=7.4 //x2=16.695 //y2=5.02
cc_544 ( N_noxref_2_c_427_p N_noxref_9_M38_noxref_d ) capacitor c=0.0138883f \
 //x=17.195 //y=7.4 //x2=16.695 //y2=5.02
cc_545 ( N_noxref_2_c_318_n N_noxref_9_M38_noxref_d ) capacitor c=4.9285e-19 \
 //x=19.24 //y=7.4 //x2=16.695 //y2=5.02
cc_546 ( N_noxref_2_M36_noxref_s N_noxref_9_M38_noxref_d ) capacitor \
 c=0.00130656f //x=15.385 //y=5.02 //x2=16.695 //y2=5.02
cc_547 ( N_noxref_2_M37_noxref_d N_noxref_9_M38_noxref_d ) capacitor \
 c=0.0664752f //x=16.255 //y=5.02 //x2=16.695 //y2=5.02
cc_548 ( N_noxref_2_M39_noxref_d N_noxref_9_M38_noxref_d ) capacitor \
 c=0.0664752f //x=17.135 //y=5.02 //x2=16.695 //y2=5.02
cc_549 ( N_noxref_2_c_320_p N_noxref_9_M40_noxref_d ) capacitor c=0.00294223f \
 //x=28.12 //y=7.4 //x2=17.575 //y2=5.02
cc_550 ( N_noxref_2_c_488_p N_noxref_9_M40_noxref_d ) capacitor c=0.0137718f \
 //x=18.075 //y=7.4 //x2=17.575 //y2=5.02
cc_551 ( N_noxref_2_c_318_n N_noxref_9_M40_noxref_d ) capacitor c=0.00939849f \
 //x=19.24 //y=7.4 //x2=17.575 //y2=5.02
cc_552 ( N_noxref_2_M39_noxref_d N_noxref_9_M40_noxref_d ) capacitor \
 c=0.0664752f //x=17.135 //y=5.02 //x2=17.575 //y2=5.02
cc_553 ( N_noxref_2_M41_noxref_d N_noxref_9_M40_noxref_d ) capacitor \
 c=0.0664752f //x=18.015 //y=5.02 //x2=17.575 //y2=5.02
cc_554 ( N_noxref_2_M42_noxref_s N_noxref_9_M40_noxref_d ) capacitor \
 c=3.57641e-19 //x=20.195 //y=5.02 //x2=17.575 //y2=5.02
cc_555 ( N_noxref_2_c_320_p N_noxref_10_c_2364_n ) capacitor c=0.00112336f \
 //x=28.12 //y=7.4 //x2=1.11 //y2=2.08
cc_556 ( N_noxref_2_c_313_n N_noxref_10_c_2364_n ) capacitor c=0.0168497f \
 //x=0.74 //y=7.4 //x2=1.11 //y2=2.08
cc_557 ( N_noxref_2_M18_noxref_s N_noxref_10_c_2364_n ) capacitor c=0.0130213f \
 //x=0.955 //y=5.02 //x2=1.11 //y2=2.08
cc_558 ( N_noxref_2_c_321_p N_noxref_10_M18_noxref_g ) capacitor c=0.00749687f \
 //x=1.885 //y=7.4 //x2=1.31 //y2=6.02
cc_559 ( N_noxref_2_M18_noxref_s N_noxref_10_M18_noxref_g ) capacitor \
 c=0.0477201f //x=0.955 //y=5.02 //x2=1.31 //y2=6.02
cc_560 ( N_noxref_2_c_321_p N_noxref_10_M19_noxref_g ) capacitor c=0.00675175f \
 //x=1.885 //y=7.4 //x2=1.75 //y2=6.02
cc_561 ( N_noxref_2_M19_noxref_d N_noxref_10_M19_noxref_g ) capacitor \
 c=0.015318f //x=1.825 //y=5.02 //x2=1.75 //y2=6.02
cc_562 ( N_noxref_2_c_313_n N_noxref_10_c_2382_n ) capacitor c=0.0076931f \
 //x=0.74 //y=7.4 //x2=1.385 //y2=4.79
cc_563 ( N_noxref_2_M18_noxref_s N_noxref_10_c_2382_n ) capacitor \
 c=0.00442959f //x=0.955 //y=5.02 //x2=1.385 //y2=4.79
cc_564 ( N_noxref_2_c_319_n N_noxref_20_c_2886_n ) capacitor c=8.81482e-19 \
 //x=24.05 //y=7.4 //x2=22.57 //y2=2.08
cc_565 ( N_noxref_2_c_572_p N_noxref_20_M46_noxref_g ) capacitor c=0.00675175f \
 //x=22.885 //y=7.4 //x2=22.31 //y2=6.02
cc_566 ( N_noxref_2_M45_noxref_d N_noxref_20_M46_noxref_g ) capacitor \
 c=0.015318f //x=21.945 //y=5.02 //x2=22.31 //y2=6.02
cc_567 ( N_noxref_2_c_572_p N_noxref_20_M47_noxref_g ) capacitor c=0.00675379f \
 //x=22.885 //y=7.4 //x2=22.75 //y2=6.02
cc_568 ( N_noxref_2_M47_noxref_d N_noxref_20_M47_noxref_g ) capacitor \
 c=0.0394719f //x=22.825 //y=5.02 //x2=22.75 //y2=6.02
cc_569 ( N_noxref_2_c_320_p N_noxref_21_c_2947_n ) capacitor c=0.00457327f \
 //x=28.12 //y=7.4 //x2=21.565 //y2=5.155
cc_570 ( N_noxref_2_c_458_p N_noxref_21_c_2947_n ) capacitor c=4.18223e-19 \
 //x=21.125 //y=7.4 //x2=21.565 //y2=5.155
cc_571 ( N_noxref_2_c_492_p N_noxref_21_c_2947_n ) capacitor c=4.18223e-19 \
 //x=22.005 //y=7.4 //x2=21.565 //y2=5.155
cc_572 ( N_noxref_2_M43_noxref_d N_noxref_21_c_2947_n ) capacitor c=0.0116565f \
 //x=21.065 //y=5.02 //x2=21.565 //y2=5.155
cc_573 ( N_noxref_2_c_318_n N_noxref_21_c_2951_n ) capacitor c=0.00863585f \
 //x=19.24 //y=7.4 //x2=20.855 //y2=5.155
cc_574 ( N_noxref_2_M42_noxref_s N_noxref_21_c_2951_n ) capacitor c=0.0831083f \
 //x=20.195 //y=5.02 //x2=20.855 //y2=5.155
cc_575 ( N_noxref_2_c_320_p N_noxref_21_c_2953_n ) capacitor c=0.00454915f \
 //x=28.12 //y=7.4 //x2=22.445 //y2=5.155
cc_576 ( N_noxref_2_c_492_p N_noxref_21_c_2953_n ) capacitor c=4.18223e-19 \
 //x=22.005 //y=7.4 //x2=22.445 //y2=5.155
cc_577 ( N_noxref_2_c_572_p N_noxref_21_c_2953_n ) capacitor c=4.18223e-19 \
 //x=22.885 //y=7.4 //x2=22.445 //y2=5.155
cc_578 ( N_noxref_2_M45_noxref_d N_noxref_21_c_2953_n ) capacitor c=0.0116565f \
 //x=21.945 //y=5.02 //x2=22.445 //y2=5.155
cc_579 ( N_noxref_2_c_320_p N_noxref_21_c_2957_n ) capacitor c=0.00450078f \
 //x=28.12 //y=7.4 //x2=23.225 //y2=5.155
cc_580 ( N_noxref_2_c_572_p N_noxref_21_c_2957_n ) capacitor c=6.98646e-19 \
 //x=22.885 //y=7.4 //x2=23.225 //y2=5.155
cc_581 ( N_noxref_2_c_588_p N_noxref_21_c_2957_n ) capacitor c=0.00179956f \
 //x=23.88 //y=7.4 //x2=23.225 //y2=5.155
cc_582 ( N_noxref_2_M47_noxref_d N_noxref_21_c_2957_n ) capacitor c=0.0116565f \
 //x=22.825 //y=5.02 //x2=23.225 //y2=5.155
cc_583 ( N_noxref_2_c_319_n N_noxref_21_c_2961_n ) capacitor c=0.0461179f \
 //x=24.05 //y=7.4 //x2=23.31 //y2=5.07
cc_584 ( N_noxref_2_c_320_p N_noxref_21_M42_noxref_d ) capacitor c=0.00294223f \
 //x=28.12 //y=7.4 //x2=20.625 //y2=5.02
cc_585 ( N_noxref_2_c_458_p N_noxref_21_M42_noxref_d ) capacitor c=0.0138437f \
 //x=21.125 //y=7.4 //x2=20.625 //y2=5.02
cc_586 ( N_noxref_2_M43_noxref_d N_noxref_21_M42_noxref_d ) capacitor \
 c=0.0664752f //x=21.065 //y=5.02 //x2=20.625 //y2=5.02
cc_587 ( N_noxref_2_c_320_p N_noxref_21_M44_noxref_d ) capacitor c=0.00294223f \
 //x=28.12 //y=7.4 //x2=21.505 //y2=5.02
cc_588 ( N_noxref_2_c_492_p N_noxref_21_M44_noxref_d ) capacitor c=0.0138437f \
 //x=22.005 //y=7.4 //x2=21.505 //y2=5.02
cc_589 ( N_noxref_2_c_319_n N_noxref_21_M44_noxref_d ) capacitor c=4.9285e-19 \
 //x=24.05 //y=7.4 //x2=21.505 //y2=5.02
cc_590 ( N_noxref_2_M42_noxref_s N_noxref_21_M44_noxref_d ) capacitor \
 c=0.00130656f //x=20.195 //y=5.02 //x2=21.505 //y2=5.02
cc_591 ( N_noxref_2_M43_noxref_d N_noxref_21_M44_noxref_d ) capacitor \
 c=0.0664752f //x=21.065 //y=5.02 //x2=21.505 //y2=5.02
cc_592 ( N_noxref_2_M45_noxref_d N_noxref_21_M44_noxref_d ) capacitor \
 c=0.0664752f //x=21.945 //y=5.02 //x2=21.505 //y2=5.02
cc_593 ( N_noxref_2_c_320_p N_noxref_21_M46_noxref_d ) capacitor c=0.00294223f \
 //x=28.12 //y=7.4 //x2=22.385 //y2=5.02
cc_594 ( N_noxref_2_c_572_p N_noxref_21_M46_noxref_d ) capacitor c=0.0137718f \
 //x=22.885 //y=7.4 //x2=22.385 //y2=5.02
cc_595 ( N_noxref_2_c_319_n N_noxref_21_M46_noxref_d ) capacitor c=0.00939849f \
 //x=24.05 //y=7.4 //x2=22.385 //y2=5.02
cc_596 ( N_noxref_2_M45_noxref_d N_noxref_21_M46_noxref_d ) capacitor \
 c=0.0664752f //x=21.945 //y=5.02 //x2=22.385 //y2=5.02
cc_597 ( N_noxref_2_M47_noxref_d N_noxref_21_M46_noxref_d ) capacitor \
 c=0.0664752f //x=22.825 //y=5.02 //x2=22.385 //y2=5.02
cc_598 ( N_noxref_2_M48_noxref_s N_noxref_21_M46_noxref_d ) capacitor \
 c=3.57641e-19 //x=25.005 //y=5.02 //x2=22.385 //y2=5.02
cc_599 ( N_noxref_2_c_320_p N_noxref_23_c_3083_n ) capacitor c=9.35768e-19 \
 //x=28.12 //y=7.4 //x2=25.16 //y2=2.08
cc_600 ( N_noxref_2_c_319_n N_noxref_23_c_3083_n ) capacitor c=0.0167484f \
 //x=24.05 //y=7.4 //x2=25.16 //y2=2.08
cc_601 ( N_noxref_2_M48_noxref_s N_noxref_23_c_3083_n ) capacitor c=0.013204f \
 //x=25.005 //y=5.02 //x2=25.16 //y2=2.08
cc_602 ( N_noxref_2_c_609_p N_noxref_23_M48_noxref_g ) capacitor c=0.00749687f \
 //x=25.935 //y=7.4 //x2=25.36 //y2=6.02
cc_603 ( N_noxref_2_M48_noxref_s N_noxref_23_M48_noxref_g ) capacitor \
 c=0.0477201f //x=25.005 //y=5.02 //x2=25.36 //y2=6.02
cc_604 ( N_noxref_2_c_609_p N_noxref_23_M49_noxref_g ) capacitor c=0.00675175f \
 //x=25.935 //y=7.4 //x2=25.8 //y2=6.02
cc_605 ( N_noxref_2_M49_noxref_d N_noxref_23_M49_noxref_g ) capacitor \
 c=0.015318f //x=25.875 //y=5.02 //x2=25.8 //y2=6.02
cc_606 ( N_noxref_2_c_319_n N_noxref_23_c_3101_n ) capacitor c=0.0076931f \
 //x=24.05 //y=7.4 //x2=25.435 //y2=4.79
cc_607 ( N_noxref_2_M48_noxref_s N_noxref_23_c_3101_n ) capacitor \
 c=0.00446175f //x=25.005 //y=5.02 //x2=25.435 //y2=4.79
cc_608 ( N_noxref_2_c_320_p N_noxref_25_c_3196_n ) capacitor c=0.00457327f \
 //x=28.12 //y=7.4 //x2=26.375 //y2=5.155
cc_609 ( N_noxref_2_c_609_p N_noxref_25_c_3196_n ) capacitor c=4.18223e-19 \
 //x=25.935 //y=7.4 //x2=26.375 //y2=5.155
cc_610 ( N_noxref_2_c_504_p N_noxref_25_c_3196_n ) capacitor c=4.18223e-19 \
 //x=26.815 //y=7.4 //x2=26.375 //y2=5.155
cc_611 ( N_noxref_2_M49_noxref_d N_noxref_25_c_3196_n ) capacitor c=0.0116565f \
 //x=25.875 //y=5.02 //x2=26.375 //y2=5.155
cc_612 ( N_noxref_2_c_319_n N_noxref_25_c_3200_n ) capacitor c=0.00863585f \
 //x=24.05 //y=7.4 //x2=25.665 //y2=5.155
cc_613 ( N_noxref_2_M48_noxref_s N_noxref_25_c_3200_n ) capacitor c=0.0831083f \
 //x=25.005 //y=5.02 //x2=25.665 //y2=5.155
cc_614 ( N_noxref_2_c_320_p N_noxref_25_c_3202_n ) capacitor c=0.00454915f \
 //x=28.12 //y=7.4 //x2=27.255 //y2=5.155
cc_615 ( N_noxref_2_c_504_p N_noxref_25_c_3202_n ) capacitor c=4.18223e-19 \
 //x=26.815 //y=7.4 //x2=27.255 //y2=5.155
cc_616 ( N_noxref_2_c_543_p N_noxref_25_c_3202_n ) capacitor c=4.18223e-19 \
 //x=27.695 //y=7.4 //x2=27.255 //y2=5.155
cc_617 ( N_noxref_2_M51_noxref_d N_noxref_25_c_3202_n ) capacitor c=0.0116565f \
 //x=26.755 //y=5.02 //x2=27.255 //y2=5.155
cc_618 ( N_noxref_2_c_320_p N_noxref_25_c_3206_n ) capacitor c=0.00637429f \
 //x=28.12 //y=7.4 //x2=28.035 //y2=5.155
cc_619 ( N_noxref_2_c_543_p N_noxref_25_c_3206_n ) capacitor c=6.98646e-19 \
 //x=27.695 //y=7.4 //x2=28.035 //y2=5.155
cc_620 ( N_noxref_2_c_314_n N_noxref_25_c_3206_n ) capacitor c=0.00179956f \
 //x=28.12 //y=7.4 //x2=28.035 //y2=5.155
cc_621 ( N_noxref_2_M53_noxref_d N_noxref_25_c_3206_n ) capacitor c=0.0119114f \
 //x=27.635 //y=5.02 //x2=28.035 //y2=5.155
cc_622 ( N_noxref_2_c_314_n N_noxref_25_c_3210_n ) capacitor c=0.046173f \
 //x=28.12 //y=7.4 //x2=28.12 //y2=5.07
cc_623 ( N_noxref_2_c_320_p N_noxref_25_M48_noxref_d ) capacitor c=0.00294223f \
 //x=28.12 //y=7.4 //x2=25.435 //y2=5.02
cc_624 ( N_noxref_2_c_609_p N_noxref_25_M48_noxref_d ) capacitor c=0.0138437f \
 //x=25.935 //y=7.4 //x2=25.435 //y2=5.02
cc_625 ( N_noxref_2_M49_noxref_d N_noxref_25_M48_noxref_d ) capacitor \
 c=0.0664752f //x=25.875 //y=5.02 //x2=25.435 //y2=5.02
cc_626 ( N_noxref_2_c_320_p N_noxref_25_M50_noxref_d ) capacitor c=0.00294223f \
 //x=28.12 //y=7.4 //x2=26.315 //y2=5.02
cc_627 ( N_noxref_2_c_504_p N_noxref_25_M50_noxref_d ) capacitor c=0.0138437f \
 //x=26.815 //y=7.4 //x2=26.315 //y2=5.02
cc_628 ( N_noxref_2_c_314_n N_noxref_25_M50_noxref_d ) capacitor c=4.9285e-19 \
 //x=28.12 //y=7.4 //x2=26.315 //y2=5.02
cc_629 ( N_noxref_2_M48_noxref_s N_noxref_25_M50_noxref_d ) capacitor \
 c=0.00130656f //x=25.005 //y=5.02 //x2=26.315 //y2=5.02
cc_630 ( N_noxref_2_M49_noxref_d N_noxref_25_M50_noxref_d ) capacitor \
 c=0.0664752f //x=25.875 //y=5.02 //x2=26.315 //y2=5.02
cc_631 ( N_noxref_2_M51_noxref_d N_noxref_25_M50_noxref_d ) capacitor \
 c=0.0664752f //x=26.755 //y=5.02 //x2=26.315 //y2=5.02
cc_632 ( N_noxref_2_c_320_p N_noxref_25_M52_noxref_d ) capacitor c=0.00293548f \
 //x=28.12 //y=7.4 //x2=27.195 //y2=5.02
cc_633 ( N_noxref_2_c_543_p N_noxref_25_M52_noxref_d ) capacitor c=0.0137718f \
 //x=27.695 //y=7.4 //x2=27.195 //y2=5.02
cc_634 ( N_noxref_2_c_314_n N_noxref_25_M52_noxref_d ) capacitor c=0.00963505f \
 //x=28.12 //y=7.4 //x2=27.195 //y2=5.02
cc_635 ( N_noxref_2_M51_noxref_d N_noxref_25_M52_noxref_d ) capacitor \
 c=0.0664752f //x=26.755 //y=5.02 //x2=27.195 //y2=5.02
cc_636 ( N_noxref_2_M53_noxref_d N_noxref_25_M52_noxref_d ) capacitor \
 c=0.0664752f //x=27.635 //y=5.02 //x2=27.195 //y2=5.02
cc_637 ( N_noxref_3_c_646_n N_noxref_4_c_882_n ) capacitor c=0.00564994f \
 //x=10.615 //y=2.59 //x2=13.805 //y2=2.59
cc_638 ( N_noxref_3_M31_noxref_g N_noxref_4_c_897_n ) capacitor c=0.0168349f \
 //x=11.37 //y=6.02 //x2=11.945 //y2=5.155
cc_639 ( N_noxref_3_M30_noxref_g N_noxref_4_c_901_n ) capacitor c=0.0213876f \
 //x=10.93 //y=6.02 //x2=11.235 //y2=5.155
cc_640 ( N_noxref_3_c_724_p N_noxref_4_c_901_n ) capacitor c=0.00428486f \
 //x=11.295 //y=4.79 //x2=11.235 //y2=5.155
cc_641 ( N_noxref_3_M31_noxref_g N_noxref_4_M30_noxref_d ) capacitor \
 c=0.0180032f //x=11.37 //y=6.02 //x2=11.005 //y2=5.02
cc_642 ( N_noxref_3_c_646_n N_noxref_5_c_1045_n ) capacitor c=0.0035915f \
 //x=10.615 //y=2.59 //x2=16.535 //y2=4.44
cc_643 ( N_noxref_3_c_651_n N_noxref_5_c_1045_n ) capacitor c=0.0232115f \
 //x=10.73 //y=2.08 //x2=16.535 //y2=4.44
cc_644 ( N_noxref_3_c_704_n N_noxref_5_c_1045_n ) capacitor c=0.0169569f \
 //x=11.005 //y=4.79 //x2=16.535 //y2=4.44
cc_645 ( N_noxref_3_c_646_n N_noxref_5_c_1056_n ) capacitor c=3.86873e-19 \
 //x=10.615 //y=2.59 //x2=7.145 //y2=4.44
cc_646 ( N_noxref_3_c_650_n N_noxref_5_c_1056_n ) capacitor c=0.00551083f \
 //x=5.92 //y=2.08 //x2=7.145 //y2=4.44
cc_647 ( N_noxref_3_c_646_n N_noxref_5_c_1043_n ) capacitor c=0.0213409f \
 //x=10.615 //y=2.59 //x2=7.03 //y2=2.08
cc_648 ( N_noxref_3_c_647_n N_noxref_5_c_1043_n ) capacitor c=9.95819e-19 \
 //x=6.035 //y=2.59 //x2=7.03 //y2=2.08
cc_649 ( N_noxref_3_c_649_n N_noxref_5_c_1043_n ) capacitor c=4.79817e-19 \
 //x=4.07 //y=2.59 //x2=7.03 //y2=2.08
cc_650 ( N_noxref_3_c_650_n N_noxref_5_c_1043_n ) capacitor c=0.0491539f \
 //x=5.92 //y=2.08 //x2=7.03 //y2=2.08
cc_651 ( N_noxref_3_c_656_n N_noxref_5_c_1043_n ) capacitor c=0.00210802f \
 //x=5.62 //y=1.915 //x2=7.03 //y2=2.08
cc_652 ( N_noxref_3_c_736_p N_noxref_5_c_1043_n ) capacitor c=0.00147352f \
 //x=6.485 //y=4.79 //x2=7.03 //y2=2.08
cc_653 ( N_noxref_3_c_702_n N_noxref_5_c_1043_n ) capacitor c=0.00141297f \
 //x=6.195 //y=4.79 //x2=7.03 //y2=2.08
cc_654 ( N_noxref_3_M24_noxref_g N_noxref_5_M26_noxref_g ) capacitor \
 c=0.0105869f //x=6.12 //y=6.02 //x2=7 //y2=6.02
cc_655 ( N_noxref_3_M25_noxref_g N_noxref_5_M26_noxref_g ) capacitor \
 c=0.10632f //x=6.56 //y=6.02 //x2=7 //y2=6.02
cc_656 ( N_noxref_3_M25_noxref_g N_noxref_5_M27_noxref_g ) capacitor \
 c=0.0101598f //x=6.56 //y=6.02 //x2=7.44 //y2=6.02
cc_657 ( N_noxref_3_c_652_n N_noxref_5_c_1084_n ) capacitor c=5.72482e-19 \
 //x=5.62 //y=0.875 //x2=6.595 //y2=0.91
cc_658 ( N_noxref_3_c_654_n N_noxref_5_c_1084_n ) capacitor c=0.00149976f \
 //x=5.62 //y=1.22 //x2=6.595 //y2=0.91
cc_659 ( N_noxref_3_c_659_n N_noxref_5_c_1084_n ) capacitor c=0.0160123f \
 //x=6.15 //y=0.875 //x2=6.595 //y2=0.91
cc_660 ( N_noxref_3_c_655_n N_noxref_5_c_1087_n ) capacitor c=0.00111227f \
 //x=5.62 //y=1.53 //x2=6.595 //y2=1.22
cc_661 ( N_noxref_3_c_661_n N_noxref_5_c_1087_n ) capacitor c=0.0124075f \
 //x=6.15 //y=1.22 //x2=6.595 //y2=1.22
cc_662 ( N_noxref_3_c_659_n N_noxref_5_c_1089_n ) capacitor c=0.00103227f \
 //x=6.15 //y=0.875 //x2=7.12 //y2=0.91
cc_663 ( N_noxref_3_c_661_n N_noxref_5_c_1090_n ) capacitor c=0.0010154f \
 //x=6.15 //y=1.22 //x2=7.12 //y2=1.22
cc_664 ( N_noxref_3_c_661_n N_noxref_5_c_1091_n ) capacitor c=9.23422e-19 \
 //x=6.15 //y=1.22 //x2=7.12 //y2=1.45
cc_665 ( N_noxref_3_c_650_n N_noxref_5_c_1092_n ) capacitor c=0.00203769f \
 //x=5.92 //y=2.08 //x2=7.12 //y2=1.915
cc_666 ( N_noxref_3_c_656_n N_noxref_5_c_1092_n ) capacitor c=0.00834532f \
 //x=5.62 //y=1.915 //x2=7.12 //y2=1.915
cc_667 ( N_noxref_3_c_650_n N_noxref_5_c_1094_n ) capacitor c=0.00183762f \
 //x=5.92 //y=2.08 //x2=7.03 //y2=4.7
cc_668 ( N_noxref_3_c_736_p N_noxref_5_c_1094_n ) capacitor c=0.0168581f \
 //x=6.485 //y=4.79 //x2=7.03 //y2=4.7
cc_669 ( N_noxref_3_c_702_n N_noxref_5_c_1094_n ) capacitor c=0.00484466f \
 //x=6.195 //y=4.79 //x2=7.03 //y2=4.7
cc_670 ( N_noxref_3_c_644_n N_noxref_6_c_1247_n ) capacitor c=0.071918f \
 //x=5.805 //y=2.59 //x2=8.765 //y2=3.33
cc_671 ( N_noxref_3_c_645_n N_noxref_6_c_1247_n ) capacitor c=0.0138373f \
 //x=4.185 //y=2.59 //x2=8.765 //y2=3.33
cc_672 ( N_noxref_3_c_646_n N_noxref_6_c_1247_n ) capacitor c=0.115668f \
 //x=10.615 //y=2.59 //x2=8.765 //y2=3.33
cc_673 ( N_noxref_3_c_647_n N_noxref_6_c_1247_n ) capacitor c=0.0125712f \
 //x=6.035 //y=2.59 //x2=8.765 //y2=3.33
cc_674 ( N_noxref_3_c_683_n N_noxref_6_c_1247_n ) capacitor c=0.00843775f \
 //x=3.985 //y=5.155 //x2=8.765 //y2=3.33
cc_675 ( N_noxref_3_c_649_n N_noxref_6_c_1247_n ) capacitor c=0.0271263f \
 //x=4.07 //y=2.59 //x2=8.765 //y2=3.33
cc_676 ( N_noxref_3_c_650_n N_noxref_6_c_1247_n ) capacitor c=0.0278638f \
 //x=5.92 //y=2.08 //x2=8.765 //y2=3.33
cc_677 ( N_noxref_3_c_679_n N_noxref_6_c_1266_n ) capacitor c=3.71839e-19 \
 //x=3.205 //y=5.155 //x2=3.445 //y2=3.33
cc_678 ( N_noxref_3_c_683_n N_noxref_6_c_1266_n ) capacitor c=5.21082e-19 \
 //x=3.985 //y=5.155 //x2=3.445 //y2=3.33
cc_679 ( N_noxref_3_c_649_n N_noxref_6_c_1266_n ) capacitor c=0.00179385f \
 //x=4.07 //y=2.59 //x2=3.445 //y2=3.33
cc_680 ( N_noxref_3_c_764_p N_noxref_6_c_1266_n ) capacitor c=4.12695e-19 \
 //x=3.29 //y=5.155 //x2=3.445 //y2=3.33
cc_681 ( N_noxref_3_c_646_n N_noxref_6_c_1248_n ) capacitor c=0.0846302f \
 //x=10.615 //y=2.59 //x2=20.235 //y2=3.33
cc_682 ( N_noxref_3_c_651_n N_noxref_6_c_1248_n ) capacitor c=0.0224325f \
 //x=10.73 //y=2.08 //x2=20.235 //y2=3.33
cc_683 ( N_noxref_3_c_646_n N_noxref_6_c_1324_n ) capacitor c=0.0120889f \
 //x=10.615 //y=2.59 //x2=8.995 //y2=3.33
cc_684 ( N_noxref_3_c_651_n N_noxref_6_c_1324_n ) capacitor c=7.01366e-19 \
 //x=10.73 //y=2.08 //x2=8.995 //y2=3.33
cc_685 ( N_noxref_3_c_645_n N_noxref_6_c_1249_n ) capacitor c=0.00687545f \
 //x=4.185 //y=2.59 //x2=3.33 //y2=2.08
cc_686 ( N_noxref_3_c_649_n N_noxref_6_c_1249_n ) capacitor c=0.0861174f \
 //x=4.07 //y=2.59 //x2=3.33 //y2=2.08
cc_687 ( N_noxref_3_c_650_n N_noxref_6_c_1249_n ) capacitor c=8.632e-19 \
 //x=5.92 //y=2.08 //x2=3.33 //y2=2.08
cc_688 ( N_noxref_3_c_764_p N_noxref_6_c_1249_n ) capacitor c=0.0179147f \
 //x=3.29 //y=5.155 //x2=3.33 //y2=2.08
cc_689 ( N_noxref_3_M25_noxref_g N_noxref_6_c_1268_n ) capacitor c=0.0192001f \
 //x=6.56 //y=6.02 //x2=7.135 //y2=5.155
cc_690 ( N_noxref_3_c_683_n N_noxref_6_c_1272_n ) capacitor c=3.10026e-19 \
 //x=3.985 //y=5.155 //x2=6.425 //y2=5.155
cc_691 ( N_noxref_3_M24_noxref_g N_noxref_6_c_1272_n ) capacitor c=0.0213876f \
 //x=6.12 //y=6.02 //x2=6.425 //y2=5.155
cc_692 ( N_noxref_3_c_736_p N_noxref_6_c_1272_n ) capacitor c=0.0044314f \
 //x=6.485 //y=4.79 //x2=6.425 //y2=5.155
cc_693 ( N_noxref_3_c_646_n N_noxref_6_c_1282_n ) capacitor c=0.0192483f \
 //x=10.615 //y=2.59 //x2=8.88 //y2=3.33
cc_694 ( N_noxref_3_c_651_n N_noxref_6_c_1282_n ) capacitor c=0.013624f \
 //x=10.73 //y=2.08 //x2=8.88 //y2=3.33
cc_695 ( N_noxref_3_c_679_n N_noxref_6_M22_noxref_g ) capacitor c=0.0205444f \
 //x=3.205 //y=5.155 //x2=3.07 //y2=6.02
cc_696 ( N_noxref_3_M22_noxref_d N_noxref_6_M22_noxref_g ) capacitor \
 c=0.0180032f //x=3.145 //y=5.02 //x2=3.07 //y2=6.02
cc_697 ( N_noxref_3_c_683_n N_noxref_6_M23_noxref_g ) capacitor c=0.0218609f \
 //x=3.985 //y=5.155 //x2=3.51 //y2=6.02
cc_698 ( N_noxref_3_M22_noxref_d N_noxref_6_M23_noxref_g ) capacitor \
 c=0.0194246f //x=3.145 //y=5.02 //x2=3.51 //y2=6.02
cc_699 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1340_n ) capacitor c=0.00217566f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=0.915
cc_700 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1341_n ) capacitor c=0.0034598f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=1.26
cc_701 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1342_n ) capacitor c=0.00546784f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=1.57
cc_702 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1343_n ) capacitor c=0.00241102f \
 //x=3.395 //y=0.915 //x2=3.695 //y2=0.76
cc_703 ( N_noxref_3_c_648_n N_noxref_6_c_1344_n ) capacitor c=0.00371277f \
 //x=3.985 //y=1.665 //x2=3.695 //y2=1.415
cc_704 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1344_n ) capacitor c=0.0138621f \
 //x=3.395 //y=0.915 //x2=3.695 //y2=1.415
cc_705 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1346_n ) capacitor c=0.00219619f \
 //x=3.395 //y=0.915 //x2=3.85 //y2=0.915
cc_706 ( N_noxref_3_c_648_n N_noxref_6_c_1347_n ) capacitor c=0.00457401f \
 //x=3.985 //y=1.665 //x2=3.85 //y2=1.26
cc_707 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1347_n ) capacitor c=0.00603828f \
 //x=3.395 //y=0.915 //x2=3.85 //y2=1.26
cc_708 ( N_noxref_3_c_649_n N_noxref_6_c_1349_n ) capacitor c=0.00709342f \
 //x=4.07 //y=2.59 //x2=3.33 //y2=2.08
cc_709 ( N_noxref_3_c_649_n N_noxref_6_c_1350_n ) capacitor c=0.00283672f \
 //x=4.07 //y=2.59 //x2=3.33 //y2=1.915
cc_710 ( N_noxref_3_M2_noxref_d N_noxref_6_c_1350_n ) capacitor c=0.00661782f \
 //x=3.395 //y=0.915 //x2=3.33 //y2=1.915
cc_711 ( N_noxref_3_c_683_n N_noxref_6_c_1352_n ) capacitor c=0.00201851f \
 //x=3.985 //y=5.155 //x2=3.33 //y2=4.7
cc_712 ( N_noxref_3_c_649_n N_noxref_6_c_1352_n ) capacitor c=0.013693f \
 //x=4.07 //y=2.59 //x2=3.33 //y2=4.7
cc_713 ( N_noxref_3_c_764_p N_noxref_6_c_1352_n ) capacitor c=0.00476349f \
 //x=3.29 //y=5.155 //x2=3.33 //y2=4.7
cc_714 ( N_noxref_3_M25_noxref_g N_noxref_6_M24_noxref_d ) capacitor \
 c=0.0180032f //x=6.56 //y=6.02 //x2=6.195 //y2=5.02
cc_715 ( N_noxref_3_c_644_n N_noxref_7_c_1511_n ) capacitor c=0.143487f \
 //x=5.805 //y=2.59 //x2=17.645 //y2=2.22
cc_716 ( N_noxref_3_c_645_n N_noxref_7_c_1511_n ) capacitor c=0.0291301f \
 //x=4.185 //y=2.59 //x2=17.645 //y2=2.22
cc_717 ( N_noxref_3_c_646_n N_noxref_7_c_1511_n ) capacitor c=0.42762f \
 //x=10.615 //y=2.59 //x2=17.645 //y2=2.22
cc_718 ( N_noxref_3_c_647_n N_noxref_7_c_1511_n ) capacitor c=0.0264401f \
 //x=6.035 //y=2.59 //x2=17.645 //y2=2.22
cc_719 ( N_noxref_3_c_803_p N_noxref_7_c_1511_n ) capacitor c=0.016327f \
 //x=3.67 //y=1.665 //x2=17.645 //y2=2.22
cc_720 ( N_noxref_3_c_649_n N_noxref_7_c_1511_n ) capacitor c=0.0215653f \
 //x=4.07 //y=2.59 //x2=17.645 //y2=2.22
cc_721 ( N_noxref_3_c_650_n N_noxref_7_c_1511_n ) capacitor c=0.021104f \
 //x=5.92 //y=2.08 //x2=17.645 //y2=2.22
cc_722 ( N_noxref_3_c_651_n N_noxref_7_c_1511_n ) capacitor c=0.021104f \
 //x=10.73 //y=2.08 //x2=17.645 //y2=2.22
cc_723 ( N_noxref_3_c_807_p N_noxref_7_c_1511_n ) capacitor c=0.0103096f \
 //x=2.41 //y=5.155 //x2=17.645 //y2=2.22
cc_724 ( N_noxref_3_c_656_n N_noxref_7_c_1511_n ) capacitor c=0.011987f \
 //x=5.62 //y=1.915 //x2=17.645 //y2=2.22
cc_725 ( N_noxref_3_c_666_n N_noxref_7_c_1511_n ) capacitor c=0.011987f \
 //x=10.43 //y=1.915 //x2=17.645 //y2=2.22
cc_726 ( N_noxref_3_c_673_n N_noxref_7_c_1522_n ) capacitor c=9.18933e-19 \
 //x=2.325 //y=5.155 //x2=2.335 //y2=2.22
cc_727 ( N_noxref_3_c_673_n N_noxref_7_c_1528_n ) capacitor c=0.0148829f \
 //x=2.325 //y=5.155 //x2=2.22 //y2=2.08
cc_728 ( N_noxref_3_c_649_n N_noxref_7_c_1528_n ) capacitor c=0.00317604f \
 //x=4.07 //y=2.59 //x2=2.22 //y2=2.08
cc_729 ( N_noxref_3_c_673_n N_noxref_7_M20_noxref_g ) capacitor c=0.0169496f \
 //x=2.325 //y=5.155 //x2=2.19 //y2=6.02
cc_730 ( N_noxref_3_M20_noxref_d N_noxref_7_M20_noxref_g ) capacitor \
 c=0.0180032f //x=2.265 //y=5.02 //x2=2.19 //y2=6.02
cc_731 ( N_noxref_3_c_679_n N_noxref_7_M21_noxref_g ) capacitor c=0.0205444f \
 //x=3.205 //y=5.155 //x2=2.63 //y2=6.02
cc_732 ( N_noxref_3_M20_noxref_d N_noxref_7_M21_noxref_g ) capacitor \
 c=0.0180032f //x=2.265 //y=5.02 //x2=2.63 //y2=6.02
cc_733 ( N_noxref_3_c_807_p N_noxref_7_c_1566_n ) capacitor c=0.00441288f \
 //x=2.41 //y=5.155 //x2=2.555 //y2=4.79
cc_734 ( N_noxref_3_c_673_n N_noxref_7_c_1567_n ) capacitor c=0.00325274f \
 //x=2.325 //y=5.155 //x2=2.22 //y2=4.7
cc_735 ( N_noxref_3_c_651_n N_noxref_8_c_1847_n ) capacitor c=0.00526349f \
 //x=10.73 //y=2.08 //x2=11.955 //y2=2.96
cc_736 ( N_noxref_3_c_646_n N_noxref_8_c_1833_n ) capacitor c=0.00311593f \
 //x=10.615 //y=2.59 //x2=11.84 //y2=2.08
cc_737 ( N_noxref_3_c_651_n N_noxref_8_c_1833_n ) capacitor c=0.0460356f \
 //x=10.73 //y=2.08 //x2=11.84 //y2=2.08
cc_738 ( N_noxref_3_c_666_n N_noxref_8_c_1833_n ) capacitor c=0.00210802f \
 //x=10.43 //y=1.915 //x2=11.84 //y2=2.08
cc_739 ( N_noxref_3_c_724_p N_noxref_8_c_1833_n ) capacitor c=0.00147352f \
 //x=11.295 //y=4.79 //x2=11.84 //y2=2.08
cc_740 ( N_noxref_3_c_704_n N_noxref_8_c_1833_n ) capacitor c=0.00142741f \
 //x=11.005 //y=4.79 //x2=11.84 //y2=2.08
cc_741 ( N_noxref_3_M30_noxref_g N_noxref_8_M32_noxref_g ) capacitor \
 c=0.0105869f //x=10.93 //y=6.02 //x2=11.81 //y2=6.02
cc_742 ( N_noxref_3_M31_noxref_g N_noxref_8_M32_noxref_g ) capacitor \
 c=0.10632f //x=11.37 //y=6.02 //x2=11.81 //y2=6.02
cc_743 ( N_noxref_3_M31_noxref_g N_noxref_8_M33_noxref_g ) capacitor \
 c=0.0101598f //x=11.37 //y=6.02 //x2=12.25 //y2=6.02
cc_744 ( N_noxref_3_c_662_n N_noxref_8_c_1856_n ) capacitor c=5.72482e-19 \
 //x=10.43 //y=0.875 //x2=11.405 //y2=0.91
cc_745 ( N_noxref_3_c_664_n N_noxref_8_c_1856_n ) capacitor c=0.00149976f \
 //x=10.43 //y=1.22 //x2=11.405 //y2=0.91
cc_746 ( N_noxref_3_c_669_n N_noxref_8_c_1856_n ) capacitor c=0.0160123f \
 //x=10.96 //y=0.875 //x2=11.405 //y2=0.91
cc_747 ( N_noxref_3_c_665_n N_noxref_8_c_1859_n ) capacitor c=0.00111227f \
 //x=10.43 //y=1.53 //x2=11.405 //y2=1.22
cc_748 ( N_noxref_3_c_671_n N_noxref_8_c_1859_n ) capacitor c=0.0124075f \
 //x=10.96 //y=1.22 //x2=11.405 //y2=1.22
cc_749 ( N_noxref_3_c_669_n N_noxref_8_c_1861_n ) capacitor c=0.00103227f \
 //x=10.96 //y=0.875 //x2=11.93 //y2=0.91
cc_750 ( N_noxref_3_c_671_n N_noxref_8_c_1862_n ) capacitor c=0.0010154f \
 //x=10.96 //y=1.22 //x2=11.93 //y2=1.22
cc_751 ( N_noxref_3_c_671_n N_noxref_8_c_1863_n ) capacitor c=9.23422e-19 \
 //x=10.96 //y=1.22 //x2=11.93 //y2=1.45
cc_752 ( N_noxref_3_c_651_n N_noxref_8_c_1864_n ) capacitor c=0.00203769f \
 //x=10.73 //y=2.08 //x2=11.93 //y2=1.915
cc_753 ( N_noxref_3_c_666_n N_noxref_8_c_1864_n ) capacitor c=0.00834532f \
 //x=10.43 //y=1.915 //x2=11.93 //y2=1.915
cc_754 ( N_noxref_3_c_651_n N_noxref_8_c_1866_n ) capacitor c=0.00183762f \
 //x=10.73 //y=2.08 //x2=11.84 //y2=4.7
cc_755 ( N_noxref_3_c_724_p N_noxref_8_c_1866_n ) capacitor c=0.0168581f \
 //x=11.295 //y=4.79 //x2=11.84 //y2=4.7
cc_756 ( N_noxref_3_c_704_n N_noxref_8_c_1866_n ) capacitor c=0.00484466f \
 //x=11.005 //y=4.79 //x2=11.84 //y2=4.7
cc_757 ( N_noxref_3_c_646_n N_noxref_9_c_2034_n ) capacitor c=0.0121818f \
 //x=10.615 //y=2.59 //x2=12.835 //y2=3.7
cc_758 ( N_noxref_3_c_651_n N_noxref_9_c_2034_n ) capacitor c=0.0220679f \
 //x=10.73 //y=2.08 //x2=12.835 //y2=3.7
cc_759 ( N_noxref_3_c_646_n N_noxref_9_c_2090_n ) capacitor c=5.84956e-19 \
 //x=10.615 //y=2.59 //x2=8.255 //y2=3.7
cc_760 ( N_noxref_3_c_646_n N_noxref_9_c_2029_n ) capacitor c=0.0203032f \
 //x=10.615 //y=2.59 //x2=8.14 //y2=2.08
cc_761 ( N_noxref_3_c_650_n N_noxref_9_c_2029_n ) capacitor c=0.00146842f \
 //x=5.92 //y=2.08 //x2=8.14 //y2=2.08
cc_762 ( N_noxref_3_c_651_n N_noxref_9_c_2029_n ) capacitor c=8.30549e-19 \
 //x=10.73 //y=2.08 //x2=8.14 //y2=2.08
cc_763 ( N_noxref_3_c_651_n N_noxref_9_c_2030_n ) capacitor c=0.00134663f \
 //x=10.73 //y=2.08 //x2=12.95 //y2=2.08
cc_764 ( N_noxref_3_c_677_n N_noxref_10_M18_noxref_g ) capacitor c=0.0213876f \
 //x=1.615 //y=5.155 //x2=1.31 //y2=6.02
cc_765 ( N_noxref_3_c_673_n N_noxref_10_M19_noxref_g ) capacitor c=0.0204065f \
 //x=2.325 //y=5.155 //x2=1.75 //y2=6.02
cc_766 ( N_noxref_3_M18_noxref_d N_noxref_10_M19_noxref_g ) capacitor \
 c=0.0180032f //x=1.385 //y=5.02 //x2=1.75 //y2=6.02
cc_767 ( N_noxref_3_c_677_n N_noxref_10_c_2387_n ) capacitor c=0.00437952f \
 //x=1.615 //y=5.155 //x2=1.675 //y2=4.79
cc_768 ( N_noxref_3_M2_noxref_d N_noxref_11_M0_noxref_s ) capacitor \
 c=0.00309936f //x=3.395 //y=0.915 //x2=0.455 //y2=0.375
cc_769 ( N_noxref_3_c_648_n N_noxref_12_c_2473_n ) capacitor c=0.00457167f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_770 ( N_noxref_3_M2_noxref_d N_noxref_12_c_2473_n ) capacitor c=0.0115903f \
 //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_771 ( N_noxref_3_c_803_p N_noxref_12_c_2484_n ) capacitor c=0.0200405f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_772 ( N_noxref_3_M2_noxref_d N_noxref_12_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_773 ( N_noxref_3_c_648_n N_noxref_12_M2_noxref_s ) capacitor c=0.0184051f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_774 ( N_noxref_3_M2_noxref_d N_noxref_12_M2_noxref_s ) capacitor \
 c=0.0426368f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
cc_775 ( N_noxref_3_c_648_n N_noxref_13_c_2537_n ) capacitor c=3.84569e-19 \
 //x=3.985 //y=1.665 //x2=5.4 //y2=1.505
cc_776 ( N_noxref_3_c_656_n N_noxref_13_c_2537_n ) capacitor c=0.0034165f \
 //x=5.62 //y=1.915 //x2=5.4 //y2=1.505
cc_777 ( N_noxref_3_c_650_n N_noxref_13_c_2521_n ) capacitor c=0.0119952f \
 //x=5.92 //y=2.08 //x2=6.285 //y2=1.59
cc_778 ( N_noxref_3_c_655_n N_noxref_13_c_2521_n ) capacitor c=0.00697148f \
 //x=5.62 //y=1.53 //x2=6.285 //y2=1.59
cc_779 ( N_noxref_3_c_656_n N_noxref_13_c_2521_n ) capacitor c=0.0204849f \
 //x=5.62 //y=1.915 //x2=6.285 //y2=1.59
cc_780 ( N_noxref_3_c_658_n N_noxref_13_c_2521_n ) capacitor c=0.00610316f \
 //x=5.995 //y=1.375 //x2=6.285 //y2=1.59
cc_781 ( N_noxref_3_c_661_n N_noxref_13_c_2521_n ) capacitor c=0.00698822f \
 //x=6.15 //y=1.22 //x2=6.285 //y2=1.59
cc_782 ( N_noxref_3_c_652_n N_noxref_13_M3_noxref_s ) capacitor c=0.0327271f \
 //x=5.62 //y=0.875 //x2=5.265 //y2=0.375
cc_783 ( N_noxref_3_c_655_n N_noxref_13_M3_noxref_s ) capacitor c=7.99997e-19 \
 //x=5.62 //y=1.53 //x2=5.265 //y2=0.375
cc_784 ( N_noxref_3_c_656_n N_noxref_13_M3_noxref_s ) capacitor c=0.00122123f \
 //x=5.62 //y=1.915 //x2=5.265 //y2=0.375
cc_785 ( N_noxref_3_c_659_n N_noxref_13_M3_noxref_s ) capacitor c=0.0121427f \
 //x=6.15 //y=0.875 //x2=5.265 //y2=0.375
cc_786 ( N_noxref_3_M2_noxref_d N_noxref_13_M3_noxref_s ) capacitor \
 c=2.55333e-19 //x=3.395 //y=0.915 //x2=5.265 //y2=0.375
cc_787 ( N_noxref_3_c_666_n N_noxref_15_c_2641_n ) capacitor c=0.0034165f \
 //x=10.43 //y=1.915 //x2=10.21 //y2=1.505
cc_788 ( N_noxref_3_c_651_n N_noxref_15_c_2625_n ) capacitor c=0.0115578f \
 //x=10.73 //y=2.08 //x2=11.095 //y2=1.59
cc_789 ( N_noxref_3_c_665_n N_noxref_15_c_2625_n ) capacitor c=0.00697148f \
 //x=10.43 //y=1.53 //x2=11.095 //y2=1.59
cc_790 ( N_noxref_3_c_666_n N_noxref_15_c_2625_n ) capacitor c=0.0204849f \
 //x=10.43 //y=1.915 //x2=11.095 //y2=1.59
cc_791 ( N_noxref_3_c_668_n N_noxref_15_c_2625_n ) capacitor c=0.00610316f \
 //x=10.805 //y=1.375 //x2=11.095 //y2=1.59
cc_792 ( N_noxref_3_c_671_n N_noxref_15_c_2625_n ) capacitor c=0.00698822f \
 //x=10.96 //y=1.22 //x2=11.095 //y2=1.59
cc_793 ( N_noxref_3_c_662_n N_noxref_15_M6_noxref_s ) capacitor c=0.0327271f \
 //x=10.43 //y=0.875 //x2=10.075 //y2=0.375
cc_794 ( N_noxref_3_c_665_n N_noxref_15_M6_noxref_s ) capacitor c=7.99997e-19 \
 //x=10.43 //y=1.53 //x2=10.075 //y2=0.375
cc_795 ( N_noxref_3_c_666_n N_noxref_15_M6_noxref_s ) capacitor c=0.00122123f \
 //x=10.43 //y=1.915 //x2=10.075 //y2=0.375
cc_796 ( N_noxref_3_c_669_n N_noxref_15_M6_noxref_s ) capacitor c=0.0121427f \
 //x=10.96 //y=0.875 //x2=10.075 //y2=0.375
cc_797 ( N_noxref_4_c_897_n N_noxref_5_c_1045_n ) capacitor c=0.032141f \
 //x=11.945 //y=5.155 //x2=16.535 //y2=4.44
cc_798 ( N_noxref_4_c_901_n N_noxref_5_c_1045_n ) capacitor c=0.0230136f \
 //x=11.235 //y=5.155 //x2=16.535 //y2=4.44
cc_799 ( N_noxref_4_c_907_n N_noxref_5_c_1045_n ) capacitor c=0.0183122f \
 //x=13.605 //y=5.155 //x2=16.535 //y2=4.44
cc_800 ( N_noxref_4_c_884_n N_noxref_5_c_1045_n ) capacitor c=0.023368f \
 //x=13.69 //y=2.59 //x2=16.535 //y2=4.44
cc_801 ( N_noxref_4_c_885_n N_noxref_5_c_1045_n ) capacitor c=0.0247443f \
 //x=15.54 //y=2.08 //x2=16.535 //y2=4.44
cc_802 ( N_noxref_4_c_919_n N_noxref_5_c_1045_n ) capacitor c=0.0171124f \
 //x=15.815 //y=4.79 //x2=16.535 //y2=4.44
cc_803 ( N_noxref_4_c_881_n N_noxref_5_c_1044_n ) capacitor c=0.00520283f \
 //x=15.425 //y=2.59 //x2=16.65 //y2=2.08
cc_804 ( N_noxref_4_c_884_n N_noxref_5_c_1044_n ) capacitor c=3.46098e-19 \
 //x=13.69 //y=2.59 //x2=16.65 //y2=2.08
cc_805 ( N_noxref_4_c_885_n N_noxref_5_c_1044_n ) capacitor c=0.0446069f \
 //x=15.54 //y=2.08 //x2=16.65 //y2=2.08
cc_806 ( N_noxref_4_c_890_n N_noxref_5_c_1044_n ) capacitor c=0.00210802f \
 //x=15.24 //y=1.915 //x2=16.65 //y2=2.08
cc_807 ( N_noxref_4_c_951_p N_noxref_5_c_1044_n ) capacitor c=0.00147352f \
 //x=16.105 //y=4.79 //x2=16.65 //y2=2.08
cc_808 ( N_noxref_4_c_919_n N_noxref_5_c_1044_n ) capacitor c=0.00141297f \
 //x=15.815 //y=4.79 //x2=16.65 //y2=2.08
cc_809 ( N_noxref_4_M36_noxref_g N_noxref_5_M38_noxref_g ) capacitor \
 c=0.0105869f //x=15.74 //y=6.02 //x2=16.62 //y2=6.02
cc_810 ( N_noxref_4_M37_noxref_g N_noxref_5_M38_noxref_g ) capacitor \
 c=0.10632f //x=16.18 //y=6.02 //x2=16.62 //y2=6.02
cc_811 ( N_noxref_4_M37_noxref_g N_noxref_5_M39_noxref_g ) capacitor \
 c=0.0101598f //x=16.18 //y=6.02 //x2=17.06 //y2=6.02
cc_812 ( N_noxref_4_c_886_n N_noxref_5_c_1112_n ) capacitor c=5.72482e-19 \
 //x=15.24 //y=0.875 //x2=16.215 //y2=0.91
cc_813 ( N_noxref_4_c_888_n N_noxref_5_c_1112_n ) capacitor c=0.00149976f \
 //x=15.24 //y=1.22 //x2=16.215 //y2=0.91
cc_814 ( N_noxref_4_c_893_n N_noxref_5_c_1112_n ) capacitor c=0.0160123f \
 //x=15.77 //y=0.875 //x2=16.215 //y2=0.91
cc_815 ( N_noxref_4_c_889_n N_noxref_5_c_1115_n ) capacitor c=0.00111227f \
 //x=15.24 //y=1.53 //x2=16.215 //y2=1.22
cc_816 ( N_noxref_4_c_895_n N_noxref_5_c_1115_n ) capacitor c=0.0124075f \
 //x=15.77 //y=1.22 //x2=16.215 //y2=1.22
cc_817 ( N_noxref_4_c_893_n N_noxref_5_c_1117_n ) capacitor c=0.00103227f \
 //x=15.77 //y=0.875 //x2=16.74 //y2=0.91
cc_818 ( N_noxref_4_c_895_n N_noxref_5_c_1118_n ) capacitor c=0.0010154f \
 //x=15.77 //y=1.22 //x2=16.74 //y2=1.22
cc_819 ( N_noxref_4_c_895_n N_noxref_5_c_1119_n ) capacitor c=9.23422e-19 \
 //x=15.77 //y=1.22 //x2=16.74 //y2=1.45
cc_820 ( N_noxref_4_c_885_n N_noxref_5_c_1120_n ) capacitor c=0.00203769f \
 //x=15.54 //y=2.08 //x2=16.74 //y2=1.915
cc_821 ( N_noxref_4_c_890_n N_noxref_5_c_1120_n ) capacitor c=0.00834532f \
 //x=15.24 //y=1.915 //x2=16.74 //y2=1.915
cc_822 ( N_noxref_4_c_885_n N_noxref_5_c_1122_n ) capacitor c=0.00183762f \
 //x=15.54 //y=2.08 //x2=16.65 //y2=4.7
cc_823 ( N_noxref_4_c_951_p N_noxref_5_c_1122_n ) capacitor c=0.0168581f \
 //x=16.105 //y=4.79 //x2=16.65 //y2=4.7
cc_824 ( N_noxref_4_c_919_n N_noxref_5_c_1122_n ) capacitor c=0.00484466f \
 //x=15.815 //y=4.79 //x2=16.65 //y2=4.7
cc_825 ( N_noxref_4_c_881_n N_noxref_6_c_1248_n ) capacitor c=0.0119023f \
 //x=15.425 //y=2.59 //x2=20.235 //y2=3.33
cc_826 ( N_noxref_4_c_882_n N_noxref_6_c_1248_n ) capacitor c=8.87672e-19 \
 //x=13.805 //y=2.59 //x2=20.235 //y2=3.33
cc_827 ( N_noxref_4_c_884_n N_noxref_6_c_1248_n ) capacitor c=0.018769f \
 //x=13.69 //y=2.59 //x2=20.235 //y2=3.33
cc_828 ( N_noxref_4_c_885_n N_noxref_6_c_1248_n ) capacitor c=0.0198064f \
 //x=15.54 //y=2.08 //x2=20.235 //y2=3.33
cc_829 ( N_noxref_4_c_901_n N_noxref_6_c_1278_n ) capacitor c=3.10026e-19 \
 //x=11.235 //y=5.155 //x2=8.795 //y2=5.155
cc_830 ( N_noxref_4_c_881_n N_noxref_7_c_1511_n ) capacitor c=0.172592f \
 //x=15.425 //y=2.59 //x2=17.645 //y2=2.22
cc_831 ( N_noxref_4_c_882_n N_noxref_7_c_1511_n ) capacitor c=0.0291301f \
 //x=13.805 //y=2.59 //x2=17.645 //y2=2.22
cc_832 ( N_noxref_4_c_976_p N_noxref_7_c_1511_n ) capacitor c=0.016327f \
 //x=13.29 //y=1.665 //x2=17.645 //y2=2.22
cc_833 ( N_noxref_4_c_884_n N_noxref_7_c_1511_n ) capacitor c=0.0215653f \
 //x=13.69 //y=2.59 //x2=17.645 //y2=2.22
cc_834 ( N_noxref_4_c_885_n N_noxref_7_c_1511_n ) capacitor c=0.021104f \
 //x=15.54 //y=2.08 //x2=17.645 //y2=2.22
cc_835 ( N_noxref_4_c_890_n N_noxref_7_c_1511_n ) capacitor c=0.011987f \
 //x=15.24 //y=1.915 //x2=17.645 //y2=2.22
cc_836 ( N_noxref_4_c_885_n N_noxref_7_c_1529_n ) capacitor c=0.00135141f \
 //x=15.54 //y=2.08 //x2=17.76 //y2=2.08
cc_837 ( N_noxref_4_c_881_n N_noxref_8_c_1827_n ) capacitor c=0.172781f \
 //x=15.425 //y=2.59 //x2=26.155 //y2=2.96
cc_838 ( N_noxref_4_c_882_n N_noxref_8_c_1827_n ) capacitor c=0.0293832f \
 //x=13.805 //y=2.59 //x2=26.155 //y2=2.96
cc_839 ( N_noxref_4_c_884_n N_noxref_8_c_1827_n ) capacitor c=0.0206007f \
 //x=13.69 //y=2.59 //x2=26.155 //y2=2.96
cc_840 ( N_noxref_4_c_885_n N_noxref_8_c_1827_n ) capacitor c=0.0216195f \
 //x=15.54 //y=2.08 //x2=26.155 //y2=2.96
cc_841 ( N_noxref_4_c_897_n N_noxref_8_c_1833_n ) capacitor c=0.0144268f \
 //x=11.945 //y=5.155 //x2=11.84 //y2=2.08
cc_842 ( N_noxref_4_c_884_n N_noxref_8_c_1833_n ) capacitor c=0.00256054f \
 //x=13.69 //y=2.59 //x2=11.84 //y2=2.08
cc_843 ( N_noxref_4_c_897_n N_noxref_8_M32_noxref_g ) capacitor c=0.0165266f \
 //x=11.945 //y=5.155 //x2=11.81 //y2=6.02
cc_844 ( N_noxref_4_M32_noxref_d N_noxref_8_M32_noxref_g ) capacitor \
 c=0.0180032f //x=11.885 //y=5.02 //x2=11.81 //y2=6.02
cc_845 ( N_noxref_4_c_903_n N_noxref_8_M33_noxref_g ) capacitor c=0.01736f \
 //x=12.825 //y=5.155 //x2=12.25 //y2=6.02
cc_846 ( N_noxref_4_M32_noxref_d N_noxref_8_M33_noxref_g ) capacitor \
 c=0.0180032f //x=11.885 //y=5.02 //x2=12.25 //y2=6.02
cc_847 ( N_noxref_4_c_991_p N_noxref_8_c_1879_n ) capacitor c=0.00426767f \
 //x=12.03 //y=5.155 //x2=12.175 //y2=4.79
cc_848 ( N_noxref_4_c_897_n N_noxref_8_c_1866_n ) capacitor c=0.00322054f \
 //x=11.945 //y=5.155 //x2=11.84 //y2=4.7
cc_849 ( N_noxref_4_c_884_n N_noxref_9_c_2035_n ) capacitor c=0.0211104f \
 //x=13.69 //y=2.59 //x2=18.385 //y2=3.7
cc_850 ( N_noxref_4_c_885_n N_noxref_9_c_2035_n ) capacitor c=0.022094f \
 //x=15.54 //y=2.08 //x2=18.385 //y2=3.7
cc_851 ( N_noxref_4_c_884_n N_noxref_9_c_2097_n ) capacitor c=0.00179385f \
 //x=13.69 //y=2.59 //x2=13.065 //y2=3.7
cc_852 ( N_noxref_4_c_882_n N_noxref_9_c_2030_n ) capacitor c=0.00456439f \
 //x=13.805 //y=2.59 //x2=12.95 //y2=2.08
cc_853 ( N_noxref_4_c_884_n N_noxref_9_c_2030_n ) capacitor c=0.0794482f \
 //x=13.69 //y=2.59 //x2=12.95 //y2=2.08
cc_854 ( N_noxref_4_c_885_n N_noxref_9_c_2030_n ) capacitor c=6.21485e-19 \
 //x=15.54 //y=2.08 //x2=12.95 //y2=2.08
cc_855 ( N_noxref_4_c_999_p N_noxref_9_c_2030_n ) capacitor c=0.016476f \
 //x=12.91 //y=5.155 //x2=12.95 //y2=2.08
cc_856 ( N_noxref_4_M37_noxref_g N_noxref_9_c_2045_n ) capacitor c=0.0168349f \
 //x=16.18 //y=6.02 //x2=16.755 //y2=5.155
cc_857 ( N_noxref_4_c_907_n N_noxref_9_c_2049_n ) capacitor c=3.10026e-19 \
 //x=13.605 //y=5.155 //x2=16.045 //y2=5.155
cc_858 ( N_noxref_4_M36_noxref_g N_noxref_9_c_2049_n ) capacitor c=0.0213876f \
 //x=15.74 //y=6.02 //x2=16.045 //y2=5.155
cc_859 ( N_noxref_4_c_951_p N_noxref_9_c_2049_n ) capacitor c=0.00428486f \
 //x=16.105 //y=4.79 //x2=16.045 //y2=5.155
cc_860 ( N_noxref_4_c_903_n N_noxref_9_M34_noxref_g ) capacitor c=0.01736f \
 //x=12.825 //y=5.155 //x2=12.69 //y2=6.02
cc_861 ( N_noxref_4_M34_noxref_d N_noxref_9_M34_noxref_g ) capacitor \
 c=0.0180032f //x=12.765 //y=5.02 //x2=12.69 //y2=6.02
cc_862 ( N_noxref_4_c_907_n N_noxref_9_M35_noxref_g ) capacitor c=0.0194981f \
 //x=13.605 //y=5.155 //x2=13.13 //y2=6.02
cc_863 ( N_noxref_4_M34_noxref_d N_noxref_9_M35_noxref_g ) capacitor \
 c=0.0194246f //x=12.765 //y=5.02 //x2=13.13 //y2=6.02
cc_864 ( N_noxref_4_M8_noxref_d N_noxref_9_c_2110_n ) capacitor c=0.00217566f \
 //x=13.015 //y=0.915 //x2=12.94 //y2=0.915
cc_865 ( N_noxref_4_M8_noxref_d N_noxref_9_c_2111_n ) capacitor c=0.0034598f \
 //x=13.015 //y=0.915 //x2=12.94 //y2=1.26
cc_866 ( N_noxref_4_M8_noxref_d N_noxref_9_c_2112_n ) capacitor c=0.00546784f \
 //x=13.015 //y=0.915 //x2=12.94 //y2=1.57
cc_867 ( N_noxref_4_M8_noxref_d N_noxref_9_c_2113_n ) capacitor c=0.00241102f \
 //x=13.015 //y=0.915 //x2=13.315 //y2=0.76
cc_868 ( N_noxref_4_c_883_n N_noxref_9_c_2114_n ) capacitor c=0.00371277f \
 //x=13.605 //y=1.665 //x2=13.315 //y2=1.415
cc_869 ( N_noxref_4_M8_noxref_d N_noxref_9_c_2114_n ) capacitor c=0.0138621f \
 //x=13.015 //y=0.915 //x2=13.315 //y2=1.415
cc_870 ( N_noxref_4_M8_noxref_d N_noxref_9_c_2116_n ) capacitor c=0.00219619f \
 //x=13.015 //y=0.915 //x2=13.47 //y2=0.915
cc_871 ( N_noxref_4_c_883_n N_noxref_9_c_2117_n ) capacitor c=0.00457401f \
 //x=13.605 //y=1.665 //x2=13.47 //y2=1.26
cc_872 ( N_noxref_4_M8_noxref_d N_noxref_9_c_2117_n ) capacitor c=0.00603828f \
 //x=13.015 //y=0.915 //x2=13.47 //y2=1.26
cc_873 ( N_noxref_4_c_884_n N_noxref_9_c_2119_n ) capacitor c=0.00731987f \
 //x=13.69 //y=2.59 //x2=12.95 //y2=2.08
cc_874 ( N_noxref_4_c_884_n N_noxref_9_c_2120_n ) capacitor c=0.00283672f \
 //x=13.69 //y=2.59 //x2=12.95 //y2=1.915
cc_875 ( N_noxref_4_M8_noxref_d N_noxref_9_c_2120_n ) capacitor c=0.00661782f \
 //x=13.015 //y=0.915 //x2=12.95 //y2=1.915
cc_876 ( N_noxref_4_c_907_n N_noxref_9_c_2122_n ) capacitor c=0.00201851f \
 //x=13.605 //y=5.155 //x2=12.95 //y2=4.7
cc_877 ( N_noxref_4_c_884_n N_noxref_9_c_2122_n ) capacitor c=0.013693f \
 //x=13.69 //y=2.59 //x2=12.95 //y2=4.7
cc_878 ( N_noxref_4_c_999_p N_noxref_9_c_2122_n ) capacitor c=0.00475601f \
 //x=12.91 //y=5.155 //x2=12.95 //y2=4.7
cc_879 ( N_noxref_4_M37_noxref_g N_noxref_9_M36_noxref_d ) capacitor \
 c=0.0180032f //x=16.18 //y=6.02 //x2=15.815 //y2=5.02
cc_880 ( N_noxref_4_M8_noxref_d N_noxref_15_M6_noxref_s ) capacitor \
 c=0.00309936f //x=13.015 //y=0.915 //x2=10.075 //y2=0.375
cc_881 ( N_noxref_4_c_883_n N_noxref_16_c_2681_n ) capacitor c=0.00457167f \
 //x=13.605 //y=1.665 //x2=13.605 //y2=0.54
cc_882 ( N_noxref_4_M8_noxref_d N_noxref_16_c_2681_n ) capacitor c=0.0115903f \
 //x=13.015 //y=0.915 //x2=13.605 //y2=0.54
cc_883 ( N_noxref_4_c_976_p N_noxref_16_c_2692_n ) capacitor c=0.0200405f \
 //x=13.29 //y=1.665 //x2=12.72 //y2=0.995
cc_884 ( N_noxref_4_M8_noxref_d N_noxref_16_M7_noxref_d ) capacitor \
 c=5.27807e-19 //x=13.015 //y=0.915 //x2=11.48 //y2=0.91
cc_885 ( N_noxref_4_c_883_n N_noxref_16_M8_noxref_s ) capacitor c=0.0184051f \
 //x=13.605 //y=1.665 //x2=12.585 //y2=0.375
cc_886 ( N_noxref_4_M8_noxref_d N_noxref_16_M8_noxref_s ) capacitor \
 c=0.0426368f //x=13.015 //y=0.915 //x2=12.585 //y2=0.375
cc_887 ( N_noxref_4_c_883_n N_noxref_17_c_2745_n ) capacitor c=3.84569e-19 \
 //x=13.605 //y=1.665 //x2=15.02 //y2=1.505
cc_888 ( N_noxref_4_c_890_n N_noxref_17_c_2745_n ) capacitor c=0.0034165f \
 //x=15.24 //y=1.915 //x2=15.02 //y2=1.505
cc_889 ( N_noxref_4_c_885_n N_noxref_17_c_2729_n ) capacitor c=0.0115578f \
 //x=15.54 //y=2.08 //x2=15.905 //y2=1.59
cc_890 ( N_noxref_4_c_889_n N_noxref_17_c_2729_n ) capacitor c=0.00697148f \
 //x=15.24 //y=1.53 //x2=15.905 //y2=1.59
cc_891 ( N_noxref_4_c_890_n N_noxref_17_c_2729_n ) capacitor c=0.0204849f \
 //x=15.24 //y=1.915 //x2=15.905 //y2=1.59
cc_892 ( N_noxref_4_c_892_n N_noxref_17_c_2729_n ) capacitor c=0.00610316f \
 //x=15.615 //y=1.375 //x2=15.905 //y2=1.59
cc_893 ( N_noxref_4_c_895_n N_noxref_17_c_2729_n ) capacitor c=0.00698822f \
 //x=15.77 //y=1.22 //x2=15.905 //y2=1.59
cc_894 ( N_noxref_4_c_886_n N_noxref_17_M9_noxref_s ) capacitor c=0.0327271f \
 //x=15.24 //y=0.875 //x2=14.885 //y2=0.375
cc_895 ( N_noxref_4_c_889_n N_noxref_17_M9_noxref_s ) capacitor c=7.99997e-19 \
 //x=15.24 //y=1.53 //x2=14.885 //y2=0.375
cc_896 ( N_noxref_4_c_890_n N_noxref_17_M9_noxref_s ) capacitor c=0.00122123f \
 //x=15.24 //y=1.915 //x2=14.885 //y2=0.375
cc_897 ( N_noxref_4_c_893_n N_noxref_17_M9_noxref_s ) capacitor c=0.0121427f \
 //x=15.77 //y=0.875 //x2=14.885 //y2=0.375
cc_898 ( N_noxref_4_M8_noxref_d N_noxref_17_M9_noxref_s ) capacitor \
 c=2.55333e-19 //x=13.015 //y=0.915 //x2=14.885 //y2=0.375
cc_899 ( N_noxref_5_c_1045_n N_noxref_6_c_1247_n ) capacitor c=0.0280154f \
 //x=16.535 //y=4.44 //x2=8.765 //y2=3.33
cc_900 ( N_noxref_5_c_1056_n N_noxref_6_c_1247_n ) capacitor c=0.00755976f \
 //x=7.145 //y=4.44 //x2=8.765 //y2=3.33
cc_901 ( N_noxref_5_c_1043_n N_noxref_6_c_1247_n ) capacitor c=0.025332f \
 //x=7.03 //y=2.08 //x2=8.765 //y2=3.33
cc_902 ( N_noxref_5_c_1045_n N_noxref_6_c_1248_n ) capacitor c=0.039007f \
 //x=16.535 //y=4.44 //x2=20.235 //y2=3.33
cc_903 ( N_noxref_5_c_1044_n N_noxref_6_c_1248_n ) capacitor c=0.0190562f \
 //x=16.65 //y=2.08 //x2=20.235 //y2=3.33
cc_904 ( N_noxref_5_c_1045_n N_noxref_6_c_1324_n ) capacitor c=3.53076e-19 \
 //x=16.535 //y=4.44 //x2=8.995 //y2=3.33
cc_905 ( N_noxref_5_c_1056_n N_noxref_6_c_1268_n ) capacitor c=0.00330099f \
 //x=7.145 //y=4.44 //x2=7.135 //y2=5.155
cc_906 ( N_noxref_5_c_1043_n N_noxref_6_c_1268_n ) capacitor c=0.0143918f \
 //x=7.03 //y=2.08 //x2=7.135 //y2=5.155
cc_907 ( N_noxref_5_M26_noxref_g N_noxref_6_c_1268_n ) capacitor c=0.016514f \
 //x=7 //y=6.02 //x2=7.135 //y2=5.155
cc_908 ( N_noxref_5_c_1094_n N_noxref_6_c_1268_n ) capacitor c=0.00322046f \
 //x=7.03 //y=4.7 //x2=7.135 //y2=5.155
cc_909 ( N_noxref_5_M27_noxref_g N_noxref_6_c_1274_n ) capacitor c=0.01736f \
 //x=7.44 //y=6.02 //x2=8.015 //y2=5.155
cc_910 ( N_noxref_5_c_1045_n N_noxref_6_c_1278_n ) capacitor c=0.0183122f \
 //x=16.535 //y=4.44 //x2=8.795 //y2=5.155
cc_911 ( N_noxref_5_c_1045_n N_noxref_6_c_1282_n ) capacitor c=0.023368f \
 //x=16.535 //y=4.44 //x2=8.88 //y2=3.33
cc_912 ( N_noxref_5_c_1043_n N_noxref_6_c_1282_n ) capacitor c=0.00275732f \
 //x=7.03 //y=2.08 //x2=8.88 //y2=3.33
cc_913 ( N_noxref_5_c_1045_n N_noxref_6_c_1375_n ) capacitor c=0.0311227f \
 //x=16.535 //y=4.44 //x2=7.22 //y2=5.155
cc_914 ( N_noxref_5_c_1140_p N_noxref_6_c_1375_n ) capacitor c=0.00426767f \
 //x=7.365 //y=4.79 //x2=7.22 //y2=5.155
cc_915 ( N_noxref_5_M26_noxref_g N_noxref_6_M26_noxref_d ) capacitor \
 c=0.0180032f //x=7 //y=6.02 //x2=7.075 //y2=5.02
cc_916 ( N_noxref_5_M27_noxref_g N_noxref_6_M26_noxref_d ) capacitor \
 c=0.0180032f //x=7.44 //y=6.02 //x2=7.075 //y2=5.02
cc_917 ( N_noxref_5_c_1043_n N_noxref_7_c_1511_n ) capacitor c=0.0193884f \
 //x=7.03 //y=2.08 //x2=17.645 //y2=2.22
cc_918 ( N_noxref_5_c_1044_n N_noxref_7_c_1511_n ) capacitor c=0.021729f \
 //x=16.65 //y=2.08 //x2=17.645 //y2=2.22
cc_919 ( N_noxref_5_c_1092_n N_noxref_7_c_1511_n ) capacitor c=0.00583058f \
 //x=7.12 //y=1.915 //x2=17.645 //y2=2.22
cc_920 ( N_noxref_5_c_1120_n N_noxref_7_c_1511_n ) capacitor c=0.00583058f \
 //x=16.74 //y=1.915 //x2=17.645 //y2=2.22
cc_921 ( N_noxref_5_c_1044_n N_noxref_7_c_1527_n ) capacitor c=0.00165648f \
 //x=16.65 //y=2.08 //x2=17.875 //y2=2.22
cc_922 ( N_noxref_5_c_1120_n N_noxref_7_c_1527_n ) capacitor c=2.3323e-19 \
 //x=16.74 //y=1.915 //x2=17.875 //y2=2.22
cc_923 ( N_noxref_5_c_1045_n N_noxref_7_c_1529_n ) capacitor c=0.00551083f \
 //x=16.535 //y=4.44 //x2=17.76 //y2=2.08
cc_924 ( N_noxref_5_c_1044_n N_noxref_7_c_1529_n ) capacitor c=0.0468207f \
 //x=16.65 //y=2.08 //x2=17.76 //y2=2.08
cc_925 ( N_noxref_5_c_1120_n N_noxref_7_c_1529_n ) capacitor c=0.00203728f \
 //x=16.74 //y=1.915 //x2=17.76 //y2=2.08
cc_926 ( N_noxref_5_c_1122_n N_noxref_7_c_1529_n ) capacitor c=0.00142741f \
 //x=16.65 //y=4.7 //x2=17.76 //y2=2.08
cc_927 ( N_noxref_5_M38_noxref_g N_noxref_7_M40_noxref_g ) capacitor \
 c=0.0101598f //x=16.62 //y=6.02 //x2=17.5 //y2=6.02
cc_928 ( N_noxref_5_M39_noxref_g N_noxref_7_M40_noxref_g ) capacitor \
 c=0.0602553f //x=17.06 //y=6.02 //x2=17.5 //y2=6.02
cc_929 ( N_noxref_5_M39_noxref_g N_noxref_7_M41_noxref_g ) capacitor \
 c=0.0101598f //x=17.06 //y=6.02 //x2=17.94 //y2=6.02
cc_930 ( N_noxref_5_c_1117_n N_noxref_7_c_1588_n ) capacitor c=0.00456962f \
 //x=16.74 //y=0.91 //x2=17.75 //y2=0.915
cc_931 ( N_noxref_5_c_1118_n N_noxref_7_c_1589_n ) capacitor c=0.00438372f \
 //x=16.74 //y=1.22 //x2=17.75 //y2=1.26
cc_932 ( N_noxref_5_c_1119_n N_noxref_7_c_1590_n ) capacitor c=0.00438372f \
 //x=16.74 //y=1.45 //x2=17.75 //y2=1.57
cc_933 ( N_noxref_5_c_1044_n N_noxref_7_c_1591_n ) capacitor c=0.00201097f \
 //x=16.65 //y=2.08 //x2=17.76 //y2=2.08
cc_934 ( N_noxref_5_c_1120_n N_noxref_7_c_1591_n ) capacitor c=0.00828003f \
 //x=16.74 //y=1.915 //x2=17.76 //y2=2.08
cc_935 ( N_noxref_5_c_1120_n N_noxref_7_c_1593_n ) capacitor c=0.00438372f \
 //x=16.74 //y=1.915 //x2=17.76 //y2=1.915
cc_936 ( N_noxref_5_c_1044_n N_noxref_7_c_1594_n ) capacitor c=0.00218014f \
 //x=16.65 //y=2.08 //x2=17.76 //y2=4.7
cc_937 ( N_noxref_5_c_1163_p N_noxref_7_c_1594_n ) capacitor c=0.0611812f \
 //x=16.985 //y=4.79 //x2=17.76 //y2=4.7
cc_938 ( N_noxref_5_c_1122_n N_noxref_7_c_1594_n ) capacitor c=0.00487508f \
 //x=16.65 //y=4.7 //x2=17.76 //y2=4.7
cc_939 ( N_noxref_5_c_1044_n N_noxref_8_c_1827_n ) capacitor c=0.021326f \
 //x=16.65 //y=2.08 //x2=26.155 //y2=2.96
cc_940 ( N_noxref_5_c_1045_n N_noxref_8_c_1833_n ) capacitor c=0.0233868f \
 //x=16.535 //y=4.44 //x2=11.84 //y2=2.08
cc_941 ( N_noxref_5_c_1045_n N_noxref_8_c_1879_n ) capacitor c=0.0085986f \
 //x=16.535 //y=4.44 //x2=12.175 //y2=4.79
cc_942 ( N_noxref_5_c_1045_n N_noxref_8_c_1866_n ) capacitor c=0.00293313f \
 //x=16.535 //y=4.44 //x2=11.84 //y2=4.7
cc_943 ( N_noxref_5_c_1045_n N_noxref_9_c_2034_n ) capacitor c=0.194918f \
 //x=16.535 //y=4.44 //x2=12.835 //y2=3.7
cc_944 ( N_noxref_5_c_1045_n N_noxref_9_c_2090_n ) capacitor c=0.0134983f \
 //x=16.535 //y=4.44 //x2=8.255 //y2=3.7
cc_945 ( N_noxref_5_c_1043_n N_noxref_9_c_2090_n ) capacitor c=0.00526349f \
 //x=7.03 //y=2.08 //x2=8.255 //y2=3.7
cc_946 ( N_noxref_5_c_1045_n N_noxref_9_c_2035_n ) capacitor c=0.162328f \
 //x=16.535 //y=4.44 //x2=18.385 //y2=3.7
cc_947 ( N_noxref_5_c_1044_n N_noxref_9_c_2035_n ) capacitor c=0.0216655f \
 //x=16.65 //y=2.08 //x2=18.385 //y2=3.7
cc_948 ( N_noxref_5_c_1163_p N_noxref_9_c_2035_n ) capacitor c=0.00525621f \
 //x=16.985 //y=4.79 //x2=18.385 //y2=3.7
cc_949 ( N_noxref_5_c_1045_n N_noxref_9_c_2097_n ) capacitor c=0.0121615f \
 //x=16.535 //y=4.44 //x2=13.065 //y2=3.7
cc_950 ( N_noxref_5_c_1045_n N_noxref_9_c_2029_n ) capacitor c=0.0226638f \
 //x=16.535 //y=4.44 //x2=8.14 //y2=2.08
cc_951 ( N_noxref_5_c_1056_n N_noxref_9_c_2029_n ) capacitor c=0.00153281f \
 //x=7.145 //y=4.44 //x2=8.14 //y2=2.08
cc_952 ( N_noxref_5_c_1043_n N_noxref_9_c_2029_n ) capacitor c=0.0469899f \
 //x=7.03 //y=2.08 //x2=8.14 //y2=2.08
cc_953 ( N_noxref_5_c_1092_n N_noxref_9_c_2029_n ) capacitor c=0.00205895f \
 //x=7.12 //y=1.915 //x2=8.14 //y2=2.08
cc_954 ( N_noxref_5_c_1094_n N_noxref_9_c_2029_n ) capacitor c=0.00142741f \
 //x=7.03 //y=4.7 //x2=8.14 //y2=2.08
cc_955 ( N_noxref_5_c_1045_n N_noxref_9_c_2030_n ) capacitor c=0.0226638f \
 //x=16.535 //y=4.44 //x2=12.95 //y2=2.08
cc_956 ( N_noxref_5_c_1045_n N_noxref_9_c_2045_n ) capacitor c=0.00241768f \
 //x=16.535 //y=4.44 //x2=16.755 //y2=5.155
cc_957 ( N_noxref_5_c_1044_n N_noxref_9_c_2045_n ) capacitor c=0.0143918f \
 //x=16.65 //y=2.08 //x2=16.755 //y2=5.155
cc_958 ( N_noxref_5_M38_noxref_g N_noxref_9_c_2045_n ) capacitor c=0.016514f \
 //x=16.62 //y=6.02 //x2=16.755 //y2=5.155
cc_959 ( N_noxref_5_c_1122_n N_noxref_9_c_2045_n ) capacitor c=0.00322046f \
 //x=16.65 //y=4.7 //x2=16.755 //y2=5.155
cc_960 ( N_noxref_5_c_1045_n N_noxref_9_c_2049_n ) capacitor c=0.0219114f \
 //x=16.535 //y=4.44 //x2=16.045 //y2=5.155
cc_961 ( N_noxref_5_M39_noxref_g N_noxref_9_c_2051_n ) capacitor c=0.019179f \
 //x=17.06 //y=6.02 //x2=17.635 //y2=5.155
cc_962 ( N_noxref_5_c_1044_n N_noxref_9_c_2059_n ) capacitor c=0.00302286f \
 //x=16.65 //y=2.08 //x2=18.5 //y2=3.7
cc_963 ( N_noxref_5_c_1045_n N_noxref_9_c_2146_n ) capacitor c=0.00101864f \
 //x=16.535 //y=4.44 //x2=16.84 //y2=5.155
cc_964 ( N_noxref_5_c_1163_p N_noxref_9_c_2146_n ) capacitor c=0.00440089f \
 //x=16.985 //y=4.79 //x2=16.84 //y2=5.155
cc_965 ( N_noxref_5_M26_noxref_g N_noxref_9_M28_noxref_g ) capacitor \
 c=0.0101598f //x=7 //y=6.02 //x2=7.88 //y2=6.02
cc_966 ( N_noxref_5_M27_noxref_g N_noxref_9_M28_noxref_g ) capacitor \
 c=0.0602553f //x=7.44 //y=6.02 //x2=7.88 //y2=6.02
cc_967 ( N_noxref_5_M27_noxref_g N_noxref_9_M29_noxref_g ) capacitor \
 c=0.0101598f //x=7.44 //y=6.02 //x2=8.32 //y2=6.02
cc_968 ( N_noxref_5_c_1089_n N_noxref_9_c_2151_n ) capacitor c=0.00456962f \
 //x=7.12 //y=0.91 //x2=8.13 //y2=0.915
cc_969 ( N_noxref_5_c_1090_n N_noxref_9_c_2152_n ) capacitor c=0.00438372f \
 //x=7.12 //y=1.22 //x2=8.13 //y2=1.26
cc_970 ( N_noxref_5_c_1091_n N_noxref_9_c_2153_n ) capacitor c=0.00438372f \
 //x=7.12 //y=1.45 //x2=8.13 //y2=1.57
cc_971 ( N_noxref_5_c_1043_n N_noxref_9_c_2154_n ) capacitor c=0.00201097f \
 //x=7.03 //y=2.08 //x2=8.14 //y2=2.08
cc_972 ( N_noxref_5_c_1092_n N_noxref_9_c_2154_n ) capacitor c=0.00828003f \
 //x=7.12 //y=1.915 //x2=8.14 //y2=2.08
cc_973 ( N_noxref_5_c_1092_n N_noxref_9_c_2156_n ) capacitor c=0.00438372f \
 //x=7.12 //y=1.915 //x2=8.14 //y2=1.915
cc_974 ( N_noxref_5_c_1045_n N_noxref_9_c_2157_n ) capacitor c=0.00988777f \
 //x=16.535 //y=4.44 //x2=8.14 //y2=4.7
cc_975 ( N_noxref_5_c_1043_n N_noxref_9_c_2157_n ) capacitor c=0.00218014f \
 //x=7.03 //y=2.08 //x2=8.14 //y2=4.7
cc_976 ( N_noxref_5_c_1140_p N_noxref_9_c_2157_n ) capacitor c=0.0611812f \
 //x=7.365 //y=4.79 //x2=8.14 //y2=4.7
cc_977 ( N_noxref_5_c_1094_n N_noxref_9_c_2157_n ) capacitor c=0.00487508f \
 //x=7.03 //y=4.7 //x2=8.14 //y2=4.7
cc_978 ( N_noxref_5_c_1045_n N_noxref_9_c_2122_n ) capacitor c=0.0111881f \
 //x=16.535 //y=4.44 //x2=12.95 //y2=4.7
cc_979 ( N_noxref_5_M38_noxref_g N_noxref_9_M38_noxref_d ) capacitor \
 c=0.0180032f //x=16.62 //y=6.02 //x2=16.695 //y2=5.02
cc_980 ( N_noxref_5_M39_noxref_g N_noxref_9_M38_noxref_d ) capacitor \
 c=0.0180032f //x=17.06 //y=6.02 //x2=16.695 //y2=5.02
cc_981 ( N_noxref_5_c_1084_n N_noxref_13_c_2528_n ) capacitor c=0.0167228f \
 //x=6.595 //y=0.91 //x2=7.255 //y2=0.54
cc_982 ( N_noxref_5_c_1089_n N_noxref_13_c_2528_n ) capacitor c=0.00534519f \
 //x=7.12 //y=0.91 //x2=7.255 //y2=0.54
cc_983 ( N_noxref_5_c_1043_n N_noxref_13_c_2551_n ) capacitor c=0.0120267f \
 //x=7.03 //y=2.08 //x2=7.255 //y2=1.59
cc_984 ( N_noxref_5_c_1087_n N_noxref_13_c_2551_n ) capacitor c=0.0157358f \
 //x=6.595 //y=1.22 //x2=7.255 //y2=1.59
cc_985 ( N_noxref_5_c_1092_n N_noxref_13_c_2551_n ) capacitor c=0.021347f \
 //x=7.12 //y=1.915 //x2=7.255 //y2=1.59
cc_986 ( N_noxref_5_c_1084_n N_noxref_13_M3_noxref_s ) capacitor c=0.00798959f \
 //x=6.595 //y=0.91 //x2=5.265 //y2=0.375
cc_987 ( N_noxref_5_c_1091_n N_noxref_13_M3_noxref_s ) capacitor c=0.00212176f \
 //x=7.12 //y=1.45 //x2=5.265 //y2=0.375
cc_988 ( N_noxref_5_c_1092_n N_noxref_13_M3_noxref_s ) capacitor c=0.00298115f \
 //x=7.12 //y=1.915 //x2=5.265 //y2=0.375
cc_989 ( N_noxref_5_c_1215_p N_noxref_14_c_2571_n ) capacitor c=2.14837e-19 \
 //x=6.965 //y=0.755 //x2=7.825 //y2=0.995
cc_990 ( N_noxref_5_c_1089_n N_noxref_14_c_2571_n ) capacitor c=0.00123426f \
 //x=7.12 //y=0.91 //x2=7.825 //y2=0.995
cc_991 ( N_noxref_5_c_1090_n N_noxref_14_c_2571_n ) capacitor c=0.0129288f \
 //x=7.12 //y=1.22 //x2=7.825 //y2=0.995
cc_992 ( N_noxref_5_c_1091_n N_noxref_14_c_2571_n ) capacitor c=0.00142359f \
 //x=7.12 //y=1.45 //x2=7.825 //y2=0.995
cc_993 ( N_noxref_5_c_1084_n N_noxref_14_M4_noxref_d ) capacitor c=0.00223875f \
 //x=6.595 //y=0.91 //x2=6.67 //y2=0.91
cc_994 ( N_noxref_5_c_1087_n N_noxref_14_M4_noxref_d ) capacitor c=0.00262485f \
 //x=6.595 //y=1.22 //x2=6.67 //y2=0.91
cc_995 ( N_noxref_5_c_1215_p N_noxref_14_M4_noxref_d ) capacitor c=0.00220746f \
 //x=6.965 //y=0.755 //x2=6.67 //y2=0.91
cc_996 ( N_noxref_5_c_1222_p N_noxref_14_M4_noxref_d ) capacitor c=0.00194798f \
 //x=6.965 //y=1.375 //x2=6.67 //y2=0.91
cc_997 ( N_noxref_5_c_1089_n N_noxref_14_M4_noxref_d ) capacitor c=0.00198465f \
 //x=7.12 //y=0.91 //x2=6.67 //y2=0.91
cc_998 ( N_noxref_5_c_1090_n N_noxref_14_M4_noxref_d ) capacitor c=0.00128384f \
 //x=7.12 //y=1.22 //x2=6.67 //y2=0.91
cc_999 ( N_noxref_5_c_1089_n N_noxref_14_M5_noxref_s ) capacitor c=7.21316e-19 \
 //x=7.12 //y=0.91 //x2=7.775 //y2=0.375
cc_1000 ( N_noxref_5_c_1090_n N_noxref_14_M5_noxref_s ) capacitor \
 c=0.00348171f //x=7.12 //y=1.22 //x2=7.775 //y2=0.375
cc_1001 ( N_noxref_5_c_1112_n N_noxref_17_c_2736_n ) capacitor c=0.0167228f \
 //x=16.215 //y=0.91 //x2=16.875 //y2=0.54
cc_1002 ( N_noxref_5_c_1117_n N_noxref_17_c_2736_n ) capacitor c=0.00534519f \
 //x=16.74 //y=0.91 //x2=16.875 //y2=0.54
cc_1003 ( N_noxref_5_c_1044_n N_noxref_17_c_2759_n ) capacitor c=0.0117694f \
 //x=16.65 //y=2.08 //x2=16.875 //y2=1.59
cc_1004 ( N_noxref_5_c_1115_n N_noxref_17_c_2759_n ) capacitor c=0.0157358f \
 //x=16.215 //y=1.22 //x2=16.875 //y2=1.59
cc_1005 ( N_noxref_5_c_1120_n N_noxref_17_c_2759_n ) capacitor c=0.021347f \
 //x=16.74 //y=1.915 //x2=16.875 //y2=1.59
cc_1006 ( N_noxref_5_c_1112_n N_noxref_17_M9_noxref_s ) capacitor \
 c=0.00798959f //x=16.215 //y=0.91 //x2=14.885 //y2=0.375
cc_1007 ( N_noxref_5_c_1119_n N_noxref_17_M9_noxref_s ) capacitor \
 c=0.00212176f //x=16.74 //y=1.45 //x2=14.885 //y2=0.375
cc_1008 ( N_noxref_5_c_1120_n N_noxref_17_M9_noxref_s ) capacitor \
 c=0.00298115f //x=16.74 //y=1.915 //x2=14.885 //y2=0.375
cc_1009 ( N_noxref_5_c_1235_p N_noxref_18_c_2779_n ) capacitor c=2.14837e-19 \
 //x=16.585 //y=0.755 //x2=17.445 //y2=0.995
cc_1010 ( N_noxref_5_c_1117_n N_noxref_18_c_2779_n ) capacitor c=0.00123426f \
 //x=16.74 //y=0.91 //x2=17.445 //y2=0.995
cc_1011 ( N_noxref_5_c_1118_n N_noxref_18_c_2779_n ) capacitor c=0.0129288f \
 //x=16.74 //y=1.22 //x2=17.445 //y2=0.995
cc_1012 ( N_noxref_5_c_1119_n N_noxref_18_c_2779_n ) capacitor c=0.00142359f \
 //x=16.74 //y=1.45 //x2=17.445 //y2=0.995
cc_1013 ( N_noxref_5_c_1112_n N_noxref_18_M10_noxref_d ) capacitor \
 c=0.00223875f //x=16.215 //y=0.91 //x2=16.29 //y2=0.91
cc_1014 ( N_noxref_5_c_1115_n N_noxref_18_M10_noxref_d ) capacitor \
 c=0.00262485f //x=16.215 //y=1.22 //x2=16.29 //y2=0.91
cc_1015 ( N_noxref_5_c_1235_p N_noxref_18_M10_noxref_d ) capacitor \
 c=0.00220746f //x=16.585 //y=0.755 //x2=16.29 //y2=0.91
cc_1016 ( N_noxref_5_c_1242_p N_noxref_18_M10_noxref_d ) capacitor \
 c=0.00194798f //x=16.585 //y=1.375 //x2=16.29 //y2=0.91
cc_1017 ( N_noxref_5_c_1117_n N_noxref_18_M10_noxref_d ) capacitor \
 c=0.00198465f //x=16.74 //y=0.91 //x2=16.29 //y2=0.91
cc_1018 ( N_noxref_5_c_1118_n N_noxref_18_M10_noxref_d ) capacitor \
 c=0.00128384f //x=16.74 //y=1.22 //x2=16.29 //y2=0.91
cc_1019 ( N_noxref_5_c_1117_n N_noxref_18_M11_noxref_s ) capacitor \
 c=7.21316e-19 //x=16.74 //y=0.91 //x2=17.395 //y2=0.375
cc_1020 ( N_noxref_5_c_1118_n N_noxref_18_M11_noxref_s ) capacitor \
 c=0.00348171f //x=16.74 //y=1.22 //x2=17.395 //y2=0.375
cc_1021 ( N_noxref_6_c_1247_n N_noxref_7_c_1511_n ) capacitor c=0.0400111f \
 //x=8.765 //y=3.33 //x2=17.645 //y2=2.22
cc_1022 ( N_noxref_6_c_1266_n N_noxref_7_c_1511_n ) capacitor c=0.00767291f \
 //x=3.445 //y=3.33 //x2=17.645 //y2=2.22
cc_1023 ( N_noxref_6_c_1248_n N_noxref_7_c_1511_n ) capacitor c=0.0561264f \
 //x=20.235 //y=3.33 //x2=17.645 //y2=2.22
cc_1024 ( N_noxref_6_c_1324_n N_noxref_7_c_1511_n ) capacitor c=3.9466e-19 \
 //x=8.995 //y=3.33 //x2=17.645 //y2=2.22
cc_1025 ( N_noxref_6_c_1249_n N_noxref_7_c_1511_n ) capacitor c=0.0225728f \
 //x=3.33 //y=2.08 //x2=17.645 //y2=2.22
cc_1026 ( N_noxref_6_c_1384_p N_noxref_7_c_1511_n ) capacitor c=0.016327f \
 //x=8.48 //y=1.665 //x2=17.645 //y2=2.22
cc_1027 ( N_noxref_6_c_1282_n N_noxref_7_c_1511_n ) capacitor c=0.0197307f \
 //x=8.88 //y=3.33 //x2=17.645 //y2=2.22
cc_1028 ( N_noxref_6_c_1344_n N_noxref_7_c_1511_n ) capacitor c=3.13485e-19 \
 //x=3.695 //y=1.415 //x2=17.645 //y2=2.22
cc_1029 ( N_noxref_6_c_1349_n N_noxref_7_c_1511_n ) capacitor c=0.00583286f \
 //x=3.33 //y=2.08 //x2=17.645 //y2=2.22
cc_1030 ( N_noxref_6_c_1249_n N_noxref_7_c_1522_n ) capacitor c=0.00165648f \
 //x=3.33 //y=2.08 //x2=2.335 //y2=2.22
cc_1031 ( N_noxref_6_c_1349_n N_noxref_7_c_1522_n ) capacitor c=2.3323e-19 \
 //x=3.33 //y=2.08 //x2=2.335 //y2=2.22
cc_1032 ( N_noxref_6_c_1248_n N_noxref_7_c_1523_n ) capacitor c=0.014255f \
 //x=20.235 //y=3.33 //x2=21.345 //y2=2.22
cc_1033 ( N_noxref_6_c_1251_n N_noxref_7_c_1523_n ) capacitor c=0.0226137f \
 //x=20.35 //y=2.08 //x2=21.345 //y2=2.22
cc_1034 ( N_noxref_6_c_1256_n N_noxref_7_c_1523_n ) capacitor c=0.0121989f \
 //x=20.05 //y=1.915 //x2=21.345 //y2=2.22
cc_1035 ( N_noxref_6_c_1248_n N_noxref_7_c_1527_n ) capacitor c=4.86139e-19 \
 //x=20.235 //y=3.33 //x2=17.875 //y2=2.22
cc_1036 ( N_noxref_6_c_1266_n N_noxref_7_c_1528_n ) capacitor c=0.00526349f \
 //x=3.445 //y=3.33 //x2=2.22 //y2=2.08
cc_1037 ( N_noxref_6_c_1249_n N_noxref_7_c_1528_n ) capacitor c=0.0539839f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=2.08
cc_1038 ( N_noxref_6_c_1349_n N_noxref_7_c_1528_n ) capacitor c=0.0019893f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=2.08
cc_1039 ( N_noxref_6_c_1352_n N_noxref_7_c_1528_n ) capacitor c=0.00219458f \
 //x=3.33 //y=4.7 //x2=2.22 //y2=2.08
cc_1040 ( N_noxref_6_c_1248_n N_noxref_7_c_1529_n ) capacitor c=0.0180187f \
 //x=20.235 //y=3.33 //x2=17.76 //y2=2.08
cc_1041 ( N_noxref_6_c_1251_n N_noxref_7_c_1529_n ) capacitor c=7.78439e-19 \
 //x=20.35 //y=2.08 //x2=17.76 //y2=2.08
cc_1042 ( N_noxref_6_c_1248_n N_noxref_7_c_1530_n ) capacitor c=0.00526349f \
 //x=20.235 //y=3.33 //x2=21.46 //y2=2.08
cc_1043 ( N_noxref_6_c_1251_n N_noxref_7_c_1530_n ) capacitor c=0.0494371f \
 //x=20.35 //y=2.08 //x2=21.46 //y2=2.08
cc_1044 ( N_noxref_6_c_1256_n N_noxref_7_c_1530_n ) capacitor c=0.00208635f \
 //x=20.05 //y=1.915 //x2=21.46 //y2=2.08
cc_1045 ( N_noxref_6_c_1403_p N_noxref_7_c_1530_n ) capacitor c=0.00147352f \
 //x=20.915 //y=4.79 //x2=21.46 //y2=2.08
cc_1046 ( N_noxref_6_c_1294_n N_noxref_7_c_1530_n ) capacitor c=0.00142741f \
 //x=20.625 //y=4.79 //x2=21.46 //y2=2.08
cc_1047 ( N_noxref_6_M22_noxref_g N_noxref_7_M20_noxref_g ) capacitor \
 c=0.0101598f //x=3.07 //y=6.02 //x2=2.19 //y2=6.02
cc_1048 ( N_noxref_6_M22_noxref_g N_noxref_7_M21_noxref_g ) capacitor \
 c=0.0602553f //x=3.07 //y=6.02 //x2=2.63 //y2=6.02
cc_1049 ( N_noxref_6_M23_noxref_g N_noxref_7_M21_noxref_g ) capacitor \
 c=0.0101598f //x=3.51 //y=6.02 //x2=2.63 //y2=6.02
cc_1050 ( N_noxref_6_M42_noxref_g N_noxref_7_M44_noxref_g ) capacitor \
 c=0.0105869f //x=20.55 //y=6.02 //x2=21.43 //y2=6.02
cc_1051 ( N_noxref_6_M43_noxref_g N_noxref_7_M44_noxref_g ) capacitor \
 c=0.10632f //x=20.99 //y=6.02 //x2=21.43 //y2=6.02
cc_1052 ( N_noxref_6_M43_noxref_g N_noxref_7_M45_noxref_g ) capacitor \
 c=0.0101598f //x=20.99 //y=6.02 //x2=21.87 //y2=6.02
cc_1053 ( N_noxref_6_c_1340_n N_noxref_7_c_1629_n ) capacitor c=0.00456962f \
 //x=3.32 //y=0.915 //x2=2.31 //y2=0.91
cc_1054 ( N_noxref_6_c_1341_n N_noxref_7_c_1630_n ) capacitor c=0.00438372f \
 //x=3.32 //y=1.26 //x2=2.31 //y2=1.22
cc_1055 ( N_noxref_6_c_1342_n N_noxref_7_c_1631_n ) capacitor c=0.00438372f \
 //x=3.32 //y=1.57 //x2=2.31 //y2=1.45
cc_1056 ( N_noxref_6_c_1249_n N_noxref_7_c_1632_n ) capacitor c=0.00205895f \
 //x=3.33 //y=2.08 //x2=2.31 //y2=1.915
cc_1057 ( N_noxref_6_c_1349_n N_noxref_7_c_1632_n ) capacitor c=0.00828003f \
 //x=3.33 //y=2.08 //x2=2.31 //y2=1.915
cc_1058 ( N_noxref_6_c_1350_n N_noxref_7_c_1632_n ) capacitor c=0.00438372f \
 //x=3.33 //y=1.915 //x2=2.31 //y2=1.915
cc_1059 ( N_noxref_6_c_1352_n N_noxref_7_c_1566_n ) capacitor c=0.0611812f \
 //x=3.33 //y=4.7 //x2=2.555 //y2=4.79
cc_1060 ( N_noxref_6_c_1252_n N_noxref_7_c_1636_n ) capacitor c=5.72482e-19 \
 //x=20.05 //y=0.875 //x2=21.025 //y2=0.91
cc_1061 ( N_noxref_6_c_1254_n N_noxref_7_c_1636_n ) capacitor c=0.00149976f \
 //x=20.05 //y=1.22 //x2=21.025 //y2=0.91
cc_1062 ( N_noxref_6_c_1259_n N_noxref_7_c_1636_n ) capacitor c=0.0160123f \
 //x=20.58 //y=0.875 //x2=21.025 //y2=0.91
cc_1063 ( N_noxref_6_c_1255_n N_noxref_7_c_1639_n ) capacitor c=0.00111227f \
 //x=20.05 //y=1.53 //x2=21.025 //y2=1.22
cc_1064 ( N_noxref_6_c_1261_n N_noxref_7_c_1639_n ) capacitor c=0.0124075f \
 //x=20.58 //y=1.22 //x2=21.025 //y2=1.22
cc_1065 ( N_noxref_6_c_1259_n N_noxref_7_c_1641_n ) capacitor c=0.00103227f \
 //x=20.58 //y=0.875 //x2=21.55 //y2=0.91
cc_1066 ( N_noxref_6_c_1261_n N_noxref_7_c_1642_n ) capacitor c=0.0010154f \
 //x=20.58 //y=1.22 //x2=21.55 //y2=1.22
cc_1067 ( N_noxref_6_c_1261_n N_noxref_7_c_1643_n ) capacitor c=9.23422e-19 \
 //x=20.58 //y=1.22 //x2=21.55 //y2=1.45
cc_1068 ( N_noxref_6_c_1251_n N_noxref_7_c_1644_n ) capacitor c=0.00203769f \
 //x=20.35 //y=2.08 //x2=21.55 //y2=1.915
cc_1069 ( N_noxref_6_c_1256_n N_noxref_7_c_1644_n ) capacitor c=0.00834532f \
 //x=20.05 //y=1.915 //x2=21.55 //y2=1.915
cc_1070 ( N_noxref_6_c_1249_n N_noxref_7_c_1567_n ) capacitor c=0.00142741f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=4.7
cc_1071 ( N_noxref_6_c_1352_n N_noxref_7_c_1567_n ) capacitor c=0.00487508f \
 //x=3.33 //y=4.7 //x2=2.22 //y2=4.7
cc_1072 ( N_noxref_6_c_1251_n N_noxref_7_c_1648_n ) capacitor c=0.00183762f \
 //x=20.35 //y=2.08 //x2=21.46 //y2=4.7
cc_1073 ( N_noxref_6_c_1403_p N_noxref_7_c_1648_n ) capacitor c=0.0168581f \
 //x=20.915 //y=4.79 //x2=21.46 //y2=4.7
cc_1074 ( N_noxref_6_c_1294_n N_noxref_7_c_1648_n ) capacitor c=0.00484466f \
 //x=20.625 //y=4.79 //x2=21.46 //y2=4.7
cc_1075 ( N_noxref_6_c_1248_n N_noxref_8_c_1827_n ) capacitor c=0.756732f \
 //x=20.235 //y=3.33 //x2=26.155 //y2=2.96
cc_1076 ( N_noxref_6_c_1251_n N_noxref_8_c_1827_n ) capacitor c=0.0238838f \
 //x=20.35 //y=2.08 //x2=26.155 //y2=2.96
cc_1077 ( N_noxref_6_c_1248_n N_noxref_8_c_1847_n ) capacitor c=0.0292094f \
 //x=20.235 //y=3.33 //x2=11.955 //y2=2.96
cc_1078 ( N_noxref_6_c_1248_n N_noxref_8_c_1833_n ) capacitor c=0.0208912f \
 //x=20.235 //y=3.33 //x2=11.84 //y2=2.08
cc_1079 ( N_noxref_6_c_1282_n N_noxref_8_c_1833_n ) capacitor c=5.12802e-19 \
 //x=8.88 //y=3.33 //x2=11.84 //y2=2.08
cc_1080 ( N_noxref_6_c_1247_n N_noxref_9_c_2034_n ) capacitor c=0.0446157f \
 //x=8.765 //y=3.33 //x2=12.835 //y2=3.7
cc_1081 ( N_noxref_6_c_1248_n N_noxref_9_c_2034_n ) capacitor c=0.340407f \
 //x=20.235 //y=3.33 //x2=12.835 //y2=3.7
cc_1082 ( N_noxref_6_c_1324_n N_noxref_9_c_2034_n ) capacitor c=0.0268386f \
 //x=8.995 //y=3.33 //x2=12.835 //y2=3.7
cc_1083 ( N_noxref_6_c_1282_n N_noxref_9_c_2034_n ) capacitor c=0.0229188f \
 //x=8.88 //y=3.33 //x2=12.835 //y2=3.7
cc_1084 ( N_noxref_6_c_1247_n N_noxref_9_c_2090_n ) capacitor c=0.029444f \
 //x=8.765 //y=3.33 //x2=8.255 //y2=3.7
cc_1085 ( N_noxref_6_c_1282_n N_noxref_9_c_2090_n ) capacitor c=0.00179385f \
 //x=8.88 //y=3.33 //x2=8.255 //y2=3.7
cc_1086 ( N_noxref_6_c_1248_n N_noxref_9_c_2035_n ) capacitor c=0.468734f \
 //x=20.235 //y=3.33 //x2=18.385 //y2=3.7
cc_1087 ( N_noxref_6_c_1248_n N_noxref_9_c_2097_n ) capacitor c=0.026734f \
 //x=20.235 //y=3.33 //x2=13.065 //y2=3.7
cc_1088 ( N_noxref_6_c_1248_n N_noxref_9_c_2028_n ) capacitor c=0.176086f \
 //x=20.235 //y=3.33 //x2=27.265 //y2=3.7
cc_1089 ( N_noxref_6_c_1251_n N_noxref_9_c_2028_n ) capacitor c=0.0263175f \
 //x=20.35 //y=2.08 //x2=27.265 //y2=3.7
cc_1090 ( N_noxref_6_c_1294_n N_noxref_9_c_2028_n ) capacitor c=0.0129605f \
 //x=20.625 //y=4.79 //x2=27.265 //y2=3.7
cc_1091 ( N_noxref_6_c_1248_n N_noxref_9_c_2042_n ) capacitor c=0.0268461f \
 //x=20.235 //y=3.33 //x2=18.615 //y2=3.7
cc_1092 ( N_noxref_6_c_1251_n N_noxref_9_c_2042_n ) capacitor c=7.01366e-19 \
 //x=20.35 //y=2.08 //x2=18.615 //y2=3.7
cc_1093 ( N_noxref_6_c_1247_n N_noxref_9_c_2029_n ) capacitor c=0.0221941f \
 //x=8.765 //y=3.33 //x2=8.14 //y2=2.08
cc_1094 ( N_noxref_6_c_1324_n N_noxref_9_c_2029_n ) capacitor c=0.00179385f \
 //x=8.995 //y=3.33 //x2=8.14 //y2=2.08
cc_1095 ( N_noxref_6_c_1282_n N_noxref_9_c_2029_n ) capacitor c=0.0802836f \
 //x=8.88 //y=3.33 //x2=8.14 //y2=2.08
cc_1096 ( N_noxref_6_c_1454_p N_noxref_9_c_2029_n ) capacitor c=0.016476f \
 //x=8.1 //y=5.155 //x2=8.14 //y2=2.08
cc_1097 ( N_noxref_6_c_1248_n N_noxref_9_c_2030_n ) capacitor c=0.0198536f \
 //x=20.235 //y=3.33 //x2=12.95 //y2=2.08
cc_1098 ( N_noxref_6_c_1248_n N_noxref_9_c_2059_n ) capacitor c=0.0212788f \
 //x=20.235 //y=3.33 //x2=18.5 //y2=3.7
cc_1099 ( N_noxref_6_c_1251_n N_noxref_9_c_2059_n ) capacitor c=0.0121179f \
 //x=20.35 //y=2.08 //x2=18.5 //y2=3.7
cc_1100 ( N_noxref_6_c_1274_n N_noxref_9_M28_noxref_g ) capacitor c=0.01736f \
 //x=8.015 //y=5.155 //x2=7.88 //y2=6.02
cc_1101 ( N_noxref_6_M28_noxref_d N_noxref_9_M28_noxref_g ) capacitor \
 c=0.0180032f //x=7.955 //y=5.02 //x2=7.88 //y2=6.02
cc_1102 ( N_noxref_6_c_1278_n N_noxref_9_M29_noxref_g ) capacitor c=0.0194981f \
 //x=8.795 //y=5.155 //x2=8.32 //y2=6.02
cc_1103 ( N_noxref_6_M28_noxref_d N_noxref_9_M29_noxref_g ) capacitor \
 c=0.0194246f //x=7.955 //y=5.02 //x2=8.32 //y2=6.02
cc_1104 ( N_noxref_6_M5_noxref_d N_noxref_9_c_2151_n ) capacitor c=0.00217566f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=0.915
cc_1105 ( N_noxref_6_M5_noxref_d N_noxref_9_c_2152_n ) capacitor c=0.0034598f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=1.26
cc_1106 ( N_noxref_6_M5_noxref_d N_noxref_9_c_2153_n ) capacitor c=0.00546784f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=1.57
cc_1107 ( N_noxref_6_M5_noxref_d N_noxref_9_c_2191_n ) capacitor c=0.00241102f \
 //x=8.205 //y=0.915 //x2=8.505 //y2=0.76
cc_1108 ( N_noxref_6_c_1250_n N_noxref_9_c_2192_n ) capacitor c=0.00371277f \
 //x=8.795 //y=1.665 //x2=8.505 //y2=1.415
cc_1109 ( N_noxref_6_M5_noxref_d N_noxref_9_c_2192_n ) capacitor c=0.0138621f \
 //x=8.205 //y=0.915 //x2=8.505 //y2=1.415
cc_1110 ( N_noxref_6_M5_noxref_d N_noxref_9_c_2194_n ) capacitor c=0.00219619f \
 //x=8.205 //y=0.915 //x2=8.66 //y2=0.915
cc_1111 ( N_noxref_6_c_1250_n N_noxref_9_c_2195_n ) capacitor c=0.00457401f \
 //x=8.795 //y=1.665 //x2=8.66 //y2=1.26
cc_1112 ( N_noxref_6_M5_noxref_d N_noxref_9_c_2195_n ) capacitor c=0.00603828f \
 //x=8.205 //y=0.915 //x2=8.66 //y2=1.26
cc_1113 ( N_noxref_6_c_1282_n N_noxref_9_c_2154_n ) capacitor c=0.00731987f \
 //x=8.88 //y=3.33 //x2=8.14 //y2=2.08
cc_1114 ( N_noxref_6_c_1282_n N_noxref_9_c_2156_n ) capacitor c=0.00283672f \
 //x=8.88 //y=3.33 //x2=8.14 //y2=1.915
cc_1115 ( N_noxref_6_M5_noxref_d N_noxref_9_c_2156_n ) capacitor c=0.00661782f \
 //x=8.205 //y=0.915 //x2=8.14 //y2=1.915
cc_1116 ( N_noxref_6_c_1278_n N_noxref_9_c_2157_n ) capacitor c=0.00201851f \
 //x=8.795 //y=5.155 //x2=8.14 //y2=4.7
cc_1117 ( N_noxref_6_c_1282_n N_noxref_9_c_2157_n ) capacitor c=0.013693f \
 //x=8.88 //y=3.33 //x2=8.14 //y2=4.7
cc_1118 ( N_noxref_6_c_1454_p N_noxref_9_c_2157_n ) capacitor c=0.00475601f \
 //x=8.1 //y=5.155 //x2=8.14 //y2=4.7
cc_1119 ( N_noxref_6_c_1249_n N_noxref_10_c_2364_n ) capacitor c=0.00175234f \
 //x=3.33 //y=2.08 //x2=1.11 //y2=2.08
cc_1120 ( N_noxref_6_c_1249_n N_noxref_12_c_2473_n ) capacitor c=0.00204385f \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_1121 ( N_noxref_6_c_1340_n N_noxref_12_c_2473_n ) capacitor c=0.0194423f \
 //x=3.32 //y=0.915 //x2=3.985 //y2=0.54
cc_1122 ( N_noxref_6_c_1346_n N_noxref_12_c_2473_n ) capacitor c=0.00656458f \
 //x=3.85 //y=0.915 //x2=3.985 //y2=0.54
cc_1123 ( N_noxref_6_c_1349_n N_noxref_12_c_2473_n ) capacitor c=2.20712e-19 \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_1124 ( N_noxref_6_c_1341_n N_noxref_12_c_2484_n ) capacitor c=0.00538829f \
 //x=3.32 //y=1.26 //x2=3.1 //y2=0.995
cc_1125 ( N_noxref_6_c_1340_n N_noxref_12_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=0.915 //x2=2.965 //y2=0.375
cc_1126 ( N_noxref_6_c_1342_n N_noxref_12_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=1.57 //x2=2.965 //y2=0.375
cc_1127 ( N_noxref_6_c_1346_n N_noxref_12_M2_noxref_s ) capacitor c=0.0143002f \
 //x=3.85 //y=0.915 //x2=2.965 //y2=0.375
cc_1128 ( N_noxref_6_c_1347_n N_noxref_12_M2_noxref_s ) capacitor \
 c=0.00290153f //x=3.85 //y=1.26 //x2=2.965 //y2=0.375
cc_1129 ( N_noxref_6_M5_noxref_d N_noxref_13_M3_noxref_s ) capacitor \
 c=0.00309936f //x=8.205 //y=0.915 //x2=5.265 //y2=0.375
cc_1130 ( N_noxref_6_c_1250_n N_noxref_14_c_2577_n ) capacitor c=0.00457167f \
 //x=8.795 //y=1.665 //x2=8.795 //y2=0.54
cc_1131 ( N_noxref_6_M5_noxref_d N_noxref_14_c_2577_n ) capacitor c=0.0115903f \
 //x=8.205 //y=0.915 //x2=8.795 //y2=0.54
cc_1132 ( N_noxref_6_c_1384_p N_noxref_14_c_2600_n ) capacitor c=0.0200405f \
 //x=8.48 //y=1.665 //x2=7.91 //y2=0.995
cc_1133 ( N_noxref_6_M5_noxref_d N_noxref_14_M4_noxref_d ) capacitor \
 c=5.27807e-19 //x=8.205 //y=0.915 //x2=6.67 //y2=0.91
cc_1134 ( N_noxref_6_c_1250_n N_noxref_14_M5_noxref_s ) capacitor c=0.0196084f \
 //x=8.795 //y=1.665 //x2=7.775 //y2=0.375
cc_1135 ( N_noxref_6_M5_noxref_d N_noxref_14_M5_noxref_s ) capacitor \
 c=0.0426368f //x=8.205 //y=0.915 //x2=7.775 //y2=0.375
cc_1136 ( N_noxref_6_c_1250_n N_noxref_15_c_2641_n ) capacitor c=3.84569e-19 \
 //x=8.795 //y=1.665 //x2=10.21 //y2=1.505
cc_1137 ( N_noxref_6_M5_noxref_d N_noxref_15_M6_noxref_s ) capacitor \
 c=2.55333e-19 //x=8.205 //y=0.915 //x2=10.075 //y2=0.375
cc_1138 ( N_noxref_6_c_1256_n N_noxref_19_c_2850_n ) capacitor c=0.0034165f \
 //x=20.05 //y=1.915 //x2=19.83 //y2=1.505
cc_1139 ( N_noxref_6_c_1251_n N_noxref_19_c_2834_n ) capacitor c=0.0119952f \
 //x=20.35 //y=2.08 //x2=20.715 //y2=1.59
cc_1140 ( N_noxref_6_c_1255_n N_noxref_19_c_2834_n ) capacitor c=0.00697148f \
 //x=20.05 //y=1.53 //x2=20.715 //y2=1.59
cc_1141 ( N_noxref_6_c_1256_n N_noxref_19_c_2834_n ) capacitor c=0.0204849f \
 //x=20.05 //y=1.915 //x2=20.715 //y2=1.59
cc_1142 ( N_noxref_6_c_1258_n N_noxref_19_c_2834_n ) capacitor c=0.00610316f \
 //x=20.425 //y=1.375 //x2=20.715 //y2=1.59
cc_1143 ( N_noxref_6_c_1261_n N_noxref_19_c_2834_n ) capacitor c=0.00698822f \
 //x=20.58 //y=1.22 //x2=20.715 //y2=1.59
cc_1144 ( N_noxref_6_c_1252_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.0327271f //x=20.05 //y=0.875 //x2=19.695 //y2=0.375
cc_1145 ( N_noxref_6_c_1255_n N_noxref_19_M12_noxref_s ) capacitor \
 c=7.99997e-19 //x=20.05 //y=1.53 //x2=19.695 //y2=0.375
cc_1146 ( N_noxref_6_c_1256_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00122123f //x=20.05 //y=1.915 //x2=19.695 //y2=0.375
cc_1147 ( N_noxref_6_c_1259_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.0121427f //x=20.58 //y=0.875 //x2=19.695 //y2=0.375
cc_1148 ( N_noxref_6_c_1251_n N_noxref_20_c_2886_n ) capacitor c=0.00135272f \
 //x=20.35 //y=2.08 //x2=22.57 //y2=2.08
cc_1149 ( N_noxref_6_M43_noxref_g N_noxref_21_c_2947_n ) capacitor \
 c=0.0186539f //x=20.99 //y=6.02 //x2=21.565 //y2=5.155
cc_1150 ( N_noxref_6_M42_noxref_g N_noxref_21_c_2951_n ) capacitor \
 c=0.0213876f //x=20.55 //y=6.02 //x2=20.855 //y2=5.155
cc_1151 ( N_noxref_6_c_1403_p N_noxref_21_c_2951_n ) capacitor c=0.0044314f \
 //x=20.915 //y=4.79 //x2=20.855 //y2=5.155
cc_1152 ( N_noxref_6_M43_noxref_g N_noxref_21_M42_noxref_d ) capacitor \
 c=0.0180032f //x=20.99 //y=6.02 //x2=20.625 //y2=5.02
cc_1153 ( N_noxref_7_c_1511_n N_noxref_8_c_1827_n ) capacitor c=0.16065f \
 //x=17.645 //y=2.22 //x2=26.155 //y2=2.96
cc_1154 ( N_noxref_7_c_1523_n N_noxref_8_c_1827_n ) capacitor c=0.16049f \
 //x=21.345 //y=2.22 //x2=26.155 //y2=2.96
cc_1155 ( N_noxref_7_c_1527_n N_noxref_8_c_1827_n ) capacitor c=0.0120222f \
 //x=17.875 //y=2.22 //x2=26.155 //y2=2.96
cc_1156 ( N_noxref_7_c_1529_n N_noxref_8_c_1827_n ) capacitor c=0.0206071f \
 //x=17.76 //y=2.08 //x2=26.155 //y2=2.96
cc_1157 ( N_noxref_7_c_1530_n N_noxref_8_c_1827_n ) capacitor c=0.0239871f \
 //x=21.46 //y=2.08 //x2=26.155 //y2=2.96
cc_1158 ( N_noxref_7_c_1644_n N_noxref_8_c_1827_n ) capacitor c=4.10467e-19 \
 //x=21.55 //y=1.915 //x2=26.155 //y2=2.96
cc_1159 ( N_noxref_7_c_1511_n N_noxref_8_c_1847_n ) capacitor c=0.0132253f \
 //x=17.645 //y=2.22 //x2=11.955 //y2=2.96
cc_1160 ( N_noxref_7_c_1511_n N_noxref_8_c_1833_n ) capacitor c=0.0220464f \
 //x=17.645 //y=2.22 //x2=11.84 //y2=2.08
cc_1161 ( N_noxref_7_c_1511_n N_noxref_8_c_1864_n ) capacitor c=0.00583058f \
 //x=17.645 //y=2.22 //x2=11.93 //y2=1.915
cc_1162 ( N_noxref_7_c_1511_n N_noxref_9_c_2034_n ) capacitor c=0.00548028f \
 //x=17.645 //y=2.22 //x2=12.835 //y2=3.7
cc_1163 ( N_noxref_7_c_1529_n N_noxref_9_c_2035_n ) capacitor c=0.0227201f \
 //x=17.76 //y=2.08 //x2=18.385 //y2=3.7
cc_1164 ( N_noxref_7_c_1594_n N_noxref_9_c_2035_n ) capacitor c=0.00684517f \
 //x=17.76 //y=4.7 //x2=18.385 //y2=3.7
cc_1165 ( N_noxref_7_c_1523_n N_noxref_9_c_2028_n ) capacitor c=0.0044763f \
 //x=21.345 //y=2.22 //x2=27.265 //y2=3.7
cc_1166 ( N_noxref_7_c_1530_n N_noxref_9_c_2028_n ) capacitor c=0.026099f \
 //x=21.46 //y=2.08 //x2=27.265 //y2=3.7
cc_1167 ( N_noxref_7_c_1665_p N_noxref_9_c_2028_n ) capacitor c=0.00535612f \
 //x=21.795 //y=4.79 //x2=27.265 //y2=3.7
cc_1168 ( N_noxref_7_c_1648_n N_noxref_9_c_2028_n ) capacitor c=0.00138305f \
 //x=21.46 //y=4.7 //x2=27.265 //y2=3.7
cc_1169 ( N_noxref_7_c_1529_n N_noxref_9_c_2042_n ) capacitor c=0.00179385f \
 //x=17.76 //y=2.08 //x2=18.615 //y2=3.7
cc_1170 ( N_noxref_7_c_1511_n N_noxref_9_c_2029_n ) capacitor c=0.0186201f \
 //x=17.645 //y=2.22 //x2=8.14 //y2=2.08
cc_1171 ( N_noxref_7_c_1511_n N_noxref_9_c_2030_n ) capacitor c=0.0209607f \
 //x=17.645 //y=2.22 //x2=12.95 //y2=2.08
cc_1172 ( N_noxref_7_M40_noxref_g N_noxref_9_c_2051_n ) capacitor c=0.019179f \
 //x=17.5 //y=6.02 //x2=17.635 //y2=5.155
cc_1173 ( N_noxref_7_M41_noxref_g N_noxref_9_c_2055_n ) capacitor c=0.0213171f \
 //x=17.94 //y=6.02 //x2=18.415 //y2=5.155
cc_1174 ( N_noxref_7_c_1594_n N_noxref_9_c_2055_n ) capacitor c=0.00201851f \
 //x=17.76 //y=4.7 //x2=18.415 //y2=5.155
cc_1175 ( N_noxref_7_c_1673_p N_noxref_9_c_2031_n ) capacitor c=0.00371277f \
 //x=18.125 //y=1.415 //x2=18.415 //y2=1.665
cc_1176 ( N_noxref_7_c_1674_p N_noxref_9_c_2031_n ) capacitor c=0.00457401f \
 //x=18.28 //y=1.26 //x2=18.415 //y2=1.665
cc_1177 ( N_noxref_7_c_1523_n N_noxref_9_c_2218_n ) capacitor c=0.016327f \
 //x=21.345 //y=2.22 //x2=18.1 //y2=1.665
cc_1178 ( N_noxref_7_c_1523_n N_noxref_9_c_2059_n ) capacitor c=0.0220713f \
 //x=21.345 //y=2.22 //x2=18.5 //y2=3.7
cc_1179 ( N_noxref_7_c_1527_n N_noxref_9_c_2059_n ) capacitor c=0.0012045f \
 //x=17.875 //y=2.22 //x2=18.5 //y2=3.7
cc_1180 ( N_noxref_7_c_1529_n N_noxref_9_c_2059_n ) capacitor c=0.0822956f \
 //x=17.76 //y=2.08 //x2=18.5 //y2=3.7
cc_1181 ( N_noxref_7_c_1530_n N_noxref_9_c_2059_n ) capacitor c=6.4072e-19 \
 //x=21.46 //y=2.08 //x2=18.5 //y2=3.7
cc_1182 ( N_noxref_7_c_1591_n N_noxref_9_c_2059_n ) capacitor c=0.00709342f \
 //x=17.76 //y=2.08 //x2=18.5 //y2=3.7
cc_1183 ( N_noxref_7_c_1593_n N_noxref_9_c_2059_n ) capacitor c=0.00283672f \
 //x=17.76 //y=1.915 //x2=18.5 //y2=3.7
cc_1184 ( N_noxref_7_c_1594_n N_noxref_9_c_2059_n ) capacitor c=0.013693f \
 //x=17.76 //y=4.7 //x2=18.5 //y2=3.7
cc_1185 ( N_noxref_7_c_1529_n N_noxref_9_c_2226_n ) capacitor c=0.0177564f \
 //x=17.76 //y=2.08 //x2=17.72 //y2=5.155
cc_1186 ( N_noxref_7_c_1594_n N_noxref_9_c_2226_n ) capacitor c=0.00476349f \
 //x=17.76 //y=4.7 //x2=17.72 //y2=5.155
cc_1187 ( N_noxref_7_c_1511_n N_noxref_9_c_2192_n ) capacitor c=3.13485e-19 \
 //x=17.645 //y=2.22 //x2=8.505 //y2=1.415
cc_1188 ( N_noxref_7_c_1511_n N_noxref_9_c_2114_n ) capacitor c=3.13485e-19 \
 //x=17.645 //y=2.22 //x2=13.315 //y2=1.415
cc_1189 ( N_noxref_7_c_1511_n N_noxref_9_c_2154_n ) capacitor c=0.00584491f \
 //x=17.645 //y=2.22 //x2=8.14 //y2=2.08
cc_1190 ( N_noxref_7_c_1511_n N_noxref_9_c_2119_n ) capacitor c=0.00584491f \
 //x=17.645 //y=2.22 //x2=12.95 //y2=2.08
cc_1191 ( N_noxref_7_c_1588_n N_noxref_9_M11_noxref_d ) capacitor \
 c=0.00217566f //x=17.75 //y=0.915 //x2=17.825 //y2=0.915
cc_1192 ( N_noxref_7_c_1589_n N_noxref_9_M11_noxref_d ) capacitor c=0.0034598f \
 //x=17.75 //y=1.26 //x2=17.825 //y2=0.915
cc_1193 ( N_noxref_7_c_1590_n N_noxref_9_M11_noxref_d ) capacitor \
 c=0.00546784f //x=17.75 //y=1.57 //x2=17.825 //y2=0.915
cc_1194 ( N_noxref_7_c_1692_p N_noxref_9_M11_noxref_d ) capacitor \
 c=0.00241102f //x=18.125 //y=0.76 //x2=17.825 //y2=0.915
cc_1195 ( N_noxref_7_c_1673_p N_noxref_9_M11_noxref_d ) capacitor c=0.0138621f \
 //x=18.125 //y=1.415 //x2=17.825 //y2=0.915
cc_1196 ( N_noxref_7_c_1694_p N_noxref_9_M11_noxref_d ) capacitor \
 c=0.00219619f //x=18.28 //y=0.915 //x2=17.825 //y2=0.915
cc_1197 ( N_noxref_7_c_1674_p N_noxref_9_M11_noxref_d ) capacitor \
 c=0.00603828f //x=18.28 //y=1.26 //x2=17.825 //y2=0.915
cc_1198 ( N_noxref_7_c_1593_n N_noxref_9_M11_noxref_d ) capacitor \
 c=0.00661782f //x=17.76 //y=1.915 //x2=17.825 //y2=0.915
cc_1199 ( N_noxref_7_M40_noxref_g N_noxref_9_M40_noxref_d ) capacitor \
 c=0.0180032f //x=17.5 //y=6.02 //x2=17.575 //y2=5.02
cc_1200 ( N_noxref_7_M41_noxref_g N_noxref_9_M40_noxref_d ) capacitor \
 c=0.0194246f //x=17.94 //y=6.02 //x2=17.575 //y2=5.02
cc_1201 ( N_noxref_7_c_1522_n N_noxref_10_c_2364_n ) capacitor c=0.00558344f \
 //x=2.335 //y=2.22 //x2=1.11 //y2=2.08
cc_1202 ( N_noxref_7_c_1528_n N_noxref_10_c_2364_n ) capacitor c=0.0564721f \
 //x=2.22 //y=2.08 //x2=1.11 //y2=2.08
cc_1203 ( N_noxref_7_c_1632_n N_noxref_10_c_2364_n ) capacitor c=0.00211714f \
 //x=2.31 //y=1.915 //x2=1.11 //y2=2.08
cc_1204 ( N_noxref_7_c_1567_n N_noxref_10_c_2364_n ) capacitor c=0.00183762f \
 //x=2.22 //y=4.7 //x2=1.11 //y2=2.08
cc_1205 ( N_noxref_7_M20_noxref_g N_noxref_10_M18_noxref_g ) capacitor \
 c=0.0105869f //x=2.19 //y=6.02 //x2=1.31 //y2=6.02
cc_1206 ( N_noxref_7_M20_noxref_g N_noxref_10_M19_noxref_g ) capacitor \
 c=0.10632f //x=2.19 //y=6.02 //x2=1.75 //y2=6.02
cc_1207 ( N_noxref_7_M21_noxref_g N_noxref_10_M19_noxref_g ) capacitor \
 c=0.0101598f //x=2.63 //y=6.02 //x2=1.75 //y2=6.02
cc_1208 ( N_noxref_7_c_1706_p N_noxref_10_c_2365_n ) capacitor c=5.72482e-19 \
 //x=1.785 //y=0.91 //x2=0.81 //y2=0.875
cc_1209 ( N_noxref_7_c_1706_p N_noxref_10_c_2367_n ) capacitor c=0.00149976f \
 //x=1.785 //y=0.91 //x2=0.81 //y2=1.22
cc_1210 ( N_noxref_7_c_1708_p N_noxref_10_c_2368_n ) capacitor c=0.00111227f \
 //x=1.785 //y=1.22 //x2=0.81 //y2=1.53
cc_1211 ( N_noxref_7_c_1522_n N_noxref_10_c_2369_n ) capacitor c=0.00341397f \
 //x=2.335 //y=2.22 //x2=0.81 //y2=1.915
cc_1212 ( N_noxref_7_c_1528_n N_noxref_10_c_2369_n ) capacitor c=0.00228225f \
 //x=2.22 //y=2.08 //x2=0.81 //y2=1.915
cc_1213 ( N_noxref_7_c_1632_n N_noxref_10_c_2369_n ) capacitor c=0.00909574f \
 //x=2.31 //y=1.915 //x2=0.81 //y2=1.915
cc_1214 ( N_noxref_7_c_1706_p N_noxref_10_c_2372_n ) capacitor c=0.0160123f \
 //x=1.785 //y=0.91 //x2=1.34 //y2=0.875
cc_1215 ( N_noxref_7_c_1629_n N_noxref_10_c_2372_n ) capacitor c=0.00103227f \
 //x=2.31 //y=0.91 //x2=1.34 //y2=0.875
cc_1216 ( N_noxref_7_c_1708_p N_noxref_10_c_2374_n ) capacitor c=0.0124075f \
 //x=1.785 //y=1.22 //x2=1.34 //y2=1.22
cc_1217 ( N_noxref_7_c_1630_n N_noxref_10_c_2374_n ) capacitor c=0.0010154f \
 //x=2.31 //y=1.22 //x2=1.34 //y2=1.22
cc_1218 ( N_noxref_7_c_1631_n N_noxref_10_c_2374_n ) capacitor c=9.23422e-19 \
 //x=2.31 //y=1.45 //x2=1.34 //y2=1.22
cc_1219 ( N_noxref_7_c_1528_n N_noxref_10_c_2387_n ) capacitor c=0.00147352f \
 //x=2.22 //y=2.08 //x2=1.675 //y2=4.79
cc_1220 ( N_noxref_7_c_1567_n N_noxref_10_c_2387_n ) capacitor c=0.0168581f \
 //x=2.22 //y=4.7 //x2=1.675 //y2=4.79
cc_1221 ( N_noxref_7_c_1528_n N_noxref_10_c_2382_n ) capacitor c=0.00142741f \
 //x=2.22 //y=2.08 //x2=1.385 //y2=4.79
cc_1222 ( N_noxref_7_c_1567_n N_noxref_10_c_2382_n ) capacitor c=0.00484466f \
 //x=2.22 //y=4.7 //x2=1.385 //y2=4.79
cc_1223 ( N_noxref_7_c_1706_p N_noxref_11_c_2428_n ) capacitor c=0.0167228f \
 //x=1.785 //y=0.91 //x2=2.445 //y2=0.54
cc_1224 ( N_noxref_7_c_1629_n N_noxref_11_c_2428_n ) capacitor c=0.00534519f \
 //x=2.31 //y=0.91 //x2=2.445 //y2=0.54
cc_1225 ( N_noxref_7_c_1511_n N_noxref_11_c_2440_n ) capacitor c=0.00380711f \
 //x=17.645 //y=2.22 //x2=2.445 //y2=1.59
cc_1226 ( N_noxref_7_c_1522_n N_noxref_11_c_2440_n ) capacitor c=0.00354473f \
 //x=2.335 //y=2.22 //x2=2.445 //y2=1.59
cc_1227 ( N_noxref_7_c_1528_n N_noxref_11_c_2440_n ) capacitor c=0.011736f \
 //x=2.22 //y=2.08 //x2=2.445 //y2=1.59
cc_1228 ( N_noxref_7_c_1708_p N_noxref_11_c_2440_n ) capacitor c=0.0153695f \
 //x=1.785 //y=1.22 //x2=2.445 //y2=1.59
cc_1229 ( N_noxref_7_c_1632_n N_noxref_11_c_2440_n ) capacitor c=0.0213278f \
 //x=2.31 //y=1.915 //x2=2.445 //y2=1.59
cc_1230 ( N_noxref_7_c_1511_n N_noxref_11_M0_noxref_s ) capacitor c=0.0058288f \
 //x=17.645 //y=2.22 //x2=0.455 //y2=0.375
cc_1231 ( N_noxref_7_c_1706_p N_noxref_11_M0_noxref_s ) capacitor \
 c=0.00798959f //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_1232 ( N_noxref_7_c_1631_n N_noxref_11_M0_noxref_s ) capacitor \
 c=0.00212176f //x=2.31 //y=1.45 //x2=0.455 //y2=0.375
cc_1233 ( N_noxref_7_c_1632_n N_noxref_11_M0_noxref_s ) capacitor \
 c=0.00298115f //x=2.31 //y=1.915 //x2=0.455 //y2=0.375
cc_1234 ( N_noxref_7_c_1511_n N_noxref_12_c_2467_n ) capacitor c=0.00608834f \
 //x=17.645 //y=2.22 //x2=3.015 //y2=0.995
cc_1235 ( N_noxref_7_c_1733_p N_noxref_12_c_2467_n ) capacitor c=2.14837e-19 \
 //x=2.155 //y=0.755 //x2=3.015 //y2=0.995
cc_1236 ( N_noxref_7_c_1629_n N_noxref_12_c_2467_n ) capacitor c=0.00123426f \
 //x=2.31 //y=0.91 //x2=3.015 //y2=0.995
cc_1237 ( N_noxref_7_c_1630_n N_noxref_12_c_2467_n ) capacitor c=0.0129288f \
 //x=2.31 //y=1.22 //x2=3.015 //y2=0.995
cc_1238 ( N_noxref_7_c_1631_n N_noxref_12_c_2467_n ) capacitor c=0.00142359f \
 //x=2.31 //y=1.45 //x2=3.015 //y2=0.995
cc_1239 ( N_noxref_7_c_1511_n N_noxref_12_c_2473_n ) capacitor c=0.00147946f \
 //x=17.645 //y=2.22 //x2=3.985 //y2=0.54
cc_1240 ( N_noxref_7_c_1706_p N_noxref_12_M1_noxref_d ) capacitor \
 c=0.00223875f //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_1241 ( N_noxref_7_c_1708_p N_noxref_12_M1_noxref_d ) capacitor \
 c=0.00262485f //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_1242 ( N_noxref_7_c_1733_p N_noxref_12_M1_noxref_d ) capacitor \
 c=0.00220746f //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_1243 ( N_noxref_7_c_1741_p N_noxref_12_M1_noxref_d ) capacitor \
 c=0.00194798f //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_1244 ( N_noxref_7_c_1629_n N_noxref_12_M1_noxref_d ) capacitor \
 c=0.00198465f //x=2.31 //y=0.91 //x2=1.86 //y2=0.91
cc_1245 ( N_noxref_7_c_1630_n N_noxref_12_M1_noxref_d ) capacitor \
 c=0.00128384f //x=2.31 //y=1.22 //x2=1.86 //y2=0.91
cc_1246 ( N_noxref_7_c_1511_n N_noxref_12_M2_noxref_s ) capacitor \
 c=0.00631802f //x=17.645 //y=2.22 //x2=2.965 //y2=0.375
cc_1247 ( N_noxref_7_c_1629_n N_noxref_12_M2_noxref_s ) capacitor \
 c=7.21316e-19 //x=2.31 //y=0.91 //x2=2.965 //y2=0.375
cc_1248 ( N_noxref_7_c_1630_n N_noxref_12_M2_noxref_s ) capacitor \
 c=0.00348171f //x=2.31 //y=1.22 //x2=2.965 //y2=0.375
cc_1249 ( N_noxref_7_c_1511_n N_noxref_13_c_2537_n ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=5.4 //y2=1.505
cc_1250 ( N_noxref_7_c_1511_n N_noxref_13_c_2521_n ) capacitor c=0.0225733f \
 //x=17.645 //y=2.22 //x2=6.285 //y2=1.59
cc_1251 ( N_noxref_7_c_1511_n N_noxref_13_c_2551_n ) capacitor c=0.0203655f \
 //x=17.645 //y=2.22 //x2=7.255 //y2=1.59
cc_1252 ( N_noxref_7_c_1511_n N_noxref_13_M3_noxref_s ) capacitor c=0.012425f \
 //x=17.645 //y=2.22 //x2=5.265 //y2=0.375
cc_1253 ( N_noxref_7_c_1511_n N_noxref_14_c_2571_n ) capacitor c=0.00657782f \
 //x=17.645 //y=2.22 //x2=7.825 //y2=0.995
cc_1254 ( N_noxref_7_c_1511_n N_noxref_14_c_2577_n ) capacitor c=0.00147946f \
 //x=17.645 //y=2.22 //x2=8.795 //y2=0.54
cc_1255 ( N_noxref_7_c_1511_n N_noxref_14_M5_noxref_s ) capacitor \
 c=0.00642985f //x=17.645 //y=2.22 //x2=7.775 //y2=0.375
cc_1256 ( N_noxref_7_c_1511_n N_noxref_15_c_2641_n ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=10.21 //y2=1.505
cc_1257 ( N_noxref_7_c_1511_n N_noxref_15_c_2625_n ) capacitor c=0.0225733f \
 //x=17.645 //y=2.22 //x2=11.095 //y2=1.59
cc_1258 ( N_noxref_7_c_1511_n N_noxref_15_c_2656_n ) capacitor c=0.0203655f \
 //x=17.645 //y=2.22 //x2=12.065 //y2=1.59
cc_1259 ( N_noxref_7_c_1511_n N_noxref_15_M6_noxref_s ) capacitor c=0.012425f \
 //x=17.645 //y=2.22 //x2=10.075 //y2=0.375
cc_1260 ( N_noxref_7_c_1511_n N_noxref_16_c_2675_n ) capacitor c=0.00657782f \
 //x=17.645 //y=2.22 //x2=12.635 //y2=0.995
cc_1261 ( N_noxref_7_c_1511_n N_noxref_16_c_2681_n ) capacitor c=0.00147946f \
 //x=17.645 //y=2.22 //x2=13.605 //y2=0.54
cc_1262 ( N_noxref_7_c_1511_n N_noxref_16_M8_noxref_s ) capacitor \
 c=0.00642985f //x=17.645 //y=2.22 //x2=12.585 //y2=0.375
cc_1263 ( N_noxref_7_c_1511_n N_noxref_17_c_2745_n ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=15.02 //y2=1.505
cc_1264 ( N_noxref_7_c_1511_n N_noxref_17_c_2729_n ) capacitor c=0.0225733f \
 //x=17.645 //y=2.22 //x2=15.905 //y2=1.59
cc_1265 ( N_noxref_7_c_1511_n N_noxref_17_c_2759_n ) capacitor c=0.0203655f \
 //x=17.645 //y=2.22 //x2=16.875 //y2=1.59
cc_1266 ( N_noxref_7_c_1511_n N_noxref_17_M9_noxref_s ) capacitor c=0.012425f \
 //x=17.645 //y=2.22 //x2=14.885 //y2=0.375
cc_1267 ( N_noxref_7_c_1511_n N_noxref_18_c_2779_n ) capacitor c=0.00657782f \
 //x=17.645 //y=2.22 //x2=17.445 //y2=0.995
cc_1268 ( N_noxref_7_c_1523_n N_noxref_18_c_2785_n ) capacitor c=7.41833e-19 \
 //x=21.345 //y=2.22 //x2=18.415 //y2=0.54
cc_1269 ( N_noxref_7_c_1527_n N_noxref_18_c_2785_n ) capacitor c=7.4531e-19 \
 //x=17.875 //y=2.22 //x2=18.415 //y2=0.54
cc_1270 ( N_noxref_7_c_1529_n N_noxref_18_c_2785_n ) capacitor c=0.00204178f \
 //x=17.76 //y=2.08 //x2=18.415 //y2=0.54
cc_1271 ( N_noxref_7_c_1588_n N_noxref_18_c_2785_n ) capacitor c=0.0194423f \
 //x=17.75 //y=0.915 //x2=18.415 //y2=0.54
cc_1272 ( N_noxref_7_c_1694_p N_noxref_18_c_2785_n ) capacitor c=0.00656458f \
 //x=18.28 //y=0.915 //x2=18.415 //y2=0.54
cc_1273 ( N_noxref_7_c_1591_n N_noxref_18_c_2785_n ) capacitor c=2.20712e-19 \
 //x=17.76 //y=2.08 //x2=18.415 //y2=0.54
cc_1274 ( N_noxref_7_c_1589_n N_noxref_18_c_2813_n ) capacitor c=0.00538829f \
 //x=17.75 //y=1.26 //x2=17.53 //y2=0.995
cc_1275 ( N_noxref_7_c_1511_n N_noxref_18_M11_noxref_s ) capacitor \
 c=0.00642985f //x=17.645 //y=2.22 //x2=17.395 //y2=0.375
cc_1276 ( N_noxref_7_c_1588_n N_noxref_18_M11_noxref_s ) capacitor \
 c=0.00538829f //x=17.75 //y=0.915 //x2=17.395 //y2=0.375
cc_1277 ( N_noxref_7_c_1590_n N_noxref_18_M11_noxref_s ) capacitor \
 c=0.00538829f //x=17.75 //y=1.57 //x2=17.395 //y2=0.375
cc_1278 ( N_noxref_7_c_1694_p N_noxref_18_M11_noxref_s ) capacitor \
 c=0.0143002f //x=18.28 //y=0.915 //x2=17.395 //y2=0.375
cc_1279 ( N_noxref_7_c_1674_p N_noxref_18_M11_noxref_s ) capacitor \
 c=0.00290153f //x=18.28 //y=1.26 //x2=17.395 //y2=0.375
cc_1280 ( N_noxref_7_c_1523_n N_noxref_19_c_2850_n ) capacitor c=0.00642985f \
 //x=21.345 //y=2.22 //x2=19.83 //y2=1.505
cc_1281 ( N_noxref_7_c_1523_n N_noxref_19_c_2834_n ) capacitor c=0.0225733f \
 //x=21.345 //y=2.22 //x2=20.715 //y2=1.59
cc_1282 ( N_noxref_7_c_1636_n N_noxref_19_c_2841_n ) capacitor c=0.0167228f \
 //x=21.025 //y=0.91 //x2=21.685 //y2=0.54
cc_1283 ( N_noxref_7_c_1641_n N_noxref_19_c_2841_n ) capacitor c=0.00534519f \
 //x=21.55 //y=0.91 //x2=21.685 //y2=0.54
cc_1284 ( N_noxref_7_c_1523_n N_noxref_19_c_2864_n ) capacitor c=0.0178105f \
 //x=21.345 //y=2.22 //x2=21.685 //y2=1.59
cc_1285 ( N_noxref_7_c_1530_n N_noxref_19_c_2864_n ) capacitor c=0.0119919f \
 //x=21.46 //y=2.08 //x2=21.685 //y2=1.59
cc_1286 ( N_noxref_7_c_1639_n N_noxref_19_c_2864_n ) capacitor c=0.0157358f \
 //x=21.025 //y=1.22 //x2=21.685 //y2=1.59
cc_1287 ( N_noxref_7_c_1644_n N_noxref_19_c_2864_n ) capacitor c=0.0215856f \
 //x=21.55 //y=1.915 //x2=21.685 //y2=1.59
cc_1288 ( N_noxref_7_c_1523_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00642985f //x=21.345 //y=2.22 //x2=19.695 //y2=0.375
cc_1289 ( N_noxref_7_c_1636_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00798959f //x=21.025 //y=0.91 //x2=19.695 //y2=0.375
cc_1290 ( N_noxref_7_c_1643_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00212176f //x=21.55 //y=1.45 //x2=19.695 //y2=0.375
cc_1291 ( N_noxref_7_c_1644_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00298115f //x=21.55 //y=1.915 //x2=19.695 //y2=0.375
cc_1292 ( N_noxref_7_c_1523_n N_noxref_20_c_2886_n ) capacitor c=0.00558344f \
 //x=21.345 //y=2.22 //x2=22.57 //y2=2.08
cc_1293 ( N_noxref_7_c_1530_n N_noxref_20_c_2886_n ) capacitor c=0.0517779f \
 //x=21.46 //y=2.08 //x2=22.57 //y2=2.08
cc_1294 ( N_noxref_7_c_1644_n N_noxref_20_c_2886_n ) capacitor c=0.00213841f \
 //x=21.55 //y=1.915 //x2=22.57 //y2=2.08
cc_1295 ( N_noxref_7_c_1648_n N_noxref_20_c_2886_n ) capacitor c=0.00142741f \
 //x=21.46 //y=4.7 //x2=22.57 //y2=2.08
cc_1296 ( N_noxref_7_M44_noxref_g N_noxref_20_M46_noxref_g ) capacitor \
 c=0.0101598f //x=21.43 //y=6.02 //x2=22.31 //y2=6.02
cc_1297 ( N_noxref_7_M45_noxref_g N_noxref_20_M46_noxref_g ) capacitor \
 c=0.0602553f //x=21.87 //y=6.02 //x2=22.31 //y2=6.02
cc_1298 ( N_noxref_7_M45_noxref_g N_noxref_20_M47_noxref_g ) capacitor \
 c=0.0101598f //x=21.87 //y=6.02 //x2=22.75 //y2=6.02
cc_1299 ( N_noxref_7_c_1641_n N_noxref_20_c_2900_n ) capacitor c=0.00456962f \
 //x=21.55 //y=0.91 //x2=22.56 //y2=0.915
cc_1300 ( N_noxref_7_c_1642_n N_noxref_20_c_2901_n ) capacitor c=0.00438372f \
 //x=21.55 //y=1.22 //x2=22.56 //y2=1.26
cc_1301 ( N_noxref_7_c_1643_n N_noxref_20_c_2902_n ) capacitor c=0.00438372f \
 //x=21.55 //y=1.45 //x2=22.56 //y2=1.57
cc_1302 ( N_noxref_7_c_1523_n N_noxref_20_c_2903_n ) capacitor c=0.00341397f \
 //x=21.345 //y=2.22 //x2=22.57 //y2=2.08
cc_1303 ( N_noxref_7_c_1530_n N_noxref_20_c_2903_n ) capacitor c=0.0021852f \
 //x=21.46 //y=2.08 //x2=22.57 //y2=2.08
cc_1304 ( N_noxref_7_c_1644_n N_noxref_20_c_2903_n ) capacitor c=0.00896806f \
 //x=21.55 //y=1.915 //x2=22.57 //y2=2.08
cc_1305 ( N_noxref_7_c_1644_n N_noxref_20_c_2906_n ) capacitor c=0.00438372f \
 //x=21.55 //y=1.915 //x2=22.57 //y2=1.915
cc_1306 ( N_noxref_7_c_1530_n N_noxref_20_c_2907_n ) capacitor c=0.00219458f \
 //x=21.46 //y=2.08 //x2=22.57 //y2=4.7
cc_1307 ( N_noxref_7_c_1665_p N_noxref_20_c_2907_n ) capacitor c=0.0611812f \
 //x=21.795 //y=4.79 //x2=22.57 //y2=4.7
cc_1308 ( N_noxref_7_c_1648_n N_noxref_20_c_2907_n ) capacitor c=0.00487508f \
 //x=21.46 //y=4.7 //x2=22.57 //y2=4.7
cc_1309 ( N_noxref_7_c_1530_n N_noxref_21_c_2947_n ) capacitor c=0.0149705f \
 //x=21.46 //y=2.08 //x2=21.565 //y2=5.155
cc_1310 ( N_noxref_7_M44_noxref_g N_noxref_21_c_2947_n ) capacitor \
 c=0.0167692f //x=21.43 //y=6.02 //x2=21.565 //y2=5.155
cc_1311 ( N_noxref_7_c_1648_n N_noxref_21_c_2947_n ) capacitor c=0.00325274f \
 //x=21.46 //y=4.7 //x2=21.565 //y2=5.155
cc_1312 ( N_noxref_7_M45_noxref_g N_noxref_21_c_2953_n ) capacitor c=0.019179f \
 //x=21.87 //y=6.02 //x2=22.445 //y2=5.155
cc_1313 ( N_noxref_7_c_1530_n N_noxref_21_c_2961_n ) capacitor c=0.00325304f \
 //x=21.46 //y=2.08 //x2=23.31 //y2=5.07
cc_1314 ( N_noxref_7_c_1665_p N_noxref_21_c_2986_n ) capacitor c=0.00441288f \
 //x=21.795 //y=4.79 //x2=21.65 //y2=5.155
cc_1315 ( N_noxref_7_M44_noxref_g N_noxref_21_M44_noxref_d ) capacitor \
 c=0.0180032f //x=21.43 //y=6.02 //x2=21.505 //y2=5.02
cc_1316 ( N_noxref_7_M45_noxref_g N_noxref_21_M44_noxref_d ) capacitor \
 c=0.0180032f //x=21.87 //y=6.02 //x2=21.505 //y2=5.02
cc_1317 ( N_noxref_7_c_1815_p N_noxref_22_c_3029_n ) capacitor c=2.14837e-19 \
 //x=21.395 //y=0.755 //x2=22.255 //y2=0.995
cc_1318 ( N_noxref_7_c_1641_n N_noxref_22_c_3029_n ) capacitor c=0.00123426f \
 //x=21.55 //y=0.91 //x2=22.255 //y2=0.995
cc_1319 ( N_noxref_7_c_1642_n N_noxref_22_c_3029_n ) capacitor c=0.0129288f \
 //x=21.55 //y=1.22 //x2=22.255 //y2=0.995
cc_1320 ( N_noxref_7_c_1643_n N_noxref_22_c_3029_n ) capacitor c=0.00142359f \
 //x=21.55 //y=1.45 //x2=22.255 //y2=0.995
cc_1321 ( N_noxref_7_c_1636_n N_noxref_22_M13_noxref_d ) capacitor \
 c=0.00223875f //x=21.025 //y=0.91 //x2=21.1 //y2=0.91
cc_1322 ( N_noxref_7_c_1639_n N_noxref_22_M13_noxref_d ) capacitor \
 c=0.00262485f //x=21.025 //y=1.22 //x2=21.1 //y2=0.91
cc_1323 ( N_noxref_7_c_1815_p N_noxref_22_M13_noxref_d ) capacitor \
 c=0.00220746f //x=21.395 //y=0.755 //x2=21.1 //y2=0.91
cc_1324 ( N_noxref_7_c_1822_p N_noxref_22_M13_noxref_d ) capacitor \
 c=0.00194798f //x=21.395 //y=1.375 //x2=21.1 //y2=0.91
cc_1325 ( N_noxref_7_c_1641_n N_noxref_22_M13_noxref_d ) capacitor \
 c=0.00198465f //x=21.55 //y=0.91 //x2=21.1 //y2=0.91
cc_1326 ( N_noxref_7_c_1642_n N_noxref_22_M13_noxref_d ) capacitor \
 c=0.00128384f //x=21.55 //y=1.22 //x2=21.1 //y2=0.91
cc_1327 ( N_noxref_7_c_1641_n N_noxref_22_M14_noxref_s ) capacitor \
 c=7.21316e-19 //x=21.55 //y=0.91 //x2=22.205 //y2=0.375
cc_1328 ( N_noxref_7_c_1642_n N_noxref_22_M14_noxref_s ) capacitor \
 c=0.00348171f //x=21.55 //y=1.22 //x2=22.205 //y2=0.375
cc_1329 ( N_noxref_8_c_1827_n N_noxref_9_c_2034_n ) capacitor c=0.0092394f \
 //x=26.155 //y=2.96 //x2=12.835 //y2=3.7
cc_1330 ( N_noxref_8_c_1847_n N_noxref_9_c_2034_n ) capacitor c=9.83937e-19 \
 //x=11.955 //y=2.96 //x2=12.835 //y2=3.7
cc_1331 ( N_noxref_8_c_1833_n N_noxref_9_c_2034_n ) capacitor c=0.0213449f \
 //x=11.84 //y=2.08 //x2=12.835 //y2=3.7
cc_1332 ( N_noxref_8_c_1827_n N_noxref_9_c_2035_n ) capacitor c=0.041794f \
 //x=26.155 //y=2.96 //x2=18.385 //y2=3.7
cc_1333 ( N_noxref_8_c_1827_n N_noxref_9_c_2097_n ) capacitor c=6.03896e-19 \
 //x=26.155 //y=2.96 //x2=13.065 //y2=3.7
cc_1334 ( N_noxref_8_c_1833_n N_noxref_9_c_2097_n ) capacitor c=0.00128547f \
 //x=11.84 //y=2.08 //x2=13.065 //y2=3.7
cc_1335 ( N_noxref_8_c_1827_n N_noxref_9_c_2028_n ) capacitor c=0.267326f \
 //x=26.155 //y=2.96 //x2=27.265 //y2=3.7
cc_1336 ( N_noxref_8_c_1834_n N_noxref_9_c_2028_n ) capacitor c=0.027702f \
 //x=26.27 //y=2.08 //x2=27.265 //y2=3.7
cc_1337 ( N_noxref_8_c_1907_p N_noxref_9_c_2028_n ) capacitor c=0.00535612f \
 //x=26.605 //y=4.79 //x2=27.265 //y2=3.7
cc_1338 ( N_noxref_8_c_1908_p N_noxref_9_c_2028_n ) capacitor c=0.00138305f \
 //x=26.27 //y=4.7 //x2=27.265 //y2=3.7
cc_1339 ( N_noxref_8_c_1827_n N_noxref_9_c_2042_n ) capacitor c=4.80612e-19 \
 //x=26.155 //y=2.96 //x2=18.615 //y2=3.7
cc_1340 ( N_noxref_8_c_1827_n N_noxref_9_c_2030_n ) capacitor c=0.0202855f \
 //x=26.155 //y=2.96 //x2=12.95 //y2=2.08
cc_1341 ( N_noxref_8_c_1847_n N_noxref_9_c_2030_n ) capacitor c=0.00128547f \
 //x=11.955 //y=2.96 //x2=12.95 //y2=2.08
cc_1342 ( N_noxref_8_c_1833_n N_noxref_9_c_2030_n ) capacitor c=0.0456719f \
 //x=11.84 //y=2.08 //x2=12.95 //y2=2.08
cc_1343 ( N_noxref_8_c_1864_n N_noxref_9_c_2030_n ) capacitor c=0.00205895f \
 //x=11.93 //y=1.915 //x2=12.95 //y2=2.08
cc_1344 ( N_noxref_8_c_1866_n N_noxref_9_c_2030_n ) capacitor c=0.00142741f \
 //x=11.84 //y=4.7 //x2=12.95 //y2=2.08
cc_1345 ( N_noxref_8_c_1827_n N_noxref_9_c_2059_n ) capacitor c=0.0210712f \
 //x=26.155 //y=2.96 //x2=18.5 //y2=3.7
cc_1346 ( N_noxref_8_c_1827_n N_noxref_9_c_2032_n ) capacitor c=0.00526349f \
 //x=26.155 //y=2.96 //x2=27.38 //y2=2.08
cc_1347 ( N_noxref_8_c_1834_n N_noxref_9_c_2032_n ) capacitor c=0.0538804f \
 //x=26.27 //y=2.08 //x2=27.38 //y2=2.08
cc_1348 ( N_noxref_8_c_1918_p N_noxref_9_c_2032_n ) capacitor c=0.0023343f \
 //x=26.36 //y=1.915 //x2=27.38 //y2=2.08
cc_1349 ( N_noxref_8_c_1908_p N_noxref_9_c_2032_n ) capacitor c=0.00142741f \
 //x=26.27 //y=4.7 //x2=27.38 //y2=2.08
cc_1350 ( N_noxref_8_M32_noxref_g N_noxref_9_M34_noxref_g ) capacitor \
 c=0.0101598f //x=11.81 //y=6.02 //x2=12.69 //y2=6.02
cc_1351 ( N_noxref_8_M33_noxref_g N_noxref_9_M34_noxref_g ) capacitor \
 c=0.0602553f //x=12.25 //y=6.02 //x2=12.69 //y2=6.02
cc_1352 ( N_noxref_8_M33_noxref_g N_noxref_9_M35_noxref_g ) capacitor \
 c=0.0101598f //x=12.25 //y=6.02 //x2=13.13 //y2=6.02
cc_1353 ( N_noxref_8_M50_noxref_g N_noxref_9_M52_noxref_g ) capacitor \
 c=0.0101598f //x=26.24 //y=6.02 //x2=27.12 //y2=6.02
cc_1354 ( N_noxref_8_M51_noxref_g N_noxref_9_M52_noxref_g ) capacitor \
 c=0.0602553f //x=26.68 //y=6.02 //x2=27.12 //y2=6.02
cc_1355 ( N_noxref_8_M51_noxref_g N_noxref_9_M53_noxref_g ) capacitor \
 c=0.0101598f //x=26.68 //y=6.02 //x2=27.56 //y2=6.02
cc_1356 ( N_noxref_8_c_1861_n N_noxref_9_c_2110_n ) capacitor c=0.00456962f \
 //x=11.93 //y=0.91 //x2=12.94 //y2=0.915
cc_1357 ( N_noxref_8_c_1862_n N_noxref_9_c_2111_n ) capacitor c=0.00438372f \
 //x=11.93 //y=1.22 //x2=12.94 //y2=1.26
cc_1358 ( N_noxref_8_c_1863_n N_noxref_9_c_2112_n ) capacitor c=0.00438372f \
 //x=11.93 //y=1.45 //x2=12.94 //y2=1.57
cc_1359 ( N_noxref_8_c_1929_p N_noxref_9_c_2272_n ) capacitor c=0.00456962f \
 //x=26.36 //y=0.91 //x2=27.37 //y2=0.915
cc_1360 ( N_noxref_8_c_1930_p N_noxref_9_c_2273_n ) capacitor c=0.00438372f \
 //x=26.36 //y=1.22 //x2=27.37 //y2=1.26
cc_1361 ( N_noxref_8_c_1931_p N_noxref_9_c_2274_n ) capacitor c=0.00438372f \
 //x=26.36 //y=1.45 //x2=27.37 //y2=1.57
cc_1362 ( N_noxref_8_c_1833_n N_noxref_9_c_2119_n ) capacitor c=0.00201097f \
 //x=11.84 //y=2.08 //x2=12.95 //y2=2.08
cc_1363 ( N_noxref_8_c_1864_n N_noxref_9_c_2119_n ) capacitor c=0.00828003f \
 //x=11.93 //y=1.915 //x2=12.95 //y2=2.08
cc_1364 ( N_noxref_8_c_1864_n N_noxref_9_c_2120_n ) capacitor c=0.00438372f \
 //x=11.93 //y=1.915 //x2=12.95 //y2=1.915
cc_1365 ( N_noxref_8_c_1833_n N_noxref_9_c_2122_n ) capacitor c=0.00219458f \
 //x=11.84 //y=2.08 //x2=12.95 //y2=4.7
cc_1366 ( N_noxref_8_c_1879_n N_noxref_9_c_2122_n ) capacitor c=0.0611812f \
 //x=12.175 //y=4.79 //x2=12.95 //y2=4.7
cc_1367 ( N_noxref_8_c_1866_n N_noxref_9_c_2122_n ) capacitor c=0.00487508f \
 //x=11.84 //y=4.7 //x2=12.95 //y2=4.7
cc_1368 ( N_noxref_8_c_1834_n N_noxref_9_c_2281_n ) capacitor c=0.00228632f \
 //x=26.27 //y=2.08 //x2=27.38 //y2=2.08
cc_1369 ( N_noxref_8_c_1918_p N_noxref_9_c_2281_n ) capacitor c=0.00933826f \
 //x=26.36 //y=1.915 //x2=27.38 //y2=2.08
cc_1370 ( N_noxref_8_c_1918_p N_noxref_9_c_2283_n ) capacitor c=0.00438372f \
 //x=26.36 //y=1.915 //x2=27.38 //y2=1.915
cc_1371 ( N_noxref_8_c_1834_n N_noxref_9_c_2284_n ) capacitor c=0.00219458f \
 //x=26.27 //y=2.08 //x2=27.38 //y2=4.7
cc_1372 ( N_noxref_8_c_1907_p N_noxref_9_c_2284_n ) capacitor c=0.0611812f \
 //x=26.605 //y=4.79 //x2=27.38 //y2=4.7
cc_1373 ( N_noxref_8_c_1908_p N_noxref_9_c_2284_n ) capacitor c=0.00487508f \
 //x=26.27 //y=4.7 //x2=27.38 //y2=4.7
cc_1374 ( N_noxref_8_c_1856_n N_noxref_15_c_2632_n ) capacitor c=0.0167228f \
 //x=11.405 //y=0.91 //x2=12.065 //y2=0.54
cc_1375 ( N_noxref_8_c_1861_n N_noxref_15_c_2632_n ) capacitor c=0.00534519f \
 //x=11.93 //y=0.91 //x2=12.065 //y2=0.54
cc_1376 ( N_noxref_8_c_1833_n N_noxref_15_c_2656_n ) capacitor c=0.0117694f \
 //x=11.84 //y=2.08 //x2=12.065 //y2=1.59
cc_1377 ( N_noxref_8_c_1859_n N_noxref_15_c_2656_n ) capacitor c=0.0157358f \
 //x=11.405 //y=1.22 //x2=12.065 //y2=1.59
cc_1378 ( N_noxref_8_c_1864_n N_noxref_15_c_2656_n ) capacitor c=0.021347f \
 //x=11.93 //y=1.915 //x2=12.065 //y2=1.59
cc_1379 ( N_noxref_8_c_1856_n N_noxref_15_M6_noxref_s ) capacitor \
 c=0.00798959f //x=11.405 //y=0.91 //x2=10.075 //y2=0.375
cc_1380 ( N_noxref_8_c_1863_n N_noxref_15_M6_noxref_s ) capacitor \
 c=0.00212176f //x=11.93 //y=1.45 //x2=10.075 //y2=0.375
cc_1381 ( N_noxref_8_c_1864_n N_noxref_15_M6_noxref_s ) capacitor \
 c=0.00298115f //x=11.93 //y=1.915 //x2=10.075 //y2=0.375
cc_1382 ( N_noxref_8_c_1952_p N_noxref_16_c_2675_n ) capacitor c=2.14837e-19 \
 //x=11.775 //y=0.755 //x2=12.635 //y2=0.995
cc_1383 ( N_noxref_8_c_1861_n N_noxref_16_c_2675_n ) capacitor c=0.00123426f \
 //x=11.93 //y=0.91 //x2=12.635 //y2=0.995
cc_1384 ( N_noxref_8_c_1862_n N_noxref_16_c_2675_n ) capacitor c=0.0129288f \
 //x=11.93 //y=1.22 //x2=12.635 //y2=0.995
cc_1385 ( N_noxref_8_c_1863_n N_noxref_16_c_2675_n ) capacitor c=0.00142359f \
 //x=11.93 //y=1.45 //x2=12.635 //y2=0.995
cc_1386 ( N_noxref_8_c_1856_n N_noxref_16_M7_noxref_d ) capacitor \
 c=0.00223875f //x=11.405 //y=0.91 //x2=11.48 //y2=0.91
cc_1387 ( N_noxref_8_c_1859_n N_noxref_16_M7_noxref_d ) capacitor \
 c=0.00262485f //x=11.405 //y=1.22 //x2=11.48 //y2=0.91
cc_1388 ( N_noxref_8_c_1952_p N_noxref_16_M7_noxref_d ) capacitor \
 c=0.00220746f //x=11.775 //y=0.755 //x2=11.48 //y2=0.91
cc_1389 ( N_noxref_8_c_1959_p N_noxref_16_M7_noxref_d ) capacitor \
 c=0.00194798f //x=11.775 //y=1.375 //x2=11.48 //y2=0.91
cc_1390 ( N_noxref_8_c_1861_n N_noxref_16_M7_noxref_d ) capacitor \
 c=0.00198465f //x=11.93 //y=0.91 //x2=11.48 //y2=0.91
cc_1391 ( N_noxref_8_c_1862_n N_noxref_16_M7_noxref_d ) capacitor \
 c=0.00128384f //x=11.93 //y=1.22 //x2=11.48 //y2=0.91
cc_1392 ( N_noxref_8_c_1861_n N_noxref_16_M8_noxref_s ) capacitor \
 c=7.21316e-19 //x=11.93 //y=0.91 //x2=12.585 //y2=0.375
cc_1393 ( N_noxref_8_c_1862_n N_noxref_16_M8_noxref_s ) capacitor \
 c=0.00348171f //x=11.93 //y=1.22 //x2=12.585 //y2=0.375
cc_1394 ( N_noxref_8_c_1827_n N_noxref_19_c_2864_n ) capacitor c=0.00152987f \
 //x=26.155 //y=2.96 //x2=21.685 //y2=1.59
cc_1395 ( N_noxref_8_c_1827_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00302917f //x=26.155 //y=2.96 //x2=19.695 //y2=0.375
cc_1396 ( N_noxref_8_c_1827_n N_noxref_20_c_2886_n ) capacitor c=0.0247864f \
 //x=26.155 //y=2.96 //x2=22.57 //y2=2.08
cc_1397 ( N_noxref_8_c_1827_n N_noxref_20_c_2903_n ) capacitor c=0.0018311f \
 //x=26.155 //y=2.96 //x2=22.57 //y2=2.08
cc_1398 ( N_noxref_8_c_1827_n N_noxref_21_c_2989_n ) capacitor c=0.00838703f \
 //x=26.155 //y=2.96 //x2=22.91 //y2=1.665
cc_1399 ( N_noxref_8_c_1827_n N_noxref_21_c_2961_n ) capacitor c=0.0261317f \
 //x=26.155 //y=2.96 //x2=23.31 //y2=5.07
cc_1400 ( N_noxref_8_c_1834_n N_noxref_21_c_2961_n ) capacitor c=4.27463e-19 \
 //x=26.27 //y=2.08 //x2=23.31 //y2=5.07
cc_1401 ( N_noxref_8_c_1827_n N_noxref_22_c_3029_n ) capacitor c=0.00383675f \
 //x=26.155 //y=2.96 //x2=22.255 //y2=0.995
cc_1402 ( N_noxref_8_c_1827_n N_noxref_22_c_3035_n ) capacitor c=6.69632e-19 \
 //x=26.155 //y=2.96 //x2=23.225 //y2=0.54
cc_1403 ( N_noxref_8_c_1827_n N_noxref_22_M14_noxref_s ) capacitor \
 c=0.00324882f //x=26.155 //y=2.96 //x2=22.205 //y2=0.375
cc_1404 ( N_noxref_8_c_1827_n N_noxref_23_c_3083_n ) capacitor c=0.0278361f \
 //x=26.155 //y=2.96 //x2=25.16 //y2=2.08
cc_1405 ( N_noxref_8_c_1834_n N_noxref_23_c_3083_n ) capacitor c=0.0533123f \
 //x=26.27 //y=2.08 //x2=25.16 //y2=2.08
cc_1406 ( N_noxref_8_c_1918_p N_noxref_23_c_3083_n ) capacitor c=0.00231304f \
 //x=26.36 //y=1.915 //x2=25.16 //y2=2.08
cc_1407 ( N_noxref_8_c_1908_p N_noxref_23_c_3083_n ) capacitor c=0.00183762f \
 //x=26.27 //y=4.7 //x2=25.16 //y2=2.08
cc_1408 ( N_noxref_8_M50_noxref_g N_noxref_23_M48_noxref_g ) capacitor \
 c=0.0105869f //x=26.24 //y=6.02 //x2=25.36 //y2=6.02
cc_1409 ( N_noxref_8_M50_noxref_g N_noxref_23_M49_noxref_g ) capacitor \
 c=0.10632f //x=26.24 //y=6.02 //x2=25.8 //y2=6.02
cc_1410 ( N_noxref_8_M51_noxref_g N_noxref_23_M49_noxref_g ) capacitor \
 c=0.0101598f //x=26.68 //y=6.02 //x2=25.8 //y2=6.02
cc_1411 ( N_noxref_8_c_1981_p N_noxref_23_c_3084_n ) capacitor c=5.72482e-19 \
 //x=25.835 //y=0.91 //x2=24.86 //y2=0.875
cc_1412 ( N_noxref_8_c_1981_p N_noxref_23_c_3086_n ) capacitor c=0.00149976f \
 //x=25.835 //y=0.91 //x2=24.86 //y2=1.22
cc_1413 ( N_noxref_8_c_1983_p N_noxref_23_c_3087_n ) capacitor c=0.00111227f \
 //x=25.835 //y=1.22 //x2=24.86 //y2=1.53
cc_1414 ( N_noxref_8_c_1827_n N_noxref_23_c_3088_n ) capacitor c=0.00546863f \
 //x=26.155 //y=2.96 //x2=24.86 //y2=1.915
cc_1415 ( N_noxref_8_c_1834_n N_noxref_23_c_3088_n ) capacitor c=0.00238338f \
 //x=26.27 //y=2.08 //x2=24.86 //y2=1.915
cc_1416 ( N_noxref_8_c_1918_p N_noxref_23_c_3088_n ) capacitor c=0.00964411f \
 //x=26.36 //y=1.915 //x2=24.86 //y2=1.915
cc_1417 ( N_noxref_8_c_1981_p N_noxref_23_c_3091_n ) capacitor c=0.0160123f \
 //x=25.835 //y=0.91 //x2=25.39 //y2=0.875
cc_1418 ( N_noxref_8_c_1929_p N_noxref_23_c_3091_n ) capacitor c=0.00103227f \
 //x=26.36 //y=0.91 //x2=25.39 //y2=0.875
cc_1419 ( N_noxref_8_c_1983_p N_noxref_23_c_3093_n ) capacitor c=0.0124075f \
 //x=25.835 //y=1.22 //x2=25.39 //y2=1.22
cc_1420 ( N_noxref_8_c_1930_p N_noxref_23_c_3093_n ) capacitor c=0.0010154f \
 //x=26.36 //y=1.22 //x2=25.39 //y2=1.22
cc_1421 ( N_noxref_8_c_1931_p N_noxref_23_c_3093_n ) capacitor c=9.23422e-19 \
 //x=26.36 //y=1.45 //x2=25.39 //y2=1.22
cc_1422 ( N_noxref_8_c_1834_n N_noxref_23_c_3121_n ) capacitor c=0.00147352f \
 //x=26.27 //y=2.08 //x2=25.725 //y2=4.79
cc_1423 ( N_noxref_8_c_1908_p N_noxref_23_c_3121_n ) capacitor c=0.0168581f \
 //x=26.27 //y=4.7 //x2=25.725 //y2=4.79
cc_1424 ( N_noxref_8_c_1834_n N_noxref_23_c_3101_n ) capacitor c=0.00142741f \
 //x=26.27 //y=2.08 //x2=25.435 //y2=4.79
cc_1425 ( N_noxref_8_c_1908_p N_noxref_23_c_3101_n ) capacitor c=0.00484466f \
 //x=26.27 //y=4.7 //x2=25.435 //y2=4.79
cc_1426 ( N_noxref_8_c_1827_n N_noxref_24_c_3158_n ) capacitor c=0.00324882f \
 //x=26.155 //y=2.96 //x2=24.64 //y2=1.505
cc_1427 ( N_noxref_8_c_1827_n N_noxref_24_c_3144_n ) capacitor c=0.0127841f \
 //x=26.155 //y=2.96 //x2=25.525 //y2=1.59
cc_1428 ( N_noxref_8_c_1981_p N_noxref_24_c_3151_n ) capacitor c=0.0167228f \
 //x=25.835 //y=0.91 //x2=26.495 //y2=0.54
cc_1429 ( N_noxref_8_c_1929_p N_noxref_24_c_3151_n ) capacitor c=0.00534519f \
 //x=26.36 //y=0.91 //x2=26.495 //y2=0.54
cc_1430 ( N_noxref_8_c_1827_n N_noxref_24_c_3162_n ) capacitor c=0.00946209f \
 //x=26.155 //y=2.96 //x2=26.495 //y2=1.59
cc_1431 ( N_noxref_8_c_1834_n N_noxref_24_c_3162_n ) capacitor c=0.0121959f \
 //x=26.27 //y=2.08 //x2=26.495 //y2=1.59
cc_1432 ( N_noxref_8_c_1983_p N_noxref_24_c_3162_n ) capacitor c=0.0153476f \
 //x=25.835 //y=1.22 //x2=26.495 //y2=1.59
cc_1433 ( N_noxref_8_c_1918_p N_noxref_24_c_3162_n ) capacitor c=0.0225008f \
 //x=26.36 //y=1.915 //x2=26.495 //y2=1.59
cc_1434 ( N_noxref_8_c_1827_n N_noxref_24_M15_noxref_s ) capacitor \
 c=0.00324882f //x=26.155 //y=2.96 //x2=24.505 //y2=0.375
cc_1435 ( N_noxref_8_c_1981_p N_noxref_24_M15_noxref_s ) capacitor \
 c=0.00798959f //x=25.835 //y=0.91 //x2=24.505 //y2=0.375
cc_1436 ( N_noxref_8_c_1931_p N_noxref_24_M15_noxref_s ) capacitor \
 c=0.00212176f //x=26.36 //y=1.45 //x2=24.505 //y2=0.375
cc_1437 ( N_noxref_8_c_1918_p N_noxref_24_M15_noxref_s ) capacitor \
 c=0.00298115f //x=26.36 //y=1.915 //x2=24.505 //y2=0.375
cc_1438 ( N_noxref_8_c_1834_n N_noxref_25_c_3196_n ) capacitor c=0.0149705f \
 //x=26.27 //y=2.08 //x2=26.375 //y2=5.155
cc_1439 ( N_noxref_8_M50_noxref_g N_noxref_25_c_3196_n ) capacitor \
 c=0.0167692f //x=26.24 //y=6.02 //x2=26.375 //y2=5.155
cc_1440 ( N_noxref_8_c_1908_p N_noxref_25_c_3196_n ) capacitor c=0.00325274f \
 //x=26.27 //y=4.7 //x2=26.375 //y2=5.155
cc_1441 ( N_noxref_8_M51_noxref_g N_noxref_25_c_3202_n ) capacitor c=0.019179f \
 //x=26.68 //y=6.02 //x2=27.255 //y2=5.155
cc_1442 ( N_noxref_8_c_1834_n N_noxref_25_c_3210_n ) capacitor c=0.00362897f \
 //x=26.27 //y=2.08 //x2=28.12 //y2=5.07
cc_1443 ( N_noxref_8_c_1907_p N_noxref_25_c_3230_n ) capacitor c=0.00441288f \
 //x=26.605 //y=4.79 //x2=26.46 //y2=5.155
cc_1444 ( N_noxref_8_M50_noxref_g N_noxref_25_M50_noxref_d ) capacitor \
 c=0.0180032f //x=26.24 //y=6.02 //x2=26.315 //y2=5.02
cc_1445 ( N_noxref_8_M51_noxref_g N_noxref_25_M50_noxref_d ) capacitor \
 c=0.0180032f //x=26.68 //y=6.02 //x2=26.315 //y2=5.02
cc_1446 ( N_noxref_8_c_2016_p N_noxref_26_c_3271_n ) capacitor c=2.14837e-19 \
 //x=26.205 //y=0.755 //x2=27.065 //y2=0.995
cc_1447 ( N_noxref_8_c_1929_p N_noxref_26_c_3271_n ) capacitor c=0.00123426f \
 //x=26.36 //y=0.91 //x2=27.065 //y2=0.995
cc_1448 ( N_noxref_8_c_1930_p N_noxref_26_c_3271_n ) capacitor c=0.0129288f \
 //x=26.36 //y=1.22 //x2=27.065 //y2=0.995
cc_1449 ( N_noxref_8_c_1931_p N_noxref_26_c_3271_n ) capacitor c=0.00142359f \
 //x=26.36 //y=1.45 //x2=27.065 //y2=0.995
cc_1450 ( N_noxref_8_c_1981_p N_noxref_26_M16_noxref_d ) capacitor \
 c=0.00223875f //x=25.835 //y=0.91 //x2=25.91 //y2=0.91
cc_1451 ( N_noxref_8_c_1983_p N_noxref_26_M16_noxref_d ) capacitor \
 c=0.00262485f //x=25.835 //y=1.22 //x2=25.91 //y2=0.91
cc_1452 ( N_noxref_8_c_2016_p N_noxref_26_M16_noxref_d ) capacitor \
 c=0.00220746f //x=26.205 //y=0.755 //x2=25.91 //y2=0.91
cc_1453 ( N_noxref_8_c_2023_p N_noxref_26_M16_noxref_d ) capacitor \
 c=0.00194798f //x=26.205 //y=1.375 //x2=25.91 //y2=0.91
cc_1454 ( N_noxref_8_c_1929_p N_noxref_26_M16_noxref_d ) capacitor \
 c=0.00198465f //x=26.36 //y=0.91 //x2=25.91 //y2=0.91
cc_1455 ( N_noxref_8_c_1930_p N_noxref_26_M16_noxref_d ) capacitor \
 c=0.00128384f //x=26.36 //y=1.22 //x2=25.91 //y2=0.91
cc_1456 ( N_noxref_8_c_1929_p N_noxref_26_M17_noxref_s ) capacitor \
 c=7.21316e-19 //x=26.36 //y=0.91 //x2=27.015 //y2=0.375
cc_1457 ( N_noxref_8_c_1930_p N_noxref_26_M17_noxref_s ) capacitor \
 c=0.00348171f //x=26.36 //y=1.22 //x2=27.015 //y2=0.375
cc_1458 ( N_noxref_9_c_2029_n N_noxref_14_c_2577_n ) capacitor c=0.00204385f \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_1459 ( N_noxref_9_c_2151_n N_noxref_14_c_2577_n ) capacitor c=0.0194423f \
 //x=8.13 //y=0.915 //x2=8.795 //y2=0.54
cc_1460 ( N_noxref_9_c_2194_n N_noxref_14_c_2577_n ) capacitor c=0.00656458f \
 //x=8.66 //y=0.915 //x2=8.795 //y2=0.54
cc_1461 ( N_noxref_9_c_2154_n N_noxref_14_c_2577_n ) capacitor c=2.20712e-19 \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_1462 ( N_noxref_9_c_2152_n N_noxref_14_c_2600_n ) capacitor c=0.00538829f \
 //x=8.13 //y=1.26 //x2=7.91 //y2=0.995
cc_1463 ( N_noxref_9_c_2151_n N_noxref_14_M5_noxref_s ) capacitor \
 c=0.00538829f //x=8.13 //y=0.915 //x2=7.775 //y2=0.375
cc_1464 ( N_noxref_9_c_2153_n N_noxref_14_M5_noxref_s ) capacitor \
 c=0.00538829f //x=8.13 //y=1.57 //x2=7.775 //y2=0.375
cc_1465 ( N_noxref_9_c_2194_n N_noxref_14_M5_noxref_s ) capacitor c=0.0143002f \
 //x=8.66 //y=0.915 //x2=7.775 //y2=0.375
cc_1466 ( N_noxref_9_c_2195_n N_noxref_14_M5_noxref_s ) capacitor \
 c=0.00290153f //x=8.66 //y=1.26 //x2=7.775 //y2=0.375
cc_1467 ( N_noxref_9_c_2030_n N_noxref_16_c_2681_n ) capacitor c=0.00204385f \
 //x=12.95 //y=2.08 //x2=13.605 //y2=0.54
cc_1468 ( N_noxref_9_c_2110_n N_noxref_16_c_2681_n ) capacitor c=0.0194423f \
 //x=12.94 //y=0.915 //x2=13.605 //y2=0.54
cc_1469 ( N_noxref_9_c_2116_n N_noxref_16_c_2681_n ) capacitor c=0.00656458f \
 //x=13.47 //y=0.915 //x2=13.605 //y2=0.54
cc_1470 ( N_noxref_9_c_2119_n N_noxref_16_c_2681_n ) capacitor c=2.20712e-19 \
 //x=12.95 //y=2.08 //x2=13.605 //y2=0.54
cc_1471 ( N_noxref_9_c_2111_n N_noxref_16_c_2692_n ) capacitor c=0.00538829f \
 //x=12.94 //y=1.26 //x2=12.72 //y2=0.995
cc_1472 ( N_noxref_9_c_2110_n N_noxref_16_M8_noxref_s ) capacitor \
 c=0.00538829f //x=12.94 //y=0.915 //x2=12.585 //y2=0.375
cc_1473 ( N_noxref_9_c_2112_n N_noxref_16_M8_noxref_s ) capacitor \
 c=0.00538829f //x=12.94 //y=1.57 //x2=12.585 //y2=0.375
cc_1474 ( N_noxref_9_c_2116_n N_noxref_16_M8_noxref_s ) capacitor c=0.0143002f \
 //x=13.47 //y=0.915 //x2=12.585 //y2=0.375
cc_1475 ( N_noxref_9_c_2117_n N_noxref_16_M8_noxref_s ) capacitor \
 c=0.00290153f //x=13.47 //y=1.26 //x2=12.585 //y2=0.375
cc_1476 ( N_noxref_9_M11_noxref_d N_noxref_17_M9_noxref_s ) capacitor \
 c=0.00309936f //x=17.825 //y=0.915 //x2=14.885 //y2=0.375
cc_1477 ( N_noxref_9_c_2031_n N_noxref_18_c_2785_n ) capacitor c=0.00457167f \
 //x=18.415 //y=1.665 //x2=18.415 //y2=0.54
cc_1478 ( N_noxref_9_M11_noxref_d N_noxref_18_c_2785_n ) capacitor \
 c=0.0115903f //x=17.825 //y=0.915 //x2=18.415 //y2=0.54
cc_1479 ( N_noxref_9_c_2218_n N_noxref_18_c_2813_n ) capacitor c=0.0200405f \
 //x=18.1 //y=1.665 //x2=17.53 //y2=0.995
cc_1480 ( N_noxref_9_M11_noxref_d N_noxref_18_M10_noxref_d ) capacitor \
 c=5.27807e-19 //x=17.825 //y=0.915 //x2=16.29 //y2=0.91
cc_1481 ( N_noxref_9_c_2031_n N_noxref_18_M11_noxref_s ) capacitor \
 c=0.0196084f //x=18.415 //y=1.665 //x2=17.395 //y2=0.375
cc_1482 ( N_noxref_9_M11_noxref_d N_noxref_18_M11_noxref_s ) capacitor \
 c=0.0426368f //x=17.825 //y=0.915 //x2=17.395 //y2=0.375
cc_1483 ( N_noxref_9_c_2031_n N_noxref_19_c_2850_n ) capacitor c=3.84569e-19 \
 //x=18.415 //y=1.665 //x2=19.83 //y2=1.505
cc_1484 ( N_noxref_9_M11_noxref_d N_noxref_19_M12_noxref_s ) capacitor \
 c=2.55333e-19 //x=17.825 //y=0.915 //x2=19.695 //y2=0.375
cc_1485 ( N_noxref_9_c_2028_n N_noxref_20_c_2886_n ) capacitor c=0.0250607f \
 //x=27.265 //y=3.7 //x2=22.57 //y2=2.08
cc_1486 ( N_noxref_9_c_2028_n N_noxref_20_c_2907_n ) capacitor c=0.00684517f \
 //x=27.265 //y=3.7 //x2=22.57 //y2=4.7
cc_1487 ( N_noxref_9_c_2028_n N_noxref_21_c_2947_n ) capacitor c=0.0194603f \
 //x=27.265 //y=3.7 //x2=21.565 //y2=5.155
cc_1488 ( N_noxref_9_c_2028_n N_noxref_21_c_2951_n ) capacitor c=0.0135617f \
 //x=27.265 //y=3.7 //x2=20.855 //y2=5.155
cc_1489 ( N_noxref_9_c_2055_n N_noxref_21_c_2951_n ) capacitor c=3.10026e-19 \
 //x=18.415 //y=5.155 //x2=20.855 //y2=5.155
cc_1490 ( N_noxref_9_c_2028_n N_noxref_21_c_2957_n ) capacitor c=0.0109339f \
 //x=27.265 //y=3.7 //x2=23.225 //y2=5.155
cc_1491 ( N_noxref_9_c_2028_n N_noxref_21_c_2961_n ) capacitor c=0.0265608f \
 //x=27.265 //y=3.7 //x2=23.31 //y2=5.07
cc_1492 ( N_noxref_9_c_2028_n N_noxref_23_c_3083_n ) capacitor c=0.0268219f \
 //x=27.265 //y=3.7 //x2=25.16 //y2=2.08
cc_1493 ( N_noxref_9_c_2032_n N_noxref_23_c_3083_n ) capacitor c=0.00145664f \
 //x=27.38 //y=2.08 //x2=25.16 //y2=2.08
cc_1494 ( N_noxref_9_c_2028_n N_noxref_23_c_3101_n ) capacitor c=0.0129605f \
 //x=27.265 //y=3.7 //x2=25.435 //y2=4.79
cc_1495 ( N_noxref_9_c_2028_n N_noxref_24_c_3162_n ) capacitor c=0.00102279f \
 //x=27.265 //y=3.7 //x2=26.495 //y2=1.59
cc_1496 ( N_noxref_9_c_2028_n N_noxref_24_M15_noxref_s ) capacitor \
 c=0.00155863f //x=27.265 //y=3.7 //x2=24.505 //y2=0.375
cc_1497 ( N_noxref_9_c_2028_n N_noxref_25_c_3196_n ) capacitor c=0.0184004f \
 //x=27.265 //y=3.7 //x2=26.375 //y2=5.155
cc_1498 ( N_noxref_9_c_2028_n N_noxref_25_c_3200_n ) capacitor c=0.0135617f \
 //x=27.265 //y=3.7 //x2=25.665 //y2=5.155
cc_1499 ( N_noxref_9_M52_noxref_g N_noxref_25_c_3202_n ) capacitor c=0.019179f \
 //x=27.12 //y=6.02 //x2=27.255 //y2=5.155
cc_1500 ( N_noxref_9_c_2028_n N_noxref_25_c_3206_n ) capacitor c=0.00151992f \
 //x=27.265 //y=3.7 //x2=28.035 //y2=5.155
cc_1501 ( N_noxref_9_M53_noxref_g N_noxref_25_c_3206_n ) capacitor \
 c=0.0225988f //x=27.56 //y=6.02 //x2=28.035 //y2=5.155
cc_1502 ( N_noxref_9_c_2284_n N_noxref_25_c_3206_n ) capacitor c=0.00201851f \
 //x=27.38 //y=4.7 //x2=28.035 //y2=5.155
cc_1503 ( N_noxref_9_c_2332_p N_noxref_25_c_3194_n ) capacitor c=0.00359704f \
 //x=27.745 //y=1.415 //x2=28.035 //y2=1.665
cc_1504 ( N_noxref_9_c_2333_p N_noxref_25_c_3194_n ) capacitor c=0.00457401f \
 //x=27.9 //y=1.26 //x2=28.035 //y2=1.665
cc_1505 ( N_noxref_9_c_2028_n N_noxref_25_c_3210_n ) capacitor c=0.00599141f \
 //x=27.265 //y=3.7 //x2=28.12 //y2=5.07
cc_1506 ( N_noxref_9_c_2032_n N_noxref_25_c_3210_n ) capacitor c=0.0911412f \
 //x=27.38 //y=2.08 //x2=28.12 //y2=5.07
cc_1507 ( N_noxref_9_c_2281_n N_noxref_25_c_3210_n ) capacitor c=0.00877984f \
 //x=27.38 //y=2.08 //x2=28.12 //y2=5.07
cc_1508 ( N_noxref_9_c_2283_n N_noxref_25_c_3210_n ) capacitor c=0.00283672f \
 //x=27.38 //y=1.915 //x2=28.12 //y2=5.07
cc_1509 ( N_noxref_9_c_2284_n N_noxref_25_c_3210_n ) capacitor c=0.013844f \
 //x=27.38 //y=4.7 //x2=28.12 //y2=5.07
cc_1510 ( N_noxref_9_c_2028_n N_noxref_25_c_3246_n ) capacitor c=5.53707e-19 \
 //x=27.265 //y=3.7 //x2=27.34 //y2=5.155
cc_1511 ( N_noxref_9_c_2032_n N_noxref_25_c_3246_n ) capacitor c=0.017024f \
 //x=27.38 //y=2.08 //x2=27.34 //y2=5.155
cc_1512 ( N_noxref_9_c_2284_n N_noxref_25_c_3246_n ) capacitor c=0.00476349f \
 //x=27.38 //y=4.7 //x2=27.34 //y2=5.155
cc_1513 ( N_noxref_9_c_2272_n N_noxref_25_M17_noxref_d ) capacitor \
 c=0.00217566f //x=27.37 //y=0.915 //x2=27.445 //y2=0.915
cc_1514 ( N_noxref_9_c_2273_n N_noxref_25_M17_noxref_d ) capacitor \
 c=0.0034598f //x=27.37 //y=1.26 //x2=27.445 //y2=0.915
cc_1515 ( N_noxref_9_c_2274_n N_noxref_25_M17_noxref_d ) capacitor \
 c=0.00544291f //x=27.37 //y=1.57 //x2=27.445 //y2=0.915
cc_1516 ( N_noxref_9_c_2345_p N_noxref_25_M17_noxref_d ) capacitor \
 c=0.00241102f //x=27.745 //y=0.76 //x2=27.445 //y2=0.915
cc_1517 ( N_noxref_9_c_2332_p N_noxref_25_M17_noxref_d ) capacitor \
 c=0.0140297f //x=27.745 //y=1.415 //x2=27.445 //y2=0.915
cc_1518 ( N_noxref_9_c_2347_p N_noxref_25_M17_noxref_d ) capacitor \
 c=0.00219619f //x=27.9 //y=0.915 //x2=27.445 //y2=0.915
cc_1519 ( N_noxref_9_c_2333_p N_noxref_25_M17_noxref_d ) capacitor \
 c=0.00603828f //x=27.9 //y=1.26 //x2=27.445 //y2=0.915
cc_1520 ( N_noxref_9_c_2283_n N_noxref_25_M17_noxref_d ) capacitor \
 c=0.00661782f //x=27.38 //y=1.915 //x2=27.445 //y2=0.915
cc_1521 ( N_noxref_9_M52_noxref_g N_noxref_25_M52_noxref_d ) capacitor \
 c=0.0180032f //x=27.12 //y=6.02 //x2=27.195 //y2=5.02
cc_1522 ( N_noxref_9_M53_noxref_g N_noxref_25_M52_noxref_d ) capacitor \
 c=0.0194246f //x=27.56 //y=6.02 //x2=27.195 //y2=5.02
cc_1523 ( N_noxref_9_c_2028_n N_noxref_26_c_3271_n ) capacitor c=0.00200649f \
 //x=27.265 //y=3.7 //x2=27.065 //y2=0.995
cc_1524 ( N_noxref_9_c_2028_n N_noxref_26_c_3276_n ) capacitor c=2.6387e-19 \
 //x=27.265 //y=3.7 //x2=28.035 //y2=0.54
cc_1525 ( N_noxref_9_c_2032_n N_noxref_26_c_3276_n ) capacitor c=0.00209081f \
 //x=27.38 //y=2.08 //x2=28.035 //y2=0.54
cc_1526 ( N_noxref_9_c_2272_n N_noxref_26_c_3276_n ) capacitor c=0.0193963f \
 //x=27.37 //y=0.915 //x2=28.035 //y2=0.54
cc_1527 ( N_noxref_9_c_2347_p N_noxref_26_c_3276_n ) capacitor c=0.00656458f \
 //x=27.9 //y=0.915 //x2=28.035 //y2=0.54
cc_1528 ( N_noxref_9_c_2281_n N_noxref_26_c_3276_n ) capacitor c=2.20712e-19 \
 //x=27.38 //y=2.08 //x2=28.035 //y2=0.54
cc_1529 ( N_noxref_9_c_2273_n N_noxref_26_c_3301_n ) capacitor c=0.00538829f \
 //x=27.37 //y=1.26 //x2=27.15 //y2=0.995
cc_1530 ( N_noxref_9_c_2028_n N_noxref_26_M17_noxref_s ) capacitor \
 c=0.0016894f //x=27.265 //y=3.7 //x2=27.015 //y2=0.375
cc_1531 ( N_noxref_9_c_2272_n N_noxref_26_M17_noxref_s ) capacitor \
 c=0.00538829f //x=27.37 //y=0.915 //x2=27.015 //y2=0.375
cc_1532 ( N_noxref_9_c_2274_n N_noxref_26_M17_noxref_s ) capacitor \
 c=0.00538829f //x=27.37 //y=1.57 //x2=27.015 //y2=0.375
cc_1533 ( N_noxref_9_c_2347_p N_noxref_26_M17_noxref_s ) capacitor \
 c=0.0143002f //x=27.9 //y=0.915 //x2=27.015 //y2=0.375
cc_1534 ( N_noxref_9_c_2333_p N_noxref_26_M17_noxref_s ) capacitor \
 c=0.00290153f //x=27.9 //y=1.26 //x2=27.015 //y2=0.375
cc_1535 ( N_noxref_10_c_2369_n N_noxref_11_c_2449_n ) capacitor c=0.0034165f \
 //x=0.81 //y=1.915 //x2=0.59 //y2=1.505
cc_1536 ( N_noxref_10_c_2364_n N_noxref_11_c_2421_n ) capacitor c=0.0122915f \
 //x=1.11 //y=2.08 //x2=1.475 //y2=1.59
cc_1537 ( N_noxref_10_c_2368_n N_noxref_11_c_2421_n ) capacitor c=0.00703864f \
 //x=0.81 //y=1.53 //x2=1.475 //y2=1.59
cc_1538 ( N_noxref_10_c_2369_n N_noxref_11_c_2421_n ) capacitor c=0.0259045f \
 //x=0.81 //y=1.915 //x2=1.475 //y2=1.59
cc_1539 ( N_noxref_10_c_2371_n N_noxref_11_c_2421_n ) capacitor c=0.00708583f \
 //x=1.185 //y=1.375 //x2=1.475 //y2=1.59
cc_1540 ( N_noxref_10_c_2374_n N_noxref_11_c_2421_n ) capacitor c=0.00698822f \
 //x=1.34 //y=1.22 //x2=1.475 //y2=1.59
cc_1541 ( N_noxref_10_c_2365_n N_noxref_11_M0_noxref_s ) capacitor \
 c=0.0327271f //x=0.81 //y=0.875 //x2=0.455 //y2=0.375
cc_1542 ( N_noxref_10_c_2368_n N_noxref_11_M0_noxref_s ) capacitor \
 c=7.99997e-19 //x=0.81 //y=1.53 //x2=0.455 //y2=0.375
cc_1543 ( N_noxref_10_c_2369_n N_noxref_11_M0_noxref_s ) capacitor \
 c=0.00122123f //x=0.81 //y=1.915 //x2=0.455 //y2=0.375
cc_1544 ( N_noxref_10_c_2372_n N_noxref_11_M0_noxref_s ) capacitor \
 c=0.0121427f //x=1.34 //y=0.875 //x2=0.455 //y2=0.375
cc_1545 ( N_noxref_11_c_2428_n N_noxref_12_c_2467_n ) capacitor c=0.0131801f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_1546 ( N_noxref_11_c_2440_n N_noxref_12_c_2467_n ) capacitor c=0.00980353f \
 //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_1547 ( N_noxref_11_M0_noxref_s N_noxref_12_c_2467_n ) capacitor \
 c=0.0221661f //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_1548 ( N_noxref_11_M0_noxref_s N_noxref_12_c_2470_n ) capacitor \
 c=0.0180035f //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_1549 ( N_noxref_11_c_2428_n N_noxref_12_M1_noxref_d ) capacitor \
 c=0.0128687f //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_1550 ( N_noxref_11_c_2440_n N_noxref_12_M1_noxref_d ) capacitor c=0.008922f \
 //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_1551 ( N_noxref_11_M0_noxref_s N_noxref_12_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_1552 ( N_noxref_11_M0_noxref_s N_noxref_12_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_1553 ( N_noxref_12_c_2476_n N_noxref_13_M3_noxref_s ) capacitor \
 c=0.00191848f //x=4.07 //y=0.625 //x2=5.265 //y2=0.375
cc_1554 ( N_noxref_13_c_2528_n N_noxref_14_c_2571_n ) capacitor c=0.0131877f \
 //x=7.255 //y=0.54 //x2=7.825 //y2=0.995
cc_1555 ( N_noxref_13_c_2551_n N_noxref_14_c_2571_n ) capacitor c=0.00981707f \
 //x=7.255 //y=1.59 //x2=7.825 //y2=0.995
cc_1556 ( N_noxref_13_M3_noxref_s N_noxref_14_c_2571_n ) capacitor \
 c=0.0221661f //x=5.265 //y=0.375 //x2=7.825 //y2=0.995
cc_1557 ( N_noxref_13_M3_noxref_s N_noxref_14_c_2574_n ) capacitor \
 c=0.0180035f //x=5.265 //y=0.375 //x2=7.91 //y2=0.625
cc_1558 ( N_noxref_13_c_2528_n N_noxref_14_M4_noxref_d ) capacitor \
 c=0.0127191f //x=7.255 //y=0.54 //x2=6.67 //y2=0.91
cc_1559 ( N_noxref_13_c_2551_n N_noxref_14_M4_noxref_d ) capacitor \
 c=0.00861161f //x=7.255 //y=1.59 //x2=6.67 //y2=0.91
cc_1560 ( N_noxref_13_M3_noxref_s N_noxref_14_M4_noxref_d ) capacitor \
 c=0.0159202f //x=5.265 //y=0.375 //x2=6.67 //y2=0.91
cc_1561 ( N_noxref_13_M3_noxref_s N_noxref_14_M5_noxref_s ) capacitor \
 c=0.0213553f //x=5.265 //y=0.375 //x2=7.775 //y2=0.375
cc_1562 ( N_noxref_14_c_2580_n N_noxref_15_M6_noxref_s ) capacitor \
 c=0.00191848f //x=8.88 //y=0.625 //x2=10.075 //y2=0.375
cc_1563 ( N_noxref_15_c_2632_n N_noxref_16_c_2675_n ) capacitor c=0.0131877f \
 //x=12.065 //y=0.54 //x2=12.635 //y2=0.995
cc_1564 ( N_noxref_15_c_2656_n N_noxref_16_c_2675_n ) capacitor c=0.00981707f \
 //x=12.065 //y=1.59 //x2=12.635 //y2=0.995
cc_1565 ( N_noxref_15_M6_noxref_s N_noxref_16_c_2675_n ) capacitor \
 c=0.0221661f //x=10.075 //y=0.375 //x2=12.635 //y2=0.995
cc_1566 ( N_noxref_15_M6_noxref_s N_noxref_16_c_2678_n ) capacitor \
 c=0.0180035f //x=10.075 //y=0.375 //x2=12.72 //y2=0.625
cc_1567 ( N_noxref_15_c_2632_n N_noxref_16_M7_noxref_d ) capacitor \
 c=0.0127191f //x=12.065 //y=0.54 //x2=11.48 //y2=0.91
cc_1568 ( N_noxref_15_c_2656_n N_noxref_16_M7_noxref_d ) capacitor \
 c=0.00861161f //x=12.065 //y=1.59 //x2=11.48 //y2=0.91
cc_1569 ( N_noxref_15_M6_noxref_s N_noxref_16_M7_noxref_d ) capacitor \
 c=0.0159202f //x=10.075 //y=0.375 //x2=11.48 //y2=0.91
cc_1570 ( N_noxref_15_M6_noxref_s N_noxref_16_M8_noxref_s ) capacitor \
 c=0.0213553f //x=10.075 //y=0.375 //x2=12.585 //y2=0.375
cc_1571 ( N_noxref_16_c_2684_n N_noxref_17_M9_noxref_s ) capacitor \
 c=0.00191848f //x=13.69 //y=0.625 //x2=14.885 //y2=0.375
cc_1572 ( N_noxref_17_c_2736_n N_noxref_18_c_2779_n ) capacitor c=0.0131877f \
 //x=16.875 //y=0.54 //x2=17.445 //y2=0.995
cc_1573 ( N_noxref_17_c_2759_n N_noxref_18_c_2779_n ) capacitor c=0.00981707f \
 //x=16.875 //y=1.59 //x2=17.445 //y2=0.995
cc_1574 ( N_noxref_17_M9_noxref_s N_noxref_18_c_2779_n ) capacitor \
 c=0.0221661f //x=14.885 //y=0.375 //x2=17.445 //y2=0.995
cc_1575 ( N_noxref_17_M9_noxref_s N_noxref_18_c_2782_n ) capacitor \
 c=0.0180035f //x=14.885 //y=0.375 //x2=17.53 //y2=0.625
cc_1576 ( N_noxref_17_c_2736_n N_noxref_18_M10_noxref_d ) capacitor \
 c=0.0127191f //x=16.875 //y=0.54 //x2=16.29 //y2=0.91
cc_1577 ( N_noxref_17_c_2759_n N_noxref_18_M10_noxref_d ) capacitor \
 c=0.00861161f //x=16.875 //y=1.59 //x2=16.29 //y2=0.91
cc_1578 ( N_noxref_17_M9_noxref_s N_noxref_18_M10_noxref_d ) capacitor \
 c=0.0159202f //x=14.885 //y=0.375 //x2=16.29 //y2=0.91
cc_1579 ( N_noxref_17_M9_noxref_s N_noxref_18_M11_noxref_s ) capacitor \
 c=0.0213553f //x=14.885 //y=0.375 //x2=17.395 //y2=0.375
cc_1580 ( N_noxref_18_c_2788_n N_noxref_19_M12_noxref_s ) capacitor \
 c=0.00191848f //x=18.5 //y=0.625 //x2=19.695 //y2=0.375
cc_1581 ( N_noxref_19_M12_noxref_s N_noxref_21_M14_noxref_d ) capacitor \
 c=0.00309936f //x=19.695 //y=0.375 //x2=22.635 //y2=0.915
cc_1582 ( N_noxref_19_c_2841_n N_noxref_22_c_3029_n ) capacitor c=0.0132328f \
 //x=21.685 //y=0.54 //x2=22.255 //y2=0.995
cc_1583 ( N_noxref_19_c_2864_n N_noxref_22_c_3029_n ) capacitor c=0.00988406f \
 //x=21.685 //y=1.59 //x2=22.255 //y2=0.995
cc_1584 ( N_noxref_19_M12_noxref_s N_noxref_22_c_3029_n ) capacitor \
 c=0.0226274f //x=19.695 //y=0.375 //x2=22.255 //y2=0.995
cc_1585 ( N_noxref_19_M12_noxref_s N_noxref_22_c_3032_n ) capacitor \
 c=0.0180035f //x=19.695 //y=0.375 //x2=22.34 //y2=0.625
cc_1586 ( N_noxref_19_c_2841_n N_noxref_22_M13_noxref_d ) capacitor \
 c=0.0127176f //x=21.685 //y=0.54 //x2=21.1 //y2=0.91
cc_1587 ( N_noxref_19_c_2864_n N_noxref_22_M13_noxref_d ) capacitor \
 c=0.0086073f //x=21.685 //y=1.59 //x2=21.1 //y2=0.91
cc_1588 ( N_noxref_19_M12_noxref_s N_noxref_22_M13_noxref_d ) capacitor \
 c=0.0159202f //x=19.695 //y=0.375 //x2=21.1 //y2=0.91
cc_1589 ( N_noxref_19_M12_noxref_s N_noxref_22_M14_noxref_s ) capacitor \
 c=0.0213553f //x=19.695 //y=0.375 //x2=22.205 //y2=0.375
cc_1590 ( N_noxref_20_M46_noxref_g N_noxref_21_c_2953_n ) capacitor \
 c=0.019179f //x=22.31 //y=6.02 //x2=22.445 //y2=5.155
cc_1591 ( N_noxref_20_M47_noxref_g N_noxref_21_c_2957_n ) capacitor \
 c=0.0213171f //x=22.75 //y=6.02 //x2=23.225 //y2=5.155
cc_1592 ( N_noxref_20_c_2907_n N_noxref_21_c_2957_n ) capacitor c=0.00201851f \
 //x=22.57 //y=4.7 //x2=23.225 //y2=5.155
cc_1593 ( N_noxref_20_c_2917_p N_noxref_21_c_2945_n ) capacitor c=0.00359704f \
 //x=22.935 //y=1.415 //x2=23.225 //y2=1.665
cc_1594 ( N_noxref_20_c_2918_p N_noxref_21_c_2945_n ) capacitor c=0.00457401f \
 //x=23.09 //y=1.26 //x2=23.225 //y2=1.665
cc_1595 ( N_noxref_20_c_2886_n N_noxref_21_c_2961_n ) capacitor c=0.0875874f \
 //x=22.57 //y=2.08 //x2=23.31 //y2=5.07
cc_1596 ( N_noxref_20_c_2903_n N_noxref_21_c_2961_n ) capacitor c=0.00772308f \
 //x=22.57 //y=2.08 //x2=23.31 //y2=5.07
cc_1597 ( N_noxref_20_c_2906_n N_noxref_21_c_2961_n ) capacitor c=0.00283672f \
 //x=22.57 //y=1.915 //x2=23.31 //y2=5.07
cc_1598 ( N_noxref_20_c_2907_n N_noxref_21_c_2961_n ) capacitor c=0.013844f \
 //x=22.57 //y=4.7 //x2=23.31 //y2=5.07
cc_1599 ( N_noxref_20_c_2886_n N_noxref_21_c_3007_n ) capacitor c=0.0171771f \
 //x=22.57 //y=2.08 //x2=22.53 //y2=5.155
cc_1600 ( N_noxref_20_c_2907_n N_noxref_21_c_3007_n ) capacitor c=0.00476349f \
 //x=22.57 //y=4.7 //x2=22.53 //y2=5.155
cc_1601 ( N_noxref_20_c_2900_n N_noxref_21_M14_noxref_d ) capacitor \
 c=0.00217566f //x=22.56 //y=0.915 //x2=22.635 //y2=0.915
cc_1602 ( N_noxref_20_c_2901_n N_noxref_21_M14_noxref_d ) capacitor \
 c=0.0034598f //x=22.56 //y=1.26 //x2=22.635 //y2=0.915
cc_1603 ( N_noxref_20_c_2902_n N_noxref_21_M14_noxref_d ) capacitor \
 c=0.00544291f //x=22.56 //y=1.57 //x2=22.635 //y2=0.915
cc_1604 ( N_noxref_20_c_2928_p N_noxref_21_M14_noxref_d ) capacitor \
 c=0.00241102f //x=22.935 //y=0.76 //x2=22.635 //y2=0.915
cc_1605 ( N_noxref_20_c_2917_p N_noxref_21_M14_noxref_d ) capacitor \
 c=0.0140297f //x=22.935 //y=1.415 //x2=22.635 //y2=0.915
cc_1606 ( N_noxref_20_c_2930_p N_noxref_21_M14_noxref_d ) capacitor \
 c=0.00219619f //x=23.09 //y=0.915 //x2=22.635 //y2=0.915
cc_1607 ( N_noxref_20_c_2918_p N_noxref_21_M14_noxref_d ) capacitor \
 c=0.00603828f //x=23.09 //y=1.26 //x2=22.635 //y2=0.915
cc_1608 ( N_noxref_20_c_2906_n N_noxref_21_M14_noxref_d ) capacitor \
 c=0.00661782f //x=22.57 //y=1.915 //x2=22.635 //y2=0.915
cc_1609 ( N_noxref_20_M46_noxref_g N_noxref_21_M46_noxref_d ) capacitor \
 c=0.0180032f //x=22.31 //y=6.02 //x2=22.385 //y2=5.02
cc_1610 ( N_noxref_20_M47_noxref_g N_noxref_21_M46_noxref_d ) capacitor \
 c=0.0194246f //x=22.75 //y=6.02 //x2=22.385 //y2=5.02
cc_1611 ( N_noxref_20_c_2886_n N_noxref_22_c_3035_n ) capacitor c=0.00207733f \
 //x=22.57 //y=2.08 //x2=23.225 //y2=0.54
cc_1612 ( N_noxref_20_c_2900_n N_noxref_22_c_3035_n ) capacitor c=0.0194423f \
 //x=22.56 //y=0.915 //x2=23.225 //y2=0.54
cc_1613 ( N_noxref_20_c_2930_p N_noxref_22_c_3035_n ) capacitor c=0.00656458f \
 //x=23.09 //y=0.915 //x2=23.225 //y2=0.54
cc_1614 ( N_noxref_20_c_2903_n N_noxref_22_c_3035_n ) capacitor c=2.20712e-19 \
 //x=22.57 //y=2.08 //x2=23.225 //y2=0.54
cc_1615 ( N_noxref_20_c_2901_n N_noxref_22_c_3071_n ) capacitor c=0.00538829f \
 //x=22.56 //y=1.26 //x2=22.34 //y2=0.995
cc_1616 ( N_noxref_20_c_2900_n N_noxref_22_M14_noxref_s ) capacitor \
 c=0.00538829f //x=22.56 //y=0.915 //x2=22.205 //y2=0.375
cc_1617 ( N_noxref_20_c_2902_n N_noxref_22_M14_noxref_s ) capacitor \
 c=0.00538829f //x=22.56 //y=1.57 //x2=22.205 //y2=0.375
cc_1618 ( N_noxref_20_c_2930_p N_noxref_22_M14_noxref_s ) capacitor \
 c=0.0143002f //x=23.09 //y=0.915 //x2=22.205 //y2=0.375
cc_1619 ( N_noxref_20_c_2918_p N_noxref_22_M14_noxref_s ) capacitor \
 c=0.00290153f //x=23.09 //y=1.26 //x2=22.205 //y2=0.375
cc_1620 ( N_noxref_20_c_2886_n N_noxref_23_c_3083_n ) capacitor c=7.46474e-19 \
 //x=22.57 //y=2.08 //x2=25.16 //y2=2.08
cc_1621 ( N_noxref_21_c_2945_n N_noxref_22_c_3035_n ) capacitor c=0.00464291f \
 //x=23.225 //y=1.665 //x2=23.225 //y2=0.54
cc_1622 ( N_noxref_21_M14_noxref_d N_noxref_22_c_3035_n ) capacitor \
 c=0.0117407f //x=22.635 //y=0.915 //x2=23.225 //y2=0.54
cc_1623 ( N_noxref_21_c_2989_n N_noxref_22_c_3071_n ) capacitor c=0.0200405f \
 //x=22.91 //y=1.665 //x2=22.34 //y2=0.995
cc_1624 ( N_noxref_21_M14_noxref_d N_noxref_22_M13_noxref_d ) capacitor \
 c=5.27807e-19 //x=22.635 //y=0.915 //x2=21.1 //y2=0.91
cc_1625 ( N_noxref_21_c_2945_n N_noxref_22_M14_noxref_s ) capacitor \
 c=0.0205269f //x=23.225 //y=1.665 //x2=22.205 //y2=0.375
cc_1626 ( N_noxref_21_M14_noxref_d N_noxref_22_M14_noxref_s ) capacitor \
 c=0.0426368f //x=22.635 //y=0.915 //x2=22.205 //y2=0.375
cc_1627 ( N_noxref_21_c_2961_n N_noxref_23_c_3083_n ) capacitor c=0.0145933f \
 //x=23.31 //y=5.07 //x2=25.16 //y2=2.08
cc_1628 ( N_noxref_21_c_2945_n N_noxref_24_c_3158_n ) capacitor c=3.84569e-19 \
 //x=23.225 //y=1.665 //x2=24.64 //y2=1.505
cc_1629 ( N_noxref_21_M14_noxref_d N_noxref_24_M15_noxref_s ) capacitor \
 c=2.55333e-19 //x=22.635 //y=0.915 //x2=24.505 //y2=0.375
cc_1630 ( N_noxref_21_c_2957_n N_noxref_25_c_3200_n ) capacitor c=3.10026e-19 \
 //x=23.225 //y=5.155 //x2=25.665 //y2=5.155
cc_1631 ( N_noxref_22_c_3038_n N_noxref_24_M15_noxref_s ) capacitor \
 c=0.00191848f //x=23.31 //y=0.625 //x2=24.505 //y2=0.375
cc_1632 ( N_noxref_23_c_3088_n N_noxref_24_c_3158_n ) capacitor c=0.0034165f \
 //x=24.86 //y=1.915 //x2=24.64 //y2=1.505
cc_1633 ( N_noxref_23_c_3083_n N_noxref_24_c_3144_n ) capacitor c=0.01197f \
 //x=25.16 //y=2.08 //x2=25.525 //y2=1.59
cc_1634 ( N_noxref_23_c_3087_n N_noxref_24_c_3144_n ) capacitor c=0.00703864f \
 //x=24.86 //y=1.53 //x2=25.525 //y2=1.59
cc_1635 ( N_noxref_23_c_3088_n N_noxref_24_c_3144_n ) capacitor c=0.0224186f \
 //x=24.86 //y=1.915 //x2=25.525 //y2=1.59
cc_1636 ( N_noxref_23_c_3090_n N_noxref_24_c_3144_n ) capacitor c=0.00708583f \
 //x=25.235 //y=1.375 //x2=25.525 //y2=1.59
cc_1637 ( N_noxref_23_c_3093_n N_noxref_24_c_3144_n ) capacitor c=0.00698822f \
 //x=25.39 //y=1.22 //x2=25.525 //y2=1.59
cc_1638 ( N_noxref_23_c_3084_n N_noxref_24_M15_noxref_s ) capacitor \
 c=0.0327271f //x=24.86 //y=0.875 //x2=24.505 //y2=0.375
cc_1639 ( N_noxref_23_c_3087_n N_noxref_24_M15_noxref_s ) capacitor \
 c=7.99997e-19 //x=24.86 //y=1.53 //x2=24.505 //y2=0.375
cc_1640 ( N_noxref_23_c_3088_n N_noxref_24_M15_noxref_s ) capacitor \
 c=0.00122123f //x=24.86 //y=1.915 //x2=24.505 //y2=0.375
cc_1641 ( N_noxref_23_c_3091_n N_noxref_24_M15_noxref_s ) capacitor \
 c=0.0121427f //x=25.39 //y=0.875 //x2=24.505 //y2=0.375
cc_1642 ( N_noxref_23_M49_noxref_g N_noxref_25_c_3196_n ) capacitor \
 c=0.0186539f //x=25.8 //y=6.02 //x2=26.375 //y2=5.155
cc_1643 ( N_noxref_23_M48_noxref_g N_noxref_25_c_3200_n ) capacitor \
 c=0.0213876f //x=25.36 //y=6.02 //x2=25.665 //y2=5.155
cc_1644 ( N_noxref_23_c_3121_n N_noxref_25_c_3200_n ) capacitor c=0.0044314f \
 //x=25.725 //y=4.79 //x2=25.665 //y2=5.155
cc_1645 ( N_noxref_23_M49_noxref_g N_noxref_25_M48_noxref_d ) capacitor \
 c=0.0180032f //x=25.8 //y=6.02 //x2=25.435 //y2=5.02
cc_1646 ( N_noxref_24_M15_noxref_s N_noxref_25_M17_noxref_d ) capacitor \
 c=0.00309936f //x=24.505 //y=0.375 //x2=27.445 //y2=0.915
cc_1647 ( N_noxref_24_c_3151_n N_noxref_26_c_3271_n ) capacitor c=0.0134007f \
 //x=26.495 //y=0.54 //x2=27.065 //y2=0.995
cc_1648 ( N_noxref_24_c_3162_n N_noxref_26_c_3271_n ) capacitor c=0.0101391f \
 //x=26.495 //y=1.59 //x2=27.065 //y2=0.995
cc_1649 ( N_noxref_24_M15_noxref_s N_noxref_26_c_3271_n ) capacitor \
 c=0.0228195f //x=24.505 //y=0.375 //x2=27.065 //y2=0.995
cc_1650 ( N_noxref_24_M15_noxref_s N_noxref_26_c_3273_n ) capacitor \
 c=0.0180035f //x=24.505 //y=0.375 //x2=27.15 //y2=0.625
cc_1651 ( N_noxref_24_c_3151_n N_noxref_26_M16_noxref_d ) capacitor \
 c=0.0128561f //x=26.495 //y=0.54 //x2=25.91 //y2=0.91
cc_1652 ( N_noxref_24_c_3162_n N_noxref_26_M16_noxref_d ) capacitor \
 c=0.00891787f //x=26.495 //y=1.59 //x2=25.91 //y2=0.91
cc_1653 ( N_noxref_24_M15_noxref_s N_noxref_26_M16_noxref_d ) capacitor \
 c=0.0159202f //x=24.505 //y=0.375 //x2=25.91 //y2=0.91
cc_1654 ( N_noxref_24_M15_noxref_s N_noxref_26_M17_noxref_s ) capacitor \
 c=0.0213553f //x=24.505 //y=0.375 //x2=27.015 //y2=0.375
cc_1655 ( N_noxref_25_c_3194_n N_noxref_26_c_3276_n ) capacitor c=0.0046926f \
 //x=28.035 //y=1.665 //x2=28.035 //y2=0.54
cc_1656 ( N_noxref_25_M17_noxref_d N_noxref_26_c_3276_n ) capacitor \
 c=0.0118457f //x=27.445 //y=0.915 //x2=28.035 //y2=0.54
cc_1657 ( N_noxref_25_c_3267_p N_noxref_26_c_3301_n ) capacitor c=0.0200405f \
 //x=27.72 //y=1.665 //x2=27.15 //y2=0.995
cc_1658 ( N_noxref_25_M17_noxref_d N_noxref_26_M16_noxref_d ) capacitor \
 c=5.27807e-19 //x=27.445 //y=0.915 //x2=25.91 //y2=0.91
cc_1659 ( N_noxref_25_c_3194_n N_noxref_26_M17_noxref_s ) capacitor \
 c=0.0212001f //x=28.035 //y=1.665 //x2=27.015 //y2=0.375
cc_1660 ( N_noxref_25_M17_noxref_d N_noxref_26_M17_noxref_s ) capacitor \
 c=0.0426368f //x=27.445 //y=0.915 //x2=27.015 //y2=0.375
