magic
tech sky130A
magscale 1 2
timestamp 1669200987
<< nwell >>
rect -87 786 5859 1550
<< pwell >>
rect -34 -34 5806 544
<< nmos >>
rect 147 290 177 351
tri 177 290 193 306 sw
rect 447 290 477 351
rect 147 260 253 290
tri 253 260 283 290 sw
rect 147 159 177 260
tri 177 244 193 260 nw
tri 237 244 253 260 ne
tri 177 159 193 175 sw
tri 237 159 253 175 se
rect 253 159 283 260
tri 342 260 372 290 se
rect 372 260 477 290
rect 342 166 372 260
tri 372 244 388 260 nw
tri 431 244 447 260 ne
tri 372 166 388 182 sw
tri 431 166 447 182 se
rect 447 166 477 260
tri 147 129 177 159 ne
rect 177 129 253 159
tri 253 129 283 159 nw
tri 342 136 372 166 ne
rect 372 136 447 166
tri 447 136 477 166 nw
rect 649 298 679 351
tri 679 298 695 314 sw
rect 649 268 755 298
tri 755 268 785 298 sw
rect 649 167 679 268
tri 679 252 695 268 nw
tri 739 252 755 268 ne
tri 679 167 695 183 sw
tri 739 167 755 183 se
rect 755 167 785 268
tri 649 137 679 167 ne
rect 679 137 755 167
tri 755 137 785 167 nw
rect 1109 290 1139 351
tri 1139 290 1155 306 sw
rect 1409 290 1439 351
rect 1109 260 1215 290
tri 1215 260 1245 290 sw
rect 1109 159 1139 260
tri 1139 244 1155 260 nw
tri 1199 244 1215 260 ne
tri 1139 159 1155 175 sw
tri 1199 159 1215 175 se
rect 1215 159 1245 260
tri 1304 260 1334 290 se
rect 1334 260 1439 290
rect 1304 166 1334 260
tri 1334 244 1350 260 nw
tri 1393 244 1409 260 ne
tri 1334 166 1350 182 sw
tri 1393 166 1409 182 se
rect 1409 166 1439 260
tri 1109 129 1139 159 ne
rect 1139 129 1215 159
tri 1215 129 1245 159 nw
tri 1304 136 1334 166 ne
rect 1334 136 1409 166
tri 1409 136 1439 166 nw
rect 1611 298 1641 351
tri 1641 298 1657 314 sw
rect 1611 268 1717 298
tri 1717 268 1747 298 sw
rect 1611 167 1641 268
tri 1641 252 1657 268 nw
tri 1701 252 1717 268 ne
tri 1641 167 1657 183 sw
tri 1701 167 1717 183 se
rect 1717 167 1747 268
tri 1611 137 1641 167 ne
rect 1641 137 1717 167
tri 1717 137 1747 167 nw
rect 2071 290 2101 351
tri 2101 290 2117 306 sw
rect 2371 290 2401 351
rect 2071 260 2177 290
tri 2177 260 2207 290 sw
rect 2071 159 2101 260
tri 2101 244 2117 260 nw
tri 2161 244 2177 260 ne
tri 2101 159 2117 175 sw
tri 2161 159 2177 175 se
rect 2177 159 2207 260
tri 2266 260 2296 290 se
rect 2296 260 2401 290
rect 2266 166 2296 260
tri 2296 244 2312 260 nw
tri 2355 244 2371 260 ne
tri 2296 166 2312 182 sw
tri 2355 166 2371 182 se
rect 2371 166 2401 260
tri 2071 129 2101 159 ne
rect 2101 129 2177 159
tri 2177 129 2207 159 nw
tri 2266 136 2296 166 ne
rect 2296 136 2371 166
tri 2371 136 2401 166 nw
rect 2573 298 2603 351
tri 2603 298 2619 314 sw
rect 2573 268 2679 298
tri 2679 268 2709 298 sw
rect 2573 167 2603 268
tri 2603 252 2619 268 nw
tri 2663 252 2679 268 ne
tri 2603 167 2619 183 sw
tri 2663 167 2679 183 se
rect 2679 167 2709 268
tri 2573 137 2603 167 ne
rect 2603 137 2679 167
tri 2679 137 2709 167 nw
rect 3033 290 3063 351
tri 3063 290 3079 306 sw
rect 3333 290 3363 351
rect 3033 260 3139 290
tri 3139 260 3169 290 sw
rect 3033 159 3063 260
tri 3063 244 3079 260 nw
tri 3123 244 3139 260 ne
tri 3063 159 3079 175 sw
tri 3123 159 3139 175 se
rect 3139 159 3169 260
tri 3228 260 3258 290 se
rect 3258 260 3363 290
rect 3228 166 3258 260
tri 3258 244 3274 260 nw
tri 3317 244 3333 260 ne
tri 3258 166 3274 182 sw
tri 3317 166 3333 182 se
rect 3333 166 3363 260
tri 3033 129 3063 159 ne
rect 3063 129 3139 159
tri 3139 129 3169 159 nw
tri 3228 136 3258 166 ne
rect 3258 136 3333 166
tri 3333 136 3363 166 nw
rect 3535 298 3565 351
tri 3565 298 3581 314 sw
rect 3535 268 3641 298
tri 3641 268 3671 298 sw
rect 3535 167 3565 268
tri 3565 252 3581 268 nw
tri 3625 252 3641 268 ne
tri 3565 167 3581 183 sw
tri 3625 167 3641 183 se
rect 3641 167 3671 268
tri 3535 137 3565 167 ne
rect 3565 137 3641 167
tri 3641 137 3671 167 nw
rect 3995 290 4025 351
tri 4025 290 4041 306 sw
rect 4295 290 4325 351
rect 3995 260 4101 290
tri 4101 260 4131 290 sw
rect 3995 159 4025 260
tri 4025 244 4041 260 nw
tri 4085 244 4101 260 ne
tri 4025 159 4041 175 sw
tri 4085 159 4101 175 se
rect 4101 159 4131 260
tri 4190 260 4220 290 se
rect 4220 260 4325 290
rect 4190 166 4220 260
tri 4220 244 4236 260 nw
tri 4279 244 4295 260 ne
tri 4220 166 4236 182 sw
tri 4279 166 4295 182 se
rect 4295 166 4325 260
tri 3995 129 4025 159 ne
rect 4025 129 4101 159
tri 4101 129 4131 159 nw
tri 4190 136 4220 166 ne
rect 4220 136 4295 166
tri 4295 136 4325 166 nw
rect 4497 298 4527 351
tri 4527 298 4543 314 sw
rect 4497 268 4603 298
tri 4603 268 4633 298 sw
rect 4497 167 4527 268
tri 4527 252 4543 268 nw
tri 4587 252 4603 268 ne
tri 4527 167 4543 183 sw
tri 4587 167 4603 183 se
rect 4603 167 4633 268
tri 4497 137 4527 167 ne
rect 4527 137 4603 167
tri 4603 137 4633 167 nw
rect 4957 290 4987 351
tri 4987 290 5003 306 sw
rect 5257 290 5287 351
rect 4957 260 5063 290
tri 5063 260 5093 290 sw
rect 4957 159 4987 260
tri 4987 244 5003 260 nw
tri 5047 244 5063 260 ne
tri 4987 159 5003 175 sw
tri 5047 159 5063 175 se
rect 5063 159 5093 260
tri 5152 260 5182 290 se
rect 5182 260 5287 290
rect 5152 166 5182 260
tri 5182 244 5198 260 nw
tri 5241 244 5257 260 ne
tri 5182 166 5198 182 sw
tri 5241 166 5257 182 se
rect 5257 166 5287 260
tri 4957 129 4987 159 ne
rect 4987 129 5063 159
tri 5063 129 5093 159 nw
tri 5152 136 5182 166 ne
rect 5182 136 5257 166
tri 5257 136 5287 166 nw
rect 5459 298 5489 351
tri 5489 298 5505 314 sw
rect 5459 268 5565 298
tri 5565 268 5595 298 sw
rect 5459 167 5489 268
tri 5489 252 5505 268 nw
tri 5549 252 5565 268 ne
tri 5489 167 5505 183 sw
tri 5549 167 5565 183 se
rect 5565 167 5595 268
tri 5459 137 5489 167 ne
rect 5489 137 5565 167
tri 5565 137 5595 167 nw
<< pmos >>
rect 247 1004 277 1404
rect 335 1004 365 1404
rect 423 1004 453 1404
rect 511 1004 541 1404
rect 599 1004 629 1404
rect 687 1004 717 1404
rect 1209 1004 1239 1404
rect 1297 1004 1327 1404
rect 1385 1004 1415 1404
rect 1473 1004 1503 1404
rect 1561 1004 1591 1404
rect 1649 1004 1679 1404
rect 2171 1004 2201 1404
rect 2259 1004 2289 1404
rect 2347 1004 2377 1404
rect 2435 1004 2465 1404
rect 2523 1004 2553 1404
rect 2611 1004 2641 1404
rect 3133 1004 3163 1404
rect 3221 1004 3251 1404
rect 3309 1004 3339 1404
rect 3397 1004 3427 1404
rect 3485 1004 3515 1404
rect 3573 1004 3603 1404
rect 4095 1004 4125 1404
rect 4183 1004 4213 1404
rect 4271 1004 4301 1404
rect 4359 1004 4389 1404
rect 4447 1004 4477 1404
rect 4535 1004 4565 1404
rect 5057 1004 5087 1404
rect 5145 1004 5175 1404
rect 5233 1004 5263 1404
rect 5321 1004 5351 1404
rect 5409 1004 5439 1404
rect 5497 1004 5527 1404
<< ndiff >>
rect 91 335 147 351
rect 91 301 101 335
rect 135 301 147 335
rect 91 263 147 301
rect 177 335 447 351
rect 177 306 198 335
tri 177 290 193 306 ne
rect 193 301 198 306
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 447 335
rect 193 290 447 301
rect 477 335 533 351
rect 477 301 489 335
rect 523 301 533 335
rect 91 229 101 263
rect 135 229 147 263
tri 253 260 283 290 ne
rect 283 263 342 290
rect 91 195 147 229
rect 91 161 101 195
rect 135 161 147 195
rect 91 129 147 161
tri 177 244 193 260 se
rect 193 244 237 260
tri 237 244 253 260 sw
rect 177 210 253 244
rect 177 176 198 210
rect 232 176 253 210
rect 177 175 253 176
tri 177 159 193 175 ne
rect 193 159 237 175
tri 237 159 253 175 nw
rect 283 229 295 263
rect 329 229 342 263
tri 342 260 372 290 nw
rect 283 195 342 229
rect 283 161 295 195
rect 329 161 342 195
tri 372 244 388 260 se
rect 388 244 431 260
tri 431 244 447 260 sw
rect 372 216 447 244
rect 372 182 393 216
rect 427 182 447 216
tri 372 166 388 182 ne
rect 388 166 431 182
tri 431 166 447 182 nw
tri 147 129 177 159 sw
tri 253 129 283 159 se
rect 283 136 342 161
tri 342 136 372 166 sw
tri 447 136 477 166 se
rect 477 136 533 301
rect 283 129 533 136
rect 91 125 533 129
rect 91 91 101 125
rect 135 91 295 125
rect 329 91 392 125
rect 426 91 489 125
rect 523 91 533 125
rect 91 75 533 91
rect 593 335 649 351
rect 593 301 603 335
rect 637 301 649 335
rect 593 263 649 301
rect 679 314 841 351
tri 679 298 695 314 ne
rect 695 298 841 314
tri 755 268 785 298 ne
rect 593 229 603 263
rect 637 229 649 263
rect 593 195 649 229
rect 593 161 603 195
rect 637 161 649 195
tri 679 252 695 268 se
rect 695 252 739 268
tri 739 252 755 268 sw
rect 679 219 755 252
rect 679 185 700 219
rect 734 185 755 219
rect 679 183 755 185
tri 679 167 695 183 ne
rect 695 167 739 183
tri 739 167 755 183 nw
rect 785 263 841 298
rect 785 229 797 263
rect 831 229 841 263
rect 785 195 841 229
rect 593 137 649 161
tri 649 137 679 167 sw
tri 755 137 785 167 se
rect 785 161 797 195
rect 831 161 841 195
rect 785 137 841 161
rect 593 125 841 137
rect 593 91 603 125
rect 637 91 700 125
rect 734 91 797 125
rect 831 91 841 125
rect 593 75 841 91
rect 1053 335 1109 351
rect 1053 301 1063 335
rect 1097 301 1109 335
rect 1053 263 1109 301
rect 1139 335 1409 351
rect 1139 306 1160 335
tri 1139 290 1155 306 ne
rect 1155 301 1160 306
rect 1194 301 1257 335
rect 1291 301 1354 335
rect 1388 301 1409 335
rect 1155 290 1409 301
rect 1439 335 1495 351
rect 1439 301 1451 335
rect 1485 301 1495 335
rect 1053 229 1063 263
rect 1097 229 1109 263
tri 1215 260 1245 290 ne
rect 1245 263 1304 290
rect 1053 195 1109 229
rect 1053 161 1063 195
rect 1097 161 1109 195
rect 1053 129 1109 161
tri 1139 244 1155 260 se
rect 1155 244 1199 260
tri 1199 244 1215 260 sw
rect 1139 210 1215 244
rect 1139 176 1160 210
rect 1194 176 1215 210
rect 1139 175 1215 176
tri 1139 159 1155 175 ne
rect 1155 159 1199 175
tri 1199 159 1215 175 nw
rect 1245 229 1257 263
rect 1291 229 1304 263
tri 1304 260 1334 290 nw
rect 1245 195 1304 229
rect 1245 161 1257 195
rect 1291 161 1304 195
tri 1334 244 1350 260 se
rect 1350 244 1393 260
tri 1393 244 1409 260 sw
rect 1334 216 1409 244
rect 1334 182 1355 216
rect 1389 182 1409 216
tri 1334 166 1350 182 ne
rect 1350 166 1393 182
tri 1393 166 1409 182 nw
tri 1109 129 1139 159 sw
tri 1215 129 1245 159 se
rect 1245 136 1304 161
tri 1304 136 1334 166 sw
tri 1409 136 1439 166 se
rect 1439 136 1495 301
rect 1245 129 1495 136
rect 1053 125 1495 129
rect 1053 91 1063 125
rect 1097 91 1257 125
rect 1291 91 1354 125
rect 1388 91 1451 125
rect 1485 91 1495 125
rect 1053 75 1495 91
rect 1555 335 1611 351
rect 1555 301 1565 335
rect 1599 301 1611 335
rect 1555 263 1611 301
rect 1641 314 1803 351
tri 1641 298 1657 314 ne
rect 1657 298 1803 314
tri 1717 268 1747 298 ne
rect 1555 229 1565 263
rect 1599 229 1611 263
rect 1555 195 1611 229
rect 1555 161 1565 195
rect 1599 161 1611 195
tri 1641 252 1657 268 se
rect 1657 252 1701 268
tri 1701 252 1717 268 sw
rect 1641 219 1717 252
rect 1641 185 1662 219
rect 1696 185 1717 219
rect 1641 183 1717 185
tri 1641 167 1657 183 ne
rect 1657 167 1701 183
tri 1701 167 1717 183 nw
rect 1747 263 1803 298
rect 1747 229 1759 263
rect 1793 229 1803 263
rect 1747 195 1803 229
rect 1555 137 1611 161
tri 1611 137 1641 167 sw
tri 1717 137 1747 167 se
rect 1747 161 1759 195
rect 1793 161 1803 195
rect 1747 137 1803 161
rect 1555 125 1803 137
rect 1555 91 1565 125
rect 1599 91 1662 125
rect 1696 91 1759 125
rect 1793 91 1803 125
rect 1555 75 1803 91
rect 2015 335 2071 351
rect 2015 301 2025 335
rect 2059 301 2071 335
rect 2015 263 2071 301
rect 2101 335 2371 351
rect 2101 306 2122 335
tri 2101 290 2117 306 ne
rect 2117 301 2122 306
rect 2156 301 2219 335
rect 2253 301 2316 335
rect 2350 301 2371 335
rect 2117 290 2371 301
rect 2401 335 2457 351
rect 2401 301 2413 335
rect 2447 301 2457 335
rect 2015 229 2025 263
rect 2059 229 2071 263
tri 2177 260 2207 290 ne
rect 2207 263 2266 290
rect 2015 195 2071 229
rect 2015 161 2025 195
rect 2059 161 2071 195
rect 2015 129 2071 161
tri 2101 244 2117 260 se
rect 2117 244 2161 260
tri 2161 244 2177 260 sw
rect 2101 210 2177 244
rect 2101 176 2122 210
rect 2156 176 2177 210
rect 2101 175 2177 176
tri 2101 159 2117 175 ne
rect 2117 159 2161 175
tri 2161 159 2177 175 nw
rect 2207 229 2219 263
rect 2253 229 2266 263
tri 2266 260 2296 290 nw
rect 2207 195 2266 229
rect 2207 161 2219 195
rect 2253 161 2266 195
tri 2296 244 2312 260 se
rect 2312 244 2355 260
tri 2355 244 2371 260 sw
rect 2296 216 2371 244
rect 2296 182 2317 216
rect 2351 182 2371 216
tri 2296 166 2312 182 ne
rect 2312 166 2355 182
tri 2355 166 2371 182 nw
tri 2071 129 2101 159 sw
tri 2177 129 2207 159 se
rect 2207 136 2266 161
tri 2266 136 2296 166 sw
tri 2371 136 2401 166 se
rect 2401 136 2457 301
rect 2207 129 2457 136
rect 2015 125 2457 129
rect 2015 91 2025 125
rect 2059 91 2219 125
rect 2253 91 2316 125
rect 2350 91 2413 125
rect 2447 91 2457 125
rect 2015 75 2457 91
rect 2517 335 2573 351
rect 2517 301 2527 335
rect 2561 301 2573 335
rect 2517 263 2573 301
rect 2603 314 2765 351
tri 2603 298 2619 314 ne
rect 2619 298 2765 314
tri 2679 268 2709 298 ne
rect 2517 229 2527 263
rect 2561 229 2573 263
rect 2517 195 2573 229
rect 2517 161 2527 195
rect 2561 161 2573 195
tri 2603 252 2619 268 se
rect 2619 252 2663 268
tri 2663 252 2679 268 sw
rect 2603 219 2679 252
rect 2603 185 2624 219
rect 2658 185 2679 219
rect 2603 183 2679 185
tri 2603 167 2619 183 ne
rect 2619 167 2663 183
tri 2663 167 2679 183 nw
rect 2709 263 2765 298
rect 2709 229 2721 263
rect 2755 229 2765 263
rect 2709 195 2765 229
rect 2517 137 2573 161
tri 2573 137 2603 167 sw
tri 2679 137 2709 167 se
rect 2709 161 2721 195
rect 2755 161 2765 195
rect 2709 137 2765 161
rect 2517 125 2765 137
rect 2517 91 2527 125
rect 2561 91 2624 125
rect 2658 91 2721 125
rect 2755 91 2765 125
rect 2517 75 2765 91
rect 2977 335 3033 351
rect 2977 301 2987 335
rect 3021 301 3033 335
rect 2977 263 3033 301
rect 3063 335 3333 351
rect 3063 306 3084 335
tri 3063 290 3079 306 ne
rect 3079 301 3084 306
rect 3118 301 3181 335
rect 3215 301 3278 335
rect 3312 301 3333 335
rect 3079 290 3333 301
rect 3363 335 3419 351
rect 3363 301 3375 335
rect 3409 301 3419 335
rect 2977 229 2987 263
rect 3021 229 3033 263
tri 3139 260 3169 290 ne
rect 3169 263 3228 290
rect 2977 195 3033 229
rect 2977 161 2987 195
rect 3021 161 3033 195
rect 2977 129 3033 161
tri 3063 244 3079 260 se
rect 3079 244 3123 260
tri 3123 244 3139 260 sw
rect 3063 210 3139 244
rect 3063 176 3084 210
rect 3118 176 3139 210
rect 3063 175 3139 176
tri 3063 159 3079 175 ne
rect 3079 159 3123 175
tri 3123 159 3139 175 nw
rect 3169 229 3181 263
rect 3215 229 3228 263
tri 3228 260 3258 290 nw
rect 3169 195 3228 229
rect 3169 161 3181 195
rect 3215 161 3228 195
tri 3258 244 3274 260 se
rect 3274 244 3317 260
tri 3317 244 3333 260 sw
rect 3258 216 3333 244
rect 3258 182 3279 216
rect 3313 182 3333 216
tri 3258 166 3274 182 ne
rect 3274 166 3317 182
tri 3317 166 3333 182 nw
tri 3033 129 3063 159 sw
tri 3139 129 3169 159 se
rect 3169 136 3228 161
tri 3228 136 3258 166 sw
tri 3333 136 3363 166 se
rect 3363 136 3419 301
rect 3169 129 3419 136
rect 2977 125 3419 129
rect 2977 91 2987 125
rect 3021 91 3181 125
rect 3215 91 3278 125
rect 3312 91 3375 125
rect 3409 91 3419 125
rect 2977 75 3419 91
rect 3479 335 3535 351
rect 3479 301 3489 335
rect 3523 301 3535 335
rect 3479 263 3535 301
rect 3565 314 3727 351
tri 3565 298 3581 314 ne
rect 3581 298 3727 314
tri 3641 268 3671 298 ne
rect 3479 229 3489 263
rect 3523 229 3535 263
rect 3479 195 3535 229
rect 3479 161 3489 195
rect 3523 161 3535 195
tri 3565 252 3581 268 se
rect 3581 252 3625 268
tri 3625 252 3641 268 sw
rect 3565 219 3641 252
rect 3565 185 3586 219
rect 3620 185 3641 219
rect 3565 183 3641 185
tri 3565 167 3581 183 ne
rect 3581 167 3625 183
tri 3625 167 3641 183 nw
rect 3671 263 3727 298
rect 3671 229 3683 263
rect 3717 229 3727 263
rect 3671 195 3727 229
rect 3479 137 3535 161
tri 3535 137 3565 167 sw
tri 3641 137 3671 167 se
rect 3671 161 3683 195
rect 3717 161 3727 195
rect 3671 137 3727 161
rect 3479 125 3727 137
rect 3479 91 3489 125
rect 3523 91 3586 125
rect 3620 91 3683 125
rect 3717 91 3727 125
rect 3479 75 3727 91
rect 3939 335 3995 351
rect 3939 301 3949 335
rect 3983 301 3995 335
rect 3939 263 3995 301
rect 4025 335 4295 351
rect 4025 306 4046 335
tri 4025 290 4041 306 ne
rect 4041 301 4046 306
rect 4080 301 4143 335
rect 4177 301 4240 335
rect 4274 301 4295 335
rect 4041 290 4295 301
rect 4325 335 4381 351
rect 4325 301 4337 335
rect 4371 301 4381 335
rect 3939 229 3949 263
rect 3983 229 3995 263
tri 4101 260 4131 290 ne
rect 4131 263 4190 290
rect 3939 195 3995 229
rect 3939 161 3949 195
rect 3983 161 3995 195
rect 3939 129 3995 161
tri 4025 244 4041 260 se
rect 4041 244 4085 260
tri 4085 244 4101 260 sw
rect 4025 210 4101 244
rect 4025 176 4046 210
rect 4080 176 4101 210
rect 4025 175 4101 176
tri 4025 159 4041 175 ne
rect 4041 159 4085 175
tri 4085 159 4101 175 nw
rect 4131 229 4143 263
rect 4177 229 4190 263
tri 4190 260 4220 290 nw
rect 4131 195 4190 229
rect 4131 161 4143 195
rect 4177 161 4190 195
tri 4220 244 4236 260 se
rect 4236 244 4279 260
tri 4279 244 4295 260 sw
rect 4220 216 4295 244
rect 4220 182 4241 216
rect 4275 182 4295 216
tri 4220 166 4236 182 ne
rect 4236 166 4279 182
tri 4279 166 4295 182 nw
tri 3995 129 4025 159 sw
tri 4101 129 4131 159 se
rect 4131 136 4190 161
tri 4190 136 4220 166 sw
tri 4295 136 4325 166 se
rect 4325 136 4381 301
rect 4131 129 4381 136
rect 3939 125 4381 129
rect 3939 91 3949 125
rect 3983 91 4143 125
rect 4177 91 4240 125
rect 4274 91 4337 125
rect 4371 91 4381 125
rect 3939 75 4381 91
rect 4441 335 4497 351
rect 4441 301 4451 335
rect 4485 301 4497 335
rect 4441 263 4497 301
rect 4527 314 4689 351
tri 4527 298 4543 314 ne
rect 4543 298 4689 314
tri 4603 268 4633 298 ne
rect 4441 229 4451 263
rect 4485 229 4497 263
rect 4441 195 4497 229
rect 4441 161 4451 195
rect 4485 161 4497 195
tri 4527 252 4543 268 se
rect 4543 252 4587 268
tri 4587 252 4603 268 sw
rect 4527 219 4603 252
rect 4527 185 4548 219
rect 4582 185 4603 219
rect 4527 183 4603 185
tri 4527 167 4543 183 ne
rect 4543 167 4587 183
tri 4587 167 4603 183 nw
rect 4633 263 4689 298
rect 4633 229 4645 263
rect 4679 229 4689 263
rect 4633 195 4689 229
rect 4441 137 4497 161
tri 4497 137 4527 167 sw
tri 4603 137 4633 167 se
rect 4633 161 4645 195
rect 4679 161 4689 195
rect 4633 137 4689 161
rect 4441 125 4689 137
rect 4441 91 4451 125
rect 4485 91 4548 125
rect 4582 91 4645 125
rect 4679 91 4689 125
rect 4441 75 4689 91
rect 4901 335 4957 351
rect 4901 301 4911 335
rect 4945 301 4957 335
rect 4901 263 4957 301
rect 4987 335 5257 351
rect 4987 306 5008 335
tri 4987 290 5003 306 ne
rect 5003 301 5008 306
rect 5042 301 5105 335
rect 5139 301 5202 335
rect 5236 301 5257 335
rect 5003 290 5257 301
rect 5287 335 5343 351
rect 5287 301 5299 335
rect 5333 301 5343 335
rect 4901 229 4911 263
rect 4945 229 4957 263
tri 5063 260 5093 290 ne
rect 5093 263 5152 290
rect 4901 195 4957 229
rect 4901 161 4911 195
rect 4945 161 4957 195
rect 4901 129 4957 161
tri 4987 244 5003 260 se
rect 5003 244 5047 260
tri 5047 244 5063 260 sw
rect 4987 210 5063 244
rect 4987 176 5008 210
rect 5042 176 5063 210
rect 4987 175 5063 176
tri 4987 159 5003 175 ne
rect 5003 159 5047 175
tri 5047 159 5063 175 nw
rect 5093 229 5105 263
rect 5139 229 5152 263
tri 5152 260 5182 290 nw
rect 5093 195 5152 229
rect 5093 161 5105 195
rect 5139 161 5152 195
tri 5182 244 5198 260 se
rect 5198 244 5241 260
tri 5241 244 5257 260 sw
rect 5182 216 5257 244
rect 5182 182 5203 216
rect 5237 182 5257 216
tri 5182 166 5198 182 ne
rect 5198 166 5241 182
tri 5241 166 5257 182 nw
tri 4957 129 4987 159 sw
tri 5063 129 5093 159 se
rect 5093 136 5152 161
tri 5152 136 5182 166 sw
tri 5257 136 5287 166 se
rect 5287 136 5343 301
rect 5093 129 5343 136
rect 4901 125 5343 129
rect 4901 91 4911 125
rect 4945 91 5105 125
rect 5139 91 5202 125
rect 5236 91 5299 125
rect 5333 91 5343 125
rect 4901 75 5343 91
rect 5403 335 5459 351
rect 5403 301 5413 335
rect 5447 301 5459 335
rect 5403 263 5459 301
rect 5489 314 5651 351
tri 5489 298 5505 314 ne
rect 5505 298 5651 314
tri 5565 268 5595 298 ne
rect 5403 229 5413 263
rect 5447 229 5459 263
rect 5403 195 5459 229
rect 5403 161 5413 195
rect 5447 161 5459 195
tri 5489 252 5505 268 se
rect 5505 252 5549 268
tri 5549 252 5565 268 sw
rect 5489 219 5565 252
rect 5489 185 5510 219
rect 5544 185 5565 219
rect 5489 183 5565 185
tri 5489 167 5505 183 ne
rect 5505 167 5549 183
tri 5549 167 5565 183 nw
rect 5595 263 5651 298
rect 5595 229 5607 263
rect 5641 229 5651 263
rect 5595 195 5651 229
rect 5403 137 5459 161
tri 5459 137 5489 167 sw
tri 5565 137 5595 167 se
rect 5595 161 5607 195
rect 5641 161 5651 195
rect 5595 137 5651 161
rect 5403 125 5651 137
rect 5403 91 5413 125
rect 5447 91 5510 125
rect 5544 91 5607 125
rect 5641 91 5651 125
rect 5403 75 5651 91
<< pdiff >>
rect 191 1366 247 1404
rect 191 1332 201 1366
rect 235 1332 247 1366
rect 191 1298 247 1332
rect 191 1264 201 1298
rect 235 1264 247 1298
rect 191 1230 247 1264
rect 191 1196 201 1230
rect 235 1196 247 1230
rect 191 1162 247 1196
rect 191 1128 201 1162
rect 235 1128 247 1162
rect 191 1093 247 1128
rect 191 1059 201 1093
rect 235 1059 247 1093
rect 191 1004 247 1059
rect 277 1366 335 1404
rect 277 1332 289 1366
rect 323 1332 335 1366
rect 277 1298 335 1332
rect 277 1264 289 1298
rect 323 1264 335 1298
rect 277 1230 335 1264
rect 277 1196 289 1230
rect 323 1196 335 1230
rect 277 1162 335 1196
rect 277 1128 289 1162
rect 323 1128 335 1162
rect 277 1093 335 1128
rect 277 1059 289 1093
rect 323 1059 335 1093
rect 277 1004 335 1059
rect 365 1366 423 1404
rect 365 1332 377 1366
rect 411 1332 423 1366
rect 365 1298 423 1332
rect 365 1264 377 1298
rect 411 1264 423 1298
rect 365 1230 423 1264
rect 365 1196 377 1230
rect 411 1196 423 1230
rect 365 1162 423 1196
rect 365 1128 377 1162
rect 411 1128 423 1162
rect 365 1004 423 1128
rect 453 1366 511 1404
rect 453 1332 465 1366
rect 499 1332 511 1366
rect 453 1298 511 1332
rect 453 1264 465 1298
rect 499 1264 511 1298
rect 453 1230 511 1264
rect 453 1196 465 1230
rect 499 1196 511 1230
rect 453 1162 511 1196
rect 453 1128 465 1162
rect 499 1128 511 1162
rect 453 1093 511 1128
rect 453 1059 465 1093
rect 499 1059 511 1093
rect 453 1004 511 1059
rect 541 1366 599 1404
rect 541 1332 553 1366
rect 587 1332 599 1366
rect 541 1298 599 1332
rect 541 1264 553 1298
rect 587 1264 599 1298
rect 541 1230 599 1264
rect 541 1196 553 1230
rect 587 1196 599 1230
rect 541 1162 599 1196
rect 541 1128 553 1162
rect 587 1128 599 1162
rect 541 1004 599 1128
rect 629 1366 687 1404
rect 629 1332 641 1366
rect 675 1332 687 1366
rect 629 1298 687 1332
rect 629 1264 641 1298
rect 675 1264 687 1298
rect 629 1230 687 1264
rect 629 1196 641 1230
rect 675 1196 687 1230
rect 629 1162 687 1196
rect 629 1128 641 1162
rect 675 1128 687 1162
rect 629 1093 687 1128
rect 629 1059 641 1093
rect 675 1059 687 1093
rect 629 1004 687 1059
rect 717 1366 771 1404
rect 717 1332 729 1366
rect 763 1332 771 1366
rect 717 1298 771 1332
rect 717 1264 729 1298
rect 763 1264 771 1298
rect 717 1230 771 1264
rect 717 1196 729 1230
rect 763 1196 771 1230
rect 717 1162 771 1196
rect 717 1128 729 1162
rect 763 1128 771 1162
rect 717 1004 771 1128
rect 1153 1366 1209 1404
rect 1153 1332 1163 1366
rect 1197 1332 1209 1366
rect 1153 1298 1209 1332
rect 1153 1264 1163 1298
rect 1197 1264 1209 1298
rect 1153 1230 1209 1264
rect 1153 1196 1163 1230
rect 1197 1196 1209 1230
rect 1153 1162 1209 1196
rect 1153 1128 1163 1162
rect 1197 1128 1209 1162
rect 1153 1093 1209 1128
rect 1153 1059 1163 1093
rect 1197 1059 1209 1093
rect 1153 1004 1209 1059
rect 1239 1366 1297 1404
rect 1239 1332 1251 1366
rect 1285 1332 1297 1366
rect 1239 1298 1297 1332
rect 1239 1264 1251 1298
rect 1285 1264 1297 1298
rect 1239 1230 1297 1264
rect 1239 1196 1251 1230
rect 1285 1196 1297 1230
rect 1239 1162 1297 1196
rect 1239 1128 1251 1162
rect 1285 1128 1297 1162
rect 1239 1093 1297 1128
rect 1239 1059 1251 1093
rect 1285 1059 1297 1093
rect 1239 1004 1297 1059
rect 1327 1366 1385 1404
rect 1327 1332 1339 1366
rect 1373 1332 1385 1366
rect 1327 1298 1385 1332
rect 1327 1264 1339 1298
rect 1373 1264 1385 1298
rect 1327 1230 1385 1264
rect 1327 1196 1339 1230
rect 1373 1196 1385 1230
rect 1327 1162 1385 1196
rect 1327 1128 1339 1162
rect 1373 1128 1385 1162
rect 1327 1004 1385 1128
rect 1415 1366 1473 1404
rect 1415 1332 1427 1366
rect 1461 1332 1473 1366
rect 1415 1298 1473 1332
rect 1415 1264 1427 1298
rect 1461 1264 1473 1298
rect 1415 1230 1473 1264
rect 1415 1196 1427 1230
rect 1461 1196 1473 1230
rect 1415 1162 1473 1196
rect 1415 1128 1427 1162
rect 1461 1128 1473 1162
rect 1415 1093 1473 1128
rect 1415 1059 1427 1093
rect 1461 1059 1473 1093
rect 1415 1004 1473 1059
rect 1503 1366 1561 1404
rect 1503 1332 1515 1366
rect 1549 1332 1561 1366
rect 1503 1298 1561 1332
rect 1503 1264 1515 1298
rect 1549 1264 1561 1298
rect 1503 1230 1561 1264
rect 1503 1196 1515 1230
rect 1549 1196 1561 1230
rect 1503 1162 1561 1196
rect 1503 1128 1515 1162
rect 1549 1128 1561 1162
rect 1503 1004 1561 1128
rect 1591 1366 1649 1404
rect 1591 1332 1603 1366
rect 1637 1332 1649 1366
rect 1591 1298 1649 1332
rect 1591 1264 1603 1298
rect 1637 1264 1649 1298
rect 1591 1230 1649 1264
rect 1591 1196 1603 1230
rect 1637 1196 1649 1230
rect 1591 1162 1649 1196
rect 1591 1128 1603 1162
rect 1637 1128 1649 1162
rect 1591 1093 1649 1128
rect 1591 1059 1603 1093
rect 1637 1059 1649 1093
rect 1591 1004 1649 1059
rect 1679 1366 1733 1404
rect 1679 1332 1691 1366
rect 1725 1332 1733 1366
rect 1679 1298 1733 1332
rect 1679 1264 1691 1298
rect 1725 1264 1733 1298
rect 1679 1230 1733 1264
rect 1679 1196 1691 1230
rect 1725 1196 1733 1230
rect 1679 1162 1733 1196
rect 1679 1128 1691 1162
rect 1725 1128 1733 1162
rect 1679 1004 1733 1128
rect 2115 1366 2171 1404
rect 2115 1332 2125 1366
rect 2159 1332 2171 1366
rect 2115 1298 2171 1332
rect 2115 1264 2125 1298
rect 2159 1264 2171 1298
rect 2115 1230 2171 1264
rect 2115 1196 2125 1230
rect 2159 1196 2171 1230
rect 2115 1162 2171 1196
rect 2115 1128 2125 1162
rect 2159 1128 2171 1162
rect 2115 1093 2171 1128
rect 2115 1059 2125 1093
rect 2159 1059 2171 1093
rect 2115 1004 2171 1059
rect 2201 1366 2259 1404
rect 2201 1332 2213 1366
rect 2247 1332 2259 1366
rect 2201 1298 2259 1332
rect 2201 1264 2213 1298
rect 2247 1264 2259 1298
rect 2201 1230 2259 1264
rect 2201 1196 2213 1230
rect 2247 1196 2259 1230
rect 2201 1162 2259 1196
rect 2201 1128 2213 1162
rect 2247 1128 2259 1162
rect 2201 1093 2259 1128
rect 2201 1059 2213 1093
rect 2247 1059 2259 1093
rect 2201 1004 2259 1059
rect 2289 1366 2347 1404
rect 2289 1332 2301 1366
rect 2335 1332 2347 1366
rect 2289 1298 2347 1332
rect 2289 1264 2301 1298
rect 2335 1264 2347 1298
rect 2289 1230 2347 1264
rect 2289 1196 2301 1230
rect 2335 1196 2347 1230
rect 2289 1162 2347 1196
rect 2289 1128 2301 1162
rect 2335 1128 2347 1162
rect 2289 1004 2347 1128
rect 2377 1366 2435 1404
rect 2377 1332 2389 1366
rect 2423 1332 2435 1366
rect 2377 1298 2435 1332
rect 2377 1264 2389 1298
rect 2423 1264 2435 1298
rect 2377 1230 2435 1264
rect 2377 1196 2389 1230
rect 2423 1196 2435 1230
rect 2377 1162 2435 1196
rect 2377 1128 2389 1162
rect 2423 1128 2435 1162
rect 2377 1093 2435 1128
rect 2377 1059 2389 1093
rect 2423 1059 2435 1093
rect 2377 1004 2435 1059
rect 2465 1366 2523 1404
rect 2465 1332 2477 1366
rect 2511 1332 2523 1366
rect 2465 1298 2523 1332
rect 2465 1264 2477 1298
rect 2511 1264 2523 1298
rect 2465 1230 2523 1264
rect 2465 1196 2477 1230
rect 2511 1196 2523 1230
rect 2465 1162 2523 1196
rect 2465 1128 2477 1162
rect 2511 1128 2523 1162
rect 2465 1004 2523 1128
rect 2553 1366 2611 1404
rect 2553 1332 2565 1366
rect 2599 1332 2611 1366
rect 2553 1298 2611 1332
rect 2553 1264 2565 1298
rect 2599 1264 2611 1298
rect 2553 1230 2611 1264
rect 2553 1196 2565 1230
rect 2599 1196 2611 1230
rect 2553 1162 2611 1196
rect 2553 1128 2565 1162
rect 2599 1128 2611 1162
rect 2553 1093 2611 1128
rect 2553 1059 2565 1093
rect 2599 1059 2611 1093
rect 2553 1004 2611 1059
rect 2641 1366 2695 1404
rect 2641 1332 2653 1366
rect 2687 1332 2695 1366
rect 2641 1298 2695 1332
rect 2641 1264 2653 1298
rect 2687 1264 2695 1298
rect 2641 1230 2695 1264
rect 2641 1196 2653 1230
rect 2687 1196 2695 1230
rect 2641 1162 2695 1196
rect 2641 1128 2653 1162
rect 2687 1128 2695 1162
rect 2641 1004 2695 1128
rect 3077 1366 3133 1404
rect 3077 1332 3087 1366
rect 3121 1332 3133 1366
rect 3077 1298 3133 1332
rect 3077 1264 3087 1298
rect 3121 1264 3133 1298
rect 3077 1230 3133 1264
rect 3077 1196 3087 1230
rect 3121 1196 3133 1230
rect 3077 1162 3133 1196
rect 3077 1128 3087 1162
rect 3121 1128 3133 1162
rect 3077 1093 3133 1128
rect 3077 1059 3087 1093
rect 3121 1059 3133 1093
rect 3077 1004 3133 1059
rect 3163 1366 3221 1404
rect 3163 1332 3175 1366
rect 3209 1332 3221 1366
rect 3163 1298 3221 1332
rect 3163 1264 3175 1298
rect 3209 1264 3221 1298
rect 3163 1230 3221 1264
rect 3163 1196 3175 1230
rect 3209 1196 3221 1230
rect 3163 1162 3221 1196
rect 3163 1128 3175 1162
rect 3209 1128 3221 1162
rect 3163 1093 3221 1128
rect 3163 1059 3175 1093
rect 3209 1059 3221 1093
rect 3163 1004 3221 1059
rect 3251 1366 3309 1404
rect 3251 1332 3263 1366
rect 3297 1332 3309 1366
rect 3251 1298 3309 1332
rect 3251 1264 3263 1298
rect 3297 1264 3309 1298
rect 3251 1230 3309 1264
rect 3251 1196 3263 1230
rect 3297 1196 3309 1230
rect 3251 1162 3309 1196
rect 3251 1128 3263 1162
rect 3297 1128 3309 1162
rect 3251 1004 3309 1128
rect 3339 1366 3397 1404
rect 3339 1332 3351 1366
rect 3385 1332 3397 1366
rect 3339 1298 3397 1332
rect 3339 1264 3351 1298
rect 3385 1264 3397 1298
rect 3339 1230 3397 1264
rect 3339 1196 3351 1230
rect 3385 1196 3397 1230
rect 3339 1162 3397 1196
rect 3339 1128 3351 1162
rect 3385 1128 3397 1162
rect 3339 1093 3397 1128
rect 3339 1059 3351 1093
rect 3385 1059 3397 1093
rect 3339 1004 3397 1059
rect 3427 1366 3485 1404
rect 3427 1332 3439 1366
rect 3473 1332 3485 1366
rect 3427 1298 3485 1332
rect 3427 1264 3439 1298
rect 3473 1264 3485 1298
rect 3427 1230 3485 1264
rect 3427 1196 3439 1230
rect 3473 1196 3485 1230
rect 3427 1162 3485 1196
rect 3427 1128 3439 1162
rect 3473 1128 3485 1162
rect 3427 1004 3485 1128
rect 3515 1366 3573 1404
rect 3515 1332 3527 1366
rect 3561 1332 3573 1366
rect 3515 1298 3573 1332
rect 3515 1264 3527 1298
rect 3561 1264 3573 1298
rect 3515 1230 3573 1264
rect 3515 1196 3527 1230
rect 3561 1196 3573 1230
rect 3515 1162 3573 1196
rect 3515 1128 3527 1162
rect 3561 1128 3573 1162
rect 3515 1093 3573 1128
rect 3515 1059 3527 1093
rect 3561 1059 3573 1093
rect 3515 1004 3573 1059
rect 3603 1366 3657 1404
rect 3603 1332 3615 1366
rect 3649 1332 3657 1366
rect 3603 1298 3657 1332
rect 3603 1264 3615 1298
rect 3649 1264 3657 1298
rect 3603 1230 3657 1264
rect 3603 1196 3615 1230
rect 3649 1196 3657 1230
rect 3603 1162 3657 1196
rect 3603 1128 3615 1162
rect 3649 1128 3657 1162
rect 3603 1004 3657 1128
rect 4039 1366 4095 1404
rect 4039 1332 4049 1366
rect 4083 1332 4095 1366
rect 4039 1298 4095 1332
rect 4039 1264 4049 1298
rect 4083 1264 4095 1298
rect 4039 1230 4095 1264
rect 4039 1196 4049 1230
rect 4083 1196 4095 1230
rect 4039 1162 4095 1196
rect 4039 1128 4049 1162
rect 4083 1128 4095 1162
rect 4039 1093 4095 1128
rect 4039 1059 4049 1093
rect 4083 1059 4095 1093
rect 4039 1004 4095 1059
rect 4125 1366 4183 1404
rect 4125 1332 4137 1366
rect 4171 1332 4183 1366
rect 4125 1298 4183 1332
rect 4125 1264 4137 1298
rect 4171 1264 4183 1298
rect 4125 1230 4183 1264
rect 4125 1196 4137 1230
rect 4171 1196 4183 1230
rect 4125 1162 4183 1196
rect 4125 1128 4137 1162
rect 4171 1128 4183 1162
rect 4125 1093 4183 1128
rect 4125 1059 4137 1093
rect 4171 1059 4183 1093
rect 4125 1004 4183 1059
rect 4213 1366 4271 1404
rect 4213 1332 4225 1366
rect 4259 1332 4271 1366
rect 4213 1298 4271 1332
rect 4213 1264 4225 1298
rect 4259 1264 4271 1298
rect 4213 1230 4271 1264
rect 4213 1196 4225 1230
rect 4259 1196 4271 1230
rect 4213 1162 4271 1196
rect 4213 1128 4225 1162
rect 4259 1128 4271 1162
rect 4213 1004 4271 1128
rect 4301 1366 4359 1404
rect 4301 1332 4313 1366
rect 4347 1332 4359 1366
rect 4301 1298 4359 1332
rect 4301 1264 4313 1298
rect 4347 1264 4359 1298
rect 4301 1230 4359 1264
rect 4301 1196 4313 1230
rect 4347 1196 4359 1230
rect 4301 1162 4359 1196
rect 4301 1128 4313 1162
rect 4347 1128 4359 1162
rect 4301 1093 4359 1128
rect 4301 1059 4313 1093
rect 4347 1059 4359 1093
rect 4301 1004 4359 1059
rect 4389 1366 4447 1404
rect 4389 1332 4401 1366
rect 4435 1332 4447 1366
rect 4389 1298 4447 1332
rect 4389 1264 4401 1298
rect 4435 1264 4447 1298
rect 4389 1230 4447 1264
rect 4389 1196 4401 1230
rect 4435 1196 4447 1230
rect 4389 1162 4447 1196
rect 4389 1128 4401 1162
rect 4435 1128 4447 1162
rect 4389 1004 4447 1128
rect 4477 1366 4535 1404
rect 4477 1332 4489 1366
rect 4523 1332 4535 1366
rect 4477 1298 4535 1332
rect 4477 1264 4489 1298
rect 4523 1264 4535 1298
rect 4477 1230 4535 1264
rect 4477 1196 4489 1230
rect 4523 1196 4535 1230
rect 4477 1162 4535 1196
rect 4477 1128 4489 1162
rect 4523 1128 4535 1162
rect 4477 1093 4535 1128
rect 4477 1059 4489 1093
rect 4523 1059 4535 1093
rect 4477 1004 4535 1059
rect 4565 1366 4619 1404
rect 4565 1332 4577 1366
rect 4611 1332 4619 1366
rect 4565 1298 4619 1332
rect 4565 1264 4577 1298
rect 4611 1264 4619 1298
rect 4565 1230 4619 1264
rect 4565 1196 4577 1230
rect 4611 1196 4619 1230
rect 4565 1162 4619 1196
rect 4565 1128 4577 1162
rect 4611 1128 4619 1162
rect 4565 1004 4619 1128
rect 5001 1366 5057 1404
rect 5001 1332 5011 1366
rect 5045 1332 5057 1366
rect 5001 1298 5057 1332
rect 5001 1264 5011 1298
rect 5045 1264 5057 1298
rect 5001 1230 5057 1264
rect 5001 1196 5011 1230
rect 5045 1196 5057 1230
rect 5001 1162 5057 1196
rect 5001 1128 5011 1162
rect 5045 1128 5057 1162
rect 5001 1093 5057 1128
rect 5001 1059 5011 1093
rect 5045 1059 5057 1093
rect 5001 1004 5057 1059
rect 5087 1366 5145 1404
rect 5087 1332 5099 1366
rect 5133 1332 5145 1366
rect 5087 1298 5145 1332
rect 5087 1264 5099 1298
rect 5133 1264 5145 1298
rect 5087 1230 5145 1264
rect 5087 1196 5099 1230
rect 5133 1196 5145 1230
rect 5087 1162 5145 1196
rect 5087 1128 5099 1162
rect 5133 1128 5145 1162
rect 5087 1093 5145 1128
rect 5087 1059 5099 1093
rect 5133 1059 5145 1093
rect 5087 1004 5145 1059
rect 5175 1366 5233 1404
rect 5175 1332 5187 1366
rect 5221 1332 5233 1366
rect 5175 1298 5233 1332
rect 5175 1264 5187 1298
rect 5221 1264 5233 1298
rect 5175 1230 5233 1264
rect 5175 1196 5187 1230
rect 5221 1196 5233 1230
rect 5175 1162 5233 1196
rect 5175 1128 5187 1162
rect 5221 1128 5233 1162
rect 5175 1004 5233 1128
rect 5263 1366 5321 1404
rect 5263 1332 5275 1366
rect 5309 1332 5321 1366
rect 5263 1298 5321 1332
rect 5263 1264 5275 1298
rect 5309 1264 5321 1298
rect 5263 1230 5321 1264
rect 5263 1196 5275 1230
rect 5309 1196 5321 1230
rect 5263 1162 5321 1196
rect 5263 1128 5275 1162
rect 5309 1128 5321 1162
rect 5263 1093 5321 1128
rect 5263 1059 5275 1093
rect 5309 1059 5321 1093
rect 5263 1004 5321 1059
rect 5351 1366 5409 1404
rect 5351 1332 5363 1366
rect 5397 1332 5409 1366
rect 5351 1298 5409 1332
rect 5351 1264 5363 1298
rect 5397 1264 5409 1298
rect 5351 1230 5409 1264
rect 5351 1196 5363 1230
rect 5397 1196 5409 1230
rect 5351 1162 5409 1196
rect 5351 1128 5363 1162
rect 5397 1128 5409 1162
rect 5351 1004 5409 1128
rect 5439 1366 5497 1404
rect 5439 1332 5451 1366
rect 5485 1332 5497 1366
rect 5439 1298 5497 1332
rect 5439 1264 5451 1298
rect 5485 1264 5497 1298
rect 5439 1230 5497 1264
rect 5439 1196 5451 1230
rect 5485 1196 5497 1230
rect 5439 1162 5497 1196
rect 5439 1128 5451 1162
rect 5485 1128 5497 1162
rect 5439 1093 5497 1128
rect 5439 1059 5451 1093
rect 5485 1059 5497 1093
rect 5439 1004 5497 1059
rect 5527 1366 5581 1404
rect 5527 1332 5539 1366
rect 5573 1332 5581 1366
rect 5527 1298 5581 1332
rect 5527 1264 5539 1298
rect 5573 1264 5581 1298
rect 5527 1230 5581 1264
rect 5527 1196 5539 1230
rect 5573 1196 5581 1230
rect 5527 1162 5581 1196
rect 5527 1128 5539 1162
rect 5573 1128 5581 1162
rect 5527 1004 5581 1128
<< ndiffc >>
rect 101 301 135 335
rect 198 301 232 335
rect 295 301 329 335
rect 392 301 426 335
rect 489 301 523 335
rect 101 229 135 263
rect 101 161 135 195
rect 198 176 232 210
rect 295 229 329 263
rect 295 161 329 195
rect 393 182 427 216
rect 101 91 135 125
rect 295 91 329 125
rect 392 91 426 125
rect 489 91 523 125
rect 603 301 637 335
rect 603 229 637 263
rect 603 161 637 195
rect 700 185 734 219
rect 797 229 831 263
rect 797 161 831 195
rect 603 91 637 125
rect 700 91 734 125
rect 797 91 831 125
rect 1063 301 1097 335
rect 1160 301 1194 335
rect 1257 301 1291 335
rect 1354 301 1388 335
rect 1451 301 1485 335
rect 1063 229 1097 263
rect 1063 161 1097 195
rect 1160 176 1194 210
rect 1257 229 1291 263
rect 1257 161 1291 195
rect 1355 182 1389 216
rect 1063 91 1097 125
rect 1257 91 1291 125
rect 1354 91 1388 125
rect 1451 91 1485 125
rect 1565 301 1599 335
rect 1565 229 1599 263
rect 1565 161 1599 195
rect 1662 185 1696 219
rect 1759 229 1793 263
rect 1759 161 1793 195
rect 1565 91 1599 125
rect 1662 91 1696 125
rect 1759 91 1793 125
rect 2025 301 2059 335
rect 2122 301 2156 335
rect 2219 301 2253 335
rect 2316 301 2350 335
rect 2413 301 2447 335
rect 2025 229 2059 263
rect 2025 161 2059 195
rect 2122 176 2156 210
rect 2219 229 2253 263
rect 2219 161 2253 195
rect 2317 182 2351 216
rect 2025 91 2059 125
rect 2219 91 2253 125
rect 2316 91 2350 125
rect 2413 91 2447 125
rect 2527 301 2561 335
rect 2527 229 2561 263
rect 2527 161 2561 195
rect 2624 185 2658 219
rect 2721 229 2755 263
rect 2721 161 2755 195
rect 2527 91 2561 125
rect 2624 91 2658 125
rect 2721 91 2755 125
rect 2987 301 3021 335
rect 3084 301 3118 335
rect 3181 301 3215 335
rect 3278 301 3312 335
rect 3375 301 3409 335
rect 2987 229 3021 263
rect 2987 161 3021 195
rect 3084 176 3118 210
rect 3181 229 3215 263
rect 3181 161 3215 195
rect 3279 182 3313 216
rect 2987 91 3021 125
rect 3181 91 3215 125
rect 3278 91 3312 125
rect 3375 91 3409 125
rect 3489 301 3523 335
rect 3489 229 3523 263
rect 3489 161 3523 195
rect 3586 185 3620 219
rect 3683 229 3717 263
rect 3683 161 3717 195
rect 3489 91 3523 125
rect 3586 91 3620 125
rect 3683 91 3717 125
rect 3949 301 3983 335
rect 4046 301 4080 335
rect 4143 301 4177 335
rect 4240 301 4274 335
rect 4337 301 4371 335
rect 3949 229 3983 263
rect 3949 161 3983 195
rect 4046 176 4080 210
rect 4143 229 4177 263
rect 4143 161 4177 195
rect 4241 182 4275 216
rect 3949 91 3983 125
rect 4143 91 4177 125
rect 4240 91 4274 125
rect 4337 91 4371 125
rect 4451 301 4485 335
rect 4451 229 4485 263
rect 4451 161 4485 195
rect 4548 185 4582 219
rect 4645 229 4679 263
rect 4645 161 4679 195
rect 4451 91 4485 125
rect 4548 91 4582 125
rect 4645 91 4679 125
rect 4911 301 4945 335
rect 5008 301 5042 335
rect 5105 301 5139 335
rect 5202 301 5236 335
rect 5299 301 5333 335
rect 4911 229 4945 263
rect 4911 161 4945 195
rect 5008 176 5042 210
rect 5105 229 5139 263
rect 5105 161 5139 195
rect 5203 182 5237 216
rect 4911 91 4945 125
rect 5105 91 5139 125
rect 5202 91 5236 125
rect 5299 91 5333 125
rect 5413 301 5447 335
rect 5413 229 5447 263
rect 5413 161 5447 195
rect 5510 185 5544 219
rect 5607 229 5641 263
rect 5607 161 5641 195
rect 5413 91 5447 125
rect 5510 91 5544 125
rect 5607 91 5641 125
<< pdiffc >>
rect 201 1332 235 1366
rect 201 1264 235 1298
rect 201 1196 235 1230
rect 201 1128 235 1162
rect 201 1059 235 1093
rect 289 1332 323 1366
rect 289 1264 323 1298
rect 289 1196 323 1230
rect 289 1128 323 1162
rect 289 1059 323 1093
rect 377 1332 411 1366
rect 377 1264 411 1298
rect 377 1196 411 1230
rect 377 1128 411 1162
rect 465 1332 499 1366
rect 465 1264 499 1298
rect 465 1196 499 1230
rect 465 1128 499 1162
rect 465 1059 499 1093
rect 553 1332 587 1366
rect 553 1264 587 1298
rect 553 1196 587 1230
rect 553 1128 587 1162
rect 641 1332 675 1366
rect 641 1264 675 1298
rect 641 1196 675 1230
rect 641 1128 675 1162
rect 641 1059 675 1093
rect 729 1332 763 1366
rect 729 1264 763 1298
rect 729 1196 763 1230
rect 729 1128 763 1162
rect 1163 1332 1197 1366
rect 1163 1264 1197 1298
rect 1163 1196 1197 1230
rect 1163 1128 1197 1162
rect 1163 1059 1197 1093
rect 1251 1332 1285 1366
rect 1251 1264 1285 1298
rect 1251 1196 1285 1230
rect 1251 1128 1285 1162
rect 1251 1059 1285 1093
rect 1339 1332 1373 1366
rect 1339 1264 1373 1298
rect 1339 1196 1373 1230
rect 1339 1128 1373 1162
rect 1427 1332 1461 1366
rect 1427 1264 1461 1298
rect 1427 1196 1461 1230
rect 1427 1128 1461 1162
rect 1427 1059 1461 1093
rect 1515 1332 1549 1366
rect 1515 1264 1549 1298
rect 1515 1196 1549 1230
rect 1515 1128 1549 1162
rect 1603 1332 1637 1366
rect 1603 1264 1637 1298
rect 1603 1196 1637 1230
rect 1603 1128 1637 1162
rect 1603 1059 1637 1093
rect 1691 1332 1725 1366
rect 1691 1264 1725 1298
rect 1691 1196 1725 1230
rect 1691 1128 1725 1162
rect 2125 1332 2159 1366
rect 2125 1264 2159 1298
rect 2125 1196 2159 1230
rect 2125 1128 2159 1162
rect 2125 1059 2159 1093
rect 2213 1332 2247 1366
rect 2213 1264 2247 1298
rect 2213 1196 2247 1230
rect 2213 1128 2247 1162
rect 2213 1059 2247 1093
rect 2301 1332 2335 1366
rect 2301 1264 2335 1298
rect 2301 1196 2335 1230
rect 2301 1128 2335 1162
rect 2389 1332 2423 1366
rect 2389 1264 2423 1298
rect 2389 1196 2423 1230
rect 2389 1128 2423 1162
rect 2389 1059 2423 1093
rect 2477 1332 2511 1366
rect 2477 1264 2511 1298
rect 2477 1196 2511 1230
rect 2477 1128 2511 1162
rect 2565 1332 2599 1366
rect 2565 1264 2599 1298
rect 2565 1196 2599 1230
rect 2565 1128 2599 1162
rect 2565 1059 2599 1093
rect 2653 1332 2687 1366
rect 2653 1264 2687 1298
rect 2653 1196 2687 1230
rect 2653 1128 2687 1162
rect 3087 1332 3121 1366
rect 3087 1264 3121 1298
rect 3087 1196 3121 1230
rect 3087 1128 3121 1162
rect 3087 1059 3121 1093
rect 3175 1332 3209 1366
rect 3175 1264 3209 1298
rect 3175 1196 3209 1230
rect 3175 1128 3209 1162
rect 3175 1059 3209 1093
rect 3263 1332 3297 1366
rect 3263 1264 3297 1298
rect 3263 1196 3297 1230
rect 3263 1128 3297 1162
rect 3351 1332 3385 1366
rect 3351 1264 3385 1298
rect 3351 1196 3385 1230
rect 3351 1128 3385 1162
rect 3351 1059 3385 1093
rect 3439 1332 3473 1366
rect 3439 1264 3473 1298
rect 3439 1196 3473 1230
rect 3439 1128 3473 1162
rect 3527 1332 3561 1366
rect 3527 1264 3561 1298
rect 3527 1196 3561 1230
rect 3527 1128 3561 1162
rect 3527 1059 3561 1093
rect 3615 1332 3649 1366
rect 3615 1264 3649 1298
rect 3615 1196 3649 1230
rect 3615 1128 3649 1162
rect 4049 1332 4083 1366
rect 4049 1264 4083 1298
rect 4049 1196 4083 1230
rect 4049 1128 4083 1162
rect 4049 1059 4083 1093
rect 4137 1332 4171 1366
rect 4137 1264 4171 1298
rect 4137 1196 4171 1230
rect 4137 1128 4171 1162
rect 4137 1059 4171 1093
rect 4225 1332 4259 1366
rect 4225 1264 4259 1298
rect 4225 1196 4259 1230
rect 4225 1128 4259 1162
rect 4313 1332 4347 1366
rect 4313 1264 4347 1298
rect 4313 1196 4347 1230
rect 4313 1128 4347 1162
rect 4313 1059 4347 1093
rect 4401 1332 4435 1366
rect 4401 1264 4435 1298
rect 4401 1196 4435 1230
rect 4401 1128 4435 1162
rect 4489 1332 4523 1366
rect 4489 1264 4523 1298
rect 4489 1196 4523 1230
rect 4489 1128 4523 1162
rect 4489 1059 4523 1093
rect 4577 1332 4611 1366
rect 4577 1264 4611 1298
rect 4577 1196 4611 1230
rect 4577 1128 4611 1162
rect 5011 1332 5045 1366
rect 5011 1264 5045 1298
rect 5011 1196 5045 1230
rect 5011 1128 5045 1162
rect 5011 1059 5045 1093
rect 5099 1332 5133 1366
rect 5099 1264 5133 1298
rect 5099 1196 5133 1230
rect 5099 1128 5133 1162
rect 5099 1059 5133 1093
rect 5187 1332 5221 1366
rect 5187 1264 5221 1298
rect 5187 1196 5221 1230
rect 5187 1128 5221 1162
rect 5275 1332 5309 1366
rect 5275 1264 5309 1298
rect 5275 1196 5309 1230
rect 5275 1128 5309 1162
rect 5275 1059 5309 1093
rect 5363 1332 5397 1366
rect 5363 1264 5397 1298
rect 5363 1196 5397 1230
rect 5363 1128 5397 1162
rect 5451 1332 5485 1366
rect 5451 1264 5485 1298
rect 5451 1196 5485 1230
rect 5451 1128 5485 1162
rect 5451 1059 5485 1093
rect 5539 1332 5573 1366
rect 5539 1264 5573 1298
rect 5539 1196 5573 1230
rect 5539 1128 5573 1162
<< psubdiff >>
rect -34 482 5806 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 928 461 996 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 928 427 945 461
rect 979 427 996 461
rect 1890 461 1958 482
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 928 313 996 353
rect 1890 427 1907 461
rect 1941 427 1958 461
rect 2852 461 2920 482
rect 1890 387 1958 427
rect 1890 353 1907 387
rect 1941 353 1958 387
rect 928 279 945 313
rect 979 279 996 313
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect -34 17 34 57
rect 928 57 945 91
rect 979 57 996 91
rect 1890 313 1958 353
rect 2852 427 2869 461
rect 2903 427 2920 461
rect 3814 461 3882 482
rect 2852 387 2920 427
rect 2852 353 2869 387
rect 2903 353 2920 387
rect 1890 279 1907 313
rect 1941 279 1958 313
rect 1890 239 1958 279
rect 1890 205 1907 239
rect 1941 205 1958 239
rect 1890 165 1958 205
rect 1890 131 1907 165
rect 1941 131 1958 165
rect 1890 91 1958 131
rect 928 17 996 57
rect 1890 57 1907 91
rect 1941 57 1958 91
rect 2852 313 2920 353
rect 3814 427 3831 461
rect 3865 427 3882 461
rect 4776 461 4844 482
rect 3814 387 3882 427
rect 3814 353 3831 387
rect 3865 353 3882 387
rect 2852 279 2869 313
rect 2903 279 2920 313
rect 2852 239 2920 279
rect 2852 205 2869 239
rect 2903 205 2920 239
rect 2852 165 2920 205
rect 2852 131 2869 165
rect 2903 131 2920 165
rect 2852 91 2920 131
rect 1890 17 1958 57
rect 2852 57 2869 91
rect 2903 57 2920 91
rect 3814 313 3882 353
rect 4776 427 4793 461
rect 4827 427 4844 461
rect 5738 461 5806 482
rect 4776 387 4844 427
rect 4776 353 4793 387
rect 4827 353 4844 387
rect 3814 279 3831 313
rect 3865 279 3882 313
rect 3814 239 3882 279
rect 3814 205 3831 239
rect 3865 205 3882 239
rect 3814 165 3882 205
rect 3814 131 3831 165
rect 3865 131 3882 165
rect 3814 91 3882 131
rect 2852 17 2920 57
rect 3814 57 3831 91
rect 3865 57 3882 91
rect 4776 313 4844 353
rect 5738 427 5755 461
rect 5789 427 5806 461
rect 5738 387 5806 427
rect 5738 353 5755 387
rect 5789 353 5806 387
rect 4776 279 4793 313
rect 4827 279 4844 313
rect 4776 239 4844 279
rect 4776 205 4793 239
rect 4827 205 4844 239
rect 4776 165 4844 205
rect 4776 131 4793 165
rect 4827 131 4844 165
rect 4776 91 4844 131
rect 3814 17 3882 57
rect 4776 57 4793 91
rect 4827 57 4844 91
rect 5738 313 5806 353
rect 5738 279 5755 313
rect 5789 279 5806 313
rect 5738 239 5806 279
rect 5738 205 5755 239
rect 5789 205 5806 239
rect 5738 165 5806 205
rect 5738 131 5755 165
rect 5789 131 5806 165
rect 5738 91 5806 131
rect 4776 17 4844 57
rect 5738 57 5755 91
rect 5789 57 5806 91
rect 5738 17 5806 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5806 17
rect -34 -34 5806 -17
<< nsubdiff >>
rect -34 1497 5806 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5806 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 928 1423 996 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 1890 1423 1958 1463
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect 928 1019 945 1053
rect 979 1019 996 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 928 979 996 1019
rect 1890 1389 1907 1423
rect 1941 1389 1958 1423
rect 2852 1423 2920 1463
rect 1890 1349 1958 1389
rect 1890 1315 1907 1349
rect 1941 1315 1958 1349
rect 1890 1275 1958 1315
rect 1890 1241 1907 1275
rect 1941 1241 1958 1275
rect 1890 1201 1958 1241
rect 1890 1167 1907 1201
rect 1941 1167 1958 1201
rect 1890 1127 1958 1167
rect 1890 1093 1907 1127
rect 1941 1093 1958 1127
rect 1890 1053 1958 1093
rect 1890 1019 1907 1053
rect 1941 1019 1958 1053
rect 928 945 945 979
rect 979 945 996 979
rect -34 871 -17 905
rect 17 884 34 905
rect 928 905 996 945
rect 1890 979 1958 1019
rect 2852 1389 2869 1423
rect 2903 1389 2920 1423
rect 3814 1423 3882 1463
rect 2852 1349 2920 1389
rect 2852 1315 2869 1349
rect 2903 1315 2920 1349
rect 2852 1275 2920 1315
rect 2852 1241 2869 1275
rect 2903 1241 2920 1275
rect 2852 1201 2920 1241
rect 2852 1167 2869 1201
rect 2903 1167 2920 1201
rect 2852 1127 2920 1167
rect 2852 1093 2869 1127
rect 2903 1093 2920 1127
rect 2852 1053 2920 1093
rect 2852 1019 2869 1053
rect 2903 1019 2920 1053
rect 1890 945 1907 979
rect 1941 945 1958 979
rect 928 884 945 905
rect 17 871 945 884
rect 979 884 996 905
rect 1890 905 1958 945
rect 2852 979 2920 1019
rect 3814 1389 3831 1423
rect 3865 1389 3882 1423
rect 4776 1423 4844 1463
rect 3814 1349 3882 1389
rect 3814 1315 3831 1349
rect 3865 1315 3882 1349
rect 3814 1275 3882 1315
rect 3814 1241 3831 1275
rect 3865 1241 3882 1275
rect 3814 1201 3882 1241
rect 3814 1167 3831 1201
rect 3865 1167 3882 1201
rect 3814 1127 3882 1167
rect 3814 1093 3831 1127
rect 3865 1093 3882 1127
rect 3814 1053 3882 1093
rect 3814 1019 3831 1053
rect 3865 1019 3882 1053
rect 2852 945 2869 979
rect 2903 945 2920 979
rect 1890 884 1907 905
rect 979 871 1907 884
rect 1941 884 1958 905
rect 2852 905 2920 945
rect 3814 979 3882 1019
rect 4776 1389 4793 1423
rect 4827 1389 4844 1423
rect 5738 1423 5806 1463
rect 4776 1349 4844 1389
rect 4776 1315 4793 1349
rect 4827 1315 4844 1349
rect 4776 1275 4844 1315
rect 4776 1241 4793 1275
rect 4827 1241 4844 1275
rect 4776 1201 4844 1241
rect 4776 1167 4793 1201
rect 4827 1167 4844 1201
rect 4776 1127 4844 1167
rect 4776 1093 4793 1127
rect 4827 1093 4844 1127
rect 4776 1053 4844 1093
rect 4776 1019 4793 1053
rect 4827 1019 4844 1053
rect 3814 945 3831 979
rect 3865 945 3882 979
rect 2852 884 2869 905
rect 1941 871 2869 884
rect 2903 884 2920 905
rect 3814 905 3882 945
rect 4776 979 4844 1019
rect 5738 1389 5755 1423
rect 5789 1389 5806 1423
rect 5738 1349 5806 1389
rect 5738 1315 5755 1349
rect 5789 1315 5806 1349
rect 5738 1275 5806 1315
rect 5738 1241 5755 1275
rect 5789 1241 5806 1275
rect 5738 1201 5806 1241
rect 5738 1167 5755 1201
rect 5789 1167 5806 1201
rect 5738 1127 5806 1167
rect 5738 1093 5755 1127
rect 5789 1093 5806 1127
rect 5738 1053 5806 1093
rect 5738 1019 5755 1053
rect 5789 1019 5806 1053
rect 4776 945 4793 979
rect 4827 945 4844 979
rect 3814 884 3831 905
rect 2903 871 3831 884
rect 3865 884 3882 905
rect 4776 905 4844 945
rect 5738 979 5806 1019
rect 5738 945 5755 979
rect 5789 945 5806 979
rect 4776 884 4793 905
rect 3865 871 4793 884
rect 4827 884 4844 905
rect 5738 905 5806 945
rect 5738 884 5755 905
rect 4827 871 5755 884
rect 5789 871 5806 905
rect -34 822 5806 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 945 427 979 461
rect 945 353 979 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1907 427 1941 461
rect 1907 353 1941 387
rect 945 279 979 313
rect 945 205 979 239
rect 945 131 979 165
rect 945 57 979 91
rect 2869 427 2903 461
rect 2869 353 2903 387
rect 1907 279 1941 313
rect 1907 205 1941 239
rect 1907 131 1941 165
rect 1907 57 1941 91
rect 3831 427 3865 461
rect 3831 353 3865 387
rect 2869 279 2903 313
rect 2869 205 2903 239
rect 2869 131 2903 165
rect 2869 57 2903 91
rect 4793 427 4827 461
rect 4793 353 4827 387
rect 3831 279 3865 313
rect 3831 205 3865 239
rect 3831 131 3865 165
rect 3831 57 3865 91
rect 5755 427 5789 461
rect 5755 353 5789 387
rect 4793 279 4827 313
rect 4793 205 4827 239
rect 4793 131 4827 165
rect 4793 57 4827 91
rect 5755 279 5789 313
rect 5755 205 5789 239
rect 5755 131 5789 165
rect 5755 57 5789 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5163 -17 5197 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5533 -17 5567 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5163 1463 5197 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5533 1463 5567 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 945 1389 979 1423
rect 945 1315 979 1349
rect 945 1241 979 1275
rect 945 1167 979 1201
rect 945 1093 979 1127
rect 945 1019 979 1053
rect -17 945 17 979
rect 1907 1389 1941 1423
rect 1907 1315 1941 1349
rect 1907 1241 1941 1275
rect 1907 1167 1941 1201
rect 1907 1093 1941 1127
rect 1907 1019 1941 1053
rect 945 945 979 979
rect -17 871 17 905
rect 2869 1389 2903 1423
rect 2869 1315 2903 1349
rect 2869 1241 2903 1275
rect 2869 1167 2903 1201
rect 2869 1093 2903 1127
rect 2869 1019 2903 1053
rect 1907 945 1941 979
rect 945 871 979 905
rect 3831 1389 3865 1423
rect 3831 1315 3865 1349
rect 3831 1241 3865 1275
rect 3831 1167 3865 1201
rect 3831 1093 3865 1127
rect 3831 1019 3865 1053
rect 2869 945 2903 979
rect 1907 871 1941 905
rect 4793 1389 4827 1423
rect 4793 1315 4827 1349
rect 4793 1241 4827 1275
rect 4793 1167 4827 1201
rect 4793 1093 4827 1127
rect 4793 1019 4827 1053
rect 3831 945 3865 979
rect 2869 871 2903 905
rect 5755 1389 5789 1423
rect 5755 1315 5789 1349
rect 5755 1241 5789 1275
rect 5755 1167 5789 1201
rect 5755 1093 5789 1127
rect 5755 1019 5789 1053
rect 4793 945 4827 979
rect 3831 871 3865 905
rect 5755 945 5789 979
rect 4793 871 4827 905
rect 5755 871 5789 905
<< poly >>
rect 247 1404 277 1430
rect 335 1404 365 1430
rect 423 1404 453 1430
rect 511 1404 541 1430
rect 599 1404 629 1430
rect 687 1404 717 1430
rect 1209 1404 1239 1430
rect 1297 1404 1327 1430
rect 1385 1404 1415 1430
rect 1473 1404 1503 1430
rect 1561 1404 1591 1430
rect 1649 1404 1679 1430
rect 247 973 277 1004
rect 335 973 365 1004
rect 423 973 453 1004
rect 511 973 541 1004
rect 195 957 365 973
rect 195 923 205 957
rect 239 943 365 957
rect 417 957 541 973
rect 239 923 249 943
rect 195 907 249 923
rect 417 923 427 957
rect 461 943 541 957
rect 599 973 629 1004
rect 687 973 717 1004
rect 599 957 717 973
rect 599 943 649 957
rect 461 923 471 943
rect 417 907 471 923
rect 639 923 649 943
rect 683 943 717 957
rect 2171 1404 2201 1430
rect 2259 1404 2289 1430
rect 2347 1404 2377 1430
rect 2435 1404 2465 1430
rect 2523 1404 2553 1430
rect 2611 1404 2641 1430
rect 1209 973 1239 1004
rect 1297 973 1327 1004
rect 1385 973 1415 1004
rect 1473 973 1503 1004
rect 683 923 693 943
rect 639 907 693 923
rect 1157 957 1327 973
rect 1157 923 1167 957
rect 1201 943 1327 957
rect 1379 957 1503 973
rect 1201 923 1211 943
rect 1157 907 1211 923
rect 1379 923 1389 957
rect 1423 943 1503 957
rect 1561 973 1591 1004
rect 1649 973 1679 1004
rect 1561 957 1679 973
rect 1561 943 1611 957
rect 1423 923 1433 943
rect 1379 907 1433 923
rect 1601 923 1611 943
rect 1645 943 1679 957
rect 3133 1404 3163 1430
rect 3221 1404 3251 1430
rect 3309 1404 3339 1430
rect 3397 1404 3427 1430
rect 3485 1404 3515 1430
rect 3573 1404 3603 1430
rect 2171 973 2201 1004
rect 2259 973 2289 1004
rect 2347 973 2377 1004
rect 2435 973 2465 1004
rect 1645 923 1655 943
rect 1601 907 1655 923
rect 2119 957 2289 973
rect 2119 923 2129 957
rect 2163 943 2289 957
rect 2341 957 2465 973
rect 2163 923 2173 943
rect 2119 907 2173 923
rect 2341 923 2351 957
rect 2385 943 2465 957
rect 2523 973 2553 1004
rect 2611 973 2641 1004
rect 2523 957 2641 973
rect 2523 943 2573 957
rect 2385 923 2395 943
rect 2341 907 2395 923
rect 2563 923 2573 943
rect 2607 943 2641 957
rect 4095 1404 4125 1430
rect 4183 1404 4213 1430
rect 4271 1404 4301 1430
rect 4359 1404 4389 1430
rect 4447 1404 4477 1430
rect 4535 1404 4565 1430
rect 3133 973 3163 1004
rect 3221 973 3251 1004
rect 3309 973 3339 1004
rect 3397 973 3427 1004
rect 2607 923 2617 943
rect 2563 907 2617 923
rect 3081 957 3251 973
rect 3081 923 3091 957
rect 3125 943 3251 957
rect 3303 957 3427 973
rect 3125 923 3135 943
rect 3081 907 3135 923
rect 3303 923 3313 957
rect 3347 943 3427 957
rect 3485 973 3515 1004
rect 3573 973 3603 1004
rect 3485 957 3603 973
rect 3485 943 3535 957
rect 3347 923 3357 943
rect 3303 907 3357 923
rect 3525 923 3535 943
rect 3569 943 3603 957
rect 5057 1404 5087 1430
rect 5145 1404 5175 1430
rect 5233 1404 5263 1430
rect 5321 1404 5351 1430
rect 5409 1404 5439 1430
rect 5497 1404 5527 1430
rect 4095 973 4125 1004
rect 4183 973 4213 1004
rect 4271 973 4301 1004
rect 4359 973 4389 1004
rect 3569 923 3579 943
rect 3525 907 3579 923
rect 4043 957 4213 973
rect 4043 923 4053 957
rect 4087 943 4213 957
rect 4265 957 4389 973
rect 4087 923 4097 943
rect 4043 907 4097 923
rect 4265 923 4275 957
rect 4309 943 4389 957
rect 4447 973 4477 1004
rect 4535 973 4565 1004
rect 4447 957 4565 973
rect 4447 943 4497 957
rect 4309 923 4319 943
rect 4265 907 4319 923
rect 4487 923 4497 943
rect 4531 943 4565 957
rect 5057 973 5087 1004
rect 5145 973 5175 1004
rect 5233 973 5263 1004
rect 5321 973 5351 1004
rect 4531 923 4541 943
rect 4487 907 4541 923
rect 5005 957 5175 973
rect 5005 923 5015 957
rect 5049 943 5175 957
rect 5227 957 5351 973
rect 5049 923 5059 943
rect 5005 907 5059 923
rect 5227 923 5237 957
rect 5271 943 5351 957
rect 5409 973 5439 1004
rect 5497 973 5527 1004
rect 5409 957 5527 973
rect 5409 943 5459 957
rect 5271 923 5281 943
rect 5227 907 5281 923
rect 5449 923 5459 943
rect 5493 943 5527 957
rect 5493 923 5503 943
rect 5449 907 5503 923
rect 195 433 249 449
rect 195 413 205 433
rect 147 399 205 413
rect 239 399 249 433
rect 147 383 249 399
rect 417 433 471 449
rect 417 399 427 433
rect 461 413 471 433
rect 639 433 693 449
rect 461 399 477 413
rect 417 383 477 399
rect 639 399 649 433
rect 683 399 693 433
rect 639 383 693 399
rect 1157 433 1211 449
rect 1157 413 1167 433
rect 147 351 177 383
rect 447 351 477 383
rect 649 351 679 383
rect 1109 399 1167 413
rect 1201 399 1211 433
rect 1109 383 1211 399
rect 1379 433 1433 449
rect 1379 399 1389 433
rect 1423 413 1433 433
rect 1601 433 1655 449
rect 1423 399 1439 413
rect 1379 383 1439 399
rect 1601 399 1611 433
rect 1645 399 1655 433
rect 1601 383 1655 399
rect 2119 433 2173 449
rect 2119 413 2129 433
rect 1109 351 1139 383
rect 1409 351 1439 383
rect 1611 351 1641 383
rect 2071 399 2129 413
rect 2163 399 2173 433
rect 2071 383 2173 399
rect 2341 433 2395 449
rect 2341 399 2351 433
rect 2385 413 2395 433
rect 2563 433 2617 449
rect 2385 399 2401 413
rect 2341 383 2401 399
rect 2563 399 2573 433
rect 2607 399 2617 433
rect 2563 383 2617 399
rect 3081 433 3135 449
rect 3081 413 3091 433
rect 2071 351 2101 383
rect 2371 351 2401 383
rect 2573 351 2603 383
rect 3033 399 3091 413
rect 3125 399 3135 433
rect 3033 383 3135 399
rect 3303 433 3357 449
rect 3303 399 3313 433
rect 3347 413 3357 433
rect 3525 433 3579 449
rect 3347 399 3363 413
rect 3303 383 3363 399
rect 3525 399 3535 433
rect 3569 399 3579 433
rect 3525 383 3579 399
rect 4043 433 4097 449
rect 4043 413 4053 433
rect 3033 351 3063 383
rect 3333 351 3363 383
rect 3535 351 3565 383
rect 3995 399 4053 413
rect 4087 399 4097 433
rect 3995 383 4097 399
rect 4265 433 4319 449
rect 4265 399 4275 433
rect 4309 413 4319 433
rect 4487 433 4541 449
rect 4309 399 4325 413
rect 4265 383 4325 399
rect 4487 399 4497 433
rect 4531 399 4541 433
rect 4487 383 4541 399
rect 5005 433 5059 449
rect 5005 413 5015 433
rect 3995 351 4025 383
rect 4295 351 4325 383
rect 4497 351 4527 383
rect 4957 399 5015 413
rect 5049 399 5059 433
rect 4957 383 5059 399
rect 5227 433 5281 449
rect 5227 399 5237 433
rect 5271 413 5281 433
rect 5449 433 5503 449
rect 5271 399 5287 413
rect 5227 383 5287 399
rect 5449 399 5459 433
rect 5493 399 5503 433
rect 5449 383 5503 399
rect 4957 351 4987 383
rect 5257 351 5287 383
rect 5459 351 5489 383
<< polycont >>
rect 205 923 239 957
rect 427 923 461 957
rect 649 923 683 957
rect 1167 923 1201 957
rect 1389 923 1423 957
rect 1611 923 1645 957
rect 2129 923 2163 957
rect 2351 923 2385 957
rect 2573 923 2607 957
rect 3091 923 3125 957
rect 3313 923 3347 957
rect 3535 923 3569 957
rect 4053 923 4087 957
rect 4275 923 4309 957
rect 4497 923 4531 957
rect 5015 923 5049 957
rect 5237 923 5271 957
rect 5459 923 5493 957
rect 205 399 239 433
rect 427 399 461 433
rect 649 399 683 433
rect 1167 399 1201 433
rect 1389 399 1423 433
rect 1611 399 1645 433
rect 2129 399 2163 433
rect 2351 399 2385 433
rect 2573 399 2607 433
rect 3091 399 3125 433
rect 3313 399 3347 433
rect 3535 399 3569 433
rect 4053 399 4087 433
rect 4275 399 4309 433
rect 4497 399 4531 433
rect 5015 399 5049 433
rect 5237 399 5271 433
rect 5459 399 5493 433
<< locali >>
rect -34 1497 5806 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5806 1497
rect -34 1446 5806 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 201 1366 235 1446
rect 201 1298 235 1332
rect 201 1230 235 1264
rect 201 1162 235 1196
rect 201 1093 235 1128
rect 201 1043 235 1059
rect 289 1366 323 1404
rect 289 1298 323 1332
rect 289 1230 323 1264
rect 289 1162 323 1196
rect 289 1093 323 1128
rect 377 1366 411 1446
rect 377 1298 411 1332
rect 377 1230 411 1264
rect 377 1162 411 1196
rect 377 1111 411 1128
rect 465 1366 499 1404
rect 465 1298 499 1332
rect 465 1230 499 1264
rect 465 1162 499 1196
rect 289 1048 323 1059
rect 465 1093 499 1128
rect 553 1366 587 1446
rect 553 1298 587 1332
rect 553 1230 587 1264
rect 553 1162 587 1196
rect 553 1111 587 1128
rect 641 1366 675 1404
rect 641 1298 675 1332
rect 641 1230 675 1264
rect 641 1162 675 1196
rect 465 1048 499 1059
rect 641 1093 675 1128
rect 729 1366 763 1446
rect 729 1298 763 1332
rect 729 1230 763 1264
rect 729 1162 763 1196
rect 729 1111 763 1128
rect 928 1423 996 1446
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 641 1048 675 1059
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect -34 979 34 1019
rect 289 1014 831 1048
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 923
rect 205 383 239 399
rect 427 957 461 973
rect 427 905 461 923
rect 427 433 461 871
rect 427 383 461 399
rect 649 957 683 973
rect 649 757 683 923
rect 649 433 683 723
rect 649 383 683 399
rect 797 610 831 1014
rect 928 1019 945 1053
rect 979 1019 996 1053
rect 1163 1366 1197 1446
rect 1163 1298 1197 1332
rect 1163 1230 1197 1264
rect 1163 1162 1197 1196
rect 1163 1093 1197 1128
rect 1163 1043 1197 1059
rect 1251 1366 1285 1404
rect 1251 1298 1285 1332
rect 1251 1230 1285 1264
rect 1251 1162 1285 1196
rect 1251 1093 1285 1128
rect 1339 1366 1373 1446
rect 1339 1298 1373 1332
rect 1339 1230 1373 1264
rect 1339 1162 1373 1196
rect 1339 1111 1373 1128
rect 1427 1366 1461 1404
rect 1427 1298 1461 1332
rect 1427 1230 1461 1264
rect 1427 1162 1461 1196
rect 1251 1048 1285 1059
rect 1427 1093 1461 1128
rect 1515 1366 1549 1446
rect 1515 1298 1549 1332
rect 1515 1230 1549 1264
rect 1515 1162 1549 1196
rect 1515 1111 1549 1128
rect 1603 1366 1637 1404
rect 1603 1298 1637 1332
rect 1603 1230 1637 1264
rect 1603 1162 1637 1196
rect 1427 1048 1461 1059
rect 1603 1093 1637 1128
rect 1691 1366 1725 1446
rect 1691 1298 1725 1332
rect 1691 1230 1725 1264
rect 1691 1162 1725 1196
rect 1691 1111 1725 1128
rect 1890 1423 1958 1446
rect 1890 1389 1907 1423
rect 1941 1389 1958 1423
rect 1890 1349 1958 1389
rect 1890 1315 1907 1349
rect 1941 1315 1958 1349
rect 1890 1275 1958 1315
rect 1890 1241 1907 1275
rect 1941 1241 1958 1275
rect 1890 1201 1958 1241
rect 1890 1167 1907 1201
rect 1941 1167 1958 1201
rect 1890 1127 1958 1167
rect 1603 1048 1637 1059
rect 1890 1093 1907 1127
rect 1941 1093 1958 1127
rect 1890 1053 1958 1093
rect 928 979 996 1019
rect 1251 1014 1793 1048
rect 928 945 945 979
rect 979 945 996 979
rect 928 905 996 945
rect 928 871 945 905
rect 979 871 996 905
rect 928 822 996 871
rect 1167 957 1201 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 101 335 135 351
rect 295 335 329 351
rect 489 335 523 351
rect 135 301 198 335
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 489 335
rect 101 263 135 301
rect 101 195 135 229
rect 295 263 329 301
rect 489 285 523 301
rect 603 335 637 351
rect 797 350 831 576
rect 1167 610 1201 923
rect 603 263 637 301
rect 101 125 135 161
rect 101 75 135 91
rect 198 210 232 226
rect -34 34 34 57
rect 198 34 232 176
rect 295 195 329 229
rect 393 216 427 232
rect 603 216 637 229
rect 427 195 637 216
rect 427 182 603 195
rect 393 166 427 182
rect 295 125 329 161
rect 700 316 831 350
rect 928 461 996 544
rect 928 427 945 461
rect 979 427 996 461
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect 1167 433 1201 576
rect 1167 383 1201 399
rect 1389 957 1423 973
rect 1389 683 1423 923
rect 1611 957 1645 973
rect 1611 847 1645 923
rect 1610 831 1645 847
rect 1644 797 1645 831
rect 1610 781 1645 797
rect 1389 433 1423 649
rect 1389 383 1423 399
rect 1611 433 1645 781
rect 1611 383 1645 399
rect 1759 757 1793 1014
rect 1890 1019 1907 1053
rect 1941 1019 1958 1053
rect 2125 1366 2159 1446
rect 2125 1298 2159 1332
rect 2125 1230 2159 1264
rect 2125 1162 2159 1196
rect 2125 1093 2159 1128
rect 2125 1043 2159 1059
rect 2213 1366 2247 1404
rect 2213 1298 2247 1332
rect 2213 1230 2247 1264
rect 2213 1162 2247 1196
rect 2213 1093 2247 1128
rect 2301 1366 2335 1446
rect 2301 1298 2335 1332
rect 2301 1230 2335 1264
rect 2301 1162 2335 1196
rect 2301 1111 2335 1128
rect 2389 1366 2423 1404
rect 2389 1298 2423 1332
rect 2389 1230 2423 1264
rect 2389 1162 2423 1196
rect 2213 1048 2247 1059
rect 2389 1093 2423 1128
rect 2477 1366 2511 1446
rect 2477 1298 2511 1332
rect 2477 1230 2511 1264
rect 2477 1162 2511 1196
rect 2477 1111 2511 1128
rect 2565 1366 2599 1404
rect 2565 1298 2599 1332
rect 2565 1230 2599 1264
rect 2565 1162 2599 1196
rect 2389 1048 2423 1059
rect 2565 1093 2599 1128
rect 2653 1366 2687 1446
rect 2653 1298 2687 1332
rect 2653 1230 2687 1264
rect 2653 1162 2687 1196
rect 2653 1111 2687 1128
rect 2852 1423 2920 1446
rect 2852 1389 2869 1423
rect 2903 1389 2920 1423
rect 2852 1349 2920 1389
rect 2852 1315 2869 1349
rect 2903 1315 2920 1349
rect 2852 1275 2920 1315
rect 2852 1241 2869 1275
rect 2903 1241 2920 1275
rect 2852 1201 2920 1241
rect 2852 1167 2869 1201
rect 2903 1167 2920 1201
rect 2852 1127 2920 1167
rect 2565 1048 2599 1059
rect 2852 1093 2869 1127
rect 2903 1093 2920 1127
rect 2852 1053 2920 1093
rect 1890 979 1958 1019
rect 2213 1014 2755 1048
rect 1890 945 1907 979
rect 1941 945 1958 979
rect 1890 905 1958 945
rect 1890 871 1907 905
rect 1941 871 1958 905
rect 1890 822 1958 871
rect 2129 957 2163 973
rect 700 219 734 316
rect 928 313 996 353
rect 928 279 945 313
rect 979 279 996 313
rect 700 169 734 185
rect 797 263 831 279
rect 797 195 831 229
rect 489 125 523 141
rect 329 91 392 125
rect 426 91 489 125
rect 295 75 329 91
rect 489 75 523 91
rect 603 125 637 161
rect 797 125 831 161
rect 637 91 700 125
rect 734 91 797 125
rect 603 75 637 91
rect 797 75 831 91
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect 928 57 945 91
rect 979 57 996 91
rect 1063 335 1097 351
rect 1257 335 1291 351
rect 1451 335 1485 351
rect 1097 301 1160 335
rect 1194 301 1257 335
rect 1291 301 1354 335
rect 1388 301 1451 335
rect 1063 263 1097 301
rect 1063 195 1097 229
rect 1257 263 1291 301
rect 1451 285 1485 301
rect 1565 335 1599 351
rect 1759 350 1793 723
rect 2129 610 2163 923
rect 1565 263 1599 301
rect 1063 125 1097 161
rect 1063 75 1097 91
rect 1160 210 1194 226
rect 928 34 996 57
rect 1160 34 1194 176
rect 1257 195 1291 229
rect 1355 216 1389 232
rect 1565 216 1599 229
rect 1389 195 1599 216
rect 1389 182 1565 195
rect 1355 166 1389 182
rect 1257 125 1291 161
rect 1662 316 1793 350
rect 1890 461 1958 544
rect 1890 427 1907 461
rect 1941 427 1958 461
rect 1890 387 1958 427
rect 1890 353 1907 387
rect 1941 353 1958 387
rect 2129 433 2163 576
rect 2129 383 2163 399
rect 2351 957 2385 973
rect 2351 536 2385 923
rect 2351 433 2385 502
rect 2351 383 2385 399
rect 2573 957 2607 973
rect 2573 831 2607 923
rect 2573 433 2607 797
rect 2573 383 2607 399
rect 2721 609 2755 1014
rect 2852 1019 2869 1053
rect 2903 1019 2920 1053
rect 3087 1366 3121 1446
rect 3087 1298 3121 1332
rect 3087 1230 3121 1264
rect 3087 1162 3121 1196
rect 3087 1093 3121 1128
rect 3087 1043 3121 1059
rect 3175 1366 3209 1404
rect 3175 1298 3209 1332
rect 3175 1230 3209 1264
rect 3175 1162 3209 1196
rect 3175 1093 3209 1128
rect 3263 1366 3297 1446
rect 3263 1298 3297 1332
rect 3263 1230 3297 1264
rect 3263 1162 3297 1196
rect 3263 1111 3297 1128
rect 3351 1366 3385 1404
rect 3351 1298 3385 1332
rect 3351 1230 3385 1264
rect 3351 1162 3385 1196
rect 3175 1048 3209 1059
rect 3351 1093 3385 1128
rect 3439 1366 3473 1446
rect 3439 1298 3473 1332
rect 3439 1230 3473 1264
rect 3439 1162 3473 1196
rect 3439 1111 3473 1128
rect 3527 1366 3561 1404
rect 3527 1298 3561 1332
rect 3527 1230 3561 1264
rect 3527 1162 3561 1196
rect 3351 1048 3385 1059
rect 3527 1093 3561 1128
rect 3615 1366 3649 1446
rect 3615 1298 3649 1332
rect 3615 1230 3649 1264
rect 3615 1162 3649 1196
rect 3615 1111 3649 1128
rect 3814 1423 3882 1446
rect 3814 1389 3831 1423
rect 3865 1389 3882 1423
rect 3814 1349 3882 1389
rect 3814 1315 3831 1349
rect 3865 1315 3882 1349
rect 3814 1275 3882 1315
rect 3814 1241 3831 1275
rect 3865 1241 3882 1275
rect 3814 1201 3882 1241
rect 3814 1167 3831 1201
rect 3865 1167 3882 1201
rect 3814 1127 3882 1167
rect 3527 1048 3561 1059
rect 3814 1093 3831 1127
rect 3865 1093 3882 1127
rect 3814 1053 3882 1093
rect 2852 979 2920 1019
rect 3175 1014 3717 1048
rect 2852 945 2869 979
rect 2903 945 2920 979
rect 2852 905 2920 945
rect 2852 871 2869 905
rect 2903 871 2920 905
rect 2852 822 2920 871
rect 3091 957 3125 973
rect 1662 219 1696 316
rect 1890 313 1958 353
rect 1890 279 1907 313
rect 1941 279 1958 313
rect 1662 169 1696 185
rect 1759 263 1793 279
rect 1759 195 1793 229
rect 1451 125 1485 141
rect 1291 91 1354 125
rect 1388 91 1451 125
rect 1257 75 1291 91
rect 1451 75 1485 91
rect 1565 125 1599 161
rect 1759 125 1793 161
rect 1599 91 1662 125
rect 1696 91 1759 125
rect 1565 75 1599 91
rect 1759 75 1793 91
rect 1890 239 1958 279
rect 1890 205 1907 239
rect 1941 205 1958 239
rect 1890 165 1958 205
rect 1890 131 1907 165
rect 1941 131 1958 165
rect 1890 91 1958 131
rect 1890 57 1907 91
rect 1941 57 1958 91
rect 2025 335 2059 351
rect 2219 335 2253 351
rect 2413 335 2447 351
rect 2059 301 2122 335
rect 2156 301 2219 335
rect 2253 301 2316 335
rect 2350 301 2413 335
rect 2025 263 2059 301
rect 2025 195 2059 229
rect 2219 263 2253 301
rect 2413 285 2447 301
rect 2527 335 2561 351
rect 2721 350 2755 575
rect 3091 609 3125 923
rect 2527 263 2561 301
rect 2025 125 2059 161
rect 2025 75 2059 91
rect 2122 210 2156 226
rect 1890 34 1958 57
rect 2122 34 2156 176
rect 2219 195 2253 229
rect 2317 216 2351 232
rect 2527 216 2561 229
rect 2351 195 2561 216
rect 2351 182 2527 195
rect 2317 166 2351 182
rect 2219 125 2253 161
rect 2624 316 2755 350
rect 2852 461 2920 544
rect 2852 427 2869 461
rect 2903 427 2920 461
rect 2852 387 2920 427
rect 2852 353 2869 387
rect 2903 353 2920 387
rect 3091 433 3125 575
rect 3091 383 3125 399
rect 3313 957 3347 973
rect 3313 683 3347 923
rect 3313 433 3347 649
rect 3313 383 3347 399
rect 3535 957 3569 973
rect 3535 905 3569 923
rect 3535 433 3569 871
rect 3535 383 3569 399
rect 3683 831 3717 1014
rect 3814 1019 3831 1053
rect 3865 1019 3882 1053
rect 4049 1366 4083 1446
rect 4049 1298 4083 1332
rect 4049 1230 4083 1264
rect 4049 1162 4083 1196
rect 4049 1093 4083 1128
rect 4049 1043 4083 1059
rect 4137 1366 4171 1404
rect 4137 1298 4171 1332
rect 4137 1230 4171 1264
rect 4137 1162 4171 1196
rect 4137 1093 4171 1128
rect 4225 1366 4259 1446
rect 4225 1298 4259 1332
rect 4225 1230 4259 1264
rect 4225 1162 4259 1196
rect 4225 1111 4259 1128
rect 4313 1366 4347 1404
rect 4313 1298 4347 1332
rect 4313 1230 4347 1264
rect 4313 1162 4347 1196
rect 4137 1048 4171 1059
rect 4313 1093 4347 1128
rect 4401 1366 4435 1446
rect 4401 1298 4435 1332
rect 4401 1230 4435 1264
rect 4401 1162 4435 1196
rect 4401 1111 4435 1128
rect 4489 1366 4523 1404
rect 4489 1298 4523 1332
rect 4489 1230 4523 1264
rect 4489 1162 4523 1196
rect 4313 1048 4347 1059
rect 4489 1093 4523 1128
rect 4577 1366 4611 1446
rect 4577 1298 4611 1332
rect 4577 1230 4611 1264
rect 4577 1162 4611 1196
rect 4577 1111 4611 1128
rect 4776 1423 4844 1446
rect 4776 1389 4793 1423
rect 4827 1389 4844 1423
rect 4776 1349 4844 1389
rect 4776 1315 4793 1349
rect 4827 1315 4844 1349
rect 4776 1275 4844 1315
rect 4776 1241 4793 1275
rect 4827 1241 4844 1275
rect 4776 1201 4844 1241
rect 4776 1167 4793 1201
rect 4827 1167 4844 1201
rect 4776 1127 4844 1167
rect 4489 1048 4523 1059
rect 4776 1093 4793 1127
rect 4827 1093 4844 1127
rect 4776 1053 4844 1093
rect 3814 979 3882 1019
rect 4137 1014 4679 1048
rect 3814 945 3831 979
rect 3865 945 3882 979
rect 3814 905 3882 945
rect 3814 871 3831 905
rect 3865 871 3882 905
rect 3814 822 3882 871
rect 4053 957 4087 973
rect 2624 219 2658 316
rect 2852 313 2920 353
rect 2852 279 2869 313
rect 2903 279 2920 313
rect 2624 169 2658 185
rect 2721 263 2755 279
rect 2721 195 2755 229
rect 2413 125 2447 141
rect 2253 91 2316 125
rect 2350 91 2413 125
rect 2219 75 2253 91
rect 2413 75 2447 91
rect 2527 125 2561 161
rect 2721 125 2755 161
rect 2561 91 2624 125
rect 2658 91 2721 125
rect 2527 75 2561 91
rect 2721 75 2755 91
rect 2852 239 2920 279
rect 2852 205 2869 239
rect 2903 205 2920 239
rect 2852 165 2920 205
rect 2852 131 2869 165
rect 2903 131 2920 165
rect 2852 91 2920 131
rect 2852 57 2869 91
rect 2903 57 2920 91
rect 2987 335 3021 351
rect 3181 335 3215 351
rect 3375 335 3409 351
rect 3021 301 3084 335
rect 3118 301 3181 335
rect 3215 301 3278 335
rect 3312 301 3375 335
rect 2987 263 3021 301
rect 2987 195 3021 229
rect 3181 263 3215 301
rect 3375 285 3409 301
rect 3489 335 3523 351
rect 3683 350 3717 797
rect 4053 757 4087 923
rect 3489 263 3523 301
rect 2987 125 3021 161
rect 2987 75 3021 91
rect 3084 210 3118 226
rect 2852 34 2920 57
rect 3084 34 3118 176
rect 3181 195 3215 229
rect 3279 216 3313 232
rect 3489 216 3523 229
rect 3313 195 3523 216
rect 3313 182 3489 195
rect 3279 166 3313 182
rect 3181 125 3215 161
rect 3586 316 3717 350
rect 3814 461 3882 544
rect 3814 427 3831 461
rect 3865 427 3882 461
rect 3814 387 3882 427
rect 3814 353 3831 387
rect 3865 353 3882 387
rect 4053 433 4087 723
rect 4053 383 4087 399
rect 4275 957 4309 973
rect 4275 905 4309 923
rect 4275 433 4309 871
rect 4275 383 4309 399
rect 4497 957 4531 973
rect 4497 757 4531 923
rect 4497 433 4531 723
rect 4497 383 4531 399
rect 4645 683 4679 1014
rect 4776 1019 4793 1053
rect 4827 1019 4844 1053
rect 5011 1366 5045 1446
rect 5011 1298 5045 1332
rect 5011 1230 5045 1264
rect 5011 1162 5045 1196
rect 5011 1093 5045 1128
rect 5011 1043 5045 1059
rect 5099 1366 5133 1404
rect 5099 1298 5133 1332
rect 5099 1230 5133 1264
rect 5099 1162 5133 1196
rect 5099 1093 5133 1128
rect 5187 1366 5221 1446
rect 5187 1298 5221 1332
rect 5187 1230 5221 1264
rect 5187 1162 5221 1196
rect 5187 1111 5221 1128
rect 5275 1366 5309 1404
rect 5275 1298 5309 1332
rect 5275 1230 5309 1264
rect 5275 1162 5309 1196
rect 5099 1048 5133 1059
rect 5275 1093 5309 1128
rect 5363 1366 5397 1446
rect 5363 1298 5397 1332
rect 5363 1230 5397 1264
rect 5363 1162 5397 1196
rect 5363 1111 5397 1128
rect 5451 1366 5485 1404
rect 5451 1298 5485 1332
rect 5451 1230 5485 1264
rect 5451 1162 5485 1196
rect 5275 1048 5309 1059
rect 5451 1093 5485 1128
rect 5539 1366 5573 1446
rect 5539 1298 5573 1332
rect 5539 1230 5573 1264
rect 5539 1162 5573 1196
rect 5539 1111 5573 1128
rect 5738 1423 5806 1446
rect 5738 1389 5755 1423
rect 5789 1389 5806 1423
rect 5738 1349 5806 1389
rect 5738 1315 5755 1349
rect 5789 1315 5806 1349
rect 5738 1275 5806 1315
rect 5738 1241 5755 1275
rect 5789 1241 5806 1275
rect 5738 1201 5806 1241
rect 5738 1167 5755 1201
rect 5789 1167 5806 1201
rect 5738 1127 5806 1167
rect 5451 1048 5485 1059
rect 5738 1093 5755 1127
rect 5789 1093 5806 1127
rect 5738 1053 5806 1093
rect 4776 979 4844 1019
rect 5099 1014 5641 1048
rect 4776 945 4793 979
rect 4827 945 4844 979
rect 4776 905 4844 945
rect 4776 871 4793 905
rect 4827 871 4844 905
rect 4776 822 4844 871
rect 5015 957 5049 973
rect 3586 219 3620 316
rect 3814 313 3882 353
rect 3814 279 3831 313
rect 3865 279 3882 313
rect 3586 169 3620 185
rect 3683 263 3717 279
rect 3683 195 3717 229
rect 3375 125 3409 141
rect 3215 91 3278 125
rect 3312 91 3375 125
rect 3181 75 3215 91
rect 3375 75 3409 91
rect 3489 125 3523 161
rect 3683 125 3717 161
rect 3523 91 3586 125
rect 3620 91 3683 125
rect 3489 75 3523 91
rect 3683 75 3717 91
rect 3814 239 3882 279
rect 3814 205 3831 239
rect 3865 205 3882 239
rect 3814 165 3882 205
rect 3814 131 3831 165
rect 3865 131 3882 165
rect 3814 91 3882 131
rect 3814 57 3831 91
rect 3865 57 3882 91
rect 3949 335 3983 351
rect 4143 335 4177 351
rect 4337 335 4371 351
rect 3983 301 4046 335
rect 4080 301 4143 335
rect 4177 301 4240 335
rect 4274 301 4337 335
rect 3949 263 3983 301
rect 3949 195 3983 229
rect 4143 263 4177 301
rect 4337 285 4371 301
rect 4451 335 4485 351
rect 4645 350 4679 649
rect 5015 683 5049 923
rect 4451 263 4485 301
rect 3949 125 3983 161
rect 3949 75 3983 91
rect 4046 210 4080 226
rect 3814 34 3882 57
rect 4046 34 4080 176
rect 4143 195 4177 229
rect 4241 216 4275 232
rect 4451 216 4485 229
rect 4275 195 4485 216
rect 4275 182 4451 195
rect 4241 166 4275 182
rect 4143 125 4177 161
rect 4548 316 4679 350
rect 4776 461 4844 544
rect 4776 427 4793 461
rect 4827 427 4844 461
rect 4776 387 4844 427
rect 4776 353 4793 387
rect 4827 353 4844 387
rect 5015 433 5049 649
rect 5015 383 5049 399
rect 5237 957 5271 973
rect 5237 535 5271 923
rect 5237 433 5271 501
rect 5237 383 5271 399
rect 5459 957 5493 973
rect 5459 831 5493 923
rect 5459 433 5493 797
rect 5459 383 5493 399
rect 5607 757 5641 1014
rect 5738 1019 5755 1053
rect 5789 1019 5806 1053
rect 5738 979 5806 1019
rect 5738 945 5755 979
rect 5789 945 5806 979
rect 5738 905 5806 945
rect 5738 871 5755 905
rect 5789 871 5806 905
rect 5738 822 5806 871
rect 4548 219 4582 316
rect 4776 313 4844 353
rect 4776 279 4793 313
rect 4827 279 4844 313
rect 4548 169 4582 185
rect 4645 263 4679 279
rect 4645 195 4679 229
rect 4337 125 4371 141
rect 4177 91 4240 125
rect 4274 91 4337 125
rect 4143 75 4177 91
rect 4337 75 4371 91
rect 4451 125 4485 161
rect 4645 125 4679 161
rect 4485 91 4548 125
rect 4582 91 4645 125
rect 4451 75 4485 91
rect 4645 75 4679 91
rect 4776 239 4844 279
rect 4776 205 4793 239
rect 4827 205 4844 239
rect 4776 165 4844 205
rect 4776 131 4793 165
rect 4827 131 4844 165
rect 4776 91 4844 131
rect 4776 57 4793 91
rect 4827 57 4844 91
rect 4911 335 4945 351
rect 5105 335 5139 351
rect 5299 335 5333 351
rect 4945 301 5008 335
rect 5042 301 5105 335
rect 5139 301 5202 335
rect 5236 301 5299 335
rect 4911 263 4945 301
rect 4911 195 4945 229
rect 5105 263 5139 301
rect 5299 285 5333 301
rect 5413 335 5447 351
rect 5607 350 5641 723
rect 5413 263 5447 301
rect 4911 125 4945 161
rect 4911 75 4945 91
rect 5008 210 5042 226
rect 4776 34 4844 57
rect 5008 34 5042 176
rect 5105 195 5139 229
rect 5203 216 5237 232
rect 5413 216 5447 229
rect 5237 195 5447 216
rect 5237 182 5413 195
rect 5203 166 5237 182
rect 5105 125 5139 161
rect 5510 316 5641 350
rect 5738 461 5806 544
rect 5738 427 5755 461
rect 5789 427 5806 461
rect 5738 387 5806 427
rect 5738 353 5755 387
rect 5789 353 5806 387
rect 5510 219 5544 316
rect 5738 313 5806 353
rect 5738 279 5755 313
rect 5789 279 5806 313
rect 5510 169 5544 185
rect 5607 263 5641 279
rect 5607 195 5641 229
rect 5299 125 5333 141
rect 5139 91 5202 125
rect 5236 91 5299 125
rect 5105 75 5139 91
rect 5299 75 5333 91
rect 5413 125 5447 161
rect 5607 125 5641 161
rect 5447 91 5510 125
rect 5544 91 5607 125
rect 5413 75 5447 91
rect 5607 75 5641 91
rect 5738 239 5806 279
rect 5738 205 5755 239
rect 5789 205 5806 239
rect 5738 165 5806 205
rect 5738 131 5755 165
rect 5789 131 5806 165
rect 5738 91 5806 131
rect 5738 57 5755 91
rect 5789 57 5806 91
rect 5738 34 5806 57
rect -34 17 5806 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5806 17
rect -34 -34 5806 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5163 1463 5197 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5533 1463 5567 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 427 871 461 905
rect 649 723 683 757
rect 797 576 831 610
rect 1167 576 1201 610
rect 1610 797 1644 831
rect 1389 649 1423 683
rect 1759 723 1793 757
rect 2129 576 2163 610
rect 2351 502 2385 536
rect 2573 797 2607 831
rect 2721 575 2755 609
rect 3091 575 3125 609
rect 3313 649 3347 683
rect 3535 871 3569 905
rect 3683 797 3717 831
rect 4053 723 4087 757
rect 4275 871 4309 905
rect 4497 723 4531 757
rect 4645 649 4679 683
rect 5015 649 5049 683
rect 5237 501 5271 535
rect 5459 797 5493 831
rect 5607 723 5641 757
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5163 -17 5197 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5533 -17 5567 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
<< metal1 >>
rect -34 1497 5806 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5806 1497
rect -34 1446 5806 1463
rect 421 905 467 911
rect 3529 905 3575 911
rect 4269 905 4315 911
rect 415 871 427 905
rect 461 871 3535 905
rect 3569 871 4275 905
rect 4309 871 4321 905
rect 421 865 467 871
rect 3529 865 3575 871
rect 4269 865 4315 871
rect 1604 831 1650 837
rect 2567 831 2613 837
rect 3677 831 3723 837
rect 5453 831 5499 837
rect 1598 797 1610 831
rect 1644 797 2573 831
rect 2607 797 3683 831
rect 3717 797 5459 831
rect 5493 797 5505 831
rect 1604 791 1650 797
rect 2567 791 2613 797
rect 3677 791 3723 797
rect 5453 791 5499 797
rect 643 757 689 763
rect 1753 757 1799 763
rect 4047 757 4093 763
rect 4491 757 4537 763
rect 5601 757 5647 763
rect 637 723 649 757
rect 683 723 1759 757
rect 1793 723 4053 757
rect 4087 723 4099 757
rect 4485 723 4497 757
rect 4531 723 5607 757
rect 5641 723 5653 757
rect 643 717 689 723
rect 1753 717 1799 723
rect 4047 717 4093 723
rect 4491 717 4537 723
rect 5601 717 5647 723
rect 1383 683 1429 689
rect 3307 683 3353 689
rect 4639 683 4685 689
rect 5009 683 5055 689
rect 1377 649 1389 683
rect 1423 649 3313 683
rect 3347 649 3359 683
rect 4633 649 4645 683
rect 4679 649 5015 683
rect 5049 649 5061 683
rect 1383 643 1429 649
rect 3307 643 3353 649
rect 4639 643 4685 649
rect 5009 643 5055 649
rect 791 610 837 616
rect 1161 610 1207 616
rect 2123 610 2169 616
rect 785 576 797 610
rect 831 576 1167 610
rect 1201 576 2129 610
rect 2163 576 2175 610
rect 2715 609 2761 615
rect 3085 609 3131 615
rect 791 570 837 576
rect 1161 570 1207 576
rect 2123 570 2169 576
rect 2709 575 2721 609
rect 2755 575 3091 609
rect 3125 575 3137 609
rect 2715 569 2761 575
rect 3085 569 3131 575
rect 2345 536 2391 542
rect 2339 502 2351 536
rect 2385 535 2421 536
rect 5231 535 5277 541
rect 2385 502 5237 535
rect 2345 496 2391 502
rect 2421 501 5237 502
rect 5271 501 5283 535
rect 5231 495 5277 501
rect -34 17 5806 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5806 17
rect -34 -34 5806 -17
<< labels >>
rlabel metal1 4645 649 4679 683 1 QN
port 1 n
rlabel metal1 205 575 239 609 1 D
port 2 n
rlabel metal1 1389 649 1423 683 1 CLK
port 3 n
rlabel metal1 427 871 461 905 1 RN
port 4 n
rlabel metal1 2351 501 2385 535 1 SN
port 5 n
rlabel metal1 4645 575 4679 609 1 QN
port 6 n
rlabel metal1 4645 427 4679 461 1 QN
port 7 n
rlabel metal1 4645 871 4679 905 1 QN
port 8 n
rlabel metal1 4645 945 4679 979 1 QN
port 9 n
rlabel metal1 5015 575 5049 609 1 QN
port 10 n
rlabel metal1 5015 649 5049 683 1 QN
port 11 n
rlabel metal1 5015 427 5049 461 1 QN
port 12 n
rlabel metal1 5015 871 5049 905 1 QN
port 13 n
rlabel metal1 205 649 239 683 1 D
port 14 n
rlabel metal1 205 723 239 757 1 D
port 15 n
rlabel metal1 205 797 239 831 1 D
port 16 n
rlabel metal1 205 871 239 905 1 D
port 17 n
rlabel metal1 205 501 239 535 1 D
port 18 n
rlabel metal1 1389 501 1423 535 1 CLK
port 19 n
rlabel metal1 1389 797 1423 831 1 CLK
port 20 n
rlabel metal1 3313 649 3347 683 1 CLK
port 21 n
rlabel metal1 3313 575 3347 609 1 CLK
port 22 n
rlabel metal1 427 797 461 831 1 RN
port 23 n
rlabel metal1 427 723 461 757 1 RN
port 24 n
rlabel metal1 427 649 461 683 1 RN
port 25 n
rlabel metal1 427 575 461 609 1 RN
port 26 n
rlabel metal1 427 501 461 535 1 RN
port 27 n
rlabel metal1 3535 649 3569 683 1 RN
port 28 n
rlabel metal1 3535 575 3569 609 1 RN
port 29 n
rlabel metal1 3535 871 3569 905 1 RN
port 30 n
rlabel metal1 4275 575 4309 609 1 RN
port 31 n
rlabel metal1 4275 649 4309 683 1 RN
port 32 n
rlabel metal1 4275 723 4309 757 1 RN
port 33 n
rlabel metal1 4275 871 4309 905 1 RN
port 34 n
rlabel metal1 -34 1446 5806 1514 1 VPWR
port 35 n
rlabel metal1 -34 -34 5806 34 1 VGND
port 36 n
rlabel nwell 57 1463 91 1497 1 VPB
port 37 n
rlabel metal1 57 -17 91 17 1 VNB
port 38 n
<< end >>
