// File: nor3x1_pcell.spi.NOR3X1_PCELL.pxi
// Created: Tue Oct 15 15:59:36 2024
// 
simulator lang=spectre
x_PM_NOR3X1_PCELL\%noxref_1 ( N_noxref_1_c_3_p N_noxref_1_c_4_p \
 N_noxref_1_c_11_p N_noxref_1_c_15_p N_noxref_1_c_19_p N_noxref_1_c_23_p \
 N_noxref_1_c_27_p N_noxref_1_c_2_p N_noxref_1_c_1_p N_noxref_1_M0_noxref_s )  \
 PM_NOR3X1_PCELL\%noxref_1
x_PM_NOR3X1_PCELL\%noxref_2 ( N_noxref_2_c_71_p N_noxref_2_c_57_p \
 N_noxref_2_c_52_n N_noxref_2_c_53_n N_noxref_2_M3_noxref_d )  \
 PM_NOR3X1_PCELL\%noxref_2
x_PM_NOR3X1_PCELL\%noxref_3 ( N_noxref_3_c_94_n N_noxref_3_c_106_n \
 N_noxref_3_M0_noxref_g N_noxref_3_M3_noxref_g N_noxref_3_M4_noxref_g \
 N_noxref_3_c_97_n N_noxref_3_c_124_p N_noxref_3_c_125_p N_noxref_3_c_99_n \
 N_noxref_3_c_101_n N_noxref_3_c_156_p N_noxref_3_c_115_p N_noxref_3_c_102_n \
 N_noxref_3_c_104_n N_noxref_3_c_113_n )  PM_NOR3X1_PCELL\%noxref_3
x_PM_NOR3X1_PCELL\%noxref_4 ( N_noxref_4_c_169_n N_noxref_4_c_159_n \
 N_noxref_4_M1_noxref_g N_noxref_4_M5_noxref_g N_noxref_4_M6_noxref_g \
 N_noxref_4_c_160_n N_noxref_4_c_179_n N_noxref_4_c_182_n N_noxref_4_c_217_p \
 N_noxref_4_c_162_n N_noxref_4_c_163_n N_noxref_4_c_164_n N_noxref_4_c_186_n \
 N_noxref_4_c_187_n N_noxref_4_c_189_n N_noxref_4_c_190_n )  \
 PM_NOR3X1_PCELL\%noxref_4
x_PM_NOR3X1_PCELL\%noxref_5 ( N_noxref_5_c_239_n N_noxref_5_c_242_n \
 N_noxref_5_c_243_n N_noxref_5_c_244_n N_noxref_5_M3_noxref_s \
 N_noxref_5_M4_noxref_d N_noxref_5_M6_noxref_d )  PM_NOR3X1_PCELL\%noxref_5
x_PM_NOR3X1_PCELL\%noxref_6 ( N_noxref_6_c_282_n N_noxref_6_M2_noxref_g \
 N_noxref_6_M7_noxref_g N_noxref_6_M8_noxref_g N_noxref_6_c_284_n \
 N_noxref_6_c_303_n N_noxref_6_c_305_n N_noxref_6_c_307_n N_noxref_6_c_286_n \
 N_noxref_6_c_287_n N_noxref_6_c_288_n N_noxref_6_c_310_n N_noxref_6_c_294_n \
 N_noxref_6_c_290_n N_noxref_6_c_313_n )  PM_NOR3X1_PCELL\%noxref_6
x_PM_NOR3X1_PCELL\%noxref_7 ( N_noxref_7_c_349_n N_noxref_7_c_374_n \
 N_noxref_7_c_353_n N_noxref_7_c_357_n N_noxref_7_c_371_n N_noxref_7_c_412_n \
 N_noxref_7_c_398_n N_noxref_7_M0_noxref_d N_noxref_7_M1_noxref_d \
 N_noxref_7_M2_noxref_d N_noxref_7_M7_noxref_d )  PM_NOR3X1_PCELL\%noxref_7
x_PM_NOR3X1_PCELL\%noxref_8 ( N_noxref_8_c_432_n N_noxref_8_c_433_n \
 N_noxref_8_c_434_n N_noxref_8_c_435_n N_noxref_8_M5_noxref_d \
 N_noxref_8_M7_noxref_s N_noxref_8_M8_noxref_d )  PM_NOR3X1_PCELL\%noxref_8
cc_1 ( N_noxref_1_c_1_p N_noxref_2_c_52_n ) capacitor c=0.00989031f //x=0.695 \
 //y=0 //x2=0.74 //y2=7.4
cc_2 ( N_noxref_1_c_2_p N_noxref_2_c_53_n ) capacitor c=0.00989031f //x=4.07 \
 //y=0 //x2=4.07 //y2=7.4
cc_3 ( N_noxref_1_c_3_p N_noxref_3_c_94_n ) capacitor c=6.7762e-19 //x=4.07 \
 //y=0 //x2=1.11 //y2=2.08
cc_4 ( N_noxref_1_c_4_p N_noxref_3_c_94_n ) capacitor c=0.00136072f //x=1.095 \
 //y=0.53 //x2=1.11 //y2=2.08
cc_5 ( N_noxref_1_c_1_p N_noxref_3_c_94_n ) capacitor c=0.0176887f //x=0.695 \
 //y=0 //x2=1.11 //y2=2.08
cc_6 ( N_noxref_1_c_4_p N_noxref_3_c_97_n ) capacitor c=0.0122371f //x=1.095 \
 //y=0.53 //x2=0.915 //y2=0.905
cc_7 ( N_noxref_1_M0_noxref_s N_noxref_3_c_97_n ) capacitor c=0.0318083f \
 //x=0.56 //y=0.365 //x2=0.915 //y2=0.905
cc_8 ( N_noxref_1_c_4_p N_noxref_3_c_99_n ) capacitor c=2.1838e-19 //x=1.095 \
 //y=0.53 //x2=0.915 //y2=1.915
cc_9 ( N_noxref_1_c_1_p N_noxref_3_c_99_n ) capacitor c=0.0198857f //x=0.695 \
 //y=0 //x2=0.915 //y2=1.915
cc_10 ( N_noxref_1_M0_noxref_s N_noxref_3_c_101_n ) capacitor c=0.00474433f \
 //x=0.56 //y=0.365 //x2=1.29 //y2=0.75
cc_11 ( N_noxref_1_c_11_p N_noxref_3_c_102_n ) capacitor c=0.0113089f //x=1.58 \
 //y=0.53 //x2=1.445 //y2=0.905
cc_12 ( N_noxref_1_M0_noxref_s N_noxref_3_c_102_n ) capacitor c=0.00514143f \
 //x=0.56 //y=0.365 //x2=1.445 //y2=0.905
cc_13 ( N_noxref_1_M0_noxref_s N_noxref_3_c_104_n ) capacitor c=8.33128e-19 \
 //x=0.56 //y=0.365 //x2=1.445 //y2=1.25
cc_14 ( N_noxref_1_c_1_p N_noxref_4_c_159_n ) capacitor c=9.2064e-19 //x=0.695 \
 //y=0 //x2=1.85 //y2=2.08
cc_15 ( N_noxref_1_c_15_p N_noxref_4_c_160_n ) capacitor c=0.01113f //x=2.065 \
 //y=0.53 //x2=1.885 //y2=0.905
cc_16 ( N_noxref_1_M0_noxref_s N_noxref_4_c_160_n ) capacitor c=0.00590563f \
 //x=0.56 //y=0.365 //x2=1.885 //y2=0.905
cc_17 ( N_noxref_1_M0_noxref_s N_noxref_4_c_162_n ) capacitor c=0.00481727f \
 //x=0.56 //y=0.365 //x2=2.26 //y2=0.75
cc_18 ( N_noxref_1_M0_noxref_s N_noxref_4_c_163_n ) capacitor c=8.38882e-19 \
 //x=0.56 //y=0.365 //x2=2.26 //y2=1.405
cc_19 ( N_noxref_1_c_19_p N_noxref_4_c_164_n ) capacitor c=0.0113819f //x=2.55 \
 //y=0.53 //x2=2.415 //y2=0.905
cc_20 ( N_noxref_1_M0_noxref_s N_noxref_4_c_164_n ) capacitor c=0.00513762f \
 //x=0.56 //y=0.365 //x2=2.415 //y2=0.905
cc_21 ( N_noxref_1_c_3_p N_noxref_6_c_282_n ) capacitor c=3.7166e-19 //x=4.07 \
 //y=0 //x2=2.96 //y2=2.08
cc_22 ( N_noxref_1_c_2_p N_noxref_6_c_282_n ) capacitor c=5.99091e-19 //x=4.07 \
 //y=0 //x2=2.96 //y2=2.08
cc_23 ( N_noxref_1_c_23_p N_noxref_6_c_284_n ) capacitor c=0.0108358f \
 //x=3.035 //y=0.53 //x2=2.855 //y2=0.905
cc_24 ( N_noxref_1_M0_noxref_s N_noxref_6_c_284_n ) capacitor c=0.00590563f \
 //x=0.56 //y=0.365 //x2=2.855 //y2=0.905
cc_25 ( N_noxref_1_M0_noxref_s N_noxref_6_c_286_n ) capacitor c=0.00452306f \
 //x=0.56 //y=0.365 //x2=3.23 //y2=0.75
cc_26 ( N_noxref_1_M0_noxref_s N_noxref_6_c_287_n ) capacitor c=0.00316186f \
 //x=0.56 //y=0.365 //x2=3.23 //y2=1.405
cc_27 ( N_noxref_1_c_27_p N_noxref_6_c_288_n ) capacitor c=0.0110876f //x=3.52 \
 //y=0.53 //x2=3.385 //y2=0.905
cc_28 ( N_noxref_1_M0_noxref_s N_noxref_6_c_288_n ) capacitor c=0.0132184f \
 //x=0.56 //y=0.365 //x2=3.385 //y2=0.905
cc_29 ( N_noxref_1_c_23_p N_noxref_6_c_290_n ) capacitor c=2.26024e-19 \
 //x=3.035 //y=0.53 //x2=2.855 //y2=2.08
cc_30 ( N_noxref_1_c_3_p N_noxref_7_c_349_n ) capacitor c=0.00359057f //x=4.07 \
 //y=0 //x2=2.065 //y2=1.655
cc_31 ( N_noxref_1_c_11_p N_noxref_7_c_349_n ) capacitor c=0.00381844f \
 //x=1.58 //y=0.53 //x2=2.065 //y2=1.655
cc_32 ( N_noxref_1_c_15_p N_noxref_7_c_349_n ) capacitor c=0.00323369f \
 //x=2.065 //y=0.53 //x2=2.065 //y2=1.655
cc_33 ( N_noxref_1_M0_noxref_s N_noxref_7_c_349_n ) capacitor c=0.0173679f \
 //x=0.56 //y=0.365 //x2=2.065 //y2=1.655
cc_34 ( N_noxref_1_c_3_p N_noxref_7_c_353_n ) capacitor c=0.00410159f //x=4.07 \
 //y=0 //x2=3.035 //y2=1.655
cc_35 ( N_noxref_1_c_19_p N_noxref_7_c_353_n ) capacitor c=0.00381844f \
 //x=2.55 //y=0.53 //x2=3.035 //y2=1.655
cc_36 ( N_noxref_1_c_23_p N_noxref_7_c_353_n ) capacitor c=0.00324961f \
 //x=3.035 //y=0.53 //x2=3.035 //y2=1.655
cc_37 ( N_noxref_1_M0_noxref_s N_noxref_7_c_353_n ) capacitor c=0.0175442f \
 //x=0.56 //y=0.365 //x2=3.035 //y2=1.655
cc_38 ( N_noxref_1_c_3_p N_noxref_7_c_357_n ) capacitor c=0.0045676f //x=4.07 \
 //y=0 //x2=3.615 //y2=1.655
cc_39 ( N_noxref_1_c_27_p N_noxref_7_c_357_n ) capacitor c=0.0047981f //x=3.52 \
 //y=0.53 //x2=3.615 //y2=1.655
cc_40 ( N_noxref_1_c_2_p N_noxref_7_c_357_n ) capacitor c=0.0296404f //x=4.07 \
 //y=0 //x2=3.615 //y2=1.655
cc_41 ( N_noxref_1_M0_noxref_s N_noxref_7_c_357_n ) capacitor c=0.0198878f \
 //x=0.56 //y=0.365 //x2=3.615 //y2=1.655
cc_42 ( N_noxref_1_c_3_p N_noxref_7_M0_noxref_d ) capacitor c=0.00175924f \
 //x=4.07 //y=0 //x2=0.99 //y2=0.905
cc_43 ( N_noxref_1_c_2_p N_noxref_7_M0_noxref_d ) capacitor c=2.31043e-19 \
 //x=4.07 //y=0 //x2=0.99 //y2=0.905
cc_44 ( N_noxref_1_c_1_p N_noxref_7_M0_noxref_d ) capacitor c=0.00419389f \
 //x=0.695 //y=0 //x2=0.99 //y2=0.905
cc_45 ( N_noxref_1_M0_noxref_s N_noxref_7_M0_noxref_d ) capacitor c=0.0775691f \
 //x=0.56 //y=0.365 //x2=0.99 //y2=0.905
cc_46 ( N_noxref_1_c_3_p N_noxref_7_M1_noxref_d ) capacitor c=0.00195394f \
 //x=4.07 //y=0 //x2=1.96 //y2=0.905
cc_47 ( N_noxref_1_c_2_p N_noxref_7_M1_noxref_d ) capacitor c=2.31043e-19 \
 //x=4.07 //y=0 //x2=1.96 //y2=0.905
cc_48 ( N_noxref_1_M0_noxref_s N_noxref_7_M1_noxref_d ) capacitor c=0.0610444f \
 //x=0.56 //y=0.365 //x2=1.96 //y2=0.905
cc_49 ( N_noxref_1_c_3_p N_noxref_7_M2_noxref_d ) capacitor c=0.00193447f \
 //x=4.07 //y=0 //x2=2.93 //y2=0.905
cc_50 ( N_noxref_1_c_2_p N_noxref_7_M2_noxref_d ) capacitor c=0.00397791f \
 //x=4.07 //y=0 //x2=2.93 //y2=0.905
cc_51 ( N_noxref_1_M0_noxref_s N_noxref_7_M2_noxref_d ) capacitor c=0.0604189f \
 //x=0.56 //y=0.365 //x2=2.93 //y2=0.905
cc_52 ( N_noxref_2_c_52_n N_noxref_3_c_94_n ) capacitor c=0.0104719f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_53 ( N_noxref_2_c_52_n N_noxref_3_c_106_n ) capacitor c=0.008636f //x=0.74 \
 //y=7.4 //x2=0.955 //y2=4.705
cc_54 ( N_noxref_2_M3_noxref_d N_noxref_3_c_106_n ) capacitor c=2.85008e-19 \
 //x=1.085 //y=5.025 //x2=0.955 //y2=4.705
cc_55 ( N_noxref_2_c_57_p N_noxref_3_M3_noxref_g ) capacitor c=0.0067918f \
 //x=1.145 //y=7.4 //x2=1.01 //y2=6.025
cc_56 ( N_noxref_2_c_52_n N_noxref_3_M3_noxref_g ) capacitor c=0.0241979f \
 //x=0.74 //y=7.4 //x2=1.01 //y2=6.025
cc_57 ( N_noxref_2_M3_noxref_d N_noxref_3_M3_noxref_g ) capacitor c=0.0156786f \
 //x=1.085 //y=5.025 //x2=1.01 //y2=6.025
cc_58 ( N_noxref_2_c_53_n N_noxref_3_M4_noxref_g ) capacitor c=0.00678153f \
 //x=4.07 //y=7.4 //x2=1.45 //y2=6.025
cc_59 ( N_noxref_2_M3_noxref_d N_noxref_3_M4_noxref_g ) capacitor c=0.019067f \
 //x=1.085 //y=5.025 //x2=1.45 //y2=6.025
cc_60 ( N_noxref_2_c_52_n N_noxref_3_c_113_n ) capacitor c=0.00890932f \
 //x=0.74 //y=7.4 //x2=0.955 //y2=4.705
cc_61 ( N_noxref_2_c_52_n N_noxref_4_c_159_n ) capacitor c=7.02327e-19 \
 //x=0.74 //y=7.4 //x2=1.85 //y2=2.08
cc_62 ( N_noxref_2_c_53_n N_noxref_4_M5_noxref_g ) capacitor c=0.00513565f \
 //x=4.07 //y=7.4 //x2=1.89 //y2=6.025
cc_63 ( N_noxref_2_c_53_n N_noxref_4_M6_noxref_g ) capacitor c=0.00512552f \
 //x=4.07 //y=7.4 //x2=2.33 //y2=6.025
cc_64 ( N_noxref_2_c_57_p N_noxref_5_c_239_n ) capacitor c=5.81484e-19 \
 //x=1.145 //y=7.4 //x2=1.585 //y2=5.21
cc_65 ( N_noxref_2_c_53_n N_noxref_5_c_239_n ) capacitor c=5.81484e-19 \
 //x=4.07 //y=7.4 //x2=1.585 //y2=5.21
cc_66 ( N_noxref_2_M3_noxref_d N_noxref_5_c_239_n ) capacitor c=0.0132432f \
 //x=1.085 //y=5.025 //x2=1.585 //y2=5.21
cc_67 ( N_noxref_2_c_52_n N_noxref_5_c_242_n ) capacitor c=0.0679103f //x=0.74 \
 //y=7.4 //x2=0.875 //y2=5.21
cc_68 ( N_noxref_2_c_53_n N_noxref_5_c_243_n ) capacitor c=0.00436083f \
 //x=4.07 //y=7.4 //x2=2.465 //y2=6.91
cc_69 ( N_noxref_2_c_71_p N_noxref_5_c_244_n ) capacitor c=0.0370274f //x=4.07 \
 //y=7.4 //x2=1.755 //y2=6.91
cc_70 ( N_noxref_2_c_53_n N_noxref_5_c_244_n ) capacitor c=0.059877f //x=4.07 \
 //y=7.4 //x2=1.755 //y2=6.91
cc_71 ( N_noxref_2_c_71_p N_noxref_5_M3_noxref_s ) capacitor c=0.00726388f \
 //x=4.07 //y=7.4 //x2=0.655 //y2=5.025
cc_72 ( N_noxref_2_c_57_p N_noxref_5_M3_noxref_s ) capacitor c=0.0141117f \
 //x=1.145 //y=7.4 //x2=0.655 //y2=5.025
cc_73 ( N_noxref_2_c_53_n N_noxref_5_M3_noxref_s ) capacitor c=0.00138926f \
 //x=4.07 //y=7.4 //x2=0.655 //y2=5.025
cc_74 ( N_noxref_2_M3_noxref_d N_noxref_5_M3_noxref_s ) capacitor c=0.0667777f \
 //x=1.085 //y=5.025 //x2=0.655 //y2=5.025
cc_75 ( N_noxref_2_c_52_n N_noxref_5_M4_noxref_d ) capacitor c=8.88629e-19 \
 //x=0.74 //y=7.4 //x2=1.525 //y2=5.025
cc_76 ( N_noxref_2_M3_noxref_d N_noxref_5_M4_noxref_d ) capacitor c=0.0659925f \
 //x=1.085 //y=5.025 //x2=1.525 //y2=5.025
cc_77 ( N_noxref_2_M3_noxref_d N_noxref_5_M6_noxref_d ) capacitor \
 c=0.00107819f //x=1.085 //y=5.025 //x2=2.405 //y2=5.025
cc_78 ( N_noxref_2_c_53_n N_noxref_6_c_282_n ) capacitor c=7.00707e-19 \
 //x=4.07 //y=7.4 //x2=2.96 //y2=2.08
cc_79 ( N_noxref_2_c_53_n N_noxref_6_M7_noxref_g ) capacitor c=0.00512552f \
 //x=4.07 //y=7.4 //x2=3.37 //y2=6.025
cc_80 ( N_noxref_2_c_53_n N_noxref_6_M8_noxref_g ) capacitor c=0.0109813f \
 //x=4.07 //y=7.4 //x2=3.81 //y2=6.025
cc_81 ( N_noxref_2_c_53_n N_noxref_6_c_294_n ) capacitor c=0.0268396f //x=4.07 \
 //y=7.4 //x2=3.735 //y2=4.795
cc_82 ( N_noxref_2_c_53_n N_noxref_7_c_371_n ) capacitor c=0.0263915f //x=4.07 \
 //y=7.4 //x2=3.7 //y2=5.125
cc_83 ( N_noxref_2_c_53_n N_noxref_7_M7_noxref_d ) capacitor c=0.00991513f \
 //x=4.07 //y=7.4 //x2=3.445 //y2=5.025
cc_84 ( N_noxref_2_c_53_n N_noxref_8_c_432_n ) capacitor c=0.00565054f \
 //x=4.07 //y=7.4 //x2=3.065 //y2=5.21
cc_85 ( N_noxref_2_c_52_n N_noxref_8_c_433_n ) capacitor c=9.33216e-19 \
 //x=0.74 //y=7.4 //x2=2.195 //y2=5.21
cc_86 ( N_noxref_2_c_53_n N_noxref_8_c_434_n ) capacitor c=0.00356149f \
 //x=4.07 //y=7.4 //x2=3.945 //y2=6.91
cc_87 ( N_noxref_2_c_71_p N_noxref_8_c_435_n ) capacitor c=0.0370274f //x=4.07 \
 //y=7.4 //x2=3.235 //y2=6.91
cc_88 ( N_noxref_2_c_53_n N_noxref_8_c_435_n ) capacitor c=0.0597427f //x=4.07 \
 //y=7.4 //x2=3.235 //y2=6.91
cc_89 ( N_noxref_2_M3_noxref_d N_noxref_8_c_435_n ) capacitor c=9.25055e-19 \
 //x=1.085 //y=5.025 //x2=3.235 //y2=6.91
cc_90 ( N_noxref_2_M3_noxref_d N_noxref_8_M5_noxref_d ) capacitor \
 c=0.00561178f //x=1.085 //y=5.025 //x2=1.965 //y2=5.025
cc_91 ( N_noxref_2_c_53_n N_noxref_8_M8_noxref_d ) capacitor c=0.0528345f \
 //x=4.07 //y=7.4 //x2=3.885 //y2=5.025
cc_92 ( N_noxref_3_c_106_n N_noxref_4_c_169_n ) capacitor c=0.0482889f \
 //x=0.955 //y=4.705 //x2=1.85 //y2=4.54
cc_93 ( N_noxref_3_c_115_p N_noxref_4_c_169_n ) capacitor c=0.00146509f \
 //x=1.375 //y=4.795 //x2=1.85 //y2=4.54
cc_94 ( N_noxref_3_c_113_n N_noxref_4_c_169_n ) capacitor c=0.00112871f \
 //x=0.955 //y=4.705 //x2=1.85 //y2=4.54
cc_95 ( N_noxref_3_c_94_n N_noxref_4_c_159_n ) capacitor c=0.0455438f //x=1.11 \
 //y=2.08 //x2=1.85 //y2=2.08
cc_96 ( N_noxref_3_c_99_n N_noxref_4_c_159_n ) capacitor c=0.00308814f \
 //x=0.915 //y=1.915 //x2=1.85 //y2=2.08
cc_97 ( N_noxref_3_M3_noxref_g N_noxref_4_M5_noxref_g ) capacitor c=0.0100243f \
 //x=1.01 //y=6.025 //x2=1.89 //y2=6.025
cc_98 ( N_noxref_3_M4_noxref_g N_noxref_4_M5_noxref_g ) capacitor c=0.107798f \
 //x=1.45 //y=6.025 //x2=1.89 //y2=6.025
cc_99 ( N_noxref_3_M4_noxref_g N_noxref_4_M6_noxref_g ) capacitor c=0.0094155f \
 //x=1.45 //y=6.025 //x2=2.33 //y2=6.025
cc_100 ( N_noxref_3_c_97_n N_noxref_4_c_160_n ) capacitor c=0.00125788f \
 //x=0.915 //y=0.905 //x2=1.885 //y2=0.905
cc_101 ( N_noxref_3_c_102_n N_noxref_4_c_160_n ) capacitor c=0.0126654f \
 //x=1.445 //y=0.905 //x2=1.885 //y2=0.905
cc_102 ( N_noxref_3_c_124_p N_noxref_4_c_179_n ) capacitor c=0.00148539f \
 //x=0.915 //y=1.25 //x2=1.885 //y2=1.255
cc_103 ( N_noxref_3_c_125_p N_noxref_4_c_179_n ) capacitor c=0.00105591f \
 //x=0.915 //y=1.56 //x2=1.885 //y2=1.255
cc_104 ( N_noxref_3_c_104_n N_noxref_4_c_179_n ) capacitor c=0.0126654f \
 //x=1.445 //y=1.25 //x2=1.885 //y2=1.255
cc_105 ( N_noxref_3_c_125_p N_noxref_4_c_182_n ) capacitor c=0.00109549f \
 //x=0.915 //y=1.56 //x2=1.885 //y2=1.56
cc_106 ( N_noxref_3_c_104_n N_noxref_4_c_182_n ) capacitor c=0.00886999f \
 //x=1.445 //y=1.25 //x2=1.885 //y2=1.56
cc_107 ( N_noxref_3_c_104_n N_noxref_4_c_163_n ) capacitor c=0.00123863f \
 //x=1.445 //y=1.25 //x2=2.26 //y2=1.405
cc_108 ( N_noxref_3_c_102_n N_noxref_4_c_164_n ) capacitor c=0.00132934f \
 //x=1.445 //y=0.905 //x2=2.415 //y2=0.905
cc_109 ( N_noxref_3_c_104_n N_noxref_4_c_186_n ) capacitor c=0.00150734f \
 //x=1.445 //y=1.25 //x2=2.415 //y2=1.255
cc_110 ( N_noxref_3_c_94_n N_noxref_4_c_187_n ) capacitor c=0.00307062f \
 //x=1.11 //y=2.08 //x2=1.85 //y2=2.08
cc_111 ( N_noxref_3_c_99_n N_noxref_4_c_187_n ) capacitor c=0.0176046f \
 //x=0.915 //y=1.915 //x2=1.85 //y2=2.08
cc_112 ( N_noxref_3_c_99_n N_noxref_4_c_189_n ) capacitor c=0.00577193f \
 //x=0.915 //y=1.915 //x2=1.85 //y2=1.915
cc_113 ( N_noxref_3_c_106_n N_noxref_4_c_190_n ) capacitor c=0.00336963f \
 //x=0.955 //y=4.705 //x2=1.885 //y2=4.705
cc_114 ( N_noxref_3_c_115_p N_noxref_4_c_190_n ) capacitor c=0.0197705f \
 //x=1.375 //y=4.795 //x2=1.885 //y2=4.705
cc_115 ( N_noxref_3_c_113_n N_noxref_4_c_190_n ) capacitor c=0.00546725f \
 //x=0.955 //y=4.705 //x2=1.885 //y2=4.705
cc_116 ( N_noxref_3_c_106_n N_noxref_5_c_239_n ) capacitor c=0.00630079f \
 //x=0.955 //y=4.705 //x2=1.585 //y2=5.21
cc_117 ( N_noxref_3_M3_noxref_g N_noxref_5_c_239_n ) capacitor c=0.0182669f \
 //x=1.01 //y=6.025 //x2=1.585 //y2=5.21
cc_118 ( N_noxref_3_M4_noxref_g N_noxref_5_c_239_n ) capacitor c=0.0204082f \
 //x=1.45 //y=6.025 //x2=1.585 //y2=5.21
cc_119 ( N_noxref_3_c_115_p N_noxref_5_c_239_n ) capacitor c=0.00365818f \
 //x=1.375 //y=4.795 //x2=1.585 //y2=5.21
cc_120 ( N_noxref_3_c_113_n N_noxref_5_c_239_n ) capacitor c=0.0017421f \
 //x=0.955 //y=4.705 //x2=1.585 //y2=5.21
cc_121 ( N_noxref_3_c_106_n N_noxref_5_c_242_n ) capacitor c=0.0118415f \
 //x=0.955 //y=4.705 //x2=0.875 //y2=5.21
cc_122 ( N_noxref_3_c_113_n N_noxref_5_c_242_n ) capacitor c=0.00613395f \
 //x=0.955 //y=4.705 //x2=0.875 //y2=5.21
cc_123 ( N_noxref_3_M3_noxref_g N_noxref_5_M3_noxref_s ) capacitor \
 c=0.0473218f //x=1.01 //y=6.025 //x2=0.655 //y2=5.025
cc_124 ( N_noxref_3_M4_noxref_g N_noxref_5_M4_noxref_d ) capacitor \
 c=0.0170604f //x=1.45 //y=6.025 //x2=1.525 //y2=5.025
cc_125 ( N_noxref_3_c_94_n N_noxref_6_c_282_n ) capacitor c=0.00219713f \
 //x=1.11 //y=2.08 //x2=2.96 //y2=2.08
cc_126 ( N_noxref_3_c_104_n N_noxref_7_c_349_n ) capacitor c=0.00431513f \
 //x=1.445 //y=1.25 //x2=2.065 //y2=1.655
cc_127 ( N_noxref_3_c_94_n N_noxref_7_c_374_n ) capacitor c=0.0112169f \
 //x=1.11 //y=2.08 //x2=1.265 //y2=1.655
cc_128 ( N_noxref_3_c_99_n N_noxref_7_c_374_n ) capacitor c=0.00589082f \
 //x=0.915 //y=1.915 //x2=1.265 //y2=1.655
cc_129 ( N_noxref_3_c_97_n N_noxref_7_M0_noxref_d ) capacitor c=0.0013184f \
 //x=0.915 //y=0.905 //x2=0.99 //y2=0.905
cc_130 ( N_noxref_3_c_124_p N_noxref_7_M0_noxref_d ) capacitor c=0.0034598f \
 //x=0.915 //y=1.25 //x2=0.99 //y2=0.905
cc_131 ( N_noxref_3_c_125_p N_noxref_7_M0_noxref_d ) capacitor c=0.00300148f \
 //x=0.915 //y=1.56 //x2=0.99 //y2=0.905
cc_132 ( N_noxref_3_c_99_n N_noxref_7_M0_noxref_d ) capacitor c=0.00274546f \
 //x=0.915 //y=1.915 //x2=0.99 //y2=0.905
cc_133 ( N_noxref_3_c_101_n N_noxref_7_M0_noxref_d ) capacitor c=0.00241102f \
 //x=1.29 //y=0.75 //x2=0.99 //y2=0.905
cc_134 ( N_noxref_3_c_156_p N_noxref_7_M0_noxref_d ) capacitor c=0.0123304f \
 //x=1.29 //y=1.405 //x2=0.99 //y2=0.905
cc_135 ( N_noxref_3_c_102_n N_noxref_7_M0_noxref_d ) capacitor c=0.00219619f \
 //x=1.445 //y=0.905 //x2=0.99 //y2=0.905
cc_136 ( N_noxref_3_c_104_n N_noxref_7_M0_noxref_d ) capacitor c=0.00603828f \
 //x=1.445 //y=1.25 //x2=0.99 //y2=0.905
cc_137 ( N_noxref_4_M5_noxref_g N_noxref_5_c_239_n ) capacitor c=0.0170604f \
 //x=1.89 //y=6.025 //x2=1.585 //y2=5.21
cc_138 ( N_noxref_4_c_190_n N_noxref_5_c_239_n ) capacitor c=2.3112e-19 \
 //x=1.885 //y=4.705 //x2=1.585 //y2=5.21
cc_139 ( N_noxref_4_c_169_n N_noxref_5_c_243_n ) capacitor c=0.00109004f \
 //x=1.85 //y=4.54 //x2=2.465 //y2=6.91
cc_140 ( N_noxref_4_M5_noxref_g N_noxref_5_c_243_n ) capacitor c=0.0148484f \
 //x=1.89 //y=6.025 //x2=2.465 //y2=6.91
cc_141 ( N_noxref_4_M6_noxref_g N_noxref_5_c_243_n ) capacitor c=0.0160244f \
 //x=2.33 //y=6.025 //x2=2.465 //y2=6.91
cc_142 ( N_noxref_4_M6_noxref_g N_noxref_5_M6_noxref_d ) capacitor \
 c=0.0216879f //x=2.33 //y=6.025 //x2=2.405 //y2=5.025
cc_143 ( N_noxref_4_c_169_n N_noxref_6_c_282_n ) capacitor c=0.00562297f \
 //x=1.85 //y=4.54 //x2=2.96 //y2=2.08
cc_144 ( N_noxref_4_c_159_n N_noxref_6_c_282_n ) capacitor c=0.0533475f \
 //x=1.85 //y=2.08 //x2=2.96 //y2=2.08
cc_145 ( N_noxref_4_c_187_n N_noxref_6_c_282_n ) capacitor c=3.80079e-19 \
 //x=1.85 //y=2.08 //x2=2.96 //y2=2.08
cc_146 ( N_noxref_4_c_190_n N_noxref_6_c_282_n ) capacitor c=4.01223e-19 \
 //x=1.885 //y=4.705 //x2=2.96 //y2=2.08
cc_147 ( N_noxref_4_M6_noxref_g N_noxref_6_M7_noxref_g ) capacitor \
 c=0.0343614f //x=2.33 //y=6.025 //x2=3.37 //y2=6.025
cc_148 ( N_noxref_4_c_160_n N_noxref_6_c_284_n ) capacitor c=0.00131574f \
 //x=1.885 //y=0.905 //x2=2.855 //y2=0.905
cc_149 ( N_noxref_4_c_164_n N_noxref_6_c_284_n ) capacitor c=0.00886682f \
 //x=2.415 //y=0.905 //x2=2.855 //y2=0.905
cc_150 ( N_noxref_4_c_179_n N_noxref_6_c_303_n ) capacitor c=0.00150456f \
 //x=1.885 //y=1.255 //x2=2.855 //y2=1.255
cc_151 ( N_noxref_4_c_186_n N_noxref_6_c_303_n ) capacitor c=0.00886682f \
 //x=2.415 //y=1.255 //x2=2.855 //y2=1.255
cc_152 ( N_noxref_4_c_182_n N_noxref_6_c_305_n ) capacitor c=0.00276257f \
 //x=1.885 //y=1.56 //x2=2.855 //y2=1.56
cc_153 ( N_noxref_4_c_163_n N_noxref_6_c_305_n ) capacitor c=0.0177628f \
 //x=2.26 //y=1.405 //x2=2.855 //y2=1.56
cc_154 ( N_noxref_4_c_189_n N_noxref_6_c_307_n ) capacitor c=0.00494016f \
 //x=1.85 //y=1.915 //x2=2.855 //y2=1.915
cc_155 ( N_noxref_4_c_163_n N_noxref_6_c_287_n ) capacitor c=0.00123863f \
 //x=2.26 //y=1.405 //x2=3.23 //y2=1.405
cc_156 ( N_noxref_4_c_164_n N_noxref_6_c_288_n ) capacitor c=0.00132934f \
 //x=2.415 //y=0.905 //x2=3.385 //y2=0.905
cc_157 ( N_noxref_4_c_186_n N_noxref_6_c_310_n ) capacitor c=0.00150456f \
 //x=2.415 //y=1.255 //x2=3.385 //y2=1.255
cc_158 ( N_noxref_4_c_159_n N_noxref_6_c_290_n ) capacitor c=0.00235136f \
 //x=1.85 //y=2.08 //x2=2.855 //y2=2.08
cc_159 ( N_noxref_4_c_187_n N_noxref_6_c_290_n ) capacitor c=0.00922588f \
 //x=1.85 //y=2.08 //x2=2.855 //y2=2.08
cc_160 ( N_noxref_4_c_169_n N_noxref_6_c_313_n ) capacitor c=0.00227279f \
 //x=1.85 //y=4.54 //x2=2.96 //y2=4.705
cc_161 ( N_noxref_4_c_217_p N_noxref_6_c_313_n ) capacitor c=0.0106154f \
 //x=2.255 //y=4.795 //x2=2.96 //y2=4.705
cc_162 ( N_noxref_4_c_190_n N_noxref_6_c_313_n ) capacitor c=0.00510965f \
 //x=1.885 //y=4.705 //x2=2.96 //y2=4.705
cc_163 ( N_noxref_4_c_159_n N_noxref_7_c_349_n ) capacitor c=0.0162392f \
 //x=1.85 //y=2.08 //x2=2.065 //y2=1.655
cc_164 ( N_noxref_4_c_182_n N_noxref_7_c_349_n ) capacitor c=0.00158038f \
 //x=1.885 //y=1.56 //x2=2.065 //y2=1.655
cc_165 ( N_noxref_4_c_187_n N_noxref_7_c_349_n ) capacitor c=0.00633758f \
 //x=1.85 //y=2.08 //x2=2.065 //y2=1.655
cc_166 ( N_noxref_4_c_189_n N_noxref_7_c_349_n ) capacitor c=0.0185539f \
 //x=1.85 //y=1.915 //x2=2.065 //y2=1.655
cc_167 ( N_noxref_4_c_163_n N_noxref_7_c_353_n ) capacitor c=0.00430135f \
 //x=2.26 //y=1.405 //x2=3.035 //y2=1.655
cc_168 ( N_noxref_4_c_159_n N_noxref_7_c_371_n ) capacitor c=0.00265434f \
 //x=1.85 //y=2.08 //x2=3.7 //y2=5.125
cc_169 ( N_noxref_4_c_182_n N_noxref_7_M0_noxref_d ) capacitor c=8.74435e-19 \
 //x=1.885 //y=1.56 //x2=0.99 //y2=0.905
cc_170 ( N_noxref_4_c_160_n N_noxref_7_M1_noxref_d ) capacitor c=0.00132426f \
 //x=1.885 //y=0.905 //x2=1.96 //y2=0.905
cc_171 ( N_noxref_4_c_179_n N_noxref_7_M1_noxref_d ) capacitor c=0.0035101f \
 //x=1.885 //y=1.255 //x2=1.96 //y2=0.905
cc_172 ( N_noxref_4_c_182_n N_noxref_7_M1_noxref_d ) capacitor c=0.00297998f \
 //x=1.885 //y=1.56 //x2=1.96 //y2=0.905
cc_173 ( N_noxref_4_c_162_n N_noxref_7_M1_noxref_d ) capacitor c=0.00241102f \
 //x=2.26 //y=0.75 //x2=1.96 //y2=0.905
cc_174 ( N_noxref_4_c_163_n N_noxref_7_M1_noxref_d ) capacitor c=0.0154425f \
 //x=2.26 //y=1.405 //x2=1.96 //y2=0.905
cc_175 ( N_noxref_4_c_164_n N_noxref_7_M1_noxref_d ) capacitor c=0.00132831f \
 //x=2.415 //y=0.905 //x2=1.96 //y2=0.905
cc_176 ( N_noxref_4_c_186_n N_noxref_7_M1_noxref_d ) capacitor c=0.0035101f \
 //x=2.415 //y=1.255 //x2=1.96 //y2=0.905
cc_177 ( N_noxref_4_M6_noxref_g N_noxref_8_c_432_n ) capacitor c=0.0222438f \
 //x=2.33 //y=6.025 //x2=3.065 //y2=5.21
cc_178 ( N_noxref_4_M5_noxref_g N_noxref_8_c_433_n ) capacitor c=0.0132989f \
 //x=1.89 //y=6.025 //x2=2.195 //y2=5.21
cc_179 ( N_noxref_4_c_217_p N_noxref_8_c_433_n ) capacitor c=0.00417892f \
 //x=2.255 //y=4.795 //x2=2.195 //y2=5.21
cc_180 ( N_noxref_4_M6_noxref_g N_noxref_8_c_435_n ) capacitor c=0.00102459f \
 //x=2.33 //y=6.025 //x2=3.235 //y2=6.91
cc_181 ( N_noxref_4_M6_noxref_g N_noxref_8_M5_noxref_d ) capacitor \
 c=0.0134276f //x=2.33 //y=6.025 //x2=1.965 //y2=5.025
cc_182 ( N_noxref_4_M6_noxref_g N_noxref_8_M7_noxref_s ) capacitor \
 c=0.00207713f //x=2.33 //y=6.025 //x2=3.015 //y2=5.025
cc_183 ( N_noxref_5_c_243_n N_noxref_6_M7_noxref_g ) capacitor c=0.00102459f \
 //x=2.465 //y=6.91 //x2=3.37 //y2=6.025
cc_184 ( N_noxref_5_c_239_n N_noxref_7_c_398_n ) capacitor c=0.00108534f \
 //x=1.585 //y=5.21 //x2=3.7 //y2=5.21
cc_185 ( N_noxref_5_M6_noxref_d N_noxref_7_M7_noxref_d ) capacitor \
 c=0.0049951f //x=2.405 //y=5.025 //x2=3.445 //y2=5.025
cc_186 ( N_noxref_5_c_243_n N_noxref_8_c_432_n ) capacitor c=0.00128698f \
 //x=2.465 //y=6.91 //x2=3.065 //y2=5.21
cc_187 ( N_noxref_5_M6_noxref_d N_noxref_8_c_432_n ) capacitor c=0.0133215f \
 //x=2.405 //y=5.025 //x2=3.065 //y2=5.21
cc_188 ( N_noxref_5_c_239_n N_noxref_8_c_433_n ) capacitor c=0.0351721f \
 //x=1.585 //y=5.21 //x2=2.195 //y2=5.21
cc_189 ( N_noxref_5_c_243_n N_noxref_8_c_435_n ) capacitor c=0.027433f \
 //x=2.465 //y=6.91 //x2=3.235 //y2=6.91
cc_190 ( N_noxref_5_c_243_n N_noxref_8_M5_noxref_d ) capacitor c=0.0118172f \
 //x=2.465 //y=6.91 //x2=1.965 //y2=5.025
cc_191 ( N_noxref_5_M3_noxref_s N_noxref_8_M5_noxref_d ) capacitor \
 c=0.00107541f //x=0.655 //y=5.025 //x2=1.965 //y2=5.025
cc_192 ( N_noxref_5_M4_noxref_d N_noxref_8_M5_noxref_d ) capacitor \
 c=0.0351721f //x=1.525 //y=5.025 //x2=1.965 //y2=5.025
cc_193 ( N_noxref_5_M6_noxref_d N_noxref_8_M5_noxref_d ) capacitor \
 c=0.0458293f //x=2.405 //y=5.025 //x2=1.965 //y2=5.025
cc_194 ( N_noxref_5_M4_noxref_d N_noxref_8_M7_noxref_s ) capacitor \
 c=0.00194853f //x=1.525 //y=5.025 //x2=3.015 //y2=5.025
cc_195 ( N_noxref_5_M6_noxref_d N_noxref_8_M7_noxref_s ) capacitor c=0.027433f \
 //x=2.405 //y=5.025 //x2=3.015 //y2=5.025
cc_196 ( N_noxref_5_M6_noxref_d N_noxref_8_M8_noxref_d ) capacitor \
 c=9.17547e-19 //x=2.405 //y=5.025 //x2=3.885 //y2=5.025
cc_197 ( N_noxref_6_c_282_n N_noxref_7_c_353_n ) capacitor c=0.0182656f \
 //x=2.96 //y=2.08 //x2=3.035 //y2=1.655
cc_198 ( N_noxref_6_c_305_n N_noxref_7_c_353_n ) capacitor c=0.0013609f \
 //x=2.855 //y=1.56 //x2=3.035 //y2=1.655
cc_199 ( N_noxref_6_c_307_n N_noxref_7_c_353_n ) capacitor c=0.0216105f \
 //x=2.855 //y=1.915 //x2=3.035 //y2=1.655
cc_200 ( N_noxref_6_c_290_n N_noxref_7_c_353_n ) capacitor c=0.003666f \
 //x=2.855 //y=2.08 //x2=3.035 //y2=1.655
cc_201 ( N_noxref_6_c_287_n N_noxref_7_c_357_n ) capacitor c=0.00777513f \
 //x=3.23 //y=1.405 //x2=3.615 //y2=1.655
cc_202 ( N_noxref_6_c_282_n N_noxref_7_c_371_n ) capacitor c=0.0935935f \
 //x=2.96 //y=2.08 //x2=3.7 //y2=5.125
cc_203 ( N_noxref_6_M7_noxref_g N_noxref_7_c_371_n ) capacitor c=0.0059988f \
 //x=3.37 //y=6.025 //x2=3.7 //y2=5.125
cc_204 ( N_noxref_6_M8_noxref_g N_noxref_7_c_371_n ) capacitor c=0.0066533f \
 //x=3.81 //y=6.025 //x2=3.7 //y2=5.125
cc_205 ( N_noxref_6_c_307_n N_noxref_7_c_371_n ) capacitor c=0.00278932f \
 //x=2.855 //y=1.915 //x2=3.7 //y2=5.125
cc_206 ( N_noxref_6_c_294_n N_noxref_7_c_371_n ) capacitor c=0.0150293f \
 //x=3.735 //y=4.795 //x2=3.7 //y2=5.125
cc_207 ( N_noxref_6_c_290_n N_noxref_7_c_371_n ) capacitor c=0.00882918f \
 //x=2.855 //y=2.08 //x2=3.7 //y2=5.125
cc_208 ( N_noxref_6_c_313_n N_noxref_7_c_371_n ) capacitor c=0.00513934f \
 //x=2.96 //y=4.705 //x2=3.7 //y2=5.125
cc_209 ( N_noxref_6_c_290_n N_noxref_7_c_412_n ) capacitor c=0.00470847f \
 //x=2.855 //y=2.08 //x2=3.12 //y2=1.655
cc_210 ( N_noxref_6_M7_noxref_g N_noxref_7_c_398_n ) capacitor c=0.0132317f \
 //x=3.37 //y=6.025 //x2=3.7 //y2=5.21
cc_211 ( N_noxref_6_M8_noxref_g N_noxref_7_c_398_n ) capacitor c=0.00775308f \
 //x=3.81 //y=6.025 //x2=3.7 //y2=5.21
cc_212 ( N_noxref_6_c_294_n N_noxref_7_c_398_n ) capacitor c=0.00303922f \
 //x=3.735 //y=4.795 //x2=3.7 //y2=5.21
cc_213 ( N_noxref_6_c_305_n N_noxref_7_M1_noxref_d ) capacitor c=0.00148728f \
 //x=2.855 //y=1.56 //x2=1.96 //y2=0.905
cc_214 ( N_noxref_6_c_284_n N_noxref_7_M2_noxref_d ) capacitor c=0.00226395f \
 //x=2.855 //y=0.905 //x2=2.93 //y2=0.905
cc_215 ( N_noxref_6_c_303_n N_noxref_7_M2_noxref_d ) capacitor c=0.0035101f \
 //x=2.855 //y=1.255 //x2=2.93 //y2=0.905
cc_216 ( N_noxref_6_c_305_n N_noxref_7_M2_noxref_d ) capacitor c=0.00484362f \
 //x=2.855 //y=1.56 //x2=2.93 //y2=0.905
cc_217 ( N_noxref_6_c_307_n N_noxref_7_M2_noxref_d ) capacitor c=3.4952e-19 \
 //x=2.855 //y=1.915 //x2=2.93 //y2=0.905
cc_218 ( N_noxref_6_c_286_n N_noxref_7_M2_noxref_d ) capacitor c=0.00241102f \
 //x=3.23 //y=0.75 //x2=2.93 //y2=0.905
cc_219 ( N_noxref_6_c_287_n N_noxref_7_M2_noxref_d ) capacitor c=0.0156879f \
 //x=3.23 //y=1.405 //x2=2.93 //y2=0.905
cc_220 ( N_noxref_6_c_288_n N_noxref_7_M2_noxref_d ) capacitor c=0.00132831f \
 //x=3.385 //y=0.905 //x2=2.93 //y2=0.905
cc_221 ( N_noxref_6_c_310_n N_noxref_7_M2_noxref_d ) capacitor c=0.0035101f \
 //x=3.385 //y=1.255 //x2=2.93 //y2=0.905
cc_222 ( N_noxref_6_M8_noxref_g N_noxref_7_M7_noxref_d ) capacitor \
 c=0.0136385f //x=3.81 //y=6.025 //x2=3.445 //y2=5.025
cc_223 ( N_noxref_6_c_282_n N_noxref_8_c_432_n ) capacitor c=0.0118924f \
 //x=2.96 //y=2.08 //x2=3.065 //y2=5.21
cc_224 ( N_noxref_6_M7_noxref_g N_noxref_8_c_432_n ) capacitor c=0.0286624f \
 //x=3.37 //y=6.025 //x2=3.065 //y2=5.21
cc_225 ( N_noxref_6_c_313_n N_noxref_8_c_432_n ) capacitor c=0.0161227f \
 //x=2.96 //y=4.705 //x2=3.065 //y2=5.21
cc_226 ( N_noxref_6_M7_noxref_g N_noxref_8_c_434_n ) capacitor c=0.016576f \
 //x=3.37 //y=6.025 //x2=3.945 //y2=6.91
cc_227 ( N_noxref_6_M8_noxref_g N_noxref_8_c_434_n ) capacitor c=0.0166873f \
 //x=3.81 //y=6.025 //x2=3.945 //y2=6.91
cc_228 ( N_noxref_6_M8_noxref_g N_noxref_8_M8_noxref_d ) capacitor \
 c=0.0351101f //x=3.81 //y=6.025 //x2=3.885 //y2=5.025
cc_229 ( N_noxref_7_c_398_n N_noxref_8_c_432_n ) capacitor c=0.0344081f \
 //x=3.7 //y=5.21 //x2=3.065 //y2=5.21
cc_230 ( N_noxref_7_c_398_n N_noxref_8_c_434_n ) capacitor c=0.0012445f \
 //x=3.7 //y=5.21 //x2=3.945 //y2=6.91
cc_231 ( N_noxref_7_M7_noxref_d N_noxref_8_c_434_n ) capacitor c=0.011849f \
 //x=3.445 //y=5.025 //x2=3.945 //y2=6.91
cc_232 ( N_noxref_7_M7_noxref_d N_noxref_8_M5_noxref_d ) capacitor \
 c=0.00101354f //x=3.445 //y=5.025 //x2=1.965 //y2=5.025
cc_233 ( N_noxref_7_M7_noxref_d N_noxref_8_M7_noxref_s ) capacitor \
 c=0.0344081f //x=3.445 //y=5.025 //x2=3.015 //y2=5.025
cc_234 ( N_noxref_7_M7_noxref_d N_noxref_8_M8_noxref_d ) capacitor \
 c=0.0458293f //x=3.445 //y=5.025 //x2=3.885 //y2=5.025
