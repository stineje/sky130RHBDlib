* SPICE3 file created from FA.ext - technology: sky130A

.subckt FA SUM COUT A B CIN VPB VNB
M1000 VPB.t9 CIN a_3461_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VPB.t7 CIN a_3027_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_575_1004.t3 a_807_943.t3 a_836_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_2795_1004.t3 a_836_182.t6 VPB.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_6791_1005.t2 a_5291_182.t3 VPB.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VNB A a_556_74.t0 nshort w=-1.605u l=1.765u
+  ad=10.9968p pd=79.06u as=0p ps=0u
M1006 a_1241_1004.t3 B VPB.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_836_182.t3 a_807_943.t4 a_575_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1241_1004.t0 a_185_182.t4 a_836_182.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPB.t3 a_5767_1004.t6 a_6401_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_2405_182.t2 a_836_182.t7 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPB.t25 B a_807_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_7511_182.t2 a_6858_181.t5 VPB.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VNB a_3027_943.t3 a_3442_74.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPB.t21 B a_5767_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPB.t15 A a_575_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPB.t2 a_836_182.t8 a_4657_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_807_943.t1 B VPB.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_4657_1004.t1 CIN VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VNB CIN a_4552_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1020 SUM a_2405_182.t3 a_3461_1004.t0 pshort w=2u l=0.15u
+  ad=1.16p pd=9.16u as=0p ps=0u
M1021 a_3027_943.t0 CIN VPB.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t28 a_5291_182.t4 a_6791_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPB.t19 A a_185_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_2795_1004.t1 a_3027_943.t4 SUM pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_4657_1004.t2 a_836_182.t9 VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_6791_1005.t0 a_6401_182.t3 a_6858_181.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPB.t24 B a_1241_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_5291_182.t2 a_4657_1004.t5 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_3461_1004.t2 CIN VPB.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPB.t26 a_6858_181.t6 a_7511_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 VNB B a_5662_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1032 SUM a_2405_182.t4 a_3442_74.t1 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.14u as=0p ps=0u
M1033 a_575_1004.t0 A VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_836_182.t1 a_185_182.t5 a_1241_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPB.t13 a_836_182.t12 a_2795_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_5767_1004.t3 B VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPB.t17 A a_5767_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VNB a_836_182.t11 a_2776_74.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPB.t30 a_836_182.t14 a_2405_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 VPB.t5 a_4657_1004.t7 a_5291_182.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_5767_1004.t1 A VPB.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VNB a_807_943.t5 a_1222_74.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_185_182.t1 A VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 SUM CIN a_2776_74.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1045 SUM a_3027_943.t5 a_2795_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPB.t6 CIN a_4657_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_6401_182.t1 a_5767_1004.t7 VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_6858_181.t1 a_6401_182.t5 a_6791_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_3461_1004.t1 a_2405_182.t5 SUM pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 A B 0.77fF
C1 A CIN 0.44fF
C2 VPB A 0.42fF
C3 B CIN 1.74fF
C4 VPB B 0.93fF
C5 VPB CIN 0.58fF
C6 SUM A 0.17fF
C7 SUM B 0.24fF
C8 SUM CIN 0.81fF
C9 VPB SUM 0.53fF
R0 a_3461_1004.n0 a_3461_1004.t1 101.66
R1 a_3461_1004.n0 a_3461_1004.t3 101.66
R2 a_3461_1004.t0 a_3461_1004.n0 14.294
R3 a_3461_1004.n0 a_3461_1004.t2 14.282
R4 VPB VPB.n765 126.832
R5 VPB.n60 VPB.n58 94.117
R6 VPB.n740 VPB.n738 94.117
R7 VPB.n681 VPB.n679 94.117
R8 VPB.n634 VPB.n632 94.117
R9 VPB.n587 VPB.n585 94.117
R10 VPB.n528 VPB.n526 94.117
R11 VPB.n470 VPB.n468 94.117
R12 VPB.n137 VPB.n135 94.117
R13 VPB.n440 VPB.n438 94.117
R14 VPB.n393 VPB.n391 94.117
R15 VPB.n330 VPB.n328 94.117
R16 VPB.n283 VPB.n281 94.117
R17 VPB.n224 VPB.n222 94.117
R18 VPB.n185 VPB.n179 76.136
R19 VPB.n185 VPB.n184 76
R20 VPB.n189 VPB.n188 76
R21 VPB.n195 VPB.n194 76
R22 VPB.n199 VPB.n198 76
R23 VPB.n226 VPB.n225 76
R24 VPB.n230 VPB.n229 76
R25 VPB.n234 VPB.n233 76
R26 VPB.n238 VPB.n237 76
R27 VPB.n243 VPB.n242 76
R28 VPB.n250 VPB.n249 76
R29 VPB.n254 VPB.n253 76
R30 VPB.n258 VPB.n257 76
R31 VPB.n285 VPB.n284 76
R32 VPB.n291 VPB.n290 76
R33 VPB.n295 VPB.n294 76
R34 VPB.n301 VPB.n300 76
R35 VPB.n305 VPB.n304 76
R36 VPB.n332 VPB.n331 76
R37 VPB.n337 VPB.n336 76
R38 VPB.n342 VPB.n341 76
R39 VPB.n349 VPB.n348 76
R40 VPB.n354 VPB.n353 76
R41 VPB.n359 VPB.n358 76
R42 VPB.n364 VPB.n363 76
R43 VPB.n368 VPB.n367 76
R44 VPB.n395 VPB.n394 76
R45 VPB.n401 VPB.n400 76
R46 VPB.n405 VPB.n404 76
R47 VPB.n411 VPB.n410 76
R48 VPB.n415 VPB.n414 76
R49 VPB.n442 VPB.n441 76
R50 VPB.n447 VPB.n446 76
R51 VPB.n452 VPB.n451 76
R52 VPB.n457 VPB.n456 76
R53 VPB.n471 VPB.n467 76
R54 VPB.n475 VPB.n474 76
R55 VPB.n479 VPB.n478 76
R56 VPB.n483 VPB.n482 76
R57 VPB.n488 VPB.n487 76
R58 VPB.n495 VPB.n494 76
R59 VPB.n499 VPB.n498 76
R60 VPB.n503 VPB.n502 76
R61 VPB.n530 VPB.n529 76
R62 VPB.n534 VPB.n533 76
R63 VPB.n538 VPB.n537 76
R64 VPB.n542 VPB.n541 76
R65 VPB.n547 VPB.n546 76
R66 VPB.n554 VPB.n553 76
R67 VPB.n558 VPB.n557 76
R68 VPB.n562 VPB.n561 76
R69 VPB.n589 VPB.n588 76
R70 VPB.n595 VPB.n594 76
R71 VPB.n599 VPB.n598 76
R72 VPB.n605 VPB.n604 76
R73 VPB.n609 VPB.n608 76
R74 VPB.n636 VPB.n635 76
R75 VPB.n642 VPB.n641 76
R76 VPB.n646 VPB.n645 76
R77 VPB.n652 VPB.n651 76
R78 VPB.n656 VPB.n655 76
R79 VPB.n683 VPB.n682 76
R80 VPB.n687 VPB.n686 76
R81 VPB.n691 VPB.n690 76
R82 VPB.n695 VPB.n694 76
R83 VPB.n700 VPB.n699 76
R84 VPB.n707 VPB.n706 76
R85 VPB.n711 VPB.n710 76
R86 VPB.n715 VPB.n714 76
R87 VPB.n742 VPB.n741 76
R88 VPB.n746 VPB.n745 76
R89 VPB.n758 VPB.n757 76
R90 VPB.n192 VPB.n191 68.979
R91 VPB.n298 VPB.n297 68.979
R92 VPB.n408 VPB.n407 68.979
R93 VPB.n141 VPB.n140 68.979
R94 VPB.n602 VPB.n601 68.979
R95 VPB.n639 VPB.n638 68.979
R96 VPB.n71 VPB.n70 68.979
R97 VPB.n46 VPB.n35 65.944
R98 VPB.n702 VPB.n701 65.944
R99 VPB.n549 VPB.n548 65.944
R100 VPB.n490 VPB.n489 65.944
R101 VPB.n182 VPB.n181 64.528
R102 VPB.n288 VPB.n287 64.528
R103 VPB.n398 VPB.n397 64.528
R104 VPB.n148 VPB.n147 64.528
R105 VPB.n592 VPB.n591 64.528
R106 VPB.n649 VPB.n648 64.528
R107 VPB.n64 VPB.n63 64.528
R108 VPB.n20 VPB.n19 61.764
R109 VPB.n722 VPB.n721 61.764
R110 VPB.n663 VPB.n662 61.764
R111 VPB.n616 VPB.n615 61.764
R112 VPB.n569 VPB.n568 61.764
R113 VPB.n510 VPB.n509 61.764
R114 VPB.n81 VPB.n80 61.764
R115 VPB.n102 VPB.n101 61.764
R116 VPB.n422 VPB.n421 61.764
R117 VPB.n375 VPB.n374 61.764
R118 VPB.n312 VPB.n311 61.764
R119 VPB.n265 VPB.n264 61.764
R120 VPB.n206 VPB.n205 61.764
R121 VPB.n74 VPB.t18 55.106
R122 VPB.n62 VPB.t19 55.106
R123 VPB.n647 VPB.t22 55.106
R124 VPB.n637 VPB.t25 55.106
R125 VPB.n600 VPB.t1 55.106
R126 VPB.n590 VPB.t30 55.106
R127 VPB.n151 VPB.t10 55.106
R128 VPB.n139 VPB.t7 55.106
R129 VPB.n127 VPB.t11 55.106
R130 VPB.n406 VPB.t12 55.106
R131 VPB.n396 VPB.t5 55.106
R132 VPB.n360 VPB.t20 55.106
R133 VPB.n296 VPB.t4 55.106
R134 VPB.n286 VPB.t3 55.106
R135 VPB.n190 VPB.t27 55.106
R136 VPB.n180 VPB.t26 55.106
R137 VPB.n443 VPB.t2 55.106
R138 VPB.n333 VPB.t17 55.106
R139 VPB.n339 VPB.n338 48.952
R140 VPB.n449 VPB.n448 48.952
R141 VPB.n247 VPB.n246 44.502
R142 VPB.n356 VPB.n355 44.502
R143 VPB.n124 VPB.n123 44.502
R144 VPB.n492 VPB.n491 44.502
R145 VPB.n551 VPB.n550 44.502
R146 VPB.n704 VPB.n703 44.502
R147 VPB.n48 VPB.n47 44.502
R148 VPB.n245 VPB.n244 41.183
R149 VPB.n118 VPB.n117 40.824
R150 VPB.n344 VPB.n343 40.824
R151 VPB.n762 VPB.n758 20.452
R152 VPB.n179 VPB.n176 20.452
R153 VPB.n346 VPB.n345 17.801
R154 VPB.n454 VPB.n453 17.801
R155 VPB.n35 VPB.t14 14.282
R156 VPB.n35 VPB.t15 14.282
R157 VPB.n701 VPB.t23 14.282
R158 VPB.n701 VPB.t24 14.282
R159 VPB.n548 VPB.t31 14.282
R160 VPB.n548 VPB.t13 14.282
R161 VPB.n489 VPB.t8 14.282
R162 VPB.n489 VPB.t9 14.282
R163 VPB.n117 VPB.t0 14.282
R164 VPB.n117 VPB.t6 14.282
R165 VPB.n343 VPB.t16 14.282
R166 VPB.n343 VPB.t21 14.282
R167 VPB.n244 VPB.t29 14.282
R168 VPB.n244 VPB.t28 14.282
R169 VPB.n179 VPB.n178 13.653
R170 VPB.n178 VPB.n177 13.653
R171 VPB.n184 VPB.n183 13.653
R172 VPB.n183 VPB.n182 13.653
R173 VPB.n188 VPB.n187 13.653
R174 VPB.n187 VPB.n186 13.653
R175 VPB.n194 VPB.n193 13.653
R176 VPB.n193 VPB.n192 13.653
R177 VPB.n198 VPB.n197 13.653
R178 VPB.n197 VPB.n196 13.653
R179 VPB.n225 VPB.n224 13.653
R180 VPB.n224 VPB.n223 13.653
R181 VPB.n229 VPB.n228 13.653
R182 VPB.n228 VPB.n227 13.653
R183 VPB.n233 VPB.n232 13.653
R184 VPB.n232 VPB.n231 13.653
R185 VPB.n237 VPB.n236 13.653
R186 VPB.n236 VPB.n235 13.653
R187 VPB.n242 VPB.n241 13.653
R188 VPB.n241 VPB.n240 13.653
R189 VPB.n249 VPB.n248 13.653
R190 VPB.n248 VPB.n247 13.653
R191 VPB.n253 VPB.n252 13.653
R192 VPB.n252 VPB.n251 13.653
R193 VPB.n257 VPB.n256 13.653
R194 VPB.n256 VPB.n255 13.653
R195 VPB.n284 VPB.n283 13.653
R196 VPB.n283 VPB.n282 13.653
R197 VPB.n290 VPB.n289 13.653
R198 VPB.n289 VPB.n288 13.653
R199 VPB.n294 VPB.n293 13.653
R200 VPB.n293 VPB.n292 13.653
R201 VPB.n300 VPB.n299 13.653
R202 VPB.n299 VPB.n298 13.653
R203 VPB.n304 VPB.n303 13.653
R204 VPB.n303 VPB.n302 13.653
R205 VPB.n331 VPB.n330 13.653
R206 VPB.n330 VPB.n329 13.653
R207 VPB.n336 VPB.n335 13.653
R208 VPB.n335 VPB.n334 13.653
R209 VPB.n341 VPB.n340 13.653
R210 VPB.n340 VPB.n339 13.653
R211 VPB.n348 VPB.n347 13.653
R212 VPB.n347 VPB.n346 13.653
R213 VPB.n353 VPB.n352 13.653
R214 VPB.n352 VPB.n351 13.653
R215 VPB.n358 VPB.n357 13.653
R216 VPB.n357 VPB.n356 13.653
R217 VPB.n363 VPB.n362 13.653
R218 VPB.n362 VPB.n361 13.653
R219 VPB.n367 VPB.n366 13.653
R220 VPB.n366 VPB.n365 13.653
R221 VPB.n394 VPB.n393 13.653
R222 VPB.n393 VPB.n392 13.653
R223 VPB.n400 VPB.n399 13.653
R224 VPB.n399 VPB.n398 13.653
R225 VPB.n404 VPB.n403 13.653
R226 VPB.n403 VPB.n402 13.653
R227 VPB.n410 VPB.n409 13.653
R228 VPB.n409 VPB.n408 13.653
R229 VPB.n414 VPB.n413 13.653
R230 VPB.n413 VPB.n412 13.653
R231 VPB.n441 VPB.n440 13.653
R232 VPB.n440 VPB.n439 13.653
R233 VPB.n446 VPB.n445 13.653
R234 VPB.n445 VPB.n444 13.653
R235 VPB.n451 VPB.n450 13.653
R236 VPB.n450 VPB.n449 13.653
R237 VPB.n456 VPB.n455 13.653
R238 VPB.n455 VPB.n454 13.653
R239 VPB.n122 VPB.n121 13.653
R240 VPB.n121 VPB.n120 13.653
R241 VPB.n126 VPB.n125 13.653
R242 VPB.n125 VPB.n124 13.653
R243 VPB.n130 VPB.n129 13.653
R244 VPB.n129 VPB.n128 13.653
R245 VPB.n133 VPB.n132 13.653
R246 VPB.n132 VPB.n131 13.653
R247 VPB.n138 VPB.n137 13.653
R248 VPB.n137 VPB.n136 13.653
R249 VPB.n143 VPB.n142 13.653
R250 VPB.n142 VPB.n141 13.653
R251 VPB.n146 VPB.n145 13.653
R252 VPB.n145 VPB.n144 13.653
R253 VPB.n150 VPB.n149 13.653
R254 VPB.n149 VPB.n148 13.653
R255 VPB.n154 VPB.n153 13.653
R256 VPB.n153 VPB.n152 13.653
R257 VPB.n471 VPB.n470 13.653
R258 VPB.n470 VPB.n469 13.653
R259 VPB.n474 VPB.n473 13.653
R260 VPB.n473 VPB.n472 13.653
R261 VPB.n478 VPB.n477 13.653
R262 VPB.n477 VPB.n476 13.653
R263 VPB.n482 VPB.n481 13.653
R264 VPB.n481 VPB.n480 13.653
R265 VPB.n487 VPB.n486 13.653
R266 VPB.n486 VPB.n485 13.653
R267 VPB.n494 VPB.n493 13.653
R268 VPB.n493 VPB.n492 13.653
R269 VPB.n498 VPB.n497 13.653
R270 VPB.n497 VPB.n496 13.653
R271 VPB.n502 VPB.n501 13.653
R272 VPB.n501 VPB.n500 13.653
R273 VPB.n529 VPB.n528 13.653
R274 VPB.n528 VPB.n527 13.653
R275 VPB.n533 VPB.n532 13.653
R276 VPB.n532 VPB.n531 13.653
R277 VPB.n537 VPB.n536 13.653
R278 VPB.n536 VPB.n535 13.653
R279 VPB.n541 VPB.n540 13.653
R280 VPB.n540 VPB.n539 13.653
R281 VPB.n546 VPB.n545 13.653
R282 VPB.n545 VPB.n544 13.653
R283 VPB.n553 VPB.n552 13.653
R284 VPB.n552 VPB.n551 13.653
R285 VPB.n557 VPB.n556 13.653
R286 VPB.n556 VPB.n555 13.653
R287 VPB.n561 VPB.n560 13.653
R288 VPB.n560 VPB.n559 13.653
R289 VPB.n588 VPB.n587 13.653
R290 VPB.n587 VPB.n586 13.653
R291 VPB.n594 VPB.n593 13.653
R292 VPB.n593 VPB.n592 13.653
R293 VPB.n598 VPB.n597 13.653
R294 VPB.n597 VPB.n596 13.653
R295 VPB.n604 VPB.n603 13.653
R296 VPB.n603 VPB.n602 13.653
R297 VPB.n608 VPB.n607 13.653
R298 VPB.n607 VPB.n606 13.653
R299 VPB.n635 VPB.n634 13.653
R300 VPB.n634 VPB.n633 13.653
R301 VPB.n641 VPB.n640 13.653
R302 VPB.n640 VPB.n639 13.653
R303 VPB.n645 VPB.n644 13.653
R304 VPB.n644 VPB.n643 13.653
R305 VPB.n651 VPB.n650 13.653
R306 VPB.n650 VPB.n649 13.653
R307 VPB.n655 VPB.n654 13.653
R308 VPB.n654 VPB.n653 13.653
R309 VPB.n682 VPB.n681 13.653
R310 VPB.n681 VPB.n680 13.653
R311 VPB.n686 VPB.n685 13.653
R312 VPB.n685 VPB.n684 13.653
R313 VPB.n690 VPB.n689 13.653
R314 VPB.n689 VPB.n688 13.653
R315 VPB.n694 VPB.n693 13.653
R316 VPB.n693 VPB.n692 13.653
R317 VPB.n699 VPB.n698 13.653
R318 VPB.n698 VPB.n697 13.653
R319 VPB.n706 VPB.n705 13.653
R320 VPB.n705 VPB.n704 13.653
R321 VPB.n710 VPB.n709 13.653
R322 VPB.n709 VPB.n708 13.653
R323 VPB.n714 VPB.n713 13.653
R324 VPB.n713 VPB.n712 13.653
R325 VPB.n741 VPB.n740 13.653
R326 VPB.n740 VPB.n739 13.653
R327 VPB.n745 VPB.n744 13.653
R328 VPB.n744 VPB.n743 13.653
R329 VPB.n38 VPB.n37 13.653
R330 VPB.n37 VPB.n36 13.653
R331 VPB.n41 VPB.n40 13.653
R332 VPB.n40 VPB.n39 13.653
R333 VPB.n45 VPB.n44 13.653
R334 VPB.n44 VPB.n43 13.653
R335 VPB.n50 VPB.n49 13.653
R336 VPB.n49 VPB.n48 13.653
R337 VPB.n53 VPB.n52 13.653
R338 VPB.n52 VPB.n51 13.653
R339 VPB.n56 VPB.n55 13.653
R340 VPB.n55 VPB.n54 13.653
R341 VPB.n61 VPB.n60 13.653
R342 VPB.n60 VPB.n59 13.653
R343 VPB.n66 VPB.n65 13.653
R344 VPB.n65 VPB.n64 13.653
R345 VPB.n69 VPB.n68 13.653
R346 VPB.n68 VPB.n67 13.653
R347 VPB.n73 VPB.n72 13.653
R348 VPB.n72 VPB.n71 13.653
R349 VPB.n758 VPB.n0 13.653
R350 VPB VPB.n0 13.653
R351 VPB.n240 VPB.n239 13.35
R352 VPB.n351 VPB.n350 13.35
R353 VPB.n120 VPB.n119 13.35
R354 VPB.n485 VPB.n484 13.35
R355 VPB.n544 VPB.n543 13.35
R356 VPB.n697 VPB.n696 13.35
R357 VPB.n43 VPB.n42 13.35
R358 VPB.n762 VPB.n761 13.276
R359 VPB.n761 VPB.n759 13.276
R360 VPB.n34 VPB.n16 13.276
R361 VPB.n16 VPB.n14 13.276
R362 VPB.n736 VPB.n718 13.276
R363 VPB.n718 VPB.n716 13.276
R364 VPB.n677 VPB.n659 13.276
R365 VPB.n659 VPB.n657 13.276
R366 VPB.n630 VPB.n612 13.276
R367 VPB.n612 VPB.n610 13.276
R368 VPB.n583 VPB.n565 13.276
R369 VPB.n565 VPB.n563 13.276
R370 VPB.n524 VPB.n506 13.276
R371 VPB.n506 VPB.n504 13.276
R372 VPB.n95 VPB.n77 13.276
R373 VPB.n77 VPB.n75 13.276
R374 VPB.n116 VPB.n98 13.276
R375 VPB.n98 VPB.n96 13.276
R376 VPB.n436 VPB.n418 13.276
R377 VPB.n418 VPB.n416 13.276
R378 VPB.n389 VPB.n371 13.276
R379 VPB.n371 VPB.n369 13.276
R380 VPB.n326 VPB.n308 13.276
R381 VPB.n308 VPB.n306 13.276
R382 VPB.n279 VPB.n261 13.276
R383 VPB.n261 VPB.n259 13.276
R384 VPB.n220 VPB.n202 13.276
R385 VPB.n202 VPB.n200 13.276
R386 VPB.n225 VPB.n221 13.276
R387 VPB.n284 VPB.n280 13.276
R388 VPB.n331 VPB.n327 13.276
R389 VPB.n394 VPB.n390 13.276
R390 VPB.n441 VPB.n437 13.276
R391 VPB.n126 VPB.n122 13.276
R392 VPB.n133 VPB.n130 13.276
R393 VPB.n134 VPB.n133 13.276
R394 VPB.n138 VPB.n134 13.276
R395 VPB.n146 VPB.n143 13.276
R396 VPB.n150 VPB.n146 13.276
R397 VPB.n155 VPB.n154 13.276
R398 VPB.n471 VPB.n155 13.276
R399 VPB.n474 VPB.n471 13.276
R400 VPB.n529 VPB.n525 13.276
R401 VPB.n588 VPB.n584 13.276
R402 VPB.n635 VPB.n631 13.276
R403 VPB.n682 VPB.n678 13.276
R404 VPB.n741 VPB.n737 13.276
R405 VPB.n41 VPB.n38 13.276
R406 VPB.n45 VPB.n41 13.276
R407 VPB.n53 VPB.n50 13.276
R408 VPB.n56 VPB.n53 13.276
R409 VPB.n57 VPB.n56 13.276
R410 VPB.n61 VPB.n57 13.276
R411 VPB.n69 VPB.n66 13.276
R412 VPB.n73 VPB.n69 13.276
R413 VPB.n176 VPB.n158 13.276
R414 VPB.n158 VPB.n156 13.276
R415 VPB.n163 VPB.n161 12.796
R416 VPB.n163 VPB.n162 12.564
R417 VPB.n172 VPB.n171 12.198
R418 VPB.n170 VPB.n169 12.198
R419 VPB.n166 VPB.n165 12.198
R420 VPB.n127 VPB.n126 11.482
R421 VPB.n139 VPB.n138 10.944
R422 VPB.n758 VPB.n74 10.944
R423 VPB.n154 VPB.n151 10.585
R424 VPB.n62 VPB.n61 10.585
R425 VPB.n46 VPB.n45 8.97
R426 VPB.n176 VPB.n175 7.5
R427 VPB.n161 VPB.n160 7.5
R428 VPB.n165 VPB.n164 7.5
R429 VPB.n169 VPB.n168 7.5
R430 VPB.n158 VPB.n157 7.5
R431 VPB.n173 VPB.n159 7.5
R432 VPB.n202 VPB.n201 7.5
R433 VPB.n215 VPB.n214 7.5
R434 VPB.n209 VPB.n208 7.5
R435 VPB.n211 VPB.n210 7.5
R436 VPB.n204 VPB.n203 7.5
R437 VPB.n220 VPB.n219 7.5
R438 VPB.n261 VPB.n260 7.5
R439 VPB.n274 VPB.n273 7.5
R440 VPB.n268 VPB.n267 7.5
R441 VPB.n270 VPB.n269 7.5
R442 VPB.n263 VPB.n262 7.5
R443 VPB.n279 VPB.n278 7.5
R444 VPB.n308 VPB.n307 7.5
R445 VPB.n321 VPB.n320 7.5
R446 VPB.n315 VPB.n314 7.5
R447 VPB.n317 VPB.n316 7.5
R448 VPB.n310 VPB.n309 7.5
R449 VPB.n326 VPB.n325 7.5
R450 VPB.n371 VPB.n370 7.5
R451 VPB.n384 VPB.n383 7.5
R452 VPB.n378 VPB.n377 7.5
R453 VPB.n380 VPB.n379 7.5
R454 VPB.n373 VPB.n372 7.5
R455 VPB.n389 VPB.n388 7.5
R456 VPB.n418 VPB.n417 7.5
R457 VPB.n431 VPB.n430 7.5
R458 VPB.n425 VPB.n424 7.5
R459 VPB.n427 VPB.n426 7.5
R460 VPB.n420 VPB.n419 7.5
R461 VPB.n436 VPB.n435 7.5
R462 VPB.n98 VPB.n97 7.5
R463 VPB.n111 VPB.n110 7.5
R464 VPB.n105 VPB.n104 7.5
R465 VPB.n107 VPB.n106 7.5
R466 VPB.n100 VPB.n99 7.5
R467 VPB.n116 VPB.n115 7.5
R468 VPB.n77 VPB.n76 7.5
R469 VPB.n90 VPB.n89 7.5
R470 VPB.n84 VPB.n83 7.5
R471 VPB.n86 VPB.n85 7.5
R472 VPB.n79 VPB.n78 7.5
R473 VPB.n95 VPB.n94 7.5
R474 VPB.n506 VPB.n505 7.5
R475 VPB.n519 VPB.n518 7.5
R476 VPB.n513 VPB.n512 7.5
R477 VPB.n515 VPB.n514 7.5
R478 VPB.n508 VPB.n507 7.5
R479 VPB.n524 VPB.n523 7.5
R480 VPB.n565 VPB.n564 7.5
R481 VPB.n578 VPB.n577 7.5
R482 VPB.n572 VPB.n571 7.5
R483 VPB.n574 VPB.n573 7.5
R484 VPB.n567 VPB.n566 7.5
R485 VPB.n583 VPB.n582 7.5
R486 VPB.n612 VPB.n611 7.5
R487 VPB.n625 VPB.n624 7.5
R488 VPB.n619 VPB.n618 7.5
R489 VPB.n621 VPB.n620 7.5
R490 VPB.n614 VPB.n613 7.5
R491 VPB.n630 VPB.n629 7.5
R492 VPB.n659 VPB.n658 7.5
R493 VPB.n672 VPB.n671 7.5
R494 VPB.n666 VPB.n665 7.5
R495 VPB.n668 VPB.n667 7.5
R496 VPB.n661 VPB.n660 7.5
R497 VPB.n677 VPB.n676 7.5
R498 VPB.n718 VPB.n717 7.5
R499 VPB.n731 VPB.n730 7.5
R500 VPB.n725 VPB.n724 7.5
R501 VPB.n727 VPB.n726 7.5
R502 VPB.n720 VPB.n719 7.5
R503 VPB.n736 VPB.n735 7.5
R504 VPB.n16 VPB.n15 7.5
R505 VPB.n29 VPB.n28 7.5
R506 VPB.n23 VPB.n22 7.5
R507 VPB.n25 VPB.n24 7.5
R508 VPB.n18 VPB.n17 7.5
R509 VPB.n34 VPB.n33 7.5
R510 VPB.n761 VPB.n760 7.5
R511 VPB.n12 VPB.n11 7.5
R512 VPB.n6 VPB.n5 7.5
R513 VPB.n8 VPB.n7 7.5
R514 VPB.n2 VPB.n1 7.5
R515 VPB.n763 VPB.n762 7.5
R516 VPB.n57 VPB.n34 7.176
R517 VPB.n737 VPB.n736 7.176
R518 VPB.n678 VPB.n677 7.176
R519 VPB.n631 VPB.n630 7.176
R520 VPB.n584 VPB.n583 7.176
R521 VPB.n525 VPB.n524 7.176
R522 VPB.n155 VPB.n95 7.176
R523 VPB.n134 VPB.n116 7.176
R524 VPB.n437 VPB.n436 7.176
R525 VPB.n390 VPB.n389 7.176
R526 VPB.n327 VPB.n326 7.176
R527 VPB.n280 VPB.n279 7.176
R528 VPB.n221 VPB.n220 7.176
R529 VPB.n122 VPB.n118 6.817
R530 VPB.n216 VPB.n213 6.729
R531 VPB.n212 VPB.n209 6.729
R532 VPB.n207 VPB.n204 6.729
R533 VPB.n275 VPB.n272 6.729
R534 VPB.n271 VPB.n268 6.729
R535 VPB.n266 VPB.n263 6.729
R536 VPB.n322 VPB.n319 6.729
R537 VPB.n318 VPB.n315 6.729
R538 VPB.n313 VPB.n310 6.729
R539 VPB.n385 VPB.n382 6.729
R540 VPB.n381 VPB.n378 6.729
R541 VPB.n376 VPB.n373 6.729
R542 VPB.n432 VPB.n429 6.729
R543 VPB.n428 VPB.n425 6.729
R544 VPB.n423 VPB.n420 6.729
R545 VPB.n112 VPB.n109 6.729
R546 VPB.n108 VPB.n105 6.729
R547 VPB.n103 VPB.n100 6.729
R548 VPB.n91 VPB.n88 6.729
R549 VPB.n87 VPB.n84 6.729
R550 VPB.n82 VPB.n79 6.729
R551 VPB.n520 VPB.n517 6.729
R552 VPB.n516 VPB.n513 6.729
R553 VPB.n511 VPB.n508 6.729
R554 VPB.n579 VPB.n576 6.729
R555 VPB.n575 VPB.n572 6.729
R556 VPB.n570 VPB.n567 6.729
R557 VPB.n626 VPB.n623 6.729
R558 VPB.n622 VPB.n619 6.729
R559 VPB.n617 VPB.n614 6.729
R560 VPB.n673 VPB.n670 6.729
R561 VPB.n669 VPB.n666 6.729
R562 VPB.n664 VPB.n661 6.729
R563 VPB.n732 VPB.n729 6.729
R564 VPB.n728 VPB.n725 6.729
R565 VPB.n723 VPB.n720 6.729
R566 VPB.n30 VPB.n27 6.729
R567 VPB.n26 VPB.n23 6.729
R568 VPB.n21 VPB.n18 6.729
R569 VPB.n13 VPB.n10 6.729
R570 VPB.n9 VPB.n6 6.729
R571 VPB.n4 VPB.n2 6.729
R572 VPB.n207 VPB.n206 6.728
R573 VPB.n212 VPB.n211 6.728
R574 VPB.n216 VPB.n215 6.728
R575 VPB.n219 VPB.n218 6.728
R576 VPB.n266 VPB.n265 6.728
R577 VPB.n271 VPB.n270 6.728
R578 VPB.n275 VPB.n274 6.728
R579 VPB.n278 VPB.n277 6.728
R580 VPB.n313 VPB.n312 6.728
R581 VPB.n318 VPB.n317 6.728
R582 VPB.n322 VPB.n321 6.728
R583 VPB.n325 VPB.n324 6.728
R584 VPB.n376 VPB.n375 6.728
R585 VPB.n381 VPB.n380 6.728
R586 VPB.n385 VPB.n384 6.728
R587 VPB.n388 VPB.n387 6.728
R588 VPB.n423 VPB.n422 6.728
R589 VPB.n428 VPB.n427 6.728
R590 VPB.n432 VPB.n431 6.728
R591 VPB.n435 VPB.n434 6.728
R592 VPB.n103 VPB.n102 6.728
R593 VPB.n108 VPB.n107 6.728
R594 VPB.n112 VPB.n111 6.728
R595 VPB.n115 VPB.n114 6.728
R596 VPB.n82 VPB.n81 6.728
R597 VPB.n87 VPB.n86 6.728
R598 VPB.n91 VPB.n90 6.728
R599 VPB.n94 VPB.n93 6.728
R600 VPB.n511 VPB.n510 6.728
R601 VPB.n516 VPB.n515 6.728
R602 VPB.n520 VPB.n519 6.728
R603 VPB.n523 VPB.n522 6.728
R604 VPB.n570 VPB.n569 6.728
R605 VPB.n575 VPB.n574 6.728
R606 VPB.n579 VPB.n578 6.728
R607 VPB.n582 VPB.n581 6.728
R608 VPB.n617 VPB.n616 6.728
R609 VPB.n622 VPB.n621 6.728
R610 VPB.n626 VPB.n625 6.728
R611 VPB.n629 VPB.n628 6.728
R612 VPB.n664 VPB.n663 6.728
R613 VPB.n669 VPB.n668 6.728
R614 VPB.n673 VPB.n672 6.728
R615 VPB.n676 VPB.n675 6.728
R616 VPB.n723 VPB.n722 6.728
R617 VPB.n728 VPB.n727 6.728
R618 VPB.n732 VPB.n731 6.728
R619 VPB.n735 VPB.n734 6.728
R620 VPB.n21 VPB.n20 6.728
R621 VPB.n26 VPB.n25 6.728
R622 VPB.n30 VPB.n29 6.728
R623 VPB.n33 VPB.n32 6.728
R624 VPB.n4 VPB.n3 6.728
R625 VPB.n9 VPB.n8 6.728
R626 VPB.n13 VPB.n12 6.728
R627 VPB.n764 VPB.n763 6.728
R628 VPB.n348 VPB.n344 6.458
R629 VPB.n175 VPB.n174 6.398
R630 VPB.n249 VPB.n245 4.305
R631 VPB.n494 VPB.n490 4.305
R632 VPB.n553 VPB.n549 4.305
R633 VPB.n706 VPB.n702 4.305
R634 VPB.n50 VPB.n46 4.305
R635 VPB.n184 VPB.n180 2.691
R636 VPB.n290 VPB.n286 2.691
R637 VPB.n400 VPB.n396 2.691
R638 VPB.n151 VPB.n150 2.691
R639 VPB.n594 VPB.n590 2.691
R640 VPB.n651 VPB.n647 2.691
R641 VPB.n66 VPB.n62 2.691
R642 VPB.n194 VPB.n190 2.332
R643 VPB.n300 VPB.n296 2.332
R644 VPB.n410 VPB.n406 2.332
R645 VPB.n143 VPB.n139 2.332
R646 VPB.n604 VPB.n600 2.332
R647 VPB.n641 VPB.n637 2.332
R648 VPB.n74 VPB.n73 2.332
R649 VPB.n363 VPB.n360 1.794
R650 VPB.n130 VPB.n127 1.794
R651 VPB.n336 VPB.n333 1.435
R652 VPB.n446 VPB.n443 1.435
R653 VPB.n173 VPB.n166 1.402
R654 VPB.n173 VPB.n167 1.402
R655 VPB.n173 VPB.n170 1.402
R656 VPB.n173 VPB.n172 1.402
R657 VPB.n174 VPB.n173 0.735
R658 VPB.n173 VPB.n163 0.735
R659 VPB.n217 VPB.n216 0.387
R660 VPB.n217 VPB.n212 0.387
R661 VPB.n217 VPB.n207 0.387
R662 VPB.n218 VPB.n217 0.387
R663 VPB.n276 VPB.n275 0.387
R664 VPB.n276 VPB.n271 0.387
R665 VPB.n276 VPB.n266 0.387
R666 VPB.n277 VPB.n276 0.387
R667 VPB.n323 VPB.n322 0.387
R668 VPB.n323 VPB.n318 0.387
R669 VPB.n323 VPB.n313 0.387
R670 VPB.n324 VPB.n323 0.387
R671 VPB.n386 VPB.n385 0.387
R672 VPB.n386 VPB.n381 0.387
R673 VPB.n386 VPB.n376 0.387
R674 VPB.n387 VPB.n386 0.387
R675 VPB.n433 VPB.n432 0.387
R676 VPB.n433 VPB.n428 0.387
R677 VPB.n433 VPB.n423 0.387
R678 VPB.n434 VPB.n433 0.387
R679 VPB.n113 VPB.n112 0.387
R680 VPB.n113 VPB.n108 0.387
R681 VPB.n113 VPB.n103 0.387
R682 VPB.n114 VPB.n113 0.387
R683 VPB.n92 VPB.n91 0.387
R684 VPB.n92 VPB.n87 0.387
R685 VPB.n92 VPB.n82 0.387
R686 VPB.n93 VPB.n92 0.387
R687 VPB.n521 VPB.n520 0.387
R688 VPB.n521 VPB.n516 0.387
R689 VPB.n521 VPB.n511 0.387
R690 VPB.n522 VPB.n521 0.387
R691 VPB.n580 VPB.n579 0.387
R692 VPB.n580 VPB.n575 0.387
R693 VPB.n580 VPB.n570 0.387
R694 VPB.n581 VPB.n580 0.387
R695 VPB.n627 VPB.n626 0.387
R696 VPB.n627 VPB.n622 0.387
R697 VPB.n627 VPB.n617 0.387
R698 VPB.n628 VPB.n627 0.387
R699 VPB.n674 VPB.n673 0.387
R700 VPB.n674 VPB.n669 0.387
R701 VPB.n674 VPB.n664 0.387
R702 VPB.n675 VPB.n674 0.387
R703 VPB.n733 VPB.n732 0.387
R704 VPB.n733 VPB.n728 0.387
R705 VPB.n733 VPB.n723 0.387
R706 VPB.n734 VPB.n733 0.387
R707 VPB.n31 VPB.n30 0.387
R708 VPB.n31 VPB.n26 0.387
R709 VPB.n31 VPB.n21 0.387
R710 VPB.n32 VPB.n31 0.387
R711 VPB.n765 VPB.n13 0.387
R712 VPB.n765 VPB.n9 0.387
R713 VPB.n765 VPB.n4 0.387
R714 VPB.n765 VPB.n764 0.387
R715 VPB.n226 VPB.n199 0.272
R716 VPB.n285 VPB.n258 0.272
R717 VPB.n332 VPB.n305 0.272
R718 VPB.n395 VPB.n368 0.272
R719 VPB.n442 VPB.n415 0.272
R720 VPB.n462 VPB.n461 0.272
R721 VPB.n467 VPB.n466 0.272
R722 VPB.n530 VPB.n503 0.272
R723 VPB.n589 VPB.n562 0.272
R724 VPB.n636 VPB.n609 0.272
R725 VPB.n683 VPB.n656 0.272
R726 VPB.n742 VPB.n715 0.272
R727 VPB.n753 VPB.n752 0.272
R728 VPB.n757 VPB 0.198
R729 VPB.n189 VPB.n185 0.136
R730 VPB.n195 VPB.n189 0.136
R731 VPB.n199 VPB.n195 0.136
R732 VPB.n230 VPB.n226 0.136
R733 VPB.n234 VPB.n230 0.136
R734 VPB.n238 VPB.n234 0.136
R735 VPB.n243 VPB.n238 0.136
R736 VPB.n250 VPB.n243 0.136
R737 VPB.n254 VPB.n250 0.136
R738 VPB.n258 VPB.n254 0.136
R739 VPB.n291 VPB.n285 0.136
R740 VPB.n295 VPB.n291 0.136
R741 VPB.n301 VPB.n295 0.136
R742 VPB.n305 VPB.n301 0.136
R743 VPB.n337 VPB.n332 0.136
R744 VPB.n342 VPB.n337 0.136
R745 VPB.n349 VPB.n342 0.136
R746 VPB.n354 VPB.n349 0.136
R747 VPB.n359 VPB.n354 0.136
R748 VPB.n364 VPB.n359 0.136
R749 VPB.n368 VPB.n364 0.136
R750 VPB.n401 VPB.n395 0.136
R751 VPB.n405 VPB.n401 0.136
R752 VPB.n411 VPB.n405 0.136
R753 VPB.n415 VPB.n411 0.136
R754 VPB.n447 VPB.n442 0.136
R755 VPB.n452 VPB.n447 0.136
R756 VPB.n457 VPB.n452 0.136
R757 VPB.n458 VPB.n457 0.136
R758 VPB.n459 VPB.n458 0.136
R759 VPB.n460 VPB.n459 0.136
R760 VPB.n461 VPB.n460 0.136
R761 VPB.n463 VPB.n462 0.136
R762 VPB.n464 VPB.n463 0.136
R763 VPB.n465 VPB.n464 0.136
R764 VPB.n466 VPB.n465 0.136
R765 VPB.n479 VPB.n475 0.136
R766 VPB.n483 VPB.n479 0.136
R767 VPB.n488 VPB.n483 0.136
R768 VPB.n495 VPB.n488 0.136
R769 VPB.n499 VPB.n495 0.136
R770 VPB.n503 VPB.n499 0.136
R771 VPB.n534 VPB.n530 0.136
R772 VPB.n538 VPB.n534 0.136
R773 VPB.n542 VPB.n538 0.136
R774 VPB.n547 VPB.n542 0.136
R775 VPB.n554 VPB.n547 0.136
R776 VPB.n558 VPB.n554 0.136
R777 VPB.n562 VPB.n558 0.136
R778 VPB.n595 VPB.n589 0.136
R779 VPB.n599 VPB.n595 0.136
R780 VPB.n605 VPB.n599 0.136
R781 VPB.n609 VPB.n605 0.136
R782 VPB.n642 VPB.n636 0.136
R783 VPB.n646 VPB.n642 0.136
R784 VPB.n652 VPB.n646 0.136
R785 VPB.n656 VPB.n652 0.136
R786 VPB.n687 VPB.n683 0.136
R787 VPB.n691 VPB.n687 0.136
R788 VPB.n695 VPB.n691 0.136
R789 VPB.n700 VPB.n695 0.136
R790 VPB.n707 VPB.n700 0.136
R791 VPB.n711 VPB.n707 0.136
R792 VPB.n715 VPB.n711 0.136
R793 VPB.n746 VPB.n742 0.136
R794 VPB.n747 VPB.n746 0.136
R795 VPB.n748 VPB.n747 0.136
R796 VPB.n749 VPB.n748 0.136
R797 VPB.n750 VPB.n749 0.136
R798 VPB.n751 VPB.n750 0.136
R799 VPB.n752 VPB.n751 0.136
R800 VPB.n754 VPB.n753 0.136
R801 VPB.n755 VPB.n754 0.136
R802 VPB.n756 VPB.n755 0.136
R803 VPB.n757 VPB.n756 0.136
R804 VPB.n467 VPB 0.068
R805 VPB.n475 VPB 0.068
R806 a_3027_943.n2 a_3027_943.t5 477.179
R807 a_3027_943.n4 a_3027_943.t3 420.747
R808 a_3027_943.n2 a_3027_943.t4 406.485
R809 a_3027_943.n3 a_3027_943.n2 211.151
R810 a_3027_943.n6 a_3027_943.n4 188.704
R811 a_3027_943.n3 a_3027_943.n1 114.038
R812 a_3027_943.n4 a_3027_943.n3 53.105
R813 a_3027_943.n6 a_3027_943.n5 30
R814 a_3027_943.n7 a_3027_943.n0 24.383
R815 a_3027_943.n7 a_3027_943.n6 23.684
R816 a_3027_943.n1 a_3027_943.t1 14.282
R817 a_3027_943.n1 a_3027_943.t0 14.282
R818 a_807_943.n2 a_807_943.t4 477.179
R819 a_807_943.n4 a_807_943.t5 420.747
R820 a_807_943.n2 a_807_943.t3 406.485
R821 a_807_943.n3 a_807_943.n2 211.151
R822 a_807_943.n6 a_807_943.n4 188.704
R823 a_807_943.n3 a_807_943.n1 114.038
R824 a_807_943.n4 a_807_943.n3 53.105
R825 a_807_943.n6 a_807_943.n5 30
R826 a_807_943.n7 a_807_943.n0 24.383
R827 a_807_943.n7 a_807_943.n6 23.684
R828 a_807_943.n1 a_807_943.t2 14.282
R829 a_807_943.n1 a_807_943.t1 14.282
R830 a_836_182.n2 a_836_182.t14 512.525
R831 a_836_182.n3 a_836_182.t6 480.392
R832 a_836_182.n6 a_836_182.t8 472.359
R833 a_836_182.n3 a_836_182.t12 403.272
R834 a_836_182.n6 a_836_182.t9 384.527
R835 a_836_182.n2 a_836_182.t7 371.139
R836 a_836_182.n4 a_836_182.t11 319.721
R837 a_836_182.n12 a_836_182.n11 242.02
R838 a_836_182.n16 a_836_182.n14 220.281
R839 a_836_182.n7 a_836_182.n6 201.031
R840 a_836_182.n5 a_836_182.n4 153.859
R841 a_836_182.n12 a_836_182.n10 148.471
R842 a_836_182.n14 a_836_182.n1 148.471
R843 a_836_182.n7 a_836_182.t10 141.018
R844 a_836_182.n8 a_836_182.t13 136.079
R845 a_836_182.n8 a_836_182.n7 107.619
R846 a_836_182.n9 a_836_182.n8 107.477
R847 a_836_182.n5 a_836_182.n2 105.194
R848 a_836_182.n13 a_836_182.n9 78.675
R849 a_836_182.n14 a_836_182.n13 78.403
R850 a_836_182.n13 a_836_182.n12 76
R851 a_836_182.n4 a_836_182.n3 55.388
R852 a_836_182.n16 a_836_182.n15 30
R853 a_836_182.n9 a_836_182.n5 26.552
R854 a_836_182.n17 a_836_182.n0 24.383
R855 a_836_182.n17 a_836_182.n16 23.684
R856 a_836_182.n10 a_836_182.t0 14.282
R857 a_836_182.n10 a_836_182.t1 14.282
R858 a_836_182.n1 a_836_182.t2 14.282
R859 a_836_182.n1 a_836_182.t3 14.282
R860 a_575_1004.t1 a_575_1004.n0 101.66
R861 a_575_1004.n0 a_575_1004.t3 101.659
R862 a_575_1004.n0 a_575_1004.t2 14.294
R863 a_575_1004.n0 a_575_1004.t0 14.282
R864 a_2795_1004.t1 a_2795_1004.n0 101.663
R865 a_2795_1004.n0 a_2795_1004.t2 101.661
R866 a_2795_1004.n0 a_2795_1004.t0 14.294
R867 a_2795_1004.n0 a_2795_1004.t3 14.282
R868 a_5291_182.n2 a_5291_182.t3 486.819
R869 a_5291_182.n2 a_5291_182.t4 384.527
R870 a_5291_182.n3 a_5291_182.t5 233.995
R871 a_5291_182.n4 a_5291_182.n1 193.696
R872 a_5291_182.n6 a_5291_182.n4 162.151
R873 a_5291_182.n4 a_5291_182.n3 157.396
R874 a_5291_182.n3 a_5291_182.n2 143.147
R875 a_5291_182.n6 a_5291_182.n5 30
R876 a_5291_182.n7 a_5291_182.n0 24.383
R877 a_5291_182.n7 a_5291_182.n6 23.684
R878 a_5291_182.n1 a_5291_182.t0 14.282
R879 a_5291_182.n1 a_5291_182.t2 14.282
R880 a_6791_1005.n0 a_6791_1005.t0 101.66
R881 a_6791_1005.n0 a_6791_1005.t1 101.66
R882 a_6791_1005.n0 a_6791_1005.t3 14.294
R883 a_6791_1005.t2 a_6791_1005.n0 14.282
R884 a_5767_1004.n4 a_5767_1004.t6 512.525
R885 a_5767_1004.n4 a_5767_1004.t7 371.139
R886 a_5767_1004.n5 a_5767_1004.t5 220.263
R887 a_5767_1004.n8 a_5767_1004.n6 194.086
R888 a_5767_1004.n6 a_5767_1004.n3 162.547
R889 a_5767_1004.n5 a_5767_1004.n4 158.3
R890 a_5767_1004.n6 a_5767_1004.n5 153.043
R891 a_5767_1004.n3 a_5767_1004.n2 76.002
R892 a_5767_1004.n8 a_5767_1004.n7 30
R893 a_5767_1004.n9 a_5767_1004.n0 24.383
R894 a_5767_1004.n9 a_5767_1004.n8 23.684
R895 a_5767_1004.n1 a_5767_1004.t2 14.282
R896 a_5767_1004.n1 a_5767_1004.t1 14.282
R897 a_5767_1004.n2 a_5767_1004.t4 14.282
R898 a_5767_1004.n2 a_5767_1004.t3 14.282
R899 a_5767_1004.n3 a_5767_1004.n1 12.85
R900 VNB VNB.n812 300.778
R901 VNB.n221 VNB.n220 199.897
R902 VNB.n293 VNB.n292 199.897
R903 VNB.n351 VNB.n350 199.897
R904 VNB.n410 VNB.n409 199.897
R905 VNB.n462 VNB.n461 199.897
R906 VNB.n115 VNB.n114 199.897
R907 VNB.n91 VNB.n90 199.897
R908 VNB.n547 VNB.n546 199.897
R909 VNB.n606 VNB.n605 199.897
R910 VNB.n664 VNB.n663 199.897
R911 VNB.n713 VNB.n712 199.897
R912 VNB.n772 VNB.n771 199.897
R913 VNB.n27 VNB.n26 199.897
R914 VNB.n322 VNB.n321 158.304
R915 VNB.n635 VNB.n634 158.304
R916 VNB.n73 VNB.n72 158.304
R917 VNB.n302 VNB.n300 154.509
R918 VNB.n230 VNB.n228 154.509
R919 VNB.n419 VNB.n417 154.509
R920 VNB.n360 VNB.n358 154.509
R921 VNB.n145 VNB.n143 154.509
R922 VNB.n471 VNB.n469 154.509
R923 VNB.n556 VNB.n554 154.509
R924 VNB.n498 VNB.n496 154.509
R925 VNB.n673 VNB.n671 154.509
R926 VNB.n615 VNB.n613 154.509
R927 VNB.n781 VNB.n779 154.509
R928 VNB.n722 VNB.n720 154.509
R929 VNB.n63 VNB.n61 154.509
R930 VNB.n257 VNB.n256 121.366
R931 VNB.n376 VNB.n375 121.366
R932 VNB.n126 VNB.n125 121.366
R933 VNB.n513 VNB.n512 121.366
R934 VNB.n572 VNB.n571 121.366
R935 VNB.n738 VNB.n737 121.366
R936 VNB.n44 VNB.n43 121.366
R937 VNB.n311 VNB.n310 105.536
R938 VNB.n624 VNB.n623 105.536
R939 VNB.n67 VNB.n66 105.536
R940 VNB.n189 VNB.n180 76.136
R941 VNB.n189 VNB.n188 76
R942 VNB.n799 VNB.n798 76
R943 VNB.n787 VNB.n786 76
R944 VNB.n783 VNB.n782 76
R945 VNB.n761 VNB.n760 76
R946 VNB.n757 VNB.n756 76
R947 VNB.n753 VNB.n752 76
R948 VNB.n742 VNB.n741 76
R949 VNB.n736 VNB.n735 76
R950 VNB.n732 VNB.n731 76
R951 VNB.n728 VNB.n727 76
R952 VNB.n724 VNB.n723 76
R953 VNB.n702 VNB.n701 76
R954 VNB.n698 VNB.n697 76
R955 VNB.n690 VNB.n689 76
R956 VNB.n683 VNB.n682 76
R957 VNB.n675 VNB.n674 76
R958 VNB.n653 VNB.n652 76
R959 VNB.n649 VNB.n648 76
R960 VNB.n639 VNB.n638 76
R961 VNB.n627 VNB.n626 76
R962 VNB.n617 VNB.n616 76
R963 VNB.n595 VNB.n594 76
R964 VNB.n591 VNB.n590 76
R965 VNB.n587 VNB.n586 76
R966 VNB.n576 VNB.n575 76
R967 VNB.n570 VNB.n569 76
R968 VNB.n566 VNB.n565 76
R969 VNB.n562 VNB.n561 76
R970 VNB.n558 VNB.n557 76
R971 VNB.n536 VNB.n535 76
R972 VNB.n532 VNB.n531 76
R973 VNB.n528 VNB.n527 76
R974 VNB.n517 VNB.n516 76
R975 VNB.n511 VNB.n510 76
R976 VNB.n507 VNB.n506 76
R977 VNB.n503 VNB.n502 76
R978 VNB.n499 VNB.n495 76
R979 VNB.n485 VNB.n484 76
R980 VNB.n481 VNB.n480 76
R981 VNB.n477 VNB.n476 76
R982 VNB.n473 VNB.n472 76
R983 VNB.n451 VNB.n450 76
R984 VNB.n447 VNB.n446 76
R985 VNB.n439 VNB.n438 76
R986 VNB.n430 VNB.n429 76
R987 VNB.n421 VNB.n420 76
R988 VNB.n399 VNB.n398 76
R989 VNB.n395 VNB.n394 76
R990 VNB.n391 VNB.n390 76
R991 VNB.n380 VNB.n379 76
R992 VNB.n374 VNB.n373 76
R993 VNB.n370 VNB.n369 76
R994 VNB.n366 VNB.n365 76
R995 VNB.n362 VNB.n361 76
R996 VNB.n340 VNB.n339 76
R997 VNB.n336 VNB.n335 76
R998 VNB.n326 VNB.n325 76
R999 VNB.n314 VNB.n313 76
R1000 VNB.n304 VNB.n303 76
R1001 VNB.n282 VNB.n281 76
R1002 VNB.n278 VNB.n277 76
R1003 VNB.n270 VNB.n269 76
R1004 VNB.n261 VNB.n260 76
R1005 VNB.n251 VNB.n250 76
R1006 VNB.n247 VNB.n246 76
R1007 VNB.n240 VNB.n239 76
R1008 VNB.n232 VNB.n231 76
R1009 VNB.n210 VNB.n209 76
R1010 VNB.n206 VNB.n205 76
R1011 VNB.n198 VNB.n197 76
R1012 VNB.n522 VNB.n521 64.194
R1013 VNB.n581 VNB.n580 64.194
R1014 VNB.n747 VNB.n746 64.194
R1015 VNB.n48 VNB.n36 64.194
R1016 VNB.n385 VNB.n384 63.835
R1017 VNB.n130 VNB.n124 63.835
R1018 VNB.n196 VNB.n195 49.896
R1019 VNB.n437 VNB.n436 49.896
R1020 VNB.n272 VNB.t6 39.412
R1021 VNB.n330 VNB.t7 39.412
R1022 VNB.n643 VNB.t5 39.412
R1023 VNB.n7 VNB.t8 39.412
R1024 VNB.n258 VNB.n257 36.937
R1025 VNB.n377 VNB.n376 36.937
R1026 VNB.n127 VNB.n126 36.937
R1027 VNB.n514 VNB.n513 36.937
R1028 VNB.n573 VNB.n572 36.937
R1029 VNB.n739 VNB.n738 36.937
R1030 VNB.n45 VNB.n44 36.937
R1031 VNB.n245 VNB.n244 36.267
R1032 VNB.n184 VNB.n183 35.01
R1033 VNB.n308 VNB.n307 35.01
R1034 VNB.n425 VNB.n424 35.01
R1035 VNB.n621 VNB.n620 35.01
R1036 VNB.n16 VNB.n15 35.01
R1037 VNB.n182 VNB.n181 29.127
R1038 VNB.n423 VNB.n422 29.127
R1039 VNB.n384 VNB.n383 28.421
R1040 VNB.n124 VNB.n123 28.421
R1041 VNB.n521 VNB.n520 28.421
R1042 VNB.n580 VNB.n579 28.421
R1043 VNB.n746 VNB.n745 28.421
R1044 VNB.n36 VNB.n35 28.421
R1045 VNB.n267 VNB.n266 27.855
R1046 VNB.n323 VNB.n320 27.855
R1047 VNB.n388 VNB.n387 27.855
R1048 VNB.n133 VNB.n132 27.855
R1049 VNB.n525 VNB.n524 27.855
R1050 VNB.n584 VNB.n583 27.855
R1051 VNB.n636 VNB.n633 27.855
R1052 VNB.n750 VNB.n749 27.855
R1053 VNB.n51 VNB.n50 27.855
R1054 VNB.n74 VNB.n71 27.855
R1055 VNB.n384 VNB.n382 25.263
R1056 VNB.n124 VNB.n122 25.263
R1057 VNB.n521 VNB.n519 25.263
R1058 VNB.n580 VNB.n578 25.263
R1059 VNB.n746 VNB.n744 25.263
R1060 VNB.n36 VNB.n34 25.263
R1061 VNB.n382 VNB.n381 24.383
R1062 VNB.n122 VNB.n121 24.383
R1063 VNB.n519 VNB.n518 24.383
R1064 VNB.n578 VNB.n577 24.383
R1065 VNB.n744 VNB.n743 24.383
R1066 VNB.n34 VNB.n33 24.383
R1067 VNB.n192 VNB.t13 20.794
R1068 VNB.n433 VNB.t1 20.794
R1069 VNB.n180 VNB.n177 20.452
R1070 VNB.n800 VNB.n799 20.452
R1071 VNB.n185 VNB.n184 20.094
R1072 VNB.n194 VNB.n193 20.094
R1073 VNB.n202 VNB.n201 20.094
R1074 VNB.n309 VNB.n308 20.094
R1075 VNB.n319 VNB.n318 20.094
R1076 VNB.n332 VNB.n331 20.094
R1077 VNB.n426 VNB.n425 20.094
R1078 VNB.n435 VNB.n434 20.094
R1079 VNB.n443 VNB.n442 20.094
R1080 VNB.n147 VNB.n104 20.094
R1081 VNB.n154 VNB.n101 20.094
R1082 VNB.n158 VNB.n99 20.094
R1083 VNB.n622 VNB.n621 20.094
R1084 VNB.n632 VNB.n631 20.094
R1085 VNB.n645 VNB.n644 20.094
R1086 VNB.n679 VNB.n678 20.094
R1087 VNB.n686 VNB.n685 20.094
R1088 VNB.n694 VNB.n693 20.094
R1089 VNB.n65 VNB.n16 20.094
R1090 VNB.n70 VNB.n12 20.094
R1091 VNB.n80 VNB.n8 20.094
R1092 VNB.n264 VNB.n263 19.735
R1093 VNB.n255 VNB.n254 19.735
R1094 VNB.n243 VNB.n242 19.735
R1095 VNB.n236 VNB.n235 19.735
R1096 VNB.n274 VNB.n273 19.735
R1097 VNB.n242 VNB.t14 19.724
R1098 VNB.n184 VNB.n182 19.017
R1099 VNB.n308 VNB.n306 19.017
R1100 VNB.n425 VNB.n423 19.017
R1101 VNB.n621 VNB.n619 19.017
R1102 VNB.n16 VNB.n14 19.017
R1103 VNB.n684 VNB.t12 18.552
R1104 VNB.n152 VNB.n151 18.269
R1105 VNB.n688 VNB.n687 18.269
R1106 VNB.n98 VNB.t2 17.595
R1107 VNB.n272 VNB.n271 17.185
R1108 VNB.n330 VNB.n329 17.185
R1109 VNB.n643 VNB.n642 17.185
R1110 VNB.n7 VNB.n6 17.185
R1111 VNB.n268 VNB.n267 16.721
R1112 VNB.n324 VNB.n323 16.721
R1113 VNB.n389 VNB.n388 16.721
R1114 VNB.n134 VNB.n133 16.721
R1115 VNB.n526 VNB.n525 16.721
R1116 VNB.n585 VNB.n584 16.721
R1117 VNB.n637 VNB.n636 16.721
R1118 VNB.n751 VNB.n750 16.721
R1119 VNB.n52 VNB.n51 16.721
R1120 VNB.n75 VNB.n74 16.721
R1121 VNB.n253 VNB.n252 13.654
R1122 VNB.n188 VNB.n187 13.653
R1123 VNB.n187 VNB.n186 13.653
R1124 VNB.n197 VNB.n196 13.653
R1125 VNB.n205 VNB.n204 13.653
R1126 VNB.n204 VNB.n203 13.653
R1127 VNB.n209 VNB.n208 13.653
R1128 VNB.n208 VNB.n207 13.653
R1129 VNB.n231 VNB.n230 13.653
R1130 VNB.n230 VNB.n229 13.653
R1131 VNB.n239 VNB.n238 13.653
R1132 VNB.n238 VNB.n237 13.653
R1133 VNB.n246 VNB.n245 13.653
R1134 VNB.n250 VNB.n249 13.653
R1135 VNB.n249 VNB.n248 13.653
R1136 VNB.n260 VNB.n259 13.653
R1137 VNB.n259 VNB.n258 13.653
R1138 VNB.n269 VNB.n268 13.653
R1139 VNB.n277 VNB.n276 13.653
R1140 VNB.n276 VNB.n275 13.653
R1141 VNB.n281 VNB.n280 13.653
R1142 VNB.n280 VNB.n279 13.653
R1143 VNB.n303 VNB.n302 13.653
R1144 VNB.n302 VNB.n301 13.653
R1145 VNB.n313 VNB.n312 13.653
R1146 VNB.n312 VNB.n311 13.653
R1147 VNB.n325 VNB.n324 13.653
R1148 VNB.n335 VNB.n334 13.653
R1149 VNB.n334 VNB.n333 13.653
R1150 VNB.n339 VNB.n338 13.653
R1151 VNB.n338 VNB.n337 13.653
R1152 VNB.n361 VNB.n360 13.653
R1153 VNB.n360 VNB.n359 13.653
R1154 VNB.n365 VNB.n364 13.653
R1155 VNB.n364 VNB.n363 13.653
R1156 VNB.n369 VNB.n368 13.653
R1157 VNB.n368 VNB.n367 13.653
R1158 VNB.n373 VNB.n372 13.653
R1159 VNB.n372 VNB.n371 13.653
R1160 VNB.n379 VNB.n378 13.653
R1161 VNB.n378 VNB.n377 13.653
R1162 VNB.n390 VNB.n389 13.653
R1163 VNB.n394 VNB.n393 13.653
R1164 VNB.n393 VNB.n392 13.653
R1165 VNB.n398 VNB.n397 13.653
R1166 VNB.n397 VNB.n396 13.653
R1167 VNB.n420 VNB.n419 13.653
R1168 VNB.n419 VNB.n418 13.653
R1169 VNB.n429 VNB.n428 13.653
R1170 VNB.n428 VNB.n427 13.653
R1171 VNB.n438 VNB.n437 13.653
R1172 VNB.n446 VNB.n445 13.653
R1173 VNB.n445 VNB.n444 13.653
R1174 VNB.n450 VNB.n449 13.653
R1175 VNB.n449 VNB.n448 13.653
R1176 VNB.n472 VNB.n471 13.653
R1177 VNB.n471 VNB.n470 13.653
R1178 VNB.n476 VNB.n475 13.653
R1179 VNB.n475 VNB.n474 13.653
R1180 VNB.n480 VNB.n479 13.653
R1181 VNB.n479 VNB.n478 13.653
R1182 VNB.n484 VNB.n483 13.653
R1183 VNB.n483 VNB.n482 13.653
R1184 VNB.n129 VNB.n128 13.653
R1185 VNB.n128 VNB.n127 13.653
R1186 VNB.n135 VNB.n134 13.653
R1187 VNB.n138 VNB.n137 13.653
R1188 VNB.n137 VNB.n136 13.653
R1189 VNB.n141 VNB.n140 13.653
R1190 VNB.n140 VNB.n139 13.653
R1191 VNB.n146 VNB.n145 13.653
R1192 VNB.n145 VNB.n144 13.653
R1193 VNB.n150 VNB.n149 13.653
R1194 VNB.n149 VNB.n148 13.653
R1195 VNB.n153 VNB.n152 13.653
R1196 VNB.n157 VNB.n156 13.653
R1197 VNB.n156 VNB.n155 13.653
R1198 VNB.n161 VNB.n160 13.653
R1199 VNB.n160 VNB.n159 13.653
R1200 VNB.n499 VNB.n498 13.653
R1201 VNB.n498 VNB.n497 13.653
R1202 VNB.n502 VNB.n501 13.653
R1203 VNB.n501 VNB.n500 13.653
R1204 VNB.n506 VNB.n505 13.653
R1205 VNB.n505 VNB.n504 13.653
R1206 VNB.n510 VNB.n509 13.653
R1207 VNB.n509 VNB.n508 13.653
R1208 VNB.n516 VNB.n515 13.653
R1209 VNB.n515 VNB.n514 13.653
R1210 VNB.n527 VNB.n526 13.653
R1211 VNB.n531 VNB.n530 13.653
R1212 VNB.n530 VNB.n529 13.653
R1213 VNB.n535 VNB.n534 13.653
R1214 VNB.n534 VNB.n533 13.653
R1215 VNB.n557 VNB.n556 13.653
R1216 VNB.n556 VNB.n555 13.653
R1217 VNB.n561 VNB.n560 13.653
R1218 VNB.n560 VNB.n559 13.653
R1219 VNB.n565 VNB.n564 13.653
R1220 VNB.n564 VNB.n563 13.653
R1221 VNB.n569 VNB.n568 13.653
R1222 VNB.n568 VNB.n567 13.653
R1223 VNB.n575 VNB.n574 13.653
R1224 VNB.n574 VNB.n573 13.653
R1225 VNB.n586 VNB.n585 13.653
R1226 VNB.n590 VNB.n589 13.653
R1227 VNB.n589 VNB.n588 13.653
R1228 VNB.n594 VNB.n593 13.653
R1229 VNB.n593 VNB.n592 13.653
R1230 VNB.n616 VNB.n615 13.653
R1231 VNB.n615 VNB.n614 13.653
R1232 VNB.n626 VNB.n625 13.653
R1233 VNB.n625 VNB.n624 13.653
R1234 VNB.n638 VNB.n637 13.653
R1235 VNB.n648 VNB.n647 13.653
R1236 VNB.n647 VNB.n646 13.653
R1237 VNB.n652 VNB.n651 13.653
R1238 VNB.n651 VNB.n650 13.653
R1239 VNB.n674 VNB.n673 13.653
R1240 VNB.n673 VNB.n672 13.653
R1241 VNB.n682 VNB.n681 13.653
R1242 VNB.n681 VNB.n680 13.653
R1243 VNB.n689 VNB.n688 13.653
R1244 VNB.n697 VNB.n696 13.653
R1245 VNB.n696 VNB.n695 13.653
R1246 VNB.n701 VNB.n700 13.653
R1247 VNB.n700 VNB.n699 13.653
R1248 VNB.n723 VNB.n722 13.653
R1249 VNB.n722 VNB.n721 13.653
R1250 VNB.n727 VNB.n726 13.653
R1251 VNB.n726 VNB.n725 13.653
R1252 VNB.n731 VNB.n730 13.653
R1253 VNB.n730 VNB.n729 13.653
R1254 VNB.n735 VNB.n734 13.653
R1255 VNB.n734 VNB.n733 13.653
R1256 VNB.n741 VNB.n740 13.653
R1257 VNB.n740 VNB.n739 13.653
R1258 VNB.n752 VNB.n751 13.653
R1259 VNB.n756 VNB.n755 13.653
R1260 VNB.n755 VNB.n754 13.653
R1261 VNB.n760 VNB.n759 13.653
R1262 VNB.n759 VNB.n758 13.653
R1263 VNB.n782 VNB.n781 13.653
R1264 VNB.n781 VNB.n780 13.653
R1265 VNB.n786 VNB.n785 13.653
R1266 VNB.n785 VNB.n784 13.653
R1267 VNB.n39 VNB.n38 13.653
R1268 VNB.n38 VNB.n37 13.653
R1269 VNB.n42 VNB.n41 13.653
R1270 VNB.n41 VNB.n40 13.653
R1271 VNB.n47 VNB.n46 13.653
R1272 VNB.n46 VNB.n45 13.653
R1273 VNB.n53 VNB.n52 13.653
R1274 VNB.n56 VNB.n55 13.653
R1275 VNB.n55 VNB.n54 13.653
R1276 VNB.n59 VNB.n58 13.653
R1277 VNB.n58 VNB.n57 13.653
R1278 VNB.n64 VNB.n63 13.653
R1279 VNB.n63 VNB.n62 13.653
R1280 VNB.n69 VNB.n68 13.653
R1281 VNB.n68 VNB.n67 13.653
R1282 VNB.n76 VNB.n75 13.653
R1283 VNB.n79 VNB.n78 13.653
R1284 VNB.n78 VNB.n77 13.653
R1285 VNB.n799 VNB.n0 13.653
R1286 VNB VNB.n0 13.653
R1287 VNB.n180 VNB.n179 13.653
R1288 VNB.n179 VNB.n178 13.653
R1289 VNB.n99 VNB.n98 13.608
R1290 VNB.n693 VNB.n692 13.608
R1291 VNB.n807 VNB.n804 13.577
R1292 VNB.n165 VNB.n163 13.276
R1293 VNB.n177 VNB.n165 13.276
R1294 VNB.n213 VNB.n211 13.276
R1295 VNB.n226 VNB.n213 13.276
R1296 VNB.n285 VNB.n283 13.276
R1297 VNB.n298 VNB.n285 13.276
R1298 VNB.n343 VNB.n341 13.276
R1299 VNB.n356 VNB.n343 13.276
R1300 VNB.n402 VNB.n400 13.276
R1301 VNB.n415 VNB.n402 13.276
R1302 VNB.n454 VNB.n452 13.276
R1303 VNB.n467 VNB.n454 13.276
R1304 VNB.n107 VNB.n105 13.276
R1305 VNB.n120 VNB.n107 13.276
R1306 VNB.n83 VNB.n81 13.276
R1307 VNB.n96 VNB.n83 13.276
R1308 VNB.n539 VNB.n537 13.276
R1309 VNB.n552 VNB.n539 13.276
R1310 VNB.n598 VNB.n596 13.276
R1311 VNB.n611 VNB.n598 13.276
R1312 VNB.n656 VNB.n654 13.276
R1313 VNB.n669 VNB.n656 13.276
R1314 VNB.n705 VNB.n703 13.276
R1315 VNB.n718 VNB.n705 13.276
R1316 VNB.n764 VNB.n762 13.276
R1317 VNB.n777 VNB.n764 13.276
R1318 VNB.n19 VNB.n17 13.276
R1319 VNB.n32 VNB.n19 13.276
R1320 VNB.n231 VNB.n227 13.276
R1321 VNB.n303 VNB.n299 13.276
R1322 VNB.n361 VNB.n357 13.276
R1323 VNB.n420 VNB.n416 13.276
R1324 VNB.n472 VNB.n468 13.276
R1325 VNB.n138 VNB.n135 13.276
R1326 VNB.n141 VNB.n138 13.276
R1327 VNB.n142 VNB.n141 13.276
R1328 VNB.n146 VNB.n142 13.276
R1329 VNB.n153 VNB.n150 13.276
R1330 VNB.n162 VNB.n161 13.276
R1331 VNB.n499 VNB.n162 13.276
R1332 VNB.n502 VNB.n499 13.276
R1333 VNB.n557 VNB.n553 13.276
R1334 VNB.n616 VNB.n612 13.276
R1335 VNB.n674 VNB.n670 13.276
R1336 VNB.n723 VNB.n719 13.276
R1337 VNB.n782 VNB.n778 13.276
R1338 VNB.n42 VNB.n39 13.276
R1339 VNB.n47 VNB.n42 13.276
R1340 VNB.n56 VNB.n53 13.276
R1341 VNB.n59 VNB.n56 13.276
R1342 VNB.n60 VNB.n59 13.276
R1343 VNB.n64 VNB.n60 13.276
R1344 VNB.n79 VNB.n76 13.276
R1345 VNB.n3 VNB.n1 13.276
R1346 VNB.n800 VNB.n3 13.276
R1347 VNB.n157 VNB.n154 13.097
R1348 VNB.n70 VNB.n69 13.097
R1349 VNB.n201 VNB.n200 12.837
R1350 VNB.n442 VNB.n441 12.837
R1351 VNB.n235 VNB.n234 11.605
R1352 VNB.n104 VNB.n103 10.853
R1353 VNB.n678 VNB.n677 10.853
R1354 VNB.n130 VNB.n129 10.764
R1355 VNB.n48 VNB.n47 10.764
R1356 VNB.n103 VNB.n102 10.417
R1357 VNB.n677 VNB.n676 10.417
R1358 VNB.n234 VNB.n233 9.809
R1359 VNB.n147 VNB.n146 9.329
R1360 VNB.n799 VNB.n80 9.329
R1361 VNB.n161 VNB.n158 8.97
R1362 VNB.n65 VNB.n64 8.97
R1363 VNB.n98 VNB.n97 7.858
R1364 VNB.n692 VNB.n691 7.858
R1365 VNB.n200 VNB.n199 7.566
R1366 VNB.n441 VNB.n440 7.566
R1367 VNB.n263 VNB.n262 7.5
R1368 VNB.n306 VNB.n305 7.5
R1369 VNB.n317 VNB.n316 7.5
R1370 VNB.n619 VNB.n618 7.5
R1371 VNB.n630 VNB.n629 7.5
R1372 VNB.n14 VNB.n13 7.5
R1373 VNB.n11 VNB.n10 7.5
R1374 VNB.n809 VNB.n808 7.5
R1375 VNB.n219 VNB.n218 7.5
R1376 VNB.n215 VNB.n214 7.5
R1377 VNB.n213 VNB.n212 7.5
R1378 VNB.n226 VNB.n225 7.5
R1379 VNB.n291 VNB.n290 7.5
R1380 VNB.n287 VNB.n286 7.5
R1381 VNB.n285 VNB.n284 7.5
R1382 VNB.n298 VNB.n297 7.5
R1383 VNB.n349 VNB.n348 7.5
R1384 VNB.n345 VNB.n344 7.5
R1385 VNB.n343 VNB.n342 7.5
R1386 VNB.n356 VNB.n355 7.5
R1387 VNB.n408 VNB.n407 7.5
R1388 VNB.n404 VNB.n403 7.5
R1389 VNB.n402 VNB.n401 7.5
R1390 VNB.n415 VNB.n414 7.5
R1391 VNB.n460 VNB.n459 7.5
R1392 VNB.n456 VNB.n455 7.5
R1393 VNB.n454 VNB.n453 7.5
R1394 VNB.n467 VNB.n466 7.5
R1395 VNB.n113 VNB.n112 7.5
R1396 VNB.n109 VNB.n108 7.5
R1397 VNB.n107 VNB.n106 7.5
R1398 VNB.n120 VNB.n119 7.5
R1399 VNB.n89 VNB.n88 7.5
R1400 VNB.n85 VNB.n84 7.5
R1401 VNB.n83 VNB.n82 7.5
R1402 VNB.n96 VNB.n95 7.5
R1403 VNB.n545 VNB.n544 7.5
R1404 VNB.n541 VNB.n540 7.5
R1405 VNB.n539 VNB.n538 7.5
R1406 VNB.n552 VNB.n551 7.5
R1407 VNB.n604 VNB.n603 7.5
R1408 VNB.n600 VNB.n599 7.5
R1409 VNB.n598 VNB.n597 7.5
R1410 VNB.n611 VNB.n610 7.5
R1411 VNB.n662 VNB.n661 7.5
R1412 VNB.n658 VNB.n657 7.5
R1413 VNB.n656 VNB.n655 7.5
R1414 VNB.n669 VNB.n668 7.5
R1415 VNB.n711 VNB.n710 7.5
R1416 VNB.n707 VNB.n706 7.5
R1417 VNB.n705 VNB.n704 7.5
R1418 VNB.n718 VNB.n717 7.5
R1419 VNB.n770 VNB.n769 7.5
R1420 VNB.n766 VNB.n765 7.5
R1421 VNB.n764 VNB.n763 7.5
R1422 VNB.n777 VNB.n776 7.5
R1423 VNB.n25 VNB.n24 7.5
R1424 VNB.n21 VNB.n20 7.5
R1425 VNB.n19 VNB.n18 7.5
R1426 VNB.n32 VNB.n31 7.5
R1427 VNB.n801 VNB.n800 7.5
R1428 VNB.n3 VNB.n2 7.5
R1429 VNB.n806 VNB.n805 7.5
R1430 VNB.n171 VNB.n170 7.5
R1431 VNB.n167 VNB.n166 7.5
R1432 VNB.n165 VNB.n164 7.5
R1433 VNB.n177 VNB.n176 7.5
R1434 VNB.n227 VNB.n226 7.176
R1435 VNB.n299 VNB.n298 7.176
R1436 VNB.n357 VNB.n356 7.176
R1437 VNB.n416 VNB.n415 7.176
R1438 VNB.n468 VNB.n467 7.176
R1439 VNB.n142 VNB.n120 7.176
R1440 VNB.n162 VNB.n96 7.176
R1441 VNB.n553 VNB.n552 7.176
R1442 VNB.n612 VNB.n611 7.176
R1443 VNB.n670 VNB.n669 7.176
R1444 VNB.n719 VNB.n718 7.176
R1445 VNB.n778 VNB.n777 7.176
R1446 VNB.n60 VNB.n32 7.176
R1447 VNB.t14 VNB.n241 7.04
R1448 VNB.n811 VNB.n809 7.011
R1449 VNB.n222 VNB.n219 7.011
R1450 VNB.n217 VNB.n215 7.011
R1451 VNB.n294 VNB.n291 7.011
R1452 VNB.n289 VNB.n287 7.011
R1453 VNB.n352 VNB.n349 7.011
R1454 VNB.n347 VNB.n345 7.011
R1455 VNB.n411 VNB.n408 7.011
R1456 VNB.n406 VNB.n404 7.011
R1457 VNB.n463 VNB.n460 7.011
R1458 VNB.n458 VNB.n456 7.011
R1459 VNB.n116 VNB.n113 7.011
R1460 VNB.n111 VNB.n109 7.011
R1461 VNB.n92 VNB.n89 7.011
R1462 VNB.n87 VNB.n85 7.011
R1463 VNB.n548 VNB.n545 7.011
R1464 VNB.n543 VNB.n541 7.011
R1465 VNB.n607 VNB.n604 7.011
R1466 VNB.n602 VNB.n600 7.011
R1467 VNB.n665 VNB.n662 7.011
R1468 VNB.n660 VNB.n658 7.011
R1469 VNB.n714 VNB.n711 7.011
R1470 VNB.n709 VNB.n707 7.011
R1471 VNB.n773 VNB.n770 7.011
R1472 VNB.n768 VNB.n766 7.011
R1473 VNB.n28 VNB.n25 7.011
R1474 VNB.n23 VNB.n21 7.011
R1475 VNB.n173 VNB.n171 7.011
R1476 VNB.n169 VNB.n167 7.011
R1477 VNB.n225 VNB.n224 7.01
R1478 VNB.n217 VNB.n216 7.01
R1479 VNB.n222 VNB.n221 7.01
R1480 VNB.n297 VNB.n296 7.01
R1481 VNB.n289 VNB.n288 7.01
R1482 VNB.n294 VNB.n293 7.01
R1483 VNB.n355 VNB.n354 7.01
R1484 VNB.n347 VNB.n346 7.01
R1485 VNB.n352 VNB.n351 7.01
R1486 VNB.n414 VNB.n413 7.01
R1487 VNB.n406 VNB.n405 7.01
R1488 VNB.n411 VNB.n410 7.01
R1489 VNB.n466 VNB.n465 7.01
R1490 VNB.n458 VNB.n457 7.01
R1491 VNB.n463 VNB.n462 7.01
R1492 VNB.n119 VNB.n118 7.01
R1493 VNB.n111 VNB.n110 7.01
R1494 VNB.n116 VNB.n115 7.01
R1495 VNB.n95 VNB.n94 7.01
R1496 VNB.n87 VNB.n86 7.01
R1497 VNB.n92 VNB.n91 7.01
R1498 VNB.n551 VNB.n550 7.01
R1499 VNB.n543 VNB.n542 7.01
R1500 VNB.n548 VNB.n547 7.01
R1501 VNB.n610 VNB.n609 7.01
R1502 VNB.n602 VNB.n601 7.01
R1503 VNB.n607 VNB.n606 7.01
R1504 VNB.n668 VNB.n667 7.01
R1505 VNB.n660 VNB.n659 7.01
R1506 VNB.n665 VNB.n664 7.01
R1507 VNB.n717 VNB.n716 7.01
R1508 VNB.n709 VNB.n708 7.01
R1509 VNB.n714 VNB.n713 7.01
R1510 VNB.n776 VNB.n775 7.01
R1511 VNB.n768 VNB.n767 7.01
R1512 VNB.n773 VNB.n772 7.01
R1513 VNB.n31 VNB.n30 7.01
R1514 VNB.n23 VNB.n22 7.01
R1515 VNB.n28 VNB.n27 7.01
R1516 VNB.n176 VNB.n175 7.01
R1517 VNB.n169 VNB.n168 7.01
R1518 VNB.n173 VNB.n172 7.01
R1519 VNB.n811 VNB.n810 7.01
R1520 VNB.n807 VNB.n806 6.788
R1521 VNB.n802 VNB.n801 6.788
R1522 VNB.n260 VNB.n255 6.638
R1523 VNB.n273 VNB.n272 6.139
R1524 VNB.n331 VNB.n330 6.139
R1525 VNB.n644 VNB.n643 6.139
R1526 VNB.n8 VNB.n7 6.139
R1527 VNB.n254 VNB.n253 5.774
R1528 VNB.n191 VNB.n190 4.551
R1529 VNB.n328 VNB.n327 4.551
R1530 VNB.n432 VNB.n431 4.551
R1531 VNB.n641 VNB.n640 4.551
R1532 VNB.n5 VNB.n4 4.551
R1533 VNB.n188 VNB.n185 4.305
R1534 VNB.n313 VNB.n309 4.305
R1535 VNB.n429 VNB.n426 4.305
R1536 VNB.n158 VNB.n157 4.305
R1537 VNB.n626 VNB.n622 4.305
R1538 VNB.n697 VNB.n694 4.305
R1539 VNB.n69 VNB.n65 4.305
R1540 VNB.n205 VNB.n202 3.947
R1541 VNB.n335 VNB.n332 3.947
R1542 VNB.n446 VNB.n443 3.947
R1543 VNB.n150 VNB.n147 3.947
R1544 VNB.n648 VNB.n645 3.947
R1545 VNB.n682 VNB.n679 3.947
R1546 VNB.n80 VNB.n79 3.947
R1547 VNB.n246 VNB.n243 2.511
R1548 VNB.n269 VNB.n264 2.511
R1549 VNB.n390 VNB.n385 2.511
R1550 VNB.n135 VNB.n130 2.511
R1551 VNB.n527 VNB.n522 2.511
R1552 VNB.n586 VNB.n581 2.511
R1553 VNB.n752 VNB.n747 2.511
R1554 VNB.n53 VNB.n48 2.511
R1555 VNB.t13 VNB.n191 2.238
R1556 VNB.t7 VNB.n328 2.238
R1557 VNB.t1 VNB.n432 2.238
R1558 VNB.t5 VNB.n641 2.238
R1559 VNB.t8 VNB.n5 2.238
R1560 VNB.n267 VNB.n265 1.99
R1561 VNB.n323 VNB.n322 1.99
R1562 VNB.n388 VNB.n386 1.99
R1563 VNB.n133 VNB.n131 1.99
R1564 VNB.n525 VNB.n523 1.99
R1565 VNB.n584 VNB.n582 1.99
R1566 VNB.n636 VNB.n635 1.99
R1567 VNB.n750 VNB.n748 1.99
R1568 VNB.n51 VNB.n49 1.99
R1569 VNB.n74 VNB.n73 1.99
R1570 VNB.n316 VNB.n315 1.935
R1571 VNB.n629 VNB.n628 1.935
R1572 VNB.n10 VNB.n9 1.935
R1573 VNB.n239 VNB.n236 1.614
R1574 VNB.n277 VNB.n274 1.614
R1575 VNB.n812 VNB.n803 0.921
R1576 VNB.n812 VNB.n807 0.476
R1577 VNB.n812 VNB.n802 0.475
R1578 VNB.n193 VNB.n192 0.358
R1579 VNB.n318 VNB.n317 0.358
R1580 VNB.n434 VNB.n433 0.358
R1581 VNB.n101 VNB.n100 0.358
R1582 VNB.n631 VNB.n630 0.358
R1583 VNB.n685 VNB.n684 0.358
R1584 VNB.n12 VNB.n11 0.358
R1585 VNB.n232 VNB.n210 0.272
R1586 VNB.n304 VNB.n282 0.272
R1587 VNB.n362 VNB.n340 0.272
R1588 VNB.n421 VNB.n399 0.272
R1589 VNB.n473 VNB.n451 0.272
R1590 VNB.n490 VNB.n489 0.272
R1591 VNB.n495 VNB.n494 0.272
R1592 VNB.n558 VNB.n536 0.272
R1593 VNB.n617 VNB.n595 0.272
R1594 VNB.n675 VNB.n653 0.272
R1595 VNB.n724 VNB.n702 0.272
R1596 VNB.n783 VNB.n761 0.272
R1597 VNB.n794 VNB.n793 0.272
R1598 VNB.n223 VNB.n217 0.246
R1599 VNB.n224 VNB.n223 0.246
R1600 VNB.n223 VNB.n222 0.246
R1601 VNB.n295 VNB.n289 0.246
R1602 VNB.n296 VNB.n295 0.246
R1603 VNB.n295 VNB.n294 0.246
R1604 VNB.n353 VNB.n347 0.246
R1605 VNB.n354 VNB.n353 0.246
R1606 VNB.n353 VNB.n352 0.246
R1607 VNB.n412 VNB.n406 0.246
R1608 VNB.n413 VNB.n412 0.246
R1609 VNB.n412 VNB.n411 0.246
R1610 VNB.n464 VNB.n458 0.246
R1611 VNB.n465 VNB.n464 0.246
R1612 VNB.n464 VNB.n463 0.246
R1613 VNB.n117 VNB.n111 0.246
R1614 VNB.n118 VNB.n117 0.246
R1615 VNB.n117 VNB.n116 0.246
R1616 VNB.n93 VNB.n87 0.246
R1617 VNB.n94 VNB.n93 0.246
R1618 VNB.n93 VNB.n92 0.246
R1619 VNB.n549 VNB.n543 0.246
R1620 VNB.n550 VNB.n549 0.246
R1621 VNB.n549 VNB.n548 0.246
R1622 VNB.n608 VNB.n602 0.246
R1623 VNB.n609 VNB.n608 0.246
R1624 VNB.n608 VNB.n607 0.246
R1625 VNB.n666 VNB.n660 0.246
R1626 VNB.n667 VNB.n666 0.246
R1627 VNB.n666 VNB.n665 0.246
R1628 VNB.n715 VNB.n709 0.246
R1629 VNB.n716 VNB.n715 0.246
R1630 VNB.n715 VNB.n714 0.246
R1631 VNB.n774 VNB.n768 0.246
R1632 VNB.n775 VNB.n774 0.246
R1633 VNB.n774 VNB.n773 0.246
R1634 VNB.n29 VNB.n23 0.246
R1635 VNB.n30 VNB.n29 0.246
R1636 VNB.n29 VNB.n28 0.246
R1637 VNB.n174 VNB.n169 0.246
R1638 VNB.n175 VNB.n174 0.246
R1639 VNB.n174 VNB.n173 0.246
R1640 VNB.n812 VNB.n811 0.246
R1641 VNB.n798 VNB 0.198
R1642 VNB.n197 VNB.n194 0.179
R1643 VNB.n325 VNB.n319 0.179
R1644 VNB.n438 VNB.n435 0.179
R1645 VNB.n154 VNB.n153 0.179
R1646 VNB.n638 VNB.n632 0.179
R1647 VNB.n689 VNB.n686 0.179
R1648 VNB.n76 VNB.n70 0.179
R1649 VNB.n198 VNB.n189 0.136
R1650 VNB.n206 VNB.n198 0.136
R1651 VNB.n210 VNB.n206 0.136
R1652 VNB.n240 VNB.n232 0.136
R1653 VNB.n247 VNB.n240 0.136
R1654 VNB.n251 VNB.n247 0.136
R1655 VNB.n261 VNB.n251 0.136
R1656 VNB.n270 VNB.n261 0.136
R1657 VNB.n278 VNB.n270 0.136
R1658 VNB.n282 VNB.n278 0.136
R1659 VNB.n314 VNB.n304 0.136
R1660 VNB.n326 VNB.n314 0.136
R1661 VNB.n336 VNB.n326 0.136
R1662 VNB.n340 VNB.n336 0.136
R1663 VNB.n366 VNB.n362 0.136
R1664 VNB.n370 VNB.n366 0.136
R1665 VNB.n374 VNB.n370 0.136
R1666 VNB.n380 VNB.n374 0.136
R1667 VNB.n391 VNB.n380 0.136
R1668 VNB.n395 VNB.n391 0.136
R1669 VNB.n399 VNB.n395 0.136
R1670 VNB.n430 VNB.n421 0.136
R1671 VNB.n439 VNB.n430 0.136
R1672 VNB.n447 VNB.n439 0.136
R1673 VNB.n451 VNB.n447 0.136
R1674 VNB.n477 VNB.n473 0.136
R1675 VNB.n481 VNB.n477 0.136
R1676 VNB.n485 VNB.n481 0.136
R1677 VNB.n486 VNB.n485 0.136
R1678 VNB.n487 VNB.n486 0.136
R1679 VNB.n488 VNB.n487 0.136
R1680 VNB.n489 VNB.n488 0.136
R1681 VNB.n491 VNB.n490 0.136
R1682 VNB.n492 VNB.n491 0.136
R1683 VNB.n493 VNB.n492 0.136
R1684 VNB.n494 VNB.n493 0.136
R1685 VNB.n507 VNB.n503 0.136
R1686 VNB.n511 VNB.n507 0.136
R1687 VNB.n517 VNB.n511 0.136
R1688 VNB.n528 VNB.n517 0.136
R1689 VNB.n532 VNB.n528 0.136
R1690 VNB.n536 VNB.n532 0.136
R1691 VNB.n562 VNB.n558 0.136
R1692 VNB.n566 VNB.n562 0.136
R1693 VNB.n570 VNB.n566 0.136
R1694 VNB.n576 VNB.n570 0.136
R1695 VNB.n587 VNB.n576 0.136
R1696 VNB.n591 VNB.n587 0.136
R1697 VNB.n595 VNB.n591 0.136
R1698 VNB.n627 VNB.n617 0.136
R1699 VNB.n639 VNB.n627 0.136
R1700 VNB.n649 VNB.n639 0.136
R1701 VNB.n653 VNB.n649 0.136
R1702 VNB.n683 VNB.n675 0.136
R1703 VNB.n690 VNB.n683 0.136
R1704 VNB.n698 VNB.n690 0.136
R1705 VNB.n702 VNB.n698 0.136
R1706 VNB.n728 VNB.n724 0.136
R1707 VNB.n732 VNB.n728 0.136
R1708 VNB.n736 VNB.n732 0.136
R1709 VNB.n742 VNB.n736 0.136
R1710 VNB.n753 VNB.n742 0.136
R1711 VNB.n757 VNB.n753 0.136
R1712 VNB.n761 VNB.n757 0.136
R1713 VNB.n787 VNB.n783 0.136
R1714 VNB.n788 VNB.n787 0.136
R1715 VNB.n789 VNB.n788 0.136
R1716 VNB.n790 VNB.n789 0.136
R1717 VNB.n791 VNB.n790 0.136
R1718 VNB.n792 VNB.n791 0.136
R1719 VNB.n793 VNB.n792 0.136
R1720 VNB.n795 VNB.n794 0.136
R1721 VNB.n796 VNB.n795 0.136
R1722 VNB.n797 VNB.n796 0.136
R1723 VNB.n798 VNB.n797 0.136
R1724 VNB.n495 VNB 0.068
R1725 VNB.n503 VNB 0.068
R1726 a_6401_182.n1 a_6401_182.t3 470.752
R1727 a_6401_182.n1 a_6401_182.t5 384.527
R1728 a_6401_182.n2 a_6401_182.t4 224.666
R1729 a_6401_182.n5 a_6401_182.n3 195.226
R1730 a_6401_182.n3 a_6401_182.n0 167.143
R1731 a_6401_182.n3 a_6401_182.n2 153.859
R1732 a_6401_182.n2 a_6401_182.n1 120.22
R1733 a_6401_182.n5 a_6401_182.n4 15.218
R1734 a_6401_182.n0 a_6401_182.t2 14.282
R1735 a_6401_182.n0 a_6401_182.t1 14.282
R1736 a_6401_182.n6 a_6401_182.n5 12.014
R1737 a_1241_1004.t2 a_1241_1004.n0 101.66
R1738 a_1241_1004.n0 a_1241_1004.t0 101.659
R1739 a_1241_1004.n0 a_1241_1004.t1 14.294
R1740 a_1241_1004.n0 a_1241_1004.t3 14.282
R1741 a_185_182.n1 a_185_182.t5 477.179
R1742 a_185_182.n1 a_185_182.t4 406.485
R1743 a_185_182.n2 a_185_182.t3 225.731
R1744 a_185_182.n3 a_185_182.n0 220.249
R1745 a_185_182.n2 a_185_182.n1 161.6
R1746 a_185_182.n3 a_185_182.n2 156.579
R1747 a_185_182.n5 a_185_182.n3 142.121
R1748 a_185_182.n5 a_185_182.n4 15.218
R1749 a_185_182.n0 a_185_182.t2 14.282
R1750 a_185_182.n0 a_185_182.t1 14.282
R1751 a_185_182.n6 a_185_182.n5 12.014
R1752 a_1222_74.t0 a_1222_74.n1 34.62
R1753 a_1222_74.t0 a_1222_74.n0 8.137
R1754 a_1222_74.t0 a_1222_74.n2 4.69
R1755 a_3442_74.n12 a_3442_74.n11 26.811
R1756 a_3442_74.n6 a_3442_74.n5 24.977
R1757 a_3442_74.n2 a_3442_74.n1 24.877
R1758 a_3442_74.t0 a_3442_74.n2 12.677
R1759 a_3442_74.t0 a_3442_74.n3 11.595
R1760 a_3442_74.t1 a_3442_74.n8 8.137
R1761 a_3442_74.t0 a_3442_74.n4 7.273
R1762 a_3442_74.t0 a_3442_74.n0 6.109
R1763 a_3442_74.t1 a_3442_74.n7 4.864
R1764 a_3442_74.t0 a_3442_74.n12 2.074
R1765 a_3442_74.n7 a_3442_74.n6 1.13
R1766 a_3442_74.n12 a_3442_74.t1 0.937
R1767 a_3442_74.t1 a_3442_74.n10 0.804
R1768 a_3442_74.n10 a_3442_74.n9 0.136
R1769 a_2405_182.n1 a_2405_182.t3 477.179
R1770 a_2405_182.n1 a_2405_182.t5 406.485
R1771 a_2405_182.n2 a_2405_182.t4 225.731
R1772 a_2405_182.n3 a_2405_182.n0 220.249
R1773 a_2405_182.n2 a_2405_182.n1 161.6
R1774 a_2405_182.n3 a_2405_182.n2 156.579
R1775 a_2405_182.n5 a_2405_182.n3 142.121
R1776 a_2405_182.n5 a_2405_182.n4 15.218
R1777 a_2405_182.n0 a_2405_182.t1 14.282
R1778 a_2405_182.n0 a_2405_182.t2 14.282
R1779 a_2405_182.n6 a_2405_182.n5 12.014
R1780 a_6858_181.n2 a_6858_181.t6 512.525
R1781 a_6858_181.n2 a_6858_181.t5 371.139
R1782 a_6858_181.n3 a_6858_181.t4 220.263
R1783 a_6858_181.n4 a_6858_181.n1 175.383
R1784 a_6858_181.n3 a_6858_181.n2 158.3
R1785 a_6858_181.n4 a_6858_181.n3 153.043
R1786 a_6858_181.n8 a_6858_181.n4 145.681
R1787 a_6858_181.n8 a_6858_181.n7 133.539
R1788 a_6858_181.n11 a_6858_181.n0 55.263
R1789 a_6858_181.n10 a_6858_181.n8 48.405
R1790 a_6858_181.n10 a_6858_181.n9 30
R1791 a_6858_181.n11 a_6858_181.n10 25.263
R1792 a_6858_181.n7 a_6858_181.n6 22.578
R1793 a_6858_181.n1 a_6858_181.t2 14.282
R1794 a_6858_181.n1 a_6858_181.t1 14.282
R1795 a_6858_181.n7 a_6858_181.n5 8.58
R1796 a_7511_182.n2 a_7511_182.n0 362.371
R1797 a_7511_182.n2 a_7511_182.n1 15.218
R1798 a_7511_182.n0 a_7511_182.t1 14.282
R1799 a_7511_182.n0 a_7511_182.t2 14.282
R1800 a_7511_182.n3 a_7511_182.n2 12.014
R1801 a_4552_73.n5 a_4552_73.n4 24.877
R1802 a_4552_73.t0 a_4552_73.n5 12.677
R1803 a_4552_73.t0 a_4552_73.n3 11.595
R1804 a_4552_73.t0 a_4552_73.n6 8.137
R1805 a_4552_73.n2 a_4552_73.n0 4.031
R1806 a_4552_73.n2 a_4552_73.n1 3.644
R1807 a_4552_73.t0 a_4552_73.n2 1.093
R1808 a_4657_1004.n4 a_4657_1004.t7 512.525
R1809 a_4657_1004.n4 a_4657_1004.t5 371.139
R1810 a_4657_1004.n5 a_4657_1004.t6 220.263
R1811 a_4657_1004.n8 a_4657_1004.n6 194.086
R1812 a_4657_1004.n6 a_4657_1004.n3 162.547
R1813 a_4657_1004.n5 a_4657_1004.n4 158.3
R1814 a_4657_1004.n6 a_4657_1004.n5 153.043
R1815 a_4657_1004.n3 a_4657_1004.n2 76.002
R1816 a_4657_1004.n9 a_4657_1004.n0 55.263
R1817 a_4657_1004.n8 a_4657_1004.n7 30
R1818 a_4657_1004.n9 a_4657_1004.n8 23.684
R1819 a_4657_1004.n1 a_4657_1004.t3 14.282
R1820 a_4657_1004.n1 a_4657_1004.t2 14.282
R1821 a_4657_1004.n2 a_4657_1004.t0 14.282
R1822 a_4657_1004.n2 a_4657_1004.t1 14.282
R1823 a_4657_1004.n3 a_4657_1004.n1 12.85
R1824 a_556_74.n12 a_556_74.n11 26.811
R1825 a_556_74.n6 a_556_74.n5 24.977
R1826 a_556_74.n2 a_556_74.n1 24.877
R1827 a_556_74.t0 a_556_74.n2 12.677
R1828 a_556_74.t0 a_556_74.n3 11.595
R1829 a_556_74.t1 a_556_74.n8 8.137
R1830 a_556_74.t0 a_556_74.n4 7.273
R1831 a_556_74.t0 a_556_74.n0 6.109
R1832 a_556_74.t1 a_556_74.n7 4.864
R1833 a_556_74.t0 a_556_74.n12 2.074
R1834 a_556_74.n7 a_556_74.n6 1.13
R1835 a_556_74.n12 a_556_74.t1 0.937
R1836 a_556_74.t1 a_556_74.n10 0.804
R1837 a_556_74.n10 a_556_74.n9 0.136
R1838 a_5662_73.t0 a_5662_73.n1 34.62
R1839 a_5662_73.t0 a_5662_73.n0 8.137
R1840 a_5662_73.t0 a_5662_73.n2 4.69
R1841 a_2776_74.t0 a_2776_74.n1 34.62
R1842 a_2776_74.t0 a_2776_74.n0 8.137
R1843 a_2776_74.t0 a_2776_74.n2 4.69
C10 VPB VNB 30.88fF
C11 a_2776_74.n0 VNB 0.05fF
C12 a_2776_74.n1 VNB 0.12fF
C13 a_2776_74.n2 VNB 0.04fF
C14 a_5662_73.n0 VNB 0.05fF
C15 a_5662_73.n1 VNB 0.12fF
C16 a_5662_73.n2 VNB 0.04fF
C17 a_556_74.n0 VNB 0.02fF
C18 a_556_74.n1 VNB 0.10fF
C19 a_556_74.n2 VNB 0.06fF
C20 a_556_74.n3 VNB 0.06fF
C21 a_556_74.n4 VNB 0.00fF
C22 a_556_74.n5 VNB 0.04fF
C23 a_556_74.n6 VNB 0.05fF
C24 a_556_74.n7 VNB 0.02fF
C25 a_556_74.n8 VNB 0.05fF
C26 a_556_74.n9 VNB 0.08fF
C27 a_556_74.n10 VNB 0.18fF
C28 a_556_74.t1 VNB 0.24fF
C29 a_556_74.n11 VNB 0.09fF
C30 a_556_74.n12 VNB 0.00fF
C31 a_4657_1004.n0 VNB 0.05fF
C32 a_4657_1004.n1 VNB 0.45fF
C33 a_4657_1004.n2 VNB 0.54fF
C34 a_4657_1004.n3 VNB 0.27fF
C35 a_4657_1004.n4 VNB 0.30fF
C36 a_4657_1004.t6 VNB 0.45fF
C37 a_4657_1004.n5 VNB 0.49fF
C38 a_4657_1004.n6 VNB 0.49fF
C39 a_4657_1004.n7 VNB 0.02fF
C40 a_4657_1004.n8 VNB 0.24fF
C41 a_4657_1004.n9 VNB 0.04fF
C42 a_4552_73.n0 VNB 0.08fF
C43 a_4552_73.n1 VNB 0.02fF
C44 a_4552_73.n2 VNB 0.01fF
C45 a_4552_73.n3 VNB 0.06fF
C46 a_4552_73.n4 VNB 0.10fF
C47 a_4552_73.n5 VNB 0.06fF
C48 a_4552_73.n6 VNB 0.05fF
C49 a_7511_182.n0 VNB 1.03fF
C50 a_7511_182.n1 VNB 0.09fF
C51 a_7511_182.n2 VNB 0.49fF
C52 a_7511_182.n3 VNB 0.05fF
C53 a_6858_181.n0 VNB 0.05fF
C54 a_6858_181.n1 VNB 0.57fF
C55 a_6858_181.n2 VNB 0.30fF
C56 a_6858_181.t4 VNB 0.43fF
C57 a_6858_181.n3 VNB 0.48fF
C58 a_6858_181.n4 VNB 0.44fF
C59 a_6858_181.n5 VNB 0.04fF
C60 a_6858_181.n6 VNB 0.05fF
C61 a_6858_181.n7 VNB 0.16fF
C62 a_6858_181.n8 VNB 0.34fF
C63 a_6858_181.n9 VNB 0.02fF
C64 a_6858_181.n10 VNB 0.08fF
C65 a_6858_181.n11 VNB 0.04fF
C66 a_2405_182.n0 VNB 1.40fF
C67 a_2405_182.n1 VNB 0.79fF
C68 a_2405_182.n2 VNB 1.62fF
C69 a_2405_182.n3 VNB 1.73fF
C70 a_2405_182.n4 VNB 0.15fF
C71 a_2405_182.n5 VNB 0.34fF
C72 a_2405_182.n6 VNB 0.08fF
C73 a_3442_74.n0 VNB 0.02fF
C74 a_3442_74.n1 VNB 0.10fF
C75 a_3442_74.n2 VNB 0.06fF
C76 a_3442_74.n3 VNB 0.06fF
C77 a_3442_74.n4 VNB 0.00fF
C78 a_3442_74.n5 VNB 0.04fF
C79 a_3442_74.n6 VNB 0.05fF
C80 a_3442_74.n7 VNB 0.02fF
C81 a_3442_74.n8 VNB 0.05fF
C82 a_3442_74.n9 VNB 0.08fF
C83 a_3442_74.n10 VNB 0.17fF
C84 a_3442_74.n11 VNB 0.09fF
C85 a_3442_74.n12 VNB 0.00fF
C86 a_1222_74.n0 VNB 0.05fF
C87 a_1222_74.n1 VNB 0.12fF
C88 a_1222_74.n2 VNB 0.04fF
C89 a_185_182.n0 VNB 1.07fF
C90 a_185_182.n1 VNB 0.60fF
C91 a_185_182.t3 VNB 0.63fF
C92 a_185_182.n2 VNB 1.24fF
C93 a_185_182.n3 VNB 1.32fF
C94 a_185_182.n4 VNB 0.11fF
C95 a_185_182.n5 VNB 0.26fF
C96 a_185_182.n6 VNB 0.06fF
C97 a_1241_1004.n0 VNB 0.52fF
C98 a_6401_182.n0 VNB 0.76fF
C99 a_6401_182.n1 VNB 0.36fF
C100 a_6401_182.t4 VNB 0.53fF
C101 a_6401_182.n2 VNB 0.63fF
C102 a_6401_182.n3 VNB 0.70fF
C103 a_6401_182.n4 VNB 0.09fF
C104 a_6401_182.n5 VNB 0.27fF
C105 a_6401_182.n6 VNB 0.05fF
C106 a_5767_1004.n0 VNB 0.04fF
C107 a_5767_1004.n1 VNB 0.48fF
C108 a_5767_1004.n2 VNB 0.57fF
C109 a_5767_1004.n3 VNB 0.29fF
C110 a_5767_1004.n4 VNB 0.32fF
C111 a_5767_1004.t5 VNB 0.47fF
C112 a_5767_1004.n5 VNB 0.52fF
C113 a_5767_1004.n6 VNB 0.51fF
C114 a_5767_1004.n7 VNB 0.03fF
C115 a_5767_1004.n8 VNB 0.25fF
C116 a_5767_1004.n9 VNB 0.05fF
C117 a_6791_1005.n0 VNB 0.55fF
C118 a_5291_182.n0 VNB 0.04fF
C119 a_5291_182.n1 VNB 0.84fF
C120 a_5291_182.n2 VNB 0.44fF
C121 a_5291_182.t5 VNB 0.54fF
C122 a_5291_182.n3 VNB 1.11fF
C123 a_5291_182.n4 VNB 1.16fF
C124 a_5291_182.n5 VNB 0.04fF
C125 a_5291_182.n6 VNB 0.26fF
C126 a_5291_182.n7 VNB 0.06fF
C127 a_2795_1004.n0 VNB 0.52fF
C128 a_575_1004.n0 VNB 0.52fF
C129 a_836_182.n0 VNB 0.06fF
C130 a_836_182.n1 VNB 1.04fF
C131 a_836_182.n2 VNB 0.46fF
C132 a_836_182.n3 VNB 0.52fF
C133 a_836_182.n4 VNB 1.01fF
C134 a_836_182.n5 VNB 0.64fF
C135 a_836_182.n6 VNB 0.71fF
C136 a_836_182.t10 VNB 0.70fF
C137 a_836_182.n7 VNB 2.22fF
C138 a_836_182.t13 VNB 0.70fF
C139 a_836_182.n8 VNB 2.06fF
C140 a_836_182.n9 VNB 0.26fF
C141 a_836_182.n10 VNB 1.04fF
C142 a_836_182.n11 VNB 0.65fF
C143 a_836_182.n12 VNB 0.75fF
C144 a_836_182.n13 VNB 1.91fF
C145 a_836_182.n14 VNB 0.71fF
C146 a_836_182.n15 VNB 0.05fF
C147 a_836_182.n16 VNB 0.50fF
C148 a_836_182.n17 VNB 0.09fF
C149 a_807_943.n0 VNB 0.07fF
C150 a_807_943.n1 VNB 1.19fF
C151 a_807_943.n2 VNB 1.29fF
C152 a_807_943.n3 VNB 1.42fF
C153 a_807_943.n4 VNB 1.61fF
C154 a_807_943.n5 VNB 0.06fF
C155 a_807_943.n6 VNB 0.48fF
C156 a_807_943.n7 VNB 0.10fF
C157 a_3027_943.n0 VNB 0.07fF
C158 a_3027_943.n1 VNB 1.23fF
C159 a_3027_943.n2 VNB 1.34fF
C160 a_3027_943.n3 VNB 1.48fF
C161 a_3027_943.n4 VNB 1.67fF
C162 a_3027_943.n5 VNB 0.06fF
C163 a_3027_943.n6 VNB 0.49fF
C164 a_3027_943.n7 VNB 0.10fF
C165 VPB.n0 VNB 0.03fF
C166 VPB.n1 VNB 0.04fF
C167 VPB.n2 VNB 0.02fF
C168 VPB.n3 VNB 0.11fF
C169 VPB.n5 VNB 0.02fF
C170 VPB.n6 VNB 0.02fF
C171 VPB.n7 VNB 0.02fF
C172 VPB.n8 VNB 0.02fF
C173 VPB.n10 VNB 0.02fF
C174 VPB.n11 VNB 0.02fF
C175 VPB.n12 VNB 0.02fF
C176 VPB.n14 VNB 0.02fF
C177 VPB.n15 VNB 0.02fF
C178 VPB.n16 VNB 0.02fF
C179 VPB.n17 VNB 0.04fF
C180 VPB.n18 VNB 0.02fF
C181 VPB.n19 VNB 0.17fF
C182 VPB.n20 VNB 0.04fF
C183 VPB.n22 VNB 0.02fF
C184 VPB.n23 VNB 0.02fF
C185 VPB.n24 VNB 0.02fF
C186 VPB.n25 VNB 0.02fF
C187 VPB.n27 VNB 0.02fF
C188 VPB.n28 VNB 0.02fF
C189 VPB.n29 VNB 0.02fF
C190 VPB.n31 VNB 0.27fF
C191 VPB.n33 VNB 0.03fF
C192 VPB.n34 VNB 0.02fF
C193 VPB.n35 VNB 0.09fF
C194 VPB.n36 VNB 0.27fF
C195 VPB.n37 VNB 0.02fF
C196 VPB.n38 VNB 0.02fF
C197 VPB.n39 VNB 0.27fF
C198 VPB.n40 VNB 0.02fF
C199 VPB.n41 VNB 0.02fF
C200 VPB.n42 VNB 0.14fF
C201 VPB.n43 VNB 0.15fF
C202 VPB.n44 VNB 0.02fF
C203 VPB.n45 VNB 0.02fF
C204 VPB.n46 VNB 0.03fF
C205 VPB.n47 VNB 0.14fF
C206 VPB.n48 VNB 0.16fF
C207 VPB.n49 VNB 0.02fF
C208 VPB.n50 VNB 0.02fF
C209 VPB.n51 VNB 0.23fF
C210 VPB.n52 VNB 0.02fF
C211 VPB.n53 VNB 0.02fF
C212 VPB.n54 VNB 0.27fF
C213 VPB.n55 VNB 0.01fF
C214 VPB.n56 VNB 0.02fF
C215 VPB.n57 VNB 0.03fF
C216 VPB.n58 VNB 0.03fF
C217 VPB.n59 VNB 0.27fF
C218 VPB.n60 VNB 0.01fF
C219 VPB.n61 VNB 0.02fF
C220 VPB.n62 VNB 0.06fF
C221 VPB.n63 VNB 0.14fF
C222 VPB.n64 VNB 0.19fF
C223 VPB.n65 VNB 0.02fF
C224 VPB.n66 VNB 0.01fF
C225 VPB.n67 VNB 0.16fF
C226 VPB.n68 VNB 0.02fF
C227 VPB.n69 VNB 0.02fF
C228 VPB.n70 VNB 0.14fF
C229 VPB.n71 VNB 0.19fF
C230 VPB.n72 VNB 0.02fF
C231 VPB.n73 VNB 0.01fF
C232 VPB.n74 VNB 0.06fF
C233 VPB.n75 VNB 0.02fF
C234 VPB.n76 VNB 0.02fF
C235 VPB.n77 VNB 0.02fF
C236 VPB.n78 VNB 0.04fF
C237 VPB.n79 VNB 0.02fF
C238 VPB.n80 VNB 0.16fF
C239 VPB.n81 VNB 0.04fF
C240 VPB.n83 VNB 0.02fF
C241 VPB.n84 VNB 0.02fF
C242 VPB.n85 VNB 0.02fF
C243 VPB.n86 VNB 0.02fF
C244 VPB.n88 VNB 0.02fF
C245 VPB.n89 VNB 0.02fF
C246 VPB.n90 VNB 0.02fF
C247 VPB.n92 VNB 0.27fF
C248 VPB.n94 VNB 0.03fF
C249 VPB.n95 VNB 0.02fF
C250 VPB.n96 VNB 0.02fF
C251 VPB.n97 VNB 0.02fF
C252 VPB.n98 VNB 0.02fF
C253 VPB.n99 VNB 0.04fF
C254 VPB.n100 VNB 0.02fF
C255 VPB.n101 VNB 0.16fF
C256 VPB.n102 VNB 0.04fF
C257 VPB.n104 VNB 0.02fF
C258 VPB.n105 VNB 0.02fF
C259 VPB.n106 VNB 0.02fF
C260 VPB.n107 VNB 0.02fF
C261 VPB.n109 VNB 0.02fF
C262 VPB.n110 VNB 0.02fF
C263 VPB.n111 VNB 0.02fF
C264 VPB.n113 VNB 0.27fF
C265 VPB.n115 VNB 0.03fF
C266 VPB.n116 VNB 0.02fF
C267 VPB.n117 VNB 0.10fF
C268 VPB.n118 VNB 0.02fF
C269 VPB.n119 VNB 0.14fF
C270 VPB.n120 VNB 0.15fF
C271 VPB.n121 VNB 0.02fF
C272 VPB.n122 VNB 0.02fF
C273 VPB.n123 VNB 0.14fF
C274 VPB.n124 VNB 0.16fF
C275 VPB.n125 VNB 0.02fF
C276 VPB.n126 VNB 0.02fF
C277 VPB.n127 VNB 0.06fF
C278 VPB.n128 VNB 0.23fF
C279 VPB.n129 VNB 0.02fF
C280 VPB.n130 VNB 0.01fF
C281 VPB.n131 VNB 0.27fF
C282 VPB.n132 VNB 0.01fF
C283 VPB.n133 VNB 0.02fF
C284 VPB.n134 VNB 0.03fF
C285 VPB.n135 VNB 0.03fF
C286 VPB.n136 VNB 0.27fF
C287 VPB.n137 VNB 0.01fF
C288 VPB.n138 VNB 0.02fF
C289 VPB.n139 VNB 0.06fF
C290 VPB.n140 VNB 0.14fF
C291 VPB.n141 VNB 0.19fF
C292 VPB.n142 VNB 0.02fF
C293 VPB.n143 VNB 0.01fF
C294 VPB.n144 VNB 0.16fF
C295 VPB.n145 VNB 0.02fF
C296 VPB.n146 VNB 0.02fF
C297 VPB.n147 VNB 0.14fF
C298 VPB.n148 VNB 0.19fF
C299 VPB.n149 VNB 0.02fF
C300 VPB.n150 VNB 0.01fF
C301 VPB.n151 VNB 0.06fF
C302 VPB.n152 VNB 0.27fF
C303 VPB.n153 VNB 0.01fF
C304 VPB.n154 VNB 0.02fF
C305 VPB.n155 VNB 0.03fF
C306 VPB.n156 VNB 0.02fF
C307 VPB.n157 VNB 0.02fF
C308 VPB.n158 VNB 0.02fF
C309 VPB.n159 VNB 0.11fF
C310 VPB.n160 VNB 0.03fF
C311 VPB.n161 VNB 0.02fF
C312 VPB.n162 VNB 0.05fF
C313 VPB.n163 VNB 0.01fF
C314 VPB.n164 VNB 0.02fF
C315 VPB.n165 VNB 0.02fF
C316 VPB.n168 VNB 0.02fF
C317 VPB.n169 VNB 0.02fF
C318 VPB.n171 VNB 0.02fF
C319 VPB.n173 VNB 0.46fF
C320 VPB.n175 VNB 0.04fF
C321 VPB.n176 VNB 0.04fF
C322 VPB.n177 VNB 0.27fF
C323 VPB.n178 VNB 0.03fF
C324 VPB.n179 VNB 0.03fF
C325 VPB.n180 VNB 0.06fF
C326 VPB.n181 VNB 0.14fF
C327 VPB.n182 VNB 0.19fF
C328 VPB.n183 VNB 0.02fF
C329 VPB.n184 VNB 0.01fF
C330 VPB.n185 VNB 0.07fF
C331 VPB.n186 VNB 0.16fF
C332 VPB.n187 VNB 0.02fF
C333 VPB.n188 VNB 0.02fF
C334 VPB.n189 VNB 0.02fF
C335 VPB.n190 VNB 0.06fF
C336 VPB.n191 VNB 0.14fF
C337 VPB.n192 VNB 0.19fF
C338 VPB.n193 VNB 0.02fF
C339 VPB.n194 VNB 0.01fF
C340 VPB.n195 VNB 0.02fF
C341 VPB.n196 VNB 0.27fF
C342 VPB.n197 VNB 0.01fF
C343 VPB.n198 VNB 0.02fF
C344 VPB.n199 VNB 0.04fF
C345 VPB.n200 VNB 0.02fF
C346 VPB.n201 VNB 0.02fF
C347 VPB.n202 VNB 0.02fF
C348 VPB.n203 VNB 0.04fF
C349 VPB.n204 VNB 0.02fF
C350 VPB.n205 VNB 0.17fF
C351 VPB.n206 VNB 0.04fF
C352 VPB.n208 VNB 0.02fF
C353 VPB.n209 VNB 0.02fF
C354 VPB.n210 VNB 0.02fF
C355 VPB.n211 VNB 0.02fF
C356 VPB.n213 VNB 0.02fF
C357 VPB.n214 VNB 0.02fF
C358 VPB.n215 VNB 0.02fF
C359 VPB.n217 VNB 0.27fF
C360 VPB.n219 VNB 0.03fF
C361 VPB.n220 VNB 0.02fF
C362 VPB.n221 VNB 0.03fF
C363 VPB.n222 VNB 0.03fF
C364 VPB.n223 VNB 0.27fF
C365 VPB.n224 VNB 0.01fF
C366 VPB.n225 VNB 0.02fF
C367 VPB.n226 VNB 0.04fF
C368 VPB.n227 VNB 0.27fF
C369 VPB.n228 VNB 0.02fF
C370 VPB.n229 VNB 0.02fF
C371 VPB.n230 VNB 0.02fF
C372 VPB.n231 VNB 0.27fF
C373 VPB.n232 VNB 0.02fF
C374 VPB.n233 VNB 0.02fF
C375 VPB.n234 VNB 0.02fF
C376 VPB.n235 VNB 0.27fF
C377 VPB.n236 VNB 0.02fF
C378 VPB.n237 VNB 0.02fF
C379 VPB.n238 VNB 0.02fF
C380 VPB.n239 VNB 0.14fF
C381 VPB.n240 VNB 0.15fF
C382 VPB.n241 VNB 0.02fF
C383 VPB.n242 VNB 0.02fF
C384 VPB.n243 VNB 0.02fF
C385 VPB.n244 VNB 0.10fF
C386 VPB.n245 VNB 0.02fF
C387 VPB.n246 VNB 0.14fF
C388 VPB.n247 VNB 0.16fF
C389 VPB.n248 VNB 0.02fF
C390 VPB.n249 VNB 0.02fF
C391 VPB.n250 VNB 0.02fF
C392 VPB.n251 VNB 0.23fF
C393 VPB.n252 VNB 0.02fF
C394 VPB.n253 VNB 0.02fF
C395 VPB.n254 VNB 0.02fF
C396 VPB.n255 VNB 0.27fF
C397 VPB.n256 VNB 0.01fF
C398 VPB.n257 VNB 0.02fF
C399 VPB.n258 VNB 0.04fF
C400 VPB.n259 VNB 0.02fF
C401 VPB.n260 VNB 0.02fF
C402 VPB.n261 VNB 0.02fF
C403 VPB.n262 VNB 0.04fF
C404 VPB.n263 VNB 0.02fF
C405 VPB.n264 VNB 0.16fF
C406 VPB.n265 VNB 0.04fF
C407 VPB.n267 VNB 0.02fF
C408 VPB.n268 VNB 0.02fF
C409 VPB.n269 VNB 0.02fF
C410 VPB.n270 VNB 0.02fF
C411 VPB.n272 VNB 0.02fF
C412 VPB.n273 VNB 0.02fF
C413 VPB.n274 VNB 0.02fF
C414 VPB.n276 VNB 0.27fF
C415 VPB.n278 VNB 0.03fF
C416 VPB.n279 VNB 0.02fF
C417 VPB.n280 VNB 0.03fF
C418 VPB.n281 VNB 0.03fF
C419 VPB.n282 VNB 0.27fF
C420 VPB.n283 VNB 0.01fF
C421 VPB.n284 VNB 0.02fF
C422 VPB.n285 VNB 0.04fF
C423 VPB.n286 VNB 0.06fF
C424 VPB.n287 VNB 0.14fF
C425 VPB.n288 VNB 0.19fF
C426 VPB.n289 VNB 0.02fF
C427 VPB.n290 VNB 0.01fF
C428 VPB.n291 VNB 0.02fF
C429 VPB.n292 VNB 0.16fF
C430 VPB.n293 VNB 0.02fF
C431 VPB.n294 VNB 0.02fF
C432 VPB.n295 VNB 0.02fF
C433 VPB.n296 VNB 0.06fF
C434 VPB.n297 VNB 0.14fF
C435 VPB.n298 VNB 0.19fF
C436 VPB.n299 VNB 0.02fF
C437 VPB.n300 VNB 0.01fF
C438 VPB.n301 VNB 0.02fF
C439 VPB.n302 VNB 0.27fF
C440 VPB.n303 VNB 0.01fF
C441 VPB.n304 VNB 0.02fF
C442 VPB.n305 VNB 0.04fF
C443 VPB.n306 VNB 0.02fF
C444 VPB.n307 VNB 0.02fF
C445 VPB.n308 VNB 0.02fF
C446 VPB.n309 VNB 0.04fF
C447 VPB.n310 VNB 0.02fF
C448 VPB.n311 VNB 0.16fF
C449 VPB.n312 VNB 0.04fF
C450 VPB.n314 VNB 0.02fF
C451 VPB.n315 VNB 0.02fF
C452 VPB.n316 VNB 0.02fF
C453 VPB.n317 VNB 0.02fF
C454 VPB.n319 VNB 0.02fF
C455 VPB.n320 VNB 0.02fF
C456 VPB.n321 VNB 0.02fF
C457 VPB.n323 VNB 0.27fF
C458 VPB.n325 VNB 0.03fF
C459 VPB.n326 VNB 0.02fF
C460 VPB.n327 VNB 0.03fF
C461 VPB.n328 VNB 0.03fF
C462 VPB.n329 VNB 0.27fF
C463 VPB.n330 VNB 0.01fF
C464 VPB.n331 VNB 0.02fF
C465 VPB.n332 VNB 0.04fF
C466 VPB.n333 VNB 0.05fF
C467 VPB.n334 VNB 0.23fF
C468 VPB.n335 VNB 0.02fF
C469 VPB.n336 VNB 0.01fF
C470 VPB.n337 VNB 0.02fF
C471 VPB.n338 VNB 0.14fF
C472 VPB.n339 VNB 0.16fF
C473 VPB.n340 VNB 0.02fF
C474 VPB.n341 VNB 0.02fF
C475 VPB.n342 VNB 0.02fF
C476 VPB.n343 VNB 0.10fF
C477 VPB.n344 VNB 0.02fF
C478 VPB.n345 VNB 0.14fF
C479 VPB.n346 VNB 0.15fF
C480 VPB.n347 VNB 0.02fF
C481 VPB.n348 VNB 0.02fF
C482 VPB.n349 VNB 0.02fF
C483 VPB.n350 VNB 0.14fF
C484 VPB.n351 VNB 0.15fF
C485 VPB.n352 VNB 0.02fF
C486 VPB.n353 VNB 0.02fF
C487 VPB.n354 VNB 0.02fF
C488 VPB.n355 VNB 0.14fF
C489 VPB.n356 VNB 0.16fF
C490 VPB.n357 VNB 0.02fF
C491 VPB.n358 VNB 0.02fF
C492 VPB.n359 VNB 0.02fF
C493 VPB.n360 VNB 0.06fF
C494 VPB.n361 VNB 0.23fF
C495 VPB.n362 VNB 0.02fF
C496 VPB.n363 VNB 0.01fF
C497 VPB.n364 VNB 0.02fF
C498 VPB.n365 VNB 0.27fF
C499 VPB.n366 VNB 0.01fF
C500 VPB.n367 VNB 0.02fF
C501 VPB.n368 VNB 0.04fF
C502 VPB.n369 VNB 0.02fF
C503 VPB.n370 VNB 0.02fF
C504 VPB.n371 VNB 0.02fF
C505 VPB.n372 VNB 0.04fF
C506 VPB.n373 VNB 0.02fF
C507 VPB.n374 VNB 0.16fF
C508 VPB.n375 VNB 0.04fF
C509 VPB.n377 VNB 0.02fF
C510 VPB.n378 VNB 0.02fF
C511 VPB.n379 VNB 0.02fF
C512 VPB.n380 VNB 0.02fF
C513 VPB.n382 VNB 0.02fF
C514 VPB.n383 VNB 0.02fF
C515 VPB.n384 VNB 0.02fF
C516 VPB.n386 VNB 0.27fF
C517 VPB.n388 VNB 0.03fF
C518 VPB.n389 VNB 0.02fF
C519 VPB.n390 VNB 0.03fF
C520 VPB.n391 VNB 0.03fF
C521 VPB.n392 VNB 0.27fF
C522 VPB.n393 VNB 0.01fF
C523 VPB.n394 VNB 0.02fF
C524 VPB.n395 VNB 0.04fF
C525 VPB.n396 VNB 0.06fF
C526 VPB.n397 VNB 0.14fF
C527 VPB.n398 VNB 0.19fF
C528 VPB.n399 VNB 0.02fF
C529 VPB.n400 VNB 0.01fF
C530 VPB.n401 VNB 0.02fF
C531 VPB.n402 VNB 0.16fF
C532 VPB.n403 VNB 0.02fF
C533 VPB.n404 VNB 0.02fF
C534 VPB.n405 VNB 0.02fF
C535 VPB.n406 VNB 0.06fF
C536 VPB.n407 VNB 0.14fF
C537 VPB.n408 VNB 0.19fF
C538 VPB.n409 VNB 0.02fF
C539 VPB.n410 VNB 0.01fF
C540 VPB.n411 VNB 0.02fF
C541 VPB.n412 VNB 0.27fF
C542 VPB.n413 VNB 0.01fF
C543 VPB.n414 VNB 0.02fF
C544 VPB.n415 VNB 0.04fF
C545 VPB.n416 VNB 0.02fF
C546 VPB.n417 VNB 0.02fF
C547 VPB.n418 VNB 0.02fF
C548 VPB.n419 VNB 0.04fF
C549 VPB.n420 VNB 0.02fF
C550 VPB.n421 VNB 0.16fF
C551 VPB.n422 VNB 0.04fF
C552 VPB.n424 VNB 0.02fF
C553 VPB.n425 VNB 0.02fF
C554 VPB.n426 VNB 0.02fF
C555 VPB.n427 VNB 0.02fF
C556 VPB.n429 VNB 0.02fF
C557 VPB.n430 VNB 0.02fF
C558 VPB.n431 VNB 0.02fF
C559 VPB.n433 VNB 0.27fF
C560 VPB.n435 VNB 0.03fF
C561 VPB.n436 VNB 0.02fF
C562 VPB.n437 VNB 0.03fF
C563 VPB.n438 VNB 0.03fF
C564 VPB.n439 VNB 0.27fF
C565 VPB.n440 VNB 0.01fF
C566 VPB.n441 VNB 0.02fF
C567 VPB.n442 VNB 0.04fF
C568 VPB.n443 VNB 0.05fF
C569 VPB.n444 VNB 0.23fF
C570 VPB.n445 VNB 0.02fF
C571 VPB.n446 VNB 0.01fF
C572 VPB.n447 VNB 0.02fF
C573 VPB.n448 VNB 0.14fF
C574 VPB.n449 VNB 0.16fF
C575 VPB.n450 VNB 0.02fF
C576 VPB.n451 VNB 0.02fF
C577 VPB.n452 VNB 0.02fF
C578 VPB.n453 VNB 0.14fF
C579 VPB.n454 VNB 0.15fF
C580 VPB.n455 VNB 0.02fF
C581 VPB.n456 VNB 0.02fF
C582 VPB.n457 VNB 0.02fF
C583 VPB.n458 VNB 0.02fF
C584 VPB.n459 VNB 0.02fF
C585 VPB.n460 VNB 0.02fF
C586 VPB.n461 VNB 0.04fF
C587 VPB.n462 VNB 0.04fF
C588 VPB.n463 VNB 0.02fF
C589 VPB.n464 VNB 0.02fF
C590 VPB.n465 VNB 0.02fF
C591 VPB.n466 VNB 0.04fF
C592 VPB.n467 VNB 0.03fF
C593 VPB.n468 VNB 0.03fF
C594 VPB.n469 VNB 0.27fF
C595 VPB.n470 VNB 0.01fF
C596 VPB.n471 VNB 0.02fF
C597 VPB.n472 VNB 0.27fF
C598 VPB.n473 VNB 0.02fF
C599 VPB.n474 VNB 0.02fF
C600 VPB.n475 VNB 0.02fF
C601 VPB.n476 VNB 0.27fF
C602 VPB.n477 VNB 0.02fF
C603 VPB.n478 VNB 0.02fF
C604 VPB.n479 VNB 0.02fF
C605 VPB.n480 VNB 0.27fF
C606 VPB.n481 VNB 0.02fF
C607 VPB.n482 VNB 0.02fF
C608 VPB.n483 VNB 0.02fF
C609 VPB.n484 VNB 0.14fF
C610 VPB.n485 VNB 0.15fF
C611 VPB.n486 VNB 0.02fF
C612 VPB.n487 VNB 0.02fF
C613 VPB.n488 VNB 0.02fF
C614 VPB.n489 VNB 0.09fF
C615 VPB.n490 VNB 0.03fF
C616 VPB.n491 VNB 0.14fF
C617 VPB.n492 VNB 0.16fF
C618 VPB.n493 VNB 0.02fF
C619 VPB.n494 VNB 0.02fF
C620 VPB.n495 VNB 0.02fF
C621 VPB.n496 VNB 0.23fF
C622 VPB.n497 VNB 0.02fF
C623 VPB.n498 VNB 0.02fF
C624 VPB.n499 VNB 0.02fF
C625 VPB.n500 VNB 0.27fF
C626 VPB.n501 VNB 0.01fF
C627 VPB.n502 VNB 0.02fF
C628 VPB.n503 VNB 0.04fF
C629 VPB.n504 VNB 0.02fF
C630 VPB.n505 VNB 0.02fF
C631 VPB.n506 VNB 0.02fF
C632 VPB.n507 VNB 0.04fF
C633 VPB.n508 VNB 0.02fF
C634 VPB.n509 VNB 0.19fF
C635 VPB.n510 VNB 0.04fF
C636 VPB.n512 VNB 0.02fF
C637 VPB.n513 VNB 0.02fF
C638 VPB.n514 VNB 0.02fF
C639 VPB.n515 VNB 0.02fF
C640 VPB.n517 VNB 0.02fF
C641 VPB.n518 VNB 0.02fF
C642 VPB.n519 VNB 0.02fF
C643 VPB.n521 VNB 0.27fF
C644 VPB.n523 VNB 0.03fF
C645 VPB.n524 VNB 0.02fF
C646 VPB.n525 VNB 0.03fF
C647 VPB.n526 VNB 0.03fF
C648 VPB.n527 VNB 0.27fF
C649 VPB.n528 VNB 0.01fF
C650 VPB.n529 VNB 0.02fF
C651 VPB.n530 VNB 0.04fF
C652 VPB.n531 VNB 0.27fF
C653 VPB.n532 VNB 0.02fF
C654 VPB.n533 VNB 0.02fF
C655 VPB.n534 VNB 0.02fF
C656 VPB.n535 VNB 0.27fF
C657 VPB.n536 VNB 0.02fF
C658 VPB.n537 VNB 0.02fF
C659 VPB.n538 VNB 0.02fF
C660 VPB.n539 VNB 0.27fF
C661 VPB.n540 VNB 0.02fF
C662 VPB.n541 VNB 0.02fF
C663 VPB.n542 VNB 0.02fF
C664 VPB.n543 VNB 0.14fF
C665 VPB.n544 VNB 0.15fF
C666 VPB.n545 VNB 0.02fF
C667 VPB.n546 VNB 0.02fF
C668 VPB.n547 VNB 0.02fF
C669 VPB.n548 VNB 0.09fF
C670 VPB.n549 VNB 0.03fF
C671 VPB.n550 VNB 0.14fF
C672 VPB.n551 VNB 0.16fF
C673 VPB.n552 VNB 0.02fF
C674 VPB.n553 VNB 0.02fF
C675 VPB.n554 VNB 0.02fF
C676 VPB.n555 VNB 0.23fF
C677 VPB.n556 VNB 0.02fF
C678 VPB.n557 VNB 0.02fF
C679 VPB.n558 VNB 0.02fF
C680 VPB.n559 VNB 0.27fF
C681 VPB.n560 VNB 0.01fF
C682 VPB.n561 VNB 0.02fF
C683 VPB.n562 VNB 0.04fF
C684 VPB.n563 VNB 0.02fF
C685 VPB.n564 VNB 0.02fF
C686 VPB.n565 VNB 0.02fF
C687 VPB.n566 VNB 0.04fF
C688 VPB.n567 VNB 0.02fF
C689 VPB.n568 VNB 0.16fF
C690 VPB.n569 VNB 0.04fF
C691 VPB.n571 VNB 0.02fF
C692 VPB.n572 VNB 0.02fF
C693 VPB.n573 VNB 0.02fF
C694 VPB.n574 VNB 0.02fF
C695 VPB.n576 VNB 0.02fF
C696 VPB.n577 VNB 0.02fF
C697 VPB.n578 VNB 0.02fF
C698 VPB.n580 VNB 0.27fF
C699 VPB.n582 VNB 0.03fF
C700 VPB.n583 VNB 0.02fF
C701 VPB.n584 VNB 0.03fF
C702 VPB.n585 VNB 0.03fF
C703 VPB.n586 VNB 0.27fF
C704 VPB.n587 VNB 0.01fF
C705 VPB.n588 VNB 0.02fF
C706 VPB.n589 VNB 0.04fF
C707 VPB.n590 VNB 0.06fF
C708 VPB.n591 VNB 0.14fF
C709 VPB.n592 VNB 0.19fF
C710 VPB.n593 VNB 0.02fF
C711 VPB.n594 VNB 0.01fF
C712 VPB.n595 VNB 0.02fF
C713 VPB.n596 VNB 0.16fF
C714 VPB.n597 VNB 0.02fF
C715 VPB.n598 VNB 0.02fF
C716 VPB.n599 VNB 0.02fF
C717 VPB.n600 VNB 0.06fF
C718 VPB.n601 VNB 0.14fF
C719 VPB.n602 VNB 0.19fF
C720 VPB.n603 VNB 0.02fF
C721 VPB.n604 VNB 0.01fF
C722 VPB.n605 VNB 0.02fF
C723 VPB.n606 VNB 0.27fF
C724 VPB.n607 VNB 0.01fF
C725 VPB.n608 VNB 0.02fF
C726 VPB.n609 VNB 0.04fF
C727 VPB.n610 VNB 0.02fF
C728 VPB.n611 VNB 0.02fF
C729 VPB.n612 VNB 0.02fF
C730 VPB.n613 VNB 0.04fF
C731 VPB.n614 VNB 0.02fF
C732 VPB.n615 VNB 0.13fF
C733 VPB.n616 VNB 0.04fF
C734 VPB.n618 VNB 0.02fF
C735 VPB.n619 VNB 0.02fF
C736 VPB.n620 VNB 0.02fF
C737 VPB.n621 VNB 0.02fF
C738 VPB.n623 VNB 0.02fF
C739 VPB.n624 VNB 0.02fF
C740 VPB.n625 VNB 0.02fF
C741 VPB.n627 VNB 0.27fF
C742 VPB.n629 VNB 0.03fF
C743 VPB.n630 VNB 0.02fF
C744 VPB.n631 VNB 0.03fF
C745 VPB.n632 VNB 0.03fF
C746 VPB.n633 VNB 0.27fF
C747 VPB.n634 VNB 0.01fF
C748 VPB.n635 VNB 0.02fF
C749 VPB.n636 VNB 0.04fF
C750 VPB.n637 VNB 0.06fF
C751 VPB.n638 VNB 0.14fF
C752 VPB.n639 VNB 0.19fF
C753 VPB.n640 VNB 0.02fF
C754 VPB.n641 VNB 0.01fF
C755 VPB.n642 VNB 0.02fF
C756 VPB.n643 VNB 0.16fF
C757 VPB.n644 VNB 0.02fF
C758 VPB.n645 VNB 0.02fF
C759 VPB.n646 VNB 0.02fF
C760 VPB.n647 VNB 0.06fF
C761 VPB.n648 VNB 0.14fF
C762 VPB.n649 VNB 0.19fF
C763 VPB.n650 VNB 0.02fF
C764 VPB.n651 VNB 0.01fF
C765 VPB.n652 VNB 0.02fF
C766 VPB.n653 VNB 0.27fF
C767 VPB.n654 VNB 0.01fF
C768 VPB.n655 VNB 0.02fF
C769 VPB.n656 VNB 0.04fF
C770 VPB.n657 VNB 0.02fF
C771 VPB.n658 VNB 0.02fF
C772 VPB.n659 VNB 0.02fF
C773 VPB.n660 VNB 0.04fF
C774 VPB.n661 VNB 0.02fF
C775 VPB.n662 VNB 0.16fF
C776 VPB.n663 VNB 0.04fF
C777 VPB.n665 VNB 0.02fF
C778 VPB.n666 VNB 0.02fF
C779 VPB.n667 VNB 0.02fF
C780 VPB.n668 VNB 0.02fF
C781 VPB.n670 VNB 0.02fF
C782 VPB.n671 VNB 0.02fF
C783 VPB.n672 VNB 0.02fF
C784 VPB.n674 VNB 0.27fF
C785 VPB.n676 VNB 0.03fF
C786 VPB.n677 VNB 0.02fF
C787 VPB.n678 VNB 0.03fF
C788 VPB.n679 VNB 0.03fF
C789 VPB.n680 VNB 0.27fF
C790 VPB.n681 VNB 0.01fF
C791 VPB.n682 VNB 0.02fF
C792 VPB.n683 VNB 0.04fF
C793 VPB.n684 VNB 0.27fF
C794 VPB.n685 VNB 0.02fF
C795 VPB.n686 VNB 0.02fF
C796 VPB.n687 VNB 0.02fF
C797 VPB.n688 VNB 0.27fF
C798 VPB.n689 VNB 0.02fF
C799 VPB.n690 VNB 0.02fF
C800 VPB.n691 VNB 0.02fF
C801 VPB.n692 VNB 0.27fF
C802 VPB.n693 VNB 0.02fF
C803 VPB.n694 VNB 0.02fF
C804 VPB.n695 VNB 0.02fF
C805 VPB.n696 VNB 0.14fF
C806 VPB.n697 VNB 0.15fF
C807 VPB.n698 VNB 0.02fF
C808 VPB.n699 VNB 0.02fF
C809 VPB.n700 VNB 0.02fF
C810 VPB.n701 VNB 0.09fF
C811 VPB.n702 VNB 0.03fF
C812 VPB.n703 VNB 0.14fF
C813 VPB.n704 VNB 0.16fF
C814 VPB.n705 VNB 0.02fF
C815 VPB.n706 VNB 0.02fF
C816 VPB.n707 VNB 0.02fF
C817 VPB.n708 VNB 0.23fF
C818 VPB.n709 VNB 0.02fF
C819 VPB.n710 VNB 0.02fF
C820 VPB.n711 VNB 0.02fF
C821 VPB.n712 VNB 0.27fF
C822 VPB.n713 VNB 0.01fF
C823 VPB.n714 VNB 0.02fF
C824 VPB.n715 VNB 0.04fF
C825 VPB.n716 VNB 0.02fF
C826 VPB.n717 VNB 0.02fF
C827 VPB.n718 VNB 0.02fF
C828 VPB.n719 VNB 0.04fF
C829 VPB.n720 VNB 0.02fF
C830 VPB.n721 VNB 0.19fF
C831 VPB.n722 VNB 0.04fF
C832 VPB.n724 VNB 0.02fF
C833 VPB.n725 VNB 0.02fF
C834 VPB.n726 VNB 0.02fF
C835 VPB.n727 VNB 0.02fF
C836 VPB.n729 VNB 0.02fF
C837 VPB.n730 VNB 0.02fF
C838 VPB.n731 VNB 0.02fF
C839 VPB.n733 VNB 0.27fF
C840 VPB.n735 VNB 0.03fF
C841 VPB.n736 VNB 0.02fF
C842 VPB.n737 VNB 0.03fF
C843 VPB.n738 VNB 0.03fF
C844 VPB.n739 VNB 0.27fF
C845 VPB.n740 VNB 0.01fF
C846 VPB.n741 VNB 0.02fF
C847 VPB.n742 VNB 0.04fF
C848 VPB.n743 VNB 0.27fF
C849 VPB.n744 VNB 0.02fF
C850 VPB.n745 VNB 0.02fF
C851 VPB.n746 VNB 0.02fF
C852 VPB.n747 VNB 0.02fF
C853 VPB.n748 VNB 0.02fF
C854 VPB.n749 VNB 0.02fF
C855 VPB.n750 VNB 0.02fF
C856 VPB.n751 VNB 0.02fF
C857 VPB.n752 VNB 0.04fF
C858 VPB.n753 VNB 0.04fF
C859 VPB.n754 VNB 0.02fF
C860 VPB.n755 VNB 0.02fF
C861 VPB.n756 VNB 0.02fF
C862 VPB.n757 VNB 0.03fF
C863 VPB.n758 VNB 0.03fF
C864 VPB.n759 VNB 0.02fF
C865 VPB.n760 VNB 0.02fF
C866 VPB.n761 VNB 0.02fF
C867 VPB.n762 VNB 0.04fF
C868 VPB.n763 VNB 0.04fF
C869 VPB.n765 VNB 0.42fF
C870 a_3461_1004.n0 VNB 0.52fF
.ends
