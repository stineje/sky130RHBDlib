magic
tech sky130A
magscale 1 2
timestamp 1651256905
<< nmos >>
tri 146 223 162 239 se
rect 162 223 192 276
tri 56 193 86 223 se
rect 86 193 192 223
rect 56 178 87 193
tri 87 178 102 193 nw
tri 146 178 161 193 ne
rect 161 178 192 193
rect 56 92 86 178
tri 86 92 102 108 sw
tri 146 92 162 108 se
rect 162 92 192 178
tri 56 62 86 92 ne
rect 86 62 162 92
tri 162 62 192 92 nw
<< ndiff >>
rect 0 239 162 276
rect 0 223 146 239
tri 146 223 162 239 nw
rect 0 188 56 223
tri 56 193 86 223 nw
rect 0 154 10 188
rect 44 154 56 188
tri 87 178 102 193 se
rect 102 178 146 193
tri 146 178 161 193 sw
rect 192 188 248 276
rect 0 120 56 154
rect 0 86 10 120
rect 44 86 56 120
rect 86 144 162 178
rect 86 110 107 144
rect 141 110 162 144
rect 86 108 162 110
tri 86 92 102 108 ne
rect 102 92 146 108
tri 146 92 162 108 nw
rect 192 154 204 188
rect 238 154 248 188
rect 192 120 248 154
rect 0 62 56 86
tri 56 62 86 92 sw
tri 162 62 192 92 se
rect 192 86 204 120
rect 238 86 248 120
rect 192 62 248 86
rect 0 50 248 62
rect 0 16 10 50
rect 44 16 107 50
rect 141 16 204 50
rect 238 16 248 50
rect 0 0 248 16
<< ndiffc >>
rect 10 154 44 188
rect 10 86 44 120
rect 107 110 141 144
rect 204 154 238 188
rect 204 86 238 120
rect 10 16 44 50
rect 107 16 141 50
rect 204 16 238 50
<< poly >>
rect 162 276 192 309
<< locali >>
rect 10 188 44 205
rect 204 188 238 205
rect 10 120 44 154
rect 107 144 141 161
rect 107 94 141 110
rect 204 120 238 154
rect 10 50 44 86
rect 204 50 238 86
rect 44 16 107 50
rect 141 16 204 50
rect 10 0 44 16
rect 204 0 238 16
<< end >>
