* SPICE3 file created from NAND3X1.ext - technology: sky130A

.subckt NAND3X1 Y A B VDD GND
M1000 Y a_599_989# a_372_210.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1001 VDD.t5 A.t0 Y.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 GND A.t1 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1003 VDD.t1 B.t0 Y.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD.t3 a_599_989# Y.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y.t6 A.t2 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y.t0 B.t2 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y.t3 a_599_989# VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 Y a_599_989# 0.26fF
C1 Y B 0.12fF
C2 Y VDD 1.77fF
C3 a_599_989# B 0.18fF
C4 Y A 0.02fF
C5 VDD a_599_989# 0.06fF
C6 VDD B 0.05fF
C7 A a_599_989# 0.02fF
C8 A B 0.18fF
C9 A VDD 0.08fF
R0 A.n0 A.t0 512.525
R1 A.n0 A.t2 371.139
R2 A.n1 A.t1 287.668
R3 A.n1 A.n0 162.713
R4 A.n2 A.n1 76
R5 A.n2 A 0.046
R6 Y.n9 Y.n4 197.352
R7 Y.n9 Y.n8 186.551
R8 Y.n3 Y.n2 79.232
R9 Y.n10 Y.n9 76
R10 Y.n4 Y.n3 63.152
R11 Y.n8 Y.n7 30
R12 Y.n6 Y.n5 24.383
R13 Y.n8 Y.n6 23.684
R14 Y.n4 Y.n0 16.08
R15 Y.n3 Y.n1 16.08
R16 Y.n0 Y.t2 14.282
R17 Y.n0 Y.t3 14.282
R18 Y.n1 Y.t1 14.282
R19 Y.n1 Y.t0 14.282
R20 Y.n2 Y.t5 14.282
R21 Y.n2 Y.t6 14.282
R22 Y.n10 Y 0.046
R23 VDD.n43 VDD.n42 76
R24 VDD.n48 VDD.n47 76
R25 VDD.n98 VDD.n97 76
R26 VDD.n93 VDD.n92 76
R27 VDD.n86 VDD.n85 76
R28 VDD.n81 VDD.n80 76
R29 VDD.n76 VDD.n75 76
R30 VDD.n72 VDD.n71 76
R31 VDD.n27 VDD.n26 64.064
R32 VDD.n83 VDD.n82 59.488
R33 VDD.n77 VDD.t4 55.106
R34 VDD.n30 VDD.t3 55.106
R35 VDD.n88 VDD.n87 40.824
R36 VDD.n41 VDD.n40 40.824
R37 VDD.n35 VDD.n34 34.942
R38 VDD.n38 VDD.n37 27.456
R39 VDD.n90 VDD.n89 22.88
R40 VDD.n71 VDD.n68 21.841
R41 VDD.n23 VDD.n20 21.841
R42 VDD.n87 VDD.t0 14.282
R43 VDD.n87 VDD.t5 14.282
R44 VDD.n40 VDD.t2 14.282
R45 VDD.n40 VDD.t1 14.282
R46 VDD.n68 VDD.n50 14.167
R47 VDD.n50 VDD.n49 14.167
R48 VDD.n20 VDD.n19 14.167
R49 VDD.n19 VDD.n17 14.167
R50 VDD.n33 VDD.n30 14.167
R51 VDD.n30 VDD.n29 14.167
R52 VDD.n95 VDD.n94 13.728
R53 VDD.n23 VDD.n22 13.653
R54 VDD.n22 VDD.n21 13.653
R55 VDD.n33 VDD.n32 13.653
R56 VDD.n32 VDD.n31 13.653
R57 VDD.n30 VDD.n25 13.653
R58 VDD.n25 VDD.n24 13.653
R59 VDD.n29 VDD.n28 13.653
R60 VDD.n28 VDD.n27 13.653
R61 VDD.n42 VDD.n39 13.653
R62 VDD.n39 VDD.n38 13.653
R63 VDD.n47 VDD.n46 13.653
R64 VDD.n46 VDD.n45 13.653
R65 VDD.n97 VDD.n96 13.653
R66 VDD.n96 VDD.n95 13.653
R67 VDD.n92 VDD.n91 13.653
R68 VDD.n91 VDD.n90 13.653
R69 VDD.n85 VDD.n84 13.653
R70 VDD.n84 VDD.n83 13.653
R71 VDD.n80 VDD.n79 13.653
R72 VDD.n79 VDD.n78 13.653
R73 VDD.n75 VDD.n74 13.653
R74 VDD.n74 VDD.n73 13.653
R75 VDD.n71 VDD.n70 13.653
R76 VDD.n70 VDD.n69 13.653
R77 VDD.n4 VDD.n2 12.915
R78 VDD.n4 VDD.n3 12.66
R79 VDD.n12 VDD.n11 12.343
R80 VDD.n10 VDD.n9 12.343
R81 VDD.n7 VDD.n6 12.343
R82 VDD.n45 VDD.n44 9.152
R83 VDD.n54 VDD.n53 7.5
R84 VDD.n57 VDD.n56 7.5
R85 VDD.n59 VDD.n58 7.5
R86 VDD.n62 VDD.n61 7.5
R87 VDD.n68 VDD.n67 7.5
R88 VDD.n20 VDD.n16 7.5
R89 VDD.n2 VDD.n1 7.5
R90 VDD.n6 VDD.n5 7.5
R91 VDD.n9 VDD.n8 7.5
R92 VDD.n19 VDD.n18 7.5
R93 VDD.n14 VDD.n0 7.5
R94 VDD.n67 VDD.n66 6.772
R95 VDD.n55 VDD.n52 6.772
R96 VDD.n60 VDD.n57 6.772
R97 VDD.n64 VDD.n62 6.772
R98 VDD.n64 VDD.n63 6.772
R99 VDD.n60 VDD.n59 6.772
R100 VDD.n55 VDD.n54 6.772
R101 VDD.n66 VDD.n51 6.772
R102 VDD.n92 VDD.n88 6.69
R103 VDD.n34 VDD.n23 6.487
R104 VDD.n34 VDD.n33 6.475
R105 VDD.n16 VDD.n15 6.458
R106 VDD.n42 VDD.n41 6.296
R107 VDD.n14 VDD.n7 1.329
R108 VDD.n14 VDD.n10 1.329
R109 VDD.n14 VDD.n12 1.329
R110 VDD.n14 VDD.n13 1.329
R111 VDD.n15 VDD.n14 0.696
R112 VDD.n14 VDD.n4 0.696
R113 VDD.n80 VDD.n77 0.393
R114 VDD.n65 VDD.n64 0.365
R115 VDD.n65 VDD.n60 0.365
R116 VDD.n65 VDD.n55 0.365
R117 VDD.n66 VDD.n65 0.365
R118 VDD.n72 VDD 0.207
R119 VDD.n36 VDD.n35 0.145
R120 VDD.n43 VDD.n36 0.145
R121 VDD.n48 VDD.n43 0.145
R122 VDD.n98 VDD.n93 0.145
R123 VDD.n93 VDD.n86 0.145
R124 VDD.n86 VDD.n81 0.145
R125 VDD.n81 VDD.n76 0.145
R126 VDD.n76 VDD.n72 0.145
R127 VDD VDD.n48 0.098
R128 VDD VDD.n98 0.098
R129 a_372_210.n10 a_372_210.n8 82.852
R130 a_372_210.n11 a_372_210.n0 49.6
R131 a_372_210.n7 a_372_210.n6 32.833
R132 a_372_210.n8 a_372_210.t1 32.416
R133 a_372_210.n10 a_372_210.n9 27.2
R134 a_372_210.n3 a_372_210.n2 23.284
R135 a_372_210.n11 a_372_210.n10 22.4
R136 a_372_210.n7 a_372_210.n4 19.017
R137 a_372_210.n6 a_372_210.n5 13.494
R138 a_372_210.t1 a_372_210.n1 7.04
R139 a_372_210.t1 a_372_210.n3 5.727
R140 a_372_210.n8 a_372_210.n7 1.435
R141 B.n0 B.t0 479.223
R142 B.n0 B.t2 375.52
R143 B.n1 B.t1 268.26
R144 B.n2 B.n1 76
R145 B.n1 B.n0 69.217
R146 B.n2 B 0.046
R147 a_91_103.t0 a_91_103.n0 117.777
R148 a_91_103.n2 a_91_103.n1 55.228
R149 a_91_103.n4 a_91_103.n3 9.111
R150 a_91_103.t0 a_91_103.n2 4.04
R151 a_91_103.n8 a_91_103.n7 2.455
R152 a_91_103.n6 a_91_103.n4 1.964
R153 a_91_103.n6 a_91_103.n5 1.964
R154 a_91_103.n8 a_91_103.n6 0.636
R155 a_91_103.t0 a_91_103.n8 0.246
R156 GND.n24 GND.n23 85.559
R157 GND.n18 GND.n17 76
R158 GND.n12 GND.n11 76
R159 GND.n15 GND.n14 76
R160 GND.n35 GND.n34 76
R161 GND.n32 GND.n31 76
R162 GND.n29 GND.n28 76
R163 GND.n26 GND.n25 76
R164 GND.n21 GND.n20 76
R165 GND.n8 GND.n7 34.942
R166 GND.n6 GND.n5 14.167
R167 GND.n5 GND.n4 14.167
R168 GND.n20 GND.n19 13.653
R169 GND.n25 GND.n22 13.653
R170 GND.n28 GND.n27 13.653
R171 GND.n31 GND.n30 13.653
R172 GND.n34 GND.n33 13.653
R173 GND.n14 GND.n13 13.653
R174 GND.n11 GND.n10 13.653
R175 GND.n4 GND.n3 13.653
R176 GND.n5 GND.n2 13.653
R177 GND.n6 GND.n1 13.653
R178 GND.n7 GND.n0 7.083
R179 GND.n7 GND.n6 6.474
R180 GND.n17 GND.n16 0.596
R181 GND.n18 GND 0.207
R182 GND.n25 GND.n24 0.196
R183 GND.n9 GND.n8 0.145
R184 GND.n12 GND.n9 0.145
R185 GND.n15 GND.n12 0.145
R186 GND.n35 GND.n32 0.145
R187 GND.n32 GND.n29 0.145
R188 GND.n29 GND.n26 0.145
R189 GND.n26 GND.n21 0.145
R190 GND.n21 GND.n18 0.145
R191 GND GND.n15 0.098
R192 GND GND.n35 0.098
C10 VDD GND 4.23fF
C11 a_91_103.n0 GND 0.03fF
C12 a_91_103.n1 GND 0.10fF
C13 a_91_103.n2 GND 0.10fF
C14 a_91_103.n3 GND 0.04fF
C15 a_91_103.n4 GND 0.03fF
C16 a_91_103.n5 GND 0.03fF
C17 a_91_103.n6 GND 0.03fF
C18 a_91_103.n7 GND 0.04fF
C19 a_372_210.n0 GND 0.02fF
C20 a_372_210.n1 GND 0.09fF
C21 a_372_210.n2 GND 0.13fF
C22 a_372_210.n3 GND 0.11fF
C23 a_372_210.n4 GND 0.09fF
C24 a_372_210.n5 GND 0.05fF
C25 a_372_210.n6 GND 0.01fF
C26 a_372_210.n7 GND 0.03fF
C27 a_372_210.n8 GND 0.11fF
C28 a_372_210.n9 GND 0.02fF
C29 a_372_210.n10 GND 0.05fF
C30 a_372_210.n11 GND 0.02fF
C31 VDD.n0 GND 0.18fF
C32 VDD.n1 GND 0.02fF
C33 VDD.n2 GND 0.02fF
C34 VDD.n3 GND 0.04fF
C35 VDD.n4 GND 0.01fF
C36 VDD.n5 GND 0.02fF
C37 VDD.n6 GND 0.02fF
C38 VDD.n8 GND 0.02fF
C39 VDD.n9 GND 0.02fF
C40 VDD.n11 GND 0.02fF
C41 VDD.n14 GND 0.41fF
C42 VDD.n16 GND 0.03fF
C43 VDD.n17 GND 0.02fF
C44 VDD.n18 GND 0.02fF
C45 VDD.n19 GND 0.02fF
C46 VDD.n20 GND 0.03fF
C47 VDD.n21 GND 0.24fF
C48 VDD.n22 GND 0.02fF
C49 VDD.n23 GND 0.03fF
C50 VDD.n24 GND 0.20fF
C51 VDD.n25 GND 0.01fF
C52 VDD.n26 GND 0.12fF
C53 VDD.n27 GND 0.15fF
C54 VDD.n28 GND 0.01fF
C55 VDD.n29 GND 0.02fF
C56 VDD.n30 GND 0.06fF
C57 VDD.n31 GND 0.24fF
C58 VDD.n32 GND 0.01fF
C59 VDD.n33 GND 0.02fF
C60 VDD.n34 GND 0.00fF
C61 VDD.n35 GND 0.08fF
C62 VDD.n36 GND 0.02fF
C63 VDD.n37 GND 0.12fF
C64 VDD.n38 GND 0.14fF
C65 VDD.n39 GND 0.01fF
C66 VDD.n40 GND 0.09fF
C67 VDD.n41 GND 0.02fF
C68 VDD.n42 GND 0.01fF
C69 VDD.n43 GND 0.02fF
C70 VDD.n44 GND 0.16fF
C71 VDD.n45 GND 0.13fF
C72 VDD.n46 GND 0.01fF
C73 VDD.n47 GND 0.02fF
C74 VDD.n48 GND 0.02fF
C75 VDD.n49 GND 0.02fF
C76 VDD.n50 GND 0.02fF
C77 VDD.n51 GND 0.02fF
C78 VDD.n52 GND 0.02fF
C79 VDD.n53 GND 0.02fF
C80 VDD.n54 GND 0.02fF
C81 VDD.n56 GND 0.02fF
C82 VDD.n57 GND 0.02fF
C83 VDD.n58 GND 0.02fF
C84 VDD.n59 GND 0.02fF
C85 VDD.n61 GND 0.03fF
C86 VDD.n62 GND 0.02fF
C87 VDD.n63 GND 0.18fF
C88 VDD.n65 GND 0.41fF
C89 VDD.n67 GND 0.03fF
C90 VDD.n68 GND 0.03fF
C91 VDD.n69 GND 0.24fF
C92 VDD.n70 GND 0.02fF
C93 VDD.n71 GND 0.03fF
C94 VDD.n72 GND 0.02fF
C95 VDD.n73 GND 0.24fF
C96 VDD.n74 GND 0.01fF
C97 VDD.n75 GND 0.02fF
C98 VDD.n76 GND 0.02fF
C99 VDD.n77 GND 0.05fF
C100 VDD.n78 GND 0.20fF
C101 VDD.n79 GND 0.01fF
C102 VDD.n80 GND 0.01fF
C103 VDD.n81 GND 0.02fF
C104 VDD.n82 GND 0.12fF
C105 VDD.n83 GND 0.15fF
C106 VDD.n84 GND 0.01fF
C107 VDD.n85 GND 0.02fF
C108 VDD.n86 GND 0.02fF
C109 VDD.n87 GND 0.09fF
C110 VDD.n88 GND 0.02fF
C111 VDD.n89 GND 0.12fF
C112 VDD.n90 GND 0.14fF
C113 VDD.n91 GND 0.01fF
C114 VDD.n92 GND 0.01fF
C115 VDD.n93 GND 0.02fF
C116 VDD.n94 GND 0.16fF
C117 VDD.n95 GND 0.13fF
C118 VDD.n96 GND 0.01fF
C119 VDD.n97 GND 0.02fF
C120 VDD.n98 GND 0.02fF
C121 Y.n0 GND 0.42fF
C122 Y.n1 GND 0.42fF
C123 Y.n2 GND 0.49fF
C124 Y.n3 GND 0.16fF
C125 Y.n4 GND 0.26fF
C126 Y.n5 GND 0.03fF
C127 Y.n6 GND 0.04fF
C128 Y.n7 GND 0.03fF
C129 Y.n8 GND 0.21fF
C130 Y.n9 GND 0.35fF
C131 Y.n10 GND 0.01fF
.ends
