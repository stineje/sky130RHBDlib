magic
tech sky130A
magscale 1 2
timestamp 1669507576
<< nwell >>
rect -87 786 2529 1550
<< pwell >>
rect -34 -34 2476 544
<< nmos >>
rect 168 288 198 349
tri 198 288 214 304 sw
rect 362 296 392 349
tri 392 296 408 312 sw
rect 168 258 274 288
tri 274 258 304 288 sw
rect 362 266 468 296
tri 468 266 498 296 sw
rect 168 157 198 258
tri 198 242 214 258 nw
tri 258 242 274 258 ne
tri 198 157 214 173 sw
tri 258 157 274 173 se
rect 274 157 304 258
rect 362 165 392 266
tri 392 250 408 266 nw
tri 452 250 468 266 ne
tri 392 165 408 181 sw
tri 452 165 468 181 se
rect 468 165 498 266
tri 168 127 198 157 ne
rect 198 127 274 157
tri 274 127 304 157 nw
tri 362 135 392 165 ne
rect 392 135 468 165
tri 468 135 498 165 nw
rect 834 296 864 349
tri 864 296 880 312 sw
rect 1028 296 1058 349
tri 1058 296 1074 312 sw
rect 834 266 940 296
tri 940 266 970 296 sw
rect 834 165 864 266
tri 864 250 880 266 nw
tri 924 250 940 266 ne
tri 864 165 880 181 sw
tri 924 165 940 181 se
rect 940 165 970 266
rect 1028 266 1134 296
tri 1134 266 1164 296 sw
rect 1028 251 1059 266
tri 1059 251 1074 266 nw
tri 1118 251 1133 266 ne
rect 1133 251 1164 266
tri 834 135 864 165 ne
rect 864 135 940 165
tri 940 135 970 165 nw
rect 1028 165 1058 251
tri 1058 165 1074 181 sw
tri 1118 165 1134 181 se
rect 1134 165 1164 251
tri 1028 135 1058 165 ne
rect 1058 135 1134 165
tri 1134 135 1164 165 nw
rect 1500 288 1530 349
tri 1530 288 1546 304 sw
rect 1694 296 1724 349
tri 1724 296 1740 312 sw
rect 1500 258 1606 288
tri 1606 258 1636 288 sw
rect 1694 266 1800 296
tri 1800 266 1830 296 sw
rect 1500 157 1530 258
tri 1530 242 1546 258 nw
tri 1590 242 1606 258 ne
tri 1530 157 1546 173 sw
tri 1590 157 1606 173 se
rect 1606 157 1636 258
rect 1694 165 1724 266
tri 1724 250 1740 266 nw
tri 1784 250 1800 266 ne
tri 1724 165 1740 181 sw
tri 1784 165 1800 181 se
rect 1800 165 1830 266
tri 1500 127 1530 157 ne
rect 1530 127 1606 157
tri 1606 127 1636 157 nw
tri 1694 135 1724 165 ne
rect 1724 135 1800 165
tri 1800 135 1830 165 nw
rect 2153 297 2183 350
tri 2183 297 2199 313 sw
rect 2153 267 2259 297
tri 2259 267 2289 297 sw
rect 2153 166 2183 267
tri 2183 251 2199 267 nw
tri 2243 251 2259 267 ne
tri 2183 166 2199 182 sw
tri 2243 166 2259 182 se
rect 2259 166 2289 267
tri 2153 136 2183 166 ne
rect 2183 136 2259 166
tri 2259 136 2289 166 nw
<< pmos >>
rect 187 1004 217 1404
rect 275 1004 305 1404
rect 363 1004 393 1404
rect 451 1004 481 1404
rect 853 1005 883 1405
rect 941 1005 971 1405
rect 1029 1005 1059 1405
rect 1117 1005 1147 1405
rect 1519 1004 1549 1404
rect 1607 1004 1637 1404
rect 1695 1004 1725 1404
rect 1783 1004 1813 1404
rect 2162 1004 2192 1404
rect 2250 1004 2280 1404
<< ndiff >>
rect 112 333 168 349
rect 112 299 122 333
rect 156 299 168 333
rect 112 261 168 299
rect 198 333 362 349
rect 198 304 219 333
tri 198 288 214 304 ne
rect 214 299 219 304
rect 253 299 316 333
rect 350 299 362 333
rect 214 288 362 299
rect 392 312 554 349
tri 392 296 408 312 ne
rect 408 296 554 312
rect 112 227 122 261
rect 156 227 168 261
tri 274 258 304 288 ne
rect 304 261 362 288
tri 468 266 498 296 ne
rect 112 193 168 227
rect 112 159 122 193
rect 156 159 168 193
rect 112 127 168 159
tri 198 242 214 258 se
rect 214 242 258 258
tri 258 242 274 258 sw
rect 198 208 274 242
rect 198 174 219 208
rect 253 174 274 208
rect 198 173 274 174
tri 198 157 214 173 ne
rect 214 157 258 173
tri 258 157 274 173 nw
rect 304 227 316 261
rect 350 227 362 261
rect 304 193 362 227
rect 304 159 316 193
rect 350 159 362 193
tri 392 250 408 266 se
rect 408 250 452 266
tri 452 250 468 266 sw
rect 392 217 468 250
rect 392 183 413 217
rect 447 183 468 217
rect 392 181 468 183
tri 392 165 408 181 ne
rect 408 165 452 181
tri 452 165 468 181 nw
rect 498 261 554 296
rect 498 227 510 261
rect 544 227 554 261
rect 498 193 554 227
tri 168 127 198 157 sw
tri 274 127 304 157 se
rect 304 135 362 159
tri 362 135 392 165 sw
tri 468 135 498 165 se
rect 498 159 510 193
rect 544 159 554 193
rect 498 135 554 159
rect 304 127 554 135
rect 112 123 554 127
rect 112 89 122 123
rect 156 89 316 123
rect 350 89 413 123
rect 447 89 510 123
rect 544 89 554 123
rect 112 73 554 89
rect 778 333 834 349
rect 778 299 788 333
rect 822 299 834 333
rect 778 261 834 299
rect 864 312 1028 349
tri 864 296 880 312 ne
rect 880 296 1028 312
rect 1058 312 1220 349
tri 1058 296 1074 312 ne
rect 1074 296 1220 312
tri 940 266 970 296 ne
rect 778 227 788 261
rect 822 227 834 261
rect 778 193 834 227
rect 778 159 788 193
rect 822 159 834 193
tri 864 250 880 266 se
rect 880 250 924 266
tri 924 250 940 266 sw
rect 864 217 940 250
rect 864 183 885 217
rect 919 183 940 217
rect 864 181 940 183
tri 864 165 880 181 ne
rect 880 165 924 181
tri 924 165 940 181 nw
rect 970 261 1028 296
tri 1134 266 1164 296 ne
rect 970 227 982 261
rect 1016 227 1028 261
tri 1059 251 1074 266 se
rect 1074 251 1118 266
tri 1118 251 1133 266 sw
rect 1164 261 1220 296
rect 970 193 1028 227
rect 778 135 834 159
tri 834 135 864 165 sw
tri 940 135 970 165 se
rect 970 159 982 193
rect 1016 159 1028 193
rect 1058 217 1134 251
rect 1058 183 1079 217
rect 1113 183 1134 217
rect 1058 181 1134 183
tri 1058 165 1074 181 ne
rect 1074 165 1118 181
tri 1118 165 1134 181 nw
rect 1164 227 1176 261
rect 1210 227 1220 261
rect 1164 193 1220 227
rect 970 135 1028 159
tri 1028 135 1058 165 sw
tri 1134 135 1164 165 se
rect 1164 159 1176 193
rect 1210 159 1220 193
rect 1164 135 1220 159
rect 778 123 1220 135
rect 778 89 788 123
rect 822 89 885 123
rect 919 89 982 123
rect 1016 89 1079 123
rect 1113 89 1176 123
rect 1210 89 1220 123
rect 778 73 1220 89
rect 1444 333 1500 349
rect 1444 299 1454 333
rect 1488 299 1500 333
rect 1444 261 1500 299
rect 1530 333 1694 349
rect 1530 304 1551 333
tri 1530 288 1546 304 ne
rect 1546 299 1551 304
rect 1585 299 1648 333
rect 1682 299 1694 333
rect 1546 288 1694 299
rect 1724 312 1886 349
tri 1724 296 1740 312 ne
rect 1740 296 1886 312
rect 1444 227 1454 261
rect 1488 227 1500 261
tri 1606 258 1636 288 ne
rect 1636 261 1694 288
tri 1800 266 1830 296 ne
rect 1444 193 1500 227
rect 1444 159 1454 193
rect 1488 159 1500 193
rect 1444 127 1500 159
tri 1530 242 1546 258 se
rect 1546 242 1590 258
tri 1590 242 1606 258 sw
rect 1530 208 1606 242
rect 1530 174 1551 208
rect 1585 174 1606 208
rect 1530 173 1606 174
tri 1530 157 1546 173 ne
rect 1546 157 1590 173
tri 1590 157 1606 173 nw
rect 1636 227 1648 261
rect 1682 227 1694 261
rect 1636 193 1694 227
rect 1636 159 1648 193
rect 1682 159 1694 193
tri 1724 250 1740 266 se
rect 1740 250 1784 266
tri 1784 250 1800 266 sw
rect 1724 217 1800 250
rect 1724 183 1745 217
rect 1779 183 1800 217
rect 1724 181 1800 183
tri 1724 165 1740 181 ne
rect 1740 165 1784 181
tri 1784 165 1800 181 nw
rect 1830 261 1886 296
rect 1830 227 1842 261
rect 1876 227 1886 261
rect 1830 193 1886 227
tri 1500 127 1530 157 sw
tri 1606 127 1636 157 se
rect 1636 135 1694 159
tri 1694 135 1724 165 sw
tri 1800 135 1830 165 se
rect 1830 159 1842 193
rect 1876 159 1886 193
rect 1830 135 1886 159
rect 1636 127 1886 135
rect 1444 123 1886 127
rect 1444 89 1454 123
rect 1488 89 1648 123
rect 1682 89 1745 123
rect 1779 89 1842 123
rect 1876 89 1886 123
rect 1444 73 1886 89
rect 2097 334 2153 350
rect 2097 300 2107 334
rect 2141 300 2153 334
rect 2097 262 2153 300
rect 2183 334 2343 350
rect 2183 313 2301 334
tri 2183 297 2199 313 ne
rect 2199 300 2301 313
rect 2335 300 2343 334
rect 2199 297 2343 300
tri 2259 267 2289 297 ne
rect 2097 228 2107 262
rect 2141 228 2153 262
rect 2097 194 2153 228
rect 2097 160 2107 194
rect 2141 160 2153 194
tri 2183 251 2199 267 se
rect 2199 251 2243 267
tri 2243 251 2259 267 sw
rect 2183 218 2259 251
rect 2183 184 2203 218
rect 2237 184 2259 218
rect 2183 182 2259 184
tri 2183 166 2199 182 ne
rect 2199 166 2243 182
tri 2243 166 2259 182 nw
rect 2289 262 2343 297
rect 2289 228 2301 262
rect 2335 228 2343 262
rect 2289 194 2343 228
rect 2097 136 2153 160
tri 2153 136 2183 166 sw
tri 2259 136 2289 166 se
rect 2289 160 2301 194
rect 2335 160 2343 194
rect 2289 136 2343 160
rect 2097 124 2343 136
rect 2097 90 2107 124
rect 2141 90 2203 124
rect 2237 90 2301 124
rect 2335 90 2343 124
rect 2097 74 2343 90
<< pdiff >>
rect 131 1366 187 1404
rect 131 1332 141 1366
rect 175 1332 187 1366
rect 131 1298 187 1332
rect 131 1264 141 1298
rect 175 1264 187 1298
rect 131 1230 187 1264
rect 131 1196 141 1230
rect 175 1196 187 1230
rect 131 1162 187 1196
rect 131 1128 141 1162
rect 175 1128 187 1162
rect 131 1093 187 1128
rect 131 1059 141 1093
rect 175 1059 187 1093
rect 131 1004 187 1059
rect 217 1366 275 1404
rect 217 1332 229 1366
rect 263 1332 275 1366
rect 217 1298 275 1332
rect 217 1264 229 1298
rect 263 1264 275 1298
rect 217 1230 275 1264
rect 217 1196 229 1230
rect 263 1196 275 1230
rect 217 1162 275 1196
rect 217 1128 229 1162
rect 263 1128 275 1162
rect 217 1093 275 1128
rect 217 1059 229 1093
rect 263 1059 275 1093
rect 217 1004 275 1059
rect 305 1366 363 1404
rect 305 1332 317 1366
rect 351 1332 363 1366
rect 305 1298 363 1332
rect 305 1264 317 1298
rect 351 1264 363 1298
rect 305 1230 363 1264
rect 305 1196 317 1230
rect 351 1196 363 1230
rect 305 1162 363 1196
rect 305 1128 317 1162
rect 351 1128 363 1162
rect 305 1004 363 1128
rect 393 1366 451 1404
rect 393 1332 405 1366
rect 439 1332 451 1366
rect 393 1298 451 1332
rect 393 1264 405 1298
rect 439 1264 451 1298
rect 393 1230 451 1264
rect 393 1196 405 1230
rect 439 1196 451 1230
rect 393 1162 451 1196
rect 393 1128 405 1162
rect 439 1128 451 1162
rect 393 1093 451 1128
rect 393 1059 405 1093
rect 439 1059 451 1093
rect 393 1004 451 1059
rect 481 1366 535 1404
rect 481 1332 493 1366
rect 527 1332 535 1366
rect 481 1298 535 1332
rect 481 1264 493 1298
rect 527 1264 535 1298
rect 481 1230 535 1264
rect 481 1196 493 1230
rect 527 1196 535 1230
rect 481 1162 535 1196
rect 481 1128 493 1162
rect 527 1128 535 1162
rect 481 1004 535 1128
rect 797 1365 853 1405
rect 797 1331 807 1365
rect 841 1331 853 1365
rect 797 1297 853 1331
rect 797 1263 807 1297
rect 841 1263 853 1297
rect 797 1229 853 1263
rect 797 1195 807 1229
rect 841 1195 853 1229
rect 797 1161 853 1195
rect 797 1127 807 1161
rect 841 1127 853 1161
rect 797 1093 853 1127
rect 797 1059 807 1093
rect 841 1059 853 1093
rect 797 1005 853 1059
rect 883 1365 941 1405
rect 883 1331 895 1365
rect 929 1331 941 1365
rect 883 1297 941 1331
rect 883 1263 895 1297
rect 929 1263 941 1297
rect 883 1229 941 1263
rect 883 1195 895 1229
rect 929 1195 941 1229
rect 883 1161 941 1195
rect 883 1127 895 1161
rect 929 1127 941 1161
rect 883 1005 941 1127
rect 971 1365 1029 1405
rect 971 1331 983 1365
rect 1017 1331 1029 1365
rect 971 1297 1029 1331
rect 971 1263 983 1297
rect 1017 1263 1029 1297
rect 971 1229 1029 1263
rect 971 1195 983 1229
rect 1017 1195 1029 1229
rect 971 1161 1029 1195
rect 971 1127 983 1161
rect 1017 1127 1029 1161
rect 971 1093 1029 1127
rect 971 1059 983 1093
rect 1017 1059 1029 1093
rect 971 1005 1029 1059
rect 1059 1297 1117 1405
rect 1059 1263 1071 1297
rect 1105 1263 1117 1297
rect 1059 1229 1117 1263
rect 1059 1195 1071 1229
rect 1105 1195 1117 1229
rect 1059 1161 1117 1195
rect 1059 1127 1071 1161
rect 1105 1127 1117 1161
rect 1059 1093 1117 1127
rect 1059 1059 1071 1093
rect 1105 1059 1117 1093
rect 1059 1005 1117 1059
rect 1147 1365 1201 1405
rect 1147 1331 1159 1365
rect 1193 1331 1201 1365
rect 1147 1297 1201 1331
rect 1147 1263 1159 1297
rect 1193 1263 1201 1297
rect 1147 1229 1201 1263
rect 1147 1195 1159 1229
rect 1193 1195 1201 1229
rect 1147 1161 1201 1195
rect 1147 1127 1159 1161
rect 1193 1127 1201 1161
rect 1147 1005 1201 1127
rect 1463 1366 1519 1404
rect 1463 1332 1473 1366
rect 1507 1332 1519 1366
rect 1463 1298 1519 1332
rect 1463 1264 1473 1298
rect 1507 1264 1519 1298
rect 1463 1230 1519 1264
rect 1463 1196 1473 1230
rect 1507 1196 1519 1230
rect 1463 1162 1519 1196
rect 1463 1128 1473 1162
rect 1507 1128 1519 1162
rect 1463 1093 1519 1128
rect 1463 1059 1473 1093
rect 1507 1059 1519 1093
rect 1463 1004 1519 1059
rect 1549 1366 1607 1404
rect 1549 1332 1561 1366
rect 1595 1332 1607 1366
rect 1549 1298 1607 1332
rect 1549 1264 1561 1298
rect 1595 1264 1607 1298
rect 1549 1230 1607 1264
rect 1549 1196 1561 1230
rect 1595 1196 1607 1230
rect 1549 1162 1607 1196
rect 1549 1128 1561 1162
rect 1595 1128 1607 1162
rect 1549 1093 1607 1128
rect 1549 1059 1561 1093
rect 1595 1059 1607 1093
rect 1549 1004 1607 1059
rect 1637 1366 1695 1404
rect 1637 1332 1649 1366
rect 1683 1332 1695 1366
rect 1637 1298 1695 1332
rect 1637 1264 1649 1298
rect 1683 1264 1695 1298
rect 1637 1230 1695 1264
rect 1637 1196 1649 1230
rect 1683 1196 1695 1230
rect 1637 1162 1695 1196
rect 1637 1128 1649 1162
rect 1683 1128 1695 1162
rect 1637 1004 1695 1128
rect 1725 1366 1783 1404
rect 1725 1332 1737 1366
rect 1771 1332 1783 1366
rect 1725 1298 1783 1332
rect 1725 1264 1737 1298
rect 1771 1264 1783 1298
rect 1725 1230 1783 1264
rect 1725 1196 1737 1230
rect 1771 1196 1783 1230
rect 1725 1162 1783 1196
rect 1725 1128 1737 1162
rect 1771 1128 1783 1162
rect 1725 1093 1783 1128
rect 1725 1059 1737 1093
rect 1771 1059 1783 1093
rect 1725 1004 1783 1059
rect 1813 1366 1867 1404
rect 1813 1332 1825 1366
rect 1859 1332 1867 1366
rect 1813 1298 1867 1332
rect 1813 1264 1825 1298
rect 1859 1264 1867 1298
rect 1813 1230 1867 1264
rect 1813 1196 1825 1230
rect 1859 1196 1867 1230
rect 1813 1162 1867 1196
rect 1813 1128 1825 1162
rect 1859 1128 1867 1162
rect 1813 1004 1867 1128
rect 2106 1366 2162 1404
rect 2106 1332 2116 1366
rect 2150 1332 2162 1366
rect 2106 1298 2162 1332
rect 2106 1264 2116 1298
rect 2150 1264 2162 1298
rect 2106 1230 2162 1264
rect 2106 1196 2116 1230
rect 2150 1196 2162 1230
rect 2106 1162 2162 1196
rect 2106 1128 2116 1162
rect 2150 1128 2162 1162
rect 2106 1093 2162 1128
rect 2106 1059 2116 1093
rect 2150 1059 2162 1093
rect 2106 1004 2162 1059
rect 2192 1366 2250 1404
rect 2192 1332 2204 1366
rect 2238 1332 2250 1366
rect 2192 1298 2250 1332
rect 2192 1264 2204 1298
rect 2238 1264 2250 1298
rect 2192 1230 2250 1264
rect 2192 1196 2204 1230
rect 2238 1196 2250 1230
rect 2192 1162 2250 1196
rect 2192 1128 2204 1162
rect 2238 1128 2250 1162
rect 2192 1093 2250 1128
rect 2192 1059 2204 1093
rect 2238 1059 2250 1093
rect 2192 1004 2250 1059
rect 2280 1366 2334 1404
rect 2280 1332 2292 1366
rect 2326 1332 2334 1366
rect 2280 1298 2334 1332
rect 2280 1264 2292 1298
rect 2326 1264 2334 1298
rect 2280 1230 2334 1264
rect 2280 1196 2292 1230
rect 2326 1196 2334 1230
rect 2280 1162 2334 1196
rect 2280 1128 2292 1162
rect 2326 1128 2334 1162
rect 2280 1093 2334 1128
rect 2280 1059 2292 1093
rect 2326 1059 2334 1093
rect 2280 1004 2334 1059
<< ndiffc >>
rect 122 299 156 333
rect 219 299 253 333
rect 316 299 350 333
rect 122 227 156 261
rect 122 159 156 193
rect 219 174 253 208
rect 316 227 350 261
rect 316 159 350 193
rect 413 183 447 217
rect 510 227 544 261
rect 510 159 544 193
rect 122 89 156 123
rect 316 89 350 123
rect 413 89 447 123
rect 510 89 544 123
rect 788 299 822 333
rect 788 227 822 261
rect 788 159 822 193
rect 885 183 919 217
rect 982 227 1016 261
rect 982 159 1016 193
rect 1079 183 1113 217
rect 1176 227 1210 261
rect 1176 159 1210 193
rect 788 89 822 123
rect 885 89 919 123
rect 982 89 1016 123
rect 1079 89 1113 123
rect 1176 89 1210 123
rect 1454 299 1488 333
rect 1551 299 1585 333
rect 1648 299 1682 333
rect 1454 227 1488 261
rect 1454 159 1488 193
rect 1551 174 1585 208
rect 1648 227 1682 261
rect 1648 159 1682 193
rect 1745 183 1779 217
rect 1842 227 1876 261
rect 1842 159 1876 193
rect 1454 89 1488 123
rect 1648 89 1682 123
rect 1745 89 1779 123
rect 1842 89 1876 123
rect 2107 300 2141 334
rect 2301 300 2335 334
rect 2107 228 2141 262
rect 2107 160 2141 194
rect 2203 184 2237 218
rect 2301 228 2335 262
rect 2301 160 2335 194
rect 2107 90 2141 124
rect 2203 90 2237 124
rect 2301 90 2335 124
<< pdiffc >>
rect 141 1332 175 1366
rect 141 1264 175 1298
rect 141 1196 175 1230
rect 141 1128 175 1162
rect 141 1059 175 1093
rect 229 1332 263 1366
rect 229 1264 263 1298
rect 229 1196 263 1230
rect 229 1128 263 1162
rect 229 1059 263 1093
rect 317 1332 351 1366
rect 317 1264 351 1298
rect 317 1196 351 1230
rect 317 1128 351 1162
rect 405 1332 439 1366
rect 405 1264 439 1298
rect 405 1196 439 1230
rect 405 1128 439 1162
rect 405 1059 439 1093
rect 493 1332 527 1366
rect 493 1264 527 1298
rect 493 1196 527 1230
rect 493 1128 527 1162
rect 807 1331 841 1365
rect 807 1263 841 1297
rect 807 1195 841 1229
rect 807 1127 841 1161
rect 807 1059 841 1093
rect 895 1331 929 1365
rect 895 1263 929 1297
rect 895 1195 929 1229
rect 895 1127 929 1161
rect 983 1331 1017 1365
rect 983 1263 1017 1297
rect 983 1195 1017 1229
rect 983 1127 1017 1161
rect 983 1059 1017 1093
rect 1071 1263 1105 1297
rect 1071 1195 1105 1229
rect 1071 1127 1105 1161
rect 1071 1059 1105 1093
rect 1159 1331 1193 1365
rect 1159 1263 1193 1297
rect 1159 1195 1193 1229
rect 1159 1127 1193 1161
rect 1473 1332 1507 1366
rect 1473 1264 1507 1298
rect 1473 1196 1507 1230
rect 1473 1128 1507 1162
rect 1473 1059 1507 1093
rect 1561 1332 1595 1366
rect 1561 1264 1595 1298
rect 1561 1196 1595 1230
rect 1561 1128 1595 1162
rect 1561 1059 1595 1093
rect 1649 1332 1683 1366
rect 1649 1264 1683 1298
rect 1649 1196 1683 1230
rect 1649 1128 1683 1162
rect 1737 1332 1771 1366
rect 1737 1264 1771 1298
rect 1737 1196 1771 1230
rect 1737 1128 1771 1162
rect 1737 1059 1771 1093
rect 1825 1332 1859 1366
rect 1825 1264 1859 1298
rect 1825 1196 1859 1230
rect 1825 1128 1859 1162
rect 2116 1332 2150 1366
rect 2116 1264 2150 1298
rect 2116 1196 2150 1230
rect 2116 1128 2150 1162
rect 2116 1059 2150 1093
rect 2204 1332 2238 1366
rect 2204 1264 2238 1298
rect 2204 1196 2238 1230
rect 2204 1128 2238 1162
rect 2204 1059 2238 1093
rect 2292 1332 2326 1366
rect 2292 1264 2326 1298
rect 2292 1196 2326 1230
rect 2292 1128 2326 1162
rect 2292 1059 2326 1093
<< psubdiff >>
rect -34 482 2476 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 632 461 700 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 632 427 649 461
rect 683 427 700 461
rect 1298 461 1366 482
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 632 313 700 353
rect 1298 427 1315 461
rect 1349 427 1366 461
rect 1964 461 2032 482
rect 1298 387 1366 427
rect 1298 353 1315 387
rect 1349 353 1366 387
rect 632 279 649 313
rect 683 279 700 313
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect -34 17 34 57
rect 632 57 649 91
rect 683 57 700 91
rect 1298 313 1366 353
rect 1964 427 1981 461
rect 2015 427 2032 461
rect 2408 461 2476 482
rect 1964 387 2032 427
rect 1964 353 1981 387
rect 2015 353 2032 387
rect 2408 427 2425 461
rect 2459 427 2476 461
rect 1298 279 1315 313
rect 1349 279 1366 313
rect 1298 239 1366 279
rect 1298 205 1315 239
rect 1349 205 1366 239
rect 1298 165 1366 205
rect 1298 131 1315 165
rect 1349 131 1366 165
rect 1298 91 1366 131
rect 632 17 700 57
rect 1298 57 1315 91
rect 1349 57 1366 91
rect 1964 313 2032 353
rect 2408 387 2476 427
rect 2408 353 2425 387
rect 2459 353 2476 387
rect 1964 279 1981 313
rect 2015 279 2032 313
rect 1964 239 2032 279
rect 1964 205 1981 239
rect 2015 205 2032 239
rect 1964 165 2032 205
rect 1964 131 1981 165
rect 2015 131 2032 165
rect 1964 91 2032 131
rect 1298 17 1366 57
rect 1964 57 1981 91
rect 2015 57 2032 91
rect 2408 313 2476 353
rect 2408 279 2425 313
rect 2459 279 2476 313
rect 2408 239 2476 279
rect 2408 205 2425 239
rect 2459 205 2476 239
rect 2408 165 2476 205
rect 2408 131 2425 165
rect 2459 131 2476 165
rect 2408 91 2476 131
rect 1964 17 2032 57
rect 2408 57 2425 91
rect 2459 57 2476 91
rect 2408 17 2476 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2476 17
rect -34 -34 2476 -17
<< nsubdiff >>
rect -34 1497 2476 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2476 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 632 1423 700 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 1298 1423 1366 1463
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 632 979 700 1019
rect 1298 1389 1315 1423
rect 1349 1389 1366 1423
rect 1964 1423 2032 1463
rect 1298 1349 1366 1389
rect 1298 1315 1315 1349
rect 1349 1315 1366 1349
rect 1298 1275 1366 1315
rect 1298 1241 1315 1275
rect 1349 1241 1366 1275
rect 1298 1201 1366 1241
rect 1298 1167 1315 1201
rect 1349 1167 1366 1201
rect 1298 1127 1366 1167
rect 1298 1093 1315 1127
rect 1349 1093 1366 1127
rect 1298 1053 1366 1093
rect 1298 1019 1315 1053
rect 1349 1019 1366 1053
rect 632 945 649 979
rect 683 945 700 979
rect -34 871 -17 905
rect 17 884 34 905
rect 632 905 700 945
rect 1298 979 1366 1019
rect 1964 1389 1981 1423
rect 2015 1389 2032 1423
rect 2408 1423 2476 1463
rect 1964 1349 2032 1389
rect 1964 1315 1981 1349
rect 2015 1315 2032 1349
rect 1964 1275 2032 1315
rect 1964 1241 1981 1275
rect 2015 1241 2032 1275
rect 1964 1201 2032 1241
rect 1964 1167 1981 1201
rect 2015 1167 2032 1201
rect 1964 1127 2032 1167
rect 1964 1093 1981 1127
rect 2015 1093 2032 1127
rect 1964 1053 2032 1093
rect 1964 1019 1981 1053
rect 2015 1019 2032 1053
rect 1298 945 1315 979
rect 1349 945 1366 979
rect 632 884 649 905
rect 17 871 649 884
rect 683 884 700 905
rect 1298 905 1366 945
rect 1964 979 2032 1019
rect 2408 1389 2425 1423
rect 2459 1389 2476 1423
rect 2408 1349 2476 1389
rect 2408 1315 2425 1349
rect 2459 1315 2476 1349
rect 2408 1275 2476 1315
rect 2408 1241 2425 1275
rect 2459 1241 2476 1275
rect 2408 1201 2476 1241
rect 2408 1167 2425 1201
rect 2459 1167 2476 1201
rect 2408 1127 2476 1167
rect 2408 1093 2425 1127
rect 2459 1093 2476 1127
rect 2408 1053 2476 1093
rect 2408 1019 2425 1053
rect 2459 1019 2476 1053
rect 1964 945 1981 979
rect 2015 945 2032 979
rect 1298 884 1315 905
rect 683 871 1315 884
rect 1349 884 1366 905
rect 1964 905 2032 945
rect 2408 979 2476 1019
rect 2408 945 2425 979
rect 2459 945 2476 979
rect 1964 884 1981 905
rect 1349 871 1981 884
rect 2015 884 2032 905
rect 2408 905 2476 945
rect 2408 884 2425 905
rect 2015 871 2425 884
rect 2459 871 2476 905
rect -34 822 2476 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 649 427 683 461
rect 649 353 683 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1315 427 1349 461
rect 1315 353 1349 387
rect 649 279 683 313
rect 649 205 683 239
rect 649 131 683 165
rect 649 57 683 91
rect 1981 427 2015 461
rect 1981 353 2015 387
rect 2425 427 2459 461
rect 1315 279 1349 313
rect 1315 205 1349 239
rect 1315 131 1349 165
rect 1315 57 1349 91
rect 2425 353 2459 387
rect 1981 279 2015 313
rect 1981 205 2015 239
rect 1981 131 2015 165
rect 1981 57 2015 91
rect 2425 279 2459 313
rect 2425 205 2459 239
rect 2425 131 2459 165
rect 2425 57 2459 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 649 1389 683 1423
rect 649 1315 683 1349
rect 649 1241 683 1275
rect 649 1167 683 1201
rect 649 1093 683 1127
rect 649 1019 683 1053
rect -17 945 17 979
rect 1315 1389 1349 1423
rect 1315 1315 1349 1349
rect 1315 1241 1349 1275
rect 1315 1167 1349 1201
rect 1315 1093 1349 1127
rect 1315 1019 1349 1053
rect 649 945 683 979
rect -17 871 17 905
rect 1981 1389 2015 1423
rect 1981 1315 2015 1349
rect 1981 1241 2015 1275
rect 1981 1167 2015 1201
rect 1981 1093 2015 1127
rect 1981 1019 2015 1053
rect 1315 945 1349 979
rect 649 871 683 905
rect 2425 1389 2459 1423
rect 2425 1315 2459 1349
rect 2425 1241 2459 1275
rect 2425 1167 2459 1201
rect 2425 1093 2459 1127
rect 2425 1019 2459 1053
rect 1981 945 2015 979
rect 1315 871 1349 905
rect 2425 945 2459 979
rect 1981 871 2015 905
rect 2425 871 2459 905
<< poly >>
rect 187 1404 217 1430
rect 275 1404 305 1430
rect 363 1404 393 1430
rect 451 1404 481 1430
rect 853 1405 883 1431
rect 941 1405 971 1431
rect 1029 1405 1059 1431
rect 1117 1405 1147 1431
rect 187 973 217 1004
rect 275 973 305 1004
rect 363 973 393 1004
rect 451 973 481 1004
rect 187 957 305 973
rect 187 943 205 957
rect 195 923 205 943
rect 239 943 305 957
rect 349 957 481 973
rect 239 923 249 943
rect 195 907 249 923
rect 349 923 359 957
rect 393 943 481 957
rect 1519 1404 1549 1430
rect 1607 1404 1637 1430
rect 1695 1404 1725 1430
rect 1783 1404 1813 1430
rect 853 974 883 1005
rect 941 974 971 1005
rect 1029 974 1059 1005
rect 1117 974 1147 1005
rect 393 923 403 943
rect 349 907 403 923
rect 830 958 971 974
rect 830 924 840 958
rect 874 944 971 958
rect 1016 958 1147 974
rect 874 924 884 944
rect 830 908 884 924
rect 1016 924 1026 958
rect 1060 944 1147 958
rect 2162 1404 2192 1430
rect 2250 1404 2280 1430
rect 1060 924 1070 944
rect 1016 908 1070 924
rect 1519 973 1549 1004
rect 1607 973 1637 1004
rect 1695 973 1725 1004
rect 1783 973 1813 1004
rect 1519 957 1637 973
rect 1519 943 1537 957
rect 1527 923 1537 943
rect 1571 943 1637 957
rect 1681 957 1813 973
rect 1571 923 1581 943
rect 1527 907 1581 923
rect 1681 923 1691 957
rect 1725 943 1813 957
rect 2162 973 2192 1004
rect 2250 973 2280 1004
rect 1725 923 1735 943
rect 1681 907 1735 923
rect 2119 957 2280 973
rect 2119 923 2129 957
rect 2163 943 2280 957
rect 2163 923 2173 943
rect 2119 907 2173 923
rect 195 433 249 449
rect 195 413 205 433
rect 168 399 205 413
rect 239 399 249 433
rect 168 383 249 399
rect 343 433 397 449
rect 343 399 353 433
rect 387 399 397 433
rect 343 383 397 399
rect 861 433 915 449
rect 861 413 871 433
rect 168 349 198 383
rect 362 349 392 383
rect 834 399 871 413
rect 905 399 915 433
rect 834 383 915 399
rect 1009 433 1063 449
rect 1009 399 1019 433
rect 1053 399 1063 433
rect 1009 383 1063 399
rect 1527 433 1581 449
rect 1527 413 1537 433
rect 834 349 864 383
rect 1028 349 1058 383
rect 1500 399 1537 413
rect 1571 399 1581 433
rect 1500 383 1581 399
rect 1675 433 1729 449
rect 1675 399 1685 433
rect 1719 399 1729 433
rect 1675 383 1729 399
rect 1500 349 1530 383
rect 1694 349 1724 383
rect 2119 434 2173 450
rect 2119 400 2129 434
rect 2163 413 2173 434
rect 2163 400 2183 413
rect 2119 384 2183 400
rect 2153 350 2183 384
<< polycont >>
rect 205 923 239 957
rect 359 923 393 957
rect 840 924 874 958
rect 1026 924 1060 958
rect 1537 923 1571 957
rect 1691 923 1725 957
rect 2129 923 2163 957
rect 205 399 239 433
rect 353 399 387 433
rect 871 399 905 433
rect 1019 399 1053 433
rect 1537 399 1571 433
rect 1685 399 1719 433
rect 2129 400 2163 434
<< locali >>
rect -34 1497 2476 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2476 1497
rect -34 1446 2476 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 141 1366 175 1446
rect 141 1298 175 1332
rect 141 1230 175 1264
rect 141 1162 175 1196
rect 141 1093 175 1128
rect 141 1027 175 1059
rect 229 1366 263 1404
rect 229 1298 263 1332
rect 229 1230 263 1264
rect 229 1162 263 1196
rect 229 1093 263 1128
rect 317 1366 351 1446
rect 317 1298 351 1332
rect 317 1230 351 1264
rect 317 1162 351 1196
rect 317 1111 351 1128
rect 405 1366 439 1404
rect 405 1298 439 1332
rect 405 1230 439 1264
rect 405 1162 439 1196
rect 229 1057 263 1059
rect 405 1093 439 1128
rect 493 1366 527 1446
rect 493 1298 527 1332
rect 493 1230 527 1264
rect 493 1162 527 1196
rect 493 1111 527 1128
rect 632 1423 700 1446
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 405 1057 439 1059
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 229 1023 535 1057
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 359 957 393 973
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 923
rect 205 383 239 399
rect 353 923 359 942
rect 353 907 393 923
rect 353 433 387 907
rect 353 383 387 399
rect 501 535 535 1023
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect 807 1365 841 1405
rect 807 1297 841 1331
rect 807 1229 841 1263
rect 807 1161 841 1195
rect 807 1093 841 1127
rect 895 1365 929 1446
rect 1298 1423 1366 1446
rect 895 1297 929 1331
rect 895 1229 929 1263
rect 895 1161 929 1195
rect 895 1111 929 1127
rect 983 1365 1193 1399
rect 983 1297 1017 1331
rect 983 1229 1017 1263
rect 983 1161 1017 1195
rect 983 1093 1017 1127
rect 807 1025 1017 1059
rect 1071 1297 1105 1313
rect 1071 1229 1105 1263
rect 1071 1161 1105 1195
rect 1071 1093 1105 1127
rect 1159 1297 1193 1331
rect 1159 1229 1193 1263
rect 1159 1161 1193 1195
rect 1159 1111 1193 1127
rect 1298 1389 1315 1423
rect 1349 1389 1366 1423
rect 1298 1349 1366 1389
rect 1298 1315 1315 1349
rect 1349 1315 1366 1349
rect 1298 1275 1366 1315
rect 1298 1241 1315 1275
rect 1349 1241 1366 1275
rect 1298 1201 1366 1241
rect 1298 1167 1315 1201
rect 1349 1167 1366 1201
rect 1298 1127 1366 1167
rect 1298 1093 1315 1127
rect 1349 1093 1366 1127
rect 1071 1025 1201 1059
rect 632 979 700 1019
rect 632 945 649 979
rect 683 945 700 979
rect 632 905 700 945
rect 840 958 874 974
rect 1026 958 1060 974
rect 874 924 905 942
rect 840 908 905 924
rect 632 871 649 905
rect 683 871 700 905
rect 632 822 700 871
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 122 333 156 349
rect 316 333 350 349
rect 501 348 535 501
rect 156 299 219 333
rect 253 299 316 333
rect 122 261 156 299
rect 122 193 156 227
rect 316 261 350 299
rect 122 123 156 159
rect 122 73 156 89
rect 219 208 253 224
rect -34 34 34 57
rect 219 34 253 174
rect 316 193 350 227
rect 413 314 535 348
rect 632 461 700 544
rect 632 427 649 461
rect 683 427 700 461
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect 871 535 905 908
rect 871 433 905 501
rect 871 383 905 399
rect 1019 924 1026 942
rect 1019 908 1060 924
rect 1019 433 1053 908
rect 1019 383 1053 399
rect 1167 535 1201 1025
rect 1298 1053 1366 1093
rect 1298 1019 1315 1053
rect 1349 1019 1366 1053
rect 1473 1366 1507 1446
rect 1473 1298 1507 1332
rect 1473 1230 1507 1264
rect 1473 1162 1507 1196
rect 1473 1093 1507 1128
rect 1473 1027 1507 1059
rect 1561 1366 1595 1404
rect 1561 1298 1595 1332
rect 1561 1230 1595 1264
rect 1561 1162 1595 1196
rect 1561 1093 1595 1128
rect 1649 1366 1683 1446
rect 1649 1298 1683 1332
rect 1649 1230 1683 1264
rect 1649 1162 1683 1196
rect 1649 1111 1683 1128
rect 1737 1366 1771 1404
rect 1737 1298 1771 1332
rect 1737 1230 1771 1264
rect 1737 1162 1771 1196
rect 1561 1057 1595 1059
rect 1737 1093 1771 1128
rect 1825 1366 1859 1446
rect 1825 1298 1859 1332
rect 1825 1230 1859 1264
rect 1825 1162 1859 1196
rect 1825 1111 1859 1128
rect 1964 1423 2032 1446
rect 1964 1389 1981 1423
rect 2015 1389 2032 1423
rect 1964 1349 2032 1389
rect 1964 1315 1981 1349
rect 2015 1315 2032 1349
rect 1964 1275 2032 1315
rect 1964 1241 1981 1275
rect 2015 1241 2032 1275
rect 1964 1201 2032 1241
rect 1964 1167 1981 1201
rect 2015 1167 2032 1201
rect 1964 1127 2032 1167
rect 1737 1057 1771 1059
rect 1964 1093 1981 1127
rect 2015 1093 2032 1127
rect 1561 1023 1867 1057
rect 1298 979 1366 1019
rect 1298 945 1315 979
rect 1349 945 1366 979
rect 1298 905 1366 945
rect 1298 871 1315 905
rect 1349 871 1366 905
rect 1298 822 1366 871
rect 1537 957 1571 973
rect 1691 957 1725 973
rect 413 217 447 314
rect 632 313 700 353
rect 632 279 649 313
rect 683 279 700 313
rect 413 167 447 183
rect 510 261 544 277
rect 510 193 544 227
rect 316 123 350 159
rect 510 123 544 159
rect 350 89 413 123
rect 447 89 510 123
rect 316 73 350 89
rect 510 73 544 89
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect 632 57 649 91
rect 683 57 700 91
rect 632 34 700 57
rect 788 333 822 349
rect 1167 348 1201 501
rect 788 261 822 299
rect 788 193 822 227
rect 885 314 1201 348
rect 1298 461 1366 544
rect 1298 427 1315 461
rect 1349 427 1366 461
rect 1298 387 1366 427
rect 1298 353 1315 387
rect 1349 353 1366 387
rect 1537 535 1571 923
rect 1537 433 1571 501
rect 1537 383 1571 399
rect 1685 923 1691 942
rect 1685 907 1725 923
rect 1685 433 1719 907
rect 1685 383 1719 399
rect 1833 535 1867 1023
rect 1964 1053 2032 1093
rect 1964 1019 1981 1053
rect 2015 1019 2032 1053
rect 2116 1366 2150 1446
rect 2116 1298 2150 1332
rect 2116 1230 2150 1264
rect 2116 1162 2150 1196
rect 2116 1093 2150 1128
rect 2116 1037 2150 1059
rect 2204 1366 2238 1404
rect 2204 1298 2238 1332
rect 2204 1230 2238 1264
rect 2204 1162 2238 1196
rect 2204 1093 2238 1128
rect 1964 979 2032 1019
rect 1964 945 1981 979
rect 2015 945 2032 979
rect 1964 905 2032 945
rect 1964 871 1981 905
rect 2015 871 2032 905
rect 1964 822 2032 871
rect 2129 957 2163 973
rect 885 217 919 314
rect 885 167 919 183
rect 982 261 1016 278
rect 982 193 1016 227
rect 788 123 822 159
rect 1079 217 1113 314
rect 1298 313 1366 353
rect 1298 279 1315 313
rect 1349 279 1366 313
rect 1079 167 1113 183
rect 1176 261 1210 278
rect 1176 193 1210 227
rect 982 123 1016 159
rect 1176 123 1210 159
rect 822 89 885 123
rect 919 89 982 123
rect 1016 89 1079 123
rect 1113 89 1176 123
rect 788 34 822 89
rect 885 34 919 89
rect 982 34 1016 89
rect 1079 34 1113 89
rect 1176 34 1210 89
rect 1298 239 1366 279
rect 1298 205 1315 239
rect 1349 205 1366 239
rect 1298 165 1366 205
rect 1298 131 1315 165
rect 1349 131 1366 165
rect 1298 91 1366 131
rect 1298 57 1315 91
rect 1349 57 1366 91
rect 1454 333 1488 349
rect 1648 333 1682 349
rect 1833 348 1867 501
rect 1488 299 1551 333
rect 1585 299 1648 333
rect 1454 261 1488 299
rect 1454 193 1488 227
rect 1648 261 1682 299
rect 1454 123 1488 159
rect 1454 73 1488 89
rect 1551 208 1585 224
rect 1298 34 1366 57
rect 1551 34 1585 174
rect 1648 193 1682 227
rect 1745 314 1867 348
rect 1964 461 2032 544
rect 1964 427 1981 461
rect 2015 427 2032 461
rect 1964 387 2032 427
rect 1964 353 1981 387
rect 2015 353 2032 387
rect 2129 535 2163 923
rect 2204 933 2238 1059
rect 2292 1366 2326 1446
rect 2292 1298 2326 1332
rect 2292 1230 2326 1264
rect 2292 1162 2326 1196
rect 2292 1093 2326 1128
rect 2292 1037 2326 1059
rect 2408 1423 2476 1446
rect 2408 1389 2425 1423
rect 2459 1389 2476 1423
rect 2408 1349 2476 1389
rect 2408 1315 2425 1349
rect 2459 1315 2476 1349
rect 2408 1275 2476 1315
rect 2408 1241 2425 1275
rect 2459 1241 2476 1275
rect 2408 1201 2476 1241
rect 2408 1167 2425 1201
rect 2459 1167 2476 1201
rect 2408 1127 2476 1167
rect 2408 1093 2425 1127
rect 2459 1093 2476 1127
rect 2408 1053 2476 1093
rect 2408 1019 2425 1053
rect 2459 1019 2476 1053
rect 2408 979 2476 1019
rect 2408 945 2425 979
rect 2459 945 2476 979
rect 2204 899 2311 933
rect 2129 434 2163 501
rect 2277 433 2311 899
rect 2408 905 2476 945
rect 2408 871 2425 905
rect 2459 871 2476 905
rect 2408 822 2476 871
rect 2129 384 2163 400
rect 2203 399 2311 433
rect 2408 461 2476 544
rect 2408 427 2425 461
rect 2459 427 2476 461
rect 1745 217 1779 314
rect 1964 313 2032 353
rect 1964 279 1981 313
rect 2015 279 2032 313
rect 1745 167 1779 183
rect 1842 261 1876 277
rect 1842 193 1876 227
rect 1648 123 1682 159
rect 1842 123 1876 159
rect 1682 89 1745 123
rect 1779 89 1842 123
rect 1648 73 1682 89
rect 1842 73 1876 89
rect 1964 239 2032 279
rect 1964 205 1981 239
rect 2015 205 2032 239
rect 1964 165 2032 205
rect 1964 131 1981 165
rect 2015 131 2032 165
rect 1964 91 2032 131
rect 1964 57 1981 91
rect 2015 57 2032 91
rect 1964 34 2032 57
rect 2107 334 2141 350
rect 2107 262 2141 300
rect 2107 194 2141 228
rect 2203 218 2237 399
rect 2408 387 2476 427
rect 2408 353 2425 387
rect 2459 353 2476 387
rect 2203 168 2237 184
rect 2301 334 2335 350
rect 2301 262 2335 300
rect 2301 194 2335 228
rect 2107 124 2141 160
rect 2301 124 2335 160
rect 2141 90 2203 124
rect 2237 90 2301 124
rect 2107 34 2141 90
rect 2204 34 2238 90
rect 2301 34 2335 90
rect 2408 313 2476 353
rect 2408 279 2425 313
rect 2459 279 2476 313
rect 2408 239 2476 279
rect 2408 205 2425 239
rect 2459 205 2476 239
rect 2408 165 2476 205
rect 2408 131 2425 165
rect 2459 131 2476 165
rect 2408 91 2476 131
rect 2408 57 2425 91
rect 2459 57 2476 91
rect 2408 34 2476 57
rect -34 17 2476 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2476 17
rect -34 -34 2476 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 501 501 535 535
rect 871 501 905 535
rect 1167 501 1201 535
rect 1537 501 1571 535
rect 1833 501 1867 535
rect 2129 501 2163 535
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
<< metal1 >>
rect -34 1497 2476 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2476 1497
rect -34 1446 2476 1463
rect 495 535 541 541
rect 865 535 911 541
rect 1161 535 1207 541
rect 1531 535 1577 541
rect 1827 535 1873 541
rect 2123 535 2169 541
rect 489 501 501 535
rect 535 501 871 535
rect 905 501 917 535
rect 1155 501 1167 535
rect 1201 501 1537 535
rect 1571 501 1583 535
rect 1821 501 1833 535
rect 1867 501 2129 535
rect 2163 501 2175 535
rect 495 495 541 501
rect 865 495 911 501
rect 1161 495 1207 501
rect 1531 495 1577 501
rect 1827 495 1873 501
rect 2123 495 2169 501
rect -34 17 2476 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2476 17
rect -34 -34 2476 -17
<< labels >>
rlabel metal1 2277 575 2311 609 1 Y
port 1 n
rlabel metal1 2277 501 2311 535 1 Y
port 2 n
rlabel metal1 2277 427 2311 461 1 Y
port 3 n
rlabel metal1 2277 649 2311 683 1 Y
port 4 n
rlabel metal1 2277 723 2311 757 1 Y
port 5 n
rlabel metal1 2277 797 2311 831 1 Y
port 6 n
rlabel metal1 2277 871 2311 905 1 Y
port 7 n
rlabel metal1 205 575 239 609 1 A
port 8 n
rlabel metal1 205 501 239 535 1 A
port 9 n
rlabel metal1 205 427 239 461 1 A
port 10 n
rlabel metal1 205 649 239 683 1 A
port 11 n
rlabel metal1 205 723 239 757 1 A
port 12 n
rlabel metal1 205 797 239 831 1 A
port 13 n
rlabel metal1 205 871 239 905 1 A
port 14 n
rlabel metal1 353 649 387 683 1 B
port 15 n
rlabel metal1 353 723 387 757 1 B
port 16 n
rlabel metal1 353 871 387 905 1 B
port 17 n
rlabel metal1 353 797 387 831 1 B
port 18 n
rlabel metal1 353 575 387 609 1 B
port 19 n
rlabel metal1 353 501 387 535 1 B
port 20 n
rlabel metal1 353 427 387 461 1 B
port 21 n
rlabel metal1 1019 723 1053 757 1 C
port 22 n
rlabel metal1 1019 797 1053 831 1 C
port 23 n
rlabel metal1 1019 871 1053 905 1 C
port 24 n
rlabel metal1 1019 649 1053 683 1 C
port 25 n
rlabel metal1 1019 575 1053 609 1 C
port 26 n
rlabel metal1 1019 501 1053 535 1 C
port 27 n
rlabel metal1 1019 427 1053 461 1 C
port 28 n
rlabel metal1 1685 797 1719 831 1 D
port 29 n
rlabel metal1 1685 723 1719 757 1 D
port 30 n
rlabel metal1 1685 649 1719 683 1 D
port 31 n
rlabel metal1 1685 575 1719 609 1 D
port 32 n
rlabel metal1 1685 501 1719 535 1 D
port 33 n
rlabel metal1 1685 427 1719 461 1 D
port 34 n
rlabel metal1 1685 871 1719 905 1 D
port 35 n
rlabel metal1 -34 1446 2476 1514 1 VPWR
port 36 n
rlabel metal1 -34 -34 2476 34 1 VGND
port 37 n
rlabel nwell 57 1463 91 1497 1 VPB
port 38 n
rlabel pwell 57 -17 91 17 1 VNB
port 39 n
<< end >>
