magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect 2174 10255 2612 10987
<< mvpmos >>
rect 2293 10321 2493 10921
<< mvpdiff >>
rect 2240 10909 2293 10921
rect 2240 10875 2248 10909
rect 2282 10875 2293 10909
rect 2240 10841 2293 10875
rect 2240 10807 2248 10841
rect 2282 10807 2293 10841
rect 2240 10773 2293 10807
rect 2240 10739 2248 10773
rect 2282 10739 2293 10773
rect 2240 10705 2293 10739
rect 2240 10671 2248 10705
rect 2282 10671 2293 10705
rect 2240 10637 2293 10671
rect 2240 10603 2248 10637
rect 2282 10603 2293 10637
rect 2240 10569 2293 10603
rect 2240 10535 2248 10569
rect 2282 10535 2293 10569
rect 2240 10501 2293 10535
rect 2240 10467 2248 10501
rect 2282 10467 2293 10501
rect 2240 10433 2293 10467
rect 2240 10399 2248 10433
rect 2282 10399 2293 10433
rect 2240 10321 2293 10399
rect 2493 10909 2546 10921
rect 2493 10875 2504 10909
rect 2538 10875 2546 10909
rect 2493 10841 2546 10875
rect 2493 10807 2504 10841
rect 2538 10807 2546 10841
rect 2493 10773 2546 10807
rect 2493 10739 2504 10773
rect 2538 10739 2546 10773
rect 2493 10705 2546 10739
rect 2493 10671 2504 10705
rect 2538 10671 2546 10705
rect 2493 10637 2546 10671
rect 2493 10603 2504 10637
rect 2538 10603 2546 10637
rect 2493 10569 2546 10603
rect 2493 10535 2504 10569
rect 2538 10535 2546 10569
rect 2493 10501 2546 10535
rect 2493 10467 2504 10501
rect 2538 10467 2546 10501
rect 2493 10433 2546 10467
rect 2493 10399 2504 10433
rect 2538 10399 2546 10433
rect 2493 10321 2546 10399
<< mvpdiffc >>
rect 2248 10875 2282 10909
rect 2248 10807 2282 10841
rect 2248 10739 2282 10773
rect 2248 10671 2282 10705
rect 2248 10603 2282 10637
rect 2248 10535 2282 10569
rect 2248 10467 2282 10501
rect 2248 10399 2282 10433
rect 2504 10875 2538 10909
rect 2504 10807 2538 10841
rect 2504 10739 2538 10773
rect 2504 10671 2538 10705
rect 2504 10603 2538 10637
rect 2504 10535 2538 10569
rect 2504 10467 2538 10501
rect 2504 10399 2538 10433
<< poly >>
rect 2293 10921 2493 10947
rect 2293 10271 2493 10321
rect 2293 10237 2309 10271
rect 2343 10237 2443 10271
rect 2477 10237 2493 10271
rect 2293 10221 2493 10237
<< polycont >>
rect 2309 10237 2343 10271
rect 2443 10237 2477 10271
<< locali >>
rect 2248 10909 2282 10925
rect 2248 10852 2282 10875
rect 2248 10773 2282 10807
rect 2248 10705 2282 10731
rect 2248 10637 2282 10644
rect 2248 10591 2282 10603
rect 2248 10503 2282 10535
rect 2248 10433 2282 10467
rect 2248 10383 2282 10399
rect 2504 10909 2538 10925
rect 2504 10841 2538 10875
rect 2504 10773 2538 10807
rect 2504 10705 2538 10739
rect 2504 10637 2538 10646
rect 2504 10569 2538 10574
rect 2504 10433 2538 10467
rect 2504 10383 2538 10399
rect 2339 10271 2447 10279
rect 2293 10245 2305 10271
rect 2293 10237 2309 10245
rect 2343 10237 2443 10271
rect 2481 10245 2493 10271
rect 2477 10237 2493 10245
rect 1713 8686 1943 8857
rect 792 7224 1045 7394
rect 12586 2220 13114 2286
rect 9652 1863 9686 1976
rect 10290 1863 10324 1976
rect 11104 1863 11138 1976
rect 11484 1863 11518 1976
rect 11770 1863 11804 1976
rect 12232 1863 12266 1976
rect 12526 1863 12560 1976
rect 12878 1863 12912 1976
rect 13230 1863 13264 1976
rect 12702 1784 12736 1822
rect 13054 1784 13088 1822
rect 9652 1594 9686 1707
rect 10290 1594 10324 1707
rect 11104 1594 11138 1707
rect 11770 1595 11804 1708
rect 12232 1595 12266 1708
rect 12526 1595 12560 1708
rect 12878 1595 12912 1708
rect 13230 1595 13264 1708
rect 12323 1318 12357 1356
rect 12409 1317 12443 1355
rect 12621 1317 12655 1355
rect 12796 1317 12830 1355
rect 12973 1317 13007 1355
rect 13153 1317 13187 1355
rect 12674 937 13114 1003
<< viali >>
rect 2248 10841 2282 10852
rect 2248 10818 2282 10841
rect 2248 10739 2282 10765
rect 2248 10731 2282 10739
rect 2248 10671 2282 10678
rect 2248 10644 2282 10671
rect 2248 10569 2282 10591
rect 2248 10557 2282 10569
rect 2248 10501 2282 10503
rect 2248 10469 2282 10501
rect 2504 10671 2538 10680
rect 2504 10646 2538 10671
rect 2504 10603 2538 10608
rect 2504 10574 2538 10603
rect 2504 10501 2538 10535
rect 2305 10271 2339 10279
rect 2447 10271 2481 10279
rect 2305 10245 2309 10271
rect 2309 10245 2339 10271
rect 2447 10245 2477 10271
rect 2477 10245 2481 10271
rect 12702 1822 12736 1856
rect 12702 1750 12736 1784
rect 13054 1822 13088 1856
rect 13054 1750 13088 1784
rect 12323 1356 12357 1390
rect 12323 1284 12357 1318
rect 12409 1355 12443 1389
rect 12409 1283 12443 1317
rect 12621 1355 12655 1389
rect 12621 1283 12655 1317
rect 12796 1355 12830 1389
rect 12796 1283 12830 1317
rect 12973 1355 13007 1389
rect 12973 1283 13007 1317
rect 13153 1355 13187 1389
rect 13153 1283 13187 1317
<< metal1 >>
tri 1728 14645 1741 14658 se
rect 1741 14645 2589 14658
rect 1650 14639 2589 14645
rect 1766 14574 2589 14639
tri 1766 14530 1810 14574 nw
rect 1650 14517 1766 14523
rect 6192 14499 6267 14545
rect 25669 14501 25704 14541
rect 3681 14418 3687 14470
rect 3739 14418 3751 14470
rect 3803 14418 3809 14470
rect 2866 14338 2872 14390
rect 2924 14338 2936 14390
rect 2988 14338 2994 14390
rect 3178 13760 3184 13812
rect 3236 13760 3248 13812
rect 3300 13760 3306 13812
tri 2240 10862 2242 10864 se
rect 2242 10862 2288 10864
tri 1620 10852 1630 10862 sw
tri 2230 10852 2240 10862 se
rect 2240 10852 2288 10862
rect 1620 10827 1630 10852
tri 1630 10827 1655 10852 sw
tri 2205 10827 2230 10852 se
rect 2230 10827 2248 10852
rect 1620 10818 2248 10827
rect 2282 10818 2288 10852
rect 1620 10785 2288 10818
rect 1620 10765 1644 10785
tri 1644 10765 1664 10785 nw
tri 2203 10765 2223 10785 ne
rect 2223 10765 2288 10785
tri 1620 10741 1644 10765 nw
tri 2223 10746 2242 10765 ne
rect 2242 10731 2248 10765
rect 2282 10731 2288 10765
rect 2242 10678 2288 10731
tri 3097 10692 3110 10705 se
rect 2242 10644 2248 10678
rect 2282 10644 2288 10678
rect 2242 10591 2288 10644
rect 2242 10557 2248 10591
rect 2282 10557 2288 10591
rect 2242 10503 2288 10557
rect 2242 10469 2248 10503
rect 2282 10469 2288 10503
rect 2498 10680 2649 10692
rect 2498 10646 2504 10680
rect 2538 10646 2649 10680
rect 2498 10640 2649 10646
rect 2650 10641 2651 10691
rect 2711 10641 2712 10691
rect 2713 10641 3110 10692
rect 2713 10640 2765 10641
tri 3074 10640 3075 10641 ne
rect 3075 10640 3110 10641
rect 2498 10608 2562 10640
rect 2498 10574 2504 10608
rect 2538 10605 2562 10608
tri 2562 10605 2597 10640 nw
tri 3075 10605 3110 10640 ne
rect 2538 10574 2544 10605
tri 2544 10587 2562 10605 nw
rect 2498 10535 2544 10574
rect 2498 10501 2504 10535
rect 2538 10501 2544 10535
rect 2498 10489 2544 10501
rect 2958 10509 3010 10515
rect 2242 10457 2288 10469
tri 3010 10502 3023 10515 sw
rect 3010 10457 3117 10502
rect 2958 10451 3117 10457
rect 2958 10445 3010 10451
tri 3010 10418 3043 10451 nw
rect 3111 10450 3117 10451
rect 3169 10450 3181 10502
rect 3233 10450 3239 10502
rect 2958 10387 3010 10393
rect 2293 10279 3254 10285
rect 2293 10245 2305 10279
rect 2339 10245 2447 10279
rect 2481 10253 3254 10279
rect 2481 10247 3200 10253
rect 2481 10245 2493 10247
rect 2293 10239 2493 10245
tri 2493 10239 2501 10247 nw
rect 3252 10247 3254 10253
rect 3200 10189 3252 10201
rect 3200 10131 3252 10137
rect 1117 7749 1478 7812
rect 26813 7501 26941 7502
rect 26356 7497 26553 7498
rect 26356 7445 26362 7497
rect 26414 7445 26429 7497
rect 26481 7445 26495 7497
rect 26547 7445 26553 7497
rect 26356 7427 26553 7445
rect 26356 7375 26362 7427
rect 26414 7375 26429 7427
rect 26481 7375 26495 7427
rect 26547 7375 26553 7427
rect 26356 7357 26553 7375
rect 26356 7305 26362 7357
rect 26414 7305 26429 7357
rect 26481 7305 26495 7357
rect 26547 7305 26553 7357
rect 26813 7449 26819 7501
rect 26871 7449 26883 7501
rect 26935 7449 26941 7501
rect 26813 7431 26941 7449
rect 26813 7379 26819 7431
rect 26871 7379 26883 7431
rect 26935 7379 26941 7431
rect 26813 7361 26941 7379
rect 26813 7309 26819 7361
rect 26871 7309 26883 7361
rect 26935 7309 26941 7361
rect 26813 7308 26941 7309
rect 26356 7304 26553 7305
rect 27219 6810 27283 6811
rect 26356 6808 26553 6809
rect 26356 6756 26362 6808
rect 26414 6756 26429 6808
rect 26481 6756 26495 6808
rect 26547 6756 26553 6808
rect 26356 6738 26553 6756
rect 26356 6686 26362 6738
rect 26414 6686 26429 6738
rect 26481 6686 26495 6738
rect 26547 6686 26553 6738
rect 26356 6668 26553 6686
rect 26356 6616 26362 6668
rect 26414 6616 26429 6668
rect 26481 6616 26495 6668
rect 26547 6616 26553 6668
rect 26356 6615 26553 6616
rect 26616 6808 26813 6809
rect 26616 6756 26622 6808
rect 26674 6756 26689 6808
rect 26741 6756 26755 6808
rect 26807 6756 26813 6808
rect 26616 6738 26813 6756
rect 26616 6686 26622 6738
rect 26674 6686 26689 6738
rect 26741 6686 26755 6738
rect 26807 6686 26813 6738
rect 26616 6668 26813 6686
rect 26616 6616 26622 6668
rect 26674 6616 26689 6668
rect 26741 6616 26755 6668
rect 26807 6616 26813 6668
rect 27219 6758 27225 6810
rect 27277 6758 27283 6810
rect 27219 6740 27283 6758
rect 27219 6688 27225 6740
rect 27277 6688 27283 6740
rect 27219 6670 27283 6688
rect 27219 6618 27225 6670
rect 27277 6618 27283 6670
rect 27219 6617 27283 6618
rect 26616 6615 26813 6616
rect 26722 4969 26868 4975
rect 26774 4917 26816 4969
rect 26722 4874 26868 4917
rect 26774 4822 26816 4874
rect 26722 4816 26868 4822
rect 26535 4469 26684 4518
tri 26684 4469 26721 4506 sw
rect 26535 4463 26868 4469
rect 26535 4411 26722 4463
rect 26774 4411 26816 4463
rect 26535 4368 26868 4411
rect 26535 4344 26722 4368
tri 26535 4310 26569 4344 ne
rect 26569 4316 26722 4344
rect 26774 4316 26816 4368
rect 26569 4310 26868 4316
tri 6752 2154 6763 2165 se
rect 6763 2154 6814 2165
rect 6535 2115 6814 2154
rect 6441 2052 6814 2115
rect 6535 1964 6814 2052
tri 6710 1963 6711 1964 ne
rect 6711 1963 6814 1964
rect 6870 2031 6876 2083
rect 6928 2031 6943 2083
rect 6995 2031 7010 2083
rect 7062 2031 7077 2083
rect 7129 2031 7144 2083
rect 7196 2031 7210 2083
rect 7262 2031 7268 2083
rect 6870 2015 7268 2031
rect 6870 1963 6876 2015
rect 6928 1963 6943 2015
rect 6995 1963 7010 2015
rect 7062 1963 7077 2015
rect 7129 1963 7144 2015
rect 7196 1963 7210 2015
rect 7262 1963 7268 2015
rect 12425 1964 12572 2165
rect 12425 1963 13276 1964
rect 12278 1935 13276 1963
rect 12425 1890 13276 1935
rect 12690 1856 13152 1862
rect 13154 1861 13190 1862
rect 12690 1822 12702 1856
rect 12736 1822 13054 1856
rect 13088 1822 13152 1856
rect 12690 1784 13152 1822
rect 12690 1750 12702 1784
rect 12736 1750 13054 1784
rect 13088 1750 13152 1784
rect 12690 1744 13152 1750
rect 13153 1745 13191 1861
rect 13154 1744 13190 1745
rect 13192 1744 13405 1862
tri 13315 1714 13345 1744 ne
rect 13345 1714 13405 1744
rect 3272 1658 3278 1710
rect 3330 1658 3342 1710
rect 3394 1658 3400 1710
rect 12278 1437 13282 1714
tri 13345 1704 13355 1714 ne
rect 12317 1397 12369 1403
rect 12317 1333 12369 1345
rect 12317 1152 12369 1281
rect 12403 1389 13193 1401
rect 12403 1355 12409 1389
rect 12443 1355 12621 1389
rect 12655 1355 12796 1389
rect 12830 1355 12973 1389
rect 13007 1355 13153 1389
rect 13187 1355 13193 1389
rect 12403 1317 13193 1355
rect 12403 1283 12409 1317
rect 12443 1283 12621 1317
rect 12655 1283 12796 1317
rect 12830 1283 12973 1317
rect 13007 1283 13153 1317
rect 13187 1283 13193 1317
rect 12403 1271 13193 1283
tri 12369 1152 12391 1174 sw
tri 12317 1078 12391 1152 ne
tri 12391 1078 12465 1152 sw
tri 12391 1014 12455 1078 ne
rect 12455 1022 12465 1078
tri 12465 1022 12521 1078 sw
rect 12455 1014 12521 1022
rect 3066 961 3072 1013
rect 3124 961 3136 1013
rect 3188 961 3194 1013
rect 10526 944 10611 982
rect 10816 962 10888 1014
tri 12455 1013 12456 1014 ne
rect 12456 1013 12521 1014
tri 12456 1004 12465 1013 ne
rect 12465 1004 12521 1013
tri 12465 1000 12469 1004 ne
rect 11943 880 12003 912
rect 12469 853 12521 1004
rect 12469 801 12475 853
rect 12527 801 12539 853
rect 12591 801 12597 853
rect 7753 749 7852 795
rect 2664 300 2917 470
rect 13355 264 13405 1714
rect 6870 189 6876 241
rect 6928 189 6943 241
rect 6995 189 7010 241
rect 7062 189 7077 241
rect 7129 189 7144 241
rect 7196 189 7210 241
rect 7262 189 7268 241
rect 13277 212 13283 264
rect 13335 212 13347 264
rect 13399 212 13405 264
rect 6870 173 7268 189
rect 6870 121 6876 173
rect 6928 121 6943 173
rect 6995 121 7010 173
rect 7062 121 7077 173
rect 7129 121 7144 173
rect 7196 121 7210 173
rect 7262 121 7268 173
<< rmetal1 >>
rect 2649 10691 2651 10692
rect 2649 10641 2650 10691
rect 2649 10640 2651 10641
rect 2711 10691 2713 10692
rect 2712 10641 2713 10691
rect 2711 10640 2713 10641
rect 13152 1861 13154 1862
rect 13190 1861 13192 1862
rect 13152 1745 13153 1861
rect 13191 1745 13192 1861
rect 13152 1744 13154 1745
rect 13190 1744 13192 1745
<< via1 >>
rect 1650 14523 1766 14639
rect 3687 14418 3739 14470
rect 3751 14418 3803 14470
rect 2872 14338 2924 14390
rect 2936 14338 2988 14390
rect 3184 13760 3236 13812
rect 3248 13760 3300 13812
rect 2958 10457 3010 10509
rect 2958 10393 3010 10445
rect 3117 10450 3169 10502
rect 3181 10450 3233 10502
rect 3200 10201 3252 10253
rect 3200 10137 3252 10189
rect 26362 7445 26414 7497
rect 26429 7445 26481 7497
rect 26495 7445 26547 7497
rect 26362 7375 26414 7427
rect 26429 7375 26481 7427
rect 26495 7375 26547 7427
rect 26362 7305 26414 7357
rect 26429 7305 26481 7357
rect 26495 7305 26547 7357
rect 26819 7449 26871 7501
rect 26883 7449 26935 7501
rect 26819 7379 26871 7431
rect 26883 7379 26935 7431
rect 26819 7309 26871 7361
rect 26883 7309 26935 7361
rect 26362 6756 26414 6808
rect 26429 6756 26481 6808
rect 26495 6756 26547 6808
rect 26362 6686 26414 6738
rect 26429 6686 26481 6738
rect 26495 6686 26547 6738
rect 26362 6616 26414 6668
rect 26429 6616 26481 6668
rect 26495 6616 26547 6668
rect 26622 6756 26674 6808
rect 26689 6756 26741 6808
rect 26755 6756 26807 6808
rect 26622 6686 26674 6738
rect 26689 6686 26741 6738
rect 26755 6686 26807 6738
rect 26622 6616 26674 6668
rect 26689 6616 26741 6668
rect 26755 6616 26807 6668
rect 27225 6758 27277 6810
rect 27225 6688 27277 6740
rect 27225 6618 27277 6670
rect 26722 4917 26774 4969
rect 26816 4917 26868 4969
rect 26722 4822 26774 4874
rect 26816 4822 26868 4874
rect 26722 4411 26774 4463
rect 26816 4411 26868 4463
rect 26722 4316 26774 4368
rect 26816 4316 26868 4368
rect 6876 2031 6928 2083
rect 6943 2031 6995 2083
rect 7010 2031 7062 2083
rect 7077 2031 7129 2083
rect 7144 2031 7196 2083
rect 7210 2031 7262 2083
rect 6876 1963 6928 2015
rect 6943 1963 6995 2015
rect 7010 1963 7062 2015
rect 7077 1963 7129 2015
rect 7144 1963 7196 2015
rect 7210 1963 7262 2015
rect 3278 1658 3330 1710
rect 3342 1658 3394 1710
rect 12317 1390 12369 1397
rect 12317 1356 12323 1390
rect 12323 1356 12357 1390
rect 12357 1356 12369 1390
rect 12317 1345 12369 1356
rect 12317 1318 12369 1333
rect 12317 1284 12323 1318
rect 12323 1284 12357 1318
rect 12357 1284 12369 1318
rect 12317 1281 12369 1284
rect 3072 961 3124 1013
rect 3136 961 3188 1013
rect 12475 801 12527 853
rect 12539 801 12591 853
rect 6876 189 6928 241
rect 6943 189 6995 241
rect 7010 189 7062 241
rect 7077 189 7129 241
rect 7144 189 7196 241
rect 7210 189 7262 241
rect 13283 212 13335 264
rect 13347 212 13399 264
rect 6876 121 6928 173
rect 6943 121 6995 173
rect 7010 121 7062 173
rect 7077 121 7129 173
rect 7144 121 7196 173
rect 7210 121 7262 173
<< metal2 >>
rect 1638 14667 1766 14676
rect 1638 14639 1674 14667
rect 1730 14639 1766 14667
rect 1638 14523 1650 14639
rect 1638 14517 1766 14523
rect 3681 14418 3687 14470
rect 3739 14418 3751 14470
rect 3803 14418 3809 14470
tri 3688 14390 3716 14418 ne
rect 2866 14338 2872 14390
rect 2924 14338 2936 14390
rect 2988 14374 3064 14390
tri 3064 14374 3080 14390 sw
rect 2988 14338 3080 14374
tri 3017 14315 3040 14338 ne
rect 2958 10509 3010 10515
rect 2958 10445 3010 10457
rect 2958 9090 3010 10393
rect 3040 9942 3080 14338
rect 3178 13812 3187 13814
rect 3243 13812 3267 13814
rect 3178 13760 3184 13812
rect 3243 13760 3248 13812
rect 3178 13758 3187 13760
rect 3243 13758 3267 13760
rect 3323 13758 3332 13814
tri 3681 10504 3716 10539 se
rect 3716 10504 3768 14418
tri 3768 14390 3796 14418 nw
rect 22063 12010 22316 12180
rect 25200 11848 25252 11903
tri 26075 11705 26097 11727 se
rect 26097 11705 26149 11751
rect 3111 10502 3768 10504
rect 3111 10450 3117 10502
rect 3169 10450 3181 10502
rect 3233 10450 3768 10502
rect 3111 10447 3768 10450
tri 26055 11685 26075 11705 se
rect 26075 11685 26107 11705
rect 26055 10354 26107 11685
tri 26107 11663 26149 11705 nw
tri 26107 10354 26192 10439 sw
rect 26055 10311 26758 10354
tri 26055 10259 26107 10311 ne
rect 26107 10259 26758 10311
rect 3199 10253 3255 10259
rect 3199 10250 3200 10253
rect 3252 10250 3255 10253
tri 26107 10251 26115 10259 ne
rect 26115 10251 26758 10259
rect 3199 10189 3255 10194
rect 3199 10170 3200 10189
rect 3252 10170 3255 10189
rect 3199 10105 3255 10114
tri 3080 9942 3097 9959 sw
rect 3040 9941 3097 9942
tri 3040 9884 3097 9941 ne
tri 3097 9884 3155 9942 sw
tri 3097 9866 3115 9884 ne
tri 3092 9691 3115 9714 se
rect 3115 9691 3155 9884
tri 3080 9679 3092 9691 se
rect 3092 9679 3143 9691
tri 3143 9679 3155 9691 nw
tri 3040 9639 3080 9679 se
rect 3040 9316 3080 9639
tri 3080 9616 3143 9679 nw
tri 3040 9309 3047 9316 ne
rect 3047 9309 3080 9316
tri 3080 9309 3101 9330 sw
tri 3047 9276 3080 9309 ne
rect 3080 9276 3101 9309
tri 3080 9255 3101 9276 ne
tri 3101 9255 3155 9309 sw
tri 3101 9201 3155 9255 ne
tri 3155 9201 3209 9255 sw
tri 3155 9187 3169 9201 ne
tri 3010 9090 3086 9166 sw
rect 2958 9034 3086 9090
rect 3169 8055 3209 9201
tri 3209 8055 3230 8076 sw
rect 3169 8046 3234 8055
rect 3169 7990 3178 8046
rect 3169 7966 3234 7990
rect 3169 7910 3178 7966
rect 3169 7901 3234 7910
rect 26356 7497 26553 7498
rect 26356 7445 26362 7497
rect 26414 7445 26429 7497
rect 26481 7445 26495 7497
rect 26547 7445 26553 7497
rect 26356 7427 26553 7445
rect 26356 7375 26362 7427
rect 26414 7375 26429 7427
rect 26481 7375 26495 7427
rect 26547 7375 26553 7427
rect 26356 7357 26553 7375
rect 26356 7305 26362 7357
rect 26414 7305 26429 7357
rect 26481 7305 26495 7357
rect 26547 7305 26553 7357
rect 26356 6808 26553 7305
rect 26356 6756 26362 6808
rect 26414 6756 26429 6808
rect 26481 6756 26495 6808
rect 26547 6756 26553 6808
rect 26356 6738 26553 6756
rect 26356 6686 26362 6738
rect 26414 6686 26429 6738
rect 26481 6686 26495 6738
rect 26547 6686 26553 6738
rect 26356 6668 26553 6686
rect 26356 6616 26362 6668
rect 26414 6616 26429 6668
rect 26481 6616 26495 6668
rect 26547 6616 26553 6668
rect 26356 6615 26553 6616
rect 26616 6810 26758 10251
rect 26813 7501 27316 7502
rect 26813 7449 26819 7501
rect 26871 7449 26883 7501
rect 26935 7449 27316 7501
rect 26813 7431 27316 7449
rect 26813 7379 26819 7431
rect 26871 7379 26883 7431
rect 26935 7379 27316 7431
rect 26813 7361 27316 7379
rect 26813 7309 26819 7361
rect 26871 7309 26883 7361
rect 26935 7309 27316 7361
rect 26813 7308 27316 7309
tri 27117 7240 27185 7308 ne
tri 26758 6810 26812 6864 sw
rect 27185 6810 27316 7308
rect 26616 6809 26812 6810
tri 26812 6809 26813 6810 sw
rect 26616 6808 26813 6809
rect 26616 6756 26622 6808
rect 26674 6756 26689 6808
rect 26741 6756 26755 6808
rect 26807 6756 26813 6808
rect 26616 6738 26813 6756
rect 26616 6686 26622 6738
rect 26674 6686 26689 6738
rect 26741 6686 26755 6738
rect 26807 6686 26813 6738
rect 26616 6668 26813 6686
rect 26616 6616 26622 6668
rect 26674 6616 26689 6668
rect 26741 6616 26755 6668
rect 26807 6616 26813 6668
rect 27185 6758 27225 6810
rect 27277 6758 27316 6810
rect 27185 6740 27316 6758
rect 27185 6688 27225 6740
rect 27277 6688 27316 6740
rect 27185 6670 27316 6688
rect 27185 6618 27225 6670
rect 27277 6618 27316 6670
rect 27185 6617 27316 6618
rect 26616 6615 26813 6616
rect 26722 4969 27083 4977
rect 26774 4917 26816 4969
rect 26868 4917 27083 4969
rect 26722 4874 27083 4917
rect 26774 4822 26816 4874
rect 26868 4822 27083 4874
rect 26722 4463 27083 4822
rect 26774 4411 26816 4463
rect 26868 4411 27083 4463
rect 26722 4368 27083 4411
rect 26774 4316 26816 4368
rect 26868 4316 27083 4368
rect 26722 2926 27083 4316
rect 26494 2917 27083 2926
rect 26550 2861 26574 2917
rect 26630 2861 26654 2917
rect 26710 2861 26734 2917
rect 26790 2861 27083 2917
rect 26494 2828 27083 2861
rect 26550 2772 26574 2828
rect 26630 2772 26654 2828
rect 26710 2772 26734 2828
rect 26790 2772 27083 2828
rect 26494 2739 27083 2772
rect 26550 2683 26574 2739
rect 26630 2683 26654 2739
rect 26710 2683 26734 2739
rect 26790 2683 27083 2739
rect 26494 2650 27083 2683
rect 26550 2594 26574 2650
rect 26630 2594 26654 2650
rect 26710 2594 26734 2650
rect 26790 2594 27083 2650
rect 26494 2560 27083 2594
rect 26550 2504 26574 2560
rect 26630 2504 26654 2560
rect 26710 2504 26734 2560
rect 26790 2504 27083 2560
rect 26494 2495 27083 2504
rect 6870 2031 6876 2083
rect 6928 2050 6943 2083
rect 6995 2050 7010 2083
rect 7062 2050 7077 2083
rect 7129 2050 7144 2083
rect 7196 2050 7210 2083
rect 6936 2031 6943 2050
rect 7196 2031 7202 2050
rect 7262 2031 7268 2083
rect 6870 2015 6880 2031
rect 6936 2015 6961 2031
rect 7017 2015 7042 2031
rect 7098 2015 7122 2031
rect 7178 2015 7202 2031
rect 7258 2015 7268 2031
rect 6870 1963 6876 2015
rect 6936 1994 6943 2015
rect 7196 1994 7202 2015
rect 6928 1963 6943 1994
rect 6995 1963 7010 1994
rect 7062 1963 7077 1994
rect 7129 1963 7144 1994
rect 7196 1963 7210 1994
rect 7262 1963 7268 2015
rect 3281 1736 3337 1745
rect 3272 1658 3278 1710
rect 3337 1680 3342 1710
rect 3330 1658 3342 1680
rect 3394 1658 3400 1710
rect 3281 1656 3337 1658
rect 3281 1591 3337 1600
rect 12317 1397 12369 1403
rect 12317 1333 12369 1345
rect 12317 1275 12369 1281
rect 3055 957 3064 1013
rect 3124 961 3136 1013
rect 3120 957 3144 961
rect 3200 957 3209 1013
tri 9764 801 9816 853 se
rect 9816 817 12475 853
rect 9816 801 9838 817
tri 9838 801 9854 817 nw
rect 12469 801 12475 817
rect 12527 801 12539 853
rect 12591 801 12597 853
tri 9742 779 9764 801 se
rect 9764 779 9816 801
tri 9816 779 9838 801 nw
tri 9727 764 9742 779 se
rect 1629 708 1638 764
rect 1694 708 1718 764
rect 1774 708 3064 764
rect 3120 708 3144 764
rect 3200 708 3209 764
tri 9671 708 9727 764 se
rect 9727 708 9742 764
tri 9668 705 9671 708 se
rect 9671 705 9742 708
tri 9742 705 9816 779 nw
tri 9594 631 9668 705 se
tri 9668 631 9742 705 nw
tri 9526 563 9594 631 se
rect 9594 563 9600 631
tri 9600 563 9668 631 nw
rect 6312 511 9548 563
tri 9548 511 9600 563 nw
rect 3389 217 3398 273
rect 3454 217 3478 273
rect 3534 252 3543 273
rect 13277 252 13283 264
rect 3534 241 3565 252
tri 3565 241 3576 252 sw
tri 3954 241 3965 252 se
rect 3965 241 6651 252
tri 6651 241 6662 252 sw
tri 7446 241 7457 252 se
rect 7457 241 13283 252
rect 3534 226 3576 241
tri 3576 226 3591 241 sw
tri 3939 226 3954 241 se
rect 3954 226 6662 241
rect 3534 224 6662 226
tri 6662 224 6679 241 sw
rect 3534 217 6679 224
rect 3389 212 6679 217
tri 3536 189 3559 212 ne
rect 3559 189 3971 212
tri 3971 189 3994 212 nw
tri 6638 189 6661 212 ne
rect 6661 199 6679 212
tri 6679 199 6704 224 sw
rect 6661 189 6704 199
tri 6704 189 6714 199 sw
rect 6870 189 6876 241
rect 6928 209 6943 241
rect 6995 209 7010 241
rect 7062 209 7077 241
rect 7129 209 7144 241
rect 7196 209 7210 241
rect 6936 189 6943 209
rect 7196 189 7202 209
rect 7262 189 7268 241
tri 7417 212 7446 241 se
rect 7446 212 13283 241
rect 13335 212 13347 264
rect 13399 212 13405 264
tri 7404 199 7417 212 se
rect 7417 199 7457 212
tri 7457 199 7470 212 nw
tri 3559 186 3562 189 ne
rect 3562 186 3968 189
tri 3968 186 3971 189 nw
tri 6661 186 6664 189 ne
rect 6664 186 6714 189
tri 6664 173 6677 186 ne
rect 6677 173 6714 186
tri 6714 173 6730 189 sw
rect 6870 173 6880 189
rect 6936 173 6961 189
rect 7017 173 7042 189
rect 7098 173 7122 189
rect 7178 173 7202 189
rect 7258 173 7268 189
tri 6677 171 6679 173 ne
rect 6679 171 6730 173
tri 6730 171 6732 173 sw
tri 6679 121 6729 171 ne
rect 6729 146 6732 171
tri 6732 146 6757 171 sw
rect 6729 121 6757 146
tri 6757 121 6782 146 sw
rect 6870 121 6876 173
rect 6936 153 6943 173
rect 7196 153 7202 173
rect 6928 121 6943 153
rect 6995 121 7010 153
rect 7062 121 7077 153
rect 7129 121 7144 153
rect 7196 121 7210 153
rect 7262 121 7268 173
tri 7351 146 7404 199 se
tri 7404 146 7457 199 nw
tri 7326 121 7351 146 se
tri 6729 118 6732 121 ne
rect 6732 118 6782 121
tri 6782 118 6785 121 sw
tri 7323 118 7326 121 se
rect 7326 118 7351 121
tri 6732 65 6785 118 ne
tri 6785 93 6810 118 sw
tri 7298 93 7323 118 se
rect 7323 93 7351 118
tri 7351 93 7404 146 nw
rect 6785 65 6810 93
tri 6810 65 6838 93 sw
tri 7270 65 7298 93 se
rect 7298 65 7323 93
tri 7323 65 7351 93 nw
tri 6785 25 6825 65 ne
rect 6825 25 7283 65
tri 7283 25 7323 65 nw
<< via2 >>
rect 1674 14639 1730 14667
rect 1674 14611 1730 14639
rect 1674 14526 1730 14582
rect 3187 13812 3243 13814
rect 3267 13812 3323 13814
rect 3187 13760 3236 13812
rect 3236 13760 3243 13812
rect 3267 13760 3300 13812
rect 3300 13760 3323 13812
rect 3187 13758 3243 13760
rect 3267 13758 3323 13760
rect 3199 10201 3200 10250
rect 3200 10201 3252 10250
rect 3252 10201 3255 10250
rect 3199 10194 3255 10201
rect 3199 10137 3200 10170
rect 3200 10137 3252 10170
rect 3252 10137 3255 10170
rect 3199 10114 3255 10137
rect 3178 7990 3234 8046
rect 3178 7910 3234 7966
rect 26494 2861 26550 2917
rect 26574 2861 26630 2917
rect 26654 2861 26710 2917
rect 26734 2861 26790 2917
rect 26494 2772 26550 2828
rect 26574 2772 26630 2828
rect 26654 2772 26710 2828
rect 26734 2772 26790 2828
rect 26494 2683 26550 2739
rect 26574 2683 26630 2739
rect 26654 2683 26710 2739
rect 26734 2683 26790 2739
rect 26494 2594 26550 2650
rect 26574 2594 26630 2650
rect 26654 2594 26710 2650
rect 26734 2594 26790 2650
rect 26494 2504 26550 2560
rect 26574 2504 26630 2560
rect 26654 2504 26710 2560
rect 26734 2504 26790 2560
rect 6880 2031 6928 2050
rect 6928 2031 6936 2050
rect 6961 2031 6995 2050
rect 6995 2031 7010 2050
rect 7010 2031 7017 2050
rect 7042 2031 7062 2050
rect 7062 2031 7077 2050
rect 7077 2031 7098 2050
rect 7122 2031 7129 2050
rect 7129 2031 7144 2050
rect 7144 2031 7178 2050
rect 7202 2031 7210 2050
rect 7210 2031 7258 2050
rect 6880 2015 6936 2031
rect 6961 2015 7017 2031
rect 7042 2015 7098 2031
rect 7122 2015 7178 2031
rect 7202 2015 7258 2031
rect 6880 1994 6928 2015
rect 6928 1994 6936 2015
rect 6961 1994 6995 2015
rect 6995 1994 7010 2015
rect 7010 1994 7017 2015
rect 7042 1994 7062 2015
rect 7062 1994 7077 2015
rect 7077 1994 7098 2015
rect 7122 1994 7129 2015
rect 7129 1994 7144 2015
rect 7144 1994 7178 2015
rect 7202 1994 7210 2015
rect 7210 1994 7258 2015
rect 3281 1710 3337 1736
rect 3281 1680 3330 1710
rect 3330 1680 3337 1710
rect 3281 1600 3337 1656
rect 3064 961 3072 1013
rect 3072 961 3120 1013
rect 3144 961 3188 1013
rect 3188 961 3200 1013
rect 3064 957 3120 961
rect 3144 957 3200 961
rect 1638 708 1694 764
rect 1718 708 1774 764
rect 3064 708 3120 764
rect 3144 708 3200 764
rect 3398 217 3454 273
rect 3478 217 3534 273
rect 6880 189 6928 209
rect 6928 189 6936 209
rect 6961 189 6995 209
rect 6995 189 7010 209
rect 7010 189 7017 209
rect 7042 189 7062 209
rect 7062 189 7077 209
rect 7077 189 7098 209
rect 7122 189 7129 209
rect 7129 189 7144 209
rect 7144 189 7178 209
rect 7202 189 7210 209
rect 7210 189 7258 209
rect 6880 173 6936 189
rect 6961 173 7017 189
rect 7042 173 7098 189
rect 7122 173 7178 189
rect 7202 173 7258 189
rect 6880 153 6928 173
rect 6928 153 6936 173
rect 6961 153 6995 173
rect 6995 153 7010 173
rect 7010 153 7017 173
rect 7042 153 7062 173
rect 7062 153 7077 173
rect 7077 153 7098 173
rect 7122 153 7129 173
rect 7129 153 7144 173
rect 7144 153 7178 173
rect 7202 153 7210 173
rect 7210 153 7258 173
<< metal3 >>
rect 1633 14667 1771 14672
rect 1633 14611 1674 14667
rect 1730 14611 1771 14667
rect 1633 14582 1771 14611
rect 1633 14526 1674 14582
rect 1730 14526 1771 14582
rect 1633 769 1771 14526
rect 3182 13814 3328 13819
rect 3182 13758 3187 13814
rect 3243 13758 3267 13814
rect 3323 13758 3328 13814
rect 3182 13753 3328 13758
rect 3182 10250 3268 13753
tri 3268 13693 3328 13753 nw
rect 3182 10194 3199 10250
rect 3255 10194 3268 10250
rect 3182 10170 3268 10194
rect 3182 10114 3199 10170
rect 3255 10114 3268 10170
rect 3182 8372 3268 10114
tri 3182 8326 3228 8372 ne
rect 3228 8326 3268 8372
tri 3268 8326 3365 8423 sw
tri 3228 8286 3268 8326 ne
rect 3268 8286 3365 8326
tri 3268 8189 3365 8286 ne
tri 3365 8189 3502 8326 sw
tri 3365 8138 3416 8189 ne
rect 3173 8046 3247 8051
rect 3173 7990 3178 8046
rect 3234 7990 3247 8046
rect 3173 7966 3247 7990
rect 3173 7910 3178 7966
rect 3234 7910 3247 7966
rect 3173 7873 3247 7910
tri 3173 7806 3240 7873 ne
rect 3240 7806 3247 7873
tri 3247 7806 3354 7913 sw
tri 3240 7799 3247 7806 ne
rect 3247 7799 3354 7806
tri 3247 7778 3268 7799 ne
rect 3268 1736 3354 7799
rect 3268 1680 3281 1736
rect 3337 1680 3354 1736
rect 3268 1656 3354 1680
rect 3268 1600 3281 1656
rect 3337 1600 3354 1656
rect 3268 1543 3354 1600
rect 3059 1013 3205 1018
rect 3059 957 3064 1013
rect 3120 957 3144 1013
rect 3200 957 3205 1013
tri 1771 769 1779 777 sw
rect 1633 764 1779 769
rect 1633 708 1638 764
rect 1694 708 1718 764
rect 1774 708 1779 764
rect 1633 703 1779 708
rect 3059 764 3205 957
rect 3059 708 3064 764
rect 3120 708 3144 764
rect 3200 708 3205 764
rect 3059 703 3205 708
rect 3416 278 3502 8189
rect 26489 2917 26795 2922
rect 26489 2861 26494 2917
rect 26550 2861 26574 2917
rect 26630 2861 26654 2917
rect 26710 2861 26734 2917
rect 26790 2861 26795 2917
rect 26489 2828 26795 2861
rect 26489 2772 26494 2828
rect 26550 2772 26574 2828
rect 26630 2772 26654 2828
rect 26710 2772 26734 2828
rect 26790 2772 26795 2828
rect 26489 2739 26795 2772
rect 26489 2683 26494 2739
rect 26550 2683 26574 2739
rect 26630 2683 26654 2739
rect 26710 2683 26734 2739
rect 26790 2683 26795 2739
rect 26489 2650 26795 2683
rect 26489 2594 26494 2650
rect 26550 2594 26574 2650
rect 26630 2594 26654 2650
rect 26710 2594 26734 2650
rect 26790 2594 26795 2650
rect 26489 2560 26795 2594
rect 26489 2504 26494 2560
rect 26550 2504 26574 2560
rect 26630 2504 26654 2560
rect 26710 2504 26734 2560
rect 26790 2504 26795 2560
rect 26489 2499 26795 2504
rect 6875 2050 7263 2085
rect 6875 1994 6880 2050
rect 6936 1994 6961 2050
rect 7017 1994 7042 2050
rect 7098 1994 7122 2050
rect 7178 1994 7202 2050
rect 7258 1994 7263 2050
rect 3393 273 3539 278
rect 3393 217 3398 273
rect 3454 217 3478 273
rect 3534 217 3539 273
rect 3393 212 3539 217
rect 6875 209 7263 1994
rect 6875 153 6880 209
rect 6936 153 6961 209
rect 7017 153 7042 209
rect 7098 153 7122 209
rect 7178 153 7202 209
rect 7258 153 7263 209
rect 6875 118 7263 153
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1645210163
transform 1 0 12702 0 1 1750
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_1
timestamp 1645210163
transform 1 0 13054 0 1 1750
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1645210163
transform 1 0 12249 0 -1 2306
box -107 21 267 1369
use sky130_fd_io__sio_tk_em1s_cdns_55959141808166  sky130_fd_io__sio_tk_em1s_cdns_55959141808166_0
timestamp 1645210163
transform 1 0 13100 0 1 1744
box 0 24 144 28
use sky130_fd_io__gpio_ovtv2_hotswap_pghspu  sky130_fd_io__gpio_ovtv2_hotswap_pghspu_0
timestamp 1645210163
transform 1 0 2662 0 1 14350
box -126 0 23503 338
use sky130_fd_pr__pfet_01v8__example_55959141808160  sky130_fd_pr__pfet_01v8__example_55959141808160_0
timestamp 1645210163
transform -1 0 2493 0 -1 10921
box -28 0 228 267
use sky130_fd_io__tk_em1o_cdns_55959141808159  sky130_fd_io__tk_em1o_cdns_55959141808159_0
timestamp 1645210163
transform -1 0 2765 0 1 10640
box 0 24 168 28
use sky130_fd_io__gpio_ovtv2_hotswap_guardrings  sky130_fd_io__gpio_ovtv2_hotswap_guardrings_0
timestamp 1645210163
transform 1 0 482 0 1 7158
box 0 0 26980 8664
use sky130_fd_io__signal_5_sym_hv_local_5term  sky130_fd_io__signal_5_sym_hv_local_5term_0
timestamp 1645210163
transform -1 0 27387 0 -1 6877
box 0 0 1591 2424
use sky130_fd_io__gpio_ovtv2_hvsbt_inv_x4  sky130_fd_io__gpio_ovtv2_hvsbt_inv_x4_0
timestamp 1645210163
transform 1 0 12543 0 -1 2307
box -107 21 795 1369
use sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix  sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix_0
timestamp 1645210163
transform 1 0 -2122 0 1 -535
box 2296 657 28371 15193
<< labels >>
flabel metal3 s 1633 14544 1771 14632 3 FreeSans 520 0 0 0 PAD
port 1 nsew
flabel metal2 s 22063 12010 22316 12180 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew
flabel metal2 s 26722 4226 27083 4289 3 FreeSans 520 0 0 0 VSSD
port 3 nsew
flabel metal2 s 3278 10449 3337 10503 3 FreeSans 520 0 0 0 PGHS_H
port 4 nsew
flabel metal2 s 25200 11848 25252 11903 3 FreeSans 520 0 0 0 P3OUT
port 5 nsew
flabel locali s 792 7224 1045 7394 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew
flabel locali s 1713 8686 1943 8857 3 FreeSans 520 0 0 0 VPB_DRVR
port 6 nsew
flabel comment s 3450 7594 3450 7594 0 FreeSans 800 90 0 0 PADLO
flabel comment s 3467 1036 3467 1036 0 FreeSans 400 0 0 0 PADLO
flabel metal1 s 13252 1744 13356 1862 3 FreeSans 520 0 0 0 PADLO
port 7 nsew
flabel metal1 s 12785 1462 13038 1632 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew
flabel metal1 s 10816 962 10888 1014 3 FreeSans 520 0 0 0 EN_H
port 8 nsew
flabel metal1 s 10526 944 10611 982 3 FreeSans 520 0 0 0 FORCE_H[1]
port 9 nsew
flabel metal1 s 11943 880 12003 912 3 FreeSans 200 0 0 0 OD_H
port 10 nsew
flabel metal1 s 7753 749 7852 795 3 FreeSans 520 0 0 0 VPWR_KA
port 11 nsew
flabel metal1 s 25669 14501 25704 14541 3 FreeSans 200 0 0 0 VCC_IO_SOFT
port 12 nsew
flabel metal1 s 6192 14499 6267 14545 3 FreeSans 200 0 0 0 TIE_HI
port 13 nsew
flabel metal1 s 1117 7749 1478 7812 3 FreeSans 520 0 0 0 VSSD
port 3 nsew
flabel metal1 s 6441 2052 6802 2115 3 FreeSans 520 0 0 0 VSSD
port 3 nsew
flabel metal1 s 2664 300 2917 470 3 FreeSans 520 0 0 0 VDDIO
port 2 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 40235080
string GDS_START 40211114
<< end >>
