magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 21 21 643 203
rect 29 -17 63 21
<< scnmos >>
rect 99 47 129 177
rect 171 47 201 177
rect 255 47 285 177
rect 443 47 473 177
rect 527 47 557 177
<< scpmoshvt >>
rect 87 297 117 497
rect 171 297 201 497
rect 347 297 377 497
rect 419 297 449 497
rect 515 297 545 497
<< ndiff >>
rect 47 163 99 177
rect 47 129 55 163
rect 89 129 99 163
rect 47 95 99 129
rect 47 61 55 95
rect 89 61 99 95
rect 47 47 99 61
rect 129 47 171 177
rect 201 163 255 177
rect 201 129 211 163
rect 245 129 255 163
rect 201 95 255 129
rect 201 61 211 95
rect 245 61 255 95
rect 201 47 255 61
rect 285 163 337 177
rect 285 129 295 163
rect 329 129 337 163
rect 285 95 337 129
rect 285 61 295 95
rect 329 61 337 95
rect 285 47 337 61
rect 391 95 443 177
rect 391 61 399 95
rect 433 61 443 95
rect 391 47 443 61
rect 473 128 527 177
rect 473 94 483 128
rect 517 94 527 128
rect 473 47 527 94
rect 557 128 617 177
rect 557 94 575 128
rect 609 94 617 128
rect 557 47 617 94
<< pdiff >>
rect 27 485 87 497
rect 27 451 43 485
rect 77 451 87 485
rect 27 297 87 451
rect 117 477 171 497
rect 117 443 127 477
rect 161 443 171 477
rect 117 409 171 443
rect 117 375 127 409
rect 161 375 171 409
rect 117 297 171 375
rect 201 475 347 497
rect 201 441 211 475
rect 245 441 303 475
rect 337 441 347 475
rect 201 297 347 441
rect 377 297 419 497
rect 449 459 515 497
rect 449 425 471 459
rect 505 425 515 459
rect 449 297 515 425
rect 545 475 617 497
rect 545 441 563 475
rect 597 441 617 475
rect 545 297 617 441
<< ndiffc >>
rect 55 129 89 163
rect 55 61 89 95
rect 211 129 245 163
rect 211 61 245 95
rect 295 129 329 163
rect 295 61 329 95
rect 399 61 433 95
rect 483 94 517 128
rect 575 94 609 128
<< pdiffc >>
rect 43 451 77 485
rect 127 443 161 477
rect 127 375 161 409
rect 211 441 245 475
rect 303 441 337 475
rect 471 425 505 459
rect 563 441 597 475
<< poly >>
rect 87 497 117 523
rect 171 497 201 523
rect 347 497 377 523
rect 419 497 449 523
rect 515 497 545 523
rect 87 265 117 297
rect 171 265 201 297
rect 347 265 377 297
rect 75 249 129 265
rect 75 215 85 249
rect 119 215 129 249
rect 75 199 129 215
rect 99 177 129 199
rect 171 249 377 265
rect 171 215 202 249
rect 236 215 270 249
rect 304 215 377 249
rect 171 199 377 215
rect 419 265 449 297
rect 515 265 545 297
rect 419 249 473 265
rect 419 215 429 249
rect 463 215 473 249
rect 419 199 473 215
rect 515 249 569 265
rect 515 215 525 249
rect 559 215 569 249
rect 515 199 569 215
rect 171 177 201 199
rect 255 177 285 199
rect 443 177 473 199
rect 527 177 557 199
rect 99 21 129 47
rect 171 21 201 47
rect 255 21 285 47
rect 443 21 473 47
rect 527 21 557 47
<< polycont >>
rect 85 215 119 249
rect 202 215 236 249
rect 270 215 304 249
rect 429 215 463 249
rect 525 215 559 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 485 77 527
rect 17 451 43 485
rect 17 425 77 451
rect 111 477 177 493
rect 111 443 127 477
rect 161 443 177 477
rect 111 409 177 443
rect 211 475 337 527
rect 245 441 303 475
rect 563 475 623 527
rect 211 425 337 441
rect 453 425 471 459
rect 505 425 529 459
rect 597 441 623 475
rect 563 425 623 441
rect 111 391 127 409
rect 17 375 127 391
rect 161 391 177 409
rect 495 391 529 425
rect 161 375 461 391
rect 17 357 461 375
rect 17 165 51 357
rect 85 289 393 323
rect 85 249 134 289
rect 119 215 134 249
rect 186 249 325 255
rect 186 215 202 249
rect 236 215 270 249
rect 304 215 325 249
rect 359 249 393 289
rect 427 317 461 357
rect 495 351 627 391
rect 427 283 559 317
rect 525 249 559 283
rect 359 215 429 249
rect 463 215 479 249
rect 85 199 134 215
rect 525 199 559 215
rect 17 163 110 165
rect 17 129 55 163
rect 89 129 110 163
rect 17 95 110 129
rect 17 61 55 95
rect 89 61 110 95
rect 17 56 110 61
rect 211 163 245 181
rect 211 95 245 129
rect 211 17 245 61
rect 279 165 461 181
rect 593 165 627 351
rect 279 163 529 165
rect 279 129 295 163
rect 329 147 529 163
rect 329 129 345 147
rect 427 131 529 147
rect 279 95 345 129
rect 483 128 529 131
rect 279 61 295 95
rect 329 61 345 95
rect 279 51 345 61
rect 379 61 399 95
rect 433 61 449 95
rect 379 17 449 61
rect 517 94 529 128
rect 483 51 529 94
rect 563 128 627 165
rect 563 94 575 128
rect 609 94 627 128
rect 563 69 627 94
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 121 289 155 323 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 581 357 615 391 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 xnor2_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 505594
string GDS_START 500290
string path 0.000 2.720 3.220 2.720 
<< end >>
