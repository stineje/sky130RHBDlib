// File: and2x1_pcell.spi.pex
// Created: Tue Oct 15 15:54:20 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_AND2X1_PCELL\%noxref_1 ( 11 15 18 23 31 34 39 43 54 58 70 71 )
c78 ( 71 0 ) capacitor c=0.0600324f //x=3.825 //y=0.37
c79 ( 70 0 ) capacitor c=0.0208404f //x=0.99 //y=0.865
c80 ( 58 0 ) capacitor c=0.10149f //x=3.33 //y=0
c81 ( 57 0 ) capacitor c=0.00440095f //x=1.18 //y=0
c82 ( 54 0 ) capacitor c=0.198211f //x=5.18 //y=0
c83 ( 52 0 ) capacitor c=0.0360689f //x=5.015 //y=0
c84 ( 46 0 ) capacitor c=0.00583665f //x=4.93 //y=0.45
c85 ( 43 0 ) capacitor c=0.00542558f //x=4.845 //y=0.535
c86 ( 42 0 ) capacitor c=0.00479856f //x=4.445 //y=0.45
c87 ( 39 0 ) capacitor c=0.0068422f //x=4.36 //y=0.535
c88 ( 34 0 ) capacitor c=0.00588377f //x=3.96 //y=0.45
c89 ( 31 0 ) capacitor c=0.0164879f //x=3.875 //y=0
c90 ( 23 0 ) capacitor c=0.0720403f //x=3.16 //y=0
c91 ( 18 0 ) capacitor c=0.179504f //x=0.74 //y=0
c92 ( 15 0 ) capacitor c=0.0426751f //x=1.095 //y=0
c93 ( 11 0 ) capacitor c=0.221897f //x=5.18 //y=0
r94 (  62 63 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.445 //y=0 //x2=4.93 //y2=0
r95 (  61 62 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=4.44 //y=0 //x2=4.445 //y2=0
r96 (  59 61 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=3.96 //y=0 //x2=4.44 //y2=0
r97 (  52 63 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.015 //y=0 //x2=4.93 //y2=0
r98 (  52 54 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=5.015 //y=0 //x2=5.18 //y2=0
r99 (  47 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=4.93 //y=0.62 //x2=4.93 //y2=0.535
r100 (  47 71 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.62 //x2=4.93 //y2=1.225
r101 (  46 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.45 //x2=4.93 //y2=0.535
r102 (  45 63 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.17 //x2=4.93 //y2=0
r103 (  45 46 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.17 //x2=4.93 //y2=0.45
r104 (  44 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.53 //y=0.535 //x2=4.445 //y2=0.535
r105 (  43 71 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.845 //y=0.535 //x2=4.93 //y2=0.535
r106 (  43 44 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.845 //y=0.535 //x2=4.53 //y2=0.535
r107 (  42 71 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.45 //x2=4.445 //y2=0.535
r108 (  41 62 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.17 //x2=4.445 //y2=0
r109 (  41 42 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.17 //x2=4.445 //y2=0.45
r110 (  40 71 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.045 //y=0.535 //x2=3.96 //y2=0.535
r111 (  39 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.36 //y=0.535 //x2=4.445 //y2=0.535
r112 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.36 //y=0.535 //x2=4.045 //y2=0.535
r113 (  35 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.62 //x2=3.96 //y2=0.535
r114 (  35 71 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.62 //x2=3.96 //y2=1.225
r115 (  34 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.45 //x2=3.96 //y2=0.535
r116 (  33 59 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.17 //x2=3.96 //y2=0
r117 (  33 34 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.17 //x2=3.96 //y2=0.45
r118 (  32 58 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.5 //y=0 //x2=3.33 //y2=0
r119 (  31 59 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.875 //y=0 //x2=3.96 //y2=0
r120 (  31 32 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=3.875 //y=0 //x2=3.5 //y2=0
r121 (  26 28 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r122 (  24 57 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.18 //y2=0
r123 (  24 26 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.85 //y2=0
r124 (  23 58 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.16 //y=0 //x2=3.33 //y2=0
r125 (  23 28 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r126 (  19 57 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r127 (  19 70 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.955
r128 (  15 57 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=1.18 //y2=0
r129 (  15 18 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=0.74 //y2=0
r130 (  11 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.18 //y=0 //x2=5.18 //y2=0
r131 (  9 61 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r132 (  9 11 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.18 //y2=0
r133 (  7 28 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r134 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r135 (  5 26 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r136 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r137 (  2 18 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r138 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_AND2X1_PCELL\%noxref_1

subckt PM_AND2X1_PCELL\%noxref_2 ( 11 23 31 55 68 72 75 78 79 80 81 82 )
c70 ( 82 0 ) capacitor c=0.0451925f //x=4.74 //y=5.02
c71 ( 81 0 ) capacitor c=0.042362f //x=3.87 //y=5.02
c72 ( 80 0 ) capacitor c=0.0382536f //x=2.405 //y=5.02
c73 ( 79 0 ) capacitor c=0.0243052f //x=1.525 //y=5.02
c74 ( 78 0 ) capacitor c=0.053196f //x=0.655 //y=5.02
c75 ( 77 0 ) capacitor c=0.00591168f //x=4.885 //y=7.4
c76 ( 76 0 ) capacitor c=0.00591168f //x=4.005 //y=7.4
c77 ( 75 0 ) capacitor c=0.110791f //x=3.33 //y=7.4
c78 ( 74 0 ) capacitor c=0.00591168f //x=2.55 //y=7.4
c79 ( 73 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c80 ( 72 0 ) capacitor c=0.24846f //x=0.74 //y=7.4
c81 ( 68 0 ) capacitor c=0.228884f //x=5.18 //y=7.4
c82 ( 55 0 ) capacitor c=0.0287207f //x=4.8 //y=7.4
c83 ( 47 0 ) capacitor c=0.0216067f //x=3.92 //y=7.4
c84 ( 41 0 ) capacitor c=0.0275781f //x=3.16 //y=7.4
c85 ( 31 0 ) capacitor c=0.0285035f //x=2.465 //y=7.4
c86 ( 23 0 ) capacitor c=0.0286367f //x=1.585 //y=7.4
c87 ( 11 0 ) capacitor c=0.232079f //x=5.18 //y=7.4
r88 (  66 77 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.97 //y=7.4 //x2=4.885 //y2=7.4
r89 (  66 68 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=4.97 //y=7.4 //x2=5.18 //y2=7.4
r90 (  59 77 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.885 //y=7.23 //x2=4.885 //y2=7.4
r91 (  59 82 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.885 //y=7.23 //x2=4.885 //y2=6.405
r92 (  56 76 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.09 //y=7.4 //x2=4.005 //y2=7.4
r93 (  56 58 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li //thickness=0.1 \
 //x=4.09 //y=7.4 //x2=4.44 //y2=7.4
r94 (  55 77 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.8 //y=7.4 //x2=4.885 //y2=7.4
r95 (  55 58 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=4.8 //y=7.4 //x2=4.44 //y2=7.4
r96 (  49 76 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.005 //y=7.23 //x2=4.005 //y2=7.4
r97 (  49 81 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.005 //y=7.23 //x2=4.005 //y2=6.405
r98 (  48 75 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r99 (  47 76 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.92 //y=7.4 //x2=4.005 //y2=7.4
r100 (  47 48 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=3.92 //y=7.4 //x2=3.5 //y2=7.4
r101 (  42 74 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.55 //y2=7.4
r102 (  42 44 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.96 //y2=7.4
r103 (  41 75 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r104 (  41 44 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r105 (  35 74 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r106 (  35 80 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.745
r107 (  32 73 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r108 (  32 34 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r109 (  31 74 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r110 (  31 34 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r111 (  25 73 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r112 (  25 79 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.745
r113 (  24 72 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r114 (  23 73 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r115 (  23 24 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r116 (  17 72 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r117 (  17 78 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.405
r118 (  11 68 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.18 //y=7.4 //x2=5.18 //y2=7.4
r119 (  9 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r120 (  9 11 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.18 //y2=7.4
r121 (  7 44 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r122 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r123 (  5 34 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r124 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r125 (  2 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r126 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_AND2X1_PCELL\%noxref_2

subckt PM_AND2X1_PCELL\%noxref_3 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 52 53 54 56 62 63 65 73 75 76 )
c132 ( 76 0 ) capacitor c=0.0220291f //x=1.965 //y=5.02
c133 ( 75 0 ) capacitor c=0.0217503f //x=1.085 //y=5.02
c134 ( 73 0 ) capacitor c=0.0084702f //x=1.96 //y=0.905
c135 ( 65 0 ) capacitor c=0.0528806f //x=4.07 //y=2.085
c136 ( 63 0 ) capacitor c=0.0435629f //x=4.71 //y=1.255
c137 ( 62 0 ) capacitor c=0.0200386f //x=4.71 //y=0.91
c138 ( 56 0 ) capacitor c=0.0152946f //x=4.555 //y=1.41
c139 ( 54 0 ) capacitor c=0.0157804f //x=4.555 //y=0.755
c140 ( 53 0 ) capacitor c=0.0524991f //x=4.3 //y=4.79
c141 ( 52 0 ) capacitor c=0.0322983f //x=4.59 //y=4.79
c142 ( 48 0 ) capacitor c=0.0290017f //x=4.18 //y=1.92
c143 ( 47 0 ) capacitor c=0.0250027f //x=4.18 //y=1.565
c144 ( 46 0 ) capacitor c=0.0234316f //x=4.18 //y=1.255
c145 ( 45 0 ) capacitor c=0.0200596f //x=4.18 //y=0.91
c146 ( 44 0 ) capacitor c=0.154218f //x=4.665 //y=6.02
c147 ( 43 0 ) capacitor c=0.154243f //x=4.225 //y=6.02
c148 ( 41 0 ) capacitor c=0.00427536f //x=2.11 //y=5.2
c149 ( 34 0 ) capacitor c=0.0944546f //x=4.07 //y=2.085
c150 ( 32 0 ) capacitor c=0.112578f //x=2.59 //y=3.33
c151 ( 28 0 ) capacitor c=0.00781917f //x=2.235 //y=1.655
c152 ( 27 0 ) capacitor c=0.0161074f //x=2.505 //y=1.655
c153 ( 25 0 ) capacitor c=0.0158072f //x=2.505 //y=5.2
c154 ( 14 0 ) capacitor c=0.00387264f //x=1.315 //y=5.2
c155 ( 13 0 ) capacitor c=0.0209922f //x=2.025 //y=5.2
c156 ( 2 0 ) capacitor c=0.0157298f //x=2.705 //y=3.33
c157 ( 1 0 ) capacitor c=0.0800687f //x=3.955 //y=3.33
r158 (  65 66 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.07 //y=2.085 //x2=4.18 //y2=2.085
r159 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.71 //y=1.255 //x2=4.67 //y2=1.41
r160 (  62 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.71 //y=0.91 //x2=4.67 //y2=0.755
r161 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.71 //y=0.91 //x2=4.71 //y2=1.255
r162 (  57 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.335 //y=1.41 //x2=4.22 //y2=1.41
r163 (  56 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.555 //y=1.41 //x2=4.67 //y2=1.41
r164 (  55 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.335 //y=0.755 //x2=4.22 //y2=0.755
r165 (  54 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.555 //y=0.755 //x2=4.67 //y2=0.755
r166 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.555 //y=0.755 //x2=4.335 //y2=0.755
r167 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.59 //y=4.79 //x2=4.665 //y2=4.865
r168 (  52 53 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=4.59 //y=4.79 //x2=4.3 //y2=4.79
r169 (  49 53 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.225 //y=4.865 //x2=4.3 //y2=4.79
r170 (  49 68 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=4.225 //y=4.865 //x2=4.07 //y2=4.7
r171 (  48 66 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.92 //x2=4.18 //y2=2.085
r172 (  47 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.565 //x2=4.22 //y2=1.41
r173 (  47 48 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.565 //x2=4.18 //y2=1.92
r174 (  46 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.255 //x2=4.22 //y2=1.41
r175 (  45 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=0.91 //x2=4.22 //y2=0.755
r176 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.18 //y=0.91 //x2=4.18 //y2=1.255
r177 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.665 //y=6.02 //x2=4.665 //y2=4.865
r178 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.225 //y=6.02 //x2=4.225 //y2=4.865
r179 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.445 //y=1.41 //x2=4.555 //y2=1.41
r180 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.445 //y=1.41 //x2=4.335 //y2=1.41
r181 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=4.7 //x2=4.07 //y2=4.7
r182 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=3.33 //x2=4.07 //y2=4.7
r183 (  34 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=2.085 //x2=4.07 //y2=2.085
r184 (  34 37 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=4.07 //y=2.085 //x2=4.07 //y2=3.33
r185 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.115 //x2=2.59 //y2=3.33
r186 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=3.33
r187 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r188 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r189 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.195 //y=5.2 //x2=2.11 //y2=5.2
r190 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.59 //y2=5.115
r191 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.195 //y2=5.2
r192 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.235 //y2=1.655
r193 (  21 73 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r194 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.2
r195 (  15 76 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.725
r196 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=2.11 //y2=5.2
r197 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=1.315 //y2=5.2
r198 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.315 //y2=5.2
r199 (  7 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.23 //y2=5.725
r200 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.33 //x2=4.07 //y2=3.33
r201 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=3.33 //x2=2.59 //y2=3.33
r202 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=3.33 //x2=2.59 //y2=3.33
r203 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.955 //y=3.33 //x2=4.07 //y2=3.33
r204 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=3.955 //y=3.33 //x2=2.705 //y2=3.33
ends PM_AND2X1_PCELL\%noxref_3

subckt PM_AND2X1_PCELL\%noxref_4 ( 2 7 8 9 10 11 12 13 17 19 22 23 33 )
c56 ( 33 0 ) capacitor c=0.0667949f //x=1.11 //y=4.7
c57 ( 23 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c58 ( 22 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c59 ( 19 0 ) capacitor c=0.0141798f //x=1.29 //y=1.365
c60 ( 17 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c61 ( 13 0 ) capacitor c=0.0860049f //x=0.915 //y=1.915
c62 ( 12 0 ) capacitor c=0.0229722f //x=0.915 //y=1.52
c63 ( 11 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c64 ( 10 0 ) capacitor c=0.0199343f //x=0.915 //y=0.865
c65 ( 9 0 ) capacitor c=0.110275f //x=1.45 //y=6.02
c66 ( 8 0 ) capacitor c=0.154305f //x=1.01 //y=6.02
c67 ( 2 0 ) capacitor c=0.116498f //x=1.11 //y=2.08
r68 (  31 33 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.7 //x2=1.11 //y2=4.7
r69 (  24 33 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=1.45 //y=4.865 //x2=1.11 //y2=4.7
r70 (  23 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r71 (  22 34 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r72 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r73 (  20 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r74 (  19 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r75 (  18 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r76 (  17 34 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r77 (  17 18 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r78 (  14 31 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.865 //x2=1.01 //y2=4.7
r79 (  13 28 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r80 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r81 (  12 13 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r82 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r83 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r84 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r85 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.02 //x2=1.45 //y2=4.865
r86 (  8 14 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.02 //x2=1.01 //y2=4.865
r87 (  7 19 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r88 (  7 20 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r89 (  5 33 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r90 (  2 28 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r91 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=4.7
ends PM_AND2X1_PCELL\%noxref_4

subckt PM_AND2X1_PCELL\%noxref_5 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c64 ( 34 0 ) capacitor c=0.034715f //x=1.88 //y=4.7
c65 ( 31 0 ) capacitor c=0.0279499f //x=1.85 //y=1.915
c66 ( 30 0 ) capacitor c=0.0437302f //x=1.85 //y=2.08
c67 ( 28 0 ) capacitor c=0.0429696f //x=2.415 //y=1.25
c68 ( 27 0 ) capacitor c=0.0192208f //x=2.415 //y=0.905
c69 ( 21 0 ) capacitor c=0.0158629f //x=2.26 //y=1.405
c70 ( 19 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c71 ( 17 0 ) capacitor c=0.0367015f //x=2.255 //y=4.79
c72 ( 12 0 ) capacitor c=0.0205163f //x=1.885 //y=1.56
c73 ( 11 0 ) capacitor c=0.0168481f //x=1.885 //y=1.25
c74 ( 10 0 ) capacitor c=0.0174783f //x=1.885 //y=0.905
c75 ( 9 0 ) capacitor c=0.15358f //x=2.33 //y=6.02
c76 ( 8 0 ) capacitor c=0.110281f //x=1.89 //y=6.02
c77 ( 3 0 ) capacitor c=0.0813556f //x=1.85 //y=2.08
c78 ( 1 0 ) capacitor c=0.00453889f //x=1.85 //y=4.535
r79 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.79 //x2=1.88 //y2=4.865
r80 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.7 //x2=1.88 //y2=4.79
r81 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r82 (  28 41 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r83 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r84 (  27 28 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r85 (  22 39 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r86 (  21 41 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r87 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r88 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r89 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r90 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.015 //y=4.79 //x2=1.88 //y2=4.79
r91 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.33 //y2=4.865
r92 (  17 18 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.015 //y2=4.79
r93 (  12 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r94 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r95 (  11 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r96 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r97 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r98 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.02 //x2=2.33 //y2=4.865
r99 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.02 //x2=1.89 //y2=4.865
r100 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r101 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r102 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.88 //y=4.7 //x2=1.88 //y2=4.7
r103 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r104 (  1 6 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.865 //y2=4.7
r105 (  1 3 ) resistor r=168.043 //w=0.187 //l=2.455 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.85 //y2=2.08
ends PM_AND2X1_PCELL\%noxref_5

subckt PM_AND2X1_PCELL\%noxref_6 ( 1 5 9 10 13 17 29 )
c50 ( 29 0 ) capacitor c=0.0633719f //x=0.56 //y=0.365
c51 ( 17 0 ) capacitor c=0.00722223f //x=2.635 //y=0.615
c52 ( 13 0 ) capacitor c=0.0154437f //x=2.55 //y=0.53
c53 ( 10 0 ) capacitor c=0.0092508f //x=1.665 //y=1.495
c54 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c55 ( 5 0 ) capacitor c=0.0255599f //x=1.58 //y=1.58
c56 ( 1 0 ) capacitor c=0.0113547f //x=0.695 //y=1.495
r57 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r58 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r59 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r60 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=2.15 //y2=0.53
r61 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r62 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.15 //y2=0.53
r63 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r64 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r65 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r66 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r67 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r68 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r69 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r70 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r71 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r72 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_AND2X1_PCELL\%noxref_6

subckt PM_AND2X1_PCELL\%noxref_7 ( 11 12 13 14 16 17 19 )
c44 ( 19 0 ) capacitor c=0.028734f //x=4.3 //y=5.02
c45 ( 17 0 ) capacitor c=0.0173218f //x=4.255 //y=0.91
c46 ( 16 0 ) capacitor c=0.105613f //x=4.81 //y=4.495
c47 ( 14 0 ) capacitor c=0.00575887f //x=4.53 //y=4.58
c48 ( 13 0 ) capacitor c=0.0136889f //x=4.725 //y=4.58
c49 ( 12 0 ) capacitor c=0.00636159f //x=4.525 //y=2.08
c50 ( 11 0 ) capacitor c=0.0140707f //x=4.725 //y=2.08
r51 (  15 16 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=4.81 //y=2.165 //x2=4.81 //y2=4.495
r52 (  13 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=4.58 //x2=4.81 //y2=4.495
r53 (  13 14 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=4.725 //y=4.58 //x2=4.53 //y2=4.58
r54 (  11 15 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=2.08 //x2=4.81 //y2=2.165
r55 (  11 12 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=4.725 //y=2.08 //x2=4.525 //y2=2.08
r56 (  5 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.445 //y=4.665 //x2=4.53 //y2=4.58
r57 (  5 19 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li //thickness=0.1 \
 //x=4.445 //y=4.665 //x2=4.445 //y2=5.725
r58 (  1 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.44 //y=1.995 //x2=4.525 //y2=2.08
r59 (  1 17 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=4.44 //y=1.995 //x2=4.44 //y2=1.005
ends PM_AND2X1_PCELL\%noxref_7

