// File: AO3X1.spi.pex
// Created: Tue Oct 15 15:44:44 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_AO3X1\%GND ( 1 16 20 23 28 39 44 48 56 60 82 86 99 119 124 131 132 \
 133 )
c122 ( 133 0 ) capacitor c=0.0597349f //x=7.155 //y=0.37
c123 ( 132 0 ) capacitor c=0.0696742f //x=3.89 //y=0.365
c124 ( 131 0 ) capacitor c=0.0208404f //x=0.99 //y=0.865
c125 ( 124 0 ) capacitor c=0.233789f //x=8.26 //y=0
c126 ( 119 0 ) capacitor c=0.0990091f //x=6.66 //y=0
c127 ( 99 0 ) capacitor c=0.107062f //x=3.33 //y=0
c128 ( 98 0 ) capacitor c=0.00440095f //x=1.18 //y=0
c129 ( 89 0 ) capacitor c=0.00587411f //x=8.26 //y=0.45
c130 ( 86 0 ) capacitor c=0.00542558f //x=8.175 //y=0.535
c131 ( 85 0 ) capacitor c=0.00479856f //x=7.775 //y=0.45
c132 ( 82 0 ) capacitor c=0.00690112f //x=7.69 //y=0.535
c133 ( 77 0 ) capacitor c=0.00592191f //x=7.29 //y=0.45
c134 ( 72 0 ) capacitor c=0.0190475f //x=7.205 //y=0
c135 ( 69 0 ) capacitor c=0.0659312f //x=6.05 //y=0
c136 ( 68 0 ) capacitor c=0.0227441f //x=6.49 //y=0
c137 ( 63 0 ) capacitor c=0.00609805f //x=5.965 //y=0.445
c138 ( 60 0 ) capacitor c=0.00508073f //x=5.88 //y=0.53
c139 ( 59 0 ) capacitor c=0.00468234f //x=5.48 //y=0.445
c140 ( 56 0 ) capacitor c=0.00556167f //x=5.395 //y=0.53
c141 ( 51 0 ) capacitor c=0.00468234f //x=4.995 //y=0.445
c142 ( 48 0 ) capacitor c=0.00556167f //x=4.91 //y=0.53
c143 ( 47 0 ) capacitor c=0.00468234f //x=4.51 //y=0.445
c144 ( 44 0 ) capacitor c=0.00692577f //x=4.425 //y=0.53
c145 ( 39 0 ) capacitor c=0.00609805f //x=4.025 //y=0.445
c146 ( 36 0 ) capacitor c=0.0227441f //x=3.94 //y=0
c147 ( 28 0 ) capacitor c=0.0751168f //x=3.16 //y=0
c148 ( 23 0 ) capacitor c=0.179504f //x=0.74 //y=0
c149 ( 20 0 ) capacitor c=0.0426751f //x=1.095 //y=0
c150 ( 16 0 ) capacitor c=0.343897f //x=8.14 //y=0
r151 (  123 124 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=8.14 //y=0 //x2=8.26 //y2=0
r152 (  121 123 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=7.775 //y=0 //x2=8.14 //y2=0
r153 (  120 121 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.29 //y=0 //x2=7.775 //y2=0
r154 (  107 108 ) resistor r=14.8796 //w=0.357 //l=0.415 //layer=li \
 //thickness=0.1 //x=5.55 //y=0 //x2=5.965 //y2=0
r155 (  105 107 ) resistor r=2.5098 //w=0.357 //l=0.07 //layer=li \
 //thickness=0.1 //x=5.48 //y=0 //x2=5.55 //y2=0
r156 (  104 105 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.995 //y=0 //x2=5.48 //y2=0
r157 (  103 104 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.51 //y=0 //x2=4.995 //y2=0
r158 (  102 103 ) resistor r=2.5098 //w=0.357 //l=0.07 //layer=li \
 //thickness=0.1 //x=4.44 //y=0 //x2=4.51 //y2=0
r159 (  100 102 ) resistor r=14.8796 //w=0.357 //l=0.415 //layer=li \
 //thickness=0.1 //x=4.025 //y=0 //x2=4.44 //y2=0
r160 (  90 133 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.26 //y=0.62 //x2=8.26 //y2=0.535
r161 (  90 133 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=8.26 //y=0.62 //x2=8.26 //y2=1.225
r162 (  89 133 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.26 //y=0.45 //x2=8.26 //y2=0.535
r163 (  88 124 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.26 //y=0.17 //x2=8.26 //y2=0
r164 (  88 89 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=8.26 //y=0.17 //x2=8.26 //y2=0.45
r165 (  87 133 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.86 //y=0.535 //x2=7.775 //y2=0.535
r166 (  86 133 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.175 //y=0.535 //x2=8.26 //y2=0.535
r167 (  86 87 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=8.175 //y=0.535 //x2=7.86 //y2=0.535
r168 (  85 133 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.775 //y=0.45 //x2=7.775 //y2=0.535
r169 (  84 121 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.775 //y=0.17 //x2=7.775 //y2=0
r170 (  84 85 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=7.775 //y=0.17 //x2=7.775 //y2=0.45
r171 (  83 133 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.375 //y=0.535 //x2=7.29 //y2=0.535
r172 (  82 133 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.69 //y=0.535 //x2=7.775 //y2=0.535
r173 (  82 83 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=7.69 //y=0.535 //x2=7.375 //y2=0.535
r174 (  78 133 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.29 //y=0.62 //x2=7.29 //y2=0.535
r175 (  78 133 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=7.29 //y=0.62 //x2=7.29 //y2=1.225
r176 (  77 133 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.29 //y=0.45 //x2=7.29 //y2=0.535
r177 (  76 120 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.29 //y=0.17 //x2=7.29 //y2=0
r178 (  76 77 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=7.29 //y=0.17 //x2=7.29 //y2=0.45
r179 (  73 119 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.83 //y=0 //x2=6.66 //y2=0
r180 (  73 75 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=6.83 //y=0 //x2=7.03 //y2=0
r181 (  72 120 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.205 //y=0 //x2=7.29 //y2=0
r182 (  72 75 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=7.205 //y=0 //x2=7.03 //y2=0
r183 (  69 108 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.05 //y=0 //x2=5.965 //y2=0
r184 (  68 119 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.49 //y=0 //x2=6.66 //y2=0
r185 (  68 69 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.49 //y=0 //x2=6.05 //y2=0
r186 (  64 132 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.615 //x2=5.965 //y2=0.53
r187 (  64 132 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.615 //x2=5.965 //y2=0.88
r188 (  63 132 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.445 //x2=5.965 //y2=0.53
r189 (  62 108 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.17 //x2=5.965 //y2=0
r190 (  62 63 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.17 //x2=5.965 //y2=0.445
r191 (  61 132 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.565 //y=0.53 //x2=5.48 //y2=0.53
r192 (  60 132 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.88 //y=0.53 //x2=5.965 //y2=0.53
r193 (  60 61 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=5.88 //y=0.53 //x2=5.565 //y2=0.53
r194 (  59 132 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.48 //y=0.445 //x2=5.48 //y2=0.53
r195 (  58 105 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.48 //y=0.17 //x2=5.48 //y2=0
r196 (  58 59 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=5.48 //y=0.17 //x2=5.48 //y2=0.445
r197 (  57 132 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=5.08 //y=0.53 //x2=4.995 //y2=0.53
r198 (  56 132 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.395 //y=0.53 //x2=5.48 //y2=0.53
r199 (  56 57 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=5.395 //y=0.53 //x2=5.08 //y2=0.53
r200 (  52 132 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=4.995 //y=0.615 //x2=4.995 //y2=0.53
r201 (  52 132 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.995 //y=0.615 //x2=4.995 //y2=0.88
r202 (  51 132 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=4.995 //y=0.445 //x2=4.995 //y2=0.53
r203 (  50 104 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.995 //y=0.17 //x2=4.995 //y2=0
r204 (  50 51 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=4.995 //y=0.17 //x2=4.995 //y2=0.445
r205 (  49 132 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.595 //y=0.53 //x2=4.51 //y2=0.53
r206 (  48 132 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=4.91 //y=0.53 //x2=4.995 //y2=0.53
r207 (  48 49 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.91 //y=0.53 //x2=4.595 //y2=0.53
r208 (  47 132 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.51 //y=0.445 //x2=4.51 //y2=0.53
r209 (  46 103 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.51 //y=0.17 //x2=4.51 //y2=0
r210 (  46 47 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=4.51 //y=0.17 //x2=4.51 //y2=0.445
r211 (  45 132 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.11 //y=0.53 //x2=4.025 //y2=0.53
r212 (  44 132 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.425 //y=0.53 //x2=4.51 //y2=0.53
r213 (  44 45 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.425 //y=0.53 //x2=4.11 //y2=0.53
r214 (  40 132 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.615 //x2=4.025 //y2=0.53
r215 (  40 132 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.615 //x2=4.025 //y2=1.22
r216 (  39 132 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.445 //x2=4.025 //y2=0.53
r217 (  38 100 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.17 //x2=4.025 //y2=0
r218 (  38 39 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.17 //x2=4.025 //y2=0.445
r219 (  37 99 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.5 //y=0 //x2=3.33 //y2=0
r220 (  36 100 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.94 //y=0 //x2=4.025 //y2=0
r221 (  36 37 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=3.94 //y=0 //x2=3.5 //y2=0
r222 (  31 33 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r223 (  29 98 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.18 //y2=0
r224 (  29 31 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.85 //y2=0
r225 (  28 99 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.16 //y=0 //x2=3.33 //y2=0
r226 (  28 33 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r227 (  24 98 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r228 (  24 131 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.955
r229 (  20 98 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=1.18 //y2=0
r230 (  20 23 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=0.74 //y2=0
r231 (  16 123 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=0 //x2=8.14 //y2=0
r232 (  14 75 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=0 //x2=7.03 //y2=0
r233 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=0 //x2=8.14 //y2=0
r234 (  12 107 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r235 (  12 14 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=7.03 //y2=0
r236 (  8 33 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r237 (  6 31 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r238 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r239 (  3 23 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r240 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r241 (  1 102 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r242 (  1 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.55 //y2=0
r243 (  1 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=2.96 //y2=0
ends PM_AO3X1\%GND

subckt PM_AO3X1\%VDD ( 1 16 28 36 52 62 78 91 94 96 99 100 101 102 103 104 105 )
c102 ( 105 0 ) capacitor c=0.0451925f //x=8.07 //y=5.02
c103 ( 104 0 ) capacitor c=0.0429364f //x=7.2 //y=5.02
c104 ( 103 0 ) capacitor c=0.0256796f //x=4.415 //y=5.025
c105 ( 102 0 ) capacitor c=0.0383753f //x=2.405 //y=5.02
c106 ( 101 0 ) capacitor c=0.0243052f //x=1.525 //y=5.02
c107 ( 100 0 ) capacitor c=0.053196f //x=0.655 //y=5.02
c108 ( 99 0 ) capacitor c=0.234796f //x=8.14 //y=7.4
c109 ( 97 0 ) capacitor c=0.00591168f //x=7.335 //y=7.4
c110 ( 96 0 ) capacitor c=0.110627f //x=6.66 //y=7.4
c111 ( 95 0 ) capacitor c=0.00591168f //x=4.56 //y=7.4
c112 ( 94 0 ) capacitor c=0.116004f //x=3.33 //y=7.4
c113 ( 93 0 ) capacitor c=0.00591168f //x=2.55 //y=7.4
c114 ( 92 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c115 ( 91 0 ) capacitor c=0.24846f //x=0.74 //y=7.4
c116 ( 78 0 ) capacitor c=0.028745f //x=8.13 //y=7.4
c117 ( 68 0 ) capacitor c=0.0216067f //x=7.25 //y=7.4
c118 ( 62 0 ) capacitor c=0.0778183f //x=6.49 //y=7.4
c119 ( 52 0 ) capacitor c=0.0465804f //x=4.475 //y=7.4
c120 ( 46 0 ) capacitor c=0.0275781f //x=3.16 //y=7.4
c121 ( 36 0 ) capacitor c=0.0285035f //x=2.465 //y=7.4
c122 ( 28 0 ) capacitor c=0.0286367f //x=1.585 //y=7.4
c123 ( 16 0 ) capacitor c=0.353989f //x=8.14 //y=7.4
r124 (  80 99 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.215 //y=7.23 //x2=8.215 //y2=7.4
r125 (  80 105 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=8.215 //y=7.23 //x2=8.215 //y2=6.405
r126 (  79 97 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.42 //y=7.4 //x2=7.335 //y2=7.4
r127 (  78 99 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.13 //y=7.4 //x2=8.215 //y2=7.4
r128 (  78 79 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.13 //y=7.4 //x2=7.42 //y2=7.4
r129 (  72 97 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.335 //y=7.23 //x2=7.335 //y2=7.4
r130 (  72 104 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=7.335 //y=7.23 //x2=7.335 //y2=6.405
r131 (  69 96 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=6.83 //y=7.4 //x2=6.66 //y2=7.4
r132 (  69 71 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=6.83 //y=7.4 //x2=7.03 //y2=7.4
r133 (  68 97 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.25 //y=7.4 //x2=7.335 //y2=7.4
r134 (  68 71 ) resistor r=7.88796 //w=0.357 //l=0.22 //layer=li \
 //thickness=0.1 //x=7.25 //y=7.4 //x2=7.03 //y2=7.4
r135 (  63 95 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.645 //y=7.4 //x2=4.56 //y2=7.4
r136 (  63 65 ) resistor r=32.4482 //w=0.357 //l=0.905 //layer=li \
 //thickness=0.1 //x=4.645 //y=7.4 //x2=5.55 //y2=7.4
r137 (  62 96 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=6.49 //y=7.4 //x2=6.66 //y2=7.4
r138 (  62 65 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=6.49 //y=7.4 //x2=5.55 //y2=7.4
r139 (  56 95 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.56 //y=7.23 //x2=4.56 //y2=7.4
r140 (  56 103 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=4.56 //y=7.23 //x2=4.56 //y2=6.74
r141 (  53 94 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r142 (  53 55 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=3.5 //y=7.4 //x2=4.44 //y2=7.4
r143 (  52 95 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.475 //y=7.4 //x2=4.56 //y2=7.4
r144 (  52 55 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=4.475 //y=7.4 //x2=4.44 //y2=7.4
r145 (  47 93 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.55 //y2=7.4
r146 (  47 49 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.96 //y2=7.4
r147 (  46 94 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r148 (  46 49 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r149 (  40 93 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r150 (  40 102 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.745
r151 (  37 92 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r152 (  37 39 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r153 (  36 93 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r154 (  36 39 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r155 (  30 92 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r156 (  30 101 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.745
r157 (  29 91 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r158 (  28 92 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r159 (  28 29 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r160 (  22 91 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r161 (  22 100 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.405
r162 (  16 99 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=7.4 //x2=8.14 //y2=7.4
r163 (  14 71 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=7.4 //x2=7.03 //y2=7.4
r164 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=7.4 //x2=8.14 //y2=7.4
r165 (  12 65 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r166 (  12 14 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=7.03 //y2=7.4
r167 (  8 49 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r168 (  6 39 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r169 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r170 (  3 91 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r171 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r172 (  1 55 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r173 (  1 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.55 //y2=7.4
r174 (  1 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=2.96 //y2=7.4
ends PM_AO3X1\%VDD

subckt PM_AO3X1\%noxref_3 ( 1 2 13 14 25 27 28 32 35 39 41 43 44 45 46 47 48 \
 49 53 55 58 60 61 66 76 78 79 )
c144 ( 79 0 ) capacitor c=0.0220291f //x=1.965 //y=5.02
c145 ( 78 0 ) capacitor c=0.0217503f //x=1.085 //y=5.02
c146 ( 76 0 ) capacitor c=0.00865153f //x=1.96 //y=0.905
c147 ( 66 0 ) capacitor c=0.04214f //x=4.285 //y=4.705
c148 ( 61 0 ) capacitor c=0.0321911f //x=4.775 //y=1.25
c149 ( 60 0 ) capacitor c=0.0185201f //x=4.775 //y=0.905
c150 ( 58 0 ) capacitor c=0.0344254f //x=4.705 //y=4.795
c151 ( 55 0 ) capacitor c=0.0133656f //x=4.62 //y=1.405
c152 ( 53 0 ) capacitor c=0.0157804f //x=4.62 //y=0.75
c153 ( 49 0 ) capacitor c=0.0785055f //x=4.245 //y=1.915
c154 ( 48 0 ) capacitor c=0.022867f //x=4.245 //y=1.56
c155 ( 47 0 ) capacitor c=0.0234318f //x=4.245 //y=1.25
c156 ( 46 0 ) capacitor c=0.0192004f //x=4.245 //y=0.905
c157 ( 45 0 ) capacitor c=0.110795f //x=4.78 //y=6.025
c158 ( 44 0 ) capacitor c=0.153847f //x=4.34 //y=6.025
c159 ( 41 0 ) capacitor c=0.00995068f //x=4.285 //y=4.705
c160 ( 39 0 ) capacitor c=0.00427536f //x=2.11 //y=5.2
c161 ( 35 0 ) capacitor c=0.0968478f //x=4.44 //y=2.08
c162 ( 32 0 ) capacitor c=0.117241f //x=2.59 //y=2.59
c163 ( 28 0 ) capacitor c=0.00781917f //x=2.235 //y=1.655
c164 ( 27 0 ) capacitor c=0.0159132f //x=2.505 //y=1.655
c165 ( 25 0 ) capacitor c=0.017841f //x=2.505 //y=5.2
c166 ( 14 0 ) capacitor c=0.00387264f //x=1.315 //y=5.2
c167 ( 13 0 ) capacitor c=0.0222171f //x=2.025 //y=5.2
c168 ( 2 0 ) capacitor c=0.0173935f //x=2.705 //y=2.59
c169 ( 1 0 ) capacitor c=0.111807f //x=4.325 //y=2.59
r170 (  68 69 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=4.285 //y=4.795 //x2=4.285 //y2=4.87
r171 (  66 68 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=4.285 //y=4.705 //x2=4.285 //y2=4.795
r172 (  61 75 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.775 //y=1.25 //x2=4.735 //y2=1.405
r173 (  60 74 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.775 //y=0.905 //x2=4.735 //y2=0.75
r174 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.775 //y=0.905 //x2=4.775 //y2=1.25
r175 (  59 68 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=4.42 //y=4.795 //x2=4.285 //y2=4.795
r176 (  58 62 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.705 //y=4.795 //x2=4.78 //y2=4.87
r177 (  58 59 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=4.705 //y=4.795 //x2=4.42 //y2=4.795
r178 (  56 73 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.4 //y=1.405 //x2=4.285 //y2=1.405
r179 (  55 75 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.62 //y=1.405 //x2=4.735 //y2=1.405
r180 (  54 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.4 //y=0.75 //x2=4.285 //y2=0.75
r181 (  53 74 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.62 //y=0.75 //x2=4.735 //y2=0.75
r182 (  53 54 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.62 //y=0.75 //x2=4.4 //y2=0.75
r183 (  49 71 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.915 //x2=4.44 //y2=2.08
r184 (  48 73 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.56 //x2=4.285 //y2=1.405
r185 (  48 49 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.56 //x2=4.245 //y2=1.915
r186 (  47 73 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.25 //x2=4.285 //y2=1.405
r187 (  46 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.245 //y=0.905 //x2=4.285 //y2=0.75
r188 (  46 47 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.245 //y=0.905 //x2=4.245 //y2=1.25
r189 (  45 62 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.78 //y=6.025 //x2=4.78 //y2=4.87
r190 (  44 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.34 //y=6.025 //x2=4.34 //y2=4.87
r191 (  43 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.51 //y=1.405 //x2=4.62 //y2=1.405
r192 (  43 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.51 //y=1.405 //x2=4.4 //y2=1.405
r193 (  41 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.285 //y=4.705 //x2=4.285 //y2=4.705
r194 (  41 42 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=4.285 //y=4.705 //x2=4.44 //y2=4.705
r195 (  35 71 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=2.08 //x2=4.44 //y2=2.08
r196 (  35 38 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.08 //x2=4.44 //y2=2.59
r197 (  33 42 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=4.44 //y=4.54 //x2=4.44 //y2=4.705
r198 (  33 38 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=4.44 //y=4.54 //x2=4.44 //y2=2.59
r199 (  30 32 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.115 //x2=2.59 //y2=2.59
r200 (  29 32 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=2.59
r201 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r202 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r203 (  26 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.195 //y=5.2 //x2=2.11 //y2=5.2
r204 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.59 //y2=5.115
r205 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.195 //y2=5.2
r206 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.235 //y2=1.655
r207 (  21 76 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r208 (  15 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.2
r209 (  15 79 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.725
r210 (  13 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=2.11 //y2=5.2
r211 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=1.315 //y2=5.2
r212 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.315 //y2=5.2
r213 (  7 78 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.23 //y2=5.725
r214 (  6 38 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=2.59 //x2=4.44 //y2=2.59
r215 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=2.59 //x2=2.59 //y2=2.59
r216 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=2.59 //x2=2.59 //y2=2.59
r217 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.325 //y=2.59 //x2=4.44 //y2=2.59
r218 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=4.325 //y=2.59 //x2=2.705 //y2=2.59
ends PM_AO3X1\%noxref_3

subckt PM_AO3X1\%noxref_4 ( 1 2 11 12 23 24 25 30 32 40 41 42 43 44 45 46 50 \
 51 52 54 60 61 63 71 72 75 )
c133 ( 75 0 ) capacitor c=0.0159573f //x=5.295 //y=5.025
c134 ( 72 0 ) capacitor c=0.00905936f //x=5.29 //y=0.905
c135 ( 71 0 ) capacitor c=0.007684f //x=4.32 //y=0.905
c136 ( 63 0 ) capacitor c=0.0517753f //x=7.4 //y=2.085
c137 ( 61 0 ) capacitor c=0.0435629f //x=8.04 //y=1.255
c138 ( 60 0 ) capacitor c=0.0200386f //x=8.04 //y=0.91
c139 ( 54 0 ) capacitor c=0.0152946f //x=7.885 //y=1.41
c140 ( 52 0 ) capacitor c=0.0157804f //x=7.885 //y=0.755
c141 ( 51 0 ) capacitor c=0.0524991f //x=7.63 //y=4.79
c142 ( 50 0 ) capacitor c=0.0322983f //x=7.92 //y=4.79
c143 ( 46 0 ) capacitor c=0.0290017f //x=7.51 //y=1.92
c144 ( 45 0 ) capacitor c=0.0250027f //x=7.51 //y=1.565
c145 ( 44 0 ) capacitor c=0.0234316f //x=7.51 //y=1.255
c146 ( 43 0 ) capacitor c=0.0200596f //x=7.51 //y=0.91
c147 ( 42 0 ) capacitor c=0.154218f //x=7.995 //y=6.02
c148 ( 41 0 ) capacitor c=0.154243f //x=7.555 //y=6.02
c149 ( 39 0 ) capacitor c=0.00710337f //x=5.48 //y=1.655
c150 ( 32 0 ) capacitor c=0.0948753f //x=7.4 //y=2.085
c151 ( 30 0 ) capacitor c=0.11371f //x=5.92 //y=2.59
c152 ( 25 0 ) capacitor c=0.0160526f //x=5.835 //y=1.655
c153 ( 24 0 ) capacitor c=0.00499395f //x=5.525 //y=5.21
c154 ( 23 0 ) capacitor c=0.0166531f //x=5.835 //y=5.21
c155 ( 12 0 ) capacitor c=0.00220849f //x=4.595 //y=1.655
c156 ( 11 0 ) capacitor c=0.0280953f //x=5.395 //y=1.655
c157 ( 2 0 ) capacitor c=0.0119578f //x=6.035 //y=2.59
c158 ( 1 0 ) capacitor c=0.093442f //x=7.285 //y=2.59
r159 (  63 64 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.4 //y=2.085 //x2=7.51 //y2=2.085
r160 (  61 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.04 //y=1.255 //x2=8 //y2=1.41
r161 (  60 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.04 //y=0.91 //x2=8 //y2=0.755
r162 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.04 //y=0.91 //x2=8.04 //y2=1.255
r163 (  55 68 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.665 //y=1.41 //x2=7.55 //y2=1.41
r164 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.885 //y=1.41 //x2=8 //y2=1.41
r165 (  53 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.665 //y=0.755 //x2=7.55 //y2=0.755
r166 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.885 //y=0.755 //x2=8 //y2=0.755
r167 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.885 //y=0.755 //x2=7.665 //y2=0.755
r168 (  50 57 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.92 //y=4.79 //x2=7.995 //y2=4.865
r169 (  50 51 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=7.92 //y=4.79 //x2=7.63 //y2=4.79
r170 (  47 51 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.555 //y=4.865 //x2=7.63 //y2=4.79
r171 (  47 66 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=7.555 //y=4.865 //x2=7.4 //y2=4.7
r172 (  46 64 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=7.51 //y=1.92 //x2=7.51 //y2=2.085
r173 (  45 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.51 //y=1.565 //x2=7.55 //y2=1.41
r174 (  45 46 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=7.51 //y=1.565 //x2=7.51 //y2=1.92
r175 (  44 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.51 //y=1.255 //x2=7.55 //y2=1.41
r176 (  43 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.51 //y=0.91 //x2=7.55 //y2=0.755
r177 (  43 44 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.51 //y=0.91 //x2=7.51 //y2=1.255
r178 (  42 57 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.995 //y=6.02 //x2=7.995 //y2=4.865
r179 (  41 47 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.555 //y=6.02 //x2=7.555 //y2=4.865
r180 (  40 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.775 //y=1.41 //x2=7.885 //y2=1.41
r181 (  40 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.775 //y=1.41 //x2=7.665 //y2=1.41
r182 (  37 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.4 //y=4.7 //x2=7.4 //y2=4.7
r183 (  35 37 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=7.4 //y=2.59 //x2=7.4 //y2=4.7
r184 (  32 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.4 //y=2.085 //x2=7.4 //y2=2.085
r185 (  32 35 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=7.4 //y=2.085 //x2=7.4 //y2=2.59
r186 (  28 30 ) resistor r=173.519 //w=0.187 //l=2.535 //layer=li \
 //thickness=0.1 //x=5.92 //y=5.125 //x2=5.92 //y2=2.59
r187 (  27 30 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=5.92 //y=1.74 //x2=5.92 //y2=2.59
r188 (  26 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.565 //y=1.655 //x2=5.48 //y2=1.655
r189 (  25 27 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.835 //y=1.655 //x2=5.92 //y2=1.74
r190 (  25 26 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=5.835 //y=1.655 //x2=5.565 //y2=1.655
r191 (  23 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.835 //y=5.21 //x2=5.92 //y2=5.125
r192 (  23 24 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=5.835 //y=5.21 //x2=5.525 //y2=5.21
r193 (  19 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.48 //y=1.57 //x2=5.48 //y2=1.655
r194 (  19 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=5.48 //y=1.57 //x2=5.48 //y2=1
r195 (  13 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.44 //y=5.295 //x2=5.525 //y2=5.21
r196 (  13 75 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=5.44 //y=5.295 //x2=5.44 //y2=5.72
r197 (  11 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.395 //y=1.655 //x2=5.48 //y2=1.655
r198 (  11 12 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=5.395 //y=1.655 //x2=4.595 //y2=1.655
r199 (  7 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.51 //y=1.57 //x2=4.595 //y2=1.655
r200 (  7 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=4.51 //y=1.57 //x2=4.51 //y2=1
r201 (  6 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=7.4 \
 //y=2.59 //x2=7.4 //y2=2.59
r202 (  4 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=2.59 //x2=5.92 //y2=2.59
r203 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=2.59 //x2=5.92 //y2=2.59
r204 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=2.59 //x2=7.4 //y2=2.59
r205 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=2.59 //x2=6.035 //y2=2.59
ends PM_AO3X1\%noxref_4

subckt PM_AO3X1\%A ( 1 2 3 4 5 6 7 9 21 22 23 24 25 26 27 31 33 36 37 47 )
c55 ( 47 0 ) capacitor c=0.0667949f //x=1.11 //y=4.7
c56 ( 37 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c57 ( 36 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c58 ( 33 0 ) capacitor c=0.0141798f //x=1.29 //y=1.365
c59 ( 31 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c60 ( 27 0 ) capacitor c=0.0860049f //x=0.915 //y=1.915
c61 ( 26 0 ) capacitor c=0.0229722f //x=0.915 //y=1.52
c62 ( 25 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c63 ( 24 0 ) capacitor c=0.0199343f //x=0.915 //y=0.865
c64 ( 23 0 ) capacitor c=0.110275f //x=1.45 //y=6.02
c65 ( 22 0 ) capacitor c=0.154305f //x=1.01 //y=6.02
c66 ( 9 0 ) capacitor c=0.116498f //x=1.11 //y=2.08
r67 (  45 47 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.7 //x2=1.11 //y2=4.7
r68 (  38 47 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=1.45 //y=4.865 //x2=1.11 //y2=4.7
r69 (  37 49 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r70 (  36 48 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r71 (  36 37 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r72 (  34 44 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r73 (  33 49 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r74 (  32 43 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r75 (  31 48 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r76 (  31 32 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r77 (  28 45 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.865 //x2=1.01 //y2=4.7
r78 (  27 42 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r79 (  26 44 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r80 (  26 27 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r81 (  25 44 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r82 (  24 43 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r83 (  24 25 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r84 (  23 38 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.02 //x2=1.45 //y2=4.865
r85 (  22 28 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.02 //x2=1.01 //y2=4.865
r86 (  21 33 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r87 (  21 34 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r88 (  19 47 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r89 (  9 42 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r90 (  7 19 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.44 //x2=1.11 //y2=4.7
r91 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r92 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r93 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r94 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r95 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r96 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.22 //x2=1.11 //y2=2.59
r97 (  1 9 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.22 //x2=1.11 //y2=2.08
ends PM_AO3X1\%A

subckt PM_AO3X1\%B ( 1 2 3 4 5 6 7 8 10 21 22 23 24 25 26 31 33 35 41 42 44 45 \
 48 )
c64 ( 48 0 ) capacitor c=0.034715f //x=1.88 //y=4.7
c65 ( 45 0 ) capacitor c=0.0279499f //x=1.85 //y=1.915
c66 ( 44 0 ) capacitor c=0.0437302f //x=1.85 //y=2.08
c67 ( 42 0 ) capacitor c=0.0429696f //x=2.415 //y=1.25
c68 ( 41 0 ) capacitor c=0.0192208f //x=2.415 //y=0.905
c69 ( 35 0 ) capacitor c=0.0158629f //x=2.26 //y=1.405
c70 ( 33 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c71 ( 31 0 ) capacitor c=0.0366192f //x=2.255 //y=4.79
c72 ( 26 0 ) capacitor c=0.0205163f //x=1.885 //y=1.56
c73 ( 25 0 ) capacitor c=0.0168481f //x=1.885 //y=1.25
c74 ( 24 0 ) capacitor c=0.0174783f //x=1.885 //y=0.905
c75 ( 23 0 ) capacitor c=0.15358f //x=2.33 //y=6.02
c76 ( 22 0 ) capacitor c=0.110281f //x=1.89 //y=6.02
c77 ( 10 0 ) capacitor c=0.0813556f //x=1.85 //y=2.08
c78 ( 8 0 ) capacitor c=0.00453889f //x=1.85 //y=4.535
r79 (  50 51 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.79 //x2=1.88 //y2=4.865
r80 (  48 50 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.7 //x2=1.88 //y2=4.79
r81 (  44 45 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r82 (  42 55 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r83 (  41 54 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r84 (  41 42 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r85 (  36 53 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r86 (  35 55 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r87 (  34 52 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r88 (  33 54 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r89 (  33 34 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r90 (  32 50 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.015 //y=4.79 //x2=1.88 //y2=4.79
r91 (  31 38 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.33 //y2=4.865
r92 (  31 32 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.015 //y2=4.79
r93 (  26 53 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r94 (  26 45 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r95 (  25 53 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r96 (  24 52 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r97 (  24 25 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r98 (  23 38 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.02 //x2=2.33 //y2=4.865
r99 (  22 51 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.02 //x2=1.89 //y2=4.865
r100 (  21 35 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r101 (  21 36 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r102 (  20 48 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.88 //y=4.7 //x2=1.88 //y2=4.7
r103 (  10 44 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r104 (  8 20 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.865 //y2=4.7
r105 (  7 8 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.44 //x2=1.85 //y2=4.535
r106 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=4.07 //x2=1.85 //y2=4.44
r107 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=3.7 //x2=1.85 //y2=4.07
r108 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=3.33 //x2=1.85 //y2=3.7
r109 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=2.96 //x2=1.85 //y2=3.33
r110 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=2.59 //x2=1.85 //y2=2.96
r111 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=2.22 //x2=1.85 //y2=2.59
r112 (  1 10 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.22 //x2=1.85 //y2=2.08
ends PM_AO3X1\%B

subckt PM_AO3X1\%noxref_7 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632971f //x=0.56 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722223f //x=2.635 //y=0.615
c53 ( 13 0 ) capacitor c=0.0154397f //x=2.55 //y=0.53
c54 ( 10 0 ) capacitor c=0.0092508f //x=1.665 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c56 ( 5 0 ) capacitor c=0.0255599f //x=1.58 //y=1.58
c57 ( 1 0 ) capacitor c=0.0113547f //x=0.695 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=2.15 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.15 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_AO3X1\%noxref_7

subckt PM_AO3X1\%C ( 1 2 3 4 5 6 7 8 10 21 22 23 24 25 26 31 33 35 41 42 44 45 \
 48 )
c71 ( 48 0 ) capacitor c=0.0369822f //x=5.215 //y=4.705
c72 ( 45 0 ) capacitor c=0.0279572f //x=5.18 //y=1.915
c73 ( 44 0 ) capacitor c=0.0422144f //x=5.18 //y=2.08
c74 ( 42 0 ) capacitor c=0.0237734f //x=5.745 //y=1.255
c75 ( 41 0 ) capacitor c=0.0191782f //x=5.745 //y=0.905
c76 ( 35 0 ) capacitor c=0.0346941f //x=5.59 //y=1.405
c77 ( 33 0 ) capacitor c=0.0157803f //x=5.59 //y=0.75
c78 ( 31 0 ) capacitor c=0.0360787f //x=5.585 //y=4.795
c79 ( 26 0 ) capacitor c=0.0199921f //x=5.215 //y=1.56
c80 ( 25 0 ) capacitor c=0.0169608f //x=5.215 //y=1.255
c81 ( 24 0 ) capacitor c=0.0185462f //x=5.215 //y=0.905
c82 ( 23 0 ) capacitor c=0.15325f //x=5.66 //y=6.025
c83 ( 22 0 ) capacitor c=0.110232f //x=5.22 //y=6.025
c84 ( 10 0 ) capacitor c=0.0800125f //x=5.18 //y=2.08
c85 ( 8 0 ) capacitor c=0.00521267f //x=5.18 //y=4.54
r86 (  50 51 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=5.215 //y=4.795 //x2=5.215 //y2=4.87
r87 (  48 50 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=5.215 //y=4.705 //x2=5.215 //y2=4.795
r88 (  44 45 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=5.18 //y=2.08 //x2=5.18 //y2=1.915
r89 (  42 55 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=5.745 //y=1.255 //x2=5.745 //y2=1.367
r90 (  41 54 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.745 //y=0.905 //x2=5.705 //y2=0.75
r91 (  41 42 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=5.745 //y=0.905 //x2=5.745 //y2=1.255
r92 (  36 53 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.37 //y=1.405 //x2=5.255 //y2=1.405
r93 (  35 55 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=5.59 //y=1.405 //x2=5.745 //y2=1.367
r94 (  34 52 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.37 //y=0.75 //x2=5.255 //y2=0.75
r95 (  33 54 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.59 //y=0.75 //x2=5.705 //y2=0.75
r96 (  33 34 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.59 //y=0.75 //x2=5.37 //y2=0.75
r97 (  32 50 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=5.35 //y=4.795 //x2=5.215 //y2=4.795
r98 (  31 38 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.585 //y=4.795 //x2=5.66 //y2=4.87
r99 (  31 32 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=5.585 //y=4.795 //x2=5.35 //y2=4.795
r100 (  26 53 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.215 //y=1.56 //x2=5.255 //y2=1.405
r101 (  26 45 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=5.215 //y=1.56 //x2=5.215 //y2=1.915
r102 (  25 53 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=5.215 //y=1.255 //x2=5.255 //y2=1.405
r103 (  24 52 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.215 //y=0.905 //x2=5.255 //y2=0.75
r104 (  24 25 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=5.215 //y=0.905 //x2=5.215 //y2=1.255
r105 (  23 38 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.66 //y=6.025 //x2=5.66 //y2=4.87
r106 (  22 51 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.22 //y=6.025 //x2=5.22 //y2=4.87
r107 (  21 35 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.48 //y=1.405 //x2=5.59 //y2=1.405
r108 (  21 36 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.48 //y=1.405 //x2=5.37 //y2=1.405
r109 (  20 48 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.215 //y=4.705 //x2=5.215 //y2=4.705
r110 (  10 44 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.18 //y=2.08 //x2=5.18 //y2=2.08
r111 (  8 20 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=5.18 //y=4.54 //x2=5.197 //y2=4.705
r112 (  7 8 ) resistor r=6.84492 //w=0.187 //l=0.1 //layer=li //thickness=0.1 \
 //x=5.18 //y=4.44 //x2=5.18 //y2=4.54
r113 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=5.18 //y=4.07 //x2=5.18 //y2=4.44
r114 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=5.18 //y=3.7 //x2=5.18 //y2=4.07
r115 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=5.18 //y=3.33 //x2=5.18 //y2=3.7
r116 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=5.18 //y=2.96 //x2=5.18 //y2=3.33
r117 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=5.18 //y=2.59 //x2=5.18 //y2=2.96
r118 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=5.18 //y=2.22 //x2=5.18 //y2=2.59
r119 (  1 10 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=5.18 //y=2.22 //x2=5.18 //y2=2.08
ends PM_AO3X1\%C

subckt PM_AO3X1\%noxref_9 ( 7 8 15 16 23 24 25 )
c43 ( 25 0 ) capacitor c=0.0308836f //x=5.735 //y=5.025
c44 ( 24 0 ) capacitor c=0.0185379f //x=4.855 //y=5.025
c45 ( 23 0 ) capacitor c=0.0409962f //x=3.985 //y=5.025
c46 ( 16 0 ) capacitor c=0.00193672f //x=5.085 //y=6.91
c47 ( 15 0 ) capacitor c=0.01354f //x=5.795 //y=6.91
c48 ( 8 0 ) capacitor c=0.00844339f //x=4.205 //y=5.21
c49 ( 7 0 ) capacitor c=0.0252644f //x=4.915 //y=5.21
r50 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.88 //y=6.825 //x2=5.88 //y2=6.74
r51 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.795 //y=6.91 //x2=5.88 //y2=6.825
r52 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.795 //y=6.91 //x2=5.085 //y2=6.91
r53 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5 //y=6.825 //x2=5.085 //y2=6.91
r54 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=5 //y=6.825 //x2=5 //y2=6.4
r55 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=5 //y=5.295 //x2=5 //y2=5.72
r56 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.915 //y=5.21 //x2=5 //y2=5.295
r57 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=4.915 //y=5.21 //x2=4.205 //y2=5.21
r58 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.12 //y=5.295 //x2=4.205 //y2=5.21
r59 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=4.12 //y=5.295 //x2=4.12 //y2=5.72
ends PM_AO3X1\%noxref_9

subckt PM_AO3X1\%Y ( 1 2 3 4 5 6 7 18 19 20 21 31 33 )
c43 ( 33 0 ) capacitor c=0.028734f //x=7.63 //y=5.02
c44 ( 31 0 ) capacitor c=0.0173218f //x=7.585 //y=0.91
c45 ( 21 0 ) capacitor c=0.00575887f //x=7.86 //y=4.58
c46 ( 20 0 ) capacitor c=0.0146395f //x=8.055 //y=4.58
c47 ( 19 0 ) capacitor c=0.00636159f //x=7.855 //y=2.08
c48 ( 18 0 ) capacitor c=0.0141837f //x=8.055 //y=2.08
c49 ( 1 0 ) capacitor c=0.105613f //x=8.14 //y=2.22
r50 (  20 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.055 //y=4.58 //x2=8.14 //y2=4.495
r51 (  20 21 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=8.055 //y=4.58 //x2=7.86 //y2=4.58
r52 (  18 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.055 //y=2.08 //x2=8.14 //y2=2.165
r53 (  18 19 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=8.055 //y=2.08 //x2=7.855 //y2=2.08
r54 (  12 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.775 //y=4.665 //x2=7.86 //y2=4.58
r55 (  12 33 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=7.775 //y=4.665 //x2=7.775 //y2=5.725
r56 (  8 19 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.77 //y=1.995 //x2=7.855 //y2=2.08
r57 (  8 31 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=7.77 //y=1.995 //x2=7.77 //y2=1.005
r58 (  7 23 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=8.14 //y=4.44 //x2=8.14 //y2=4.495
r59 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=8.14 //y=4.07 //x2=8.14 //y2=4.44
r60 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=8.14 //y=3.7 //x2=8.14 //y2=4.07
r61 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=8.14 //y=3.33 //x2=8.14 //y2=3.7
r62 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=8.14 //y=2.96 //x2=8.14 //y2=3.33
r63 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=8.14 //y=2.59 //x2=8.14 //y2=2.96
r64 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=8.14 //y=2.22 //x2=8.14 //y2=2.59
r65 (  1 22 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.22 //x2=8.14 //y2=2.165
ends PM_AO3X1\%Y

