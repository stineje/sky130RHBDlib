* SPICE3 file created from DLATCH.ext - technology: sky130A

.subckt DLATCH Q D GATE VPB VNB
M1000 VPB.t7 GATE a_661_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VPB.t15 a_1295_182.t3 a_2795_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPB.t3 D a_1771_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_661_1004.t2 GATE VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1771_1004.t0 D VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_2405_182.t1 a_1771_1004.t5 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VNB GATE a_1666_73.t0 nshort w=-1.605u l=1.765u
+  ad=7.6538p pd=53.32u as=0p ps=0u
M1007 Q a_3007_383.t4 a_2795_1005.t2 pshort w=2u l=0.15u
+  ad=0.58p pd=4.58u as=0p ps=0u
M1008 a_3461_1005.t3 a_2405_182.t4 a_3007_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_661_1004.t3 a_185_182.t3 VPB.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1771_1004.t4 GATE VPB.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPB.t1 Q a_3461_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_2795_1005.t0 a_1295_182.t4 VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 Q a_1295_182.t5 VNB.t3 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.15u as=0p ps=0u
M1014 VPB.t4 D a_185_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPB.t14 a_661_1004.t5 a_1295_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 Q a_3007_383.t5 VNB.t1 nshort w=-1.83u l=2.06u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t16 a_185_182.t5 a_661_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPB.t9 GATE a_1771_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VNB a_185_182.t4 a_556_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_3007_383.t2 a_2405_182.t5 a_3461_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPB.t17 a_1771_1004.t7 a_2405_182.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_2795_1005.t3 a_3007_383.t6 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_185_182.t0 D VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1295_182.t1 a_661_1004.t7 VPB.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_3461_1005.t0 Q VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 Q VPB 0.34fF
C1 VPB D 0.62fF
C2 GATE D 0.58fF
C3 GATE VPB 0.15fF
R0 a_556_73.t0 a_556_73.n1 93.333
R1 a_556_73.n4 a_556_73.n2 55.07
R2 a_556_73.t0 a_556_73.n0 8.137
R3 a_556_73.n4 a_556_73.n3 4.619
R4 a_556_73.t0 a_556_73.n4 0.071
R5 a_661_1004.n4 a_661_1004.t5 512.525
R6 a_661_1004.n4 a_661_1004.t7 371.139
R7 a_661_1004.n5 a_661_1004.t6 220.263
R8 a_661_1004.n8 a_661_1004.n6 194.086
R9 a_661_1004.n6 a_661_1004.n3 162.547
R10 a_661_1004.n5 a_661_1004.n4 158.3
R11 a_661_1004.n6 a_661_1004.n5 153.043
R12 a_661_1004.n3 a_661_1004.n2 76.002
R13 a_661_1004.n9 a_661_1004.n0 55.263
R14 a_661_1004.n8 a_661_1004.n7 30
R15 a_661_1004.n9 a_661_1004.n8 23.684
R16 a_661_1004.n1 a_661_1004.t0 14.282
R17 a_661_1004.n1 a_661_1004.t2 14.282
R18 a_661_1004.n2 a_661_1004.t4 14.282
R19 a_661_1004.n2 a_661_1004.t3 14.282
R20 a_661_1004.n3 a_661_1004.n1 12.85
R21 VPB VPB.n400 126.832
R22 VPB.n63 VPB.n61 94.117
R23 VPB.n374 VPB.n372 94.117
R24 VPB.n327 VPB.n325 94.117
R25 VPB.n157 VPB.n155 94.117
R26 VPB.n136 VPB.n134 94.117
R27 VPB.n239 VPB.n237 94.117
R28 VPB.n199 VPB.n198 76
R29 VPB.n206 VPB.n205 76
R30 VPB.n210 VPB.n209 76
R31 VPB.n214 VPB.n213 76
R32 VPB.n241 VPB.n240 76
R33 VPB.n245 VPB.n244 76
R34 VPB.n249 VPB.n248 76
R35 VPB.n253 VPB.n252 76
R36 VPB.n258 VPB.n257 76
R37 VPB.n271 VPB.n268 76
R38 VPB.n276 VPB.n78 76
R39 VPB.n283 VPB.n282 76
R40 VPB.n288 VPB.n287 76
R41 VPB.n293 VPB.n292 76
R42 VPB.n298 VPB.n297 76
R43 VPB.n302 VPB.n301 76
R44 VPB.n329 VPB.n328 76
R45 VPB.n335 VPB.n334 76
R46 VPB.n339 VPB.n338 76
R47 VPB.n345 VPB.n344 76
R48 VPB.n349 VPB.n348 76
R49 VPB.n376 VPB.n375 76
R50 VPB.n381 VPB.n380 76
R51 VPB.n393 VPB.n392 76
R52 VPB.n147 VPB.n146 68.979
R53 VPB.n342 VPB.n341 68.979
R54 VPB.n74 VPB.n73 68.979
R55 VPB.n140 VPB.n139 64.528
R56 VPB.n332 VPB.n331 64.528
R57 VPB.n67 VPB.n66 64.528
R58 VPB.n20 VPB.n19 61.764
R59 VPB.n356 VPB.n355 61.764
R60 VPB.n309 VPB.n308 61.764
R61 VPB.n85 VPB.n84 61.764
R62 VPB.n106 VPB.n105 61.764
R63 VPB.n221 VPB.n220 61.764
R64 VPB.n77 VPB.t5 55.106
R65 VPB.n65 VPB.t4 55.106
R66 VPB.n53 VPB.t10 55.106
R67 VPB.n340 VPB.t13 55.106
R68 VPB.n330 VPB.t14 55.106
R69 VPB.n294 VPB.t8 55.106
R70 VPB.n150 VPB.t12 55.106
R71 VPB.n138 VPB.t17 55.106
R72 VPB.n377 VPB.t7 55.106
R73 VPB.n272 VPB.t3 55.106
R74 VPB.n274 VPB.n273 48.952
R75 VPB.n37 VPB.n36 48.952
R76 VPB.n203 VPB.n202 44.502
R77 VPB.n124 VPB.n123 44.502
R78 VPB.n290 VPB.n289 44.502
R79 VPB.n50 VPB.n49 44.502
R80 VPB.n122 VPB.n121 41.183
R81 VPB.n201 VPB.n200 41.183
R82 VPB.n44 VPB.n35 40.824
R83 VPB.n278 VPB.n277 40.824
R84 VPB.n193 VPB.n192 35.118
R85 VPB.n397 VPB.n393 20.452
R86 VPB.n182 VPB.n179 20.452
R87 VPB.n280 VPB.n279 17.801
R88 VPB.n41 VPB.n40 17.801
R89 VPB.n35 VPB.t6 14.282
R90 VPB.n35 VPB.t16 14.282
R91 VPB.n277 VPB.t2 14.282
R92 VPB.n277 VPB.t9 14.282
R93 VPB.n121 VPB.t11 14.282
R94 VPB.n121 VPB.t15 14.282
R95 VPB.n200 VPB.t0 14.282
R96 VPB.n200 VPB.t1 14.282
R97 VPB.n182 VPB.n181 13.653
R98 VPB.n181 VPB.n180 13.653
R99 VPB.n191 VPB.n190 13.653
R100 VPB.n190 VPB.n189 13.653
R101 VPB.n188 VPB.n187 13.653
R102 VPB.n187 VPB.n186 13.653
R103 VPB.n185 VPB.n184 13.653
R104 VPB.n184 VPB.n183 13.653
R105 VPB.n198 VPB.n197 13.653
R106 VPB.n197 VPB.n196 13.653
R107 VPB.n205 VPB.n204 13.653
R108 VPB.n204 VPB.n203 13.653
R109 VPB.n209 VPB.n208 13.653
R110 VPB.n208 VPB.n207 13.653
R111 VPB.n213 VPB.n212 13.653
R112 VPB.n212 VPB.n211 13.653
R113 VPB.n240 VPB.n239 13.653
R114 VPB.n239 VPB.n238 13.653
R115 VPB.n244 VPB.n243 13.653
R116 VPB.n243 VPB.n242 13.653
R117 VPB.n248 VPB.n247 13.653
R118 VPB.n247 VPB.n246 13.653
R119 VPB.n252 VPB.n251 13.653
R120 VPB.n251 VPB.n250 13.653
R121 VPB.n257 VPB.n256 13.653
R122 VPB.n256 VPB.n255 13.653
R123 VPB.n126 VPB.n125 13.653
R124 VPB.n125 VPB.n124 13.653
R125 VPB.n129 VPB.n128 13.653
R126 VPB.n128 VPB.n127 13.653
R127 VPB.n132 VPB.n131 13.653
R128 VPB.n131 VPB.n130 13.653
R129 VPB.n137 VPB.n136 13.653
R130 VPB.n136 VPB.n135 13.653
R131 VPB.n142 VPB.n141 13.653
R132 VPB.n141 VPB.n140 13.653
R133 VPB.n145 VPB.n144 13.653
R134 VPB.n144 VPB.n143 13.653
R135 VPB.n149 VPB.n148 13.653
R136 VPB.n148 VPB.n147 13.653
R137 VPB.n153 VPB.n152 13.653
R138 VPB.n152 VPB.n151 13.653
R139 VPB.n158 VPB.n157 13.653
R140 VPB.n157 VPB.n156 13.653
R141 VPB.n271 VPB.n270 13.653
R142 VPB.n270 VPB.n269 13.653
R143 VPB.n276 VPB.n275 13.653
R144 VPB.n275 VPB.n274 13.653
R145 VPB.n282 VPB.n281 13.653
R146 VPB.n281 VPB.n280 13.653
R147 VPB.n287 VPB.n286 13.653
R148 VPB.n286 VPB.n285 13.653
R149 VPB.n292 VPB.n291 13.653
R150 VPB.n291 VPB.n290 13.653
R151 VPB.n297 VPB.n296 13.653
R152 VPB.n296 VPB.n295 13.653
R153 VPB.n301 VPB.n300 13.653
R154 VPB.n300 VPB.n299 13.653
R155 VPB.n328 VPB.n327 13.653
R156 VPB.n327 VPB.n326 13.653
R157 VPB.n334 VPB.n333 13.653
R158 VPB.n333 VPB.n332 13.653
R159 VPB.n338 VPB.n337 13.653
R160 VPB.n337 VPB.n336 13.653
R161 VPB.n344 VPB.n343 13.653
R162 VPB.n343 VPB.n342 13.653
R163 VPB.n348 VPB.n347 13.653
R164 VPB.n347 VPB.n346 13.653
R165 VPB.n375 VPB.n374 13.653
R166 VPB.n374 VPB.n373 13.653
R167 VPB.n380 VPB.n379 13.653
R168 VPB.n379 VPB.n378 13.653
R169 VPB.n39 VPB.n38 13.653
R170 VPB.n38 VPB.n37 13.653
R171 VPB.n43 VPB.n42 13.653
R172 VPB.n42 VPB.n41 13.653
R173 VPB.n48 VPB.n47 13.653
R174 VPB.n47 VPB.n46 13.653
R175 VPB.n52 VPB.n51 13.653
R176 VPB.n51 VPB.n50 13.653
R177 VPB.n56 VPB.n55 13.653
R178 VPB.n55 VPB.n54 13.653
R179 VPB.n59 VPB.n58 13.653
R180 VPB.n58 VPB.n57 13.653
R181 VPB.n64 VPB.n63 13.653
R182 VPB.n63 VPB.n62 13.653
R183 VPB.n69 VPB.n68 13.653
R184 VPB.n68 VPB.n67 13.653
R185 VPB.n72 VPB.n71 13.653
R186 VPB.n71 VPB.n70 13.653
R187 VPB.n76 VPB.n75 13.653
R188 VPB.n75 VPB.n74 13.653
R189 VPB.n393 VPB.n0 13.653
R190 VPB VPB.n0 13.653
R191 VPB.n196 VPB.n195 13.35
R192 VPB.n255 VPB.n254 13.35
R193 VPB.n285 VPB.n284 13.35
R194 VPB.n46 VPB.n45 13.35
R195 VPB.n397 VPB.n396 13.276
R196 VPB.n396 VPB.n394 13.276
R197 VPB.n34 VPB.n16 13.276
R198 VPB.n16 VPB.n14 13.276
R199 VPB.n370 VPB.n352 13.276
R200 VPB.n352 VPB.n350 13.276
R201 VPB.n323 VPB.n305 13.276
R202 VPB.n305 VPB.n303 13.276
R203 VPB.n99 VPB.n81 13.276
R204 VPB.n81 VPB.n79 13.276
R205 VPB.n120 VPB.n102 13.276
R206 VPB.n102 VPB.n100 13.276
R207 VPB.n235 VPB.n217 13.276
R208 VPB.n217 VPB.n215 13.276
R209 VPB.n191 VPB.n188 13.276
R210 VPB.n188 VPB.n185 13.276
R211 VPB.n240 VPB.n236 13.276
R212 VPB.n129 VPB.n126 13.276
R213 VPB.n132 VPB.n129 13.276
R214 VPB.n133 VPB.n132 13.276
R215 VPB.n137 VPB.n133 13.276
R216 VPB.n145 VPB.n142 13.276
R217 VPB.n149 VPB.n145 13.276
R218 VPB.n154 VPB.n153 13.276
R219 VPB.n158 VPB.n154 13.276
R220 VPB.n271 VPB.n158 13.276
R221 VPB.n282 VPB.n276 13.276
R222 VPB.n328 VPB.n324 13.276
R223 VPB.n375 VPB.n371 13.276
R224 VPB.n43 VPB.n39 13.276
R225 VPB.n52 VPB.n48 13.276
R226 VPB.n59 VPB.n56 13.276
R227 VPB.n60 VPB.n59 13.276
R228 VPB.n64 VPB.n60 13.276
R229 VPB.n72 VPB.n69 13.276
R230 VPB.n76 VPB.n72 13.276
R231 VPB.n179 VPB.n161 13.276
R232 VPB.n161 VPB.n159 13.276
R233 VPB.n166 VPB.n164 12.796
R234 VPB.n166 VPB.n165 12.564
R235 VPB.n174 VPB.n173 12.198
R236 VPB.n170 VPB.n169 12.198
R237 VPB.n174 VPB.n171 12.198
R238 VPB.n276 VPB.n272 11.841
R239 VPB.n53 VPB.n52 11.482
R240 VPB.n153 VPB.n150 10.944
R241 VPB.n393 VPB.n77 10.944
R242 VPB.n138 VPB.n137 10.585
R243 VPB.n65 VPB.n64 10.585
R244 VPB.n179 VPB.n178 7.5
R245 VPB.n164 VPB.n163 7.5
R246 VPB.n169 VPB.n168 7.5
R247 VPB.n173 VPB.n172 7.5
R248 VPB.n161 VPB.n160 7.5
R249 VPB.n176 VPB.n162 7.5
R250 VPB.n217 VPB.n216 7.5
R251 VPB.n230 VPB.n229 7.5
R252 VPB.n224 VPB.n223 7.5
R253 VPB.n226 VPB.n225 7.5
R254 VPB.n219 VPB.n218 7.5
R255 VPB.n235 VPB.n234 7.5
R256 VPB.n102 VPB.n101 7.5
R257 VPB.n115 VPB.n114 7.5
R258 VPB.n109 VPB.n108 7.5
R259 VPB.n111 VPB.n110 7.5
R260 VPB.n104 VPB.n103 7.5
R261 VPB.n120 VPB.n119 7.5
R262 VPB.n81 VPB.n80 7.5
R263 VPB.n94 VPB.n93 7.5
R264 VPB.n88 VPB.n87 7.5
R265 VPB.n90 VPB.n89 7.5
R266 VPB.n83 VPB.n82 7.5
R267 VPB.n99 VPB.n98 7.5
R268 VPB.n305 VPB.n304 7.5
R269 VPB.n318 VPB.n317 7.5
R270 VPB.n312 VPB.n311 7.5
R271 VPB.n314 VPB.n313 7.5
R272 VPB.n307 VPB.n306 7.5
R273 VPB.n323 VPB.n322 7.5
R274 VPB.n352 VPB.n351 7.5
R275 VPB.n365 VPB.n364 7.5
R276 VPB.n359 VPB.n358 7.5
R277 VPB.n361 VPB.n360 7.5
R278 VPB.n354 VPB.n353 7.5
R279 VPB.n370 VPB.n369 7.5
R280 VPB.n16 VPB.n15 7.5
R281 VPB.n29 VPB.n28 7.5
R282 VPB.n23 VPB.n22 7.5
R283 VPB.n25 VPB.n24 7.5
R284 VPB.n18 VPB.n17 7.5
R285 VPB.n34 VPB.n33 7.5
R286 VPB.n396 VPB.n395 7.5
R287 VPB.n12 VPB.n11 7.5
R288 VPB.n6 VPB.n5 7.5
R289 VPB.n8 VPB.n7 7.5
R290 VPB.n2 VPB.n1 7.5
R291 VPB.n398 VPB.n397 7.5
R292 VPB.n60 VPB.n34 7.176
R293 VPB.n371 VPB.n370 7.176
R294 VPB.n324 VPB.n323 7.176
R295 VPB.n154 VPB.n99 7.176
R296 VPB.n133 VPB.n120 7.176
R297 VPB.n236 VPB.n235 7.176
R298 VPB.n48 VPB.n44 6.817
R299 VPB.n231 VPB.n228 6.729
R300 VPB.n227 VPB.n224 6.729
R301 VPB.n222 VPB.n219 6.729
R302 VPB.n116 VPB.n113 6.729
R303 VPB.n112 VPB.n109 6.729
R304 VPB.n107 VPB.n104 6.729
R305 VPB.n95 VPB.n92 6.729
R306 VPB.n91 VPB.n88 6.729
R307 VPB.n86 VPB.n83 6.729
R308 VPB.n319 VPB.n316 6.729
R309 VPB.n315 VPB.n312 6.729
R310 VPB.n310 VPB.n307 6.729
R311 VPB.n366 VPB.n363 6.729
R312 VPB.n362 VPB.n359 6.729
R313 VPB.n357 VPB.n354 6.729
R314 VPB.n30 VPB.n27 6.729
R315 VPB.n26 VPB.n23 6.729
R316 VPB.n21 VPB.n18 6.729
R317 VPB.n13 VPB.n10 6.729
R318 VPB.n9 VPB.n6 6.729
R319 VPB.n4 VPB.n2 6.729
R320 VPB.n222 VPB.n221 6.728
R321 VPB.n227 VPB.n226 6.728
R322 VPB.n231 VPB.n230 6.728
R323 VPB.n234 VPB.n233 6.728
R324 VPB.n107 VPB.n106 6.728
R325 VPB.n112 VPB.n111 6.728
R326 VPB.n116 VPB.n115 6.728
R327 VPB.n119 VPB.n118 6.728
R328 VPB.n86 VPB.n85 6.728
R329 VPB.n91 VPB.n90 6.728
R330 VPB.n95 VPB.n94 6.728
R331 VPB.n98 VPB.n97 6.728
R332 VPB.n310 VPB.n309 6.728
R333 VPB.n315 VPB.n314 6.728
R334 VPB.n319 VPB.n318 6.728
R335 VPB.n322 VPB.n321 6.728
R336 VPB.n357 VPB.n356 6.728
R337 VPB.n362 VPB.n361 6.728
R338 VPB.n366 VPB.n365 6.728
R339 VPB.n369 VPB.n368 6.728
R340 VPB.n21 VPB.n20 6.728
R341 VPB.n26 VPB.n25 6.728
R342 VPB.n30 VPB.n29 6.728
R343 VPB.n33 VPB.n32 6.728
R344 VPB.n4 VPB.n3 6.728
R345 VPB.n9 VPB.n8 6.728
R346 VPB.n13 VPB.n12 6.728
R347 VPB.n399 VPB.n398 6.728
R348 VPB.n282 VPB.n278 6.458
R349 VPB.n44 VPB.n43 6.458
R350 VPB.n178 VPB.n177 6.398
R351 VPB.n192 VPB.n182 6.112
R352 VPB.n192 VPB.n191 6.101
R353 VPB.n205 VPB.n201 4.305
R354 VPB.n126 VPB.n122 4.305
R355 VPB.n142 VPB.n138 2.691
R356 VPB.n334 VPB.n330 2.691
R357 VPB.n69 VPB.n65 2.691
R358 VPB.n150 VPB.n149 2.332
R359 VPB.n344 VPB.n340 2.332
R360 VPB.n77 VPB.n76 2.332
R361 VPB.n297 VPB.n294 1.794
R362 VPB.n56 VPB.n53 1.794
R363 VPB.n272 VPB.n271 1.435
R364 VPB.n380 VPB.n377 1.435
R365 VPB.n176 VPB.n167 1.402
R366 VPB.n176 VPB.n170 1.402
R367 VPB.n176 VPB.n174 1.402
R368 VPB.n176 VPB.n175 1.402
R369 VPB.n177 VPB.n176 0.735
R370 VPB.n176 VPB.n166 0.735
R371 VPB.n232 VPB.n231 0.387
R372 VPB.n232 VPB.n227 0.387
R373 VPB.n232 VPB.n222 0.387
R374 VPB.n233 VPB.n232 0.387
R375 VPB.n117 VPB.n116 0.387
R376 VPB.n117 VPB.n112 0.387
R377 VPB.n117 VPB.n107 0.387
R378 VPB.n118 VPB.n117 0.387
R379 VPB.n96 VPB.n95 0.387
R380 VPB.n96 VPB.n91 0.387
R381 VPB.n96 VPB.n86 0.387
R382 VPB.n97 VPB.n96 0.387
R383 VPB.n320 VPB.n319 0.387
R384 VPB.n320 VPB.n315 0.387
R385 VPB.n320 VPB.n310 0.387
R386 VPB.n321 VPB.n320 0.387
R387 VPB.n367 VPB.n366 0.387
R388 VPB.n367 VPB.n362 0.387
R389 VPB.n367 VPB.n357 0.387
R390 VPB.n368 VPB.n367 0.387
R391 VPB.n31 VPB.n30 0.387
R392 VPB.n31 VPB.n26 0.387
R393 VPB.n31 VPB.n21 0.387
R394 VPB.n32 VPB.n31 0.387
R395 VPB.n400 VPB.n13 0.387
R396 VPB.n400 VPB.n9 0.387
R397 VPB.n400 VPB.n4 0.387
R398 VPB.n400 VPB.n399 0.387
R399 VPB.n241 VPB.n214 0.272
R400 VPB.n262 VPB.n261 0.272
R401 VPB.n267 VPB.n266 0.272
R402 VPB.n329 VPB.n302 0.272
R403 VPB.n376 VPB.n349 0.272
R404 VPB.n388 VPB.n387 0.272
R405 VPB.n392 VPB 0.198
R406 VPB.n194 VPB.n193 0.136
R407 VPB.n199 VPB.n194 0.136
R408 VPB.n206 VPB.n199 0.136
R409 VPB.n210 VPB.n206 0.136
R410 VPB.n214 VPB.n210 0.136
R411 VPB.n245 VPB.n241 0.136
R412 VPB.n249 VPB.n245 0.136
R413 VPB.n253 VPB.n249 0.136
R414 VPB.n258 VPB.n253 0.136
R415 VPB.n259 VPB.n258 0.136
R416 VPB.n260 VPB.n259 0.136
R417 VPB.n261 VPB.n260 0.136
R418 VPB.n263 VPB.n262 0.136
R419 VPB.n264 VPB.n263 0.136
R420 VPB.n265 VPB.n264 0.136
R421 VPB.n266 VPB.n265 0.136
R422 VPB.n268 VPB.n267 0.136
R423 VPB.n268 VPB.n78 0.136
R424 VPB.n283 VPB.n78 0.136
R425 VPB.n288 VPB.n283 0.136
R426 VPB.n293 VPB.n288 0.136
R427 VPB.n298 VPB.n293 0.136
R428 VPB.n302 VPB.n298 0.136
R429 VPB.n335 VPB.n329 0.136
R430 VPB.n339 VPB.n335 0.136
R431 VPB.n345 VPB.n339 0.136
R432 VPB.n349 VPB.n345 0.136
R433 VPB.n381 VPB.n376 0.136
R434 VPB.n382 VPB.n381 0.136
R435 VPB.n383 VPB.n382 0.136
R436 VPB.n384 VPB.n383 0.136
R437 VPB.n385 VPB.n384 0.136
R438 VPB.n386 VPB.n385 0.136
R439 VPB.n387 VPB.n386 0.136
R440 VPB.n389 VPB.n388 0.136
R441 VPB.n390 VPB.n389 0.136
R442 VPB.n391 VPB.n390 0.136
R443 VPB.n392 VPB.n391 0.136
R444 a_1295_182.n2 a_1295_182.t4 486.819
R445 a_1295_182.n2 a_1295_182.t3 384.527
R446 a_1295_182.n3 a_1295_182.t5 287.101
R447 a_1295_182.n6 a_1295_182.n4 215.257
R448 a_1295_182.n4 a_1295_182.n3 157.396
R449 a_1295_182.n4 a_1295_182.n1 140.59
R450 a_1295_182.n3 a_1295_182.n2 90.041
R451 a_1295_182.n6 a_1295_182.n5 30
R452 a_1295_182.n7 a_1295_182.n0 24.383
R453 a_1295_182.n7 a_1295_182.n6 23.684
R454 a_1295_182.n1 a_1295_182.t2 14.282
R455 a_1295_182.n1 a_1295_182.t1 14.282
R456 a_2795_1005.t1 a_2795_1005.n0 101.66
R457 a_2795_1005.n0 a_2795_1005.t3 101.659
R458 a_2795_1005.n0 a_2795_1005.t2 14.294
R459 a_2795_1005.n0 a_2795_1005.t0 14.282
R460 a_1771_1004.n4 a_1771_1004.t7 512.525
R461 a_1771_1004.n4 a_1771_1004.t5 371.139
R462 a_1771_1004.n5 a_1771_1004.t6 220.263
R463 a_1771_1004.n8 a_1771_1004.n6 194.086
R464 a_1771_1004.n6 a_1771_1004.n3 162.547
R465 a_1771_1004.n5 a_1771_1004.n4 158.3
R466 a_1771_1004.n6 a_1771_1004.n5 153.043
R467 a_1771_1004.n3 a_1771_1004.n2 76.002
R468 a_1771_1004.n8 a_1771_1004.n7 30
R469 a_1771_1004.n9 a_1771_1004.n0 24.383
R470 a_1771_1004.n9 a_1771_1004.n8 23.684
R471 a_1771_1004.n1 a_1771_1004.t1 14.282
R472 a_1771_1004.n1 a_1771_1004.t0 14.282
R473 a_1771_1004.n2 a_1771_1004.t3 14.282
R474 a_1771_1004.n2 a_1771_1004.t4 14.282
R475 a_1771_1004.n3 a_1771_1004.n1 12.85
R476 a_1666_73.t0 a_1666_73.n1 93.333
R477 a_1666_73.n4 a_1666_73.n2 55.07
R478 a_1666_73.t0 a_1666_73.n0 8.137
R479 a_1666_73.n4 a_1666_73.n3 4.619
R480 a_1666_73.t0 a_1666_73.n4 0.071
R481 VNB VNB.n420 300.778
R482 VNB.n241 VNB.n240 199.897
R483 VNB.n114 VNB.n113 199.897
R484 VNB.n85 VNB.n84 199.897
R485 VNB.n328 VNB.n327 199.897
R486 VNB.n380 VNB.n379 199.897
R487 VNB.n27 VNB.n26 199.897
R488 VNB.n147 VNB.n146 158.304
R489 VNB.n66 VNB.n65 158.304
R490 VNB.n250 VNB.n248 154.509
R491 VNB.n161 VNB.n159 154.509
R492 VNB.n137 VNB.n135 154.509
R493 VNB.n389 VNB.n387 154.509
R494 VNB.n337 VNB.n335 154.509
R495 VNB.n56 VNB.n54 154.509
R496 VNB.n205 VNB.n204 121.366
R497 VNB.n141 VNB.n140 105.536
R498 VNB.n60 VNB.n59 105.536
R499 VNB.n305 VNB.n304 84.842
R500 VNB.n43 VNB.n33 84.842
R501 VNB.n188 VNB.n180 76.136
R502 VNB.n188 VNB.n187 76
R503 VNB.n295 VNB.n74 76
R504 VNB.n407 VNB.n406 76
R505 VNB.n395 VNB.n394 76
R506 VNB.n391 VNB.n390 76
R507 VNB.n369 VNB.n368 76
R508 VNB.n365 VNB.n364 76
R509 VNB.n357 VNB.n356 76
R510 VNB.n348 VNB.n347 76
R511 VNB.n339 VNB.n338 76
R512 VNB.n317 VNB.n316 76
R513 VNB.n313 VNB.n312 76
R514 VNB.n309 VNB.n308 76
R515 VNB.n303 VNB.n302 76
R516 VNB.n299 VNB.n298 76
R517 VNB.n292 VNB.n289 76
R518 VNB.n279 VNB.n278 76
R519 VNB.n271 VNB.n270 76
R520 VNB.n267 VNB.n266 76
R521 VNB.n260 VNB.n259 76
R522 VNB.n252 VNB.n251 76
R523 VNB.n230 VNB.n229 76
R524 VNB.n226 VNB.n225 76
R525 VNB.n218 VNB.n217 76
R526 VNB.n209 VNB.n208 76
R527 VNB.n199 VNB.n198 76
R528 VNB.n195 VNB.n194 76
R529 VNB.n355 VNB.n354 49.896
R530 VNB.n220 VNB.t0 39.412
R531 VNB.n94 VNB.t2 39.412
R532 VNB.n7 VNB.t5 39.412
R533 VNB.n206 VNB.n205 36.937
R534 VNB.n276 VNB.n275 36.937
R535 VNB.n307 VNB.n306 36.678
R536 VNB.n45 VNB.n44 36.678
R537 VNB.n193 VNB.n192 36.267
R538 VNB.n265 VNB.n264 36.267
R539 VNB.n103 VNB.n102 35.01
R540 VNB.n343 VNB.n342 35.01
R541 VNB.n16 VNB.n15 35.01
R542 VNB.n341 VNB.n340 29.127
R543 VNB.n215 VNB.n214 27.855
R544 VNB.n148 VNB.n145 27.855
R545 VNB.n67 VNB.n64 27.855
R546 VNB.n351 VNB.t7 20.794
R547 VNB.n180 VNB.n177 20.452
R548 VNB.n408 VNB.n407 20.452
R549 VNB.n139 VNB.n103 20.094
R550 VNB.n144 VNB.n99 20.094
R551 VNB.n154 VNB.n95 20.094
R552 VNB.n344 VNB.n343 20.094
R553 VNB.n353 VNB.n352 20.094
R554 VNB.n361 VNB.n360 20.094
R555 VNB.n58 VNB.n16 20.094
R556 VNB.n63 VNB.n12 20.094
R557 VNB.n73 VNB.n8 20.094
R558 VNB.n212 VNB.n211 19.735
R559 VNB.n203 VNB.n202 19.735
R560 VNB.n191 VNB.n190 19.735
R561 VNB.n184 VNB.n183 19.735
R562 VNB.n222 VNB.n221 19.735
R563 VNB.n124 VNB.n123 19.735
R564 VNB.n274 VNB.n273 19.735
R565 VNB.n263 VNB.n262 19.735
R566 VNB.n256 VNB.n255 19.735
R567 VNB.n130 VNB.n122 19.735
R568 VNB.n190 VNB.t4 19.724
R569 VNB.n262 VNB.t1 19.724
R570 VNB.n103 VNB.n101 19.017
R571 VNB.n343 VNB.n341 19.017
R572 VNB.n16 VNB.n14 19.017
R573 VNB.n121 VNB.t3 17.353
R574 VNB.n220 VNB.n219 17.185
R575 VNB.n94 VNB.n93 17.185
R576 VNB.n7 VNB.n6 17.185
R577 VNB.n216 VNB.n215 16.721
R578 VNB.n149 VNB.n148 16.721
R579 VNB.n68 VNB.n67 16.721
R580 VNB.n201 VNB.n200 13.654
R581 VNB.n187 VNB.n186 13.653
R582 VNB.n186 VNB.n185 13.653
R583 VNB.n194 VNB.n193 13.653
R584 VNB.n198 VNB.n197 13.653
R585 VNB.n197 VNB.n196 13.653
R586 VNB.n208 VNB.n207 13.653
R587 VNB.n207 VNB.n206 13.653
R588 VNB.n217 VNB.n216 13.653
R589 VNB.n225 VNB.n224 13.653
R590 VNB.n224 VNB.n223 13.653
R591 VNB.n229 VNB.n228 13.653
R592 VNB.n228 VNB.n227 13.653
R593 VNB.n251 VNB.n250 13.653
R594 VNB.n250 VNB.n249 13.653
R595 VNB.n259 VNB.n258 13.653
R596 VNB.n258 VNB.n257 13.653
R597 VNB.n266 VNB.n265 13.653
R598 VNB.n270 VNB.n269 13.653
R599 VNB.n269 VNB.n268 13.653
R600 VNB.n278 VNB.n277 13.653
R601 VNB.n277 VNB.n276 13.653
R602 VNB.n126 VNB.n125 13.653
R603 VNB.n129 VNB.n128 13.653
R604 VNB.n128 VNB.n127 13.653
R605 VNB.n133 VNB.n132 13.653
R606 VNB.n132 VNB.n131 13.653
R607 VNB.n138 VNB.n137 13.653
R608 VNB.n137 VNB.n136 13.653
R609 VNB.n143 VNB.n142 13.653
R610 VNB.n142 VNB.n141 13.653
R611 VNB.n150 VNB.n149 13.653
R612 VNB.n153 VNB.n152 13.653
R613 VNB.n152 VNB.n151 13.653
R614 VNB.n157 VNB.n156 13.653
R615 VNB.n156 VNB.n155 13.653
R616 VNB.n162 VNB.n161 13.653
R617 VNB.n161 VNB.n160 13.653
R618 VNB.n292 VNB.n291 13.653
R619 VNB.n291 VNB.n290 13.653
R620 VNB.n295 VNB.n294 13.653
R621 VNB.n294 VNB.n293 13.653
R622 VNB.n298 VNB.n297 13.653
R623 VNB.n297 VNB.n296 13.653
R624 VNB.n302 VNB.n301 13.653
R625 VNB.n301 VNB.n300 13.653
R626 VNB.n308 VNB.n307 13.653
R627 VNB.n312 VNB.n311 13.653
R628 VNB.n311 VNB.n310 13.653
R629 VNB.n316 VNB.n315 13.653
R630 VNB.n315 VNB.n314 13.653
R631 VNB.n338 VNB.n337 13.653
R632 VNB.n337 VNB.n336 13.653
R633 VNB.n347 VNB.n346 13.653
R634 VNB.n346 VNB.n345 13.653
R635 VNB.n356 VNB.n355 13.653
R636 VNB.n364 VNB.n363 13.653
R637 VNB.n363 VNB.n362 13.653
R638 VNB.n368 VNB.n367 13.653
R639 VNB.n367 VNB.n366 13.653
R640 VNB.n390 VNB.n389 13.653
R641 VNB.n389 VNB.n388 13.653
R642 VNB.n394 VNB.n393 13.653
R643 VNB.n393 VNB.n392 13.653
R644 VNB.n36 VNB.n35 13.653
R645 VNB.n35 VNB.n34 13.653
R646 VNB.n39 VNB.n38 13.653
R647 VNB.n38 VNB.n37 13.653
R648 VNB.n42 VNB.n41 13.653
R649 VNB.n41 VNB.n40 13.653
R650 VNB.n46 VNB.n45 13.653
R651 VNB.n49 VNB.n48 13.653
R652 VNB.n48 VNB.n47 13.653
R653 VNB.n52 VNB.n51 13.653
R654 VNB.n51 VNB.n50 13.653
R655 VNB.n57 VNB.n56 13.653
R656 VNB.n56 VNB.n55 13.653
R657 VNB.n62 VNB.n61 13.653
R658 VNB.n61 VNB.n60 13.653
R659 VNB.n69 VNB.n68 13.653
R660 VNB.n72 VNB.n71 13.653
R661 VNB.n71 VNB.n70 13.653
R662 VNB.n407 VNB.n0 13.653
R663 VNB VNB.n0 13.653
R664 VNB.n180 VNB.n179 13.653
R665 VNB.n179 VNB.n178 13.653
R666 VNB.n415 VNB.n412 13.577
R667 VNB.n165 VNB.n163 13.276
R668 VNB.n177 VNB.n165 13.276
R669 VNB.n233 VNB.n231 13.276
R670 VNB.n246 VNB.n233 13.276
R671 VNB.n106 VNB.n104 13.276
R672 VNB.n119 VNB.n106 13.276
R673 VNB.n77 VNB.n75 13.276
R674 VNB.n90 VNB.n77 13.276
R675 VNB.n320 VNB.n318 13.276
R676 VNB.n333 VNB.n320 13.276
R677 VNB.n372 VNB.n370 13.276
R678 VNB.n385 VNB.n372 13.276
R679 VNB.n19 VNB.n17 13.276
R680 VNB.n32 VNB.n19 13.276
R681 VNB.n251 VNB.n247 13.276
R682 VNB.n129 VNB.n126 13.276
R683 VNB.n134 VNB.n133 13.276
R684 VNB.n138 VNB.n134 13.276
R685 VNB.n153 VNB.n150 13.276
R686 VNB.n158 VNB.n157 13.276
R687 VNB.n162 VNB.n158 13.276
R688 VNB.n292 VNB.n162 13.276
R689 VNB.n295 VNB.n292 13.276
R690 VNB.n298 VNB.n295 13.276
R691 VNB.n338 VNB.n334 13.276
R692 VNB.n390 VNB.n386 13.276
R693 VNB.n39 VNB.n36 13.276
R694 VNB.n42 VNB.n39 13.276
R695 VNB.n49 VNB.n46 13.276
R696 VNB.n52 VNB.n49 13.276
R697 VNB.n53 VNB.n52 13.276
R698 VNB.n57 VNB.n53 13.276
R699 VNB.n72 VNB.n69 13.276
R700 VNB.n3 VNB.n1 13.276
R701 VNB.n408 VNB.n3 13.276
R702 VNB.n144 VNB.n143 13.097
R703 VNB.n63 VNB.n62 13.097
R704 VNB.n122 VNB.n121 12.837
R705 VNB.n360 VNB.n359 12.837
R706 VNB.n133 VNB.n130 11.661
R707 VNB.n183 VNB.n182 11.605
R708 VNB.n255 VNB.n254 11.605
R709 VNB.n43 VNB.n42 10.764
R710 VNB.n182 VNB.n181 9.809
R711 VNB.n254 VNB.n253 9.809
R712 VNB.n157 VNB.n154 9.329
R713 VNB.n407 VNB.n73 9.329
R714 VNB.n139 VNB.n138 8.97
R715 VNB.n58 VNB.n57 8.97
R716 VNB.n121 VNB.n120 7.566
R717 VNB.n359 VNB.n358 7.566
R718 VNB.n211 VNB.n210 7.5
R719 VNB.n101 VNB.n100 7.5
R720 VNB.n98 VNB.n97 7.5
R721 VNB.n14 VNB.n13 7.5
R722 VNB.n11 VNB.n10 7.5
R723 VNB.n417 VNB.n416 7.5
R724 VNB.n239 VNB.n238 7.5
R725 VNB.n235 VNB.n234 7.5
R726 VNB.n233 VNB.n232 7.5
R727 VNB.n246 VNB.n245 7.5
R728 VNB.n112 VNB.n111 7.5
R729 VNB.n108 VNB.n107 7.5
R730 VNB.n106 VNB.n105 7.5
R731 VNB.n119 VNB.n118 7.5
R732 VNB.n83 VNB.n82 7.5
R733 VNB.n79 VNB.n78 7.5
R734 VNB.n77 VNB.n76 7.5
R735 VNB.n90 VNB.n89 7.5
R736 VNB.n326 VNB.n325 7.5
R737 VNB.n322 VNB.n321 7.5
R738 VNB.n320 VNB.n319 7.5
R739 VNB.n333 VNB.n332 7.5
R740 VNB.n378 VNB.n377 7.5
R741 VNB.n374 VNB.n373 7.5
R742 VNB.n372 VNB.n371 7.5
R743 VNB.n385 VNB.n384 7.5
R744 VNB.n25 VNB.n24 7.5
R745 VNB.n21 VNB.n20 7.5
R746 VNB.n19 VNB.n18 7.5
R747 VNB.n32 VNB.n31 7.5
R748 VNB.n409 VNB.n408 7.5
R749 VNB.n3 VNB.n2 7.5
R750 VNB.n414 VNB.n413 7.5
R751 VNB.n171 VNB.n170 7.5
R752 VNB.n167 VNB.n166 7.5
R753 VNB.n165 VNB.n164 7.5
R754 VNB.n177 VNB.n176 7.5
R755 VNB.n247 VNB.n246 7.176
R756 VNB.n134 VNB.n119 7.176
R757 VNB.n158 VNB.n90 7.176
R758 VNB.n334 VNB.n333 7.176
R759 VNB.n386 VNB.n385 7.176
R760 VNB.n53 VNB.n32 7.176
R761 VNB.t4 VNB.n189 7.04
R762 VNB.t1 VNB.n261 7.04
R763 VNB.n419 VNB.n417 7.011
R764 VNB.n242 VNB.n239 7.011
R765 VNB.n237 VNB.n235 7.011
R766 VNB.n115 VNB.n112 7.011
R767 VNB.n110 VNB.n108 7.011
R768 VNB.n86 VNB.n83 7.011
R769 VNB.n81 VNB.n79 7.011
R770 VNB.n329 VNB.n326 7.011
R771 VNB.n324 VNB.n322 7.011
R772 VNB.n381 VNB.n378 7.011
R773 VNB.n376 VNB.n374 7.011
R774 VNB.n28 VNB.n25 7.011
R775 VNB.n23 VNB.n21 7.011
R776 VNB.n173 VNB.n171 7.011
R777 VNB.n169 VNB.n167 7.011
R778 VNB.n245 VNB.n244 7.01
R779 VNB.n237 VNB.n236 7.01
R780 VNB.n242 VNB.n241 7.01
R781 VNB.n118 VNB.n117 7.01
R782 VNB.n110 VNB.n109 7.01
R783 VNB.n115 VNB.n114 7.01
R784 VNB.n89 VNB.n88 7.01
R785 VNB.n81 VNB.n80 7.01
R786 VNB.n86 VNB.n85 7.01
R787 VNB.n332 VNB.n331 7.01
R788 VNB.n324 VNB.n323 7.01
R789 VNB.n329 VNB.n328 7.01
R790 VNB.n384 VNB.n383 7.01
R791 VNB.n376 VNB.n375 7.01
R792 VNB.n381 VNB.n380 7.01
R793 VNB.n31 VNB.n30 7.01
R794 VNB.n23 VNB.n22 7.01
R795 VNB.n28 VNB.n27 7.01
R796 VNB.n176 VNB.n175 7.01
R797 VNB.n169 VNB.n168 7.01
R798 VNB.n173 VNB.n172 7.01
R799 VNB.n419 VNB.n418 7.01
R800 VNB.n415 VNB.n414 6.788
R801 VNB.n410 VNB.n409 6.788
R802 VNB.n208 VNB.n203 6.638
R803 VNB.n278 VNB.n274 6.638
R804 VNB.n221 VNB.n220 6.139
R805 VNB.n95 VNB.n94 6.139
R806 VNB.n8 VNB.n7 6.139
R807 VNB.n202 VNB.n201 5.774
R808 VNB.n273 VNB.n272 5.774
R809 VNB.n92 VNB.n91 4.551
R810 VNB.n350 VNB.n349 4.551
R811 VNB.n5 VNB.n4 4.551
R812 VNB.n143 VNB.n139 4.305
R813 VNB.n347 VNB.n344 4.305
R814 VNB.n62 VNB.n58 4.305
R815 VNB.n154 VNB.n153 3.947
R816 VNB.n364 VNB.n361 3.947
R817 VNB.n73 VNB.n72 3.947
R818 VNB.n194 VNB.n191 2.511
R819 VNB.n217 VNB.n212 2.511
R820 VNB.n266 VNB.n263 2.511
R821 VNB.n126 VNB.n124 2.511
R822 VNB.n308 VNB.n305 2.511
R823 VNB.n46 VNB.n43 2.511
R824 VNB.t2 VNB.n92 2.238
R825 VNB.t7 VNB.n350 2.238
R826 VNB.t5 VNB.n5 2.238
R827 VNB.n215 VNB.n213 1.99
R828 VNB.n148 VNB.n147 1.99
R829 VNB.n67 VNB.n66 1.99
R830 VNB.n97 VNB.n96 1.935
R831 VNB.n10 VNB.n9 1.935
R832 VNB.n187 VNB.n184 1.614
R833 VNB.n225 VNB.n222 1.614
R834 VNB.n259 VNB.n256 1.614
R835 VNB.n130 VNB.n129 1.614
R836 VNB.n420 VNB.n411 0.921
R837 VNB.n420 VNB.n415 0.476
R838 VNB.n420 VNB.n410 0.475
R839 VNB.n99 VNB.n98 0.358
R840 VNB.n352 VNB.n351 0.358
R841 VNB.n12 VNB.n11 0.358
R842 VNB.n252 VNB.n230 0.272
R843 VNB.n283 VNB.n282 0.272
R844 VNB.n288 VNB.n287 0.272
R845 VNB.n339 VNB.n317 0.272
R846 VNB.n391 VNB.n369 0.272
R847 VNB.n402 VNB.n401 0.272
R848 VNB.n243 VNB.n237 0.246
R849 VNB.n244 VNB.n243 0.246
R850 VNB.n243 VNB.n242 0.246
R851 VNB.n116 VNB.n110 0.246
R852 VNB.n117 VNB.n116 0.246
R853 VNB.n116 VNB.n115 0.246
R854 VNB.n87 VNB.n81 0.246
R855 VNB.n88 VNB.n87 0.246
R856 VNB.n87 VNB.n86 0.246
R857 VNB.n330 VNB.n324 0.246
R858 VNB.n331 VNB.n330 0.246
R859 VNB.n330 VNB.n329 0.246
R860 VNB.n382 VNB.n376 0.246
R861 VNB.n383 VNB.n382 0.246
R862 VNB.n382 VNB.n381 0.246
R863 VNB.n29 VNB.n23 0.246
R864 VNB.n30 VNB.n29 0.246
R865 VNB.n29 VNB.n28 0.246
R866 VNB.n174 VNB.n169 0.246
R867 VNB.n175 VNB.n174 0.246
R868 VNB.n174 VNB.n173 0.246
R869 VNB.n420 VNB.n419 0.246
R870 VNB.n406 VNB 0.198
R871 VNB.n150 VNB.n144 0.179
R872 VNB.n356 VNB.n353 0.179
R873 VNB.n69 VNB.n63 0.179
R874 VNB.n195 VNB.n188 0.136
R875 VNB.n199 VNB.n195 0.136
R876 VNB.n209 VNB.n199 0.136
R877 VNB.n218 VNB.n209 0.136
R878 VNB.n226 VNB.n218 0.136
R879 VNB.n230 VNB.n226 0.136
R880 VNB.n260 VNB.n252 0.136
R881 VNB.n267 VNB.n260 0.136
R882 VNB.n271 VNB.n267 0.136
R883 VNB.n279 VNB.n271 0.136
R884 VNB.n280 VNB.n279 0.136
R885 VNB.n281 VNB.n280 0.136
R886 VNB.n282 VNB.n281 0.136
R887 VNB.n284 VNB.n283 0.136
R888 VNB.n285 VNB.n284 0.136
R889 VNB.n286 VNB.n285 0.136
R890 VNB.n287 VNB.n286 0.136
R891 VNB.n289 VNB.n288 0.136
R892 VNB.n289 VNB.n74 0.136
R893 VNB.n299 VNB.n74 0.136
R894 VNB.n303 VNB.n299 0.136
R895 VNB.n309 VNB.n303 0.136
R896 VNB.n313 VNB.n309 0.136
R897 VNB.n317 VNB.n313 0.136
R898 VNB.n348 VNB.n339 0.136
R899 VNB.n357 VNB.n348 0.136
R900 VNB.n365 VNB.n357 0.136
R901 VNB.n369 VNB.n365 0.136
R902 VNB.n395 VNB.n391 0.136
R903 VNB.n396 VNB.n395 0.136
R904 VNB.n397 VNB.n396 0.136
R905 VNB.n398 VNB.n397 0.136
R906 VNB.n399 VNB.n398 0.136
R907 VNB.n400 VNB.n399 0.136
R908 VNB.n401 VNB.n400 0.136
R909 VNB.n403 VNB.n402 0.136
R910 VNB.n404 VNB.n403 0.136
R911 VNB.n405 VNB.n404 0.136
R912 VNB.n406 VNB.n405 0.136
R913 a_2405_182.n1 a_2405_182.t4 470.752
R914 a_2405_182.n1 a_2405_182.t5 384.527
R915 a_2405_182.n2 a_2405_182.t3 277.772
R916 a_2405_182.n5 a_2405_182.n3 248.332
R917 a_2405_182.n3 a_2405_182.n2 156.307
R918 a_2405_182.n3 a_2405_182.n0 114.038
R919 a_2405_182.n2 a_2405_182.n1 67.114
R920 a_2405_182.n5 a_2405_182.n4 15.218
R921 a_2405_182.n0 a_2405_182.t0 14.282
R922 a_2405_182.n0 a_2405_182.t1 14.282
R923 a_2405_182.n6 a_2405_182.n5 12.014
R924 a_3007_383.n1 a_3007_383.t6 470.752
R925 a_3007_383.n1 a_3007_383.t4 384.527
R926 a_3007_383.n2 a_3007_383.t5 251.219
R927 a_3007_383.n7 a_3007_383.n3 172.234
R928 a_3007_383.n3 a_3007_383.n2 154.947
R929 a_3007_383.n3 a_3007_383.n0 148.83
R930 a_3007_383.n7 a_3007_383.n6 133.539
R931 a_3007_383.n2 a_3007_383.n1 93.667
R932 a_3007_383.n9 a_3007_383.n7 55.263
R933 a_3007_383.n6 a_3007_383.n5 22.578
R934 a_3007_383.n9 a_3007_383.n8 15.001
R935 a_3007_383.n0 a_3007_383.t1 14.282
R936 a_3007_383.n0 a_3007_383.t2 14.282
R937 a_3007_383.n10 a_3007_383.n9 12.632
R938 a_3007_383.n6 a_3007_383.n4 8.58
R939 a_3461_1005.t1 a_3461_1005.n0 101.66
R940 a_3461_1005.n0 a_3461_1005.t3 101.659
R941 a_3461_1005.n0 a_3461_1005.t2 14.294
R942 a_3461_1005.n0 a_3461_1005.t0 14.282
R943 a_185_182.n1 a_185_182.t5 480.392
R944 a_185_182.n1 a_185_182.t3 403.272
R945 a_185_182.n2 a_185_182.t4 293.527
R946 a_185_182.n5 a_185_182.n3 221.779
R947 a_185_182.n3 a_185_182.n2 153.315
R948 a_185_182.n3 a_185_182.n0 140.59
R949 a_185_182.n2 a_185_182.n1 81.941
R950 a_185_182.n5 a_185_182.n4 15.218
R951 a_185_182.n0 a_185_182.t1 14.282
R952 a_185_182.n0 a_185_182.t0 14.282
R953 a_185_182.n6 a_185_182.n5 12.014
C4 VPB VNB 16.40fF
C5 a_185_182.n0 VNB 0.68fF
C6 a_185_182.n1 VNB 0.35fF
C7 a_185_182.n2 VNB 0.55fF
C8 a_185_182.n3 VNB 0.60fF
C9 a_185_182.n4 VNB 0.08fF
C10 a_185_182.n5 VNB 0.28fF
C11 a_185_182.n6 VNB 0.04fF
C12 a_3461_1005.n0 VNB 0.52fF
C13 a_3007_383.n0 VNB 0.74fF
C14 a_3007_383.n1 VNB 0.36fF
C15 a_3007_383.n2 VNB 0.84fF
C16 a_3007_383.n3 VNB 0.84fF
C17 a_3007_383.n4 VNB 0.05fF
C18 a_3007_383.n5 VNB 0.06fF
C19 a_3007_383.n6 VNB 0.22fF
C20 a_3007_383.n7 VNB 0.51fF
C21 a_3007_383.n8 VNB 0.09fF
C22 a_3007_383.n9 VNB 0.09fF
C23 a_3007_383.n10 VNB 0.05fF
C24 a_2405_182.n0 VNB 0.82fF
C25 a_2405_182.n1 VNB 0.35fF
C26 a_2405_182.t3 VNB 0.70fF
C27 a_2405_182.n2 VNB 1.08fF
C28 a_2405_182.n3 VNB 1.16fF
C29 a_2405_182.n4 VNB 0.10fF
C30 a_2405_182.n5 VNB 0.39fF
C31 a_2405_182.n6 VNB 0.06fF
C32 a_1666_73.n0 VNB 0.05fF
C33 a_1666_73.n1 VNB 0.02fF
C34 a_1666_73.n2 VNB 0.12fF
C35 a_1666_73.n3 VNB 0.04fF
C36 a_1666_73.n4 VNB 0.17fF
C37 a_1771_1004.n0 VNB 0.04fF
C38 a_1771_1004.n1 VNB 0.47fF
C39 a_1771_1004.n2 VNB 0.56fF
C40 a_1771_1004.n3 VNB 0.28fF
C41 a_1771_1004.n4 VNB 0.32fF
C42 a_1771_1004.t6 VNB 0.46fF
C43 a_1771_1004.n5 VNB 0.51fF
C44 a_1771_1004.n6 VNB 0.51fF
C45 a_1771_1004.n7 VNB 0.03fF
C46 a_1771_1004.n8 VNB 0.25fF
C47 a_1771_1004.n9 VNB 0.05fF
C48 a_2795_1005.n0 VNB 0.55fF
C49 a_1295_182.n0 VNB 0.05fF
C50 a_1295_182.n1 VNB 0.87fF
C51 a_1295_182.n2 VNB 0.41fF
C52 a_1295_182.n3 VNB 1.27fF
C53 a_1295_182.n4 VNB 1.31fF
C54 a_1295_182.n5 VNB 0.04fF
C55 a_1295_182.n6 VNB 0.37fF
C56 a_1295_182.n7 VNB 0.07fF
C57 VPB.n0 VNB 0.03fF
C58 VPB.n1 VNB 0.04fF
C59 VPB.n2 VNB 0.02fF
C60 VPB.n3 VNB 0.10fF
C61 VPB.n5 VNB 0.02fF
C62 VPB.n6 VNB 0.02fF
C63 VPB.n7 VNB 0.02fF
C64 VPB.n8 VNB 0.02fF
C65 VPB.n10 VNB 0.02fF
C66 VPB.n11 VNB 0.02fF
C67 VPB.n12 VNB 0.02fF
C68 VPB.n14 VNB 0.02fF
C69 VPB.n15 VNB 0.02fF
C70 VPB.n16 VNB 0.02fF
C71 VPB.n17 VNB 0.04fF
C72 VPB.n18 VNB 0.02fF
C73 VPB.n19 VNB 0.16fF
C74 VPB.n20 VNB 0.04fF
C75 VPB.n22 VNB 0.02fF
C76 VPB.n23 VNB 0.02fF
C77 VPB.n24 VNB 0.02fF
C78 VPB.n25 VNB 0.02fF
C79 VPB.n27 VNB 0.02fF
C80 VPB.n28 VNB 0.02fF
C81 VPB.n29 VNB 0.02fF
C82 VPB.n31 VNB 0.27fF
C83 VPB.n33 VNB 0.03fF
C84 VPB.n34 VNB 0.02fF
C85 VPB.n35 VNB 0.10fF
C86 VPB.n36 VNB 0.13fF
C87 VPB.n37 VNB 0.16fF
C88 VPB.n38 VNB 0.02fF
C89 VPB.n39 VNB 0.02fF
C90 VPB.n40 VNB 0.13fF
C91 VPB.n41 VNB 0.15fF
C92 VPB.n42 VNB 0.02fF
C93 VPB.n43 VNB 0.02fF
C94 VPB.n44 VNB 0.02fF
C95 VPB.n45 VNB 0.13fF
C96 VPB.n46 VNB 0.15fF
C97 VPB.n47 VNB 0.02fF
C98 VPB.n48 VNB 0.02fF
C99 VPB.n49 VNB 0.13fF
C100 VPB.n50 VNB 0.16fF
C101 VPB.n51 VNB 0.02fF
C102 VPB.n52 VNB 0.02fF
C103 VPB.n53 VNB 0.06fF
C104 VPB.n54 VNB 0.23fF
C105 VPB.n55 VNB 0.02fF
C106 VPB.n56 VNB 0.01fF
C107 VPB.n57 VNB 0.27fF
C108 VPB.n58 VNB 0.01fF
C109 VPB.n59 VNB 0.02fF
C110 VPB.n60 VNB 0.03fF
C111 VPB.n61 VNB 0.03fF
C112 VPB.n62 VNB 0.27fF
C113 VPB.n63 VNB 0.01fF
C114 VPB.n64 VNB 0.02fF
C115 VPB.n65 VNB 0.06fF
C116 VPB.n66 VNB 0.13fF
C117 VPB.n67 VNB 0.19fF
C118 VPB.n68 VNB 0.02fF
C119 VPB.n69 VNB 0.01fF
C120 VPB.n70 VNB 0.16fF
C121 VPB.n71 VNB 0.02fF
C122 VPB.n72 VNB 0.02fF
C123 VPB.n73 VNB 0.13fF
C124 VPB.n74 VNB 0.19fF
C125 VPB.n75 VNB 0.02fF
C126 VPB.n76 VNB 0.01fF
C127 VPB.n77 VNB 0.06fF
C128 VPB.n78 VNB 0.02fF
C129 VPB.n79 VNB 0.02fF
C130 VPB.n80 VNB 0.02fF
C131 VPB.n81 VNB 0.02fF
C132 VPB.n82 VNB 0.04fF
C133 VPB.n83 VNB 0.02fF
C134 VPB.n84 VNB 0.16fF
C135 VPB.n85 VNB 0.04fF
C136 VPB.n87 VNB 0.02fF
C137 VPB.n88 VNB 0.02fF
C138 VPB.n89 VNB 0.02fF
C139 VPB.n90 VNB 0.02fF
C140 VPB.n92 VNB 0.02fF
C141 VPB.n93 VNB 0.02fF
C142 VPB.n94 VNB 0.02fF
C143 VPB.n96 VNB 0.27fF
C144 VPB.n98 VNB 0.03fF
C145 VPB.n99 VNB 0.02fF
C146 VPB.n100 VNB 0.02fF
C147 VPB.n101 VNB 0.02fF
C148 VPB.n102 VNB 0.02fF
C149 VPB.n103 VNB 0.04fF
C150 VPB.n104 VNB 0.02fF
C151 VPB.n105 VNB 0.16fF
C152 VPB.n106 VNB 0.04fF
C153 VPB.n108 VNB 0.02fF
C154 VPB.n109 VNB 0.02fF
C155 VPB.n110 VNB 0.02fF
C156 VPB.n111 VNB 0.02fF
C157 VPB.n113 VNB 0.02fF
C158 VPB.n114 VNB 0.02fF
C159 VPB.n115 VNB 0.02fF
C160 VPB.n117 VNB 0.27fF
C161 VPB.n119 VNB 0.03fF
C162 VPB.n120 VNB 0.02fF
C163 VPB.n121 VNB 0.10fF
C164 VPB.n122 VNB 0.02fF
C165 VPB.n123 VNB 0.13fF
C166 VPB.n124 VNB 0.16fF
C167 VPB.n125 VNB 0.02fF
C168 VPB.n126 VNB 0.02fF
C169 VPB.n127 VNB 0.23fF
C170 VPB.n128 VNB 0.02fF
C171 VPB.n129 VNB 0.02fF
C172 VPB.n130 VNB 0.27fF
C173 VPB.n131 VNB 0.01fF
C174 VPB.n132 VNB 0.02fF
C175 VPB.n133 VNB 0.03fF
C176 VPB.n134 VNB 0.03fF
C177 VPB.n135 VNB 0.27fF
C178 VPB.n136 VNB 0.01fF
C179 VPB.n137 VNB 0.02fF
C180 VPB.n138 VNB 0.06fF
C181 VPB.n139 VNB 0.13fF
C182 VPB.n140 VNB 0.19fF
C183 VPB.n141 VNB 0.02fF
C184 VPB.n142 VNB 0.01fF
C185 VPB.n143 VNB 0.16fF
C186 VPB.n144 VNB 0.02fF
C187 VPB.n145 VNB 0.02fF
C188 VPB.n146 VNB 0.13fF
C189 VPB.n147 VNB 0.19fF
C190 VPB.n148 VNB 0.02fF
C191 VPB.n149 VNB 0.01fF
C192 VPB.n150 VNB 0.06fF
C193 VPB.n151 VNB 0.27fF
C194 VPB.n152 VNB 0.01fF
C195 VPB.n153 VNB 0.02fF
C196 VPB.n154 VNB 0.03fF
C197 VPB.n155 VNB 0.03fF
C198 VPB.n156 VNB 0.27fF
C199 VPB.n157 VNB 0.01fF
C200 VPB.n158 VNB 0.02fF
C201 VPB.n159 VNB 0.02fF
C202 VPB.n160 VNB 0.02fF
C203 VPB.n161 VNB 0.02fF
C204 VPB.n162 VNB 0.14fF
C205 VPB.n163 VNB 0.03fF
C206 VPB.n164 VNB 0.02fF
C207 VPB.n165 VNB 0.05fF
C208 VPB.n166 VNB 0.01fF
C209 VPB.n168 VNB 0.02fF
C210 VPB.n169 VNB 0.02fF
C211 VPB.n171 VNB 0.02fF
C212 VPB.n172 VNB 0.02fF
C213 VPB.n173 VNB 0.02fF
C214 VPB.n176 VNB 0.45fF
C215 VPB.n178 VNB 0.04fF
C216 VPB.n179 VNB 0.04fF
C217 VPB.n180 VNB 0.27fF
C218 VPB.n181 VNB 0.03fF
C219 VPB.n182 VNB 0.03fF
C220 VPB.n183 VNB 0.27fF
C221 VPB.n184 VNB 0.02fF
C222 VPB.n185 VNB 0.02fF
C223 VPB.n186 VNB 0.27fF
C224 VPB.n187 VNB 0.02fF
C225 VPB.n188 VNB 0.02fF
C226 VPB.n189 VNB 0.27fF
C227 VPB.n190 VNB 0.02fF
C228 VPB.n191 VNB 0.02fF
C229 VPB.n192 VNB 0.00fF
C230 VPB.n193 VNB 0.09fF
C231 VPB.n194 VNB 0.02fF
C232 VPB.n195 VNB 0.13fF
C233 VPB.n196 VNB 0.15fF
C234 VPB.n197 VNB 0.02fF
C235 VPB.n198 VNB 0.02fF
C236 VPB.n199 VNB 0.02fF
C237 VPB.n200 VNB 0.10fF
C238 VPB.n201 VNB 0.02fF
C239 VPB.n202 VNB 0.13fF
C240 VPB.n203 VNB 0.16fF
C241 VPB.n204 VNB 0.02fF
C242 VPB.n205 VNB 0.02fF
C243 VPB.n206 VNB 0.02fF
C244 VPB.n207 VNB 0.23fF
C245 VPB.n208 VNB 0.02fF
C246 VPB.n209 VNB 0.02fF
C247 VPB.n210 VNB 0.02fF
C248 VPB.n211 VNB 0.27fF
C249 VPB.n212 VNB 0.01fF
C250 VPB.n213 VNB 0.02fF
C251 VPB.n214 VNB 0.04fF
C252 VPB.n215 VNB 0.02fF
C253 VPB.n216 VNB 0.02fF
C254 VPB.n217 VNB 0.02fF
C255 VPB.n218 VNB 0.04fF
C256 VPB.n219 VNB 0.02fF
C257 VPB.n220 VNB 0.20fF
C258 VPB.n221 VNB 0.04fF
C259 VPB.n223 VNB 0.02fF
C260 VPB.n224 VNB 0.02fF
C261 VPB.n225 VNB 0.02fF
C262 VPB.n226 VNB 0.02fF
C263 VPB.n228 VNB 0.02fF
C264 VPB.n229 VNB 0.02fF
C265 VPB.n230 VNB 0.02fF
C266 VPB.n232 VNB 0.27fF
C267 VPB.n234 VNB 0.03fF
C268 VPB.n235 VNB 0.02fF
C269 VPB.n236 VNB 0.03fF
C270 VPB.n237 VNB 0.03fF
C271 VPB.n238 VNB 0.27fF
C272 VPB.n239 VNB 0.01fF
C273 VPB.n240 VNB 0.02fF
C274 VPB.n241 VNB 0.04fF
C275 VPB.n242 VNB 0.27fF
C276 VPB.n243 VNB 0.02fF
C277 VPB.n244 VNB 0.02fF
C278 VPB.n245 VNB 0.02fF
C279 VPB.n246 VNB 0.27fF
C280 VPB.n247 VNB 0.02fF
C281 VPB.n248 VNB 0.02fF
C282 VPB.n249 VNB 0.02fF
C283 VPB.n250 VNB 0.27fF
C284 VPB.n251 VNB 0.02fF
C285 VPB.n252 VNB 0.02fF
C286 VPB.n253 VNB 0.02fF
C287 VPB.n254 VNB 0.13fF
C288 VPB.n255 VNB 0.15fF
C289 VPB.n256 VNB 0.02fF
C290 VPB.n257 VNB 0.02fF
C291 VPB.n258 VNB 0.02fF
C292 VPB.n259 VNB 0.02fF
C293 VPB.n260 VNB 0.02fF
C294 VPB.n261 VNB 0.04fF
C295 VPB.n262 VNB 0.04fF
C296 VPB.n263 VNB 0.02fF
C297 VPB.n264 VNB 0.02fF
C298 VPB.n265 VNB 0.02fF
C299 VPB.n266 VNB 0.04fF
C300 VPB.n267 VNB 0.04fF
C301 VPB.n268 VNB 0.02fF
C302 VPB.n269 VNB 0.23fF
C303 VPB.n270 VNB 0.02fF
C304 VPB.n271 VNB 0.01fF
C305 VPB.n272 VNB 0.05fF
C306 VPB.n273 VNB 0.13fF
C307 VPB.n274 VNB 0.16fF
C308 VPB.n275 VNB 0.02fF
C309 VPB.n276 VNB 0.02fF
C310 VPB.n277 VNB 0.10fF
C311 VPB.n278 VNB 0.02fF
C312 VPB.n279 VNB 0.13fF
C313 VPB.n280 VNB 0.15fF
C314 VPB.n281 VNB 0.02fF
C315 VPB.n282 VNB 0.02fF
C316 VPB.n283 VNB 0.02fF
C317 VPB.n284 VNB 0.13fF
C318 VPB.n285 VNB 0.15fF
C319 VPB.n286 VNB 0.02fF
C320 VPB.n287 VNB 0.02fF
C321 VPB.n288 VNB 0.02fF
C322 VPB.n289 VNB 0.13fF
C323 VPB.n290 VNB 0.16fF
C324 VPB.n291 VNB 0.02fF
C325 VPB.n292 VNB 0.02fF
C326 VPB.n293 VNB 0.02fF
C327 VPB.n294 VNB 0.06fF
C328 VPB.n295 VNB 0.23fF
C329 VPB.n296 VNB 0.02fF
C330 VPB.n297 VNB 0.01fF
C331 VPB.n298 VNB 0.02fF
C332 VPB.n299 VNB 0.27fF
C333 VPB.n300 VNB 0.01fF
C334 VPB.n301 VNB 0.02fF
C335 VPB.n302 VNB 0.04fF
C336 VPB.n303 VNB 0.02fF
C337 VPB.n304 VNB 0.02fF
C338 VPB.n305 VNB 0.02fF
C339 VPB.n306 VNB 0.04fF
C340 VPB.n307 VNB 0.02fF
C341 VPB.n308 VNB 0.16fF
C342 VPB.n309 VNB 0.04fF
C343 VPB.n311 VNB 0.02fF
C344 VPB.n312 VNB 0.02fF
C345 VPB.n313 VNB 0.02fF
C346 VPB.n314 VNB 0.02fF
C347 VPB.n316 VNB 0.02fF
C348 VPB.n317 VNB 0.02fF
C349 VPB.n318 VNB 0.02fF
C350 VPB.n320 VNB 0.27fF
C351 VPB.n322 VNB 0.03fF
C352 VPB.n323 VNB 0.02fF
C353 VPB.n324 VNB 0.03fF
C354 VPB.n325 VNB 0.03fF
C355 VPB.n326 VNB 0.27fF
C356 VPB.n327 VNB 0.01fF
C357 VPB.n328 VNB 0.02fF
C358 VPB.n329 VNB 0.04fF
C359 VPB.n330 VNB 0.06fF
C360 VPB.n331 VNB 0.13fF
C361 VPB.n332 VNB 0.19fF
C362 VPB.n333 VNB 0.02fF
C363 VPB.n334 VNB 0.01fF
C364 VPB.n335 VNB 0.02fF
C365 VPB.n336 VNB 0.16fF
C366 VPB.n337 VNB 0.02fF
C367 VPB.n338 VNB 0.02fF
C368 VPB.n339 VNB 0.02fF
C369 VPB.n340 VNB 0.06fF
C370 VPB.n341 VNB 0.13fF
C371 VPB.n342 VNB 0.19fF
C372 VPB.n343 VNB 0.02fF
C373 VPB.n344 VNB 0.01fF
C374 VPB.n345 VNB 0.02fF
C375 VPB.n346 VNB 0.27fF
C376 VPB.n347 VNB 0.01fF
C377 VPB.n348 VNB 0.02fF
C378 VPB.n349 VNB 0.04fF
C379 VPB.n350 VNB 0.02fF
C380 VPB.n351 VNB 0.02fF
C381 VPB.n352 VNB 0.02fF
C382 VPB.n353 VNB 0.04fF
C383 VPB.n354 VNB 0.02fF
C384 VPB.n355 VNB 0.16fF
C385 VPB.n356 VNB 0.04fF
C386 VPB.n358 VNB 0.02fF
C387 VPB.n359 VNB 0.02fF
C388 VPB.n360 VNB 0.02fF
C389 VPB.n361 VNB 0.02fF
C390 VPB.n363 VNB 0.02fF
C391 VPB.n364 VNB 0.02fF
C392 VPB.n365 VNB 0.02fF
C393 VPB.n367 VNB 0.27fF
C394 VPB.n369 VNB 0.03fF
C395 VPB.n370 VNB 0.02fF
C396 VPB.n371 VNB 0.03fF
C397 VPB.n372 VNB 0.03fF
C398 VPB.n373 VNB 0.27fF
C399 VPB.n374 VNB 0.01fF
C400 VPB.n375 VNB 0.02fF
C401 VPB.n376 VNB 0.04fF
C402 VPB.n377 VNB 0.05fF
C403 VPB.n378 VNB 0.23fF
C404 VPB.n379 VNB 0.02fF
C405 VPB.n380 VNB 0.01fF
C406 VPB.n381 VNB 0.02fF
C407 VPB.n382 VNB 0.02fF
C408 VPB.n383 VNB 0.02fF
C409 VPB.n384 VNB 0.02fF
C410 VPB.n385 VNB 0.02fF
C411 VPB.n386 VNB 0.02fF
C412 VPB.n387 VNB 0.04fF
C413 VPB.n388 VNB 0.04fF
C414 VPB.n389 VNB 0.02fF
C415 VPB.n390 VNB 0.02fF
C416 VPB.n391 VNB 0.02fF
C417 VPB.n392 VNB 0.03fF
C418 VPB.n393 VNB 0.03fF
C419 VPB.n394 VNB 0.02fF
C420 VPB.n395 VNB 0.02fF
C421 VPB.n396 VNB 0.02fF
C422 VPB.n397 VNB 0.04fF
C423 VPB.n398 VNB 0.04fF
C424 VPB.n400 VNB 0.42fF
C425 a_661_1004.n0 VNB 0.05fF
C426 a_661_1004.n1 VNB 0.50fF
C427 a_661_1004.n2 VNB 0.59fF
C428 a_661_1004.n3 VNB 0.30fF
C429 a_661_1004.n4 VNB 0.33fF
C430 a_661_1004.t6 VNB 0.49fF
C431 a_661_1004.n5 VNB 0.54fF
C432 a_661_1004.n6 VNB 0.53fF
C433 a_661_1004.n7 VNB 0.02fF
C434 a_661_1004.n8 VNB 0.26fF
C435 a_661_1004.n9 VNB 0.04fF
C436 a_556_73.n0 VNB 0.05fF
C437 a_556_73.n1 VNB 0.02fF
C438 a_556_73.n2 VNB 0.12fF
C439 a_556_73.n3 VNB 0.04fF
C440 a_556_73.n4 VNB 0.17fF
.ends
