// File: OR2X1.spi.OR2X1.pxi
// Created: Tue Oct 15 15:50:42 2024
// 
simulator lang=spectre
x_PM_OR2X1\%GND ( GND N_GND_c_4_p N_GND_c_48_p N_GND_c_13_p N_GND_c_14_p \
 N_GND_c_17_p N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p N_GND_c_31_p N_GND_c_2_p \
 N_GND_c_1_p N_GND_c_3_p N_GND_M0_noxref_s N_GND_M2_noxref_s )  PM_OR2X1\%GND
x_PM_OR2X1\%VDD ( VDD N_VDD_c_78_p N_VDD_c_106_p N_VDD_c_75_n N_VDD_c_83_p \
 N_VDD_c_91_p N_VDD_c_76_n N_VDD_c_77_n N_VDD_M3_noxref_d N_VDD_M7_noxref_s \
 N_VDD_M8_noxref_d )  PM_OR2X1\%VDD
x_PM_OR2X1\%noxref_3 ( N_noxref_3_c_147_n N_noxref_3_c_153_n \
 N_noxref_3_c_155_n N_noxref_3_c_214_p N_noxref_3_c_194_n N_noxref_3_c_196_n \
 N_noxref_3_c_159_n N_noxref_3_c_164_n N_noxref_3_c_165_n \
 N_noxref_3_M2_noxref_g N_noxref_3_M7_noxref_g N_noxref_3_M8_noxref_g \
 N_noxref_3_c_170_n N_noxref_3_c_271_p N_noxref_3_c_272_p N_noxref_3_c_172_n \
 N_noxref_3_c_208_n N_noxref_3_c_209_n N_noxref_3_c_173_n N_noxref_3_c_263_p \
 N_noxref_3_c_174_n N_noxref_3_c_176_n N_noxref_3_c_177_n \
 N_noxref_3_M0_noxref_d N_noxref_3_M1_noxref_d N_noxref_3_M5_noxref_d )  \
 PM_OR2X1\%noxref_3
x_PM_OR2X1\%A ( A A A A A A A N_A_c_283_n N_A_c_295_n N_A_M0_noxref_g \
 N_A_M3_noxref_g N_A_M4_noxref_g N_A_c_286_n N_A_c_307_n N_A_c_308_n \
 N_A_c_288_n N_A_c_290_n N_A_c_312_n N_A_c_317_p N_A_c_291_n N_A_c_293_n \
 N_A_c_303_n )  PM_OR2X1\%A
x_PM_OR2X1\%B ( B B B B B B B N_B_c_362_n N_B_c_349_n N_B_M1_noxref_g \
 N_B_M5_noxref_g N_B_M6_noxref_g N_B_c_351_n N_B_c_371_n N_B_c_372_n \
 N_B_c_375_n N_B_c_353_n N_B_c_354_n N_B_c_355_n N_B_c_381_n N_B_c_382_n \
 N_B_c_384_n N_B_c_387_n )  PM_OR2X1\%B
x_PM_OR2X1\%noxref_6 ( N_noxref_6_c_418_n N_noxref_6_c_423_n \
 N_noxref_6_c_424_n N_noxref_6_c_425_n N_noxref_6_M3_noxref_s \
 N_noxref_6_M4_noxref_d N_noxref_6_M6_noxref_d )  PM_OR2X1\%noxref_6
x_PM_OR2X1\%Y ( Y Y Y Y Y Y Y N_Y_c_460_n N_Y_c_484_n N_Y_c_470_n N_Y_c_473_n \
 N_Y_M2_noxref_d N_Y_M7_noxref_d )  PM_OR2X1\%Y
cc_1 ( N_GND_c_1_p N_VDD_c_75_n ) capacitor c=0.00989031f //x=0.695 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_76_n ) capacitor c=0.00989031f //x=5.18 //y=0 \
 //x2=5.18 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_77_n ) capacitor c=0.00855708f //x=3.33 //y=0 \
 //x2=3.33 //y2=7.4
cc_4 ( N_GND_c_4_p N_noxref_3_c_147_n ) capacitor c=0.0116078f //x=5.18 //y=0 \
 //x2=3.955 //y2=3.33
cc_5 ( N_GND_c_5_p N_noxref_3_c_147_n ) capacitor c=0.00136402f //x=3.16 //y=0 \
 //x2=3.955 //y2=3.33
cc_6 ( N_GND_c_6_p N_noxref_3_c_147_n ) capacitor c=0.00110325f //x=3.875 \
 //y=0 //x2=3.955 //y2=3.33
cc_7 ( N_GND_c_7_p N_noxref_3_c_147_n ) capacitor c=2.76195e-19 //x=4.36 \
 //y=0.535 //x2=3.955 //y2=3.33
cc_8 ( N_GND_c_3_p N_noxref_3_c_147_n ) capacitor c=0.00820844f //x=3.33 //y=0 \
 //x2=3.955 //y2=3.33
cc_9 ( N_GND_M2_noxref_s N_noxref_3_c_147_n ) capacitor c=0.00164577f \
 //x=3.825 //y=0.37 //x2=3.955 //y2=3.33
cc_10 ( N_GND_c_4_p N_noxref_3_c_153_n ) capacitor c=0.00192312f //x=5.18 \
 //y=0 //x2=2.705 //y2=3.33
cc_11 ( N_GND_M0_noxref_s N_noxref_3_c_153_n ) capacitor c=6.50479e-19 \
 //x=0.56 //y=0.365 //x2=2.705 //y2=3.33
cc_12 ( N_GND_c_4_p N_noxref_3_c_155_n ) capacitor c=0.00359057f //x=5.18 \
 //y=0 //x2=2.065 //y2=1.655
cc_13 ( N_GND_c_13_p N_noxref_3_c_155_n ) capacitor c=0.00381844f //x=1.58 \
 //y=0.53 //x2=2.065 //y2=1.655
cc_14 ( N_GND_c_14_p N_noxref_3_c_155_n ) capacitor c=0.00323369f //x=2.065 \
 //y=0.53 //x2=2.065 //y2=1.655
cc_15 ( N_GND_M0_noxref_s N_noxref_3_c_155_n ) capacitor c=0.0173679f //x=0.56 \
 //y=0.365 //x2=2.065 //y2=1.655
cc_16 ( N_GND_c_4_p N_noxref_3_c_159_n ) capacitor c=0.00197099f //x=5.18 \
 //y=0 //x2=2.505 //y2=1.655
cc_17 ( N_GND_c_17_p N_noxref_3_c_159_n ) capacitor c=0.00479136f //x=2.55 \
 //y=0.53 //x2=2.505 //y2=1.655
cc_18 ( N_GND_c_3_p N_noxref_3_c_159_n ) capacitor c=0.0464456f //x=3.33 //y=0 \
 //x2=2.505 //y2=1.655
cc_19 ( N_GND_M0_noxref_s N_noxref_3_c_159_n ) capacitor c=0.0158743f //x=0.56 \
 //y=0.365 //x2=2.505 //y2=1.655
cc_20 ( N_GND_M2_noxref_s N_noxref_3_c_159_n ) capacitor c=3.53679e-19 \
 //x=3.825 //y=0.37 //x2=2.505 //y2=1.655
cc_21 ( N_GND_c_1_p N_noxref_3_c_164_n ) capacitor c=0.00101801f //x=0.695 \
 //y=0 //x2=2.59 //y2=3.33
cc_22 ( N_GND_c_4_p N_noxref_3_c_165_n ) capacitor c=0.00184963f //x=5.18 \
 //y=0 //x2=4.07 //y2=2.085
cc_23 ( N_GND_c_7_p N_noxref_3_c_165_n ) capacitor c=7.87839e-19 //x=4.36 \
 //y=0.535 //x2=4.07 //y2=2.085
cc_24 ( N_GND_c_2_p N_noxref_3_c_165_n ) capacitor c=0.00118981f //x=5.18 \
 //y=0 //x2=4.07 //y2=2.085
cc_25 ( N_GND_c_3_p N_noxref_3_c_165_n ) capacitor c=0.029021f //x=3.33 //y=0 \
 //x2=4.07 //y2=2.085
cc_26 ( N_GND_M2_noxref_s N_noxref_3_c_165_n ) capacitor c=0.0108503f \
 //x=3.825 //y=0.37 //x2=4.07 //y2=2.085
cc_27 ( N_GND_c_7_p N_noxref_3_c_170_n ) capacitor c=0.0121757f //x=4.36 \
 //y=0.535 //x2=4.18 //y2=0.91
cc_28 ( N_GND_M2_noxref_s N_noxref_3_c_170_n ) capacitor c=0.0317181f \
 //x=3.825 //y=0.37 //x2=4.18 //y2=0.91
cc_29 ( N_GND_c_3_p N_noxref_3_c_172_n ) capacitor c=0.00552709f //x=3.33 \
 //y=0 //x2=4.18 //y2=1.92
cc_30 ( N_GND_M2_noxref_s N_noxref_3_c_173_n ) capacitor c=0.00483274f \
 //x=3.825 //y=0.37 //x2=4.555 //y2=0.755
cc_31 ( N_GND_c_31_p N_noxref_3_c_174_n ) capacitor c=0.0118602f //x=4.845 \
 //y=0.535 //x2=4.71 //y2=0.91
cc_32 ( N_GND_M2_noxref_s N_noxref_3_c_174_n ) capacitor c=0.0143355f \
 //x=3.825 //y=0.37 //x2=4.71 //y2=0.91
cc_33 ( N_GND_M2_noxref_s N_noxref_3_c_176_n ) capacitor c=0.0074042f \
 //x=3.825 //y=0.37 //x2=4.71 //y2=1.255
cc_34 ( N_GND_c_7_p N_noxref_3_c_177_n ) capacitor c=2.1838e-19 //x=4.36 \
 //y=0.535 //x2=4.07 //y2=2.085
cc_35 ( N_GND_c_3_p N_noxref_3_c_177_n ) capacitor c=0.0108179f //x=3.33 //y=0 \
 //x2=4.07 //y2=2.085
cc_36 ( N_GND_M2_noxref_s N_noxref_3_c_177_n ) capacitor c=0.00655738f \
 //x=3.825 //y=0.37 //x2=4.07 //y2=2.085
cc_37 ( N_GND_c_4_p N_noxref_3_M0_noxref_d ) capacitor c=0.00175924f //x=5.18 \
 //y=0 //x2=0.99 //y2=0.905
cc_38 ( N_GND_c_2_p N_noxref_3_M0_noxref_d ) capacitor c=2.31043e-19 //x=5.18 \
 //y=0 //x2=0.99 //y2=0.905
cc_39 ( N_GND_c_1_p N_noxref_3_M0_noxref_d ) capacitor c=0.00416273f //x=0.695 \
 //y=0 //x2=0.99 //y2=0.905
cc_40 ( N_GND_c_3_p N_noxref_3_M0_noxref_d ) capacitor c=2.57516e-19 //x=3.33 \
 //y=0 //x2=0.99 //y2=0.905
cc_41 ( N_GND_M0_noxref_s N_noxref_3_M0_noxref_d ) capacitor c=0.0770866f \
 //x=0.56 //y=0.365 //x2=0.99 //y2=0.905
cc_42 ( N_GND_c_4_p N_noxref_3_M1_noxref_d ) capacitor c=0.00195394f //x=5.18 \
 //y=0 //x2=1.96 //y2=0.905
cc_43 ( N_GND_c_2_p N_noxref_3_M1_noxref_d ) capacitor c=2.31043e-19 //x=5.18 \
 //y=0 //x2=1.96 //y2=0.905
cc_44 ( N_GND_c_3_p N_noxref_3_M1_noxref_d ) capacitor c=0.00609243f //x=3.33 \
 //y=0 //x2=1.96 //y2=0.905
cc_45 ( N_GND_M0_noxref_s N_noxref_3_M1_noxref_d ) capacitor c=0.0610175f \
 //x=0.56 //y=0.365 //x2=1.96 //y2=0.905
cc_46 ( N_GND_M2_noxref_s N_noxref_3_M1_noxref_d ) capacitor c=2.04477e-19 \
 //x=3.825 //y=0.37 //x2=1.96 //y2=0.905
cc_47 ( N_GND_c_4_p N_A_c_283_n ) capacitor c=6.7762e-19 //x=5.18 //y=0 \
 //x2=1.11 //y2=2.08
cc_48 ( N_GND_c_48_p N_A_c_283_n ) capacitor c=0.00136072f //x=1.095 //y=0.53 \
 //x2=1.11 //y2=2.08
cc_49 ( N_GND_c_1_p N_A_c_283_n ) capacitor c=0.0176887f //x=0.695 //y=0 \
 //x2=1.11 //y2=2.08
cc_50 ( N_GND_c_48_p N_A_c_286_n ) capacitor c=0.0122371f //x=1.095 //y=0.53 \
 //x2=0.915 //y2=0.905
cc_51 ( N_GND_M0_noxref_s N_A_c_286_n ) capacitor c=0.0318086f //x=0.56 \
 //y=0.365 //x2=0.915 //y2=0.905
cc_52 ( N_GND_c_48_p N_A_c_288_n ) capacitor c=2.1838e-19 //x=1.095 //y=0.53 \
 //x2=0.915 //y2=1.915
cc_53 ( N_GND_c_1_p N_A_c_288_n ) capacitor c=0.0196165f //x=0.695 //y=0 \
 //x2=0.915 //y2=1.915
cc_54 ( N_GND_M0_noxref_s N_A_c_290_n ) capacitor c=0.00474433f //x=0.56 \
 //y=0.365 //x2=1.29 //y2=0.75
cc_55 ( N_GND_c_13_p N_A_c_291_n ) capacitor c=0.0113089f //x=1.58 //y=0.53 \
 //x2=1.445 //y2=0.905
cc_56 ( N_GND_M0_noxref_s N_A_c_291_n ) capacitor c=0.00514143f //x=0.56 \
 //y=0.365 //x2=1.445 //y2=0.905
cc_57 ( N_GND_M0_noxref_s N_A_c_293_n ) capacitor c=8.33128e-19 //x=0.56 \
 //y=0.365 //x2=1.445 //y2=1.25
cc_58 ( N_GND_c_1_p N_B_c_349_n ) capacitor c=9.2064e-19 //x=0.695 //y=0 \
 //x2=1.85 //y2=2.08
cc_59 ( N_GND_c_3_p N_B_c_349_n ) capacitor c=9.53263e-19 //x=3.33 //y=0 \
 //x2=1.85 //y2=2.08
cc_60 ( N_GND_c_14_p N_B_c_351_n ) capacitor c=0.0109802f //x=2.065 //y=0.53 \
 //x2=1.885 //y2=0.905
cc_61 ( N_GND_M0_noxref_s N_B_c_351_n ) capacitor c=0.00590563f //x=0.56 \
 //y=0.365 //x2=1.885 //y2=0.905
cc_62 ( N_GND_M0_noxref_s N_B_c_353_n ) capacitor c=0.00466751f //x=0.56 \
 //y=0.365 //x2=2.26 //y2=0.75
cc_63 ( N_GND_M0_noxref_s N_B_c_354_n ) capacitor c=0.00316186f //x=0.56 \
 //y=0.365 //x2=2.26 //y2=1.405
cc_64 ( N_GND_c_17_p N_B_c_355_n ) capacitor c=0.0112321f //x=2.55 //y=0.53 \
 //x2=2.415 //y2=0.905
cc_65 ( N_GND_M0_noxref_s N_B_c_355_n ) capacitor c=0.0142835f //x=0.56 \
 //y=0.365 //x2=2.415 //y2=0.905
cc_66 ( N_GND_c_3_p Y ) capacitor c=8.10282e-19 //x=3.33 //y=0 //x2=4.81 \
 //y2=2.22
cc_67 ( N_GND_c_4_p N_Y_c_460_n ) capacitor c=0.00180637f //x=5.18 //y=0 \
 //x2=4.725 //y2=2.08
cc_68 ( N_GND_c_2_p N_Y_c_460_n ) capacitor c=0.0301661f //x=5.18 //y=0 \
 //x2=4.725 //y2=2.08
cc_69 ( N_GND_M2_noxref_s N_Y_c_460_n ) capacitor c=0.00999304f //x=3.825 \
 //y=0.37 //x2=4.725 //y2=2.08
cc_70 ( N_GND_c_4_p N_Y_M2_noxref_d ) capacitor c=0.00194883f //x=5.18 //y=0 \
 //x2=4.255 //y2=0.91
cc_71 ( N_GND_c_7_p N_Y_M2_noxref_d ) capacitor c=0.0146043f //x=4.36 \
 //y=0.535 //x2=4.255 //y2=0.91
cc_72 ( N_GND_c_2_p N_Y_M2_noxref_d ) capacitor c=0.00973758f //x=5.18 //y=0 \
 //x2=4.255 //y2=0.91
cc_73 ( N_GND_c_3_p N_Y_M2_noxref_d ) capacitor c=0.00924905f //x=3.33 //y=0 \
 //x2=4.255 //y2=0.91
cc_74 ( N_GND_M2_noxref_s N_Y_M2_noxref_d ) capacitor c=0.076995f //x=3.825 \
 //y=0.37 //x2=4.255 //y2=0.91
cc_75 ( N_VDD_c_78_p N_noxref_3_c_147_n ) capacitor c=0.00920603f //x=5.18 \
 //y=7.4 //x2=3.955 //y2=3.33
cc_76 ( N_VDD_c_77_n N_noxref_3_c_147_n ) capacitor c=0.0069465f //x=3.33 \
 //y=7.4 //x2=3.955 //y2=3.33
cc_77 ( N_VDD_M7_noxref_s N_noxref_3_c_147_n ) capacitor c=0.00106085f \
 //x=3.87 //y=5.02 //x2=3.955 //y2=3.33
cc_78 ( N_VDD_c_78_p N_noxref_3_c_153_n ) capacitor c=0.0014539f //x=5.18 \
 //y=7.4 //x2=2.705 //y2=3.33
cc_79 ( N_VDD_c_78_p N_noxref_3_c_194_n ) capacitor c=0.00178185f //x=5.18 \
 //y=7.4 //x2=2.505 //y2=5.21
cc_80 ( N_VDD_c_83_p N_noxref_3_c_194_n ) capacitor c=0.00136949f //x=3.16 \
 //y=7.4 //x2=2.505 //y2=5.21
cc_81 ( N_VDD_c_75_n N_noxref_3_c_196_n ) capacitor c=8.9933e-19 //x=0.74 \
 //y=7.4 //x2=2.195 //y2=5.21
cc_82 ( N_VDD_c_75_n N_noxref_3_c_164_n ) capacitor c=0.00163766f //x=0.74 \
 //y=7.4 //x2=2.59 //y2=3.33
cc_83 ( N_VDD_c_77_n N_noxref_3_c_164_n ) capacitor c=0.0462234f //x=3.33 \
 //y=7.4 //x2=2.59 //y2=3.33
cc_84 ( N_VDD_c_78_p N_noxref_3_c_165_n ) capacitor c=0.00160122f //x=5.18 \
 //y=7.4 //x2=4.07 //y2=2.085
cc_85 ( N_VDD_c_76_n N_noxref_3_c_165_n ) capacitor c=0.00144809f //x=5.18 \
 //y=7.4 //x2=4.07 //y2=2.085
cc_86 ( N_VDD_c_77_n N_noxref_3_c_165_n ) capacitor c=0.0272885f //x=3.33 \
 //y=7.4 //x2=4.07 //y2=2.085
cc_87 ( N_VDD_M7_noxref_s N_noxref_3_c_165_n ) capacitor c=0.00971593f \
 //x=3.87 //y=5.02 //x2=4.07 //y2=2.085
cc_88 ( N_VDD_c_91_p N_noxref_3_M7_noxref_g ) capacitor c=0.00748034f //x=4.8 \
 //y=7.4 //x2=4.225 //y2=6.02
cc_89 ( N_VDD_c_77_n N_noxref_3_M7_noxref_g ) capacitor c=0.0102569f //x=3.33 \
 //y=7.4 //x2=4.225 //y2=6.02
cc_90 ( N_VDD_M7_noxref_s N_noxref_3_M7_noxref_g ) capacitor c=0.0528676f \
 //x=3.87 //y=5.02 //x2=4.225 //y2=6.02
cc_91 ( N_VDD_c_91_p N_noxref_3_M8_noxref_g ) capacitor c=0.00697478f //x=4.8 \
 //y=7.4 //x2=4.665 //y2=6.02
cc_92 ( N_VDD_M8_noxref_d N_noxref_3_M8_noxref_g ) capacitor c=0.0528676f \
 //x=4.74 //y=5.02 //x2=4.665 //y2=6.02
cc_93 ( N_VDD_c_76_n N_noxref_3_c_208_n ) capacitor c=0.0287802f //x=5.18 \
 //y=7.4 //x2=4.59 //y2=4.79
cc_94 ( N_VDD_c_77_n N_noxref_3_c_209_n ) capacitor c=0.011132f //x=3.33 \
 //y=7.4 //x2=4.3 //y2=4.79
cc_95 ( N_VDD_M7_noxref_s N_noxref_3_c_209_n ) capacitor c=0.00527247f \
 //x=3.87 //y=5.02 //x2=4.3 //y2=4.79
cc_96 ( N_VDD_c_77_n N_noxref_3_M5_noxref_d ) capacitor c=0.00966019f //x=3.33 \
 //y=7.4 //x2=1.965 //y2=5.025
cc_97 ( N_VDD_M3_noxref_d N_noxref_3_M5_noxref_d ) capacitor c=0.00561178f \
 //x=1.085 //y=5.025 //x2=1.965 //y2=5.025
cc_98 ( N_VDD_M7_noxref_s N_noxref_3_M5_noxref_d ) capacitor c=4.94992e-19 \
 //x=3.87 //y=5.02 //x2=1.965 //y2=5.025
cc_99 ( N_VDD_c_75_n N_A_c_283_n ) capacitor c=0.0104719f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_100 ( N_VDD_c_78_p N_A_c_295_n ) capacitor c=3.36335e-19 //x=5.18 //y=7.4 \
 //x2=0.955 //y2=4.705
cc_101 ( N_VDD_c_75_n N_A_c_295_n ) capacitor c=0.008636f //x=0.74 //y=7.4 \
 //x2=0.955 //y2=4.705
cc_102 ( N_VDD_M3_noxref_d N_A_c_295_n ) capacitor c=2.82936e-19 //x=1.085 \
 //y=5.025 //x2=0.955 //y2=4.705
cc_103 ( N_VDD_c_106_p N_A_M3_noxref_g ) capacitor c=0.0067918f //x=1.145 \
 //y=7.4 //x2=1.01 //y2=6.025
cc_104 ( N_VDD_c_75_n N_A_M3_noxref_g ) capacitor c=0.0237757f //x=0.74 \
 //y=7.4 //x2=1.01 //y2=6.025
cc_105 ( N_VDD_M3_noxref_d N_A_M3_noxref_g ) capacitor c=0.0156786f //x=1.085 \
 //y=5.025 //x2=1.01 //y2=6.025
cc_106 ( N_VDD_c_83_p N_A_M4_noxref_g ) capacitor c=0.00678153f //x=3.16 \
 //y=7.4 //x2=1.45 //y2=6.025
cc_107 ( N_VDD_M3_noxref_d N_A_M4_noxref_g ) capacitor c=0.0183011f //x=1.085 \
 //y=5.025 //x2=1.45 //y2=6.025
cc_108 ( N_VDD_c_75_n N_A_c_303_n ) capacitor c=0.00890932f //x=0.74 //y=7.4 \
 //x2=0.955 //y2=4.705
cc_109 ( N_VDD_c_75_n N_B_c_349_n ) capacitor c=7.02327e-19 //x=0.74 //y=7.4 \
 //x2=1.85 //y2=2.08
cc_110 ( N_VDD_c_77_n N_B_c_349_n ) capacitor c=6.16704e-19 //x=3.33 //y=7.4 \
 //x2=1.85 //y2=2.08
cc_111 ( N_VDD_c_83_p N_B_M5_noxref_g ) capacitor c=0.00513565f //x=3.16 \
 //y=7.4 //x2=1.89 //y2=6.025
cc_112 ( N_VDD_c_83_p N_B_M6_noxref_g ) capacitor c=0.00512552f //x=3.16 \
 //y=7.4 //x2=2.33 //y2=6.025
cc_113 ( N_VDD_c_77_n N_B_M6_noxref_g ) capacitor c=0.0120232f //x=3.33 \
 //y=7.4 //x2=2.33 //y2=6.025
cc_114 ( N_VDD_c_78_p N_noxref_6_c_418_n ) capacitor c=0.00568164f //x=5.18 \
 //y=7.4 //x2=1.585 //y2=5.21
cc_115 ( N_VDD_c_106_p N_noxref_6_c_418_n ) capacitor c=4.37585e-19 //x=1.145 \
 //y=7.4 //x2=1.585 //y2=5.21
cc_116 ( N_VDD_c_83_p N_noxref_6_c_418_n ) capacitor c=4.37585e-19 //x=3.16 \
 //y=7.4 //x2=1.585 //y2=5.21
cc_117 ( N_VDD_c_77_n N_noxref_6_c_418_n ) capacitor c=0.00289291f //x=3.33 \
 //y=7.4 //x2=1.585 //y2=5.21
cc_118 ( N_VDD_M3_noxref_d N_noxref_6_c_418_n ) capacitor c=0.0130894f \
 //x=1.085 //y=5.025 //x2=1.585 //y2=5.21
cc_119 ( N_VDD_c_75_n N_noxref_6_c_423_n ) capacitor c=0.0679103f //x=0.74 \
 //y=7.4 //x2=0.875 //y2=5.21
cc_120 ( N_VDD_c_76_n N_noxref_6_c_424_n ) capacitor c=0.00359315f //x=5.18 \
 //y=7.4 //x2=2.465 //y2=6.91
cc_121 ( N_VDD_c_78_p N_noxref_6_c_425_n ) capacitor c=0.0351698f //x=5.18 \
 //y=7.4 //x2=1.755 //y2=6.91
cc_122 ( N_VDD_c_83_p N_noxref_6_c_425_n ) capacitor c=0.0586694f //x=3.16 \
 //y=7.4 //x2=1.755 //y2=6.91
cc_123 ( N_VDD_c_76_n N_noxref_6_c_425_n ) capacitor c=0.00118659f //x=5.18 \
 //y=7.4 //x2=1.755 //y2=6.91
cc_124 ( N_VDD_c_78_p N_noxref_6_M3_noxref_s ) capacitor c=0.00712902f \
 //x=5.18 //y=7.4 //x2=0.655 //y2=5.025
cc_125 ( N_VDD_c_106_p N_noxref_6_M3_noxref_s ) capacitor c=0.0141117f \
 //x=1.145 //y=7.4 //x2=0.655 //y2=5.025
cc_126 ( N_VDD_c_76_n N_noxref_6_M3_noxref_s ) capacitor c=0.00138926f \
 //x=5.18 //y=7.4 //x2=0.655 //y2=5.025
cc_127 ( N_VDD_M3_noxref_d N_noxref_6_M3_noxref_s ) capacitor c=0.0667021f \
 //x=1.085 //y=5.025 //x2=0.655 //y2=5.025
cc_128 ( N_VDD_c_75_n N_noxref_6_M4_noxref_d ) capacitor c=8.88629e-19 \
 //x=0.74 //y=7.4 //x2=1.525 //y2=5.025
cc_129 ( N_VDD_M3_noxref_d N_noxref_6_M4_noxref_d ) capacitor c=0.0659925f \
 //x=1.085 //y=5.025 //x2=1.525 //y2=5.025
cc_130 ( N_VDD_c_77_n N_noxref_6_M6_noxref_d ) capacitor c=0.0520312f //x=3.33 \
 //y=7.4 //x2=2.405 //y2=5.025
cc_131 ( N_VDD_M3_noxref_d N_noxref_6_M6_noxref_d ) capacitor c=0.00107819f \
 //x=1.085 //y=5.025 //x2=2.405 //y2=5.025
cc_132 ( N_VDD_M7_noxref_s N_noxref_6_M6_noxref_d ) capacitor c=0.00226909f \
 //x=3.87 //y=5.02 //x2=2.405 //y2=5.025
cc_133 ( N_VDD_c_76_n Y ) capacitor c=0.0232778f //x=5.18 //y=7.4 //x2=4.81 \
 //y2=2.22
cc_134 ( N_VDD_c_77_n Y ) capacitor c=4.80934e-19 //x=3.33 //y=7.4 //x2=4.81 \
 //y2=2.22
cc_135 ( N_VDD_c_78_p N_Y_c_470_n ) capacitor c=0.00190861f //x=5.18 //y=7.4 \
 //x2=4.725 //y2=4.58
cc_136 ( N_VDD_c_91_p N_Y_c_470_n ) capacitor c=8.8179e-19 //x=4.8 //y=7.4 \
 //x2=4.725 //y2=4.58
cc_137 ( N_VDD_M8_noxref_d N_Y_c_470_n ) capacitor c=0.00641434f //x=4.74 \
 //y=5.02 //x2=4.725 //y2=4.58
cc_138 ( N_VDD_c_77_n N_Y_c_473_n ) capacitor c=0.017572f //x=3.33 //y=7.4 \
 //x2=4.53 //y2=4.58
cc_139 ( N_VDD_c_78_p N_Y_M7_noxref_d ) capacitor c=0.00708604f //x=5.18 \
 //y=7.4 //x2=4.3 //y2=5.02
cc_140 ( N_VDD_c_91_p N_Y_M7_noxref_d ) capacitor c=0.0139004f //x=4.8 //y=7.4 \
 //x2=4.3 //y2=5.02
cc_141 ( N_VDD_c_76_n N_Y_M7_noxref_d ) capacitor c=0.0219131f //x=5.18 \
 //y=7.4 //x2=4.3 //y2=5.02
cc_142 ( N_VDD_M7_noxref_s N_Y_M7_noxref_d ) capacitor c=0.0843065f //x=3.87 \
 //y=5.02 //x2=4.3 //y2=5.02
cc_143 ( N_VDD_M8_noxref_d N_Y_M7_noxref_d ) capacitor c=0.0832641f //x=4.74 \
 //y=5.02 //x2=4.3 //y2=5.02
cc_144 ( N_noxref_3_c_214_p N_A_c_283_n ) capacitor c=0.0112169f //x=1.265 \
 //y=1.655 //x2=1.11 //y2=2.08
cc_145 ( N_noxref_3_c_164_n N_A_c_283_n ) capacitor c=0.00392263f //x=2.59 \
 //y=3.33 //x2=1.11 //y2=2.08
cc_146 ( N_noxref_3_M0_noxref_d N_A_c_286_n ) capacitor c=0.0013184f //x=0.99 \
 //y=0.905 //x2=0.915 //y2=0.905
cc_147 ( N_noxref_3_M0_noxref_d N_A_c_307_n ) capacitor c=0.0034598f //x=0.99 \
 //y=0.905 //x2=0.915 //y2=1.25
cc_148 ( N_noxref_3_M0_noxref_d N_A_c_308_n ) capacitor c=0.00300148f //x=0.99 \
 //y=0.905 //x2=0.915 //y2=1.56
cc_149 ( N_noxref_3_c_214_p N_A_c_288_n ) capacitor c=0.00589082f //x=1.265 \
 //y=1.655 //x2=0.915 //y2=1.915
cc_150 ( N_noxref_3_M0_noxref_d N_A_c_288_n ) capacitor c=0.00273686f //x=0.99 \
 //y=0.905 //x2=0.915 //y2=1.915
cc_151 ( N_noxref_3_M0_noxref_d N_A_c_290_n ) capacitor c=0.00241102f //x=0.99 \
 //y=0.905 //x2=1.29 //y2=0.75
cc_152 ( N_noxref_3_M0_noxref_d N_A_c_312_n ) capacitor c=0.0123304f //x=0.99 \
 //y=0.905 //x2=1.29 //y2=1.405
cc_153 ( N_noxref_3_M0_noxref_d N_A_c_291_n ) capacitor c=0.00219619f //x=0.99 \
 //y=0.905 //x2=1.445 //y2=0.905
cc_154 ( N_noxref_3_c_155_n N_A_c_293_n ) capacitor c=0.00431513f //x=2.065 \
 //y=1.655 //x2=1.445 //y2=1.25
cc_155 ( N_noxref_3_M0_noxref_d N_A_c_293_n ) capacitor c=0.00603828f //x=0.99 \
 //y=0.905 //x2=1.445 //y2=1.25
cc_156 ( N_noxref_3_c_164_n N_B_c_362_n ) capacitor c=0.0102183f //x=2.59 \
 //y=3.33 //x2=1.85 //y2=4.54
cc_157 ( N_noxref_3_c_153_n N_B_c_349_n ) capacitor c=0.00717888f //x=2.705 \
 //y=3.33 //x2=1.85 //y2=2.08
cc_158 ( N_noxref_3_c_155_n N_B_c_349_n ) capacitor c=0.0162392f //x=2.065 \
 //y=1.655 //x2=1.85 //y2=2.08
cc_159 ( N_noxref_3_c_164_n N_B_c_349_n ) capacitor c=0.0815617f //x=2.59 \
 //y=3.33 //x2=1.85 //y2=2.08
cc_160 ( N_noxref_3_c_165_n N_B_c_349_n ) capacitor c=0.00126776f //x=4.07 \
 //y=2.085 //x2=1.85 //y2=2.08
cc_161 ( N_noxref_3_c_196_n N_B_M5_noxref_g ) capacitor c=0.0132788f //x=2.195 \
 //y=5.21 //x2=1.89 //y2=6.025
cc_162 ( N_noxref_3_c_194_n N_B_M6_noxref_g ) capacitor c=0.0217686f //x=2.505 \
 //y=5.21 //x2=2.33 //y2=6.025
cc_163 ( N_noxref_3_M5_noxref_d N_B_M6_noxref_g ) capacitor c=0.0136385f \
 //x=1.965 //y=5.025 //x2=2.33 //y2=6.025
cc_164 ( N_noxref_3_M1_noxref_d N_B_c_351_n ) capacitor c=0.00226395f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=0.905
cc_165 ( N_noxref_3_M1_noxref_d N_B_c_371_n ) capacitor c=0.0035101f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.255
cc_166 ( N_noxref_3_c_155_n N_B_c_372_n ) capacitor c=0.00218915f //x=2.065 \
 //y=1.655 //x2=1.885 //y2=1.56
cc_167 ( N_noxref_3_M0_noxref_d N_B_c_372_n ) capacitor c=0.00148728f //x=0.99 \
 //y=0.905 //x2=1.885 //y2=1.56
cc_168 ( N_noxref_3_M1_noxref_d N_B_c_372_n ) capacitor c=0.00546704f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.56
cc_169 ( N_noxref_3_c_196_n N_B_c_375_n ) capacitor c=0.00410596f //x=2.195 \
 //y=5.21 //x2=2.255 //y2=4.795
cc_170 ( N_noxref_3_c_164_n N_B_c_375_n ) capacitor c=0.0144455f //x=2.59 \
 //y=3.33 //x2=2.255 //y2=4.795
cc_171 ( N_noxref_3_M1_noxref_d N_B_c_353_n ) capacitor c=0.00241102f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=0.75
cc_172 ( N_noxref_3_c_159_n N_B_c_354_n ) capacitor c=0.00801563f //x=2.505 \
 //y=1.655 //x2=2.26 //y2=1.405
cc_173 ( N_noxref_3_M1_noxref_d N_B_c_354_n ) capacitor c=0.0158021f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=1.405
cc_174 ( N_noxref_3_M1_noxref_d N_B_c_355_n ) capacitor c=0.00132831f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=0.905
cc_175 ( N_noxref_3_M1_noxref_d N_B_c_381_n ) capacitor c=0.0035101f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=1.255
cc_176 ( N_noxref_3_c_155_n N_B_c_382_n ) capacitor c=0.00633758f //x=2.065 \
 //y=1.655 //x2=1.85 //y2=2.08
cc_177 ( N_noxref_3_c_164_n N_B_c_382_n ) capacitor c=0.00877984f //x=2.59 \
 //y=3.33 //x2=1.85 //y2=2.08
cc_178 ( N_noxref_3_c_155_n N_B_c_384_n ) capacitor c=0.0189958f //x=2.065 \
 //y=1.655 //x2=1.85 //y2=1.915
cc_179 ( N_noxref_3_c_164_n N_B_c_384_n ) capacitor c=0.00306024f //x=2.59 \
 //y=3.33 //x2=1.85 //y2=1.915
cc_180 ( N_noxref_3_M1_noxref_d N_B_c_384_n ) capacitor c=3.4952e-19 //x=1.96 \
 //y=0.905 //x2=1.85 //y2=1.915
cc_181 ( N_noxref_3_c_164_n N_B_c_387_n ) capacitor c=0.00537091f //x=2.59 \
 //y=3.33 //x2=1.885 //y2=4.705
cc_182 ( N_noxref_3_c_196_n N_noxref_6_c_418_n ) capacitor c=0.0348754f \
 //x=2.195 //y=5.21 //x2=1.585 //y2=5.21
cc_183 ( N_noxref_3_c_194_n N_noxref_6_c_424_n ) capacitor c=0.00173777f \
 //x=2.505 //y=5.21 //x2=2.465 //y2=6.91
cc_184 ( N_noxref_3_M5_noxref_d N_noxref_6_c_424_n ) capacitor c=0.0118172f \
 //x=1.965 //y=5.025 //x2=2.465 //y2=6.91
cc_185 ( N_noxref_3_M5_noxref_d N_noxref_6_M3_noxref_s ) capacitor \
 c=0.00107541f //x=1.965 //y=5.025 //x2=0.655 //y2=5.025
cc_186 ( N_noxref_3_M5_noxref_d N_noxref_6_M4_noxref_d ) capacitor \
 c=0.0348754f //x=1.965 //y=5.025 //x2=1.525 //y2=5.025
cc_187 ( N_noxref_3_c_194_n N_noxref_6_M6_noxref_d ) capacitor c=0.015774f \
 //x=2.505 //y=5.21 //x2=2.405 //y2=5.025
cc_188 ( N_noxref_3_M5_noxref_d N_noxref_6_M6_noxref_d ) capacitor \
 c=0.0458293f //x=1.965 //y=5.025 //x2=2.405 //y2=5.025
cc_189 ( N_noxref_3_c_147_n Y ) capacitor c=0.00582634f //x=3.955 //y=3.33 \
 //x2=4.81 //y2=2.22
cc_190 ( N_noxref_3_c_164_n Y ) capacitor c=0.00126776f //x=2.59 //y=3.33 \
 //x2=4.81 //y2=2.22
cc_191 ( N_noxref_3_c_165_n Y ) capacitor c=0.0711303f //x=4.07 //y=2.085 \
 //x2=4.81 //y2=2.22
cc_192 ( N_noxref_3_c_177_n Y ) capacitor c=8.49451e-19 //x=4.07 //y=2.085 \
 //x2=4.81 //y2=2.22
cc_193 ( N_noxref_3_c_263_p N_Y_c_460_n ) capacitor c=0.0023507f //x=4.555 \
 //y=1.41 //x2=4.725 //y2=2.08
cc_194 ( N_noxref_3_c_177_n N_Y_c_484_n ) capacitor c=0.0167852f //x=4.07 \
 //y=2.085 //x2=4.525 //y2=2.08
cc_195 ( N_noxref_3_c_208_n N_Y_c_470_n ) capacitor c=0.0101013f //x=4.59 \
 //y=4.79 //x2=4.725 //y2=4.58
cc_196 ( N_noxref_3_c_165_n N_Y_c_473_n ) capacitor c=0.0250878f //x=4.07 \
 //y=2.085 //x2=4.53 //y2=4.58
cc_197 ( N_noxref_3_c_209_n N_Y_c_473_n ) capacitor c=0.00962086f //x=4.3 \
 //y=4.79 //x2=4.53 //y2=4.58
cc_198 ( N_noxref_3_c_164_n N_Y_M2_noxref_d ) capacitor c=3.35192e-19 //x=2.59 \
 //y=3.33 //x2=4.255 //y2=0.91
cc_199 ( N_noxref_3_c_165_n N_Y_M2_noxref_d ) capacitor c=0.0175773f //x=4.07 \
 //y=2.085 //x2=4.255 //y2=0.91
cc_200 ( N_noxref_3_c_170_n N_Y_M2_noxref_d ) capacitor c=0.00218556f //x=4.18 \
 //y=0.91 //x2=4.255 //y2=0.91
cc_201 ( N_noxref_3_c_271_p N_Y_M2_noxref_d ) capacitor c=0.00347355f //x=4.18 \
 //y=1.255 //x2=4.255 //y2=0.91
cc_202 ( N_noxref_3_c_272_p N_Y_M2_noxref_d ) capacitor c=0.00742431f //x=4.18 \
 //y=1.565 //x2=4.255 //y2=0.91
cc_203 ( N_noxref_3_c_172_n N_Y_M2_noxref_d ) capacitor c=0.00957707f //x=4.18 \
 //y=1.92 //x2=4.255 //y2=0.91
cc_204 ( N_noxref_3_c_173_n N_Y_M2_noxref_d ) capacitor c=0.00220879f \
 //x=4.555 //y=0.755 //x2=4.255 //y2=0.91
cc_205 ( N_noxref_3_c_263_p N_Y_M2_noxref_d ) capacitor c=0.0138447f //x=4.555 \
 //y=1.41 //x2=4.255 //y2=0.91
cc_206 ( N_noxref_3_c_174_n N_Y_M2_noxref_d ) capacitor c=0.00218624f //x=4.71 \
 //y=0.91 //x2=4.255 //y2=0.91
cc_207 ( N_noxref_3_c_176_n N_Y_M2_noxref_d ) capacitor c=0.00601286f //x=4.71 \
 //y=1.255 //x2=4.255 //y2=0.91
cc_208 ( N_noxref_3_c_164_n N_Y_M7_noxref_d ) capacitor c=6.2839e-19 //x=2.59 \
 //y=3.33 //x2=4.3 //y2=5.02
cc_209 ( N_noxref_3_M7_noxref_g N_Y_M7_noxref_d ) capacitor c=0.0219309f \
 //x=4.225 //y=6.02 //x2=4.3 //y2=5.02
cc_210 ( N_noxref_3_M8_noxref_g N_Y_M7_noxref_d ) capacitor c=0.021902f \
 //x=4.665 //y=6.02 //x2=4.3 //y2=5.02
cc_211 ( N_noxref_3_c_208_n N_Y_M7_noxref_d ) capacitor c=0.0148755f //x=4.59 \
 //y=4.79 //x2=4.3 //y2=5.02
cc_212 ( N_noxref_3_c_209_n N_Y_M7_noxref_d ) capacitor c=0.00307344f //x=4.3 \
 //y=4.79 //x2=4.3 //y2=5.02
cc_213 ( N_A_c_295_n N_B_c_362_n ) capacitor c=0.0480335f //x=0.955 //y=4.705 \
 //x2=1.85 //y2=4.54
cc_214 ( N_A_c_317_p N_B_c_362_n ) capacitor c=0.00146509f //x=1.375 //y=4.795 \
 //x2=1.85 //y2=4.54
cc_215 ( N_A_c_303_n N_B_c_362_n ) capacitor c=0.00112871f //x=0.955 //y=4.705 \
 //x2=1.85 //y2=4.54
cc_216 ( N_A_c_283_n N_B_c_349_n ) capacitor c=0.0452884f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_217 ( N_A_c_288_n N_B_c_349_n ) capacitor c=0.00308814f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_218 ( N_A_M3_noxref_g N_B_M5_noxref_g ) capacitor c=0.0100243f //x=1.01 \
 //y=6.025 //x2=1.89 //y2=6.025
cc_219 ( N_A_M4_noxref_g N_B_M5_noxref_g ) capacitor c=0.107798f //x=1.45 \
 //y=6.025 //x2=1.89 //y2=6.025
cc_220 ( N_A_M4_noxref_g N_B_M6_noxref_g ) capacitor c=0.0094155f //x=1.45 \
 //y=6.025 //x2=2.33 //y2=6.025
cc_221 ( N_A_c_286_n N_B_c_351_n ) capacitor c=0.00125788f //x=0.915 //y=0.905 \
 //x2=1.885 //y2=0.905
cc_222 ( N_A_c_291_n N_B_c_351_n ) capacitor c=0.0126654f //x=1.445 //y=0.905 \
 //x2=1.885 //y2=0.905
cc_223 ( N_A_c_307_n N_B_c_371_n ) capacitor c=0.00148539f //x=0.915 //y=1.25 \
 //x2=1.885 //y2=1.255
cc_224 ( N_A_c_308_n N_B_c_371_n ) capacitor c=0.00105591f //x=0.915 //y=1.56 \
 //x2=1.885 //y2=1.255
cc_225 ( N_A_c_293_n N_B_c_371_n ) capacitor c=0.0126654f //x=1.445 //y=1.25 \
 //x2=1.885 //y2=1.255
cc_226 ( N_A_c_308_n N_B_c_372_n ) capacitor c=0.00109549f //x=0.915 //y=1.56 \
 //x2=1.885 //y2=1.56
cc_227 ( N_A_c_293_n N_B_c_372_n ) capacitor c=0.00886999f //x=1.445 //y=1.25 \
 //x2=1.885 //y2=1.56
cc_228 ( N_A_c_293_n N_B_c_354_n ) capacitor c=0.00123863f //x=1.445 //y=1.25 \
 //x2=2.26 //y2=1.405
cc_229 ( N_A_c_291_n N_B_c_355_n ) capacitor c=0.00132934f //x=1.445 //y=0.905 \
 //x2=2.415 //y2=0.905
cc_230 ( N_A_c_293_n N_B_c_381_n ) capacitor c=0.00150734f //x=1.445 //y=1.25 \
 //x2=2.415 //y2=1.255
cc_231 ( N_A_c_283_n N_B_c_382_n ) capacitor c=0.00307062f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_232 ( N_A_c_288_n N_B_c_382_n ) capacitor c=0.0179092f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_233 ( N_A_c_288_n N_B_c_384_n ) capacitor c=0.00577193f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=1.915
cc_234 ( N_A_c_295_n N_B_c_387_n ) capacitor c=0.00336963f //x=0.955 //y=4.705 \
 //x2=1.885 //y2=4.705
cc_235 ( N_A_c_317_p N_B_c_387_n ) capacitor c=0.020271f //x=1.375 //y=4.795 \
 //x2=1.885 //y2=4.705
cc_236 ( N_A_c_303_n N_B_c_387_n ) capacitor c=0.00546725f //x=0.955 //y=4.705 \
 //x2=1.885 //y2=4.705
cc_237 ( N_A_c_295_n N_noxref_6_c_418_n ) capacitor c=0.00628365f //x=0.955 \
 //y=4.705 //x2=1.585 //y2=5.21
cc_238 ( N_A_M3_noxref_g N_noxref_6_c_418_n ) capacitor c=0.0182391f //x=1.01 \
 //y=6.025 //x2=1.585 //y2=5.21
cc_239 ( N_A_M4_noxref_g N_noxref_6_c_418_n ) capacitor c=0.0203804f //x=1.45 \
 //y=6.025 //x2=1.585 //y2=5.21
cc_240 ( N_A_c_317_p N_noxref_6_c_418_n ) capacitor c=0.00343485f //x=1.375 \
 //y=4.795 //x2=1.585 //y2=5.21
cc_241 ( N_A_c_303_n N_noxref_6_c_418_n ) capacitor c=0.0017421f //x=0.955 \
 //y=4.705 //x2=1.585 //y2=5.21
cc_242 ( N_A_c_295_n N_noxref_6_c_423_n ) capacitor c=0.0120346f //x=0.955 \
 //y=4.705 //x2=0.875 //y2=5.21
cc_243 ( N_A_c_303_n N_noxref_6_c_423_n ) capacitor c=0.00518332f //x=0.955 \
 //y=4.705 //x2=0.875 //y2=5.21
cc_244 ( N_A_M3_noxref_g N_noxref_6_M3_noxref_s ) capacitor c=0.0473218f \
 //x=1.01 //y=6.025 //x2=0.655 //y2=5.025
cc_245 ( N_A_M4_noxref_g N_noxref_6_M4_noxref_d ) capacitor c=0.0170604f \
 //x=1.45 //y=6.025 //x2=1.525 //y2=5.025
cc_246 ( N_B_M5_noxref_g N_noxref_6_c_418_n ) capacitor c=0.0170604f //x=1.89 \
 //y=6.025 //x2=1.585 //y2=5.21
cc_247 ( N_B_c_387_n N_noxref_6_c_418_n ) capacitor c=2.24869e-19 //x=1.885 \
 //y=4.705 //x2=1.585 //y2=5.21
cc_248 ( N_B_c_362_n N_noxref_6_c_424_n ) capacitor c=8.92402e-19 //x=1.85 \
 //y=4.54 //x2=2.465 //y2=6.91
cc_249 ( N_B_M5_noxref_g N_noxref_6_c_424_n ) capacitor c=0.0148484f //x=1.89 \
 //y=6.025 //x2=2.465 //y2=6.91
cc_250 ( N_B_M6_noxref_g N_noxref_6_c_424_n ) capacitor c=0.0163196f //x=2.33 \
 //y=6.025 //x2=2.465 //y2=6.91
cc_251 ( N_B_M6_noxref_g N_noxref_6_M6_noxref_d ) capacitor c=0.0351101f \
 //x=2.33 //y=6.025 //x2=2.405 //y2=5.025
