magic
tech sky130A
magscale 1 2
timestamp 1670281657
<< nwell >>
rect -87 786 309 1550
<< pwell >>
rect -34 -34 256 544
<< psubdiff >>
rect -34 482 256 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 17 34 57
rect 188 461 256 482
rect 188 427 205 461
rect 239 427 256 461
rect 188 387 256 427
rect 188 353 205 387
rect 239 353 256 387
rect 188 313 256 353
rect 188 279 205 313
rect 239 279 256 313
rect 188 239 256 279
rect 188 205 205 239
rect 239 205 256 239
rect 188 165 256 205
rect 188 131 205 165
rect 239 131 256 165
rect 188 91 256 131
rect 188 57 205 91
rect 239 57 256 91
rect 188 17 256 57
rect -34 -17 94 17
rect 128 -17 256 17
rect -34 -34 256 -17
<< nsubdiff >>
rect -34 1497 256 1514
rect -34 1463 94 1497
rect 128 1463 256 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 884 34 905
rect 188 1423 256 1463
rect 188 1389 205 1423
rect 239 1389 256 1423
rect 188 1349 256 1389
rect 188 1315 205 1349
rect 239 1315 256 1349
rect 188 1275 256 1315
rect 188 1241 205 1275
rect 239 1241 256 1275
rect 188 1201 256 1241
rect 188 1167 205 1201
rect 239 1167 256 1201
rect 188 1127 256 1167
rect 188 1093 205 1127
rect 239 1093 256 1127
rect 188 1053 256 1093
rect 188 1019 205 1053
rect 239 1019 256 1053
rect 188 979 256 1019
rect 188 945 205 979
rect 239 945 256 979
rect 188 905 256 945
rect 188 884 205 905
rect 17 871 205 884
rect 239 871 256 905
rect -34 822 256 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 205 427 239 461
rect 205 353 239 387
rect 205 279 239 313
rect 205 205 239 239
rect 205 131 239 165
rect 205 57 239 91
rect 94 -17 128 17
<< nsubdiffcont >>
rect 94 1463 128 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect -17 945 17 979
rect -17 871 17 905
rect 205 1389 239 1423
rect 205 1315 239 1349
rect 205 1241 239 1275
rect 205 1167 239 1201
rect 205 1093 239 1127
rect 205 1019 239 1053
rect 205 945 239 979
rect 205 871 239 905
<< locali >>
rect -34 1497 256 1514
rect -34 1463 94 1497
rect 128 1463 256 1497
rect -34 1446 256 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 188 1423 256 1446
rect 188 1389 205 1423
rect 239 1389 256 1423
rect 188 1349 256 1389
rect 188 1315 205 1349
rect 239 1315 256 1349
rect 188 1275 256 1315
rect 188 1241 205 1275
rect 239 1241 256 1275
rect 188 1201 256 1241
rect 188 1167 205 1201
rect 239 1167 256 1201
rect 188 1127 256 1167
rect 188 1093 205 1127
rect 239 1093 256 1127
rect 188 1053 256 1093
rect 188 1019 205 1053
rect 239 1019 256 1053
rect 188 979 256 1019
rect 188 945 205 979
rect 239 945 256 979
rect 188 905 256 945
rect 188 871 205 905
rect 239 871 256 905
rect 188 822 256 871
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 188 461 256 544
rect 188 427 205 461
rect 239 427 256 461
rect 188 387 256 427
rect 188 353 205 387
rect 239 353 256 387
rect 188 313 256 353
rect 188 279 205 313
rect 239 279 256 313
rect 188 239 256 279
rect 188 205 205 239
rect 239 205 256 239
rect 188 165 256 205
rect 188 131 205 165
rect 239 131 256 165
rect 188 91 256 131
rect 188 57 205 91
rect 239 57 256 91
rect 188 34 256 57
rect -34 17 256 34
rect -34 -17 94 17
rect 128 -17 256 17
rect -34 -34 256 -17
<< metal1 >>
rect -34 1446 256 1514
rect -34 -34 256 34
<< labels >>
rlabel metal1 -34 1446 256 1514 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 -34 -34 256 34 1 GND
port 2 nsew ground bidirectional abutment
<< end >>
