// File: MUX2X1.spi.MUX2X1.pxi
// Created: Tue Oct 15 15:49:38 2024
// 
simulator lang=spectre
x_PM_MUX2X1\%GND ( GND N_GND_c_6_p N_GND_c_7_p N_GND_c_24_p N_GND_c_114_p \
 N_GND_c_8_p N_GND_c_9_p N_GND_c_33_p N_GND_c_46_p N_GND_c_53_p N_GND_c_66_p \
 N_GND_c_5_p N_GND_c_1_p N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p N_GND_M0_noxref_s \
 N_GND_M1_noxref_d N_GND_M3_noxref_d N_GND_M5_noxref_d )  PM_MUX2X1\%GND
x_PM_MUX2X1\%VDD ( VDD N_VDD_c_171_p N_VDD_c_181_p N_VDD_c_179_p N_VDD_c_226_p \
 N_VDD_c_210_p N_VDD_c_264_p N_VDD_c_237_p N_VDD_c_276_p N_VDD_c_166_n \
 N_VDD_c_167_n N_VDD_c_168_n N_VDD_c_169_n N_VDD_c_170_n N_VDD_M7_noxref_s \
 N_VDD_M8_noxref_d N_VDD_M9_noxref_s N_VDD_M10_noxref_d N_VDD_M12_noxref_d \
 N_VDD_M13_noxref_s N_VDD_M14_noxref_d N_VDD_M16_noxref_d N_VDD_M17_noxref_s \
 N_VDD_M18_noxref_d N_VDD_M20_noxref_d )  PM_MUX2X1\%VDD
x_PM_MUX2X1\%S ( N_S_c_329_n N_S_c_335_n S S S S S S S S S S S S S N_S_c_337_n \
 N_S_c_342_n N_S_M0_noxref_g N_S_M1_noxref_g N_S_M7_noxref_g N_S_M8_noxref_g \
 N_S_M9_noxref_g N_S_M10_noxref_g N_S_c_343_n N_S_c_404_p N_S_c_405_p \
 N_S_c_345_n N_S_c_381_n N_S_c_382_n N_S_c_346_n N_S_c_391_p N_S_c_347_n \
 N_S_c_349_n N_S_c_350_n N_S_c_352_n N_S_c_433_p N_S_c_353_n N_S_c_354_n \
 N_S_c_355_n N_S_c_356_n N_S_c_358_n N_S_c_359_n N_S_c_384_n )  PM_MUX2X1\%S
x_PM_MUX2X1\%noxref_4 ( N_noxref_4_c_456_n N_noxref_4_c_486_n \
 N_noxref_4_c_458_n N_noxref_4_c_515_n N_noxref_4_c_488_n N_noxref_4_c_491_n \
 N_noxref_4_c_461_n N_noxref_4_c_462_n N_noxref_4_M3_noxref_g \
 N_noxref_4_M13_noxref_g N_noxref_4_M14_noxref_g N_noxref_4_c_463_n \
 N_noxref_4_c_465_n N_noxref_4_c_466_n N_noxref_4_c_467_n N_noxref_4_c_468_n \
 N_noxref_4_c_469_n N_noxref_4_c_470_n N_noxref_4_c_472_n N_noxref_4_c_501_n \
 N_noxref_4_M0_noxref_d N_noxref_4_M7_noxref_d )  PM_MUX2X1\%noxref_4
x_PM_MUX2X1\%noxref_5 ( N_noxref_5_c_595_n N_noxref_5_c_602_n \
 N_noxref_5_c_620_n N_noxref_5_c_624_n N_noxref_5_c_626_n N_noxref_5_c_603_n \
 N_noxref_5_c_667_n N_noxref_5_c_604_n N_noxref_5_c_605_n N_noxref_5_c_714_p \
 N_noxref_5_M5_noxref_g N_noxref_5_M17_noxref_g N_noxref_5_M18_noxref_g \
 N_noxref_5_c_606_n N_noxref_5_c_608_n N_noxref_5_c_609_n N_noxref_5_c_610_n \
 N_noxref_5_c_611_n N_noxref_5_c_612_n N_noxref_5_c_613_n N_noxref_5_c_615_n \
 N_noxref_5_c_639_n N_noxref_5_M2_noxref_d N_noxref_5_M9_noxref_d \
 N_noxref_5_M11_noxref_d )  PM_MUX2X1\%noxref_5
x_PM_MUX2X1\%noxref_6 ( N_noxref_6_c_763_n N_noxref_6_c_774_n \
 N_noxref_6_c_776_n N_noxref_6_c_780_n N_noxref_6_c_782_n N_noxref_6_c_764_n \
 N_noxref_6_c_822_n N_noxref_6_c_765_n N_noxref_6_c_826_n N_noxref_6_c_766_n \
 N_noxref_6_c_860_p N_noxref_6_M6_noxref_g N_noxref_6_M19_noxref_g \
 N_noxref_6_M20_noxref_g N_noxref_6_c_834_n N_noxref_6_c_837_n \
 N_noxref_6_c_839_n N_noxref_6_c_882_p N_noxref_6_c_898_p N_noxref_6_c_892_p \
 N_noxref_6_c_842_n N_noxref_6_c_843_n N_noxref_6_c_844_n N_noxref_6_c_884_p \
 N_noxref_6_c_846_n N_noxref_6_M4_noxref_d N_noxref_6_M13_noxref_d \
 N_noxref_6_M15_noxref_d )  PM_MUX2X1\%noxref_6
x_PM_MUX2X1\%A0 ( A0 A0 A0 A0 A0 A0 N_A0_c_927_n N_A0_c_918_n N_A0_M2_noxref_g \
 N_A0_M11_noxref_g N_A0_M12_noxref_g N_A0_c_935_n N_A0_c_938_n N_A0_c_940_n \
 N_A0_c_964_n N_A0_c_966_n N_A0_c_967_n N_A0_c_943_n N_A0_c_944_n N_A0_c_945_n \
 N_A0_c_973_n N_A0_c_947_n )  PM_MUX2X1\%A0
x_PM_MUX2X1\%noxref_8 ( N_noxref_8_c_986_n N_noxref_8_c_987_n \
 N_noxref_8_c_991_n N_noxref_8_c_995_n N_noxref_8_c_996_n N_noxref_8_c_999_n \
 N_noxref_8_M1_noxref_s )  PM_MUX2X1\%noxref_8
x_PM_MUX2X1\%A1 ( A1 A1 A1 A1 A1 A1 N_A1_c_1052_n N_A1_c_1043_n \
 N_A1_M4_noxref_g N_A1_M15_noxref_g N_A1_M16_noxref_g N_A1_c_1060_n \
 N_A1_c_1063_n N_A1_c_1065_n N_A1_c_1090_n N_A1_c_1092_n N_A1_c_1093_n \
 N_A1_c_1068_n N_A1_c_1069_n N_A1_c_1070_n N_A1_c_1099_n N_A1_c_1072_n )  \
 PM_MUX2X1\%A1
x_PM_MUX2X1\%noxref_10 ( N_noxref_10_c_1134_n N_noxref_10_c_1112_n \
 N_noxref_10_c_1116_n N_noxref_10_c_1120_n N_noxref_10_c_1121_n \
 N_noxref_10_c_1124_n N_noxref_10_M3_noxref_s )  PM_MUX2X1\%noxref_10
x_PM_MUX2X1\%Y ( Y Y Y Y Y Y Y Y N_Y_c_1174_n N_Y_c_1178_n N_Y_c_1180_n \
 N_Y_c_1168_n N_Y_c_1226_p N_Y_c_1215_n N_Y_M6_noxref_d N_Y_M17_noxref_d \
 N_Y_M19_noxref_d )  PM_MUX2X1\%Y
x_PM_MUX2X1\%noxref_12 ( N_noxref_12_c_1249_n N_noxref_12_c_1232_n \
 N_noxref_12_c_1236_n N_noxref_12_c_1239_n N_noxref_12_c_1240_n \
 N_noxref_12_c_1242_n N_noxref_12_M5_noxref_s )  PM_MUX2X1\%noxref_12
cc_1 ( N_GND_c_1_p N_VDD_c_166_n ) capacitor c=0.00989031f //x=0.63 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_167_n ) capacitor c=0.00829849f //x=2.22 //y=0 \
 //x2=2.22 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_168_n ) capacitor c=0.00829849f //x=5.55 //y=0 \
 //x2=5.55 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_169_n ) capacitor c=0.00829849f //x=8.88 //y=0 \
 //x2=8.88 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_170_n ) capacitor c=0.00989031f //x=11.47 //y=0 \
 //x2=11.47 //y2=7.4
cc_6 ( N_GND_c_6_p N_S_c_329_n ) capacitor c=0.0211888f //x=11.47 //y=0 \
 //x2=3.215 //y2=2.96
cc_7 ( N_GND_c_7_p N_S_c_329_n ) capacitor c=0.00114872f //x=1.03 //y=0.535 \
 //x2=3.215 //y2=2.96
cc_8 ( N_GND_c_8_p N_S_c_329_n ) capacitor c=0.00129597f //x=2.05 //y=0 \
 //x2=3.215 //y2=2.96
cc_9 ( N_GND_c_9_p N_S_c_329_n ) capacitor c=0.00230184f //x=3.315 //y=0 \
 //x2=3.215 //y2=2.96
cc_10 ( N_GND_c_2_p N_S_c_329_n ) capacitor c=0.0144849f //x=2.22 //y=0 \
 //x2=3.215 //y2=2.96
cc_11 ( N_GND_M0_noxref_s N_S_c_329_n ) capacitor c=0.00258314f //x=0.495 \
 //y=0.37 //x2=3.215 //y2=2.96
cc_12 ( N_GND_c_6_p N_S_c_335_n ) capacitor c=0.00206599f //x=11.47 //y=0 \
 //x2=0.855 //y2=2.96
cc_13 ( N_GND_M0_noxref_s N_S_c_335_n ) capacitor c=0.00142333f //x=0.495 \
 //y=0.37 //x2=0.855 //y2=2.96
cc_14 ( N_GND_c_6_p N_S_c_337_n ) capacitor c=0.00183756f //x=11.47 //y=0 \
 //x2=0.74 //y2=2.085
cc_15 ( N_GND_c_7_p N_S_c_337_n ) capacitor c=7.8474e-19 //x=1.03 //y=0.535 \
 //x2=0.74 //y2=2.085
cc_16 ( N_GND_c_1_p N_S_c_337_n ) capacitor c=0.0293771f //x=0.63 //y=0 \
 //x2=0.74 //y2=2.085
cc_17 ( N_GND_c_2_p N_S_c_337_n ) capacitor c=0.00118911f //x=2.22 //y=0 \
 //x2=0.74 //y2=2.085
cc_18 ( N_GND_M0_noxref_s N_S_c_337_n ) capacitor c=0.0102424f //x=0.495 \
 //y=0.37 //x2=0.74 //y2=2.085
cc_19 ( N_GND_c_2_p N_S_c_342_n ) capacitor c=0.0179404f //x=2.22 //y=0 \
 //x2=3.33 //y2=2.08
cc_20 ( N_GND_c_7_p N_S_c_343_n ) capacitor c=0.0123171f //x=1.03 //y=0.535 \
 //x2=0.85 //y2=0.91
cc_21 ( N_GND_M0_noxref_s N_S_c_343_n ) capacitor c=0.0316657f //x=0.495 \
 //y=0.37 //x2=0.85 //y2=0.91
cc_22 ( N_GND_c_1_p N_S_c_345_n ) capacitor c=0.0124051f //x=0.63 //y=0 \
 //x2=0.85 //y2=1.92
cc_23 ( N_GND_M0_noxref_s N_S_c_346_n ) capacitor c=0.00489f //x=0.495 \
 //y=0.37 //x2=1.225 //y2=0.755
cc_24 ( N_GND_c_24_p N_S_c_347_n ) capacitor c=0.0119174f //x=1.515 //y=0.535 \
 //x2=1.38 //y2=0.91
cc_25 ( N_GND_M0_noxref_s N_S_c_347_n ) capacitor c=0.0143355f //x=0.495 \
 //y=0.37 //x2=1.38 //y2=0.91
cc_26 ( N_GND_M0_noxref_s N_S_c_349_n ) capacitor c=0.0074042f //x=0.495 \
 //y=0.37 //x2=1.38 //y2=1.255
cc_27 ( N_GND_c_9_p N_S_c_350_n ) capacitor c=0.00135046f //x=3.315 //y=0 \
 //x2=3.135 //y2=0.865
cc_28 ( N_GND_M1_noxref_d N_S_c_350_n ) capacitor c=0.00220047f //x=3.21 \
 //y=0.865 //x2=3.135 //y2=0.865
cc_29 ( N_GND_M1_noxref_d N_S_c_352_n ) capacitor c=0.00255985f //x=3.21 \
 //y=0.865 //x2=3.135 //y2=1.21
cc_30 ( N_GND_c_2_p N_S_c_353_n ) capacitor c=0.0114883f //x=2.22 //y=0 \
 //x2=3.135 //y2=1.915
cc_31 ( N_GND_M1_noxref_d N_S_c_354_n ) capacitor c=0.0131326f //x=3.21 \
 //y=0.865 //x2=3.51 //y2=0.71
cc_32 ( N_GND_M1_noxref_d N_S_c_355_n ) capacitor c=0.00193127f //x=3.21 \
 //y=0.865 //x2=3.51 //y2=1.365
cc_33 ( N_GND_c_33_p N_S_c_356_n ) capacitor c=0.00130622f //x=5.38 //y=0 \
 //x2=3.665 //y2=0.865
cc_34 ( N_GND_M1_noxref_d N_S_c_356_n ) capacitor c=0.00257848f //x=3.21 \
 //y=0.865 //x2=3.665 //y2=0.865
cc_35 ( N_GND_M1_noxref_d N_S_c_358_n ) capacitor c=0.00255985f //x=3.21 \
 //y=0.865 //x2=3.665 //y2=1.21
cc_36 ( N_GND_c_7_p N_S_c_359_n ) capacitor c=2.1838e-19 //x=1.03 //y=0.535 \
 //x2=0.74 //y2=2.085
cc_37 ( N_GND_c_1_p N_S_c_359_n ) capacitor c=0.0108179f //x=0.63 //y=0 \
 //x2=0.74 //y2=2.085
cc_38 ( N_GND_M0_noxref_s N_S_c_359_n ) capacitor c=0.00652836f //x=0.495 \
 //y=0.37 //x2=0.74 //y2=2.085
cc_39 ( N_GND_c_6_p N_noxref_4_c_456_n ) capacitor c=0.0249003f //x=11.47 \
 //y=0 //x2=6.545 //y2=3.33
cc_40 ( N_GND_c_33_p N_noxref_4_c_456_n ) capacitor c=5.39691e-19 //x=5.38 \
 //y=0 //x2=6.545 //y2=3.33
cc_41 ( N_GND_c_6_p N_noxref_4_c_458_n ) capacitor c=0.00130393f //x=11.47 \
 //y=0 //x2=1.395 //y2=2.08
cc_42 ( N_GND_c_2_p N_noxref_4_c_458_n ) capacitor c=0.0296841f //x=2.22 //y=0 \
 //x2=1.395 //y2=2.08
cc_43 ( N_GND_M0_noxref_s N_noxref_4_c_458_n ) capacitor c=0.00967469f \
 //x=0.495 //y=0.37 //x2=1.395 //y2=2.08
cc_44 ( N_GND_c_1_p N_noxref_4_c_461_n ) capacitor c=8.10282e-19 //x=0.63 \
 //y=0 //x2=1.48 //y2=3.33
cc_45 ( N_GND_c_3_p N_noxref_4_c_462_n ) capacitor c=0.0179404f //x=5.55 //y=0 \
 //x2=6.66 //y2=2.08
cc_46 ( N_GND_c_46_p N_noxref_4_c_463_n ) capacitor c=0.00135046f //x=6.645 \
 //y=0 //x2=6.465 //y2=0.865
cc_47 ( N_GND_M3_noxref_d N_noxref_4_c_463_n ) capacitor c=0.00220047f \
 //x=6.54 //y=0.865 //x2=6.465 //y2=0.865
cc_48 ( N_GND_M3_noxref_d N_noxref_4_c_465_n ) capacitor c=0.00255985f \
 //x=6.54 //y=0.865 //x2=6.465 //y2=1.21
cc_49 ( N_GND_c_3_p N_noxref_4_c_466_n ) capacitor c=0.0018059f //x=5.55 //y=0 \
 //x2=6.465 //y2=1.52
cc_50 ( N_GND_c_3_p N_noxref_4_c_467_n ) capacitor c=0.0114883f //x=5.55 //y=0 \
 //x2=6.465 //y2=1.915
cc_51 ( N_GND_M3_noxref_d N_noxref_4_c_468_n ) capacitor c=0.0131326f //x=6.54 \
 //y=0.865 //x2=6.84 //y2=0.71
cc_52 ( N_GND_M3_noxref_d N_noxref_4_c_469_n ) capacitor c=0.00193127f \
 //x=6.54 //y=0.865 //x2=6.84 //y2=1.365
cc_53 ( N_GND_c_53_p N_noxref_4_c_470_n ) capacitor c=0.00130622f //x=8.71 \
 //y=0 //x2=6.995 //y2=0.865
cc_54 ( N_GND_M3_noxref_d N_noxref_4_c_470_n ) capacitor c=0.00257848f \
 //x=6.54 //y=0.865 //x2=6.995 //y2=0.865
cc_55 ( N_GND_M3_noxref_d N_noxref_4_c_472_n ) capacitor c=0.00255985f \
 //x=6.54 //y=0.865 //x2=6.995 //y2=1.21
cc_56 ( N_GND_c_6_p N_noxref_4_M0_noxref_d ) capacitor c=0.00124113f //x=11.47 \
 //y=0 //x2=0.925 //y2=0.91
cc_57 ( N_GND_c_7_p N_noxref_4_M0_noxref_d ) capacitor c=0.0150482f //x=1.03 \
 //y=0.535 //x2=0.925 //y2=0.91
cc_58 ( N_GND_c_5_p N_noxref_4_M0_noxref_d ) capacitor c=2.29264e-19 //x=11.47 \
 //y=0 //x2=0.925 //y2=0.91
cc_59 ( N_GND_c_1_p N_noxref_4_M0_noxref_d ) capacitor c=0.0094373f //x=0.63 \
 //y=0 //x2=0.925 //y2=0.91
cc_60 ( N_GND_c_2_p N_noxref_4_M0_noxref_d ) capacitor c=0.00949241f //x=2.22 \
 //y=0 //x2=0.925 //y2=0.91
cc_61 ( N_GND_M0_noxref_s N_noxref_4_M0_noxref_d ) capacitor c=0.076995f \
 //x=0.495 //y=0.37 //x2=0.925 //y2=0.91
cc_62 ( N_GND_c_6_p N_noxref_5_c_595_n ) capacitor c=0.0412892f //x=11.47 \
 //y=0 //x2=9.875 //y2=2.96
cc_63 ( N_GND_c_33_p N_noxref_5_c_595_n ) capacitor c=0.00191528f //x=5.38 \
 //y=0 //x2=9.875 //y2=2.96
cc_64 ( N_GND_c_46_p N_noxref_5_c_595_n ) capacitor c=0.00233429f //x=6.645 \
 //y=0 //x2=9.875 //y2=2.96
cc_65 ( N_GND_c_53_p N_noxref_5_c_595_n ) capacitor c=0.00272473f //x=8.71 \
 //y=0 //x2=9.875 //y2=2.96
cc_66 ( N_GND_c_66_p N_noxref_5_c_595_n ) capacitor c=0.00230184f //x=9.975 \
 //y=0 //x2=9.875 //y2=2.96
cc_67 ( N_GND_c_3_p N_noxref_5_c_595_n ) capacitor c=0.0144849f //x=5.55 //y=0 \
 //x2=9.875 //y2=2.96
cc_68 ( N_GND_c_4_p N_noxref_5_c_595_n ) capacitor c=0.0144849f //x=8.88 //y=0 \
 //x2=9.875 //y2=2.96
cc_69 ( N_GND_c_6_p N_noxref_5_c_602_n ) capacitor c=0.00194856f //x=11.47 \
 //y=0 //x2=4.925 //y2=2.96
cc_70 ( N_GND_c_3_p N_noxref_5_c_603_n ) capacitor c=0.0462817f //x=5.55 //y=0 \
 //x2=4.725 //y2=1.655
cc_71 ( N_GND_c_2_p N_noxref_5_c_604_n ) capacitor c=0.00101801f //x=2.22 \
 //y=0 //x2=4.81 //y2=2.96
cc_72 ( N_GND_c_4_p N_noxref_5_c_605_n ) capacitor c=0.0179404f //x=8.88 //y=0 \
 //x2=9.99 //y2=2.08
cc_73 ( N_GND_c_66_p N_noxref_5_c_606_n ) capacitor c=0.00135046f //x=9.975 \
 //y=0 //x2=9.795 //y2=0.865
cc_74 ( N_GND_M5_noxref_d N_noxref_5_c_606_n ) capacitor c=0.00220047f \
 //x=9.87 //y=0.865 //x2=9.795 //y2=0.865
cc_75 ( N_GND_M5_noxref_d N_noxref_5_c_608_n ) capacitor c=0.00255985f \
 //x=9.87 //y=0.865 //x2=9.795 //y2=1.21
cc_76 ( N_GND_c_4_p N_noxref_5_c_609_n ) capacitor c=0.0018059f //x=8.88 //y=0 \
 //x2=9.795 //y2=1.52
cc_77 ( N_GND_c_4_p N_noxref_5_c_610_n ) capacitor c=0.0114883f //x=8.88 //y=0 \
 //x2=9.795 //y2=1.915
cc_78 ( N_GND_M5_noxref_d N_noxref_5_c_611_n ) capacitor c=0.0131326f //x=9.87 \
 //y=0.865 //x2=10.17 //y2=0.71
cc_79 ( N_GND_M5_noxref_d N_noxref_5_c_612_n ) capacitor c=0.00193127f \
 //x=9.87 //y=0.865 //x2=10.17 //y2=1.365
cc_80 ( N_GND_c_5_p N_noxref_5_c_613_n ) capacitor c=0.00130622f //x=11.47 \
 //y=0 //x2=10.325 //y2=0.865
cc_81 ( N_GND_M5_noxref_d N_noxref_5_c_613_n ) capacitor c=0.00257848f \
 //x=9.87 //y=0.865 //x2=10.325 //y2=0.865
cc_82 ( N_GND_M5_noxref_d N_noxref_5_c_615_n ) capacitor c=0.00255985f \
 //x=9.87 //y=0.865 //x2=10.325 //y2=1.21
cc_83 ( N_GND_c_2_p N_noxref_5_M2_noxref_d ) capacitor c=8.58106e-19 //x=2.22 \
 //y=0 //x2=4.18 //y2=0.905
cc_84 ( N_GND_c_3_p N_noxref_5_M2_noxref_d ) capacitor c=0.00616547f //x=5.55 \
 //y=0 //x2=4.18 //y2=0.905
cc_85 ( N_GND_M1_noxref_d N_noxref_5_M2_noxref_d ) capacitor c=0.00143464f \
 //x=3.21 //y=0.865 //x2=4.18 //y2=0.905
cc_86 ( N_GND_c_6_p N_noxref_6_c_763_n ) capacitor c=0.0138525f //x=11.47 \
 //y=0 //x2=10.615 //y2=3.33
cc_87 ( N_GND_c_4_p N_noxref_6_c_764_n ) capacitor c=0.0462817f //x=8.88 //y=0 \
 //x2=8.055 //y2=1.655
cc_88 ( N_GND_c_3_p N_noxref_6_c_765_n ) capacitor c=9.64732e-19 //x=5.55 \
 //y=0 //x2=8.14 //y2=3.33
cc_89 ( N_GND_c_5_p N_noxref_6_c_766_n ) capacitor c=9.53263e-19 //x=11.47 \
 //y=0 //x2=10.73 //y2=2.08
cc_90 ( N_GND_c_4_p N_noxref_6_c_766_n ) capacitor c=9.2064e-19 //x=8.88 //y=0 \
 //x2=10.73 //y2=2.08
cc_91 ( N_GND_c_3_p N_noxref_6_M4_noxref_d ) capacitor c=8.58106e-19 //x=5.55 \
 //y=0 //x2=7.51 //y2=0.905
cc_92 ( N_GND_c_4_p N_noxref_6_M4_noxref_d ) capacitor c=0.00616547f //x=8.88 \
 //y=0 //x2=7.51 //y2=0.905
cc_93 ( N_GND_M3_noxref_d N_noxref_6_M4_noxref_d ) capacitor c=0.00143464f \
 //x=6.54 //y=0.865 //x2=7.51 //y2=0.905
cc_94 ( N_GND_c_2_p N_A0_c_918_n ) capacitor c=9.2064e-19 //x=2.22 //y=0 \
 //x2=4.07 //y2=2.08
cc_95 ( N_GND_c_3_p N_A0_c_918_n ) capacitor c=9.53263e-19 //x=5.55 //y=0 \
 //x2=4.07 //y2=2.08
cc_96 ( N_GND_M0_noxref_s N_noxref_8_c_986_n ) capacitor c=0.0013253f \
 //x=0.495 //y=0.37 //x2=2.915 //y2=1.495
cc_97 ( N_GND_c_6_p N_noxref_8_c_987_n ) capacitor c=0.00546052f //x=11.47 \
 //y=0 //x2=3.8 //y2=1.58
cc_98 ( N_GND_c_9_p N_noxref_8_c_987_n ) capacitor c=0.00112963f //x=3.315 \
 //y=0 //x2=3.8 //y2=1.58
cc_99 ( N_GND_c_33_p N_noxref_8_c_987_n ) capacitor c=0.0018242f //x=5.38 \
 //y=0 //x2=3.8 //y2=1.58
cc_100 ( N_GND_M1_noxref_d N_noxref_8_c_987_n ) capacitor c=0.00890221f \
 //x=3.21 //y=0.865 //x2=3.8 //y2=1.58
cc_101 ( N_GND_c_6_p N_noxref_8_c_991_n ) capacitor c=0.00293348f //x=11.47 \
 //y=0 //x2=3.885 //y2=0.615
cc_102 ( N_GND_c_33_p N_noxref_8_c_991_n ) capacitor c=0.0149357f //x=5.38 \
 //y=0 //x2=3.885 //y2=0.615
cc_103 ( N_GND_c_5_p N_noxref_8_c_991_n ) capacitor c=0.00145873f //x=11.47 \
 //y=0 //x2=3.885 //y2=0.615
cc_104 ( N_GND_M1_noxref_d N_noxref_8_c_991_n ) capacitor c=0.033812f //x=3.21 \
 //y=0.865 //x2=3.885 //y2=0.615
cc_105 ( N_GND_c_2_p N_noxref_8_c_995_n ) capacitor c=2.91423e-19 //x=2.22 \
 //y=0 //x2=3.885 //y2=1.495
cc_106 ( N_GND_c_6_p N_noxref_8_c_996_n ) capacitor c=0.0119856f //x=11.47 \
 //y=0 //x2=4.77 //y2=0.53
cc_107 ( N_GND_c_33_p N_noxref_8_c_996_n ) capacitor c=0.0375343f //x=5.38 \
 //y=0 //x2=4.77 //y2=0.53
cc_108 ( N_GND_c_5_p N_noxref_8_c_996_n ) capacitor c=0.00199095f //x=11.47 \
 //y=0 //x2=4.77 //y2=0.53
cc_109 ( N_GND_c_6_p N_noxref_8_c_999_n ) capacitor c=0.00282055f //x=11.47 \
 //y=0 //x2=4.855 //y2=0.615
cc_110 ( N_GND_c_33_p N_noxref_8_c_999_n ) capacitor c=0.0147946f //x=5.38 \
 //y=0 //x2=4.855 //y2=0.615
cc_111 ( N_GND_c_5_p N_noxref_8_c_999_n ) capacitor c=0.00145015f //x=11.47 \
 //y=0 //x2=4.855 //y2=0.615
cc_112 ( N_GND_c_3_p N_noxref_8_c_999_n ) capacitor c=0.0431718f //x=5.55 \
 //y=0 //x2=4.855 //y2=0.615
cc_113 ( N_GND_c_6_p N_noxref_8_M1_noxref_s ) capacitor c=0.00282937f \
 //x=11.47 //y=0 //x2=2.78 //y2=0.365
cc_114 ( N_GND_c_114_p N_noxref_8_M1_noxref_s ) capacitor c=0.0013253f //x=1.6 \
 //y=0.45 //x2=2.78 //y2=0.365
cc_115 ( N_GND_c_9_p N_noxref_8_M1_noxref_s ) capacitor c=0.0148639f //x=3.315 \
 //y=0 //x2=2.78 //y2=0.365
cc_116 ( N_GND_c_5_p N_noxref_8_M1_noxref_s ) capacitor c=0.00145873f \
 //x=11.47 //y=0 //x2=2.78 //y2=0.365
cc_117 ( N_GND_c_2_p N_noxref_8_M1_noxref_s ) capacitor c=0.058339f //x=2.22 \
 //y=0 //x2=2.78 //y2=0.365
cc_118 ( N_GND_c_3_p N_noxref_8_M1_noxref_s ) capacitor c=0.00198043f //x=5.55 \
 //y=0 //x2=2.78 //y2=0.365
cc_119 ( N_GND_M1_noxref_d N_noxref_8_M1_noxref_s ) capacitor c=0.0334197f \
 //x=3.21 //y=0.865 //x2=2.78 //y2=0.365
cc_120 ( N_GND_c_3_p N_A1_c_1043_n ) capacitor c=9.2064e-19 //x=5.55 //y=0 \
 //x2=7.4 //y2=2.08
cc_121 ( N_GND_c_4_p N_A1_c_1043_n ) capacitor c=9.53263e-19 //x=8.88 //y=0 \
 //x2=7.4 //y2=2.08
cc_122 ( N_GND_c_6_p N_noxref_10_c_1112_n ) capacitor c=0.00542069f //x=11.47 \
 //y=0 //x2=7.13 //y2=1.58
cc_123 ( N_GND_c_46_p N_noxref_10_c_1112_n ) capacitor c=0.00112963f //x=6.645 \
 //y=0 //x2=7.13 //y2=1.58
cc_124 ( N_GND_c_53_p N_noxref_10_c_1112_n ) capacitor c=0.00182382f //x=8.71 \
 //y=0 //x2=7.13 //y2=1.58
cc_125 ( N_GND_M3_noxref_d N_noxref_10_c_1112_n ) capacitor c=0.00890129f \
 //x=6.54 //y=0.865 //x2=7.13 //y2=1.58
cc_126 ( N_GND_c_6_p N_noxref_10_c_1116_n ) capacitor c=0.00282937f //x=11.47 \
 //y=0 //x2=7.215 //y2=0.615
cc_127 ( N_GND_c_53_p N_noxref_10_c_1116_n ) capacitor c=0.0148639f //x=8.71 \
 //y=0 //x2=7.215 //y2=0.615
cc_128 ( N_GND_c_5_p N_noxref_10_c_1116_n ) capacitor c=0.00145873f //x=11.47 \
 //y=0 //x2=7.215 //y2=0.615
cc_129 ( N_GND_M3_noxref_d N_noxref_10_c_1116_n ) capacitor c=0.033812f \
 //x=6.54 //y=0.865 //x2=7.215 //y2=0.615
cc_130 ( N_GND_c_3_p N_noxref_10_c_1120_n ) capacitor c=2.91423e-19 //x=5.55 \
 //y=0 //x2=7.215 //y2=1.495
cc_131 ( N_GND_c_6_p N_noxref_10_c_1121_n ) capacitor c=0.0116329f //x=11.47 \
 //y=0 //x2=8.1 //y2=0.53
cc_132 ( N_GND_c_53_p N_noxref_10_c_1121_n ) capacitor c=0.0375167f //x=8.71 \
 //y=0 //x2=8.1 //y2=0.53
cc_133 ( N_GND_c_5_p N_noxref_10_c_1121_n ) capacitor c=0.00199095f //x=11.47 \
 //y=0 //x2=8.1 //y2=0.53
cc_134 ( N_GND_c_6_p N_noxref_10_c_1124_n ) capacitor c=0.00282863f //x=11.47 \
 //y=0 //x2=8.185 //y2=0.615
cc_135 ( N_GND_c_53_p N_noxref_10_c_1124_n ) capacitor c=0.0148003f //x=8.71 \
 //y=0 //x2=8.185 //y2=0.615
cc_136 ( N_GND_c_5_p N_noxref_10_c_1124_n ) capacitor c=0.00145015f //x=11.47 \
 //y=0 //x2=8.185 //y2=0.615
cc_137 ( N_GND_c_4_p N_noxref_10_c_1124_n ) capacitor c=0.0431718f //x=8.88 \
 //y=0 //x2=8.185 //y2=0.615
cc_138 ( N_GND_c_6_p N_noxref_10_M3_noxref_s ) capacitor c=0.00282937f \
 //x=11.47 //y=0 //x2=6.11 //y2=0.365
cc_139 ( N_GND_c_46_p N_noxref_10_M3_noxref_s ) capacitor c=0.0148639f \
 //x=6.645 //y=0 //x2=6.11 //y2=0.365
cc_140 ( N_GND_c_5_p N_noxref_10_M3_noxref_s ) capacitor c=0.00145873f \
 //x=11.47 //y=0 //x2=6.11 //y2=0.365
cc_141 ( N_GND_c_3_p N_noxref_10_M3_noxref_s ) capacitor c=0.058339f //x=5.55 \
 //y=0 //x2=6.11 //y2=0.365
cc_142 ( N_GND_c_4_p N_noxref_10_M3_noxref_s ) capacitor c=0.00198043f \
 //x=8.88 //y=0 //x2=6.11 //y2=0.365
cc_143 ( N_GND_M3_noxref_d N_noxref_10_M3_noxref_s ) capacitor c=0.0334197f \
 //x=6.54 //y=0.865 //x2=6.11 //y2=0.365
cc_144 ( N_GND_c_4_p Y ) capacitor c=9.64732e-19 //x=8.88 //y=0 //x2=11.47 \
 //y2=2.22
cc_145 ( N_GND_c_5_p N_Y_c_1168_n ) capacitor c=0.0468439f //x=11.47 //y=0 \
 //x2=11.385 //y2=1.655
cc_146 ( N_GND_c_5_p N_Y_M6_noxref_d ) capacitor c=0.00618259f //x=11.47 //y=0 \
 //x2=10.84 //y2=0.905
cc_147 ( N_GND_c_4_p N_Y_M6_noxref_d ) capacitor c=8.58106e-19 //x=8.88 //y=0 \
 //x2=10.84 //y2=0.905
cc_148 ( N_GND_M5_noxref_d N_Y_M6_noxref_d ) capacitor c=0.00143464f //x=9.87 \
 //y=0.865 //x2=10.84 //y2=0.905
cc_149 ( N_GND_c_6_p N_noxref_12_c_1232_n ) capacitor c=0.00546052f //x=11.47 \
 //y=0 //x2=10.46 //y2=1.58
cc_150 ( N_GND_c_66_p N_noxref_12_c_1232_n ) capacitor c=0.00112963f //x=9.975 \
 //y=0 //x2=10.46 //y2=1.58
cc_151 ( N_GND_c_5_p N_noxref_12_c_1232_n ) capacitor c=0.0018242f //x=11.47 \
 //y=0 //x2=10.46 //y2=1.58
cc_152 ( N_GND_M5_noxref_d N_noxref_12_c_1232_n ) capacitor c=0.00890221f \
 //x=9.87 //y=0.865 //x2=10.46 //y2=1.58
cc_153 ( N_GND_c_6_p N_noxref_12_c_1236_n ) capacitor c=0.00293276f //x=11.47 \
 //y=0 //x2=10.545 //y2=0.615
cc_154 ( N_GND_c_5_p N_noxref_12_c_1236_n ) capacitor c=0.0163939f //x=11.47 \
 //y=0 //x2=10.545 //y2=0.615
cc_155 ( N_GND_M5_noxref_d N_noxref_12_c_1236_n ) capacitor c=0.033812f \
 //x=9.87 //y=0.865 //x2=10.545 //y2=0.615
cc_156 ( N_GND_c_4_p N_noxref_12_c_1239_n ) capacitor c=2.91423e-19 //x=8.88 \
 //y=0 //x2=10.545 //y2=1.495
cc_157 ( N_GND_c_6_p N_noxref_12_c_1240_n ) capacitor c=0.0172036f //x=11.47 \
 //y=0 //x2=11.43 //y2=0.53
cc_158 ( N_GND_c_5_p N_noxref_12_c_1240_n ) capacitor c=0.0393339f //x=11.47 \
 //y=0 //x2=11.43 //y2=0.53
cc_159 ( N_GND_c_6_p N_noxref_12_c_1242_n ) capacitor c=0.00719615f //x=11.47 \
 //y=0 //x2=11.515 //y2=0.615
cc_160 ( N_GND_c_5_p N_noxref_12_c_1242_n ) capacitor c=0.0598581f //x=11.47 \
 //y=0 //x2=11.515 //y2=0.615
cc_161 ( N_GND_c_6_p N_noxref_12_M5_noxref_s ) capacitor c=0.00282937f \
 //x=11.47 //y=0 //x2=9.44 //y2=0.365
cc_162 ( N_GND_c_66_p N_noxref_12_M5_noxref_s ) capacitor c=0.0148639f \
 //x=9.975 //y=0 //x2=9.44 //y2=0.365
cc_163 ( N_GND_c_5_p N_noxref_12_M5_noxref_s ) capacitor c=0.00344356f \
 //x=11.47 //y=0 //x2=9.44 //y2=0.365
cc_164 ( N_GND_c_4_p N_noxref_12_M5_noxref_s ) capacitor c=0.058339f //x=8.88 \
 //y=0 //x2=9.44 //y2=0.365
cc_165 ( N_GND_M5_noxref_d N_noxref_12_M5_noxref_s ) capacitor c=0.0334197f \
 //x=9.87 //y=0.865 //x2=9.44 //y2=0.365
cc_166 ( N_VDD_c_171_p N_S_c_329_n ) capacitor c=0.00802055f //x=11.47 //y=7.4 \
 //x2=3.215 //y2=2.96
cc_167 ( N_VDD_c_171_p N_S_c_335_n ) capacitor c=0.0014834f //x=11.47 //y=7.4 \
 //x2=0.855 //y2=2.96
cc_168 ( N_VDD_M7_noxref_s N_S_c_335_n ) capacitor c=7.86045e-19 //x=0.54 \
 //y=5.02 //x2=0.855 //y2=2.96
cc_169 ( N_VDD_c_171_p N_S_c_337_n ) capacitor c=0.00161202f //x=11.47 //y=7.4 \
 //x2=0.74 //y2=2.085
cc_170 ( N_VDD_c_166_n N_S_c_337_n ) capacitor c=0.0276175f //x=0.74 //y=7.4 \
 //x2=0.74 //y2=2.085
cc_171 ( N_VDD_c_167_n N_S_c_337_n ) capacitor c=0.00144308f //x=2.22 //y=7.4 \
 //x2=0.74 //y2=2.085
cc_172 ( N_VDD_M7_noxref_s N_S_c_337_n ) capacitor c=0.00978508f //x=0.54 \
 //y=5.02 //x2=0.74 //y2=2.085
cc_173 ( N_VDD_c_171_p N_S_c_342_n ) capacitor c=0.00127895f //x=11.47 //y=7.4 \
 //x2=3.33 //y2=2.08
cc_174 ( N_VDD_c_179_p N_S_c_342_n ) capacitor c=2.63811e-19 //x=3.805 //y=7.4 \
 //x2=3.33 //y2=2.08
cc_175 ( N_VDD_c_167_n N_S_c_342_n ) capacitor c=0.0167437f //x=2.22 //y=7.4 \
 //x2=3.33 //y2=2.08
cc_176 ( N_VDD_c_181_p N_S_M7_noxref_g ) capacitor c=0.00748034f //x=1.47 \
 //y=7.4 //x2=0.895 //y2=6.02
cc_177 ( N_VDD_c_166_n N_S_M7_noxref_g ) capacitor c=0.0241676f //x=0.74 \
 //y=7.4 //x2=0.895 //y2=6.02
cc_178 ( N_VDD_M7_noxref_s N_S_M7_noxref_g ) capacitor c=0.0528676f //x=0.54 \
 //y=5.02 //x2=0.895 //y2=6.02
cc_179 ( N_VDD_c_181_p N_S_M8_noxref_g ) capacitor c=0.00697478f //x=1.47 \
 //y=7.4 //x2=1.335 //y2=6.02
cc_180 ( N_VDD_M8_noxref_d N_S_M8_noxref_g ) capacitor c=0.0528676f //x=1.41 \
 //y=5.02 //x2=1.335 //y2=6.02
cc_181 ( N_VDD_c_179_p N_S_M9_noxref_g ) capacitor c=0.00726866f //x=3.805 \
 //y=7.4 //x2=3.23 //y2=6.02
cc_182 ( N_VDD_M9_noxref_s N_S_M9_noxref_g ) capacitor c=0.054195f //x=2.875 \
 //y=5.02 //x2=3.23 //y2=6.02
cc_183 ( N_VDD_c_179_p N_S_M10_noxref_g ) capacitor c=0.00672952f //x=3.805 \
 //y=7.4 //x2=3.67 //y2=6.02
cc_184 ( N_VDD_M10_noxref_d N_S_M10_noxref_g ) capacitor c=0.015318f //x=3.745 \
 //y=5.02 //x2=3.67 //y2=6.02
cc_185 ( N_VDD_c_167_n N_S_c_381_n ) capacitor c=0.0110053f //x=2.22 //y=7.4 \
 //x2=1.26 //y2=4.79
cc_186 ( N_VDD_c_166_n N_S_c_382_n ) capacitor c=0.011132f //x=0.74 //y=7.4 \
 //x2=0.97 //y2=4.79
cc_187 ( N_VDD_M7_noxref_s N_S_c_382_n ) capacitor c=0.00527247f //x=0.54 \
 //y=5.02 //x2=0.97 //y2=4.79
cc_188 ( N_VDD_c_167_n N_S_c_384_n ) capacitor c=0.012849f //x=2.22 //y=7.4 \
 //x2=3.33 //y2=4.7
cc_189 ( N_VDD_c_171_p N_noxref_4_c_456_n ) capacitor c=0.0304223f //x=11.47 \
 //y=7.4 //x2=6.545 //y2=3.33
cc_190 ( N_VDD_c_167_n N_noxref_4_c_456_n ) capacitor c=0.0069465f //x=2.22 \
 //y=7.4 //x2=6.545 //y2=3.33
cc_191 ( N_VDD_c_168_n N_noxref_4_c_456_n ) capacitor c=0.0069465f //x=5.55 \
 //y=7.4 //x2=6.545 //y2=3.33
cc_192 ( N_VDD_M8_noxref_d N_noxref_4_c_456_n ) capacitor c=5.17699e-19 \
 //x=1.41 //y=5.02 //x2=6.545 //y2=3.33
cc_193 ( N_VDD_M9_noxref_s N_noxref_4_c_456_n ) capacitor c=0.00204557f \
 //x=2.875 //y=5.02 //x2=6.545 //y2=3.33
cc_194 ( N_VDD_M12_noxref_d N_noxref_4_c_456_n ) capacitor c=3.2832e-19 \
 //x=4.625 //y=5.02 //x2=6.545 //y2=3.33
cc_195 ( N_VDD_M13_noxref_s N_noxref_4_c_456_n ) capacitor c=0.00204557f \
 //x=6.205 //y=5.02 //x2=6.545 //y2=3.33
cc_196 ( N_VDD_c_171_p N_noxref_4_c_486_n ) capacitor c=0.00163324f //x=11.47 \
 //y=7.4 //x2=1.595 //y2=3.33
cc_197 ( N_VDD_M8_noxref_d N_noxref_4_c_486_n ) capacitor c=7.33386e-19 \
 //x=1.41 //y=5.02 //x2=1.595 //y2=3.33
cc_198 ( N_VDD_c_171_p N_noxref_4_c_488_n ) capacitor c=0.00128923f //x=11.47 \
 //y=7.4 //x2=1.395 //y2=4.58
cc_199 ( N_VDD_c_181_p N_noxref_4_c_488_n ) capacitor c=8.8179e-19 //x=1.47 \
 //y=7.4 //x2=1.395 //y2=4.58
cc_200 ( N_VDD_M8_noxref_d N_noxref_4_c_488_n ) capacitor c=0.00627485f \
 //x=1.41 //y=5.02 //x2=1.395 //y2=4.58
cc_201 ( N_VDD_c_166_n N_noxref_4_c_491_n ) capacitor c=0.0179238f //x=0.74 \
 //y=7.4 //x2=1.2 //y2=4.58
cc_202 ( N_VDD_c_166_n N_noxref_4_c_461_n ) capacitor c=4.80934e-19 //x=0.74 \
 //y=7.4 //x2=1.48 //y2=3.33
cc_203 ( N_VDD_c_167_n N_noxref_4_c_461_n ) capacitor c=0.0228983f //x=2.22 \
 //y=7.4 //x2=1.48 //y2=3.33
cc_204 ( N_VDD_c_171_p N_noxref_4_c_462_n ) capacitor c=0.00127831f //x=11.47 \
 //y=7.4 //x2=6.66 //y2=2.08
cc_205 ( N_VDD_c_210_p N_noxref_4_c_462_n ) capacitor c=2.63811e-19 //x=7.135 \
 //y=7.4 //x2=6.66 //y2=2.08
cc_206 ( N_VDD_c_168_n N_noxref_4_c_462_n ) capacitor c=0.0167437f //x=5.55 \
 //y=7.4 //x2=6.66 //y2=2.08
cc_207 ( N_VDD_c_210_p N_noxref_4_M13_noxref_g ) capacitor c=0.00726866f \
 //x=7.135 //y=7.4 //x2=6.56 //y2=6.02
cc_208 ( N_VDD_M13_noxref_s N_noxref_4_M13_noxref_g ) capacitor c=0.054195f \
 //x=6.205 //y=5.02 //x2=6.56 //y2=6.02
cc_209 ( N_VDD_c_210_p N_noxref_4_M14_noxref_g ) capacitor c=0.00672952f \
 //x=7.135 //y=7.4 //x2=7 //y2=6.02
cc_210 ( N_VDD_M14_noxref_d N_noxref_4_M14_noxref_g ) capacitor c=0.015318f \
 //x=7.075 //y=5.02 //x2=7 //y2=6.02
cc_211 ( N_VDD_c_168_n N_noxref_4_c_501_n ) capacitor c=0.0150435f //x=5.55 \
 //y=7.4 //x2=6.66 //y2=4.7
cc_212 ( N_VDD_c_171_p N_noxref_4_M7_noxref_d ) capacitor c=0.00585331f \
 //x=11.47 //y=7.4 //x2=0.97 //y2=5.02
cc_213 ( N_VDD_c_181_p N_noxref_4_M7_noxref_d ) capacitor c=0.0139004f \
 //x=1.47 //y=7.4 //x2=0.97 //y2=5.02
cc_214 ( N_VDD_c_167_n N_noxref_4_M7_noxref_d ) capacitor c=0.0204591f \
 //x=2.22 //y=7.4 //x2=0.97 //y2=5.02
cc_215 ( N_VDD_c_170_n N_noxref_4_M7_noxref_d ) capacitor c=0.00135976f \
 //x=11.47 //y=7.4 //x2=0.97 //y2=5.02
cc_216 ( N_VDD_M7_noxref_s N_noxref_4_M7_noxref_d ) capacitor c=0.0843065f \
 //x=0.54 //y=5.02 //x2=0.97 //y2=5.02
cc_217 ( N_VDD_M8_noxref_d N_noxref_4_M7_noxref_d ) capacitor c=0.0832641f \
 //x=1.41 //y=5.02 //x2=0.97 //y2=5.02
cc_218 ( N_VDD_c_171_p N_noxref_5_c_595_n ) capacitor c=0.016877f //x=11.47 \
 //y=7.4 //x2=9.875 //y2=2.96
cc_219 ( N_VDD_c_171_p N_noxref_5_c_620_n ) capacitor c=0.00471288f //x=11.47 \
 //y=7.4 //x2=4.245 //y2=5.2
cc_220 ( N_VDD_c_179_p N_noxref_5_c_620_n ) capacitor c=4.3394e-19 //x=3.805 \
 //y=7.4 //x2=4.245 //y2=5.2
cc_221 ( N_VDD_c_226_p N_noxref_5_c_620_n ) capacitor c=4.3394e-19 //x=4.685 \
 //y=7.4 //x2=4.245 //y2=5.2
cc_222 ( N_VDD_M10_noxref_d N_noxref_5_c_620_n ) capacitor c=0.0129494f \
 //x=3.745 //y=5.02 //x2=4.245 //y2=5.2
cc_223 ( N_VDD_c_167_n N_noxref_5_c_624_n ) capacitor c=0.00985474f //x=2.22 \
 //y=7.4 //x2=3.535 //y2=5.2
cc_224 ( N_VDD_M9_noxref_s N_noxref_5_c_624_n ) capacitor c=0.087833f \
 //x=2.875 //y=5.02 //x2=3.535 //y2=5.2
cc_225 ( N_VDD_c_171_p N_noxref_5_c_626_n ) capacitor c=0.00316347f //x=11.47 \
 //y=7.4 //x2=4.725 //y2=5.2
cc_226 ( N_VDD_c_226_p N_noxref_5_c_626_n ) capacitor c=7.21492e-19 //x=4.685 \
 //y=7.4 //x2=4.725 //y2=5.2
cc_227 ( N_VDD_M12_noxref_d N_noxref_5_c_626_n ) capacitor c=0.0164758f \
 //x=4.625 //y=5.02 //x2=4.725 //y2=5.2
cc_228 ( N_VDD_M13_noxref_s N_noxref_5_c_626_n ) capacitor c=2.44532e-19 \
 //x=6.205 //y=5.02 //x2=4.725 //y2=5.2
cc_229 ( N_VDD_c_167_n N_noxref_5_c_604_n ) capacitor c=0.00159771f //x=2.22 \
 //y=7.4 //x2=4.81 //y2=2.96
cc_230 ( N_VDD_c_168_n N_noxref_5_c_604_n ) capacitor c=0.0462955f //x=5.55 \
 //y=7.4 //x2=4.81 //y2=2.96
cc_231 ( N_VDD_c_171_p N_noxref_5_c_605_n ) capacitor c=0.00127895f //x=11.47 \
 //y=7.4 //x2=9.99 //y2=2.08
cc_232 ( N_VDD_c_237_p N_noxref_5_c_605_n ) capacitor c=2.63811e-19 //x=10.465 \
 //y=7.4 //x2=9.99 //y2=2.08
cc_233 ( N_VDD_c_169_n N_noxref_5_c_605_n ) capacitor c=0.0167437f //x=8.88 \
 //y=7.4 //x2=9.99 //y2=2.08
cc_234 ( N_VDD_c_237_p N_noxref_5_M17_noxref_g ) capacitor c=0.00726866f \
 //x=10.465 //y=7.4 //x2=9.89 //y2=6.02
cc_235 ( N_VDD_M17_noxref_s N_noxref_5_M17_noxref_g ) capacitor c=0.054195f \
 //x=9.535 //y=5.02 //x2=9.89 //y2=6.02
cc_236 ( N_VDD_c_237_p N_noxref_5_M18_noxref_g ) capacitor c=0.00672952f \
 //x=10.465 //y=7.4 //x2=10.33 //y2=6.02
cc_237 ( N_VDD_M18_noxref_d N_noxref_5_M18_noxref_g ) capacitor c=0.015318f \
 //x=10.405 //y=5.02 //x2=10.33 //y2=6.02
cc_238 ( N_VDD_c_169_n N_noxref_5_c_639_n ) capacitor c=0.0150435f //x=8.88 \
 //y=7.4 //x2=9.99 //y2=4.7
cc_239 ( N_VDD_c_171_p N_noxref_5_M9_noxref_d ) capacitor c=0.00574621f \
 //x=11.47 //y=7.4 //x2=3.305 //y2=5.02
cc_240 ( N_VDD_c_179_p N_noxref_5_M9_noxref_d ) capacitor c=0.0138103f \
 //x=3.805 //y=7.4 //x2=3.305 //y2=5.02
cc_241 ( N_VDD_c_168_n N_noxref_5_M9_noxref_d ) capacitor c=6.94454e-19 \
 //x=5.55 //y=7.4 //x2=3.305 //y2=5.02
cc_242 ( N_VDD_c_170_n N_noxref_5_M9_noxref_d ) capacitor c=0.00135231f \
 //x=11.47 //y=7.4 //x2=3.305 //y2=5.02
cc_243 ( N_VDD_M10_noxref_d N_noxref_5_M9_noxref_d ) capacitor c=0.0664752f \
 //x=3.745 //y=5.02 //x2=3.305 //y2=5.02
cc_244 ( N_VDD_c_171_p N_noxref_5_M11_noxref_d ) capacitor c=0.00574621f \
 //x=11.47 //y=7.4 //x2=4.185 //y2=5.02
cc_245 ( N_VDD_c_226_p N_noxref_5_M11_noxref_d ) capacitor c=0.0138379f \
 //x=4.685 //y=7.4 //x2=4.185 //y2=5.02
cc_246 ( N_VDD_c_168_n N_noxref_5_M11_noxref_d ) capacitor c=0.0120541f \
 //x=5.55 //y=7.4 //x2=4.185 //y2=5.02
cc_247 ( N_VDD_c_170_n N_noxref_5_M11_noxref_d ) capacitor c=0.00135231f \
 //x=11.47 //y=7.4 //x2=4.185 //y2=5.02
cc_248 ( N_VDD_M9_noxref_s N_noxref_5_M11_noxref_d ) capacitor c=0.00111971f \
 //x=2.875 //y=5.02 //x2=4.185 //y2=5.02
cc_249 ( N_VDD_M10_noxref_d N_noxref_5_M11_noxref_d ) capacitor c=0.0664752f \
 //x=3.745 //y=5.02 //x2=4.185 //y2=5.02
cc_250 ( N_VDD_M12_noxref_d N_noxref_5_M11_noxref_d ) capacitor c=0.0664752f \
 //x=4.625 //y=5.02 //x2=4.185 //y2=5.02
cc_251 ( N_VDD_M13_noxref_s N_noxref_5_M11_noxref_d ) capacitor c=4.54516e-19 \
 //x=6.205 //y=5.02 //x2=4.185 //y2=5.02
cc_252 ( N_VDD_c_171_p N_noxref_6_c_763_n ) capacitor c=0.0155621f //x=11.47 \
 //y=7.4 //x2=10.615 //y2=3.33
cc_253 ( N_VDD_c_169_n N_noxref_6_c_763_n ) capacitor c=0.0069465f //x=8.88 \
 //y=7.4 //x2=10.615 //y2=3.33
cc_254 ( N_VDD_M17_noxref_s N_noxref_6_c_763_n ) capacitor c=0.00204557f \
 //x=9.535 //y=5.02 //x2=10.615 //y2=3.33
cc_255 ( N_VDD_c_171_p N_noxref_6_c_774_n ) capacitor c=0.00161874f //x=11.47 \
 //y=7.4 //x2=8.255 //y2=3.33
cc_256 ( N_VDD_M16_noxref_d N_noxref_6_c_774_n ) capacitor c=3.3085e-19 \
 //x=7.955 //y=5.02 //x2=8.255 //y2=3.33
cc_257 ( N_VDD_c_171_p N_noxref_6_c_776_n ) capacitor c=0.0047626f //x=11.47 \
 //y=7.4 //x2=7.575 //y2=5.2
cc_258 ( N_VDD_c_210_p N_noxref_6_c_776_n ) capacitor c=4.3394e-19 //x=7.135 \
 //y=7.4 //x2=7.575 //y2=5.2
cc_259 ( N_VDD_c_264_p N_noxref_6_c_776_n ) capacitor c=4.3394e-19 //x=8.015 \
 //y=7.4 //x2=7.575 //y2=5.2
cc_260 ( N_VDD_M14_noxref_d N_noxref_6_c_776_n ) capacitor c=0.0130143f \
 //x=7.075 //y=5.02 //x2=7.575 //y2=5.2
cc_261 ( N_VDD_c_168_n N_noxref_6_c_780_n ) capacitor c=0.00985474f //x=5.55 \
 //y=7.4 //x2=6.865 //y2=5.2
cc_262 ( N_VDD_M13_noxref_s N_noxref_6_c_780_n ) capacitor c=0.087833f \
 //x=6.205 //y=5.02 //x2=6.865 //y2=5.2
cc_263 ( N_VDD_c_171_p N_noxref_6_c_782_n ) capacitor c=0.00318278f //x=11.47 \
 //y=7.4 //x2=8.055 //y2=5.2
cc_264 ( N_VDD_c_264_p N_noxref_6_c_782_n ) capacitor c=7.21492e-19 //x=8.015 \
 //y=7.4 //x2=8.055 //y2=5.2
cc_265 ( N_VDD_M16_noxref_d N_noxref_6_c_782_n ) capacitor c=0.016468f \
 //x=7.955 //y=5.02 //x2=8.055 //y2=5.2
cc_266 ( N_VDD_M17_noxref_s N_noxref_6_c_782_n ) capacitor c=2.44532e-19 \
 //x=9.535 //y=5.02 //x2=8.055 //y2=5.2
cc_267 ( N_VDD_c_168_n N_noxref_6_c_765_n ) capacitor c=0.00151618f //x=5.55 \
 //y=7.4 //x2=8.14 //y2=3.33
cc_268 ( N_VDD_c_169_n N_noxref_6_c_765_n ) capacitor c=0.0462955f //x=8.88 \
 //y=7.4 //x2=8.14 //y2=3.33
cc_269 ( N_VDD_c_169_n N_noxref_6_c_766_n ) capacitor c=6.61004e-19 //x=8.88 \
 //y=7.4 //x2=10.73 //y2=2.08
cc_270 ( N_VDD_c_170_n N_noxref_6_c_766_n ) capacitor c=6.09526e-19 //x=11.47 \
 //y=7.4 //x2=10.73 //y2=2.08
cc_271 ( N_VDD_c_276_p N_noxref_6_M19_noxref_g ) capacitor c=0.00673971f \
 //x=11.345 //y=7.4 //x2=10.77 //y2=6.02
cc_272 ( N_VDD_M18_noxref_d N_noxref_6_M19_noxref_g ) capacitor c=0.015318f \
 //x=10.405 //y=5.02 //x2=10.77 //y2=6.02
cc_273 ( N_VDD_c_276_p N_noxref_6_M20_noxref_g ) capacitor c=0.00672952f \
 //x=11.345 //y=7.4 //x2=11.21 //y2=6.02
cc_274 ( N_VDD_c_170_n N_noxref_6_M20_noxref_g ) capacitor c=0.024326f \
 //x=11.47 //y=7.4 //x2=11.21 //y2=6.02
cc_275 ( N_VDD_M20_noxref_d N_noxref_6_M20_noxref_g ) capacitor c=0.0430452f \
 //x=11.285 //y=5.02 //x2=11.21 //y2=6.02
cc_276 ( N_VDD_c_171_p N_noxref_6_M13_noxref_d ) capacitor c=0.00577138f \
 //x=11.47 //y=7.4 //x2=6.635 //y2=5.02
cc_277 ( N_VDD_c_210_p N_noxref_6_M13_noxref_d ) capacitor c=0.0138103f \
 //x=7.135 //y=7.4 //x2=6.635 //y2=5.02
cc_278 ( N_VDD_c_169_n N_noxref_6_M13_noxref_d ) capacitor c=6.94454e-19 \
 //x=8.88 //y=7.4 //x2=6.635 //y2=5.02
cc_279 ( N_VDD_c_170_n N_noxref_6_M13_noxref_d ) capacitor c=0.00135231f \
 //x=11.47 //y=7.4 //x2=6.635 //y2=5.02
cc_280 ( N_VDD_M14_noxref_d N_noxref_6_M13_noxref_d ) capacitor c=0.0664752f \
 //x=7.075 //y=5.02 //x2=6.635 //y2=5.02
cc_281 ( N_VDD_c_171_p N_noxref_6_M15_noxref_d ) capacitor c=0.00582647f \
 //x=11.47 //y=7.4 //x2=7.515 //y2=5.02
cc_282 ( N_VDD_c_264_p N_noxref_6_M15_noxref_d ) capacitor c=0.0138379f \
 //x=8.015 //y=7.4 //x2=7.515 //y2=5.02
cc_283 ( N_VDD_c_169_n N_noxref_6_M15_noxref_d ) capacitor c=0.0120541f \
 //x=8.88 //y=7.4 //x2=7.515 //y2=5.02
cc_284 ( N_VDD_c_170_n N_noxref_6_M15_noxref_d ) capacitor c=0.00135231f \
 //x=11.47 //y=7.4 //x2=7.515 //y2=5.02
cc_285 ( N_VDD_M13_noxref_s N_noxref_6_M15_noxref_d ) capacitor c=0.00111971f \
 //x=6.205 //y=5.02 //x2=7.515 //y2=5.02
cc_286 ( N_VDD_M14_noxref_d N_noxref_6_M15_noxref_d ) capacitor c=0.0664752f \
 //x=7.075 //y=5.02 //x2=7.515 //y2=5.02
cc_287 ( N_VDD_M16_noxref_d N_noxref_6_M15_noxref_d ) capacitor c=0.0664752f \
 //x=7.955 //y=5.02 //x2=7.515 //y2=5.02
cc_288 ( N_VDD_M17_noxref_s N_noxref_6_M15_noxref_d ) capacitor c=4.54516e-19 \
 //x=9.535 //y=5.02 //x2=7.515 //y2=5.02
cc_289 ( N_VDD_c_167_n N_A0_c_918_n ) capacitor c=6.61004e-19 //x=2.22 //y=7.4 \
 //x2=4.07 //y2=2.08
cc_290 ( N_VDD_c_168_n N_A0_c_918_n ) capacitor c=6.09526e-19 //x=5.55 //y=7.4 \
 //x2=4.07 //y2=2.08
cc_291 ( N_VDD_c_226_p N_A0_M11_noxref_g ) capacitor c=0.00673971f //x=4.685 \
 //y=7.4 //x2=4.11 //y2=6.02
cc_292 ( N_VDD_M10_noxref_d N_A0_M11_noxref_g ) capacitor c=0.015318f \
 //x=3.745 //y=5.02 //x2=4.11 //y2=6.02
cc_293 ( N_VDD_c_226_p N_A0_M12_noxref_g ) capacitor c=0.00672952f //x=4.685 \
 //y=7.4 //x2=4.55 //y2=6.02
cc_294 ( N_VDD_c_168_n N_A0_M12_noxref_g ) capacitor c=0.00864163f //x=5.55 \
 //y=7.4 //x2=4.55 //y2=6.02
cc_295 ( N_VDD_M12_noxref_d N_A0_M12_noxref_g ) capacitor c=0.0430452f \
 //x=4.625 //y=5.02 //x2=4.55 //y2=6.02
cc_296 ( N_VDD_c_168_n N_A1_c_1043_n ) capacitor c=6.61004e-19 //x=5.55 \
 //y=7.4 //x2=7.4 //y2=2.08
cc_297 ( N_VDD_c_169_n N_A1_c_1043_n ) capacitor c=6.09526e-19 //x=8.88 \
 //y=7.4 //x2=7.4 //y2=2.08
cc_298 ( N_VDD_c_264_p N_A1_M15_noxref_g ) capacitor c=0.00673971f //x=8.015 \
 //y=7.4 //x2=7.44 //y2=6.02
cc_299 ( N_VDD_M14_noxref_d N_A1_M15_noxref_g ) capacitor c=0.015318f \
 //x=7.075 //y=5.02 //x2=7.44 //y2=6.02
cc_300 ( N_VDD_c_264_p N_A1_M16_noxref_g ) capacitor c=0.00672952f //x=8.015 \
 //y=7.4 //x2=7.88 //y2=6.02
cc_301 ( N_VDD_c_169_n N_A1_M16_noxref_g ) capacitor c=0.00864163f //x=8.88 \
 //y=7.4 //x2=7.88 //y2=6.02
cc_302 ( N_VDD_M16_noxref_d N_A1_M16_noxref_g ) capacitor c=0.0430452f \
 //x=7.955 //y=5.02 //x2=7.88 //y2=6.02
cc_303 ( N_VDD_c_169_n Y ) capacitor c=0.00151618f //x=8.88 //y=7.4 //x2=11.47 \
 //y2=2.22
cc_304 ( N_VDD_c_170_n Y ) capacitor c=0.0468798f //x=11.47 //y=7.4 //x2=11.47 \
 //y2=2.22
cc_305 ( N_VDD_c_171_p N_Y_c_1174_n ) capacitor c=0.00471133f //x=11.47 \
 //y=7.4 //x2=10.905 //y2=5.2
cc_306 ( N_VDD_c_237_p N_Y_c_1174_n ) capacitor c=4.3394e-19 //x=10.465 \
 //y=7.4 //x2=10.905 //y2=5.2
cc_307 ( N_VDD_c_276_p N_Y_c_1174_n ) capacitor c=4.3394e-19 //x=11.345 \
 //y=7.4 //x2=10.905 //y2=5.2
cc_308 ( N_VDD_M18_noxref_d N_Y_c_1174_n ) capacitor c=0.0129484f //x=10.405 \
 //y=5.02 //x2=10.905 //y2=5.2
cc_309 ( N_VDD_c_169_n N_Y_c_1178_n ) capacitor c=0.00985474f //x=8.88 //y=7.4 \
 //x2=10.195 //y2=5.2
cc_310 ( N_VDD_M17_noxref_s N_Y_c_1178_n ) capacitor c=0.087833f //x=9.535 \
 //y=5.02 //x2=10.195 //y2=5.2
cc_311 ( N_VDD_c_171_p N_Y_c_1180_n ) capacitor c=0.00445413f //x=11.47 \
 //y=7.4 //x2=11.385 //y2=5.2
cc_312 ( N_VDD_c_276_p N_Y_c_1180_n ) capacitor c=7.21492e-19 //x=11.345 \
 //y=7.4 //x2=11.385 //y2=5.2
cc_313 ( N_VDD_M20_noxref_d N_Y_c_1180_n ) capacitor c=0.0165872f //x=11.285 \
 //y=5.02 //x2=11.385 //y2=5.2
cc_314 ( N_VDD_c_171_p N_Y_M17_noxref_d ) capacitor c=0.00574621f //x=11.47 \
 //y=7.4 //x2=9.965 //y2=5.02
cc_315 ( N_VDD_c_237_p N_Y_M17_noxref_d ) capacitor c=0.0138103f //x=10.465 \
 //y=7.4 //x2=9.965 //y2=5.02
cc_316 ( N_VDD_c_170_n N_Y_M17_noxref_d ) capacitor c=0.00204676f //x=11.47 \
 //y=7.4 //x2=9.965 //y2=5.02
cc_317 ( N_VDD_M18_noxref_d N_Y_M17_noxref_d ) capacitor c=0.0664752f \
 //x=10.405 //y=5.02 //x2=9.965 //y2=5.02
cc_318 ( N_VDD_c_171_p N_Y_M19_noxref_d ) capacitor c=0.00706239f //x=11.47 \
 //y=7.4 //x2=10.845 //y2=5.02
cc_319 ( N_VDD_c_276_p N_Y_M19_noxref_d ) capacitor c=0.0138379f //x=11.345 \
 //y=7.4 //x2=10.845 //y2=5.02
cc_320 ( N_VDD_c_170_n N_Y_M19_noxref_d ) capacitor c=0.0136712f //x=11.47 \
 //y=7.4 //x2=10.845 //y2=5.02
cc_321 ( N_VDD_M17_noxref_s N_Y_M19_noxref_d ) capacitor c=0.00111971f \
 //x=9.535 //y=5.02 //x2=10.845 //y2=5.02
cc_322 ( N_VDD_M18_noxref_d N_Y_M19_noxref_d ) capacitor c=0.0664752f \
 //x=10.405 //y=5.02 //x2=10.845 //y2=5.02
cc_323 ( N_VDD_M20_noxref_d N_Y_M19_noxref_d ) capacitor c=0.0664752f \
 //x=11.285 //y=5.02 //x2=10.845 //y2=5.02
cc_324 ( N_S_c_329_n N_noxref_4_c_456_n ) capacitor c=0.173644f //x=3.215 \
 //y=2.96 //x2=6.545 //y2=3.33
cc_325 ( N_S_c_342_n N_noxref_4_c_456_n ) capacitor c=0.0260635f //x=3.33 \
 //y=2.08 //x2=6.545 //y2=3.33
cc_326 ( N_S_c_329_n N_noxref_4_c_486_n ) capacitor c=0.029061f //x=3.215 \
 //y=2.96 //x2=1.595 //y2=3.33
cc_327 ( N_S_c_337_n N_noxref_4_c_486_n ) capacitor c=0.00599141f //x=0.74 \
 //y=2.085 //x2=1.595 //y2=3.33
cc_328 ( N_S_c_342_n N_noxref_4_c_486_n ) capacitor c=5.96166e-19 //x=3.33 \
 //y=2.08 //x2=1.595 //y2=3.33
cc_329 ( N_S_c_342_n N_noxref_4_c_458_n ) capacitor c=0.0138358f //x=3.33 \
 //y=2.08 //x2=1.395 //y2=2.08
cc_330 ( N_S_c_391_p N_noxref_4_c_458_n ) capacitor c=0.0023507f //x=1.225 \
 //y=1.41 //x2=1.395 //y2=2.08
cc_331 ( N_S_c_329_n N_noxref_4_c_515_n ) capacitor c=0.00763858f //x=3.215 \
 //y=2.96 //x2=1.195 //y2=2.08
cc_332 ( N_S_c_359_n N_noxref_4_c_515_n ) capacitor c=0.0167852f //x=0.74 \
 //y=2.085 //x2=1.195 //y2=2.08
cc_333 ( N_S_c_381_n N_noxref_4_c_488_n ) capacitor c=0.0101013f //x=1.26 \
 //y=4.79 //x2=1.395 //y2=4.58
cc_334 ( N_S_c_329_n N_noxref_4_c_491_n ) capacitor c=0.00318102f //x=3.215 \
 //y=2.96 //x2=1.2 //y2=4.58
cc_335 ( N_S_c_337_n N_noxref_4_c_491_n ) capacitor c=0.0250789f //x=0.74 \
 //y=2.085 //x2=1.2 //y2=4.58
cc_336 ( N_S_c_382_n N_noxref_4_c_491_n ) capacitor c=0.00962086f //x=0.97 \
 //y=4.79 //x2=1.2 //y2=4.58
cc_337 ( N_S_c_329_n N_noxref_4_c_461_n ) capacitor c=0.025579f //x=3.215 \
 //y=2.96 //x2=1.48 //y2=3.33
cc_338 ( N_S_c_335_n N_noxref_4_c_461_n ) capacitor c=0.00101501f //x=0.855 \
 //y=2.96 //x2=1.48 //y2=3.33
cc_339 ( N_S_c_337_n N_noxref_4_c_461_n ) capacitor c=0.0685954f //x=0.74 \
 //y=2.085 //x2=1.48 //y2=3.33
cc_340 ( N_S_c_359_n N_noxref_4_c_461_n ) capacitor c=8.49451e-19 //x=0.74 \
 //y=2.085 //x2=1.48 //y2=3.33
cc_341 ( N_S_c_337_n N_noxref_4_M0_noxref_d ) capacitor c=0.0175773f //x=0.74 \
 //y=2.085 //x2=0.925 //y2=0.91
cc_342 ( N_S_c_343_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218556f //x=0.85 \
 //y=0.91 //x2=0.925 //y2=0.91
cc_343 ( N_S_c_404_p N_noxref_4_M0_noxref_d ) capacitor c=0.00347355f //x=0.85 \
 //y=1.255 //x2=0.925 //y2=0.91
cc_344 ( N_S_c_405_p N_noxref_4_M0_noxref_d ) capacitor c=0.00742431f //x=0.85 \
 //y=1.565 //x2=0.925 //y2=0.91
cc_345 ( N_S_c_345_n N_noxref_4_M0_noxref_d ) capacitor c=0.00957707f //x=0.85 \
 //y=1.92 //x2=0.925 //y2=0.91
cc_346 ( N_S_c_346_n N_noxref_4_M0_noxref_d ) capacitor c=0.00220879f \
 //x=1.225 //y=0.755 //x2=0.925 //y2=0.91
cc_347 ( N_S_c_391_p N_noxref_4_M0_noxref_d ) capacitor c=0.0138447f //x=1.225 \
 //y=1.41 //x2=0.925 //y2=0.91
cc_348 ( N_S_c_347_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218624f //x=1.38 \
 //y=0.91 //x2=0.925 //y2=0.91
cc_349 ( N_S_c_349_n N_noxref_4_M0_noxref_d ) capacitor c=0.00601286f //x=1.38 \
 //y=1.255 //x2=0.925 //y2=0.91
cc_350 ( N_S_M7_noxref_g N_noxref_4_M7_noxref_d ) capacitor c=0.0219309f \
 //x=0.895 //y=6.02 //x2=0.97 //y2=5.02
cc_351 ( N_S_M8_noxref_g N_noxref_4_M7_noxref_d ) capacitor c=0.021902f \
 //x=1.335 //y=6.02 //x2=0.97 //y2=5.02
cc_352 ( N_S_c_381_n N_noxref_4_M7_noxref_d ) capacitor c=0.0148755f //x=1.26 \
 //y=4.79 //x2=0.97 //y2=5.02
cc_353 ( N_S_c_382_n N_noxref_4_M7_noxref_d ) capacitor c=0.00307344f //x=0.97 \
 //y=4.79 //x2=0.97 //y2=5.02
cc_354 ( N_S_c_329_n N_noxref_5_c_602_n ) capacitor c=0.0114735f //x=3.215 \
 //y=2.96 //x2=4.925 //y2=2.96
cc_355 ( N_S_M10_noxref_g N_noxref_5_c_620_n ) capacitor c=0.0192312f //x=3.67 \
 //y=6.02 //x2=4.245 //y2=5.2
cc_356 ( N_S_c_342_n N_noxref_5_c_624_n ) capacitor c=0.0056116f //x=3.33 \
 //y=2.08 //x2=3.535 //y2=5.2
cc_357 ( N_S_M9_noxref_g N_noxref_5_c_624_n ) capacitor c=0.0177326f //x=3.23 \
 //y=6.02 //x2=3.535 //y2=5.2
cc_358 ( N_S_c_384_n N_noxref_5_c_624_n ) capacitor c=0.00589848f //x=3.33 \
 //y=4.7 //x2=3.535 //y2=5.2
cc_359 ( N_S_c_342_n N_noxref_5_c_604_n ) capacitor c=0.0036353f //x=3.33 \
 //y=2.08 //x2=4.81 //y2=2.96
cc_360 ( N_S_M10_noxref_g N_noxref_5_M9_noxref_d ) capacitor c=0.0173476f \
 //x=3.67 //y=6.02 //x2=3.305 //y2=5.02
cc_361 ( N_S_c_342_n N_A0_c_927_n ) capacitor c=0.00400249f //x=3.33 //y=2.08 \
 //x2=4.07 //y2=4.535
cc_362 ( N_S_c_384_n N_A0_c_927_n ) capacitor c=0.00417994f //x=3.33 //y=4.7 \
 //x2=4.07 //y2=4.535
cc_363 ( N_S_c_329_n N_A0_c_918_n ) capacitor c=0.00317669f //x=3.215 //y=2.96 \
 //x2=4.07 //y2=2.08
cc_364 ( N_S_c_342_n N_A0_c_918_n ) capacitor c=0.0845408f //x=3.33 //y=2.08 \
 //x2=4.07 //y2=2.08
cc_365 ( N_S_c_353_n N_A0_c_918_n ) capacitor c=0.00308814f //x=3.135 \
 //y=1.915 //x2=4.07 //y2=2.08
cc_366 ( N_S_M9_noxref_g N_A0_M11_noxref_g ) capacitor c=0.0104611f //x=3.23 \
 //y=6.02 //x2=4.11 //y2=6.02
cc_367 ( N_S_M10_noxref_g N_A0_M11_noxref_g ) capacitor c=0.106811f //x=3.67 \
 //y=6.02 //x2=4.11 //y2=6.02
cc_368 ( N_S_M10_noxref_g N_A0_M12_noxref_g ) capacitor c=0.0100341f //x=3.67 \
 //y=6.02 //x2=4.55 //y2=6.02
cc_369 ( N_S_c_350_n N_A0_c_935_n ) capacitor c=4.86506e-19 //x=3.135 \
 //y=0.865 //x2=4.105 //y2=0.905
cc_370 ( N_S_c_352_n N_A0_c_935_n ) capacitor c=0.00152104f //x=3.135 //y=1.21 \
 //x2=4.105 //y2=0.905
cc_371 ( N_S_c_356_n N_A0_c_935_n ) capacitor c=0.0151475f //x=3.665 //y=0.865 \
 //x2=4.105 //y2=0.905
cc_372 ( N_S_c_433_p N_A0_c_938_n ) capacitor c=0.00109982f //x=3.135 //y=1.52 \
 //x2=4.105 //y2=1.25
cc_373 ( N_S_c_358_n N_A0_c_938_n ) capacitor c=0.0111064f //x=3.665 //y=1.21 \
 //x2=4.105 //y2=1.25
cc_374 ( N_S_c_433_p N_A0_c_940_n ) capacitor c=9.57794e-19 //x=3.135 //y=1.52 \
 //x2=4.105 //y2=1.56
cc_375 ( N_S_c_353_n N_A0_c_940_n ) capacitor c=0.00662747f //x=3.135 \
 //y=1.915 //x2=4.105 //y2=1.56
cc_376 ( N_S_c_358_n N_A0_c_940_n ) capacitor c=0.00862358f //x=3.665 //y=1.21 \
 //x2=4.105 //y2=1.56
cc_377 ( N_S_c_356_n N_A0_c_943_n ) capacitor c=0.00124821f //x=3.665 \
 //y=0.865 //x2=4.635 //y2=0.905
cc_378 ( N_S_c_358_n N_A0_c_944_n ) capacitor c=0.00200715f //x=3.665 //y=1.21 \
 //x2=4.635 //y2=1.25
cc_379 ( N_S_c_342_n N_A0_c_945_n ) capacitor c=0.00307062f //x=3.33 //y=2.08 \
 //x2=4.07 //y2=2.08
cc_380 ( N_S_c_353_n N_A0_c_945_n ) capacitor c=0.0179092f //x=3.135 //y=1.915 \
 //x2=4.07 //y2=2.08
cc_381 ( N_S_c_342_n N_A0_c_947_n ) capacitor c=0.00344981f //x=3.33 //y=2.08 \
 //x2=4.1 //y2=4.7
cc_382 ( N_S_c_384_n N_A0_c_947_n ) capacitor c=0.0293367f //x=3.33 //y=4.7 \
 //x2=4.1 //y2=4.7
cc_383 ( N_S_c_329_n N_noxref_8_c_986_n ) capacitor c=0.00321948f //x=3.215 \
 //y=2.96 //x2=2.915 //y2=1.495
cc_384 ( N_S_c_353_n N_noxref_8_c_986_n ) capacitor c=0.0034165f //x=3.135 \
 //y=1.915 //x2=2.915 //y2=1.495
cc_385 ( N_S_c_329_n N_noxref_8_c_987_n ) capacitor c=0.00765882f //x=3.215 \
 //y=2.96 //x2=3.8 //y2=1.58
cc_386 ( N_S_c_342_n N_noxref_8_c_987_n ) capacitor c=0.0115783f //x=3.33 \
 //y=2.08 //x2=3.8 //y2=1.58
cc_387 ( N_S_c_433_p N_noxref_8_c_987_n ) capacitor c=0.00703567f //x=3.135 \
 //y=1.52 //x2=3.8 //y2=1.58
cc_388 ( N_S_c_353_n N_noxref_8_c_987_n ) capacitor c=0.01939f //x=3.135 \
 //y=1.915 //x2=3.8 //y2=1.58
cc_389 ( N_S_c_355_n N_noxref_8_c_987_n ) capacitor c=0.00780629f //x=3.51 \
 //y=1.365 //x2=3.8 //y2=1.58
cc_390 ( N_S_c_358_n N_noxref_8_c_987_n ) capacitor c=0.00339872f //x=3.665 \
 //y=1.21 //x2=3.8 //y2=1.58
cc_391 ( N_S_c_353_n N_noxref_8_c_995_n ) capacitor c=6.71402e-19 //x=3.135 \
 //y=1.915 //x2=3.885 //y2=1.495
cc_392 ( N_S_c_350_n N_noxref_8_M1_noxref_s ) capacitor c=0.0326577f //x=3.135 \
 //y=0.865 //x2=2.78 //y2=0.365
cc_393 ( N_S_c_433_p N_noxref_8_M1_noxref_s ) capacitor c=3.48408e-19 \
 //x=3.135 //y=1.52 //x2=2.78 //y2=0.365
cc_394 ( N_S_c_356_n N_noxref_8_M1_noxref_s ) capacitor c=0.0120759f //x=3.665 \
 //y=0.865 //x2=2.78 //y2=0.365
cc_395 ( N_noxref_4_c_456_n N_noxref_5_c_595_n ) capacitor c=0.173506f \
 //x=6.545 //y=3.33 //x2=9.875 //y2=2.96
cc_396 ( N_noxref_4_c_462_n N_noxref_5_c_595_n ) capacitor c=0.0250048f \
 //x=6.66 //y=2.08 //x2=9.875 //y2=2.96
cc_397 ( N_noxref_4_c_467_n N_noxref_5_c_595_n ) capacitor c=0.0044801f \
 //x=6.465 //y=1.915 //x2=9.875 //y2=2.96
cc_398 ( N_noxref_4_c_456_n N_noxref_5_c_602_n ) capacitor c=0.0293964f \
 //x=6.545 //y=3.33 //x2=4.925 //y2=2.96
cc_399 ( N_noxref_4_c_462_n N_noxref_5_c_602_n ) capacitor c=5.96166e-19 \
 //x=6.66 //y=2.08 //x2=4.925 //y2=2.96
cc_400 ( N_noxref_4_c_456_n N_noxref_5_c_620_n ) capacitor c=0.0087538f \
 //x=6.545 //y=3.33 //x2=4.245 //y2=5.2
cc_401 ( N_noxref_4_c_456_n N_noxref_5_c_624_n ) capacitor c=0.00851197f \
 //x=6.545 //y=3.33 //x2=3.535 //y2=5.2
cc_402 ( N_noxref_4_c_456_n N_noxref_5_c_667_n ) capacitor c=0.00488601f \
 //x=6.545 //y=3.33 //x2=4.455 //y2=1.655
cc_403 ( N_noxref_4_c_456_n N_noxref_5_c_604_n ) capacitor c=0.0268499f \
 //x=6.545 //y=3.33 //x2=4.81 //y2=2.96
cc_404 ( N_noxref_4_c_462_n N_noxref_5_c_604_n ) capacitor c=0.0139161f \
 //x=6.66 //y=2.08 //x2=4.81 //y2=2.96
cc_405 ( N_noxref_4_c_456_n N_noxref_6_c_774_n ) capacitor c=0.0114735f \
 //x=6.545 //y=3.33 //x2=8.255 //y2=3.33
cc_406 ( N_noxref_4_M14_noxref_g N_noxref_6_c_776_n ) capacitor c=0.0195934f \
 //x=7 //y=6.02 //x2=7.575 //y2=5.2
cc_407 ( N_noxref_4_c_456_n N_noxref_6_c_780_n ) capacitor c=7.64123e-19 \
 //x=6.545 //y=3.33 //x2=6.865 //y2=5.2
cc_408 ( N_noxref_4_c_462_n N_noxref_6_c_780_n ) capacitor c=0.00560864f \
 //x=6.66 //y=2.08 //x2=6.865 //y2=5.2
cc_409 ( N_noxref_4_M13_noxref_g N_noxref_6_c_780_n ) capacitor c=0.0177326f \
 //x=6.56 //y=6.02 //x2=6.865 //y2=5.2
cc_410 ( N_noxref_4_c_501_n N_noxref_6_c_780_n ) capacitor c=0.00589848f \
 //x=6.66 //y=4.7 //x2=6.865 //y2=5.2
cc_411 ( N_noxref_4_c_462_n N_noxref_6_c_765_n ) capacitor c=0.0036353f \
 //x=6.66 //y=2.08 //x2=8.14 //y2=3.33
cc_412 ( N_noxref_4_M14_noxref_g N_noxref_6_M13_noxref_d ) capacitor \
 c=0.0173476f //x=7 //y=6.02 //x2=6.635 //y2=5.02
cc_413 ( N_noxref_4_c_456_n N_A0_c_927_n ) capacitor c=9.89359e-19 //x=6.545 \
 //y=3.33 //x2=4.07 //y2=4.535
cc_414 ( N_noxref_4_c_456_n N_A0_c_918_n ) capacitor c=0.0276573f //x=6.545 \
 //y=3.33 //x2=4.07 //y2=2.08
cc_415 ( N_noxref_4_c_461_n N_A0_c_918_n ) capacitor c=0.00116216f //x=1.48 \
 //y=3.33 //x2=4.07 //y2=2.08
cc_416 ( N_noxref_4_c_462_n N_A0_c_918_n ) capacitor c=0.00116216f //x=6.66 \
 //y=2.08 //x2=4.07 //y2=2.08
cc_417 ( N_noxref_4_c_456_n N_noxref_8_c_987_n ) capacitor c=0.00379932f \
 //x=6.545 //y=3.33 //x2=3.8 //y2=1.58
cc_418 ( N_noxref_4_c_456_n N_noxref_8_c_995_n ) capacitor c=0.00224213f \
 //x=6.545 //y=3.33 //x2=3.885 //y2=1.495
cc_419 ( N_noxref_4_c_456_n N_noxref_8_c_996_n ) capacitor c=5.79678e-19 \
 //x=6.545 //y=3.33 //x2=4.77 //y2=0.53
cc_420 ( N_noxref_4_c_462_n N_A1_c_1052_n ) capacitor c=0.00400249f //x=6.66 \
 //y=2.08 //x2=7.4 //y2=4.535
cc_421 ( N_noxref_4_c_501_n N_A1_c_1052_n ) capacitor c=0.00417994f //x=6.66 \
 //y=4.7 //x2=7.4 //y2=4.535
cc_422 ( N_noxref_4_c_456_n N_A1_c_1043_n ) capacitor c=0.00318578f //x=6.545 \
 //y=3.33 //x2=7.4 //y2=2.08
cc_423 ( N_noxref_4_c_462_n N_A1_c_1043_n ) capacitor c=0.0845408f //x=6.66 \
 //y=2.08 //x2=7.4 //y2=2.08
cc_424 ( N_noxref_4_c_467_n N_A1_c_1043_n ) capacitor c=0.00308814f //x=6.465 \
 //y=1.915 //x2=7.4 //y2=2.08
cc_425 ( N_noxref_4_M13_noxref_g N_A1_M15_noxref_g ) capacitor c=0.0104611f \
 //x=6.56 //y=6.02 //x2=7.44 //y2=6.02
cc_426 ( N_noxref_4_M14_noxref_g N_A1_M15_noxref_g ) capacitor c=0.106811f \
 //x=7 //y=6.02 //x2=7.44 //y2=6.02
cc_427 ( N_noxref_4_M14_noxref_g N_A1_M16_noxref_g ) capacitor c=0.0100341f \
 //x=7 //y=6.02 //x2=7.88 //y2=6.02
cc_428 ( N_noxref_4_c_463_n N_A1_c_1060_n ) capacitor c=4.86506e-19 //x=6.465 \
 //y=0.865 //x2=7.435 //y2=0.905
cc_429 ( N_noxref_4_c_465_n N_A1_c_1060_n ) capacitor c=0.00152104f //x=6.465 \
 //y=1.21 //x2=7.435 //y2=0.905
cc_430 ( N_noxref_4_c_470_n N_A1_c_1060_n ) capacitor c=0.0151475f //x=6.995 \
 //y=0.865 //x2=7.435 //y2=0.905
cc_431 ( N_noxref_4_c_466_n N_A1_c_1063_n ) capacitor c=0.00109982f //x=6.465 \
 //y=1.52 //x2=7.435 //y2=1.25
cc_432 ( N_noxref_4_c_472_n N_A1_c_1063_n ) capacitor c=0.0111064f //x=6.995 \
 //y=1.21 //x2=7.435 //y2=1.25
cc_433 ( N_noxref_4_c_466_n N_A1_c_1065_n ) capacitor c=9.57794e-19 //x=6.465 \
 //y=1.52 //x2=7.435 //y2=1.56
cc_434 ( N_noxref_4_c_467_n N_A1_c_1065_n ) capacitor c=0.00662747f //x=6.465 \
 //y=1.915 //x2=7.435 //y2=1.56
cc_435 ( N_noxref_4_c_472_n N_A1_c_1065_n ) capacitor c=0.00862358f //x=6.995 \
 //y=1.21 //x2=7.435 //y2=1.56
cc_436 ( N_noxref_4_c_470_n N_A1_c_1068_n ) capacitor c=0.00124821f //x=6.995 \
 //y=0.865 //x2=7.965 //y2=0.905
cc_437 ( N_noxref_4_c_472_n N_A1_c_1069_n ) capacitor c=0.00200715f //x=6.995 \
 //y=1.21 //x2=7.965 //y2=1.25
cc_438 ( N_noxref_4_c_462_n N_A1_c_1070_n ) capacitor c=0.00307062f //x=6.66 \
 //y=2.08 //x2=7.4 //y2=2.08
cc_439 ( N_noxref_4_c_467_n N_A1_c_1070_n ) capacitor c=0.0179092f //x=6.465 \
 //y=1.915 //x2=7.4 //y2=2.08
cc_440 ( N_noxref_4_c_462_n N_A1_c_1072_n ) capacitor c=0.00344981f //x=6.66 \
 //y=2.08 //x2=7.43 //y2=4.7
cc_441 ( N_noxref_4_c_501_n N_A1_c_1072_n ) capacitor c=0.0293367f //x=6.66 \
 //y=4.7 //x2=7.43 //y2=4.7
cc_442 ( N_noxref_4_c_467_n N_noxref_10_c_1134_n ) capacitor c=0.0034165f \
 //x=6.465 //y=1.915 //x2=6.245 //y2=1.495
cc_443 ( N_noxref_4_c_462_n N_noxref_10_c_1112_n ) capacitor c=0.0115894f \
 //x=6.66 //y=2.08 //x2=7.13 //y2=1.58
cc_444 ( N_noxref_4_c_466_n N_noxref_10_c_1112_n ) capacitor c=0.00703567f \
 //x=6.465 //y=1.52 //x2=7.13 //y2=1.58
cc_445 ( N_noxref_4_c_467_n N_noxref_10_c_1112_n ) capacitor c=0.01939f \
 //x=6.465 //y=1.915 //x2=7.13 //y2=1.58
cc_446 ( N_noxref_4_c_469_n N_noxref_10_c_1112_n ) capacitor c=0.00780629f \
 //x=6.84 //y=1.365 //x2=7.13 //y2=1.58
cc_447 ( N_noxref_4_c_472_n N_noxref_10_c_1112_n ) capacitor c=0.00339872f \
 //x=6.995 //y=1.21 //x2=7.13 //y2=1.58
cc_448 ( N_noxref_4_c_467_n N_noxref_10_c_1120_n ) capacitor c=6.71402e-19 \
 //x=6.465 //y=1.915 //x2=7.215 //y2=1.495
cc_449 ( N_noxref_4_c_463_n N_noxref_10_M3_noxref_s ) capacitor c=0.0326577f \
 //x=6.465 //y=0.865 //x2=6.11 //y2=0.365
cc_450 ( N_noxref_4_c_466_n N_noxref_10_M3_noxref_s ) capacitor c=3.48408e-19 \
 //x=6.465 //y=1.52 //x2=6.11 //y2=0.365
cc_451 ( N_noxref_4_c_470_n N_noxref_10_M3_noxref_s ) capacitor c=0.0120759f \
 //x=6.995 //y=0.865 //x2=6.11 //y2=0.365
cc_452 ( N_noxref_5_c_595_n N_noxref_6_c_763_n ) capacitor c=0.1737f //x=9.875 \
 //y=2.96 //x2=10.615 //y2=3.33
cc_453 ( N_noxref_5_c_605_n N_noxref_6_c_763_n ) capacitor c=0.0270785f \
 //x=9.99 //y=2.08 //x2=10.615 //y2=3.33
cc_454 ( N_noxref_5_c_595_n N_noxref_6_c_774_n ) capacitor c=0.0292689f \
 //x=9.875 //y=2.96 //x2=8.255 //y2=3.33
cc_455 ( N_noxref_5_c_605_n N_noxref_6_c_774_n ) capacitor c=3.78304e-19 \
 //x=9.99 //y=2.08 //x2=8.255 //y2=3.33
cc_456 ( N_noxref_5_c_595_n N_noxref_6_c_776_n ) capacitor c=0.00681665f \
 //x=9.875 //y=2.96 //x2=7.575 //y2=5.2
cc_457 ( N_noxref_5_c_595_n N_noxref_6_c_780_n ) capacitor c=0.0065469f \
 //x=9.875 //y=2.96 //x2=6.865 //y2=5.2
cc_458 ( N_noxref_5_c_595_n N_noxref_6_c_822_n ) capacitor c=0.00745069f \
 //x=9.875 //y=2.96 //x2=7.785 //y2=1.655
cc_459 ( N_noxref_5_c_595_n N_noxref_6_c_765_n ) capacitor c=0.026264f \
 //x=9.875 //y=2.96 //x2=8.14 //y2=3.33
cc_460 ( N_noxref_5_c_604_n N_noxref_6_c_765_n ) capacitor c=3.49822e-19 \
 //x=4.81 //y=2.96 //x2=8.14 //y2=3.33
cc_461 ( N_noxref_5_c_605_n N_noxref_6_c_765_n ) capacitor c=0.0139777f \
 //x=9.99 //y=2.08 //x2=8.14 //y2=3.33
cc_462 ( N_noxref_5_c_605_n N_noxref_6_c_826_n ) capacitor c=0.00400249f \
 //x=9.99 //y=2.08 //x2=10.73 //y2=4.535
cc_463 ( N_noxref_5_c_639_n N_noxref_6_c_826_n ) capacitor c=0.00417994f \
 //x=9.99 //y=4.7 //x2=10.73 //y2=4.535
cc_464 ( N_noxref_5_c_595_n N_noxref_6_c_766_n ) capacitor c=0.00735597f \
 //x=9.875 //y=2.96 //x2=10.73 //y2=2.08
cc_465 ( N_noxref_5_c_605_n N_noxref_6_c_766_n ) capacitor c=0.0840234f \
 //x=9.99 //y=2.08 //x2=10.73 //y2=2.08
cc_466 ( N_noxref_5_c_610_n N_noxref_6_c_766_n ) capacitor c=0.00308814f \
 //x=9.795 //y=1.915 //x2=10.73 //y2=2.08
cc_467 ( N_noxref_5_M17_noxref_g N_noxref_6_M19_noxref_g ) capacitor \
 c=0.0104611f //x=9.89 //y=6.02 //x2=10.77 //y2=6.02
cc_468 ( N_noxref_5_M18_noxref_g N_noxref_6_M19_noxref_g ) capacitor \
 c=0.106811f //x=10.33 //y=6.02 //x2=10.77 //y2=6.02
cc_469 ( N_noxref_5_M18_noxref_g N_noxref_6_M20_noxref_g ) capacitor \
 c=0.0100341f //x=10.33 //y=6.02 //x2=11.21 //y2=6.02
cc_470 ( N_noxref_5_c_606_n N_noxref_6_c_834_n ) capacitor c=4.86506e-19 \
 //x=9.795 //y=0.865 //x2=10.765 //y2=0.905
cc_471 ( N_noxref_5_c_608_n N_noxref_6_c_834_n ) capacitor c=0.00152104f \
 //x=9.795 //y=1.21 //x2=10.765 //y2=0.905
cc_472 ( N_noxref_5_c_613_n N_noxref_6_c_834_n ) capacitor c=0.0151475f \
 //x=10.325 //y=0.865 //x2=10.765 //y2=0.905
cc_473 ( N_noxref_5_c_609_n N_noxref_6_c_837_n ) capacitor c=0.00109982f \
 //x=9.795 //y=1.52 //x2=10.765 //y2=1.25
cc_474 ( N_noxref_5_c_615_n N_noxref_6_c_837_n ) capacitor c=0.0111064f \
 //x=10.325 //y=1.21 //x2=10.765 //y2=1.25
cc_475 ( N_noxref_5_c_609_n N_noxref_6_c_839_n ) capacitor c=9.57794e-19 \
 //x=9.795 //y=1.52 //x2=10.765 //y2=1.56
cc_476 ( N_noxref_5_c_610_n N_noxref_6_c_839_n ) capacitor c=0.00662747f \
 //x=9.795 //y=1.915 //x2=10.765 //y2=1.56
cc_477 ( N_noxref_5_c_615_n N_noxref_6_c_839_n ) capacitor c=0.00862358f \
 //x=10.325 //y=1.21 //x2=10.765 //y2=1.56
cc_478 ( N_noxref_5_c_613_n N_noxref_6_c_842_n ) capacitor c=0.00124821f \
 //x=10.325 //y=0.865 //x2=11.295 //y2=0.905
cc_479 ( N_noxref_5_c_615_n N_noxref_6_c_843_n ) capacitor c=0.00200715f \
 //x=10.325 //y=1.21 //x2=11.295 //y2=1.25
cc_480 ( N_noxref_5_c_605_n N_noxref_6_c_844_n ) capacitor c=0.00307062f \
 //x=9.99 //y=2.08 //x2=10.73 //y2=2.08
cc_481 ( N_noxref_5_c_610_n N_noxref_6_c_844_n ) capacitor c=0.0179092f \
 //x=9.795 //y=1.915 //x2=10.73 //y2=2.08
cc_482 ( N_noxref_5_c_605_n N_noxref_6_c_846_n ) capacitor c=0.00344981f \
 //x=9.99 //y=2.08 //x2=10.76 //y2=4.7
cc_483 ( N_noxref_5_c_639_n N_noxref_6_c_846_n ) capacitor c=0.0293367f \
 //x=9.99 //y=4.7 //x2=10.76 //y2=4.7
cc_484 ( N_noxref_5_c_620_n N_A0_c_927_n ) capacitor c=0.0131334f //x=4.245 \
 //y=5.2 //x2=4.07 //y2=4.535
cc_485 ( N_noxref_5_c_604_n N_A0_c_927_n ) capacitor c=0.0101284f //x=4.81 \
 //y=2.96 //x2=4.07 //y2=4.535
cc_486 ( N_noxref_5_c_602_n N_A0_c_918_n ) capacitor c=0.00318578f //x=4.925 \
 //y=2.96 //x2=4.07 //y2=2.08
cc_487 ( N_noxref_5_c_604_n N_A0_c_918_n ) capacitor c=0.0793882f //x=4.81 \
 //y=2.96 //x2=4.07 //y2=2.08
cc_488 ( N_noxref_5_c_620_n N_A0_M11_noxref_g ) capacitor c=0.0166421f \
 //x=4.245 //y=5.2 //x2=4.11 //y2=6.02
cc_489 ( N_noxref_5_M11_noxref_d N_A0_M11_noxref_g ) capacitor c=0.0173476f \
 //x=4.185 //y=5.02 //x2=4.11 //y2=6.02
cc_490 ( N_noxref_5_c_626_n N_A0_M12_noxref_g ) capacitor c=0.021201f \
 //x=4.725 //y=5.2 //x2=4.55 //y2=6.02
cc_491 ( N_noxref_5_M11_noxref_d N_A0_M12_noxref_g ) capacitor c=0.0179769f \
 //x=4.185 //y=5.02 //x2=4.55 //y2=6.02
cc_492 ( N_noxref_5_M2_noxref_d N_A0_c_935_n ) capacitor c=0.00217566f \
 //x=4.18 //y=0.905 //x2=4.105 //y2=0.905
cc_493 ( N_noxref_5_M2_noxref_d N_A0_c_938_n ) capacitor c=0.0034598f //x=4.18 \
 //y=0.905 //x2=4.105 //y2=1.25
cc_494 ( N_noxref_5_M2_noxref_d N_A0_c_940_n ) capacitor c=0.0065582f //x=4.18 \
 //y=0.905 //x2=4.105 //y2=1.56
cc_495 ( N_noxref_5_c_604_n N_A0_c_964_n ) capacitor c=0.0142673f //x=4.81 \
 //y=2.96 //x2=4.475 //y2=4.79
cc_496 ( N_noxref_5_c_714_p N_A0_c_964_n ) capacitor c=0.00421574f //x=4.33 \
 //y=5.2 //x2=4.475 //y2=4.79
cc_497 ( N_noxref_5_M2_noxref_d N_A0_c_966_n ) capacitor c=0.00241102f \
 //x=4.18 //y=0.905 //x2=4.48 //y2=0.75
cc_498 ( N_noxref_5_c_603_n N_A0_c_967_n ) capacitor c=0.00359704f //x=4.725 \
 //y=1.655 //x2=4.48 //y2=1.405
cc_499 ( N_noxref_5_M2_noxref_d N_A0_c_967_n ) capacitor c=0.0138845f //x=4.18 \
 //y=0.905 //x2=4.48 //y2=1.405
cc_500 ( N_noxref_5_M2_noxref_d N_A0_c_943_n ) capacitor c=0.00132245f \
 //x=4.18 //y=0.905 //x2=4.635 //y2=0.905
cc_501 ( N_noxref_5_c_603_n N_A0_c_944_n ) capacitor c=0.00457401f //x=4.725 \
 //y=1.655 //x2=4.635 //y2=1.25
cc_502 ( N_noxref_5_M2_noxref_d N_A0_c_944_n ) capacitor c=0.00566463f \
 //x=4.18 //y=0.905 //x2=4.635 //y2=1.25
cc_503 ( N_noxref_5_c_604_n N_A0_c_945_n ) capacitor c=0.00877984f //x=4.81 \
 //y=2.96 //x2=4.07 //y2=2.08
cc_504 ( N_noxref_5_c_604_n N_A0_c_973_n ) capacitor c=0.00306024f //x=4.81 \
 //y=2.96 //x2=4.07 //y2=1.915
cc_505 ( N_noxref_5_M2_noxref_d N_A0_c_973_n ) capacitor c=0.00660593f \
 //x=4.18 //y=0.905 //x2=4.07 //y2=1.915
cc_506 ( N_noxref_5_c_620_n N_A0_c_947_n ) capacitor c=0.00345427f //x=4.245 \
 //y=5.2 //x2=4.1 //y2=4.7
cc_507 ( N_noxref_5_c_604_n N_A0_c_947_n ) capacitor c=0.00533692f //x=4.81 \
 //y=2.96 //x2=4.1 //y2=4.7
cc_508 ( N_noxref_5_c_667_n N_noxref_8_c_986_n ) capacitor c=3.15806e-19 \
 //x=4.455 //y=1.655 //x2=2.915 //y2=1.495
cc_509 ( N_noxref_5_c_667_n N_noxref_8_c_995_n ) capacitor c=0.0201674f \
 //x=4.455 //y=1.655 //x2=3.885 //y2=1.495
cc_510 ( N_noxref_5_c_603_n N_noxref_8_c_996_n ) capacitor c=0.00465585f \
 //x=4.725 //y=1.655 //x2=4.77 //y2=0.53
cc_511 ( N_noxref_5_M2_noxref_d N_noxref_8_c_996_n ) capacitor c=0.0117692f \
 //x=4.18 //y=0.905 //x2=4.77 //y2=0.53
cc_512 ( N_noxref_5_c_595_n N_noxref_8_M1_noxref_s ) capacitor c=2.01804e-19 \
 //x=9.875 //y=2.96 //x2=2.78 //y2=0.365
cc_513 ( N_noxref_5_c_602_n N_noxref_8_M1_noxref_s ) capacitor c=4.48477e-19 \
 //x=4.925 //y=2.96 //x2=2.78 //y2=0.365
cc_514 ( N_noxref_5_c_603_n N_noxref_8_M1_noxref_s ) capacitor c=0.0140125f \
 //x=4.725 //y=1.655 //x2=2.78 //y2=0.365
cc_515 ( N_noxref_5_M2_noxref_d N_noxref_8_M1_noxref_s ) capacitor \
 c=0.0437911f //x=4.18 //y=0.905 //x2=2.78 //y2=0.365
cc_516 ( N_noxref_5_c_595_n N_A1_c_1052_n ) capacitor c=8.80769e-19 //x=9.875 \
 //y=2.96 //x2=7.4 //y2=4.535
cc_517 ( N_noxref_5_c_595_n N_A1_c_1043_n ) capacitor c=0.0270593f //x=9.875 \
 //y=2.96 //x2=7.4 //y2=2.08
cc_518 ( N_noxref_5_c_604_n N_A1_c_1043_n ) capacitor c=0.00116216f //x=4.81 \
 //y=2.96 //x2=7.4 //y2=2.08
cc_519 ( N_noxref_5_c_605_n N_A1_c_1043_n ) capacitor c=0.00116216f //x=9.99 \
 //y=2.08 //x2=7.4 //y2=2.08
cc_520 ( N_noxref_5_c_595_n N_A1_c_1070_n ) capacitor c=0.00172252f //x=9.875 \
 //y=2.96 //x2=7.4 //y2=2.08
cc_521 ( N_noxref_5_c_595_n N_noxref_10_c_1134_n ) capacitor c=0.00321948f \
 //x=9.875 //y=2.96 //x2=6.245 //y2=1.495
cc_522 ( N_noxref_5_c_603_n N_noxref_10_c_1134_n ) capacitor c=3.22188e-19 \
 //x=4.725 //y=1.655 //x2=6.245 //y2=1.495
cc_523 ( N_noxref_5_c_595_n N_noxref_10_c_1112_n ) capacitor c=0.0126309f \
 //x=9.875 //y=2.96 //x2=7.13 //y2=1.58
cc_524 ( N_noxref_5_c_595_n N_noxref_10_c_1120_n ) capacitor c=0.00307759f \
 //x=9.875 //y=2.96 //x2=7.215 //y2=1.495
cc_525 ( N_noxref_5_c_595_n N_noxref_10_c_1121_n ) capacitor c=7.29507e-19 \
 //x=9.875 //y=2.96 //x2=8.1 //y2=0.53
cc_526 ( N_noxref_5_c_595_n N_noxref_10_M3_noxref_s ) capacitor c=6.20367e-19 \
 //x=9.875 //y=2.96 //x2=6.11 //y2=0.365
cc_527 ( N_noxref_5_c_605_n Y ) capacitor c=0.00425321f //x=9.99 //y=2.08 \
 //x2=11.47 //y2=2.22
cc_528 ( N_noxref_5_M18_noxref_g N_Y_c_1174_n ) capacitor c=0.0192312f \
 //x=10.33 //y=6.02 //x2=10.905 //y2=5.2
cc_529 ( N_noxref_5_c_605_n N_Y_c_1178_n ) capacitor c=0.0056116f //x=9.99 \
 //y=2.08 //x2=10.195 //y2=5.2
cc_530 ( N_noxref_5_M17_noxref_g N_Y_c_1178_n ) capacitor c=0.0177326f \
 //x=9.89 //y=6.02 //x2=10.195 //y2=5.2
cc_531 ( N_noxref_5_c_639_n N_Y_c_1178_n ) capacitor c=0.00589848f //x=9.99 \
 //y=4.7 //x2=10.195 //y2=5.2
cc_532 ( N_noxref_5_M18_noxref_g N_Y_M17_noxref_d ) capacitor c=0.0173476f \
 //x=10.33 //y=6.02 //x2=9.965 //y2=5.02
cc_533 ( N_noxref_5_c_595_n N_noxref_12_c_1249_n ) capacitor c=0.00321948f \
 //x=9.875 //y=2.96 //x2=9.575 //y2=1.495
cc_534 ( N_noxref_5_c_610_n N_noxref_12_c_1249_n ) capacitor c=0.0034165f \
 //x=9.795 //y=1.915 //x2=9.575 //y2=1.495
cc_535 ( N_noxref_5_c_595_n N_noxref_12_c_1232_n ) capacitor c=0.00765882f \
 //x=9.875 //y=2.96 //x2=10.46 //y2=1.58
cc_536 ( N_noxref_5_c_605_n N_noxref_12_c_1232_n ) capacitor c=0.0115783f \
 //x=9.99 //y=2.08 //x2=10.46 //y2=1.58
cc_537 ( N_noxref_5_c_609_n N_noxref_12_c_1232_n ) capacitor c=0.00703567f \
 //x=9.795 //y=1.52 //x2=10.46 //y2=1.58
cc_538 ( N_noxref_5_c_610_n N_noxref_12_c_1232_n ) capacitor c=0.01939f \
 //x=9.795 //y=1.915 //x2=10.46 //y2=1.58
cc_539 ( N_noxref_5_c_612_n N_noxref_12_c_1232_n ) capacitor c=0.00780629f \
 //x=10.17 //y=1.365 //x2=10.46 //y2=1.58
cc_540 ( N_noxref_5_c_615_n N_noxref_12_c_1232_n ) capacitor c=0.00339872f \
 //x=10.325 //y=1.21 //x2=10.46 //y2=1.58
cc_541 ( N_noxref_5_c_610_n N_noxref_12_c_1239_n ) capacitor c=6.71402e-19 \
 //x=9.795 //y=1.915 //x2=10.545 //y2=1.495
cc_542 ( N_noxref_5_c_606_n N_noxref_12_M5_noxref_s ) capacitor c=0.0326577f \
 //x=9.795 //y=0.865 //x2=9.44 //y2=0.365
cc_543 ( N_noxref_5_c_609_n N_noxref_12_M5_noxref_s ) capacitor c=3.48408e-19 \
 //x=9.795 //y=1.52 //x2=9.44 //y2=0.365
cc_544 ( N_noxref_5_c_613_n N_noxref_12_M5_noxref_s ) capacitor c=0.0120759f \
 //x=10.325 //y=0.865 //x2=9.44 //y2=0.365
cc_545 ( N_noxref_6_c_776_n N_A1_c_1052_n ) capacitor c=0.0131536f //x=7.575 \
 //y=5.2 //x2=7.4 //y2=4.535
cc_546 ( N_noxref_6_c_765_n N_A1_c_1052_n ) capacitor c=0.0101284f //x=8.14 \
 //y=3.33 //x2=7.4 //y2=4.535
cc_547 ( N_noxref_6_c_774_n N_A1_c_1043_n ) capacitor c=0.00317669f //x=8.255 \
 //y=3.33 //x2=7.4 //y2=2.08
cc_548 ( N_noxref_6_c_765_n N_A1_c_1043_n ) capacitor c=0.0793882f //x=8.14 \
 //y=3.33 //x2=7.4 //y2=2.08
cc_549 ( N_noxref_6_c_776_n N_A1_M15_noxref_g ) capacitor c=0.0166421f \
 //x=7.575 //y=5.2 //x2=7.44 //y2=6.02
cc_550 ( N_noxref_6_M15_noxref_d N_A1_M15_noxref_g ) capacitor c=0.0173476f \
 //x=7.515 //y=5.02 //x2=7.44 //y2=6.02
cc_551 ( N_noxref_6_c_782_n N_A1_M16_noxref_g ) capacitor c=0.0215633f \
 //x=8.055 //y=5.2 //x2=7.88 //y2=6.02
cc_552 ( N_noxref_6_M15_noxref_d N_A1_M16_noxref_g ) capacitor c=0.0179769f \
 //x=7.515 //y=5.02 //x2=7.88 //y2=6.02
cc_553 ( N_noxref_6_M4_noxref_d N_A1_c_1060_n ) capacitor c=0.00217566f \
 //x=7.51 //y=0.905 //x2=7.435 //y2=0.905
cc_554 ( N_noxref_6_M4_noxref_d N_A1_c_1063_n ) capacitor c=0.0034598f \
 //x=7.51 //y=0.905 //x2=7.435 //y2=1.25
cc_555 ( N_noxref_6_M4_noxref_d N_A1_c_1065_n ) capacitor c=0.0065582f \
 //x=7.51 //y=0.905 //x2=7.435 //y2=1.56
cc_556 ( N_noxref_6_c_765_n N_A1_c_1090_n ) capacitor c=0.0142673f //x=8.14 \
 //y=3.33 //x2=7.805 //y2=4.79
cc_557 ( N_noxref_6_c_860_p N_A1_c_1090_n ) capacitor c=0.00421574f //x=7.66 \
 //y=5.2 //x2=7.805 //y2=4.79
cc_558 ( N_noxref_6_M4_noxref_d N_A1_c_1092_n ) capacitor c=0.00241102f \
 //x=7.51 //y=0.905 //x2=7.81 //y2=0.75
cc_559 ( N_noxref_6_c_764_n N_A1_c_1093_n ) capacitor c=0.00359704f //x=8.055 \
 //y=1.655 //x2=7.81 //y2=1.405
cc_560 ( N_noxref_6_M4_noxref_d N_A1_c_1093_n ) capacitor c=0.0138845f \
 //x=7.51 //y=0.905 //x2=7.81 //y2=1.405
cc_561 ( N_noxref_6_M4_noxref_d N_A1_c_1068_n ) capacitor c=0.00132245f \
 //x=7.51 //y=0.905 //x2=7.965 //y2=0.905
cc_562 ( N_noxref_6_c_764_n N_A1_c_1069_n ) capacitor c=0.00457401f //x=8.055 \
 //y=1.655 //x2=7.965 //y2=1.25
cc_563 ( N_noxref_6_M4_noxref_d N_A1_c_1069_n ) capacitor c=0.00566463f \
 //x=7.51 //y=0.905 //x2=7.965 //y2=1.25
cc_564 ( N_noxref_6_c_765_n N_A1_c_1070_n ) capacitor c=0.00877984f //x=8.14 \
 //y=3.33 //x2=7.4 //y2=2.08
cc_565 ( N_noxref_6_c_765_n N_A1_c_1099_n ) capacitor c=0.00306024f //x=8.14 \
 //y=3.33 //x2=7.4 //y2=1.915
cc_566 ( N_noxref_6_M4_noxref_d N_A1_c_1099_n ) capacitor c=0.00660593f \
 //x=7.51 //y=0.905 //x2=7.4 //y2=1.915
cc_567 ( N_noxref_6_c_776_n N_A1_c_1072_n ) capacitor c=0.00345427f //x=7.575 \
 //y=5.2 //x2=7.43 //y2=4.7
cc_568 ( N_noxref_6_c_765_n N_A1_c_1072_n ) capacitor c=0.00533692f //x=8.14 \
 //y=3.33 //x2=7.43 //y2=4.7
cc_569 ( N_noxref_6_c_822_n N_noxref_10_c_1134_n ) capacitor c=3.15806e-19 \
 //x=7.785 //y=1.655 //x2=6.245 //y2=1.495
cc_570 ( N_noxref_6_c_822_n N_noxref_10_c_1120_n ) capacitor c=0.0203424f \
 //x=7.785 //y=1.655 //x2=7.215 //y2=1.495
cc_571 ( N_noxref_6_c_764_n N_noxref_10_c_1121_n ) capacitor c=0.00464204f \
 //x=8.055 //y=1.655 //x2=8.1 //y2=0.53
cc_572 ( N_noxref_6_M4_noxref_d N_noxref_10_c_1121_n ) capacitor c=0.0117318f \
 //x=7.51 //y=0.905 //x2=8.1 //y2=0.53
cc_573 ( N_noxref_6_c_764_n N_noxref_10_M3_noxref_s ) capacitor c=0.0140283f \
 //x=8.055 //y=1.655 //x2=6.11 //y2=0.365
cc_574 ( N_noxref_6_M4_noxref_d N_noxref_10_M3_noxref_s ) capacitor \
 c=0.043966f //x=7.51 //y=0.905 //x2=6.11 //y2=0.365
cc_575 ( N_noxref_6_c_763_n Y ) capacitor c=0.00549673f //x=10.615 //y=3.33 \
 //x2=11.47 //y2=2.22
cc_576 ( N_noxref_6_c_765_n Y ) capacitor c=3.49822e-19 //x=8.14 //y=3.33 \
 //x2=11.47 //y2=2.22
cc_577 ( N_noxref_6_c_826_n Y ) capacitor c=0.0101115f //x=10.73 //y=4.535 \
 //x2=11.47 //y2=2.22
cc_578 ( N_noxref_6_c_766_n Y ) capacitor c=0.0813921f //x=10.73 //y=2.08 \
 //x2=11.47 //y2=2.22
cc_579 ( N_noxref_6_c_882_p Y ) capacitor c=0.0142673f //x=11.135 //y=4.79 \
 //x2=11.47 //y2=2.22
cc_580 ( N_noxref_6_c_844_n Y ) capacitor c=0.00877984f //x=10.73 //y=2.08 \
 //x2=11.47 //y2=2.22
cc_581 ( N_noxref_6_c_884_p Y ) capacitor c=0.00306024f //x=10.73 //y=1.915 \
 //x2=11.47 //y2=2.22
cc_582 ( N_noxref_6_c_846_n Y ) capacitor c=0.00533692f //x=10.76 //y=4.7 \
 //x2=11.47 //y2=2.22
cc_583 ( N_noxref_6_c_763_n N_Y_c_1174_n ) capacitor c=0.00113909f //x=10.615 \
 //y=3.33 //x2=10.905 //y2=5.2
cc_584 ( N_noxref_6_c_826_n N_Y_c_1174_n ) capacitor c=0.0131311f //x=10.73 \
 //y=4.535 //x2=10.905 //y2=5.2
cc_585 ( N_noxref_6_M19_noxref_g N_Y_c_1174_n ) capacitor c=0.0166421f \
 //x=10.77 //y=6.02 //x2=10.905 //y2=5.2
cc_586 ( N_noxref_6_c_846_n N_Y_c_1174_n ) capacitor c=0.00345427f //x=10.76 \
 //y=4.7 //x2=10.905 //y2=5.2
cc_587 ( N_noxref_6_c_763_n N_Y_c_1178_n ) capacitor c=0.008207f //x=10.615 \
 //y=3.33 //x2=10.195 //y2=5.2
cc_588 ( N_noxref_6_M20_noxref_g N_Y_c_1180_n ) capacitor c=0.0223536f \
 //x=11.21 //y=6.02 //x2=11.385 //y2=5.2
cc_589 ( N_noxref_6_c_892_p N_Y_c_1168_n ) capacitor c=0.00359704f //x=11.14 \
 //y=1.405 //x2=11.385 //y2=1.655
cc_590 ( N_noxref_6_c_843_n N_Y_c_1168_n ) capacitor c=0.00457401f //x=11.295 \
 //y=1.25 //x2=11.385 //y2=1.655
cc_591 ( N_noxref_6_c_882_p N_Y_c_1215_n ) capacitor c=0.00414324f //x=11.135 \
 //y=4.79 //x2=10.99 //y2=5.2
cc_592 ( N_noxref_6_c_834_n N_Y_M6_noxref_d ) capacitor c=0.00217566f \
 //x=10.765 //y=0.905 //x2=10.84 //y2=0.905
cc_593 ( N_noxref_6_c_837_n N_Y_M6_noxref_d ) capacitor c=0.0034598f \
 //x=10.765 //y=1.25 //x2=10.84 //y2=0.905
cc_594 ( N_noxref_6_c_839_n N_Y_M6_noxref_d ) capacitor c=0.0065582f \
 //x=10.765 //y=1.56 //x2=10.84 //y2=0.905
cc_595 ( N_noxref_6_c_898_p N_Y_M6_noxref_d ) capacitor c=0.00241102f \
 //x=11.14 //y=0.75 //x2=10.84 //y2=0.905
cc_596 ( N_noxref_6_c_892_p N_Y_M6_noxref_d ) capacitor c=0.0138845f //x=11.14 \
 //y=1.405 //x2=10.84 //y2=0.905
cc_597 ( N_noxref_6_c_842_n N_Y_M6_noxref_d ) capacitor c=0.00132245f \
 //x=11.295 //y=0.905 //x2=10.84 //y2=0.905
cc_598 ( N_noxref_6_c_843_n N_Y_M6_noxref_d ) capacitor c=0.00566463f \
 //x=11.295 //y=1.25 //x2=10.84 //y2=0.905
cc_599 ( N_noxref_6_c_884_p N_Y_M6_noxref_d ) capacitor c=0.00660593f \
 //x=10.73 //y=1.915 //x2=10.84 //y2=0.905
cc_600 ( N_noxref_6_M19_noxref_g N_Y_M19_noxref_d ) capacitor c=0.0173476f \
 //x=10.77 //y=6.02 //x2=10.845 //y2=5.02
cc_601 ( N_noxref_6_M20_noxref_g N_Y_M19_noxref_d ) capacitor c=0.0179769f \
 //x=11.21 //y=6.02 //x2=10.845 //y2=5.02
cc_602 ( N_noxref_6_c_764_n N_noxref_12_c_1249_n ) capacitor c=3.22188e-19 \
 //x=8.055 //y=1.655 //x2=9.575 //y2=1.495
cc_603 ( N_noxref_6_c_763_n N_noxref_12_c_1232_n ) capacitor c=0.00379932f \
 //x=10.615 //y=3.33 //x2=10.46 //y2=1.58
cc_604 ( N_noxref_6_c_763_n N_noxref_12_c_1239_n ) capacitor c=0.0022567f \
 //x=10.615 //y=3.33 //x2=10.545 //y2=1.495
cc_605 ( N_noxref_6_c_839_n N_noxref_12_c_1239_n ) capacitor c=0.00623646f \
 //x=10.765 //y=1.56 //x2=10.545 //y2=1.495
cc_606 ( N_noxref_6_c_844_n N_noxref_12_c_1239_n ) capacitor c=0.00176439f \
 //x=10.73 //y=2.08 //x2=10.545 //y2=1.495
cc_607 ( N_noxref_6_c_763_n N_noxref_12_c_1240_n ) capacitor c=2.75166e-19 \
 //x=10.615 //y=3.33 //x2=11.43 //y2=0.53
cc_608 ( N_noxref_6_c_766_n N_noxref_12_c_1240_n ) capacitor c=0.00159853f \
 //x=10.73 //y=2.08 //x2=11.43 //y2=0.53
cc_609 ( N_noxref_6_c_834_n N_noxref_12_c_1240_n ) capacitor c=0.018734f \
 //x=10.765 //y=0.905 //x2=11.43 //y2=0.53
cc_610 ( N_noxref_6_c_842_n N_noxref_12_c_1240_n ) capacitor c=0.00656458f \
 //x=11.295 //y=0.905 //x2=11.43 //y2=0.53
cc_611 ( N_noxref_6_c_844_n N_noxref_12_c_1240_n ) capacitor c=2.1838e-19 \
 //x=10.73 //y=2.08 //x2=11.43 //y2=0.53
cc_612 ( N_noxref_6_c_834_n N_noxref_12_M5_noxref_s ) capacitor c=0.00623646f \
 //x=10.765 //y=0.905 //x2=9.44 //y2=0.365
cc_613 ( N_noxref_6_c_842_n N_noxref_12_M5_noxref_s ) capacitor c=0.0143002f \
 //x=11.295 //y=0.905 //x2=9.44 //y2=0.365
cc_614 ( N_noxref_6_c_843_n N_noxref_12_M5_noxref_s ) capacitor c=0.00290153f \
 //x=11.295 //y=1.25 //x2=9.44 //y2=0.365
cc_615 ( N_A0_c_940_n N_noxref_8_c_995_n ) capacitor c=0.00623646f //x=4.105 \
 //y=1.56 //x2=3.885 //y2=1.495
cc_616 ( N_A0_c_945_n N_noxref_8_c_995_n ) capacitor c=0.00176439f //x=4.07 \
 //y=2.08 //x2=3.885 //y2=1.495
cc_617 ( N_A0_c_918_n N_noxref_8_c_996_n ) capacitor c=0.00159897f //x=4.07 \
 //y=2.08 //x2=4.77 //y2=0.53
cc_618 ( N_A0_c_935_n N_noxref_8_c_996_n ) capacitor c=0.0188655f //x=4.105 \
 //y=0.905 //x2=4.77 //y2=0.53
cc_619 ( N_A0_c_943_n N_noxref_8_c_996_n ) capacitor c=0.00656458f //x=4.635 \
 //y=0.905 //x2=4.77 //y2=0.53
cc_620 ( N_A0_c_945_n N_noxref_8_c_996_n ) capacitor c=2.1838e-19 //x=4.07 \
 //y=2.08 //x2=4.77 //y2=0.53
cc_621 ( N_A0_c_935_n N_noxref_8_M1_noxref_s ) capacitor c=0.00623646f \
 //x=4.105 //y=0.905 //x2=2.78 //y2=0.365
cc_622 ( N_A0_c_943_n N_noxref_8_M1_noxref_s ) capacitor c=0.0143002f \
 //x=4.635 //y=0.905 //x2=2.78 //y2=0.365
cc_623 ( N_A0_c_944_n N_noxref_8_M1_noxref_s ) capacitor c=0.00290153f \
 //x=4.635 //y=1.25 //x2=2.78 //y2=0.365
cc_624 ( N_noxref_8_c_999_n N_noxref_10_M3_noxref_s ) capacitor c=0.00174327f \
 //x=4.855 //y=0.615 //x2=6.11 //y2=0.365
cc_625 ( N_A1_c_1065_n N_noxref_10_c_1120_n ) capacitor c=0.00623646f \
 //x=7.435 //y=1.56 //x2=7.215 //y2=1.495
cc_626 ( N_A1_c_1070_n N_noxref_10_c_1120_n ) capacitor c=0.00174428f //x=7.4 \
 //y=2.08 //x2=7.215 //y2=1.495
cc_627 ( N_A1_c_1043_n N_noxref_10_c_1121_n ) capacitor c=0.00159235f //x=7.4 \
 //y=2.08 //x2=8.1 //y2=0.53
cc_628 ( N_A1_c_1060_n N_noxref_10_c_1121_n ) capacitor c=0.0188655f //x=7.435 \
 //y=0.905 //x2=8.1 //y2=0.53
cc_629 ( N_A1_c_1068_n N_noxref_10_c_1121_n ) capacitor c=0.00656458f \
 //x=7.965 //y=0.905 //x2=8.1 //y2=0.53
cc_630 ( N_A1_c_1070_n N_noxref_10_c_1121_n ) capacitor c=2.1838e-19 //x=7.4 \
 //y=2.08 //x2=8.1 //y2=0.53
cc_631 ( N_A1_c_1060_n N_noxref_10_M3_noxref_s ) capacitor c=0.00623646f \
 //x=7.435 //y=0.905 //x2=6.11 //y2=0.365
cc_632 ( N_A1_c_1068_n N_noxref_10_M3_noxref_s ) capacitor c=0.0143002f \
 //x=7.965 //y=0.905 //x2=6.11 //y2=0.365
cc_633 ( N_A1_c_1069_n N_noxref_10_M3_noxref_s ) capacitor c=0.00290153f \
 //x=7.965 //y=1.25 //x2=6.11 //y2=0.365
cc_634 ( N_noxref_10_c_1124_n N_noxref_12_M5_noxref_s ) capacitor \
 c=0.00174327f //x=8.185 //y=0.615 //x2=9.44 //y2=0.365
cc_635 ( N_Y_c_1226_p N_noxref_12_c_1249_n ) capacitor c=3.15806e-19 \
 //x=11.115 //y=1.655 //x2=9.575 //y2=1.495
cc_636 ( N_Y_c_1226_p N_noxref_12_c_1239_n ) capacitor c=0.0203424f //x=11.115 \
 //y=1.655 //x2=10.545 //y2=1.495
cc_637 ( N_Y_c_1168_n N_noxref_12_c_1240_n ) capacitor c=0.00469114f \
 //x=11.385 //y=1.655 //x2=11.43 //y2=0.53
cc_638 ( N_Y_M6_noxref_d N_noxref_12_c_1240_n ) capacitor c=0.0118355f \
 //x=10.84 //y=0.905 //x2=11.43 //y2=0.53
cc_639 ( N_Y_c_1168_n N_noxref_12_M5_noxref_s ) capacitor c=0.0144625f \
 //x=11.385 //y=1.655 //x2=9.44 //y2=0.365
cc_640 ( N_Y_M6_noxref_d N_noxref_12_M5_noxref_s ) capacitor c=0.043966f \
 //x=10.84 //y=0.905 //x2=9.44 //y2=0.365
