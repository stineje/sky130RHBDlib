* SPICE3 file created from AO3X1.ext - technology: sky130A

.subckt AO3X1 Y A B C VDD GND
X0 Y ao3x1_pcell_0/m1_1201_501# GND GND nshort w=3 l=0.15
X1 VDD ao3x1_pcell_0/m1_1201_501# Y VDD pshort w=2 l=0.15
X2 GND A ao3x1_pcell_0/aoi3x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X3 ao3x1_pcell_0/aoi3x1_pcell_0/m1_537_501# B ao3x1_pcell_0/aoi3x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X4 VDD A ao3x1_pcell_0/aoi3x1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X5 VDD B ao3x1_pcell_0/aoi3x1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X6 VDD ao3x1_pcell_0/aoi3x1_pcell_0/m1_537_501# ao3x1_pcell_0/aoi3x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X7 ao3x1_pcell_0/m1_1201_501# C ao3x1_pcell_0/aoi3x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X8 ao3x1_pcell_0/m1_1201_501# ao3x1_pcell_0/aoi3x1_pcell_0/m1_537_501# GND GND nshort w=3 l=0.15
X9 ao3x1_pcell_0/m1_1201_501# C GND GND nshort w=3 l=0.15
C0 VDD GND 3.35fF
.ends
