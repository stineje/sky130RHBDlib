* SPICE3 file created from XOR2X1.ext - technology: sky130A

.subckt XOR2X1 Y A B VDD GND
X0 Y a_807_943 a_575_1004 VDD pshort w=2 l=0.15 M=2
X1 a_1241_1004 a_185_182 Y VDD pshort w=2 l=0.15 M=2
X2 GND A a_556_74 GND nshort w=3 l=0.15
X3 VDD B a_807_943 VDD pshort w=2 l=0.15 M=2
X4 a_185_182 A GND GND nshort w=3 l=0.15
X5 VDD A a_575_1004 VDD pshort w=2 l=0.15 M=2
X6 Y a_185_182 a_1222_74 GND nshort w=3 l=0.15
X7 VDD A a_185_182 VDD pshort w=2 l=0.15 M=2
X8 a_807_943 B GND GND nshort w=3 l=0.15
X9 VDD B a_1241_1004 VDD pshort w=2 l=0.15 M=2
X10 Y B a_556_74 GND nshort w=3 l=0.15
X11 GND a_807_943 a_1222_74 GND nshort w=3 l=0.15
C0 B a_807_943 2.23fF
C1 VDD GND 5.63fF
.ends
