// File: AND2X1.spi.AND2X1.pxi
// Created: Tue Oct 15 15:44:19 2024
// 
simulator lang=spectre
x_PM_AND2X1\%GND ( GND N_GND_c_4_p N_GND_c_34_p N_GND_c_2_p N_GND_c_5_p \
 N_GND_c_6_p N_GND_c_60_p N_GND_c_7_p N_GND_c_23_p N_GND_c_1_p N_GND_c_3_p \
 N_GND_M0_noxref_d N_GND_M2_noxref_s )  PM_AND2X1\%GND
x_PM_AND2X1\%VDD ( VDD N_VDD_c_82_p N_VDD_c_88_p N_VDD_c_89_p N_VDD_c_102_p \
 N_VDD_c_79_n N_VDD_c_80_n N_VDD_c_81_n N_VDD_M3_noxref_s N_VDD_M4_noxref_d \
 N_VDD_M6_noxref_d N_VDD_M7_noxref_s N_VDD_M8_noxref_d )  PM_AND2X1\%VDD
x_PM_AND2X1\%noxref_3 ( N_noxref_3_c_149_n N_noxref_3_c_155_n \
 N_noxref_3_c_183_n N_noxref_3_c_187_n N_noxref_3_c_189_n N_noxref_3_c_156_n \
 N_noxref_3_c_250_p N_noxref_3_c_158_n N_noxref_3_c_159_n N_noxref_3_c_238_p \
 N_noxref_3_M2_noxref_g N_noxref_3_M7_noxref_g N_noxref_3_M8_noxref_g \
 N_noxref_3_c_164_n N_noxref_3_c_269_p N_noxref_3_c_270_p N_noxref_3_c_166_n \
 N_noxref_3_c_203_n N_noxref_3_c_204_n N_noxref_3_c_167_n N_noxref_3_c_261_p \
 N_noxref_3_c_168_n N_noxref_3_c_170_n N_noxref_3_c_171_n \
 N_noxref_3_M1_noxref_d N_noxref_3_M3_noxref_d N_noxref_3_M5_noxref_d )  \
 PM_AND2X1\%noxref_3
x_PM_AND2X1\%A ( A A A A A A A N_A_c_281_n N_A_M0_noxref_g N_A_M3_noxref_g \
 N_A_M4_noxref_g N_A_c_282_n N_A_c_284_n N_A_c_285_n N_A_c_286_n N_A_c_287_n \
 N_A_c_288_n N_A_c_289_n N_A_c_291_n N_A_c_299_n )  PM_AND2X1\%A
x_PM_AND2X1\%B ( B B B B B B B N_B_c_346_n N_B_c_337_n N_B_M1_noxref_g \
 N_B_M5_noxref_g N_B_M6_noxref_g N_B_c_355_n N_B_c_356_n N_B_c_357_n \
 N_B_c_358_n N_B_c_360_n N_B_c_361_n N_B_c_363_n N_B_c_364_n N_B_c_366_n \
 N_B_c_367_n N_B_c_369_n )  PM_AND2X1\%B
x_PM_AND2X1\%noxref_6 ( N_noxref_6_c_425_n N_noxref_6_c_401_n \
 N_noxref_6_c_405_n N_noxref_6_c_409_n N_noxref_6_c_410_n N_noxref_6_c_413_n \
 N_noxref_6_M0_noxref_s )  PM_AND2X1\%noxref_6
x_PM_AND2X1\%Y ( Y Y Y Y Y Y Y N_Y_c_452_n N_Y_c_476_n N_Y_c_462_n N_Y_c_465_n \
 N_Y_M2_noxref_d N_Y_M7_noxref_d )  PM_AND2X1\%Y
cc_1 ( N_GND_c_1_p N_VDD_c_79_n ) capacitor c=0.00989031f //x=5.18 //y=0 \
 //x2=5.18 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_80_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_81_n ) capacitor c=0.00855708f //x=3.33 //y=0 \
 //x2=3.33 //y2=7.4
cc_4 ( N_GND_c_4_p N_noxref_3_c_149_n ) capacitor c=0.011611f //x=5.18 //y=0 \
 //x2=3.955 //y2=3.33
cc_5 ( N_GND_c_5_p N_noxref_3_c_149_n ) capacitor c=0.00157139f //x=3.16 //y=0 \
 //x2=3.955 //y2=3.33
cc_6 ( N_GND_c_6_p N_noxref_3_c_149_n ) capacitor c=0.00110325f //x=3.875 \
 //y=0 //x2=3.955 //y2=3.33
cc_7 ( N_GND_c_7_p N_noxref_3_c_149_n ) capacitor c=2.76195e-19 //x=4.36 \
 //y=0.535 //x2=3.955 //y2=3.33
cc_8 ( N_GND_c_3_p N_noxref_3_c_149_n ) capacitor c=0.00820844f //x=3.33 //y=0 \
 //x2=3.955 //y2=3.33
cc_9 ( N_GND_M2_noxref_s N_noxref_3_c_149_n ) capacitor c=0.00164577f \
 //x=3.825 //y=0.37 //x2=3.955 //y2=3.33
cc_10 ( N_GND_c_4_p N_noxref_3_c_155_n ) capacitor c=0.00174211f //x=5.18 \
 //y=0 //x2=2.705 //y2=3.33
cc_11 ( N_GND_c_3_p N_noxref_3_c_156_n ) capacitor c=0.0461206f //x=3.33 //y=0 \
 //x2=2.505 //y2=1.655
cc_12 ( N_GND_M2_noxref_s N_noxref_3_c_156_n ) capacitor c=3.37896e-19 \
 //x=3.825 //y=0.37 //x2=2.505 //y2=1.655
cc_13 ( N_GND_c_2_p N_noxref_3_c_158_n ) capacitor c=0.00101801f //x=0.74 \
 //y=0 //x2=2.59 //y2=3.33
cc_14 ( N_GND_c_4_p N_noxref_3_c_159_n ) capacitor c=0.00184963f //x=5.18 \
 //y=0 //x2=4.07 //y2=2.085
cc_15 ( N_GND_c_7_p N_noxref_3_c_159_n ) capacitor c=7.87839e-19 //x=4.36 \
 //y=0.535 //x2=4.07 //y2=2.085
cc_16 ( N_GND_c_1_p N_noxref_3_c_159_n ) capacitor c=0.00118981f //x=5.18 \
 //y=0 //x2=4.07 //y2=2.085
cc_17 ( N_GND_c_3_p N_noxref_3_c_159_n ) capacitor c=0.029021f //x=3.33 //y=0 \
 //x2=4.07 //y2=2.085
cc_18 ( N_GND_M2_noxref_s N_noxref_3_c_159_n ) capacitor c=0.0108503f \
 //x=3.825 //y=0.37 //x2=4.07 //y2=2.085
cc_19 ( N_GND_c_7_p N_noxref_3_c_164_n ) capacitor c=0.0121757f //x=4.36 \
 //y=0.535 //x2=4.18 //y2=0.91
cc_20 ( N_GND_M2_noxref_s N_noxref_3_c_164_n ) capacitor c=0.0317689f \
 //x=3.825 //y=0.37 //x2=4.18 //y2=0.91
cc_21 ( N_GND_c_3_p N_noxref_3_c_166_n ) capacitor c=0.00562003f //x=3.33 \
 //y=0 //x2=4.18 //y2=1.92
cc_22 ( N_GND_M2_noxref_s N_noxref_3_c_167_n ) capacitor c=0.00483274f \
 //x=3.825 //y=0.37 //x2=4.555 //y2=0.755
cc_23 ( N_GND_c_23_p N_noxref_3_c_168_n ) capacitor c=0.0118602f //x=4.845 \
 //y=0.535 //x2=4.71 //y2=0.91
cc_24 ( N_GND_M2_noxref_s N_noxref_3_c_168_n ) capacitor c=0.0143355f \
 //x=3.825 //y=0.37 //x2=4.71 //y2=0.91
cc_25 ( N_GND_M2_noxref_s N_noxref_3_c_170_n ) capacitor c=0.0074042f \
 //x=3.825 //y=0.37 //x2=4.71 //y2=1.255
cc_26 ( N_GND_c_7_p N_noxref_3_c_171_n ) capacitor c=2.1838e-19 //x=4.36 \
 //y=0.535 //x2=4.07 //y2=2.085
cc_27 ( N_GND_c_3_p N_noxref_3_c_171_n ) capacitor c=0.0108179f //x=3.33 //y=0 \
 //x2=4.07 //y2=2.085
cc_28 ( N_GND_M2_noxref_s N_noxref_3_c_171_n ) capacitor c=0.00655738f \
 //x=3.825 //y=0.37 //x2=4.07 //y2=2.085
cc_29 ( N_GND_c_2_p N_noxref_3_M1_noxref_d ) capacitor c=8.58106e-19 //x=0.74 \
 //y=0 //x2=1.96 //y2=0.905
cc_30 ( N_GND_c_3_p N_noxref_3_M1_noxref_d ) capacitor c=0.00616547f //x=3.33 \
 //y=0 //x2=1.96 //y2=0.905
cc_31 ( N_GND_M0_noxref_d N_noxref_3_M1_noxref_d ) capacitor c=0.00143464f \
 //x=0.99 //y=0.865 //x2=1.96 //y2=0.905
cc_32 ( N_GND_M2_noxref_s N_noxref_3_M1_noxref_d ) capacitor c=2.09402e-19 \
 //x=3.825 //y=0.37 //x2=1.96 //y2=0.905
cc_33 ( N_GND_c_2_p N_A_c_281_n ) capacitor c=0.0180518f //x=0.74 //y=0 \
 //x2=1.11 //y2=2.08
cc_34 ( N_GND_c_34_p N_A_c_282_n ) capacitor c=0.00135046f //x=1.095 //y=0 \
 //x2=0.915 //y2=0.865
cc_35 ( N_GND_M0_noxref_d N_A_c_282_n ) capacitor c=0.00220047f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=0.865
cc_36 ( N_GND_M0_noxref_d N_A_c_284_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=1.21
cc_37 ( N_GND_c_2_p N_A_c_285_n ) capacitor c=0.00264481f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.52
cc_38 ( N_GND_c_2_p N_A_c_286_n ) capacitor c=0.0121947f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.915
cc_39 ( N_GND_M0_noxref_d N_A_c_287_n ) capacitor c=0.0131326f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=0.71
cc_40 ( N_GND_M0_noxref_d N_A_c_288_n ) capacitor c=0.00193127f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=1.365
cc_41 ( N_GND_c_5_p N_A_c_289_n ) capacitor c=0.00130622f //x=3.16 //y=0 \
 //x2=1.445 //y2=0.865
cc_42 ( N_GND_M0_noxref_d N_A_c_289_n ) capacitor c=0.00257848f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=0.865
cc_43 ( N_GND_M0_noxref_d N_A_c_291_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=1.21
cc_44 ( N_GND_c_2_p N_B_c_337_n ) capacitor c=9.2064e-19 //x=0.74 //y=0 \
 //x2=1.85 //y2=2.08
cc_45 ( N_GND_c_3_p N_B_c_337_n ) capacitor c=9.53263e-19 //x=3.33 //y=0 \
 //x2=1.85 //y2=2.08
cc_46 ( N_GND_c_4_p N_noxref_6_c_401_n ) capacitor c=0.00710948f //x=5.18 \
 //y=0 //x2=1.58 //y2=1.58
cc_47 ( N_GND_c_34_p N_noxref_6_c_401_n ) capacitor c=0.00111428f //x=1.095 \
 //y=0 //x2=1.58 //y2=1.58
cc_48 ( N_GND_c_5_p N_noxref_6_c_401_n ) capacitor c=0.00180846f //x=3.16 \
 //y=0 //x2=1.58 //y2=1.58
cc_49 ( N_GND_M0_noxref_d N_noxref_6_c_401_n ) capacitor c=0.0090983f //x=0.99 \
 //y=0.865 //x2=1.58 //y2=1.58
cc_50 ( N_GND_c_4_p N_noxref_6_c_405_n ) capacitor c=0.00723598f //x=5.18 \
 //y=0 //x2=1.665 //y2=0.615
cc_51 ( N_GND_c_5_p N_noxref_6_c_405_n ) capacitor c=0.0146208f //x=3.16 //y=0 \
 //x2=1.665 //y2=0.615
cc_52 ( N_GND_c_1_p N_noxref_6_c_405_n ) capacitor c=0.00145873f //x=5.18 \
 //y=0 //x2=1.665 //y2=0.615
cc_53 ( N_GND_M0_noxref_d N_noxref_6_c_405_n ) capacitor c=0.033812f //x=0.99 \
 //y=0.865 //x2=1.665 //y2=0.615
cc_54 ( N_GND_c_2_p N_noxref_6_c_409_n ) capacitor c=2.91423e-19 //x=0.74 \
 //y=0 //x2=1.665 //y2=1.495
cc_55 ( N_GND_c_4_p N_noxref_6_c_410_n ) capacitor c=0.0182925f //x=5.18 //y=0 \
 //x2=2.55 //y2=0.53
cc_56 ( N_GND_c_5_p N_noxref_6_c_410_n ) capacitor c=0.0373121f //x=3.16 //y=0 \
 //x2=2.55 //y2=0.53
cc_57 ( N_GND_c_1_p N_noxref_6_c_410_n ) capacitor c=0.00198448f //x=5.18 \
 //y=0 //x2=2.55 //y2=0.53
cc_58 ( N_GND_c_4_p N_noxref_6_c_413_n ) capacitor c=0.00292576f //x=5.18 \
 //y=0 //x2=2.635 //y2=0.615
cc_59 ( N_GND_c_5_p N_noxref_6_c_413_n ) capacitor c=0.0148673f //x=3.16 //y=0 \
 //x2=2.635 //y2=0.615
cc_60 ( N_GND_c_60_p N_noxref_6_c_413_n ) capacitor c=9.77746e-19 //x=3.96 \
 //y=0.45 //x2=2.635 //y2=0.615
cc_61 ( N_GND_c_1_p N_noxref_6_c_413_n ) capacitor c=0.00145015f //x=5.18 \
 //y=0 //x2=2.635 //y2=0.615
cc_62 ( N_GND_c_3_p N_noxref_6_c_413_n ) capacitor c=0.0431718f //x=3.33 //y=0 \
 //x2=2.635 //y2=0.615
cc_63 ( N_GND_c_4_p N_noxref_6_M0_noxref_s ) capacitor c=0.00723598f //x=5.18 \
 //y=0 //x2=0.56 //y2=0.365
cc_64 ( N_GND_c_34_p N_noxref_6_M0_noxref_s ) capacitor c=0.0146208f //x=1.095 \
 //y=0 //x2=0.56 //y2=0.365
cc_65 ( N_GND_c_2_p N_noxref_6_M0_noxref_s ) capacitor c=0.0594057f //x=0.74 \
 //y=0 //x2=0.56 //y2=0.365
cc_66 ( N_GND_c_1_p N_noxref_6_M0_noxref_s ) capacitor c=0.00145873f //x=5.18 \
 //y=0 //x2=0.56 //y2=0.365
cc_67 ( N_GND_c_3_p N_noxref_6_M0_noxref_s ) capacitor c=0.00198098f //x=3.33 \
 //y=0 //x2=0.56 //y2=0.365
cc_68 ( N_GND_M0_noxref_d N_noxref_6_M0_noxref_s ) capacitor c=0.0334197f \
 //x=0.99 //y=0.865 //x2=0.56 //y2=0.365
cc_69 ( N_GND_M2_noxref_s N_noxref_6_M0_noxref_s ) capacitor c=9.77746e-19 \
 //x=3.825 //y=0.37 //x2=0.56 //y2=0.365
cc_70 ( N_GND_c_3_p Y ) capacitor c=8.10282e-19 //x=3.33 //y=0 //x2=4.81 \
 //y2=2.22
cc_71 ( N_GND_c_4_p N_Y_c_452_n ) capacitor c=0.00180637f //x=5.18 //y=0 \
 //x2=4.725 //y2=2.08
cc_72 ( N_GND_c_1_p N_Y_c_452_n ) capacitor c=0.0301661f //x=5.18 //y=0 \
 //x2=4.725 //y2=2.08
cc_73 ( N_GND_M2_noxref_s N_Y_c_452_n ) capacitor c=0.00999304f //x=3.825 \
 //y=0.37 //x2=4.725 //y2=2.08
cc_74 ( N_GND_c_4_p N_Y_M2_noxref_d ) capacitor c=0.00194883f //x=5.18 //y=0 \
 //x2=4.255 //y2=0.91
cc_75 ( N_GND_c_7_p N_Y_M2_noxref_d ) capacitor c=0.0146043f //x=4.36 \
 //y=0.535 //x2=4.255 //y2=0.91
cc_76 ( N_GND_c_1_p N_Y_M2_noxref_d ) capacitor c=0.00973758f //x=5.18 //y=0 \
 //x2=4.255 //y2=0.91
cc_77 ( N_GND_c_3_p N_Y_M2_noxref_d ) capacitor c=0.00924905f //x=3.33 //y=0 \
 //x2=4.255 //y2=0.91
cc_78 ( N_GND_M2_noxref_s N_Y_M2_noxref_d ) capacitor c=0.076995f //x=3.825 \
 //y=0.37 //x2=4.255 //y2=0.91
cc_79 ( N_VDD_c_82_p N_noxref_3_c_149_n ) capacitor c=0.00920603f //x=5.18 \
 //y=7.4 //x2=3.955 //y2=3.33
cc_80 ( N_VDD_c_81_n N_noxref_3_c_149_n ) capacitor c=0.0069465f //x=3.33 \
 //y=7.4 //x2=3.955 //y2=3.33
cc_81 ( N_VDD_M7_noxref_s N_noxref_3_c_149_n ) capacitor c=0.00106085f \
 //x=3.87 //y=5.02 //x2=3.955 //y2=3.33
cc_82 ( N_VDD_c_82_p N_noxref_3_c_155_n ) capacitor c=0.00161874f //x=5.18 \
 //y=7.4 //x2=2.705 //y2=3.33
cc_83 ( N_VDD_M6_noxref_d N_noxref_3_c_155_n ) capacitor c=3.3085e-19 \
 //x=2.405 //y=5.02 //x2=2.705 //y2=3.33
cc_84 ( N_VDD_c_82_p N_noxref_3_c_183_n ) capacitor c=0.00596529f //x=5.18 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_85 ( N_VDD_c_88_p N_noxref_3_c_183_n ) capacitor c=4.3394e-19 //x=1.585 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_86 ( N_VDD_c_89_p N_noxref_3_c_183_n ) capacitor c=4.3394e-19 //x=2.465 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_87 ( N_VDD_M4_noxref_d N_noxref_3_c_183_n ) capacitor c=0.0131293f \
 //x=1.525 //y=5.02 //x2=2.025 //y2=5.2
cc_88 ( N_VDD_c_80_n N_noxref_3_c_187_n ) capacitor c=0.00989999f //x=0.74 \
 //y=7.4 //x2=1.315 //y2=5.2
cc_89 ( N_VDD_M3_noxref_s N_noxref_3_c_187_n ) capacitor c=0.087833f //x=0.655 \
 //y=5.02 //x2=1.315 //y2=5.2
cc_90 ( N_VDD_c_82_p N_noxref_3_c_189_n ) capacitor c=0.00362183f //x=5.18 \
 //y=7.4 //x2=2.505 //y2=5.2
cc_91 ( N_VDD_c_89_p N_noxref_3_c_189_n ) capacitor c=7.21492e-19 //x=2.465 \
 //y=7.4 //x2=2.505 //y2=5.2
cc_92 ( N_VDD_M6_noxref_d N_noxref_3_c_189_n ) capacitor c=0.016468f //x=2.405 \
 //y=5.02 //x2=2.505 //y2=5.2
cc_93 ( N_VDD_c_80_n N_noxref_3_c_158_n ) capacitor c=0.00159771f //x=0.74 \
 //y=7.4 //x2=2.59 //y2=3.33
cc_94 ( N_VDD_c_81_n N_noxref_3_c_158_n ) capacitor c=0.0461201f //x=3.33 \
 //y=7.4 //x2=2.59 //y2=3.33
cc_95 ( N_VDD_c_82_p N_noxref_3_c_159_n ) capacitor c=0.00160122f //x=5.18 \
 //y=7.4 //x2=4.07 //y2=2.085
cc_96 ( N_VDD_c_79_n N_noxref_3_c_159_n ) capacitor c=0.00144809f //x=5.18 \
 //y=7.4 //x2=4.07 //y2=2.085
cc_97 ( N_VDD_c_81_n N_noxref_3_c_159_n ) capacitor c=0.0272885f //x=3.33 \
 //y=7.4 //x2=4.07 //y2=2.085
cc_98 ( N_VDD_M7_noxref_s N_noxref_3_c_159_n ) capacitor c=0.00971593f \
 //x=3.87 //y=5.02 //x2=4.07 //y2=2.085
cc_99 ( N_VDD_c_102_p N_noxref_3_M7_noxref_g ) capacitor c=0.00748034f //x=4.8 \
 //y=7.4 //x2=4.225 //y2=6.02
cc_100 ( N_VDD_c_81_n N_noxref_3_M7_noxref_g ) capacitor c=0.00895557f \
 //x=3.33 //y=7.4 //x2=4.225 //y2=6.02
cc_101 ( N_VDD_M7_noxref_s N_noxref_3_M7_noxref_g ) capacitor c=0.0528676f \
 //x=3.87 //y=5.02 //x2=4.225 //y2=6.02
cc_102 ( N_VDD_c_102_p N_noxref_3_M8_noxref_g ) capacitor c=0.00697478f \
 //x=4.8 //y=7.4 //x2=4.665 //y2=6.02
cc_103 ( N_VDD_M8_noxref_d N_noxref_3_M8_noxref_g ) capacitor c=0.0528676f \
 //x=4.74 //y=5.02 //x2=4.665 //y2=6.02
cc_104 ( N_VDD_c_79_n N_noxref_3_c_203_n ) capacitor c=0.0287802f //x=5.18 \
 //y=7.4 //x2=4.59 //y2=4.79
cc_105 ( N_VDD_c_81_n N_noxref_3_c_204_n ) capacitor c=0.011132f //x=3.33 \
 //y=7.4 //x2=4.3 //y2=4.79
cc_106 ( N_VDD_M7_noxref_s N_noxref_3_c_204_n ) capacitor c=0.00527247f \
 //x=3.87 //y=5.02 //x2=4.3 //y2=4.79
cc_107 ( N_VDD_c_82_p N_noxref_3_M3_noxref_d ) capacitor c=0.00706239f \
 //x=5.18 //y=7.4 //x2=1.085 //y2=5.02
cc_108 ( N_VDD_c_88_p N_noxref_3_M3_noxref_d ) capacitor c=0.0138103f \
 //x=1.585 //y=7.4 //x2=1.085 //y2=5.02
cc_109 ( N_VDD_c_79_n N_noxref_3_M3_noxref_d ) capacitor c=0.00135231f \
 //x=5.18 //y=7.4 //x2=1.085 //y2=5.02
cc_110 ( N_VDD_c_81_n N_noxref_3_M3_noxref_d ) capacitor c=6.94454e-19 \
 //x=3.33 //y=7.4 //x2=1.085 //y2=5.02
cc_111 ( N_VDD_M4_noxref_d N_noxref_3_M3_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.085 //y2=5.02
cc_112 ( N_VDD_c_82_p N_noxref_3_M5_noxref_d ) capacitor c=0.00706239f \
 //x=5.18 //y=7.4 //x2=1.965 //y2=5.02
cc_113 ( N_VDD_c_89_p N_noxref_3_M5_noxref_d ) capacitor c=0.0138379f \
 //x=2.465 //y=7.4 //x2=1.965 //y2=5.02
cc_114 ( N_VDD_c_79_n N_noxref_3_M5_noxref_d ) capacitor c=0.00135231f \
 //x=5.18 //y=7.4 //x2=1.965 //y2=5.02
cc_115 ( N_VDD_c_81_n N_noxref_3_M5_noxref_d ) capacitor c=0.0120541f //x=3.33 \
 //y=7.4 //x2=1.965 //y2=5.02
cc_116 ( N_VDD_M3_noxref_s N_noxref_3_M5_noxref_d ) capacitor c=0.00111971f \
 //x=0.655 //y=5.02 //x2=1.965 //y2=5.02
cc_117 ( N_VDD_M4_noxref_d N_noxref_3_M5_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.965 //y2=5.02
cc_118 ( N_VDD_M6_noxref_d N_noxref_3_M5_noxref_d ) capacitor c=0.0664752f \
 //x=2.405 //y=5.02 //x2=1.965 //y2=5.02
cc_119 ( N_VDD_M7_noxref_s N_noxref_3_M5_noxref_d ) capacitor c=5.1407e-19 \
 //x=3.87 //y=5.02 //x2=1.965 //y2=5.02
cc_120 ( N_VDD_c_82_p N_A_c_281_n ) capacitor c=0.00140404f //x=5.18 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_121 ( N_VDD_c_88_p N_A_c_281_n ) capacitor c=2.63811e-19 //x=1.585 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_122 ( N_VDD_c_80_n N_A_c_281_n ) capacitor c=0.016845f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_123 ( N_VDD_c_88_p N_A_M3_noxref_g ) capacitor c=0.00726866f //x=1.585 \
 //y=7.4 //x2=1.01 //y2=6.02
cc_124 ( N_VDD_M3_noxref_s N_A_M3_noxref_g ) capacitor c=0.054195f //x=0.655 \
 //y=5.02 //x2=1.01 //y2=6.02
cc_125 ( N_VDD_c_88_p N_A_M4_noxref_g ) capacitor c=0.00672952f //x=1.585 \
 //y=7.4 //x2=1.45 //y2=6.02
cc_126 ( N_VDD_M4_noxref_d N_A_M4_noxref_g ) capacitor c=0.015318f //x=1.525 \
 //y=5.02 //x2=1.45 //y2=6.02
cc_127 ( N_VDD_c_80_n N_A_c_299_n ) capacitor c=0.0292267f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=4.7
cc_128 ( N_VDD_c_80_n N_B_c_337_n ) capacitor c=6.61004e-19 //x=0.74 //y=7.4 \
 //x2=1.85 //y2=2.08
cc_129 ( N_VDD_c_81_n N_B_c_337_n ) capacitor c=6.09526e-19 //x=3.33 //y=7.4 \
 //x2=1.85 //y2=2.08
cc_130 ( N_VDD_c_89_p N_B_M5_noxref_g ) capacitor c=0.00673971f //x=2.465 \
 //y=7.4 //x2=1.89 //y2=6.02
cc_131 ( N_VDD_M4_noxref_d N_B_M5_noxref_g ) capacitor c=0.015318f //x=1.525 \
 //y=5.02 //x2=1.89 //y2=6.02
cc_132 ( N_VDD_c_89_p N_B_M6_noxref_g ) capacitor c=0.00672952f //x=2.465 \
 //y=7.4 //x2=2.33 //y2=6.02
cc_133 ( N_VDD_c_81_n N_B_M6_noxref_g ) capacitor c=0.00904525f //x=3.33 \
 //y=7.4 //x2=2.33 //y2=6.02
cc_134 ( N_VDD_M6_noxref_d N_B_M6_noxref_g ) capacitor c=0.0430452f //x=2.405 \
 //y=5.02 //x2=2.33 //y2=6.02
cc_135 ( N_VDD_c_79_n Y ) capacitor c=0.0232778f //x=5.18 //y=7.4 //x2=4.81 \
 //y2=2.22
cc_136 ( N_VDD_c_81_n Y ) capacitor c=4.80934e-19 //x=3.33 //y=7.4 //x2=4.81 \
 //y2=2.22
cc_137 ( N_VDD_c_82_p N_Y_c_462_n ) capacitor c=0.00190861f //x=5.18 //y=7.4 \
 //x2=4.725 //y2=4.58
cc_138 ( N_VDD_c_102_p N_Y_c_462_n ) capacitor c=8.8179e-19 //x=4.8 //y=7.4 \
 //x2=4.725 //y2=4.58
cc_139 ( N_VDD_M8_noxref_d N_Y_c_462_n ) capacitor c=0.00641434f //x=4.74 \
 //y=5.02 //x2=4.725 //y2=4.58
cc_140 ( N_VDD_c_81_n N_Y_c_465_n ) capacitor c=0.017572f //x=3.33 //y=7.4 \
 //x2=4.53 //y2=4.58
cc_141 ( N_VDD_c_82_p N_Y_M7_noxref_d ) capacitor c=0.00708604f //x=5.18 \
 //y=7.4 //x2=4.3 //y2=5.02
cc_142 ( N_VDD_c_102_p N_Y_M7_noxref_d ) capacitor c=0.0139004f //x=4.8 \
 //y=7.4 //x2=4.3 //y2=5.02
cc_143 ( N_VDD_c_79_n N_Y_M7_noxref_d ) capacitor c=0.0219131f //x=5.18 \
 //y=7.4 //x2=4.3 //y2=5.02
cc_144 ( N_VDD_M7_noxref_s N_Y_M7_noxref_d ) capacitor c=0.0843065f //x=3.87 \
 //y=5.02 //x2=4.3 //y2=5.02
cc_145 ( N_VDD_M8_noxref_d N_Y_M7_noxref_d ) capacitor c=0.0832641f //x=4.74 \
 //y=5.02 //x2=4.3 //y2=5.02
cc_146 ( N_noxref_3_c_187_n N_A_c_281_n ) capacitor c=0.00569255f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=2.08
cc_147 ( N_noxref_3_c_158_n N_A_c_281_n ) capacitor c=0.00407922f //x=2.59 \
 //y=3.33 //x2=1.11 //y2=2.08
cc_148 ( N_noxref_3_c_187_n N_A_M3_noxref_g ) capacitor c=0.0177326f //x=1.315 \
 //y=5.2 //x2=1.01 //y2=6.02
cc_149 ( N_noxref_3_c_183_n N_A_M4_noxref_g ) capacitor c=0.0203837f //x=2.025 \
 //y=5.2 //x2=1.45 //y2=6.02
cc_150 ( N_noxref_3_M3_noxref_d N_A_M4_noxref_g ) capacitor c=0.0173476f \
 //x=1.085 //y=5.02 //x2=1.45 //y2=6.02
cc_151 ( N_noxref_3_c_187_n N_A_c_299_n ) capacitor c=0.00571434f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=4.7
cc_152 ( N_noxref_3_c_183_n N_B_c_346_n ) capacitor c=0.0130171f //x=2.025 \
 //y=5.2 //x2=1.85 //y2=4.535
cc_153 ( N_noxref_3_c_158_n N_B_c_346_n ) capacitor c=0.0101115f //x=2.59 \
 //y=3.33 //x2=1.85 //y2=4.535
cc_154 ( N_noxref_3_c_155_n N_B_c_337_n ) capacitor c=0.00717888f //x=2.705 \
 //y=3.33 //x2=1.85 //y2=2.08
cc_155 ( N_noxref_3_c_158_n N_B_c_337_n ) capacitor c=0.0813981f //x=2.59 \
 //y=3.33 //x2=1.85 //y2=2.08
cc_156 ( N_noxref_3_c_159_n N_B_c_337_n ) capacitor c=0.00126776f //x=4.07 \
 //y=2.085 //x2=1.85 //y2=2.08
cc_157 ( N_noxref_3_c_183_n N_B_M5_noxref_g ) capacitor c=0.0166421f //x=2.025 \
 //y=5.2 //x2=1.89 //y2=6.02
cc_158 ( N_noxref_3_M5_noxref_d N_B_M5_noxref_g ) capacitor c=0.0173476f \
 //x=1.965 //y=5.02 //x2=1.89 //y2=6.02
cc_159 ( N_noxref_3_c_189_n N_B_M6_noxref_g ) capacitor c=0.0223536f //x=2.505 \
 //y=5.2 //x2=2.33 //y2=6.02
cc_160 ( N_noxref_3_M5_noxref_d N_B_M6_noxref_g ) capacitor c=0.0179769f \
 //x=1.965 //y=5.02 //x2=2.33 //y2=6.02
cc_161 ( N_noxref_3_M1_noxref_d N_B_c_355_n ) capacitor c=0.00217566f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=0.905
cc_162 ( N_noxref_3_M1_noxref_d N_B_c_356_n ) capacitor c=0.0034598f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.25
cc_163 ( N_noxref_3_M1_noxref_d N_B_c_357_n ) capacitor c=0.0065582f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.56
cc_164 ( N_noxref_3_c_158_n N_B_c_358_n ) capacitor c=0.0142673f //x=2.59 \
 //y=3.33 //x2=2.255 //y2=4.79
cc_165 ( N_noxref_3_c_238_p N_B_c_358_n ) capacitor c=0.00414324f //x=2.11 \
 //y=5.2 //x2=2.255 //y2=4.79
cc_166 ( N_noxref_3_M1_noxref_d N_B_c_360_n ) capacitor c=0.00241102f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=0.75
cc_167 ( N_noxref_3_c_156_n N_B_c_361_n ) capacitor c=0.00359704f //x=2.505 \
 //y=1.655 //x2=2.26 //y2=1.405
cc_168 ( N_noxref_3_M1_noxref_d N_B_c_361_n ) capacitor c=0.0138845f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=1.405
cc_169 ( N_noxref_3_M1_noxref_d N_B_c_363_n ) capacitor c=0.00132245f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=0.905
cc_170 ( N_noxref_3_c_156_n N_B_c_364_n ) capacitor c=0.00457401f //x=2.505 \
 //y=1.655 //x2=2.415 //y2=1.25
cc_171 ( N_noxref_3_M1_noxref_d N_B_c_364_n ) capacitor c=0.00566463f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=1.25
cc_172 ( N_noxref_3_c_158_n N_B_c_366_n ) capacitor c=0.00877984f //x=2.59 \
 //y=3.33 //x2=1.85 //y2=2.08
cc_173 ( N_noxref_3_c_158_n N_B_c_367_n ) capacitor c=0.00306024f //x=2.59 \
 //y=3.33 //x2=1.85 //y2=1.915
cc_174 ( N_noxref_3_M1_noxref_d N_B_c_367_n ) capacitor c=0.00660593f //x=1.96 \
 //y=0.905 //x2=1.85 //y2=1.915
cc_175 ( N_noxref_3_c_183_n N_B_c_369_n ) capacitor c=0.00344394f //x=2.025 \
 //y=5.2 //x2=1.88 //y2=4.7
cc_176 ( N_noxref_3_c_158_n N_B_c_369_n ) capacitor c=0.00533692f //x=2.59 \
 //y=3.33 //x2=1.88 //y2=4.7
cc_177 ( N_noxref_3_c_250_p N_noxref_6_c_425_n ) capacitor c=3.15806e-19 \
 //x=2.235 //y=1.655 //x2=0.695 //y2=1.495
cc_178 ( N_noxref_3_c_250_p N_noxref_6_c_409_n ) capacitor c=0.0201674f \
 //x=2.235 //y=1.655 //x2=1.665 //y2=1.495
cc_179 ( N_noxref_3_c_156_n N_noxref_6_c_410_n ) capacitor c=0.0046844f \
 //x=2.505 //y=1.655 //x2=2.55 //y2=0.53
cc_180 ( N_noxref_3_M1_noxref_d N_noxref_6_c_410_n ) capacitor c=0.0118355f \
 //x=1.96 //y=0.905 //x2=2.55 //y2=0.53
cc_181 ( N_noxref_3_c_155_n N_noxref_6_M0_noxref_s ) capacitor c=3.12455e-19 \
 //x=2.705 //y=3.33 //x2=0.56 //y2=0.365
cc_182 ( N_noxref_3_c_156_n N_noxref_6_M0_noxref_s ) capacitor c=0.0141735f \
 //x=2.505 //y=1.655 //x2=0.56 //y2=0.365
cc_183 ( N_noxref_3_M1_noxref_d N_noxref_6_M0_noxref_s ) capacitor \
 c=0.0437911f //x=1.96 //y=0.905 //x2=0.56 //y2=0.365
cc_184 ( N_noxref_3_c_149_n Y ) capacitor c=0.00582634f //x=3.955 //y=3.33 \
 //x2=4.81 //y2=2.22
cc_185 ( N_noxref_3_c_158_n Y ) capacitor c=0.00126776f //x=2.59 //y=3.33 \
 //x2=4.81 //y2=2.22
cc_186 ( N_noxref_3_c_159_n Y ) capacitor c=0.0711303f //x=4.07 //y=2.085 \
 //x2=4.81 //y2=2.22
cc_187 ( N_noxref_3_c_171_n Y ) capacitor c=8.49451e-19 //x=4.07 //y=2.085 \
 //x2=4.81 //y2=2.22
cc_188 ( N_noxref_3_c_261_p N_Y_c_452_n ) capacitor c=0.0023507f //x=4.555 \
 //y=1.41 //x2=4.725 //y2=2.08
cc_189 ( N_noxref_3_c_171_n N_Y_c_476_n ) capacitor c=0.0167852f //x=4.07 \
 //y=2.085 //x2=4.525 //y2=2.08
cc_190 ( N_noxref_3_c_203_n N_Y_c_462_n ) capacitor c=0.0101013f //x=4.59 \
 //y=4.79 //x2=4.725 //y2=4.58
cc_191 ( N_noxref_3_c_159_n N_Y_c_465_n ) capacitor c=0.0250789f //x=4.07 \
 //y=2.085 //x2=4.53 //y2=4.58
cc_192 ( N_noxref_3_c_204_n N_Y_c_465_n ) capacitor c=0.00962086f //x=4.3 \
 //y=4.79 //x2=4.53 //y2=4.58
cc_193 ( N_noxref_3_c_158_n N_Y_M2_noxref_d ) capacitor c=3.35192e-19 //x=2.59 \
 //y=3.33 //x2=4.255 //y2=0.91
cc_194 ( N_noxref_3_c_159_n N_Y_M2_noxref_d ) capacitor c=0.0175773f //x=4.07 \
 //y=2.085 //x2=4.255 //y2=0.91
cc_195 ( N_noxref_3_c_164_n N_Y_M2_noxref_d ) capacitor c=0.00218556f //x=4.18 \
 //y=0.91 //x2=4.255 //y2=0.91
cc_196 ( N_noxref_3_c_269_p N_Y_M2_noxref_d ) capacitor c=0.00347355f //x=4.18 \
 //y=1.255 //x2=4.255 //y2=0.91
cc_197 ( N_noxref_3_c_270_p N_Y_M2_noxref_d ) capacitor c=0.00742431f //x=4.18 \
 //y=1.565 //x2=4.255 //y2=0.91
cc_198 ( N_noxref_3_c_166_n N_Y_M2_noxref_d ) capacitor c=0.00957707f //x=4.18 \
 //y=1.92 //x2=4.255 //y2=0.91
cc_199 ( N_noxref_3_c_167_n N_Y_M2_noxref_d ) capacitor c=0.00220879f \
 //x=4.555 //y=0.755 //x2=4.255 //y2=0.91
cc_200 ( N_noxref_3_c_261_p N_Y_M2_noxref_d ) capacitor c=0.0138447f //x=4.555 \
 //y=1.41 //x2=4.255 //y2=0.91
cc_201 ( N_noxref_3_c_168_n N_Y_M2_noxref_d ) capacitor c=0.00218624f //x=4.71 \
 //y=0.91 //x2=4.255 //y2=0.91
cc_202 ( N_noxref_3_c_170_n N_Y_M2_noxref_d ) capacitor c=0.00601286f //x=4.71 \
 //y=1.255 //x2=4.255 //y2=0.91
cc_203 ( N_noxref_3_c_158_n N_Y_M7_noxref_d ) capacitor c=6.3502e-19 //x=2.59 \
 //y=3.33 //x2=4.3 //y2=5.02
cc_204 ( N_noxref_3_M7_noxref_g N_Y_M7_noxref_d ) capacitor c=0.0219309f \
 //x=4.225 //y=6.02 //x2=4.3 //y2=5.02
cc_205 ( N_noxref_3_M8_noxref_g N_Y_M7_noxref_d ) capacitor c=0.021902f \
 //x=4.665 //y=6.02 //x2=4.3 //y2=5.02
cc_206 ( N_noxref_3_c_203_n N_Y_M7_noxref_d ) capacitor c=0.0148755f //x=4.59 \
 //y=4.79 //x2=4.3 //y2=5.02
cc_207 ( N_noxref_3_c_204_n N_Y_M7_noxref_d ) capacitor c=0.00307344f //x=4.3 \
 //y=4.79 //x2=4.3 //y2=5.02
cc_208 ( N_A_c_281_n N_B_c_346_n ) capacitor c=0.00400249f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=4.535
cc_209 ( N_A_c_299_n N_B_c_346_n ) capacitor c=0.00417994f //x=1.11 //y=4.7 \
 //x2=1.85 //y2=4.535
cc_210 ( N_A_c_281_n N_B_c_337_n ) capacitor c=0.0887263f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_211 ( N_A_c_286_n N_B_c_337_n ) capacitor c=0.00308814f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_212 ( N_A_M3_noxref_g N_B_M5_noxref_g ) capacitor c=0.0104611f //x=1.01 \
 //y=6.02 //x2=1.89 //y2=6.02
cc_213 ( N_A_M4_noxref_g N_B_M5_noxref_g ) capacitor c=0.106811f //x=1.45 \
 //y=6.02 //x2=1.89 //y2=6.02
cc_214 ( N_A_M4_noxref_g N_B_M6_noxref_g ) capacitor c=0.0100341f //x=1.45 \
 //y=6.02 //x2=2.33 //y2=6.02
cc_215 ( N_A_c_282_n N_B_c_355_n ) capacitor c=4.86506e-19 //x=0.915 //y=0.865 \
 //x2=1.885 //y2=0.905
cc_216 ( N_A_c_284_n N_B_c_355_n ) capacitor c=0.00152104f //x=0.915 //y=1.21 \
 //x2=1.885 //y2=0.905
cc_217 ( N_A_c_289_n N_B_c_355_n ) capacitor c=0.0151475f //x=1.445 //y=0.865 \
 //x2=1.885 //y2=0.905
cc_218 ( N_A_c_285_n N_B_c_356_n ) capacitor c=0.00109982f //x=0.915 //y=1.52 \
 //x2=1.885 //y2=1.25
cc_219 ( N_A_c_291_n N_B_c_356_n ) capacitor c=0.0111064f //x=1.445 //y=1.21 \
 //x2=1.885 //y2=1.25
cc_220 ( N_A_c_285_n N_B_c_357_n ) capacitor c=9.57794e-19 //x=0.915 //y=1.52 \
 //x2=1.885 //y2=1.56
cc_221 ( N_A_c_286_n N_B_c_357_n ) capacitor c=0.00662747f //x=0.915 //y=1.915 \
 //x2=1.885 //y2=1.56
cc_222 ( N_A_c_291_n N_B_c_357_n ) capacitor c=0.00862358f //x=1.445 //y=1.21 \
 //x2=1.885 //y2=1.56
cc_223 ( N_A_c_289_n N_B_c_363_n ) capacitor c=0.00124821f //x=1.445 //y=0.865 \
 //x2=2.415 //y2=0.905
cc_224 ( N_A_c_291_n N_B_c_364_n ) capacitor c=0.00200715f //x=1.445 //y=1.21 \
 //x2=2.415 //y2=1.25
cc_225 ( N_A_c_281_n N_B_c_366_n ) capacitor c=0.00307062f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_226 ( N_A_c_286_n N_B_c_366_n ) capacitor c=0.0179092f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_227 ( N_A_c_281_n N_B_c_369_n ) capacitor c=0.00344981f //x=1.11 //y=2.08 \
 //x2=1.88 //y2=4.7
cc_228 ( N_A_c_299_n N_B_c_369_n ) capacitor c=0.0293367f //x=1.11 //y=4.7 \
 //x2=1.88 //y2=4.7
cc_229 ( N_A_c_286_n N_noxref_6_c_425_n ) capacitor c=0.0034165f //x=0.915 \
 //y=1.915 //x2=0.695 //y2=1.495
cc_230 ( N_A_c_281_n N_noxref_6_c_401_n ) capacitor c=0.0118986f //x=1.11 \
 //y=2.08 //x2=1.58 //y2=1.58
cc_231 ( N_A_c_285_n N_noxref_6_c_401_n ) capacitor c=0.00703567f //x=0.915 \
 //y=1.52 //x2=1.58 //y2=1.58
cc_232 ( N_A_c_286_n N_noxref_6_c_401_n ) capacitor c=0.0216532f //x=0.915 \
 //y=1.915 //x2=1.58 //y2=1.58
cc_233 ( N_A_c_288_n N_noxref_6_c_401_n ) capacitor c=0.00780629f //x=1.29 \
 //y=1.365 //x2=1.58 //y2=1.58
cc_234 ( N_A_c_291_n N_noxref_6_c_401_n ) capacitor c=0.00339872f //x=1.445 \
 //y=1.21 //x2=1.58 //y2=1.58
cc_235 ( N_A_c_286_n N_noxref_6_c_409_n ) capacitor c=6.71402e-19 //x=0.915 \
 //y=1.915 //x2=1.665 //y2=1.495
cc_236 ( N_A_c_282_n N_noxref_6_M0_noxref_s ) capacitor c=0.0326577f //x=0.915 \
 //y=0.865 //x2=0.56 //y2=0.365
cc_237 ( N_A_c_285_n N_noxref_6_M0_noxref_s ) capacitor c=3.48408e-19 \
 //x=0.915 //y=1.52 //x2=0.56 //y2=0.365
cc_238 ( N_A_c_289_n N_noxref_6_M0_noxref_s ) capacitor c=0.0120759f //x=1.445 \
 //y=0.865 //x2=0.56 //y2=0.365
cc_239 ( N_B_c_357_n N_noxref_6_c_409_n ) capacitor c=0.00623646f //x=1.885 \
 //y=1.56 //x2=1.665 //y2=1.495
cc_240 ( N_B_c_366_n N_noxref_6_c_409_n ) capacitor c=0.00172768f //x=1.85 \
 //y=2.08 //x2=1.665 //y2=1.495
cc_241 ( N_B_c_337_n N_noxref_6_c_410_n ) capacitor c=0.00161845f //x=1.85 \
 //y=2.08 //x2=2.55 //y2=0.53
cc_242 ( N_B_c_355_n N_noxref_6_c_410_n ) capacitor c=0.0186143f //x=1.885 \
 //y=0.905 //x2=2.55 //y2=0.53
cc_243 ( N_B_c_363_n N_noxref_6_c_410_n ) capacitor c=0.00656458f //x=2.415 \
 //y=0.905 //x2=2.55 //y2=0.53
cc_244 ( N_B_c_366_n N_noxref_6_c_410_n ) capacitor c=2.1838e-19 //x=1.85 \
 //y=2.08 //x2=2.55 //y2=0.53
cc_245 ( N_B_c_355_n N_noxref_6_M0_noxref_s ) capacitor c=0.00623646f \
 //x=1.885 //y=0.905 //x2=0.56 //y2=0.365
cc_246 ( N_B_c_363_n N_noxref_6_M0_noxref_s ) capacitor c=0.0143002f //x=2.415 \
 //y=0.905 //x2=0.56 //y2=0.365
cc_247 ( N_B_c_364_n N_noxref_6_M0_noxref_s ) capacitor c=0.00290153f \
 //x=2.415 //y=1.25 //x2=0.56 //y2=0.365
