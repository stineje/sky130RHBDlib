* SPICE3 file created from DLATCH.ext - technology: sky130A

.subckt DLATCH Q D GATE VDD GND
X0 m1_349_723# D GND GND nshort w=3 l=0.15
X1 VDD D m1_349_723# VDD pshort w=2 l=0.15
X2 m1_1459_723# and2x1_pcell_0/m1_547_649# GND GND nshort w=3 l=0.15
X3 VDD and2x1_pcell_0/m1_547_649# m1_1459_723# VDD pshort w=2 l=0.15
X4 GND m1_349_723# and2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X5 and2x1_pcell_0/m1_547_649# GATE and2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X6 VDD m1_349_723# and2x1_pcell_0/m1_547_649# VDD pshort w=2 l=0.15
X7 VDD GATE and2x1_pcell_0/m1_547_649# VDD pshort w=2 l=0.15
X8 m1_2569_797# and2x1_pcell_1/m1_547_649# GND GND nshort w=3 l=0.15
X9 VDD and2x1_pcell_1/m1_547_649# m1_2569_797# VDD pshort w=2 l=0.15
X10 GND GATE and2x1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X11 and2x1_pcell_1/m1_547_649# D and2x1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X12 VDD GATE and2x1_pcell_1/m1_547_649# VDD pshort w=2 l=0.15
X13 VDD D and2x1_pcell_1/m1_547_649# VDD pshort w=2 l=0.15
X14 VDD m1_1459_723# nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X15 Q m1_3087_723# nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X16 Q m1_1459_723# GND GND nshort w=3 l=0.15
X17 Q m1_3087_723# GND GND nshort w=3 l=0.15
X18 VDD Q nor2x1_pcell_1/a_317_1331# VDD pshort w=2 l=0.15
X19 m1_3087_723# m1_2569_797# nor2x1_pcell_1/a_317_1331# VDD pshort w=2 l=0.15
X20 m1_3087_723# Q GND GND nshort w=3 l=0.15
X21 m1_3087_723# m1_2569_797# GND GND nshort w=3 l=0.15
.ends
