* SPICE3 file created from TMRDFFQX1.ext - technology: sky130A

.subckt TMRDFFQX1 Q D CLK VDD GND
X0 VDD CLK a_277_1004 VDD pshort w=2 l=0.15 M=2
X1 a_3177_1004 a_3303_383 a_3072_73 GND nshort w=3 l=0.15
X2 a_13757_1005 a_7595_383 a_13268_181 VDD pshort w=2 l=0.15 M=2
X3 a_3177_1004 a_3303_383 VDD VDD pshort w=2 l=0.15 M=2
X4 a_4439_159 CLK a_6698_73 GND nshort w=3 l=0.15
X5 a_6137_1004 a_4439_159 a_6032_73 GND nshort w=3 l=0.15
X6 GND a_147_159 a_91_75 GND nshort w=3 l=0.15
X7 VDD CLK a_147_159 VDD pshort w=2 l=0.15 M=2
X8 a_8956_182 CLK a_8675_75 GND nshort w=3 l=0.15
X9 a_11887_383 a_8731_159 VDD VDD pshort w=2 l=0.15 M=2
X10 VDD a_11887_383 a_11761_1004 VDD pshort w=2 l=0.15 M=2
X11 a_13268_181 a_7595_383 a_14320_73 GND nshort w=3 l=0.15
X12 GND a_8861_1004 a_11656_73 GND nshort w=3 l=0.15
X13 VDD CLK a_4439_159 VDD pshort w=2 l=0.15 M=2
X14 a_9183_943 D VDD VDD pshort w=2 l=0.15 M=2
X15 GND a_10429_1004 a_10990_73 GND nshort w=3 l=0.15
X16 GND a_4439_159 a_4383_75 GND nshort w=3 l=0.15
X17 a_3303_383 a_3177_1004 VDD VDD pshort w=2 l=0.15 M=2
X18 VDD a_599_943 a_277_1004 VDD pshort w=2 l=0.15 M=2
X19 VDD a_277_1004 a_599_943 VDD pshort w=2 l=0.15 M=2
X20 a_8731_159 a_10429_1004 VDD VDD pshort w=2 l=0.15 M=2
X21 a_4569_1004 a_4891_943 VDD VDD pshort w=2 l=0.15 M=2
X22 a_13757_1005 a_3303_383 a_13268_181 VDD pshort w=2 l=0.15 M=2
X23 VDD a_147_159 a_3303_383 VDD pshort w=2 l=0.15 M=2
X24 VDD a_9183_943 a_10429_1004 VDD pshort w=2 l=0.15 M=2
X25 a_7595_383 a_7469_1004 VDD VDD pshort w=2 l=0.15 M=2
X26 VDD a_4569_1004 a_7469_1004 VDD pshort w=2 l=0.15 M=2
X27 a_1845_1004 a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X28 a_8861_1004 a_9183_943 VDD VDD pshort w=2 l=0.15 M=2
X29 VDD a_4439_159 a_4569_1004 VDD pshort w=2 l=0.15 M=2
X30 a_7595_383 a_4439_159 a_8030_73 GND nshort w=3 l=0.15
X31 GND a_4569_1004 a_5366_73 GND nshort w=3 l=0.15
X32 GND a_599_943 a_1740_73 GND nshort w=3 l=0.15
X33 a_6137_1004 a_4439_159 VDD VDD pshort w=2 l=0.15 M=2
X34 a_372_182 CLK a_91_75 GND nshort w=3 l=0.15
X35 a_9183_943 a_8861_1004 VDD VDD pshort w=2 l=0.15 M=2
X36 GND a_11887_383 a_13654_73 GND nshort w=3 l=0.15
X37 a_13093_1005 a_3303_383 a_13757_1005 VDD pshort w=2 l=0.15 M=2
X38 VDD a_7595_383 a_13093_1005 VDD pshort w=2 l=0.15 M=2
X39 GND a_11887_383 a_12988_73 GND nshort w=3 l=0.15
X40 VDD D a_599_943 VDD pshort w=2 l=0.15 M=2
X41 a_8731_159 CLK VDD VDD pshort w=2 l=0.15 M=2
X42 a_13757_1005 a_11887_383 a_13093_1005 VDD pshort w=2 l=0.15 M=2
X43 VDD a_8731_159 a_10429_1004 VDD pshort w=2 l=0.15 M=2
X44 a_4439_159 a_6137_1004 VDD VDD pshort w=2 l=0.15 M=2
X45 a_147_159 CLK a_2406_73 GND nshort w=3 l=0.15
X46 a_277_1004 a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X47 a_4664_182 CLK a_4383_75 GND nshort w=3 l=0.15
X48 VDD a_7595_383 a_7469_1004 VDD pshort w=2 l=0.15 M=2
X49 VDD CLK a_4569_1004 VDD pshort w=2 l=0.15 M=2
X50 a_9183_943 D a_9658_73 GND nshort w=3 l=0.15
X51 VDD a_599_943 a_1845_1004 VDD pshort w=2 l=0.15 M=2
X52 GND a_4569_1004 a_7364_73 GND nshort w=3 l=0.15
X53 GND a_3177_1004 a_3738_73 GND nshort w=3 l=0.15
X54 a_11761_1004 a_8861_1004 VDD VDD pshort w=2 l=0.15 M=2
X55 GND a_9183_943 a_10324_73 GND nshort w=3 l=0.15
X56 VDD a_11887_383 a_13093_1005 VDD pshort w=2 l=0.15 M=2
X57 a_4891_943 D VDD VDD pshort w=2 l=0.15 M=2
X58 a_8861_1004 a_9183_943 a_8956_182 GND nshort w=3 l=0.15
X59 a_11761_1004 a_11887_383 a_11656_73 GND nshort w=3 l=0.15
X60 GND a_277_1004 a_1074_73 GND nshort w=3 l=0.15
X61 VDD a_277_1004 a_3177_1004 VDD pshort w=2 l=0.15 M=2
X62 a_8731_159 CLK a_10990_73 GND nshort w=3 l=0.15
X63 VDD a_13268_181 Q VDD pshort w=2 l=0.15 M=2
X64 VDD a_11761_1004 a_11887_383 VDD pshort w=2 l=0.15 M=2
X65 a_4891_943 a_4569_1004 VDD VDD pshort w=2 l=0.15 M=2
X66 Q a_13268_181 GND GND nshort w=3 l=0.15
X67 a_1845_1004 a_147_159 a_1740_73 GND nshort w=3 l=0.15
X68 a_7595_383 a_4439_159 VDD VDD pshort w=2 l=0.15 M=2
X69 GND a_11761_1004 a_12322_73 GND nshort w=3 l=0.15
X70 a_8861_1004 a_8731_159 VDD VDD pshort w=2 l=0.15 M=2
X71 a_4891_943 D a_5366_73 GND nshort w=3 l=0.15
X72 a_147_159 a_1845_1004 VDD VDD pshort w=2 l=0.15 M=2
X73 VDD CLK a_8861_1004 VDD pshort w=2 l=0.15 M=2
X74 a_13268_181 a_3303_383 a_13654_73 GND nshort w=3 l=0.15
X75 VDD a_4891_943 a_6137_1004 VDD pshort w=2 l=0.15 M=2
X76 GND a_6137_1004 a_6698_73 GND nshort w=3 l=0.15
X77 GND a_277_1004 a_3072_73 GND nshort w=3 l=0.15
X78 a_13268_181 a_7595_383 a_12988_73 GND nshort w=3 l=0.15
X79 GND a_4891_943 a_6032_73 GND nshort w=3 l=0.15
X80 GND a_3303_383 a_14320_73 GND nshort w=3 l=0.15
X81 a_3303_383 a_147_159 a_3738_73 GND nshort w=3 l=0.15
X82 a_7469_1004 a_7595_383 a_7364_73 GND nshort w=3 l=0.15
X83 a_10429_1004 a_8731_159 a_10324_73 GND nshort w=3 l=0.15
X84 GND a_8731_159 a_8675_75 GND nshort w=3 l=0.15
X85 GND a_7469_1004 a_8030_73 GND nshort w=3 l=0.15
X86 a_599_943 D a_1074_73 GND nshort w=3 l=0.15
X87 a_11887_383 a_8731_159 a_12322_73 GND nshort w=3 l=0.15
X88 GND a_1845_1004 a_2406_73 GND nshort w=3 l=0.15
X89 a_277_1004 a_599_943 a_372_182 GND nshort w=3 l=0.15
X90 GND a_8861_1004 a_9658_73 GND nshort w=3 l=0.15
X91 a_4569_1004 a_4891_943 a_4664_182 GND nshort w=3 l=0.15
C0 VDD a_13093_1005 2.02fF
C1 a_277_1004 a_147_159 3.00fF
C2 a_147_159 CLK 4.49fF
C3 a_4569_1004 VDD 2.49fF
C4 a_277_1004 VDD 2.32fF
C5 a_3303_383 VDD 2.67fF
C6 D a_7595_383 2.68fF
C7 CLK VDD 5.18fF
C8 CLK a_8731_159 3.25fF
C9 a_147_159 VDD 3.05fF
C10 VDD a_11887_383 2.41fF
C11 a_4439_159 a_4569_1004 3.00fF
C12 a_3303_383 a_7595_383 2.76fF
C13 VDD a_8731_159 3.06fF
C14 a_4439_159 CLK 4.81fF
C15 a_3303_383 D 7.42fF
C16 a_7595_383 VDD 2.61fF
C17 a_4439_159 VDD 3.02fF
C18 VDD a_8861_1004 2.49fF
C19 a_8731_159 a_8861_1004 3.00fF
C20 VDD GND 36.40fF
C21 a_7595_383 GND 2.24fF **FLOATING
C22 a_3303_383 GND 3.31fF **FLOATING
.ends
