// File: DFFRNQNX1.spi.DFFRNQNX1.pxi
// Created: Tue Oct 15 15:46:14 2024
// 
simulator lang=spectre
x_PM_DFFRNQNX1\%GND ( GND N_GND_c_8_p N_GND_c_117_p N_GND_c_1_p N_GND_c_9_p \
 N_GND_c_10_p N_GND_c_58_p N_GND_c_17_p N_GND_c_24_p N_GND_c_32_p N_GND_c_39_p \
 N_GND_c_61_p N_GND_c_68_p N_GND_c_92_p N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p \
 N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p N_GND_M0_noxref_d N_GND_M3_noxref_d \
 N_GND_M6_noxref_d N_GND_M8_noxref_d N_GND_M11_noxref_d N_GND_M14_noxref_d )  \
 PM_DFFRNQNX1\%GND
x_PM_DFFRNQNX1\%VDD ( VDD N_VDD_c_301_p N_VDD_c_293_n N_VDD_c_405_p \
 N_VDD_c_396_p N_VDD_c_319_p N_VDD_c_375_p N_VDD_c_376_p N_VDD_c_302_p \
 N_VDD_c_303_p N_VDD_c_309_p N_VDD_c_313_p N_VDD_c_379_p N_VDD_c_317_p \
 N_VDD_c_345_p N_VDD_c_381_p N_VDD_c_382_p N_VDD_c_357_p N_VDD_c_400_p \
 N_VDD_c_460_p N_VDD_c_516_p N_VDD_c_517_p N_VDD_c_429_p N_VDD_c_464_p \
 N_VDD_c_477_p N_VDD_c_481_p N_VDD_c_520_p N_VDD_c_484_p N_VDD_c_560_p \
 N_VDD_c_294_n N_VDD_c_295_n N_VDD_c_296_n N_VDD_c_297_n N_VDD_c_298_n \
 N_VDD_c_299_n N_VDD_M16_noxref_s N_VDD_M17_noxref_d N_VDD_M19_noxref_d \
 N_VDD_M21_noxref_d N_VDD_M22_noxref_s N_VDD_M23_noxref_d N_VDD_M25_noxref_d \
 N_VDD_M27_noxref_d N_VDD_M28_noxref_s N_VDD_M29_noxref_d N_VDD_M31_noxref_d \
 N_VDD_M32_noxref_s N_VDD_M33_noxref_d N_VDD_M35_noxref_d N_VDD_M37_noxref_d \
 N_VDD_M38_noxref_s N_VDD_M39_noxref_d N_VDD_M41_noxref_d N_VDD_M43_noxref_d \
 N_VDD_M44_noxref_s N_VDD_M45_noxref_d N_VDD_M47_noxref_d )  PM_DFFRNQNX1\%VDD
x_PM_DFFRNQNX1\%noxref_3 ( N_noxref_3_c_616_n N_noxref_3_c_620_n \
 N_noxref_3_c_621_n N_noxref_3_c_719_p N_noxref_3_c_622_n N_noxref_3_c_637_n \
 N_noxref_3_c_641_n N_noxref_3_c_643_n N_noxref_3_c_647_n N_noxref_3_c_623_n \
 N_noxref_3_c_757_p N_noxref_3_c_651_n N_noxref_3_c_624_n N_noxref_3_c_836_p \
 N_noxref_3_c_767_p N_noxref_3_M2_noxref_g N_noxref_3_M6_noxref_g \
 N_noxref_3_M20_noxref_g N_noxref_3_M21_noxref_g N_noxref_3_M28_noxref_g \
 N_noxref_3_M29_noxref_g N_noxref_3_c_705_p N_noxref_3_c_706_p \
 N_noxref_3_c_707_p N_noxref_3_c_747_p N_noxref_3_c_727_p N_noxref_3_c_749_p \
 N_noxref_3_c_728_p N_noxref_3_c_625_n N_noxref_3_c_627_n N_noxref_3_c_628_n \
 N_noxref_3_c_629_n N_noxref_3_c_630_n N_noxref_3_c_631_n N_noxref_3_c_632_n \
 N_noxref_3_c_634_n N_noxref_3_c_700_p N_noxref_3_c_710_p N_noxref_3_c_695_p \
 N_noxref_3_c_663_n N_noxref_3_M5_noxref_d N_noxref_3_M22_noxref_d \
 N_noxref_3_M24_noxref_d N_noxref_3_M26_noxref_d )  PM_DFFRNQNX1\%noxref_3
x_PM_DFFRNQNX1\%noxref_4 ( N_noxref_4_c_862_n N_noxref_4_c_910_n \
 N_noxref_4_c_879_n N_noxref_4_c_883_n N_noxref_4_c_885_n N_noxref_4_c_863_n \
 N_noxref_4_c_951_p N_noxref_4_c_864_n N_noxref_4_c_865_n N_noxref_4_c_978_p \
 N_noxref_4_M8_noxref_g N_noxref_4_M32_noxref_g N_noxref_4_M33_noxref_g \
 N_noxref_4_c_866_n N_noxref_4_c_868_n N_noxref_4_c_869_n N_noxref_4_c_870_n \
 N_noxref_4_c_871_n N_noxref_4_c_872_n N_noxref_4_c_873_n N_noxref_4_c_875_n \
 N_noxref_4_c_927_p N_noxref_4_c_897_n N_noxref_4_M7_noxref_d \
 N_noxref_4_M28_noxref_d N_noxref_4_M30_noxref_d )  PM_DFFRNQNX1\%noxref_4
x_PM_DFFRNQNX1\%CLK ( N_CLK_c_1011_n N_CLK_c_1028_n CLK CLK CLK CLK CLK CLK \
 CLK CLK CLK N_CLK_c_1009_n N_CLK_c_1010_n N_CLK_M1_noxref_g N_CLK_M9_noxref_g \
 N_CLK_M18_noxref_g N_CLK_M19_noxref_g N_CLK_M34_noxref_g N_CLK_M35_noxref_g \
 N_CLK_c_1163_p N_CLK_c_1165_p N_CLK_c_1189_p N_CLK_c_1196_p N_CLK_c_1059_n \
 N_CLK_c_1060_n N_CLK_c_1061_n N_CLK_c_1062_n N_CLK_c_1065_n N_CLK_c_1082_n \
 N_CLK_c_1085_n N_CLK_c_1212_p N_CLK_c_1219_p N_CLK_c_1087_n N_CLK_c_1088_n \
 N_CLK_c_1089_n N_CLK_c_1090_n N_CLK_c_1134_p N_CLK_c_1066_n N_CLK_c_1092_n )  \
 PM_DFFRNQNX1\%CLK
x_PM_DFFRNQNX1\%noxref_6 ( N_noxref_6_c_1297_n N_noxref_6_c_1298_n \
 N_noxref_6_c_1224_n N_noxref_6_c_1305_n N_noxref_6_c_1249_n \
 N_noxref_6_c_1253_n N_noxref_6_c_1255_n N_noxref_6_c_1259_n \
 N_noxref_6_c_1225_n N_noxref_6_c_1312_n N_noxref_6_c_1263_n \
 N_noxref_6_c_1226_n N_noxref_6_c_1227_n N_noxref_6_c_1355_n \
 N_noxref_6_c_1321_n N_noxref_6_M3_noxref_g N_noxref_6_M11_noxref_g \
 N_noxref_6_M22_noxref_g N_noxref_6_M23_noxref_g N_noxref_6_M38_noxref_g \
 N_noxref_6_M39_noxref_g N_noxref_6_c_1228_n N_noxref_6_c_1230_n \
 N_noxref_6_c_1231_n N_noxref_6_c_1232_n N_noxref_6_c_1233_n \
 N_noxref_6_c_1234_n N_noxref_6_c_1235_n N_noxref_6_c_1237_n \
 N_noxref_6_c_1326_n N_noxref_6_c_1278_n N_noxref_6_c_1238_n \
 N_noxref_6_c_1240_n N_noxref_6_c_1241_n N_noxref_6_c_1242_n \
 N_noxref_6_c_1243_n N_noxref_6_c_1244_n N_noxref_6_c_1245_n \
 N_noxref_6_c_1247_n N_noxref_6_c_1373_p N_noxref_6_c_1280_n \
 N_noxref_6_M2_noxref_d N_noxref_6_M16_noxref_d N_noxref_6_M18_noxref_d \
 N_noxref_6_M20_noxref_d )  PM_DFFRNQNX1\%noxref_6
x_PM_DFFRNQNX1\%RN ( N_RN_c_1470_n N_RN_c_1478_n N_RN_c_1480_n N_RN_c_1484_n \
 RN RN RN RN RN RN RN RN RN RN RN RN RN RN N_RN_c_1485_n N_RN_c_1486_n \
 N_RN_c_1487_n N_RN_M5_noxref_g N_RN_M10_noxref_g N_RN_M12_noxref_g \
 N_RN_M26_noxref_g N_RN_M27_noxref_g N_RN_M36_noxref_g N_RN_M37_noxref_g \
 N_RN_M40_noxref_g N_RN_M41_noxref_g N_RN_c_1522_n N_RN_c_1523_n N_RN_c_1524_n \
 N_RN_c_1525_n N_RN_c_1526_n N_RN_c_1528_n N_RN_c_1529_n N_RN_c_1556_n \
 N_RN_c_1557_n N_RN_c_1558_n N_RN_c_1640_p N_RN_c_1623_p N_RN_c_1642_p \
 N_RN_c_1624_p N_RN_c_1584_n N_RN_c_1587_n N_RN_c_1727_p N_RN_c_1734_p \
 N_RN_c_1589_n N_RN_c_1590_n N_RN_c_1591_n N_RN_c_1592_n N_RN_c_1602_p \
 N_RN_c_1531_n N_RN_c_1532_n N_RN_c_1534_n N_RN_c_1560_n N_RN_c_1562_n \
 N_RN_c_1563_n N_RN_c_1594_n )  PM_DFFRNQNX1\%RN
x_PM_DFFRNQNX1\%QN ( N_QN_c_1739_n N_QN_c_1743_n QN QN QN QN QN QN QN QN QN QN \
 QN N_QN_c_1758_n N_QN_c_1762_n N_QN_c_1764_n N_QN_c_1768_n N_QN_c_1744_n \
 N_QN_c_1842_p N_QN_c_1745_n N_QN_c_1804_n N_QN_c_1848_p N_QN_M14_noxref_g \
 N_QN_M44_noxref_g N_QN_M45_noxref_g N_QN_c_1746_n N_QN_c_1748_n N_QN_c_1749_n \
 N_QN_c_1750_n N_QN_c_1751_n N_QN_c_1752_n N_QN_c_1753_n N_QN_c_1755_n \
 N_QN_c_1779_n N_QN_M13_noxref_d N_QN_M38_noxref_d N_QN_M40_noxref_d \
 N_QN_M42_noxref_d )  PM_DFFRNQNX1\%QN
x_PM_DFFRNQNX1\%noxref_9 ( N_noxref_9_c_1895_n N_noxref_9_c_1896_n \
 N_noxref_9_c_1922_n N_noxref_9_c_1998_n N_noxref_9_c_1897_n \
 N_noxref_9_c_1935_n N_noxref_9_c_1898_n N_noxref_9_c_2000_n \
 N_noxref_9_c_1899_n N_noxref_9_c_1943_n N_noxref_9_c_1947_n \
 N_noxref_9_c_1949_n N_noxref_9_c_1953_n N_noxref_9_c_1901_n \
 N_noxref_9_c_2144_n N_noxref_9_c_1957_n N_noxref_9_c_2175_n \
 N_noxref_9_c_1902_n N_noxref_9_c_2080_n N_noxref_9_c_2152_n \
 N_noxref_9_M0_noxref_g N_noxref_9_M7_noxref_g N_noxref_9_M15_noxref_g \
 N_noxref_9_M16_noxref_g N_noxref_9_M17_noxref_g N_noxref_9_M30_noxref_g \
 N_noxref_9_M31_noxref_g N_noxref_9_M46_noxref_g N_noxref_9_M47_noxref_g \
 N_noxref_9_c_1904_n N_noxref_9_c_1906_n N_noxref_9_c_1907_n \
 N_noxref_9_c_1908_n N_noxref_9_c_1909_n N_noxref_9_c_1910_n \
 N_noxref_9_c_1911_n N_noxref_9_c_1913_n N_noxref_9_c_2095_n \
 N_noxref_9_c_1974_n N_noxref_9_c_2009_n N_noxref_9_c_2012_n \
 N_noxref_9_c_2014_n N_noxref_9_c_2044_n N_noxref_9_c_2046_n \
 N_noxref_9_c_2047_n N_noxref_9_c_2017_n N_noxref_9_c_2018_n \
 N_noxref_9_c_2184_n N_noxref_9_c_2187_n N_noxref_9_c_2189_n \
 N_noxref_9_c_2200_p N_noxref_9_c_2224_p N_noxref_9_c_2210_p \
 N_noxref_9_c_2192_n N_noxref_9_c_2193_n N_noxref_9_c_2019_n \
 N_noxref_9_c_2053_n N_noxref_9_c_2021_n N_noxref_9_c_2194_n \
 N_noxref_9_c_2217_p N_noxref_9_c_2196_n N_noxref_9_M10_noxref_d \
 N_noxref_9_M32_noxref_d N_noxref_9_M34_noxref_d N_noxref_9_M36_noxref_d )  \
 PM_DFFRNQNX1\%noxref_9
x_PM_DFFRNQNX1\%noxref_10 ( N_noxref_10_c_2279_n N_noxref_10_c_2280_n \
 N_noxref_10_c_2281_n N_noxref_10_c_2290_n N_noxref_10_c_2294_n \
 N_noxref_10_c_2296_n N_noxref_10_c_2282_n N_noxref_10_c_2413_p \
 N_noxref_10_c_2283_n N_noxref_10_c_2392_n N_noxref_10_M13_noxref_g \
 N_noxref_10_M42_noxref_g N_noxref_10_M43_noxref_g N_noxref_10_c_2325_n \
 N_noxref_10_c_2326_n N_noxref_10_c_2327_n N_noxref_10_c_2358_n \
 N_noxref_10_c_2359_n N_noxref_10_c_2361_n N_noxref_10_c_2362_n \
 N_noxref_10_c_2328_n N_noxref_10_c_2331_n N_noxref_10_c_2332_n \
 N_noxref_10_M15_noxref_d N_noxref_10_M44_noxref_d N_noxref_10_M46_noxref_d )  \
 PM_DFFRNQNX1\%noxref_10
x_PM_DFFRNQNX1\%noxref_11 ( N_noxref_11_c_2448_n N_noxref_11_c_2423_n \
 N_noxref_11_c_2427_n N_noxref_11_c_2430_n N_noxref_11_c_2441_n \
 N_noxref_11_M0_noxref_s )  PM_DFFRNQNX1\%noxref_11
x_PM_DFFRNQNX1\%noxref_12 ( N_noxref_12_c_2470_n N_noxref_12_c_2472_n \
 N_noxref_12_c_2475_n N_noxref_12_c_2478_n N_noxref_12_c_2489_n \
 N_noxref_12_M1_noxref_d N_noxref_12_M2_noxref_s )  PM_DFFRNQNX1\%noxref_12
x_PM_DFFRNQNX1\%D ( D D N_D_c_2523_n N_D_M4_noxref_g N_D_M24_noxref_g \
 N_D_M25_noxref_g N_D_c_2552_n N_D_c_2555_n N_D_c_2591_p N_D_c_2598_p \
 N_D_c_2557_n N_D_c_2558_n N_D_c_2559_n N_D_c_2560_n N_D_c_2537_n N_D_c_2538_n \
 )  PM_DFFRNQNX1\%D
x_PM_DFFRNQNX1\%noxref_14 ( N_noxref_14_c_2619_n N_noxref_14_c_2603_n \
 N_noxref_14_c_2607_n N_noxref_14_c_2610_n N_noxref_14_c_2621_n \
 N_noxref_14_M3_noxref_s )  PM_DFFRNQNX1\%noxref_14
x_PM_DFFRNQNX1\%noxref_15 ( N_noxref_15_c_2653_n N_noxref_15_c_2655_n \
 N_noxref_15_c_2658_n N_noxref_15_c_2661_n N_noxref_15_c_2670_n \
 N_noxref_15_M4_noxref_d N_noxref_15_M5_noxref_s )  PM_DFFRNQNX1\%noxref_15
x_PM_DFFRNQNX1\%noxref_16 ( N_noxref_16_c_2726_n N_noxref_16_c_2707_n \
 N_noxref_16_c_2711_n N_noxref_16_c_2714_n N_noxref_16_c_2715_n \
 N_noxref_16_c_2718_n N_noxref_16_M6_noxref_s )  PM_DFFRNQNX1\%noxref_16
x_PM_DFFRNQNX1\%noxref_17 ( N_noxref_17_c_2775_n N_noxref_17_c_2759_n \
 N_noxref_17_c_2763_n N_noxref_17_c_2766_n N_noxref_17_c_2789_n \
 N_noxref_17_M8_noxref_s )  PM_DFFRNQNX1\%noxref_17
x_PM_DFFRNQNX1\%noxref_18 ( N_noxref_18_c_2809_n N_noxref_18_c_2811_n \
 N_noxref_18_c_2814_n N_noxref_18_c_2817_n N_noxref_18_c_2842_n \
 N_noxref_18_M9_noxref_d N_noxref_18_M10_noxref_s )  PM_DFFRNQNX1\%noxref_18
x_PM_DFFRNQNX1\%noxref_19 ( N_noxref_19_c_2879_n N_noxref_19_c_2863_n \
 N_noxref_19_c_2867_n N_noxref_19_c_2870_n N_noxref_19_c_2893_n \
 N_noxref_19_M11_noxref_s )  PM_DFFRNQNX1\%noxref_19
x_PM_DFFRNQNX1\%noxref_20 ( N_noxref_20_c_2915_n N_noxref_20_c_2917_n \
 N_noxref_20_c_2920_n N_noxref_20_c_2923_n N_noxref_20_c_2943_n \
 N_noxref_20_M12_noxref_d N_noxref_20_M13_noxref_s )  PM_DFFRNQNX1\%noxref_20
x_PM_DFFRNQNX1\%noxref_21 ( N_noxref_21_c_2984_n N_noxref_21_c_2967_n \
 N_noxref_21_c_2971_n N_noxref_21_c_2974_n N_noxref_21_c_2975_n \
 N_noxref_21_c_2977_n N_noxref_21_M14_noxref_s )  PM_DFFRNQNX1\%noxref_21
cc_1 ( N_GND_c_1_p N_VDD_c_293_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_294_n ) capacitor c=0.00989031f //x=25.53 //y=0 \
 //x2=25.53 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_295_n ) capacitor c=0.00500587f //x=4.81 //y=0 \
 //x2=4.81 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_296_n ) capacitor c=0.00500587f //x=9.62 //y=0 \
 //x2=9.62 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_297_n ) capacitor c=0.00500587f //x=12.95 //y=0 \
 //x2=12.95 //y2=7.4
cc_6 ( N_GND_c_6_p N_VDD_c_298_n ) capacitor c=0.00524516f //x=17.76 //y=0 \
 //x2=17.76 //y2=7.4
cc_7 ( N_GND_c_7_p N_VDD_c_299_n ) capacitor c=0.00500587f //x=22.57 //y=0 \
 //x2=22.57 //y2=7.4
cc_8 ( N_GND_c_8_p N_noxref_3_c_616_n ) capacitor c=0.0324991f //x=25.53 //y=0 \
 //x2=8.765 //y2=3.33
cc_9 ( N_GND_c_9_p N_noxref_3_c_616_n ) capacitor c=0.00174514f //x=4.64 //y=0 \
 //x2=8.765 //y2=3.33
cc_10 ( N_GND_c_10_p N_noxref_3_c_616_n ) capacitor c=0.00152503f //x=5.8 \
 //y=0 //x2=8.765 //y2=3.33
cc_11 ( N_GND_c_3_p N_noxref_3_c_616_n ) capacitor c=0.00820844f //x=4.81 \
 //y=0 //x2=8.765 //y2=3.33
cc_12 ( N_GND_c_8_p N_noxref_3_c_620_n ) capacitor c=0.00172266f //x=25.53 \
 //y=0 //x2=3.445 //y2=3.33
cc_13 ( N_GND_c_4_p N_noxref_3_c_621_n ) capacitor c=0.00582294f //x=9.62 \
 //y=0 //x2=10.615 //y2=3.33
cc_14 ( N_GND_c_3_p N_noxref_3_c_622_n ) capacitor c=9.53263e-19 //x=4.81 \
 //y=0 //x2=3.33 //y2=2.08
cc_15 ( N_GND_c_4_p N_noxref_3_c_623_n ) capacitor c=0.0432238f //x=9.62 //y=0 \
 //x2=8.795 //y2=1.665
cc_16 ( N_GND_c_4_p N_noxref_3_c_624_n ) capacitor c=0.0156446f //x=9.62 //y=0 \
 //x2=10.73 //y2=2.08
cc_17 ( N_GND_c_17_p N_noxref_3_c_625_n ) capacitor c=0.00135046f //x=10.715 \
 //y=0 //x2=10.535 //y2=0.865
cc_18 ( N_GND_M6_noxref_d N_noxref_3_c_625_n ) capacitor c=0.00220047f \
 //x=10.61 //y=0.865 //x2=10.535 //y2=0.865
cc_19 ( N_GND_M6_noxref_d N_noxref_3_c_627_n ) capacitor c=0.00255985f \
 //x=10.61 //y=0.865 //x2=10.535 //y2=1.21
cc_20 ( N_GND_c_4_p N_noxref_3_c_628_n ) capacitor c=0.00189421f //x=9.62 \
 //y=0 //x2=10.535 //y2=1.52
cc_21 ( N_GND_c_4_p N_noxref_3_c_629_n ) capacitor c=0.00992619f //x=9.62 \
 //y=0 //x2=10.535 //y2=1.915
cc_22 ( N_GND_M6_noxref_d N_noxref_3_c_630_n ) capacitor c=0.0131326f \
 //x=10.61 //y=0.865 //x2=10.91 //y2=0.71
cc_23 ( N_GND_M6_noxref_d N_noxref_3_c_631_n ) capacitor c=0.00193127f \
 //x=10.61 //y=0.865 //x2=10.91 //y2=1.365
cc_24 ( N_GND_c_24_p N_noxref_3_c_632_n ) capacitor c=0.00130622f //x=12.78 \
 //y=0 //x2=11.065 //y2=0.865
cc_25 ( N_GND_M6_noxref_d N_noxref_3_c_632_n ) capacitor c=0.00257848f \
 //x=10.61 //y=0.865 //x2=11.065 //y2=0.865
cc_26 ( N_GND_M6_noxref_d N_noxref_3_c_634_n ) capacitor c=0.00255985f \
 //x=10.61 //y=0.865 //x2=11.065 //y2=1.21
cc_27 ( N_GND_c_4_p N_noxref_3_M5_noxref_d ) capacitor c=0.00591582f //x=9.62 \
 //y=0 //x2=8.205 //y2=0.915
cc_28 ( N_GND_c_5_p N_noxref_4_c_862_n ) capacitor c=0.00582294f //x=12.95 \
 //y=0 //x2=13.945 //y2=3.33
cc_29 ( N_GND_c_5_p N_noxref_4_c_863_n ) capacitor c=0.0436242f //x=12.95 \
 //y=0 //x2=12.125 //y2=1.655
cc_30 ( N_GND_c_4_p N_noxref_4_c_864_n ) capacitor c=9.64732e-19 //x=9.62 \
 //y=0 //x2=12.21 //y2=3.33
cc_31 ( N_GND_c_5_p N_noxref_4_c_865_n ) capacitor c=0.0156442f //x=12.95 \
 //y=0 //x2=14.06 //y2=2.08
cc_32 ( N_GND_c_32_p N_noxref_4_c_866_n ) capacitor c=0.00132755f //x=13.94 \
 //y=0 //x2=13.76 //y2=0.875
cc_33 ( N_GND_M8_noxref_d N_noxref_4_c_866_n ) capacitor c=0.00211996f \
 //x=13.835 //y=0.875 //x2=13.76 //y2=0.875
cc_34 ( N_GND_M8_noxref_d N_noxref_4_c_868_n ) capacitor c=0.00255985f \
 //x=13.835 //y=0.875 //x2=13.76 //y2=1.22
cc_35 ( N_GND_c_5_p N_noxref_4_c_869_n ) capacitor c=0.00195164f //x=12.95 \
 //y=0 //x2=13.76 //y2=1.53
cc_36 ( N_GND_c_5_p N_noxref_4_c_870_n ) capacitor c=0.0110952f //x=12.95 \
 //y=0 //x2=13.76 //y2=1.915
cc_37 ( N_GND_M8_noxref_d N_noxref_4_c_871_n ) capacitor c=0.0131341f \
 //x=13.835 //y=0.875 //x2=14.135 //y2=0.72
cc_38 ( N_GND_M8_noxref_d N_noxref_4_c_872_n ) capacitor c=0.00193146f \
 //x=13.835 //y=0.875 //x2=14.135 //y2=1.375
cc_39 ( N_GND_c_39_p N_noxref_4_c_873_n ) capacitor c=0.00129018f //x=17.59 \
 //y=0 //x2=14.29 //y2=0.875
cc_40 ( N_GND_M8_noxref_d N_noxref_4_c_873_n ) capacitor c=0.00257848f \
 //x=13.835 //y=0.875 //x2=14.29 //y2=0.875
cc_41 ( N_GND_M8_noxref_d N_noxref_4_c_875_n ) capacitor c=0.00255985f \
 //x=13.835 //y=0.875 //x2=14.29 //y2=1.22
cc_42 ( N_GND_c_4_p N_noxref_4_M7_noxref_d ) capacitor c=8.58106e-19 //x=9.62 \
 //y=0 //x2=11.58 //y2=0.905
cc_43 ( N_GND_c_5_p N_noxref_4_M7_noxref_d ) capacitor c=0.00616547f //x=12.95 \
 //y=0 //x2=11.58 //y2=0.905
cc_44 ( N_GND_M6_noxref_d N_noxref_4_M7_noxref_d ) capacitor c=0.00143464f \
 //x=10.61 //y=0.865 //x2=11.58 //y2=0.905
cc_45 ( N_GND_c_1_p N_CLK_c_1009_n ) capacitor c=7.64246e-19 //x=0.74 //y=0 \
 //x2=2.22 //y2=2.08
cc_46 ( N_GND_c_5_p N_CLK_c_1010_n ) capacitor c=6.04789e-19 //x=12.95 //y=0 \
 //x2=15.17 //y2=2.08
cc_47 ( N_GND_c_6_p N_noxref_6_c_1224_n ) capacitor c=0.00390249f //x=17.76 \
 //y=0 //x2=18.755 //y2=3.7
cc_48 ( N_GND_c_3_p N_noxref_6_c_1225_n ) capacitor c=0.0459494f //x=4.81 \
 //y=0 //x2=3.985 //y2=1.665
cc_49 ( N_GND_c_3_p N_noxref_6_c_1226_n ) capacitor c=0.0178133f //x=4.81 \
 //y=0 //x2=5.92 //y2=2.08
cc_50 ( N_GND_c_6_p N_noxref_6_c_1227_n ) capacitor c=0.0155796f //x=17.76 \
 //y=0 //x2=18.87 //y2=2.08
cc_51 ( N_GND_c_10_p N_noxref_6_c_1228_n ) capacitor c=0.00132755f //x=5.8 \
 //y=0 //x2=5.62 //y2=0.875
cc_52 ( N_GND_M3_noxref_d N_noxref_6_c_1228_n ) capacitor c=0.00211996f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=0.875
cc_53 ( N_GND_M3_noxref_d N_noxref_6_c_1230_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=1.22
cc_54 ( N_GND_c_3_p N_noxref_6_c_1231_n ) capacitor c=0.00204716f //x=4.81 \
 //y=0 //x2=5.62 //y2=1.53
cc_55 ( N_GND_c_3_p N_noxref_6_c_1232_n ) capacitor c=0.0118433f //x=4.81 \
 //y=0 //x2=5.62 //y2=1.915
cc_56 ( N_GND_M3_noxref_d N_noxref_6_c_1233_n ) capacitor c=0.0131341f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=0.72
cc_57 ( N_GND_M3_noxref_d N_noxref_6_c_1234_n ) capacitor c=0.00193146f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=1.375
cc_58 ( N_GND_c_58_p N_noxref_6_c_1235_n ) capacitor c=0.00129018f //x=9.45 \
 //y=0 //x2=6.15 //y2=0.875
cc_59 ( N_GND_M3_noxref_d N_noxref_6_c_1235_n ) capacitor c=0.00257848f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=0.875
cc_60 ( N_GND_M3_noxref_d N_noxref_6_c_1237_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=1.22
cc_61 ( N_GND_c_61_p N_noxref_6_c_1238_n ) capacitor c=0.00132755f //x=18.75 \
 //y=0 //x2=18.57 //y2=0.875
cc_62 ( N_GND_M11_noxref_d N_noxref_6_c_1238_n ) capacitor c=0.00211996f \
 //x=18.645 //y=0.875 //x2=18.57 //y2=0.875
cc_63 ( N_GND_M11_noxref_d N_noxref_6_c_1240_n ) capacitor c=0.00255985f \
 //x=18.645 //y=0.875 //x2=18.57 //y2=1.22
cc_64 ( N_GND_c_6_p N_noxref_6_c_1241_n ) capacitor c=0.00204716f //x=17.76 \
 //y=0 //x2=18.57 //y2=1.53
cc_65 ( N_GND_c_6_p N_noxref_6_c_1242_n ) capacitor c=0.0110952f //x=17.76 \
 //y=0 //x2=18.57 //y2=1.915
cc_66 ( N_GND_M11_noxref_d N_noxref_6_c_1243_n ) capacitor c=0.0131341f \
 //x=18.645 //y=0.875 //x2=18.945 //y2=0.72
cc_67 ( N_GND_M11_noxref_d N_noxref_6_c_1244_n ) capacitor c=0.00193146f \
 //x=18.645 //y=0.875 //x2=18.945 //y2=1.375
cc_68 ( N_GND_c_68_p N_noxref_6_c_1245_n ) capacitor c=0.00129018f //x=22.4 \
 //y=0 //x2=19.1 //y2=0.875
cc_69 ( N_GND_M11_noxref_d N_noxref_6_c_1245_n ) capacitor c=0.00257848f \
 //x=18.645 //y=0.875 //x2=19.1 //y2=0.875
cc_70 ( N_GND_M11_noxref_d N_noxref_6_c_1247_n ) capacitor c=0.00255985f \
 //x=18.645 //y=0.875 //x2=19.1 //y2=1.22
cc_71 ( N_GND_c_3_p N_noxref_6_M2_noxref_d ) capacitor c=0.00591582f //x=4.81 \
 //y=0 //x2=3.395 //y2=0.915
cc_72 ( N_GND_c_8_p N_RN_c_1470_n ) capacitor c=0.0754427f //x=25.53 //y=0 \
 //x2=16.165 //y2=2.22
cc_73 ( N_GND_c_58_p N_RN_c_1470_n ) capacitor c=0.00318526f //x=9.45 //y=0 \
 //x2=16.165 //y2=2.22
cc_74 ( N_GND_c_17_p N_RN_c_1470_n ) capacitor c=0.00347653f //x=10.715 //y=0 \
 //x2=16.165 //y2=2.22
cc_75 ( N_GND_c_24_p N_RN_c_1470_n ) capacitor c=0.00411932f //x=12.78 //y=0 \
 //x2=16.165 //y2=2.22
cc_76 ( N_GND_c_32_p N_RN_c_1470_n ) capacitor c=0.00274252f //x=13.94 //y=0 \
 //x2=16.165 //y2=2.22
cc_77 ( N_GND_c_39_p N_RN_c_1470_n ) capacitor c=0.00111309f //x=17.59 //y=0 \
 //x2=16.165 //y2=2.22
cc_78 ( N_GND_c_4_p N_RN_c_1470_n ) capacitor c=0.0418918f //x=9.62 //y=0 \
 //x2=16.165 //y2=2.22
cc_79 ( N_GND_c_5_p N_RN_c_1470_n ) capacitor c=0.0418918f //x=12.95 //y=0 \
 //x2=16.165 //y2=2.22
cc_80 ( N_GND_c_8_p N_RN_c_1478_n ) capacitor c=0.00221055f //x=25.53 //y=0 \
 //x2=8.255 //y2=2.22
cc_81 ( N_GND_c_58_p N_RN_c_1478_n ) capacitor c=4.19033e-19 //x=9.45 //y=0 \
 //x2=8.255 //y2=2.22
cc_82 ( N_GND_c_8_p N_RN_c_1480_n ) capacitor c=0.0355717f //x=25.53 //y=0 \
 //x2=19.865 //y2=2.22
cc_83 ( N_GND_c_39_p N_RN_c_1480_n ) capacitor c=0.00318526f //x=17.59 //y=0 \
 //x2=19.865 //y2=2.22
cc_84 ( N_GND_c_61_p N_RN_c_1480_n ) capacitor c=0.00274252f //x=18.75 //y=0 \
 //x2=19.865 //y2=2.22
cc_85 ( N_GND_c_6_p N_RN_c_1480_n ) capacitor c=0.0430854f //x=17.76 //y=0 \
 //x2=19.865 //y2=2.22
cc_86 ( N_GND_c_8_p N_RN_c_1484_n ) capacitor c=0.00195247f //x=25.53 //y=0 \
 //x2=16.395 //y2=2.22
cc_87 ( N_GND_c_4_p N_RN_c_1485_n ) capacitor c=8.37259e-19 //x=9.62 //y=0 \
 //x2=8.14 //y2=2.08
cc_88 ( N_GND_c_6_p N_RN_c_1486_n ) capacitor c=8.37259e-19 //x=17.76 //y=0 \
 //x2=16.28 //y2=2.08
cc_89 ( N_GND_c_6_p N_RN_c_1487_n ) capacitor c=5.94159e-19 //x=17.76 //y=0 \
 //x2=19.98 //y2=2.08
cc_90 ( N_GND_c_8_p N_QN_c_1739_n ) capacitor c=0.0143872f //x=25.53 //y=0 \
 //x2=23.565 //y2=3.33
cc_91 ( N_GND_c_68_p N_QN_c_1739_n ) capacitor c=0.0016229f //x=22.4 //y=0 \
 //x2=23.565 //y2=3.33
cc_92 ( N_GND_c_92_p N_QN_c_1739_n ) capacitor c=0.00189853f //x=23.665 //y=0 \
 //x2=23.565 //y2=3.33
cc_93 ( N_GND_c_7_p N_QN_c_1739_n ) capacitor c=0.00820844f //x=22.57 //y=0 \
 //x2=23.565 //y2=3.33
cc_94 ( N_GND_c_8_p N_QN_c_1743_n ) capacitor c=0.0017709f //x=25.53 //y=0 \
 //x2=21.945 //y2=3.33
cc_95 ( N_GND_c_7_p N_QN_c_1744_n ) capacitor c=0.0455978f //x=22.57 //y=0 \
 //x2=21.745 //y2=1.665
cc_96 ( N_GND_c_7_p N_QN_c_1745_n ) capacitor c=0.0179404f //x=22.57 //y=0 \
 //x2=23.68 //y2=2.08
cc_97 ( N_GND_c_92_p N_QN_c_1746_n ) capacitor c=0.00135046f //x=23.665 //y=0 \
 //x2=23.485 //y2=0.865
cc_98 ( N_GND_M14_noxref_d N_QN_c_1746_n ) capacitor c=0.00220047f //x=23.56 \
 //y=0.865 //x2=23.485 //y2=0.865
cc_99 ( N_GND_M14_noxref_d N_QN_c_1748_n ) capacitor c=0.00255985f //x=23.56 \
 //y=0.865 //x2=23.485 //y2=1.21
cc_100 ( N_GND_c_7_p N_QN_c_1749_n ) capacitor c=0.00189421f //x=22.57 //y=0 \
 //x2=23.485 //y2=1.52
cc_101 ( N_GND_c_7_p N_QN_c_1750_n ) capacitor c=0.0106743f //x=22.57 //y=0 \
 //x2=23.485 //y2=1.915
cc_102 ( N_GND_M14_noxref_d N_QN_c_1751_n ) capacitor c=0.0131326f //x=23.56 \
 //y=0.865 //x2=23.86 //y2=0.71
cc_103 ( N_GND_M14_noxref_d N_QN_c_1752_n ) capacitor c=0.00193127f //x=23.56 \
 //y=0.865 //x2=23.86 //y2=1.365
cc_104 ( N_GND_c_2_p N_QN_c_1753_n ) capacitor c=0.00130622f //x=25.53 //y=0 \
 //x2=24.015 //y2=0.865
cc_105 ( N_GND_M14_noxref_d N_QN_c_1753_n ) capacitor c=0.00257848f //x=23.56 \
 //y=0.865 //x2=24.015 //y2=0.865
cc_106 ( N_GND_M14_noxref_d N_QN_c_1755_n ) capacitor c=0.00255985f //x=23.56 \
 //y=0.865 //x2=24.015 //y2=1.21
cc_107 ( N_GND_c_7_p N_QN_M13_noxref_d ) capacitor c=0.00591582f //x=22.57 \
 //y=0 //x2=21.155 //y2=0.915
cc_108 ( N_GND_c_8_p N_noxref_9_c_1895_n ) capacitor c=0.0122686f //x=25.53 \
 //y=0 //x2=11.355 //y2=4.07
cc_109 ( N_GND_c_8_p N_noxref_9_c_1896_n ) capacitor c=0.0015877f //x=25.53 \
 //y=0 //x2=1.225 //y2=4.07
cc_110 ( N_GND_c_8_p N_noxref_9_c_1897_n ) capacitor c=0.010852f //x=25.53 \
 //y=0 //x2=24.305 //y2=4.07
cc_111 ( N_GND_c_1_p N_noxref_9_c_1898_n ) capacitor c=0.0180363f //x=0.74 \
 //y=0 //x2=1.11 //y2=2.08
cc_112 ( N_GND_c_4_p N_noxref_9_c_1899_n ) capacitor c=7.4738e-19 //x=9.62 \
 //y=0 //x2=11.47 //y2=2.08
cc_113 ( N_GND_c_5_p N_noxref_9_c_1899_n ) capacitor c=7.76678e-19 //x=12.95 \
 //y=0 //x2=11.47 //y2=2.08
cc_114 ( N_GND_c_6_p N_noxref_9_c_1901_n ) capacitor c=0.0430857f //x=17.76 \
 //y=0 //x2=16.935 //y2=1.665
cc_115 ( N_GND_c_2_p N_noxref_9_c_1902_n ) capacitor c=9.53263e-19 //x=25.53 \
 //y=0 //x2=24.42 //y2=2.08
cc_116 ( N_GND_c_7_p N_noxref_9_c_1902_n ) capacitor c=9.2064e-19 //x=22.57 \
 //y=0 //x2=24.42 //y2=2.08
cc_117 ( N_GND_c_117_p N_noxref_9_c_1904_n ) capacitor c=0.00132755f //x=0.99 \
 //y=0 //x2=0.81 //y2=0.875
cc_118 ( N_GND_M0_noxref_d N_noxref_9_c_1904_n ) capacitor c=0.00211996f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=0.875
cc_119 ( N_GND_M0_noxref_d N_noxref_9_c_1906_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=1.22
cc_120 ( N_GND_c_1_p N_noxref_9_c_1907_n ) capacitor c=0.00295461f //x=0.74 \
 //y=0 //x2=0.81 //y2=1.53
cc_121 ( N_GND_c_1_p N_noxref_9_c_1908_n ) capacitor c=0.0134214f //x=0.74 \
 //y=0 //x2=0.81 //y2=1.915
cc_122 ( N_GND_M0_noxref_d N_noxref_9_c_1909_n ) capacitor c=0.0131341f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=0.72
cc_123 ( N_GND_M0_noxref_d N_noxref_9_c_1910_n ) capacitor c=0.00193146f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=1.375
cc_124 ( N_GND_c_9_p N_noxref_9_c_1911_n ) capacitor c=0.00129018f //x=4.64 \
 //y=0 //x2=1.34 //y2=0.875
cc_125 ( N_GND_M0_noxref_d N_noxref_9_c_1911_n ) capacitor c=0.00257848f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=0.875
cc_126 ( N_GND_M0_noxref_d N_noxref_9_c_1913_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=1.22
cc_127 ( N_GND_c_6_p N_noxref_9_M10_noxref_d ) capacitor c=0.00591582f \
 //x=17.76 //y=0 //x2=16.345 //y2=0.915
cc_128 ( N_GND_c_8_p N_noxref_10_c_2279_n ) capacitor c=0.0185866f //x=25.53 \
 //y=0 //x2=25.045 //y2=3.7
cc_129 ( N_GND_c_8_p N_noxref_10_c_2280_n ) capacitor c=0.00154647f //x=25.53 \
 //y=0 //x2=21.205 //y2=3.7
cc_130 ( N_GND_c_7_p N_noxref_10_c_2281_n ) capacitor c=0.00128267f //x=22.57 \
 //y=0 //x2=21.09 //y2=2.08
cc_131 ( N_GND_c_2_p N_noxref_10_c_2282_n ) capacitor c=0.0468439f //x=25.53 \
 //y=0 //x2=25.075 //y2=1.655
cc_132 ( N_GND_c_7_p N_noxref_10_c_2283_n ) capacitor c=9.64732e-19 //x=22.57 \
 //y=0 //x2=25.16 //y2=3.7
cc_133 ( N_GND_c_2_p N_noxref_10_M15_noxref_d ) capacitor c=0.00618259f \
 //x=25.53 //y=0 //x2=24.53 //y2=0.905
cc_134 ( N_GND_c_7_p N_noxref_10_M15_noxref_d ) capacitor c=8.58106e-19 \
 //x=22.57 //y=0 //x2=24.53 //y2=0.905
cc_135 ( N_GND_M14_noxref_d N_noxref_10_M15_noxref_d ) capacitor c=0.00143464f \
 //x=23.56 //y=0.865 //x2=24.53 //y2=0.905
cc_136 ( N_GND_c_8_p N_noxref_11_c_2423_n ) capacitor c=0.00618812f //x=25.53 \
 //y=0 //x2=1.475 //y2=1.59
cc_137 ( N_GND_c_117_p N_noxref_11_c_2423_n ) capacitor c=0.00110021f //x=0.99 \
 //y=0 //x2=1.475 //y2=1.59
cc_138 ( N_GND_c_9_p N_noxref_11_c_2423_n ) capacitor c=0.00179185f //x=4.64 \
 //y=0 //x2=1.475 //y2=1.59
cc_139 ( N_GND_M0_noxref_d N_noxref_11_c_2423_n ) capacitor c=0.00894788f \
 //x=0.885 //y=0.875 //x2=1.475 //y2=1.59
cc_140 ( N_GND_c_8_p N_noxref_11_c_2427_n ) capacitor c=0.00575184f //x=25.53 \
 //y=0 //x2=1.56 //y2=0.625
cc_141 ( N_GND_c_9_p N_noxref_11_c_2427_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=1.56 //y2=0.625
cc_142 ( N_GND_M0_noxref_d N_noxref_11_c_2427_n ) capacitor c=0.033954f \
 //x=0.885 //y=0.875 //x2=1.56 //y2=0.625
cc_143 ( N_GND_c_8_p N_noxref_11_c_2430_n ) capacitor c=0.0139021f //x=25.53 \
 //y=0 //x2=2.445 //y2=0.54
cc_144 ( N_GND_c_9_p N_noxref_11_c_2430_n ) capacitor c=0.0356078f //x=4.64 \
 //y=0 //x2=2.445 //y2=0.54
cc_145 ( N_GND_c_2_p N_noxref_11_c_2430_n ) capacitor c=0.00177266f //x=25.53 \
 //y=0 //x2=2.445 //y2=0.54
cc_146 ( N_GND_c_8_p N_noxref_11_M0_noxref_s ) capacitor c=0.0125336f \
 //x=25.53 //y=0 //x2=0.455 //y2=0.375
cc_147 ( N_GND_c_117_p N_noxref_11_M0_noxref_s ) capacitor c=0.0140218f \
 //x=0.99 //y=0 //x2=0.455 //y2=0.375
cc_148 ( N_GND_c_1_p N_noxref_11_M0_noxref_s ) capacitor c=0.0712607f //x=0.74 \
 //y=0 //x2=0.455 //y2=0.375
cc_149 ( N_GND_c_9_p N_noxref_11_M0_noxref_s ) capacitor c=0.0131422f //x=4.64 \
 //y=0 //x2=0.455 //y2=0.375
cc_150 ( N_GND_c_3_p N_noxref_11_M0_noxref_s ) capacitor c=3.31601e-19 \
 //x=4.81 //y=0 //x2=0.455 //y2=0.375
cc_151 ( N_GND_M0_noxref_d N_noxref_11_M0_noxref_s ) capacitor c=0.033718f \
 //x=0.885 //y=0.875 //x2=0.455 //y2=0.375
cc_152 ( N_GND_c_8_p N_noxref_12_c_2470_n ) capacitor c=0.00402784f //x=25.53 \
 //y=0 //x2=3.015 //y2=0.995
cc_153 ( N_GND_c_9_p N_noxref_12_c_2470_n ) capacitor c=0.00829979f //x=4.64 \
 //y=0 //x2=3.015 //y2=0.995
cc_154 ( N_GND_c_8_p N_noxref_12_c_2472_n ) capacitor c=0.00575184f //x=25.53 \
 //y=0 //x2=3.1 //y2=0.625
cc_155 ( N_GND_c_9_p N_noxref_12_c_2472_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=3.1 //y2=0.625
cc_156 ( N_GND_M0_noxref_d N_noxref_12_c_2472_n ) capacitor c=6.21394e-19 \
 //x=0.885 //y=0.875 //x2=3.1 //y2=0.625
cc_157 ( N_GND_c_8_p N_noxref_12_c_2475_n ) capacitor c=0.0118365f //x=25.53 \
 //y=0 //x2=3.985 //y2=0.54
cc_158 ( N_GND_c_9_p N_noxref_12_c_2475_n ) capacitor c=0.0365413f //x=4.64 \
 //y=0 //x2=3.985 //y2=0.54
cc_159 ( N_GND_c_2_p N_noxref_12_c_2475_n ) capacitor c=0.00189358f //x=25.53 \
 //y=0 //x2=3.985 //y2=0.54
cc_160 ( N_GND_c_8_p N_noxref_12_c_2478_n ) capacitor c=0.00287549f //x=25.53 \
 //y=0 //x2=4.07 //y2=0.625
cc_161 ( N_GND_c_9_p N_noxref_12_c_2478_n ) capacitor c=0.0142658f //x=4.64 \
 //y=0 //x2=4.07 //y2=0.625
cc_162 ( N_GND_c_3_p N_noxref_12_c_2478_n ) capacitor c=0.0404137f //x=4.81 \
 //y=0 //x2=4.07 //y2=0.625
cc_163 ( N_GND_M0_noxref_d N_noxref_12_M1_noxref_d ) capacitor c=0.00162435f \
 //x=0.885 //y=0.875 //x2=1.86 //y2=0.91
cc_164 ( N_GND_c_1_p N_noxref_12_M2_noxref_s ) capacitor c=8.16352e-19 \
 //x=0.74 //y=0 //x2=2.965 //y2=0.375
cc_165 ( N_GND_c_3_p N_noxref_12_M2_noxref_s ) capacitor c=0.00183204f \
 //x=4.81 //y=0 //x2=2.965 //y2=0.375
cc_166 ( N_GND_c_3_p N_D_c_2523_n ) capacitor c=8.54129e-19 //x=4.81 //y=0 \
 //x2=7.03 //y2=2.08
cc_167 ( N_GND_c_8_p N_noxref_14_c_2603_n ) capacitor c=0.00551063f //x=25.53 \
 //y=0 //x2=6.285 //y2=1.59
cc_168 ( N_GND_c_10_p N_noxref_14_c_2603_n ) capacitor c=0.00111576f //x=5.8 \
 //y=0 //x2=6.285 //y2=1.59
cc_169 ( N_GND_c_58_p N_noxref_14_c_2603_n ) capacitor c=0.0018074f //x=9.45 \
 //y=0 //x2=6.285 //y2=1.59
cc_170 ( N_GND_M3_noxref_d N_noxref_14_c_2603_n ) capacitor c=0.00887549f \
 //x=5.695 //y=0.875 //x2=6.285 //y2=1.59
cc_171 ( N_GND_c_8_p N_noxref_14_c_2607_n ) capacitor c=0.00287639f //x=25.53 \
 //y=0 //x2=6.37 //y2=0.625
cc_172 ( N_GND_c_58_p N_noxref_14_c_2607_n ) capacitor c=0.014327f //x=9.45 \
 //y=0 //x2=6.37 //y2=0.625
cc_173 ( N_GND_M3_noxref_d N_noxref_14_c_2607_n ) capacitor c=0.033954f \
 //x=5.695 //y=0.875 //x2=6.37 //y2=0.625
cc_174 ( N_GND_c_8_p N_noxref_14_c_2610_n ) capacitor c=0.0117685f //x=25.53 \
 //y=0 //x2=7.255 //y2=0.54
cc_175 ( N_GND_c_58_p N_noxref_14_c_2610_n ) capacitor c=0.0362073f //x=9.45 \
 //y=0 //x2=7.255 //y2=0.54
cc_176 ( N_GND_c_2_p N_noxref_14_c_2610_n ) capacitor c=0.00177266f //x=25.53 \
 //y=0 //x2=7.255 //y2=0.54
cc_177 ( N_GND_c_8_p N_noxref_14_M3_noxref_s ) capacitor c=0.00575103f \
 //x=25.53 //y=0 //x2=5.265 //y2=0.375
cc_178 ( N_GND_c_10_p N_noxref_14_M3_noxref_s ) capacitor c=0.014327f //x=5.8 \
 //y=0 //x2=5.265 //y2=0.375
cc_179 ( N_GND_c_58_p N_noxref_14_M3_noxref_s ) capacitor c=0.0133864f \
 //x=9.45 //y=0 //x2=5.265 //y2=0.375
cc_180 ( N_GND_c_3_p N_noxref_14_M3_noxref_s ) capacitor c=0.0696963f //x=4.81 \
 //y=0 //x2=5.265 //y2=0.375
cc_181 ( N_GND_c_4_p N_noxref_14_M3_noxref_s ) capacitor c=3.31601e-19 \
 //x=9.62 //y=0 //x2=5.265 //y2=0.375
cc_182 ( N_GND_M3_noxref_d N_noxref_14_M3_noxref_s ) capacitor c=0.033718f \
 //x=5.695 //y=0.875 //x2=5.265 //y2=0.375
cc_183 ( N_GND_c_8_p N_noxref_15_c_2653_n ) capacitor c=0.00385233f //x=25.53 \
 //y=0 //x2=7.825 //y2=0.995
cc_184 ( N_GND_c_58_p N_noxref_15_c_2653_n ) capacitor c=0.0094913f //x=9.45 \
 //y=0 //x2=7.825 //y2=0.995
cc_185 ( N_GND_c_8_p N_noxref_15_c_2655_n ) capacitor c=0.00287639f //x=25.53 \
 //y=0 //x2=7.91 //y2=0.625
cc_186 ( N_GND_c_58_p N_noxref_15_c_2655_n ) capacitor c=0.014327f //x=9.45 \
 //y=0 //x2=7.91 //y2=0.625
cc_187 ( N_GND_M3_noxref_d N_noxref_15_c_2655_n ) capacitor c=6.21394e-19 \
 //x=5.695 //y=0.875 //x2=7.91 //y2=0.625
cc_188 ( N_GND_c_8_p N_noxref_15_c_2658_n ) capacitor c=0.0105197f //x=25.53 \
 //y=0 //x2=8.795 //y2=0.54
cc_189 ( N_GND_c_58_p N_noxref_15_c_2658_n ) capacitor c=0.036368f //x=9.45 \
 //y=0 //x2=8.795 //y2=0.54
cc_190 ( N_GND_c_2_p N_noxref_15_c_2658_n ) capacitor c=0.00189358f //x=25.53 \
 //y=0 //x2=8.795 //y2=0.54
cc_191 ( N_GND_c_8_p N_noxref_15_c_2661_n ) capacitor c=0.00254232f //x=25.53 \
 //y=0 //x2=8.88 //y2=0.625
cc_192 ( N_GND_c_58_p N_noxref_15_c_2661_n ) capacitor c=0.0140304f //x=9.45 \
 //y=0 //x2=8.88 //y2=0.625
cc_193 ( N_GND_c_4_p N_noxref_15_c_2661_n ) capacitor c=0.0404137f //x=9.62 \
 //y=0 //x2=8.88 //y2=0.625
cc_194 ( N_GND_M3_noxref_d N_noxref_15_M4_noxref_d ) capacitor c=0.00162435f \
 //x=5.695 //y=0.875 //x2=6.67 //y2=0.91
cc_195 ( N_GND_c_3_p N_noxref_15_M5_noxref_s ) capacitor c=8.16352e-19 \
 //x=4.81 //y=0 //x2=7.775 //y2=0.375
cc_196 ( N_GND_c_4_p N_noxref_15_M5_noxref_s ) capacitor c=0.00183576f \
 //x=9.62 //y=0 //x2=7.775 //y2=0.375
cc_197 ( N_GND_c_8_p N_noxref_16_c_2707_n ) capacitor c=0.00517234f //x=25.53 \
 //y=0 //x2=11.2 //y2=1.58
cc_198 ( N_GND_c_17_p N_noxref_16_c_2707_n ) capacitor c=0.00112872f \
 //x=10.715 //y=0 //x2=11.2 //y2=1.58
cc_199 ( N_GND_c_24_p N_noxref_16_c_2707_n ) capacitor c=0.0018229f //x=12.78 \
 //y=0 //x2=11.2 //y2=1.58
cc_200 ( N_GND_M6_noxref_d N_noxref_16_c_2707_n ) capacitor c=0.008625f \
 //x=10.61 //y=0.865 //x2=11.2 //y2=1.58
cc_201 ( N_GND_c_8_p N_noxref_16_c_2711_n ) capacitor c=0.00259029f //x=25.53 \
 //y=0 //x2=11.285 //y2=0.615
cc_202 ( N_GND_c_24_p N_noxref_16_c_2711_n ) capacitor c=0.0146901f //x=12.78 \
 //y=0 //x2=11.285 //y2=0.615
cc_203 ( N_GND_M6_noxref_d N_noxref_16_c_2711_n ) capacitor c=0.033812f \
 //x=10.61 //y=0.865 //x2=11.285 //y2=0.615
cc_204 ( N_GND_c_4_p N_noxref_16_c_2714_n ) capacitor c=2.91423e-19 //x=9.62 \
 //y=0 //x2=11.285 //y2=1.495
cc_205 ( N_GND_c_8_p N_noxref_16_c_2715_n ) capacitor c=0.0106919f //x=25.53 \
 //y=0 //x2=12.17 //y2=0.53
cc_206 ( N_GND_c_24_p N_noxref_16_c_2715_n ) capacitor c=0.0374253f //x=12.78 \
 //y=0 //x2=12.17 //y2=0.53
cc_207 ( N_GND_c_2_p N_noxref_16_c_2715_n ) capacitor c=0.00198372f //x=25.53 \
 //y=0 //x2=12.17 //y2=0.53
cc_208 ( N_GND_c_8_p N_noxref_16_c_2718_n ) capacitor c=0.00258845f //x=25.53 \
 //y=0 //x2=12.255 //y2=0.615
cc_209 ( N_GND_c_24_p N_noxref_16_c_2718_n ) capacitor c=0.0146256f //x=12.78 \
 //y=0 //x2=12.255 //y2=0.615
cc_210 ( N_GND_c_5_p N_noxref_16_c_2718_n ) capacitor c=0.0431718f //x=12.95 \
 //y=0 //x2=12.255 //y2=0.615
cc_211 ( N_GND_c_8_p N_noxref_16_M6_noxref_s ) capacitor c=0.00259029f \
 //x=25.53 //y=0 //x2=10.18 //y2=0.365
cc_212 ( N_GND_c_17_p N_noxref_16_M6_noxref_s ) capacitor c=0.0146901f \
 //x=10.715 //y=0 //x2=10.18 //y2=0.365
cc_213 ( N_GND_c_4_p N_noxref_16_M6_noxref_s ) capacitor c=0.0583534f //x=9.62 \
 //y=0 //x2=10.18 //y2=0.365
cc_214 ( N_GND_c_5_p N_noxref_16_M6_noxref_s ) capacitor c=0.00198098f \
 //x=12.95 //y=0 //x2=10.18 //y2=0.365
cc_215 ( N_GND_M6_noxref_d N_noxref_16_M6_noxref_s ) capacitor c=0.0334197f \
 //x=10.61 //y=0.865 //x2=10.18 //y2=0.365
cc_216 ( N_GND_c_8_p N_noxref_17_c_2759_n ) capacitor c=0.00517576f //x=25.53 \
 //y=0 //x2=14.425 //y2=1.59
cc_217 ( N_GND_c_32_p N_noxref_17_c_2759_n ) capacitor c=0.00111448f //x=13.94 \
 //y=0 //x2=14.425 //y2=1.59
cc_218 ( N_GND_c_39_p N_noxref_17_c_2759_n ) capacitor c=0.00180612f //x=17.59 \
 //y=0 //x2=14.425 //y2=1.59
cc_219 ( N_GND_M8_noxref_d N_noxref_17_c_2759_n ) capacitor c=0.00853078f \
 //x=13.835 //y=0.875 //x2=14.425 //y2=1.59
cc_220 ( N_GND_c_8_p N_noxref_17_c_2763_n ) capacitor c=0.00254475f //x=25.53 \
 //y=0 //x2=14.51 //y2=0.625
cc_221 ( N_GND_c_39_p N_noxref_17_c_2763_n ) capacitor c=0.0140928f //x=17.59 \
 //y=0 //x2=14.51 //y2=0.625
cc_222 ( N_GND_M8_noxref_d N_noxref_17_c_2763_n ) capacitor c=0.033954f \
 //x=13.835 //y=0.875 //x2=14.51 //y2=0.625
cc_223 ( N_GND_c_8_p N_noxref_17_c_2766_n ) capacitor c=0.0104506f //x=25.53 \
 //y=0 //x2=15.395 //y2=0.54
cc_224 ( N_GND_c_39_p N_noxref_17_c_2766_n ) capacitor c=0.0360726f //x=17.59 \
 //y=0 //x2=15.395 //y2=0.54
cc_225 ( N_GND_c_2_p N_noxref_17_c_2766_n ) capacitor c=0.00177266f //x=25.53 \
 //y=0 //x2=15.395 //y2=0.54
cc_226 ( N_GND_c_8_p N_noxref_17_M8_noxref_s ) capacitor c=0.00507657f \
 //x=25.53 //y=0 //x2=13.405 //y2=0.375
cc_227 ( N_GND_c_32_p N_noxref_17_M8_noxref_s ) capacitor c=0.0140928f \
 //x=13.94 //y=0 //x2=13.405 //y2=0.375
cc_228 ( N_GND_c_39_p N_noxref_17_M8_noxref_s ) capacitor c=0.0131437f \
 //x=17.59 //y=0 //x2=13.405 //y2=0.375
cc_229 ( N_GND_c_5_p N_noxref_17_M8_noxref_s ) capacitor c=0.0696963f \
 //x=12.95 //y=0 //x2=13.405 //y2=0.375
cc_230 ( N_GND_c_6_p N_noxref_17_M8_noxref_s ) capacitor c=3.31601e-19 \
 //x=17.76 //y=0 //x2=13.405 //y2=0.375
cc_231 ( N_GND_M8_noxref_d N_noxref_17_M8_noxref_s ) capacitor c=0.033718f \
 //x=13.835 //y=0.875 //x2=13.405 //y2=0.375
cc_232 ( N_GND_c_8_p N_noxref_18_c_2809_n ) capacitor c=0.00352952f //x=25.53 \
 //y=0 //x2=15.965 //y2=0.995
cc_233 ( N_GND_c_39_p N_noxref_18_c_2809_n ) capacitor c=0.00934524f //x=17.59 \
 //y=0 //x2=15.965 //y2=0.995
cc_234 ( N_GND_c_8_p N_noxref_18_c_2811_n ) capacitor c=0.00254475f //x=25.53 \
 //y=0 //x2=16.05 //y2=0.625
cc_235 ( N_GND_c_39_p N_noxref_18_c_2811_n ) capacitor c=0.0140928f //x=17.59 \
 //y=0 //x2=16.05 //y2=0.625
cc_236 ( N_GND_M8_noxref_d N_noxref_18_c_2811_n ) capacitor c=6.21394e-19 \
 //x=13.835 //y=0.875 //x2=16.05 //y2=0.625
cc_237 ( N_GND_c_8_p N_noxref_18_c_2814_n ) capacitor c=0.0105197f //x=25.53 \
 //y=0 //x2=16.935 //y2=0.54
cc_238 ( N_GND_c_39_p N_noxref_18_c_2814_n ) capacitor c=0.0364139f //x=17.59 \
 //y=0 //x2=16.935 //y2=0.54
cc_239 ( N_GND_c_2_p N_noxref_18_c_2814_n ) capacitor c=0.00189358f //x=25.53 \
 //y=0 //x2=16.935 //y2=0.54
cc_240 ( N_GND_c_8_p N_noxref_18_c_2817_n ) capacitor c=0.00254232f //x=25.53 \
 //y=0 //x2=17.02 //y2=0.625
cc_241 ( N_GND_c_39_p N_noxref_18_c_2817_n ) capacitor c=0.0140304f //x=17.59 \
 //y=0 //x2=17.02 //y2=0.625
cc_242 ( N_GND_c_6_p N_noxref_18_c_2817_n ) capacitor c=0.0404137f //x=17.76 \
 //y=0 //x2=17.02 //y2=0.625
cc_243 ( N_GND_M8_noxref_d N_noxref_18_M9_noxref_d ) capacitor c=0.00162435f \
 //x=13.835 //y=0.875 //x2=14.81 //y2=0.91
cc_244 ( N_GND_c_5_p N_noxref_18_M10_noxref_s ) capacitor c=8.16352e-19 \
 //x=12.95 //y=0 //x2=15.915 //y2=0.375
cc_245 ( N_GND_c_6_p N_noxref_18_M10_noxref_s ) capacitor c=0.00183204f \
 //x=17.76 //y=0 //x2=15.915 //y2=0.375
cc_246 ( N_GND_c_8_p N_noxref_19_c_2863_n ) capacitor c=0.00517576f //x=25.53 \
 //y=0 //x2=19.235 //y2=1.59
cc_247 ( N_GND_c_61_p N_noxref_19_c_2863_n ) capacitor c=0.00111448f //x=18.75 \
 //y=0 //x2=19.235 //y2=1.59
cc_248 ( N_GND_c_68_p N_noxref_19_c_2863_n ) capacitor c=0.00180612f //x=22.4 \
 //y=0 //x2=19.235 //y2=1.59
cc_249 ( N_GND_M11_noxref_d N_noxref_19_c_2863_n ) capacitor c=0.00853078f \
 //x=18.645 //y=0.875 //x2=19.235 //y2=1.59
cc_250 ( N_GND_c_8_p N_noxref_19_c_2867_n ) capacitor c=0.00254475f //x=25.53 \
 //y=0 //x2=19.32 //y2=0.625
cc_251 ( N_GND_c_68_p N_noxref_19_c_2867_n ) capacitor c=0.0140928f //x=22.4 \
 //y=0 //x2=19.32 //y2=0.625
cc_252 ( N_GND_M11_noxref_d N_noxref_19_c_2867_n ) capacitor c=0.033954f \
 //x=18.645 //y=0.875 //x2=19.32 //y2=0.625
cc_253 ( N_GND_c_8_p N_noxref_19_c_2870_n ) capacitor c=0.0113218f //x=25.53 \
 //y=0 //x2=20.205 //y2=0.54
cc_254 ( N_GND_c_68_p N_noxref_19_c_2870_n ) capacitor c=0.0358495f //x=22.4 \
 //y=0 //x2=20.205 //y2=0.54
cc_255 ( N_GND_c_2_p N_noxref_19_c_2870_n ) capacitor c=0.00177266f //x=25.53 \
 //y=0 //x2=20.205 //y2=0.54
cc_256 ( N_GND_c_8_p N_noxref_19_M11_noxref_s ) capacitor c=0.00798327f \
 //x=25.53 //y=0 //x2=18.215 //y2=0.375
cc_257 ( N_GND_c_61_p N_noxref_19_M11_noxref_s ) capacitor c=0.0140928f \
 //x=18.75 //y=0 //x2=18.215 //y2=0.375
cc_258 ( N_GND_c_68_p N_noxref_19_M11_noxref_s ) capacitor c=0.0131422f \
 //x=22.4 //y=0 //x2=18.215 //y2=0.375
cc_259 ( N_GND_c_6_p N_noxref_19_M11_noxref_s ) capacitor c=0.0696963f \
 //x=17.76 //y=0 //x2=18.215 //y2=0.375
cc_260 ( N_GND_c_7_p N_noxref_19_M11_noxref_s ) capacitor c=3.31601e-19 \
 //x=22.57 //y=0 //x2=18.215 //y2=0.375
cc_261 ( N_GND_M11_noxref_d N_noxref_19_M11_noxref_s ) capacitor c=0.033718f \
 //x=18.645 //y=0.875 //x2=18.215 //y2=0.375
cc_262 ( N_GND_c_8_p N_noxref_20_c_2915_n ) capacitor c=0.00402784f //x=25.53 \
 //y=0 //x2=20.775 //y2=0.995
cc_263 ( N_GND_c_68_p N_noxref_20_c_2915_n ) capacitor c=0.00829979f //x=22.4 \
 //y=0 //x2=20.775 //y2=0.995
cc_264 ( N_GND_c_8_p N_noxref_20_c_2917_n ) capacitor c=0.00575184f //x=25.53 \
 //y=0 //x2=20.86 //y2=0.625
cc_265 ( N_GND_c_68_p N_noxref_20_c_2917_n ) capacitor c=0.0140218f //x=22.4 \
 //y=0 //x2=20.86 //y2=0.625
cc_266 ( N_GND_M11_noxref_d N_noxref_20_c_2917_n ) capacitor c=6.21394e-19 \
 //x=18.645 //y=0.875 //x2=20.86 //y2=0.625
cc_267 ( N_GND_c_8_p N_noxref_20_c_2920_n ) capacitor c=0.0121783f //x=25.53 \
 //y=0 //x2=21.745 //y2=0.54
cc_268 ( N_GND_c_68_p N_noxref_20_c_2920_n ) capacitor c=0.0362762f //x=22.4 \
 //y=0 //x2=21.745 //y2=0.54
cc_269 ( N_GND_c_2_p N_noxref_20_c_2920_n ) capacitor c=0.00189358f //x=25.53 \
 //y=0 //x2=21.745 //y2=0.54
cc_270 ( N_GND_c_8_p N_noxref_20_c_2923_n ) capacitor c=0.00286759f //x=25.53 \
 //y=0 //x2=21.83 //y2=0.625
cc_271 ( N_GND_c_68_p N_noxref_20_c_2923_n ) capacitor c=0.0142605f //x=22.4 \
 //y=0 //x2=21.83 //y2=0.625
cc_272 ( N_GND_c_7_p N_noxref_20_c_2923_n ) capacitor c=0.0404137f //x=22.57 \
 //y=0 //x2=21.83 //y2=0.625
cc_273 ( N_GND_M11_noxref_d N_noxref_20_M12_noxref_d ) capacitor c=0.00162435f \
 //x=18.645 //y=0.875 //x2=19.62 //y2=0.91
cc_274 ( N_GND_c_6_p N_noxref_20_M13_noxref_s ) capacitor c=8.16352e-19 \
 //x=17.76 //y=0 //x2=20.725 //y2=0.375
cc_275 ( N_GND_c_7_p N_noxref_20_M13_noxref_s ) capacitor c=0.00183576f \
 //x=22.57 //y=0 //x2=20.725 //y2=0.375
cc_276 ( N_GND_c_8_p N_noxref_21_c_2967_n ) capacitor c=0.00556119f //x=25.53 \
 //y=0 //x2=24.15 //y2=1.58
cc_277 ( N_GND_c_92_p N_noxref_21_c_2967_n ) capacitor c=0.00113001f \
 //x=23.665 //y=0 //x2=24.15 //y2=1.58
cc_278 ( N_GND_c_2_p N_noxref_21_c_2967_n ) capacitor c=0.00180846f //x=25.53 \
 //y=0 //x2=24.15 //y2=1.58
cc_279 ( N_GND_M14_noxref_d N_noxref_21_c_2967_n ) capacitor c=0.00897268f \
 //x=23.56 //y=0.865 //x2=24.15 //y2=1.58
cc_280 ( N_GND_c_8_p N_noxref_21_c_2971_n ) capacitor c=0.00302994f //x=25.53 \
 //y=0 //x2=24.235 //y2=0.615
cc_281 ( N_GND_c_2_p N_noxref_21_c_2971_n ) capacitor c=0.0146208f //x=25.53 \
 //y=0 //x2=24.235 //y2=0.615
cc_282 ( N_GND_M14_noxref_d N_noxref_21_c_2971_n ) capacitor c=0.033812f \
 //x=23.56 //y=0.865 //x2=24.235 //y2=0.615
cc_283 ( N_GND_c_7_p N_noxref_21_c_2974_n ) capacitor c=2.91423e-19 //x=22.57 \
 //y=0 //x2=24.235 //y2=1.495
cc_284 ( N_GND_c_8_p N_noxref_21_c_2975_n ) capacitor c=0.0124196f //x=25.53 \
 //y=0 //x2=25.12 //y2=0.53
cc_285 ( N_GND_c_2_p N_noxref_21_c_2975_n ) capacitor c=0.0390872f //x=25.53 \
 //y=0 //x2=25.12 //y2=0.53
cc_286 ( N_GND_c_8_p N_noxref_21_c_2977_n ) capacitor c=0.00302319f //x=25.53 \
 //y=0 //x2=25.205 //y2=0.615
cc_287 ( N_GND_c_2_p N_noxref_21_c_2977_n ) capacitor c=0.0584079f //x=25.53 \
 //y=0 //x2=25.205 //y2=0.615
cc_288 ( N_GND_c_8_p N_noxref_21_M14_noxref_s ) capacitor c=0.00293348f \
 //x=25.53 //y=0 //x2=23.13 //y2=0.365
cc_289 ( N_GND_c_92_p N_noxref_21_M14_noxref_s ) capacitor c=0.0149357f \
 //x=23.665 //y=0 //x2=23.13 //y2=0.365
cc_290 ( N_GND_c_2_p N_noxref_21_M14_noxref_s ) capacitor c=0.00198482f \
 //x=25.53 //y=0 //x2=23.13 //y2=0.365
cc_291 ( N_GND_c_7_p N_noxref_21_M14_noxref_s ) capacitor c=0.0583534f \
 //x=22.57 //y=0 //x2=23.13 //y2=0.365
cc_292 ( N_GND_M14_noxref_d N_noxref_21_M14_noxref_s ) capacitor c=0.0334197f \
 //x=23.56 //y=0.865 //x2=23.13 //y2=0.365
cc_293 ( N_VDD_c_295_n N_noxref_3_c_622_n ) capacitor c=6.58823e-19 //x=4.81 \
 //y=7.4 //x2=3.33 //y2=2.08
cc_294 ( N_VDD_c_301_p N_noxref_3_c_637_n ) capacitor c=0.00444892f //x=25.53 \
 //y=7.4 //x2=7.135 //y2=5.155
cc_295 ( N_VDD_c_302_p N_noxref_3_c_637_n ) capacitor c=4.31931e-19 //x=6.695 \
 //y=7.4 //x2=7.135 //y2=5.155
cc_296 ( N_VDD_c_303_p N_noxref_3_c_637_n ) capacitor c=4.31931e-19 //x=7.575 \
 //y=7.4 //x2=7.135 //y2=5.155
cc_297 ( N_VDD_M23_noxref_d N_noxref_3_c_637_n ) capacitor c=0.0112985f \
 //x=6.635 //y=5.02 //x2=7.135 //y2=5.155
cc_298 ( N_VDD_c_295_n N_noxref_3_c_641_n ) capacitor c=0.00863585f //x=4.81 \
 //y=7.4 //x2=6.425 //y2=5.155
cc_299 ( N_VDD_M22_noxref_s N_noxref_3_c_641_n ) capacitor c=0.0831083f \
 //x=5.765 //y=5.02 //x2=6.425 //y2=5.155
cc_300 ( N_VDD_c_301_p N_noxref_3_c_643_n ) capacitor c=0.0044221f //x=25.53 \
 //y=7.4 //x2=8.015 //y2=5.155
cc_301 ( N_VDD_c_303_p N_noxref_3_c_643_n ) capacitor c=4.31931e-19 //x=7.575 \
 //y=7.4 //x2=8.015 //y2=5.155
cc_302 ( N_VDD_c_309_p N_noxref_3_c_643_n ) capacitor c=4.31931e-19 //x=8.455 \
 //y=7.4 //x2=8.015 //y2=5.155
cc_303 ( N_VDD_M25_noxref_d N_noxref_3_c_643_n ) capacitor c=0.0112985f \
 //x=7.515 //y=5.02 //x2=8.015 //y2=5.155
cc_304 ( N_VDD_c_301_p N_noxref_3_c_647_n ) capacitor c=0.00434174f //x=25.53 \
 //y=7.4 //x2=8.795 //y2=5.155
cc_305 ( N_VDD_c_309_p N_noxref_3_c_647_n ) capacitor c=7.46626e-19 //x=8.455 \
 //y=7.4 //x2=8.795 //y2=5.155
cc_306 ( N_VDD_c_313_p N_noxref_3_c_647_n ) capacitor c=0.00198565f //x=9.45 \
 //y=7.4 //x2=8.795 //y2=5.155
cc_307 ( N_VDD_M27_noxref_d N_noxref_3_c_647_n ) capacitor c=0.0112985f \
 //x=8.395 //y=5.02 //x2=8.795 //y2=5.155
cc_308 ( N_VDD_c_296_n N_noxref_3_c_651_n ) capacitor c=0.0426864f //x=9.62 \
 //y=7.4 //x2=8.88 //y2=3.33
cc_309 ( N_VDD_c_301_p N_noxref_3_c_624_n ) capacitor c=0.00125279f //x=25.53 \
 //y=7.4 //x2=10.73 //y2=2.08
cc_310 ( N_VDD_c_317_p N_noxref_3_c_624_n ) capacitor c=2.87256e-19 //x=11.205 \
 //y=7.4 //x2=10.73 //y2=2.08
cc_311 ( N_VDD_c_296_n N_noxref_3_c_624_n ) capacitor c=0.0134208f //x=9.62 \
 //y=7.4 //x2=10.73 //y2=2.08
cc_312 ( N_VDD_c_319_p N_noxref_3_M20_noxref_g ) capacitor c=0.00675175f \
 //x=3.645 //y=7.4 //x2=3.07 //y2=6.02
cc_313 ( N_VDD_M19_noxref_d N_noxref_3_M20_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=3.07 //y2=6.02
cc_314 ( N_VDD_c_319_p N_noxref_3_M21_noxref_g ) capacitor c=0.00675379f \
 //x=3.645 //y=7.4 //x2=3.51 //y2=6.02
cc_315 ( N_VDD_M21_noxref_d N_noxref_3_M21_noxref_g ) capacitor c=0.0394719f \
 //x=3.585 //y=5.02 //x2=3.51 //y2=6.02
cc_316 ( N_VDD_c_317_p N_noxref_3_M28_noxref_g ) capacitor c=0.00726866f \
 //x=11.205 //y=7.4 //x2=10.63 //y2=6.02
cc_317 ( N_VDD_M28_noxref_s N_noxref_3_M28_noxref_g ) capacitor c=0.054195f \
 //x=10.275 //y=5.02 //x2=10.63 //y2=6.02
cc_318 ( N_VDD_c_317_p N_noxref_3_M29_noxref_g ) capacitor c=0.00672952f \
 //x=11.205 //y=7.4 //x2=11.07 //y2=6.02
cc_319 ( N_VDD_M29_noxref_d N_noxref_3_M29_noxref_g ) capacitor c=0.015318f \
 //x=11.145 //y=5.02 //x2=11.07 //y2=6.02
cc_320 ( N_VDD_c_296_n N_noxref_3_c_663_n ) capacitor c=0.0154093f //x=9.62 \
 //y=7.4 //x2=10.73 //y2=4.7
cc_321 ( N_VDD_c_301_p N_noxref_3_M22_noxref_d ) capacitor c=0.00275235f \
 //x=25.53 //y=7.4 //x2=6.195 //y2=5.02
cc_322 ( N_VDD_c_302_p N_noxref_3_M22_noxref_d ) capacitor c=0.014035f \
 //x=6.695 //y=7.4 //x2=6.195 //y2=5.02
cc_323 ( N_VDD_M23_noxref_d N_noxref_3_M22_noxref_d ) capacitor c=0.0664752f \
 //x=6.635 //y=5.02 //x2=6.195 //y2=5.02
cc_324 ( N_VDD_c_301_p N_noxref_3_M24_noxref_d ) capacitor c=0.00275235f \
 //x=25.53 //y=7.4 //x2=7.075 //y2=5.02
cc_325 ( N_VDD_c_303_p N_noxref_3_M24_noxref_d ) capacitor c=0.014035f \
 //x=7.575 //y=7.4 //x2=7.075 //y2=5.02
cc_326 ( N_VDD_c_296_n N_noxref_3_M24_noxref_d ) capacitor c=4.9285e-19 \
 //x=9.62 //y=7.4 //x2=7.075 //y2=5.02
cc_327 ( N_VDD_M22_noxref_s N_noxref_3_M24_noxref_d ) capacitor c=0.00130656f \
 //x=5.765 //y=5.02 //x2=7.075 //y2=5.02
cc_328 ( N_VDD_M23_noxref_d N_noxref_3_M24_noxref_d ) capacitor c=0.0664752f \
 //x=6.635 //y=5.02 //x2=7.075 //y2=5.02
cc_329 ( N_VDD_M25_noxref_d N_noxref_3_M24_noxref_d ) capacitor c=0.0664752f \
 //x=7.515 //y=5.02 //x2=7.075 //y2=5.02
cc_330 ( N_VDD_c_301_p N_noxref_3_M26_noxref_d ) capacitor c=0.00275235f \
 //x=25.53 //y=7.4 //x2=7.955 //y2=5.02
cc_331 ( N_VDD_c_309_p N_noxref_3_M26_noxref_d ) capacitor c=0.014035f \
 //x=8.455 //y=7.4 //x2=7.955 //y2=5.02
cc_332 ( N_VDD_c_296_n N_noxref_3_M26_noxref_d ) capacitor c=0.00939849f \
 //x=9.62 //y=7.4 //x2=7.955 //y2=5.02
cc_333 ( N_VDD_M25_noxref_d N_noxref_3_M26_noxref_d ) capacitor c=0.0664752f \
 //x=7.515 //y=5.02 //x2=7.955 //y2=5.02
cc_334 ( N_VDD_M27_noxref_d N_noxref_3_M26_noxref_d ) capacitor c=0.0664752f \
 //x=8.395 //y=5.02 //x2=7.955 //y2=5.02
cc_335 ( N_VDD_M28_noxref_s N_noxref_3_M26_noxref_d ) capacitor c=4.52683e-19 \
 //x=10.275 //y=5.02 //x2=7.955 //y2=5.02
cc_336 ( N_VDD_c_301_p N_noxref_4_c_879_n ) capacitor c=0.00453663f //x=25.53 \
 //y=7.4 //x2=11.645 //y2=5.2
cc_337 ( N_VDD_c_317_p N_noxref_4_c_879_n ) capacitor c=4.48391e-19 //x=11.205 \
 //y=7.4 //x2=11.645 //y2=5.2
cc_338 ( N_VDD_c_345_p N_noxref_4_c_879_n ) capacitor c=4.48391e-19 //x=12.085 \
 //y=7.4 //x2=11.645 //y2=5.2
cc_339 ( N_VDD_M29_noxref_d N_noxref_4_c_879_n ) capacitor c=0.0124542f \
 //x=11.145 //y=5.02 //x2=11.645 //y2=5.2
cc_340 ( N_VDD_c_296_n N_noxref_4_c_883_n ) capacitor c=0.00985474f //x=9.62 \
 //y=7.4 //x2=10.935 //y2=5.2
cc_341 ( N_VDD_M28_noxref_s N_noxref_4_c_883_n ) capacitor c=0.087833f \
 //x=10.275 //y=5.02 //x2=10.935 //y2=5.2
cc_342 ( N_VDD_c_301_p N_noxref_4_c_885_n ) capacitor c=0.00301575f //x=25.53 \
 //y=7.4 //x2=12.125 //y2=5.2
cc_343 ( N_VDD_c_345_p N_noxref_4_c_885_n ) capacitor c=7.72068e-19 //x=12.085 \
 //y=7.4 //x2=12.125 //y2=5.2
cc_344 ( N_VDD_M31_noxref_d N_noxref_4_c_885_n ) capacitor c=0.0158515f \
 //x=12.025 //y=5.02 //x2=12.125 //y2=5.2
cc_345 ( N_VDD_c_296_n N_noxref_4_c_864_n ) capacitor c=0.00151618f //x=9.62 \
 //y=7.4 //x2=12.21 //y2=3.33
cc_346 ( N_VDD_c_297_n N_noxref_4_c_864_n ) capacitor c=0.0428942f //x=12.95 \
 //y=7.4 //x2=12.21 //y2=3.33
cc_347 ( N_VDD_c_301_p N_noxref_4_c_865_n ) capacitor c=9.10347e-19 //x=25.53 \
 //y=7.4 //x2=14.06 //y2=2.08
cc_348 ( N_VDD_c_297_n N_noxref_4_c_865_n ) capacitor c=0.0133749f //x=12.95 \
 //y=7.4 //x2=14.06 //y2=2.08
cc_349 ( N_VDD_M32_noxref_s N_noxref_4_c_865_n ) capacitor c=0.0125322f \
 //x=13.905 //y=5.02 //x2=14.06 //y2=2.08
cc_350 ( N_VDD_c_357_p N_noxref_4_M32_noxref_g ) capacitor c=0.00749687f \
 //x=14.835 //y=7.4 //x2=14.26 //y2=6.02
cc_351 ( N_VDD_M32_noxref_s N_noxref_4_M32_noxref_g ) capacitor c=0.0477201f \
 //x=13.905 //y=5.02 //x2=14.26 //y2=6.02
cc_352 ( N_VDD_c_357_p N_noxref_4_M33_noxref_g ) capacitor c=0.00675175f \
 //x=14.835 //y=7.4 //x2=14.7 //y2=6.02
cc_353 ( N_VDD_M33_noxref_d N_noxref_4_M33_noxref_g ) capacitor c=0.015318f \
 //x=14.775 //y=5.02 //x2=14.7 //y2=6.02
cc_354 ( N_VDD_c_297_n N_noxref_4_c_897_n ) capacitor c=0.00757682f //x=12.95 \
 //y=7.4 //x2=14.335 //y2=4.79
cc_355 ( N_VDD_M32_noxref_s N_noxref_4_c_897_n ) capacitor c=0.00444914f \
 //x=13.905 //y=5.02 //x2=14.335 //y2=4.79
cc_356 ( N_VDD_c_301_p N_noxref_4_M28_noxref_d ) capacitor c=0.00275225f \
 //x=25.53 //y=7.4 //x2=10.705 //y2=5.02
cc_357 ( N_VDD_c_317_p N_noxref_4_M28_noxref_d ) capacitor c=0.0140317f \
 //x=11.205 //y=7.4 //x2=10.705 //y2=5.02
cc_358 ( N_VDD_c_297_n N_noxref_4_M28_noxref_d ) capacitor c=6.94454e-19 \
 //x=12.95 //y=7.4 //x2=10.705 //y2=5.02
cc_359 ( N_VDD_M29_noxref_d N_noxref_4_M28_noxref_d ) capacitor c=0.0664752f \
 //x=11.145 //y=5.02 //x2=10.705 //y2=5.02
cc_360 ( N_VDD_c_301_p N_noxref_4_M30_noxref_d ) capacitor c=0.00275225f \
 //x=25.53 //y=7.4 //x2=11.585 //y2=5.02
cc_361 ( N_VDD_c_345_p N_noxref_4_M30_noxref_d ) capacitor c=0.0140317f \
 //x=12.085 //y=7.4 //x2=11.585 //y2=5.02
cc_362 ( N_VDD_c_297_n N_noxref_4_M30_noxref_d ) capacitor c=0.0120541f \
 //x=12.95 //y=7.4 //x2=11.585 //y2=5.02
cc_363 ( N_VDD_M28_noxref_s N_noxref_4_M30_noxref_d ) capacitor c=0.00111971f \
 //x=10.275 //y=5.02 //x2=11.585 //y2=5.02
cc_364 ( N_VDD_M29_noxref_d N_noxref_4_M30_noxref_d ) capacitor c=0.0664752f \
 //x=11.145 //y=5.02 //x2=11.585 //y2=5.02
cc_365 ( N_VDD_M31_noxref_d N_noxref_4_M30_noxref_d ) capacitor c=0.0664752f \
 //x=12.025 //y=5.02 //x2=11.585 //y2=5.02
cc_366 ( N_VDD_M32_noxref_s N_noxref_4_M30_noxref_d ) capacitor c=3.73257e-19 \
 //x=13.905 //y=5.02 //x2=11.585 //y2=5.02
cc_367 ( N_VDD_c_301_p N_CLK_c_1011_n ) capacitor c=0.0971263f //x=25.53 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_368 ( N_VDD_c_375_p N_CLK_c_1011_n ) capacitor c=0.00258496f //x=4.64 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_369 ( N_VDD_c_376_p N_CLK_c_1011_n ) capacitor c=0.00328994f //x=5.815 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_370 ( N_VDD_c_302_p N_CLK_c_1011_n ) capacitor c=0.00135925f //x=6.695 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_371 ( N_VDD_c_313_p N_CLK_c_1011_n ) capacitor c=0.00258496f //x=9.45 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_372 ( N_VDD_c_379_p N_CLK_c_1011_n ) capacitor c=0.00209689f //x=10.325 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_373 ( N_VDD_c_317_p N_CLK_c_1011_n ) capacitor c=7.81728e-19 //x=11.205 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_374 ( N_VDD_c_381_p N_CLK_c_1011_n ) capacitor c=0.00205475f //x=12.78 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_375 ( N_VDD_c_382_p N_CLK_c_1011_n ) capacitor c=0.00328994f //x=13.955 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_376 ( N_VDD_c_357_p N_CLK_c_1011_n ) capacitor c=0.00135925f //x=14.835 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_377 ( N_VDD_c_295_n N_CLK_c_1011_n ) capacitor c=0.0389825f //x=4.81 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_378 ( N_VDD_c_296_n N_CLK_c_1011_n ) capacitor c=0.0389825f //x=9.62 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_379 ( N_VDD_c_297_n N_CLK_c_1011_n ) capacitor c=0.0389825f //x=12.95 \
 //y=7.4 //x2=15.055 //y2=4.44
cc_380 ( N_VDD_M22_noxref_s N_CLK_c_1011_n ) capacitor c=0.00179496f //x=5.765 \
 //y=5.02 //x2=15.055 //y2=4.44
cc_381 ( N_VDD_M28_noxref_s N_CLK_c_1011_n ) capacitor c=0.00541054f \
 //x=10.275 //y=5.02 //x2=15.055 //y2=4.44
cc_382 ( N_VDD_M31_noxref_d N_CLK_c_1011_n ) capacitor c=6.7165e-19 //x=12.025 \
 //y=5.02 //x2=15.055 //y2=4.44
cc_383 ( N_VDD_M32_noxref_s N_CLK_c_1011_n ) capacitor c=0.00179496f \
 //x=13.905 //y=5.02 //x2=15.055 //y2=4.44
cc_384 ( N_VDD_c_301_p N_CLK_c_1028_n ) capacitor c=0.00146064f //x=25.53 \
 //y=7.4 //x2=2.335 //y2=4.44
cc_385 ( N_VDD_c_301_p N_CLK_c_1009_n ) capacitor c=2.03287e-19 //x=25.53 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_386 ( N_VDD_c_293_n N_CLK_c_1009_n ) capacitor c=9.53425e-19 //x=0.74 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_387 ( N_VDD_c_301_p N_CLK_c_1010_n ) capacitor c=2.03287e-19 //x=25.53 \
 //y=7.4 //x2=15.17 //y2=2.08
cc_388 ( N_VDD_c_297_n N_CLK_c_1010_n ) capacitor c=6.15921e-19 //x=12.95 \
 //y=7.4 //x2=15.17 //y2=2.08
cc_389 ( N_VDD_c_396_p N_CLK_M18_noxref_g ) capacitor c=0.00676195f //x=2.765 \
 //y=7.4 //x2=2.19 //y2=6.02
cc_390 ( N_VDD_M17_noxref_d N_CLK_M18_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=2.19 //y2=6.02
cc_391 ( N_VDD_c_396_p N_CLK_M19_noxref_g ) capacitor c=0.00675175f //x=2.765 \
 //y=7.4 //x2=2.63 //y2=6.02
cc_392 ( N_VDD_M19_noxref_d N_CLK_M19_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=2.63 //y2=6.02
cc_393 ( N_VDD_c_400_p N_CLK_M34_noxref_g ) capacitor c=0.00676195f //x=15.715 \
 //y=7.4 //x2=15.14 //y2=6.02
cc_394 ( N_VDD_M33_noxref_d N_CLK_M34_noxref_g ) capacitor c=0.015318f \
 //x=14.775 //y=5.02 //x2=15.14 //y2=6.02
cc_395 ( N_VDD_c_400_p N_CLK_M35_noxref_g ) capacitor c=0.00675175f //x=15.715 \
 //y=7.4 //x2=15.58 //y2=6.02
cc_396 ( N_VDD_M35_noxref_d N_CLK_M35_noxref_g ) capacitor c=0.015318f \
 //x=15.655 //y=5.02 //x2=15.58 //y2=6.02
cc_397 ( N_VDD_c_301_p N_noxref_6_c_1249_n ) capacitor c=0.00449316f //x=25.53 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_398 ( N_VDD_c_405_p N_noxref_6_c_1249_n ) capacitor c=4.32228e-19 //x=1.885 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_399 ( N_VDD_c_396_p N_noxref_6_c_1249_n ) capacitor c=4.31906e-19 //x=2.765 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_400 ( N_VDD_M17_noxref_d N_noxref_6_c_1249_n ) capacitor c=0.0115147f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_401 ( N_VDD_c_293_n N_noxref_6_c_1253_n ) capacitor c=0.00880189f //x=0.74 \
 //y=7.4 //x2=1.615 //y2=5.155
cc_402 ( N_VDD_M16_noxref_s N_noxref_6_c_1253_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_403 ( N_VDD_c_301_p N_noxref_6_c_1255_n ) capacitor c=0.0044221f //x=25.53 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_404 ( N_VDD_c_396_p N_noxref_6_c_1255_n ) capacitor c=4.31931e-19 //x=2.765 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_405 ( N_VDD_c_319_p N_noxref_6_c_1255_n ) capacitor c=4.31931e-19 //x=3.645 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_406 ( N_VDD_M19_noxref_d N_noxref_6_c_1255_n ) capacitor c=0.0112985f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_407 ( N_VDD_c_301_p N_noxref_6_c_1259_n ) capacitor c=0.00434174f //x=25.53 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_408 ( N_VDD_c_319_p N_noxref_6_c_1259_n ) capacitor c=7.46626e-19 //x=3.645 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_409 ( N_VDD_c_375_p N_noxref_6_c_1259_n ) capacitor c=0.00198565f //x=4.64 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_410 ( N_VDD_M21_noxref_d N_noxref_6_c_1259_n ) capacitor c=0.0112985f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_411 ( N_VDD_c_295_n N_noxref_6_c_1263_n ) capacitor c=0.0427116f //x=4.81 \
 //y=7.4 //x2=4.07 //y2=3.7
cc_412 ( N_VDD_c_301_p N_noxref_6_c_1226_n ) capacitor c=9.10347e-19 //x=25.53 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_413 ( N_VDD_c_295_n N_noxref_6_c_1226_n ) capacitor c=0.0134711f //x=4.81 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_414 ( N_VDD_M22_noxref_s N_noxref_6_c_1226_n ) capacitor c=0.0120327f \
 //x=5.765 //y=5.02 //x2=5.92 //y2=2.08
cc_415 ( N_VDD_c_301_p N_noxref_6_c_1227_n ) capacitor c=9.23542e-19 //x=25.53 \
 //y=7.4 //x2=18.87 //y2=2.08
cc_416 ( N_VDD_c_298_n N_noxref_6_c_1227_n ) capacitor c=0.0160182f //x=17.76 \
 //y=7.4 //x2=18.87 //y2=2.08
cc_417 ( N_VDD_M38_noxref_s N_noxref_6_c_1227_n ) capacitor c=0.0123142f \
 //x=18.715 //y=5.02 //x2=18.87 //y2=2.08
cc_418 ( N_VDD_c_302_p N_noxref_6_M22_noxref_g ) capacitor c=0.00749687f \
 //x=6.695 //y=7.4 //x2=6.12 //y2=6.02
cc_419 ( N_VDD_M22_noxref_s N_noxref_6_M22_noxref_g ) capacitor c=0.0477201f \
 //x=5.765 //y=5.02 //x2=6.12 //y2=6.02
cc_420 ( N_VDD_c_302_p N_noxref_6_M23_noxref_g ) capacitor c=0.00675175f \
 //x=6.695 //y=7.4 //x2=6.56 //y2=6.02
cc_421 ( N_VDD_M23_noxref_d N_noxref_6_M23_noxref_g ) capacitor c=0.015318f \
 //x=6.635 //y=5.02 //x2=6.56 //y2=6.02
cc_422 ( N_VDD_c_429_p N_noxref_6_M38_noxref_g ) capacitor c=0.00749687f \
 //x=19.645 //y=7.4 //x2=19.07 //y2=6.02
cc_423 ( N_VDD_M38_noxref_s N_noxref_6_M38_noxref_g ) capacitor c=0.0477201f \
 //x=18.715 //y=5.02 //x2=19.07 //y2=6.02
cc_424 ( N_VDD_c_429_p N_noxref_6_M39_noxref_g ) capacitor c=0.00675175f \
 //x=19.645 //y=7.4 //x2=19.51 //y2=6.02
cc_425 ( N_VDD_M39_noxref_d N_noxref_6_M39_noxref_g ) capacitor c=0.015318f \
 //x=19.585 //y=5.02 //x2=19.51 //y2=6.02
cc_426 ( N_VDD_c_295_n N_noxref_6_c_1278_n ) capacitor c=0.00757682f //x=4.81 \
 //y=7.4 //x2=6.195 //y2=4.79
cc_427 ( N_VDD_M22_noxref_s N_noxref_6_c_1278_n ) capacitor c=0.00444914f \
 //x=5.765 //y=5.02 //x2=6.195 //y2=4.79
cc_428 ( N_VDD_c_298_n N_noxref_6_c_1280_n ) capacitor c=0.00757682f //x=17.76 \
 //y=7.4 //x2=19.145 //y2=4.79
cc_429 ( N_VDD_M38_noxref_s N_noxref_6_c_1280_n ) capacitor c=0.00445134f \
 //x=18.715 //y=5.02 //x2=19.145 //y2=4.79
cc_430 ( N_VDD_c_301_p N_noxref_6_M16_noxref_d ) capacitor c=0.00285091f \
 //x=25.53 //y=7.4 //x2=1.385 //y2=5.02
cc_431 ( N_VDD_c_405_p N_noxref_6_M16_noxref_d ) capacitor c=0.0141016f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_432 ( N_VDD_M17_noxref_d N_noxref_6_M16_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_433 ( N_VDD_c_301_p N_noxref_6_M18_noxref_d ) capacitor c=0.00275186f \
 //x=25.53 //y=7.4 //x2=2.265 //y2=5.02
cc_434 ( N_VDD_c_396_p N_noxref_6_M18_noxref_d ) capacitor c=0.0140346f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_435 ( N_VDD_c_295_n N_noxref_6_M18_noxref_d ) capacitor c=4.9285e-19 \
 //x=4.81 //y=7.4 //x2=2.265 //y2=5.02
cc_436 ( N_VDD_M16_noxref_s N_noxref_6_M18_noxref_d ) capacitor c=0.00130656f \
 //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_437 ( N_VDD_M17_noxref_d N_noxref_6_M18_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_438 ( N_VDD_M19_noxref_d N_noxref_6_M18_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_439 ( N_VDD_c_301_p N_noxref_6_M20_noxref_d ) capacitor c=0.00275235f \
 //x=25.53 //y=7.4 //x2=3.145 //y2=5.02
cc_440 ( N_VDD_c_319_p N_noxref_6_M20_noxref_d ) capacitor c=0.0137384f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_441 ( N_VDD_c_295_n N_noxref_6_M20_noxref_d ) capacitor c=0.00939849f \
 //x=4.81 //y=7.4 //x2=3.145 //y2=5.02
cc_442 ( N_VDD_M19_noxref_d N_noxref_6_M20_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_443 ( N_VDD_M21_noxref_d N_noxref_6_M20_noxref_d ) capacitor c=0.0664752f \
 //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_444 ( N_VDD_M22_noxref_s N_noxref_6_M20_noxref_d ) capacitor c=3.57641e-19 \
 //x=5.765 //y=5.02 //x2=3.145 //y2=5.02
cc_445 ( N_VDD_c_296_n N_RN_c_1485_n ) capacitor c=6.09414e-19 //x=9.62 \
 //y=7.4 //x2=8.14 //y2=2.08
cc_446 ( N_VDD_c_298_n N_RN_c_1486_n ) capacitor c=0.00120861f //x=17.76 \
 //y=7.4 //x2=16.28 //y2=2.08
cc_447 ( N_VDD_c_301_p N_RN_c_1487_n ) capacitor c=2.05828e-19 //x=25.53 \
 //y=7.4 //x2=19.98 //y2=2.08
cc_448 ( N_VDD_c_298_n N_RN_c_1487_n ) capacitor c=7.30063e-19 //x=17.76 \
 //y=7.4 //x2=19.98 //y2=2.08
cc_449 ( N_VDD_c_309_p N_RN_M26_noxref_g ) capacitor c=0.00675175f //x=8.455 \
 //y=7.4 //x2=7.88 //y2=6.02
cc_450 ( N_VDD_M25_noxref_d N_RN_M26_noxref_g ) capacitor c=0.015318f \
 //x=7.515 //y=5.02 //x2=7.88 //y2=6.02
cc_451 ( N_VDD_c_309_p N_RN_M27_noxref_g ) capacitor c=0.00675379f //x=8.455 \
 //y=7.4 //x2=8.32 //y2=6.02
cc_452 ( N_VDD_M27_noxref_d N_RN_M27_noxref_g ) capacitor c=0.0394719f \
 //x=8.395 //y=5.02 //x2=8.32 //y2=6.02
cc_453 ( N_VDD_c_460_p N_RN_M36_noxref_g ) capacitor c=0.00675175f //x=16.595 \
 //y=7.4 //x2=16.02 //y2=6.02
cc_454 ( N_VDD_M35_noxref_d N_RN_M36_noxref_g ) capacitor c=0.015318f \
 //x=15.655 //y=5.02 //x2=16.02 //y2=6.02
cc_455 ( N_VDD_c_460_p N_RN_M37_noxref_g ) capacitor c=0.00675379f //x=16.595 \
 //y=7.4 //x2=16.46 //y2=6.02
cc_456 ( N_VDD_M37_noxref_d N_RN_M37_noxref_g ) capacitor c=0.0394719f \
 //x=16.535 //y=5.02 //x2=16.46 //y2=6.02
cc_457 ( N_VDD_c_464_p N_RN_M40_noxref_g ) capacitor c=0.00676195f //x=20.525 \
 //y=7.4 //x2=19.95 //y2=6.02
cc_458 ( N_VDD_M39_noxref_d N_RN_M40_noxref_g ) capacitor c=0.015318f \
 //x=19.585 //y=5.02 //x2=19.95 //y2=6.02
cc_459 ( N_VDD_c_464_p N_RN_M41_noxref_g ) capacitor c=0.00675175f //x=20.525 \
 //y=7.4 //x2=20.39 //y2=6.02
cc_460 ( N_VDD_M41_noxref_d N_RN_M41_noxref_g ) capacitor c=0.015318f \
 //x=20.465 //y=5.02 //x2=20.39 //y2=6.02
cc_461 ( N_VDD_c_299_n QN ) capacitor c=0.0452986f //x=22.57 //y=7.4 \
 //x2=21.83 //y2=2.22
cc_462 ( N_VDD_c_301_p N_QN_c_1758_n ) capacitor c=0.004515f //x=25.53 //y=7.4 \
 //x2=20.085 //y2=5.155
cc_463 ( N_VDD_c_429_p N_QN_c_1758_n ) capacitor c=4.32228e-19 //x=19.645 \
 //y=7.4 //x2=20.085 //y2=5.155
cc_464 ( N_VDD_c_464_p N_QN_c_1758_n ) capacitor c=4.32228e-19 //x=20.525 \
 //y=7.4 //x2=20.085 //y2=5.155
cc_465 ( N_VDD_M39_noxref_d N_QN_c_1758_n ) capacitor c=0.0115147f //x=19.585 \
 //y=5.02 //x2=20.085 //y2=5.155
cc_466 ( N_VDD_c_298_n N_QN_c_1762_n ) capacitor c=0.00863585f //x=17.76 \
 //y=7.4 //x2=19.375 //y2=5.155
cc_467 ( N_VDD_M38_noxref_s N_QN_c_1762_n ) capacitor c=0.0831083f //x=18.715 \
 //y=5.02 //x2=19.375 //y2=5.155
cc_468 ( N_VDD_c_301_p N_QN_c_1764_n ) capacitor c=0.00448996f //x=25.53 \
 //y=7.4 //x2=20.965 //y2=5.155
cc_469 ( N_VDD_c_464_p N_QN_c_1764_n ) capacitor c=4.32228e-19 //x=20.525 \
 //y=7.4 //x2=20.965 //y2=5.155
cc_470 ( N_VDD_c_477_p N_QN_c_1764_n ) capacitor c=4.32228e-19 //x=21.405 \
 //y=7.4 //x2=20.965 //y2=5.155
cc_471 ( N_VDD_M41_noxref_d N_QN_c_1764_n ) capacitor c=0.0115147f //x=20.465 \
 //y=5.02 //x2=20.965 //y2=5.155
cc_472 ( N_VDD_c_301_p N_QN_c_1768_n ) capacitor c=0.00442621f //x=25.53 \
 //y=7.4 //x2=21.745 //y2=5.155
cc_473 ( N_VDD_c_477_p N_QN_c_1768_n ) capacitor c=7.47666e-19 //x=21.405 \
 //y=7.4 //x2=21.745 //y2=5.155
cc_474 ( N_VDD_c_481_p N_QN_c_1768_n ) capacitor c=0.00198981f //x=22.4 \
 //y=7.4 //x2=21.745 //y2=5.155
cc_475 ( N_VDD_M43_noxref_d N_QN_c_1768_n ) capacitor c=0.0115147f //x=21.345 \
 //y=5.02 //x2=21.745 //y2=5.155
cc_476 ( N_VDD_c_301_p N_QN_c_1745_n ) capacitor c=0.00126216f //x=25.53 \
 //y=7.4 //x2=23.68 //y2=2.08
cc_477 ( N_VDD_c_484_p N_QN_c_1745_n ) capacitor c=2.87813e-19 //x=24.155 \
 //y=7.4 //x2=23.68 //y2=2.08
cc_478 ( N_VDD_c_299_n N_QN_c_1745_n ) capacitor c=0.0160121f //x=22.57 \
 //y=7.4 //x2=23.68 //y2=2.08
cc_479 ( N_VDD_c_484_p N_QN_M44_noxref_g ) capacitor c=0.00726866f //x=24.155 \
 //y=7.4 //x2=23.58 //y2=6.02
cc_480 ( N_VDD_M44_noxref_s N_QN_M44_noxref_g ) capacitor c=0.054195f \
 //x=23.225 //y=5.02 //x2=23.58 //y2=6.02
cc_481 ( N_VDD_c_484_p N_QN_M45_noxref_g ) capacitor c=0.00672952f //x=24.155 \
 //y=7.4 //x2=24.02 //y2=6.02
cc_482 ( N_VDD_M45_noxref_d N_QN_M45_noxref_g ) capacitor c=0.015318f \
 //x=24.095 //y=5.02 //x2=24.02 //y2=6.02
cc_483 ( N_VDD_c_299_n N_QN_c_1779_n ) capacitor c=0.0154093f //x=22.57 \
 //y=7.4 //x2=23.68 //y2=4.7
cc_484 ( N_VDD_c_301_p N_QN_M38_noxref_d ) capacitor c=0.00285091f //x=25.53 \
 //y=7.4 //x2=19.145 //y2=5.02
cc_485 ( N_VDD_c_429_p N_QN_M38_noxref_d ) capacitor c=0.0141016f //x=19.645 \
 //y=7.4 //x2=19.145 //y2=5.02
cc_486 ( N_VDD_M39_noxref_d N_QN_M38_noxref_d ) capacitor c=0.0664752f \
 //x=19.585 //y=5.02 //x2=19.145 //y2=5.02
cc_487 ( N_VDD_c_301_p N_QN_M40_noxref_d ) capacitor c=0.00285091f //x=25.53 \
 //y=7.4 //x2=20.025 //y2=5.02
cc_488 ( N_VDD_c_464_p N_QN_M40_noxref_d ) capacitor c=0.0141016f //x=20.525 \
 //y=7.4 //x2=20.025 //y2=5.02
cc_489 ( N_VDD_c_299_n N_QN_M40_noxref_d ) capacitor c=4.9285e-19 //x=22.57 \
 //y=7.4 //x2=20.025 //y2=5.02
cc_490 ( N_VDD_M38_noxref_s N_QN_M40_noxref_d ) capacitor c=0.00130656f \
 //x=18.715 //y=5.02 //x2=20.025 //y2=5.02
cc_491 ( N_VDD_M39_noxref_d N_QN_M40_noxref_d ) capacitor c=0.0664752f \
 //x=19.585 //y=5.02 //x2=20.025 //y2=5.02
cc_492 ( N_VDD_M41_noxref_d N_QN_M40_noxref_d ) capacitor c=0.0664752f \
 //x=20.465 //y=5.02 //x2=20.025 //y2=5.02
cc_493 ( N_VDD_c_301_p N_QN_M42_noxref_d ) capacitor c=0.00285091f //x=25.53 \
 //y=7.4 //x2=20.905 //y2=5.02
cc_494 ( N_VDD_c_477_p N_QN_M42_noxref_d ) capacitor c=0.0138051f //x=21.405 \
 //y=7.4 //x2=20.905 //y2=5.02
cc_495 ( N_VDD_c_299_n N_QN_M42_noxref_d ) capacitor c=0.00939849f //x=22.57 \
 //y=7.4 //x2=20.905 //y2=5.02
cc_496 ( N_VDD_M41_noxref_d N_QN_M42_noxref_d ) capacitor c=0.0664752f \
 //x=20.465 //y=5.02 //x2=20.905 //y2=5.02
cc_497 ( N_VDD_M43_noxref_d N_QN_M42_noxref_d ) capacitor c=0.0664752f \
 //x=21.345 //y=5.02 //x2=20.905 //y2=5.02
cc_498 ( N_VDD_M44_noxref_s N_QN_M42_noxref_d ) capacitor c=4.52683e-19 \
 //x=23.225 //y=5.02 //x2=20.905 //y2=5.02
cc_499 ( N_VDD_c_301_p N_noxref_9_c_1895_n ) capacitor c=0.0425735f //x=25.53 \
 //y=7.4 //x2=11.355 //y2=4.07
cc_500 ( N_VDD_c_405_p N_noxref_9_c_1895_n ) capacitor c=0.00113322f //x=1.885 \
 //y=7.4 //x2=11.355 //y2=4.07
cc_501 ( N_VDD_c_295_n N_noxref_9_c_1895_n ) capacitor c=0.0140578f //x=4.81 \
 //y=7.4 //x2=11.355 //y2=4.07
cc_502 ( N_VDD_c_296_n N_noxref_9_c_1895_n ) capacitor c=0.0140578f //x=9.62 \
 //y=7.4 //x2=11.355 //y2=4.07
cc_503 ( N_VDD_c_301_p N_noxref_9_c_1896_n ) capacitor c=0.00189266f //x=25.53 \
 //y=7.4 //x2=1.225 //y2=4.07
cc_504 ( N_VDD_c_293_n N_noxref_9_c_1896_n ) capacitor c=0.0017219f //x=0.74 \
 //y=7.4 //x2=1.225 //y2=4.07
cc_505 ( N_VDD_M16_noxref_s N_noxref_9_c_1896_n ) capacitor c=0.00128242f \
 //x=0.955 //y=5.02 //x2=1.225 //y2=4.07
cc_506 ( N_VDD_c_301_p N_noxref_9_c_1922_n ) capacitor c=0.0256485f //x=25.53 \
 //y=7.4 //x2=16.905 //y2=4.07
cc_507 ( N_VDD_c_297_n N_noxref_9_c_1922_n ) capacitor c=0.0140578f //x=12.95 \
 //y=7.4 //x2=16.905 //y2=4.07
cc_508 ( N_VDD_c_301_p N_noxref_9_c_1897_n ) capacitor c=0.0509002f //x=25.53 \
 //y=7.4 //x2=24.305 //y2=4.07
cc_509 ( N_VDD_c_516_p N_noxref_9_c_1897_n ) capacitor c=0.0016229f //x=17.59 \
 //y=7.4 //x2=24.305 //y2=4.07
cc_510 ( N_VDD_c_517_p N_noxref_9_c_1897_n ) capacitor c=0.0027159f //x=18.765 \
 //y=7.4 //x2=24.305 //y2=4.07
cc_511 ( N_VDD_c_429_p N_noxref_9_c_1897_n ) capacitor c=0.00113459f \
 //x=19.645 //y=7.4 //x2=24.305 //y2=4.07
cc_512 ( N_VDD_c_481_p N_noxref_9_c_1897_n ) capacitor c=0.00214241f //x=22.4 \
 //y=7.4 //x2=24.305 //y2=4.07
cc_513 ( N_VDD_c_520_p N_noxref_9_c_1897_n ) capacitor c=0.00172186f \
 //x=23.275 //y=7.4 //x2=24.305 //y2=4.07
cc_514 ( N_VDD_c_484_p N_noxref_9_c_1897_n ) capacitor c=6.61469e-19 \
 //x=24.155 //y=7.4 //x2=24.305 //y2=4.07
cc_515 ( N_VDD_c_298_n N_noxref_9_c_1897_n ) capacitor c=0.0269494f //x=17.76 \
 //y=7.4 //x2=24.305 //y2=4.07
cc_516 ( N_VDD_c_299_n N_noxref_9_c_1897_n ) capacitor c=0.0269494f //x=22.57 \
 //y=7.4 //x2=24.305 //y2=4.07
cc_517 ( N_VDD_M38_noxref_s N_noxref_9_c_1897_n ) capacitor c=0.00122826f \
 //x=18.715 //y=5.02 //x2=24.305 //y2=4.07
cc_518 ( N_VDD_M44_noxref_s N_noxref_9_c_1897_n ) capacitor c=0.00363031f \
 //x=23.225 //y=5.02 //x2=24.305 //y2=4.07
cc_519 ( N_VDD_c_301_p N_noxref_9_c_1935_n ) capacitor c=0.00175338f //x=25.53 \
 //y=7.4 //x2=17.135 //y2=4.07
cc_520 ( N_VDD_c_516_p N_noxref_9_c_1935_n ) capacitor c=5.20513e-19 //x=17.59 \
 //y=7.4 //x2=17.135 //y2=4.07
cc_521 ( N_VDD_c_298_n N_noxref_9_c_1935_n ) capacitor c=0.00104972f //x=17.76 \
 //y=7.4 //x2=17.135 //y2=4.07
cc_522 ( N_VDD_c_301_p N_noxref_9_c_1898_n ) capacitor c=9.2251e-19 //x=25.53 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_523 ( N_VDD_c_293_n N_noxref_9_c_1898_n ) capacitor c=0.0159723f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_524 ( N_VDD_M16_noxref_s N_noxref_9_c_1898_n ) capacitor c=0.0122951f \
 //x=0.955 //y=5.02 //x2=1.11 //y2=2.08
cc_525 ( N_VDD_c_296_n N_noxref_9_c_1899_n ) capacitor c=4.57806e-19 //x=9.62 \
 //y=7.4 //x2=11.47 //y2=2.08
cc_526 ( N_VDD_c_297_n N_noxref_9_c_1899_n ) capacitor c=3.21957e-19 //x=12.95 \
 //y=7.4 //x2=11.47 //y2=2.08
cc_527 ( N_VDD_c_301_p N_noxref_9_c_1943_n ) capacitor c=0.00444751f //x=25.53 \
 //y=7.4 //x2=15.275 //y2=5.155
cc_528 ( N_VDD_c_357_p N_noxref_9_c_1943_n ) capacitor c=4.31931e-19 \
 //x=14.835 //y=7.4 //x2=15.275 //y2=5.155
cc_529 ( N_VDD_c_400_p N_noxref_9_c_1943_n ) capacitor c=4.31906e-19 \
 //x=15.715 //y=7.4 //x2=15.275 //y2=5.155
cc_530 ( N_VDD_M33_noxref_d N_noxref_9_c_1943_n ) capacitor c=0.0112985f \
 //x=14.775 //y=5.02 //x2=15.275 //y2=5.155
cc_531 ( N_VDD_c_297_n N_noxref_9_c_1947_n ) capacitor c=0.00863585f //x=12.95 \
 //y=7.4 //x2=14.565 //y2=5.155
cc_532 ( N_VDD_M32_noxref_s N_noxref_9_c_1947_n ) capacitor c=0.0831083f \
 //x=13.905 //y=5.02 //x2=14.565 //y2=5.155
cc_533 ( N_VDD_c_301_p N_noxref_9_c_1949_n ) capacitor c=0.00448996f //x=25.53 \
 //y=7.4 //x2=16.155 //y2=5.155
cc_534 ( N_VDD_c_400_p N_noxref_9_c_1949_n ) capacitor c=4.32228e-19 \
 //x=15.715 //y=7.4 //x2=16.155 //y2=5.155
cc_535 ( N_VDD_c_460_p N_noxref_9_c_1949_n ) capacitor c=4.32228e-19 \
 //x=16.595 //y=7.4 //x2=16.155 //y2=5.155
cc_536 ( N_VDD_M35_noxref_d N_noxref_9_c_1949_n ) capacitor c=0.0115147f \
 //x=15.655 //y=5.02 //x2=16.155 //y2=5.155
cc_537 ( N_VDD_c_301_p N_noxref_9_c_1953_n ) capacitor c=0.00442469f //x=25.53 \
 //y=7.4 //x2=16.935 //y2=5.155
cc_538 ( N_VDD_c_460_p N_noxref_9_c_1953_n ) capacitor c=7.47666e-19 \
 //x=16.595 //y=7.4 //x2=16.935 //y2=5.155
cc_539 ( N_VDD_c_516_p N_noxref_9_c_1953_n ) capacitor c=0.00198959f //x=17.59 \
 //y=7.4 //x2=16.935 //y2=5.155
cc_540 ( N_VDD_M37_noxref_d N_noxref_9_c_1953_n ) capacitor c=0.0115147f \
 //x=16.535 //y=5.02 //x2=16.935 //y2=5.155
cc_541 ( N_VDD_c_298_n N_noxref_9_c_1957_n ) capacitor c=0.0452313f //x=17.76 \
 //y=7.4 //x2=17.02 //y2=4.07
cc_542 ( N_VDD_c_294_n N_noxref_9_c_1902_n ) capacitor c=6.61994e-19 //x=25.53 \
 //y=7.4 //x2=24.42 //y2=2.08
cc_543 ( N_VDD_c_299_n N_noxref_9_c_1902_n ) capacitor c=6.2696e-19 //x=22.57 \
 //y=7.4 //x2=24.42 //y2=2.08
cc_544 ( N_VDD_c_405_p N_noxref_9_M16_noxref_g ) capacitor c=0.00749687f \
 //x=1.885 //y=7.4 //x2=1.31 //y2=6.02
cc_545 ( N_VDD_M16_noxref_s N_noxref_9_M16_noxref_g ) capacitor c=0.0477201f \
 //x=0.955 //y=5.02 //x2=1.31 //y2=6.02
cc_546 ( N_VDD_c_405_p N_noxref_9_M17_noxref_g ) capacitor c=0.00675175f \
 //x=1.885 //y=7.4 //x2=1.75 //y2=6.02
cc_547 ( N_VDD_M17_noxref_d N_noxref_9_M17_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=1.75 //y2=6.02
cc_548 ( N_VDD_c_345_p N_noxref_9_M30_noxref_g ) capacitor c=0.00673971f \
 //x=12.085 //y=7.4 //x2=11.51 //y2=6.02
cc_549 ( N_VDD_M29_noxref_d N_noxref_9_M30_noxref_g ) capacitor c=0.015318f \
 //x=11.145 //y=5.02 //x2=11.51 //y2=6.02
cc_550 ( N_VDD_c_345_p N_noxref_9_M31_noxref_g ) capacitor c=0.00672952f \
 //x=12.085 //y=7.4 //x2=11.95 //y2=6.02
cc_551 ( N_VDD_c_297_n N_noxref_9_M31_noxref_g ) capacitor c=0.00928743f \
 //x=12.95 //y=7.4 //x2=11.95 //y2=6.02
cc_552 ( N_VDD_M31_noxref_d N_noxref_9_M31_noxref_g ) capacitor c=0.0430452f \
 //x=12.025 //y=5.02 //x2=11.95 //y2=6.02
cc_553 ( N_VDD_c_560_p N_noxref_9_M46_noxref_g ) capacitor c=0.00673971f \
 //x=25.035 //y=7.4 //x2=24.46 //y2=6.02
cc_554 ( N_VDD_M45_noxref_d N_noxref_9_M46_noxref_g ) capacitor c=0.015318f \
 //x=24.095 //y=5.02 //x2=24.46 //y2=6.02
cc_555 ( N_VDD_c_560_p N_noxref_9_M47_noxref_g ) capacitor c=0.00672952f \
 //x=25.035 //y=7.4 //x2=24.9 //y2=6.02
cc_556 ( N_VDD_c_294_n N_noxref_9_M47_noxref_g ) capacitor c=0.024326f \
 //x=25.53 //y=7.4 //x2=24.9 //y2=6.02
cc_557 ( N_VDD_M47_noxref_d N_noxref_9_M47_noxref_g ) capacitor c=0.0430452f \
 //x=24.975 //y=5.02 //x2=24.9 //y2=6.02
cc_558 ( N_VDD_c_293_n N_noxref_9_c_1974_n ) capacitor c=0.00757682f //x=0.74 \
 //y=7.4 //x2=1.385 //y2=4.79
cc_559 ( N_VDD_M16_noxref_s N_noxref_9_c_1974_n ) capacitor c=0.00445117f \
 //x=0.955 //y=5.02 //x2=1.385 //y2=4.79
cc_560 ( N_VDD_c_301_p N_noxref_9_M32_noxref_d ) capacitor c=0.00275235f \
 //x=25.53 //y=7.4 //x2=14.335 //y2=5.02
cc_561 ( N_VDD_c_357_p N_noxref_9_M32_noxref_d ) capacitor c=0.014035f \
 //x=14.835 //y=7.4 //x2=14.335 //y2=5.02
cc_562 ( N_VDD_M33_noxref_d N_noxref_9_M32_noxref_d ) capacitor c=0.0664752f \
 //x=14.775 //y=5.02 //x2=14.335 //y2=5.02
cc_563 ( N_VDD_c_301_p N_noxref_9_M34_noxref_d ) capacitor c=0.00282723f \
 //x=25.53 //y=7.4 //x2=15.215 //y2=5.02
cc_564 ( N_VDD_c_400_p N_noxref_9_M34_noxref_d ) capacitor c=0.0140856f \
 //x=15.715 //y=7.4 //x2=15.215 //y2=5.02
cc_565 ( N_VDD_c_298_n N_noxref_9_M34_noxref_d ) capacitor c=4.9285e-19 \
 //x=17.76 //y=7.4 //x2=15.215 //y2=5.02
cc_566 ( N_VDD_M32_noxref_s N_noxref_9_M34_noxref_d ) capacitor c=0.00130656f \
 //x=13.905 //y=5.02 //x2=15.215 //y2=5.02
cc_567 ( N_VDD_M33_noxref_d N_noxref_9_M34_noxref_d ) capacitor c=0.0664752f \
 //x=14.775 //y=5.02 //x2=15.215 //y2=5.02
cc_568 ( N_VDD_M35_noxref_d N_noxref_9_M34_noxref_d ) capacitor c=0.0664752f \
 //x=15.655 //y=5.02 //x2=15.215 //y2=5.02
cc_569 ( N_VDD_c_301_p N_noxref_9_M36_noxref_d ) capacitor c=0.00285091f \
 //x=25.53 //y=7.4 //x2=16.095 //y2=5.02
cc_570 ( N_VDD_c_460_p N_noxref_9_M36_noxref_d ) capacitor c=0.0138051f \
 //x=16.595 //y=7.4 //x2=16.095 //y2=5.02
cc_571 ( N_VDD_c_298_n N_noxref_9_M36_noxref_d ) capacitor c=0.00939849f \
 //x=17.76 //y=7.4 //x2=16.095 //y2=5.02
cc_572 ( N_VDD_M35_noxref_d N_noxref_9_M36_noxref_d ) capacitor c=0.0664752f \
 //x=15.655 //y=5.02 //x2=16.095 //y2=5.02
cc_573 ( N_VDD_M37_noxref_d N_noxref_9_M36_noxref_d ) capacitor c=0.0664752f \
 //x=16.535 //y=5.02 //x2=16.095 //y2=5.02
cc_574 ( N_VDD_M38_noxref_s N_noxref_9_M36_noxref_d ) capacitor c=3.57641e-19 \
 //x=18.715 //y=5.02 //x2=16.095 //y2=5.02
cc_575 ( N_VDD_c_301_p N_noxref_10_c_2279_n ) capacitor c=0.0163609f //x=25.53 \
 //y=7.4 //x2=25.045 //y2=3.7
cc_576 ( N_VDD_M47_noxref_d N_noxref_10_c_2279_n ) capacitor c=4.05358e-19 \
 //x=24.975 //y=5.02 //x2=25.045 //y2=3.7
cc_577 ( N_VDD_c_299_n N_noxref_10_c_2281_n ) capacitor c=8.5347e-19 //x=22.57 \
 //y=7.4 //x2=21.09 //y2=2.08
cc_578 ( N_VDD_c_301_p N_noxref_10_c_2290_n ) capacitor c=0.00459955f \
 //x=25.53 //y=7.4 //x2=24.595 //y2=5.2
cc_579 ( N_VDD_c_484_p N_noxref_10_c_2290_n ) capacitor c=4.48705e-19 \
 //x=24.155 //y=7.4 //x2=24.595 //y2=5.2
cc_580 ( N_VDD_c_560_p N_noxref_10_c_2290_n ) capacitor c=4.48693e-19 \
 //x=25.035 //y=7.4 //x2=24.595 //y2=5.2
cc_581 ( N_VDD_M45_noxref_d N_noxref_10_c_2290_n ) capacitor c=0.01269f \
 //x=24.095 //y=5.02 //x2=24.595 //y2=5.2
cc_582 ( N_VDD_c_299_n N_noxref_10_c_2294_n ) capacitor c=0.00985474f \
 //x=22.57 //y=7.4 //x2=23.885 //y2=5.2
cc_583 ( N_VDD_M44_noxref_s N_noxref_10_c_2294_n ) capacitor c=0.087833f \
 //x=23.225 //y=5.02 //x2=23.885 //y2=5.2
cc_584 ( N_VDD_c_301_p N_noxref_10_c_2296_n ) capacitor c=0.00311875f \
 //x=25.53 //y=7.4 //x2=25.075 //y2=5.2
cc_585 ( N_VDD_c_560_p N_noxref_10_c_2296_n ) capacitor c=7.21492e-19 \
 //x=25.035 //y=7.4 //x2=25.075 //y2=5.2
cc_586 ( N_VDD_M47_noxref_d N_noxref_10_c_2296_n ) capacitor c=0.0163364f \
 //x=24.975 //y=5.02 //x2=25.075 //y2=5.2
cc_587 ( N_VDD_c_294_n N_noxref_10_c_2283_n ) capacitor c=0.0466813f //x=25.53 \
 //y=7.4 //x2=25.16 //y2=3.7
cc_588 ( N_VDD_c_299_n N_noxref_10_c_2283_n ) capacitor c=0.00151618f \
 //x=22.57 //y=7.4 //x2=25.16 //y2=3.7
cc_589 ( N_VDD_c_477_p N_noxref_10_M42_noxref_g ) capacitor c=0.00675175f \
 //x=21.405 //y=7.4 //x2=20.83 //y2=6.02
cc_590 ( N_VDD_M41_noxref_d N_noxref_10_M42_noxref_g ) capacitor c=0.015318f \
 //x=20.465 //y=5.02 //x2=20.83 //y2=6.02
cc_591 ( N_VDD_c_477_p N_noxref_10_M43_noxref_g ) capacitor c=0.00675379f \
 //x=21.405 //y=7.4 //x2=21.27 //y2=6.02
cc_592 ( N_VDD_M43_noxref_d N_noxref_10_M43_noxref_g ) capacitor c=0.0394719f \
 //x=21.345 //y=5.02 //x2=21.27 //y2=6.02
cc_593 ( N_VDD_c_301_p N_noxref_10_M44_noxref_d ) capacitor c=0.00285083f \
 //x=25.53 //y=7.4 //x2=23.655 //y2=5.02
cc_594 ( N_VDD_c_484_p N_noxref_10_M44_noxref_d ) capacitor c=0.0140984f \
 //x=24.155 //y=7.4 //x2=23.655 //y2=5.02
cc_595 ( N_VDD_c_294_n N_noxref_10_M44_noxref_d ) capacitor c=6.94454e-19 \
 //x=25.53 //y=7.4 //x2=23.655 //y2=5.02
cc_596 ( N_VDD_M45_noxref_d N_noxref_10_M44_noxref_d ) capacitor c=0.0664752f \
 //x=24.095 //y=5.02 //x2=23.655 //y2=5.02
cc_597 ( N_VDD_c_301_p N_noxref_10_M46_noxref_d ) capacitor c=0.00294217f \
 //x=25.53 //y=7.4 //x2=24.535 //y2=5.02
cc_598 ( N_VDD_c_560_p N_noxref_10_M46_noxref_d ) capacitor c=0.0138379f \
 //x=25.035 //y=7.4 //x2=24.535 //y2=5.02
cc_599 ( N_VDD_c_294_n N_noxref_10_M46_noxref_d ) capacitor c=0.0123189f \
 //x=25.53 //y=7.4 //x2=24.535 //y2=5.02
cc_600 ( N_VDD_M44_noxref_s N_noxref_10_M46_noxref_d ) capacitor c=0.00111971f \
 //x=23.225 //y=5.02 //x2=24.535 //y2=5.02
cc_601 ( N_VDD_M45_noxref_d N_noxref_10_M46_noxref_d ) capacitor c=0.0664752f \
 //x=24.095 //y=5.02 //x2=24.535 //y2=5.02
cc_602 ( N_VDD_M47_noxref_d N_noxref_10_M46_noxref_d ) capacitor c=0.0664752f \
 //x=24.975 //y=5.02 //x2=24.535 //y2=5.02
cc_603 ( N_VDD_c_301_p N_D_c_2523_n ) capacitor c=2.03486e-19 //x=25.53 \
 //y=7.4 //x2=7.03 //y2=2.08
cc_604 ( N_VDD_c_295_n N_D_c_2523_n ) capacitor c=5.89117e-19 //x=4.81 //y=7.4 \
 //x2=7.03 //y2=2.08
cc_605 ( N_VDD_c_303_p N_D_M24_noxref_g ) capacitor c=0.00676195f //x=7.575 \
 //y=7.4 //x2=7 //y2=6.02
cc_606 ( N_VDD_M23_noxref_d N_D_M24_noxref_g ) capacitor c=0.015318f //x=6.635 \
 //y=5.02 //x2=7 //y2=6.02
cc_607 ( N_VDD_c_303_p N_D_M25_noxref_g ) capacitor c=0.00675175f //x=7.575 \
 //y=7.4 //x2=7.44 //y2=6.02
cc_608 ( N_VDD_M25_noxref_d N_D_M25_noxref_g ) capacitor c=0.015318f //x=7.515 \
 //y=5.02 //x2=7.44 //y2=6.02
cc_609 ( N_noxref_3_c_621_n N_noxref_4_c_910_n ) capacitor c=0.011463f \
 //x=10.615 //y=3.33 //x2=12.325 //y2=3.33
cc_610 ( N_noxref_3_M29_noxref_g N_noxref_4_c_879_n ) capacitor c=0.0169521f \
 //x=11.07 //y=6.02 //x2=11.645 //y2=5.2
cc_611 ( N_noxref_3_c_624_n N_noxref_4_c_883_n ) capacitor c=0.00539951f \
 //x=10.73 //y=2.08 //x2=10.935 //y2=5.2
cc_612 ( N_noxref_3_M28_noxref_g N_noxref_4_c_883_n ) capacitor c=0.0177326f \
 //x=10.63 //y=6.02 //x2=10.935 //y2=5.2
cc_613 ( N_noxref_3_c_663_n N_noxref_4_c_883_n ) capacitor c=0.00581252f \
 //x=10.73 //y=4.7 //x2=10.935 //y2=5.2
cc_614 ( N_noxref_3_c_651_n N_noxref_4_c_864_n ) capacitor c=3.52729e-19 \
 //x=8.88 //y=3.33 //x2=12.21 //y2=3.33
cc_615 ( N_noxref_3_c_624_n N_noxref_4_c_864_n ) capacitor c=0.00292364f \
 //x=10.73 //y=2.08 //x2=12.21 //y2=3.33
cc_616 ( N_noxref_3_M29_noxref_g N_noxref_4_M28_noxref_d ) capacitor \
 c=0.0173476f //x=11.07 //y=6.02 //x2=10.705 //y2=5.02
cc_617 ( N_noxref_3_c_616_n N_CLK_c_1011_n ) capacitor c=0.00360213f //x=8.765 \
 //y=3.33 //x2=15.055 //y2=4.44
cc_618 ( N_noxref_3_c_620_n N_CLK_c_1011_n ) capacitor c=4.49102e-19 //x=3.445 \
 //y=3.33 //x2=15.055 //y2=4.44
cc_619 ( N_noxref_3_c_622_n N_CLK_c_1011_n ) capacitor c=0.0200057f //x=3.33 \
 //y=2.08 //x2=15.055 //y2=4.44
cc_620 ( N_noxref_3_c_637_n N_CLK_c_1011_n ) capacitor c=0.032141f //x=7.135 \
 //y=5.155 //x2=15.055 //y2=4.44
cc_621 ( N_noxref_3_c_641_n N_CLK_c_1011_n ) capacitor c=0.0230136f //x=6.425 \
 //y=5.155 //x2=15.055 //y2=4.44
cc_622 ( N_noxref_3_c_647_n N_CLK_c_1011_n ) capacitor c=0.0183122f //x=8.795 \
 //y=5.155 //x2=15.055 //y2=4.44
cc_623 ( N_noxref_3_c_651_n N_CLK_c_1011_n ) capacitor c=0.0210274f //x=8.88 \
 //y=3.33 //x2=15.055 //y2=4.44
cc_624 ( N_noxref_3_c_624_n N_CLK_c_1011_n ) capacitor c=0.0198304f //x=10.73 \
 //y=2.08 //x2=15.055 //y2=4.44
cc_625 ( N_noxref_3_c_695_p N_CLK_c_1011_n ) capacitor c=0.0111881f //x=3.33 \
 //y=4.7 //x2=15.055 //y2=4.44
cc_626 ( N_noxref_3_c_663_n N_CLK_c_1011_n ) capacitor c=0.0107057f //x=10.73 \
 //y=4.7 //x2=15.055 //y2=4.44
cc_627 ( N_noxref_3_c_622_n N_CLK_c_1028_n ) capacitor c=0.00153281f //x=3.33 \
 //y=2.08 //x2=2.335 //y2=4.44
cc_628 ( N_noxref_3_c_620_n N_CLK_c_1009_n ) capacitor c=0.00526349f //x=3.445 \
 //y=3.33 //x2=2.22 //y2=2.08
cc_629 ( N_noxref_3_c_622_n N_CLK_c_1009_n ) capacitor c=0.0511464f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_630 ( N_noxref_3_c_700_p N_CLK_c_1009_n ) capacitor c=0.00228632f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_631 ( N_noxref_3_c_695_p N_CLK_c_1009_n ) capacitor c=0.00218014f //x=3.33 \
 //y=4.7 //x2=2.22 //y2=2.08
cc_632 ( N_noxref_3_M20_noxref_g N_CLK_M18_noxref_g ) capacitor c=0.0101598f \
 //x=3.07 //y=6.02 //x2=2.19 //y2=6.02
cc_633 ( N_noxref_3_M20_noxref_g N_CLK_M19_noxref_g ) capacitor c=0.0602553f \
 //x=3.07 //y=6.02 //x2=2.63 //y2=6.02
cc_634 ( N_noxref_3_M21_noxref_g N_CLK_M19_noxref_g ) capacitor c=0.0101598f \
 //x=3.51 //y=6.02 //x2=2.63 //y2=6.02
cc_635 ( N_noxref_3_c_705_p N_CLK_c_1059_n ) capacitor c=0.00456962f //x=3.32 \
 //y=0.915 //x2=2.31 //y2=0.91
cc_636 ( N_noxref_3_c_706_p N_CLK_c_1060_n ) capacitor c=0.00438372f //x=3.32 \
 //y=1.26 //x2=2.31 //y2=1.22
cc_637 ( N_noxref_3_c_707_p N_CLK_c_1061_n ) capacitor c=0.00438372f //x=3.32 \
 //y=1.57 //x2=2.31 //y2=1.45
cc_638 ( N_noxref_3_c_622_n N_CLK_c_1062_n ) capacitor c=0.0023343f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_639 ( N_noxref_3_c_700_p N_CLK_c_1062_n ) capacitor c=0.00933826f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_640 ( N_noxref_3_c_710_p N_CLK_c_1062_n ) capacitor c=0.00438372f //x=3.33 \
 //y=1.915 //x2=2.31 //y2=1.915
cc_641 ( N_noxref_3_c_695_p N_CLK_c_1065_n ) capacitor c=0.0611812f //x=3.33 \
 //y=4.7 //x2=2.555 //y2=4.79
cc_642 ( N_noxref_3_c_622_n N_CLK_c_1066_n ) capacitor c=0.00142741f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=4.7
cc_643 ( N_noxref_3_c_695_p N_CLK_c_1066_n ) capacitor c=0.00487508f //x=3.33 \
 //y=4.7 //x2=2.22 //y2=4.7
cc_644 ( N_noxref_3_c_616_n N_noxref_6_c_1297_n ) capacitor c=0.146539f \
 //x=8.765 //y=3.33 //x2=5.805 //y2=3.7
cc_645 ( N_noxref_3_c_616_n N_noxref_6_c_1298_n ) capacitor c=0.0294746f \
 //x=8.765 //y=3.33 //x2=4.185 //y2=3.7
cc_646 ( N_noxref_3_c_622_n N_noxref_6_c_1298_n ) capacitor c=0.00687545f \
 //x=3.33 //y=2.08 //x2=4.185 //y2=3.7
cc_647 ( N_noxref_3_c_616_n N_noxref_6_c_1224_n ) capacitor c=0.238435f \
 //x=8.765 //y=3.33 //x2=18.755 //y2=3.7
cc_648 ( N_noxref_3_c_621_n N_noxref_6_c_1224_n ) capacitor c=0.175734f \
 //x=10.615 //y=3.33 //x2=18.755 //y2=3.7
cc_649 ( N_noxref_3_c_719_p N_noxref_6_c_1224_n ) capacitor c=0.0268386f \
 //x=8.995 //y=3.33 //x2=18.755 //y2=3.7
cc_650 ( N_noxref_3_c_651_n N_noxref_6_c_1224_n ) capacitor c=0.0206044f \
 //x=8.88 //y=3.33 //x2=18.755 //y2=3.7
cc_651 ( N_noxref_3_c_624_n N_noxref_6_c_1224_n ) capacitor c=0.0205831f \
 //x=10.73 //y=2.08 //x2=18.755 //y2=3.7
cc_652 ( N_noxref_3_c_616_n N_noxref_6_c_1305_n ) capacitor c=0.0266966f \
 //x=8.765 //y=3.33 //x2=6.035 //y2=3.7
cc_653 ( N_noxref_3_M20_noxref_g N_noxref_6_c_1255_n ) capacitor c=0.01736f \
 //x=3.07 //y=6.02 //x2=3.205 //y2=5.155
cc_654 ( N_noxref_3_c_641_n N_noxref_6_c_1259_n ) capacitor c=3.10026e-19 \
 //x=6.425 //y=5.155 //x2=3.985 //y2=5.155
cc_655 ( N_noxref_3_M21_noxref_g N_noxref_6_c_1259_n ) capacitor c=0.0194981f \
 //x=3.51 //y=6.02 //x2=3.985 //y2=5.155
cc_656 ( N_noxref_3_c_695_p N_noxref_6_c_1259_n ) capacitor c=0.00201851f \
 //x=3.33 //y=4.7 //x2=3.985 //y2=5.155
cc_657 ( N_noxref_3_c_727_p N_noxref_6_c_1225_n ) capacitor c=0.00359704f \
 //x=3.695 //y=1.415 //x2=3.985 //y2=1.665
cc_658 ( N_noxref_3_c_728_p N_noxref_6_c_1225_n ) capacitor c=0.00457401f \
 //x=3.85 //y=1.26 //x2=3.985 //y2=1.665
cc_659 ( N_noxref_3_c_616_n N_noxref_6_c_1312_n ) capacitor c=0.00628992f \
 //x=8.765 //y=3.33 //x2=3.67 //y2=1.665
cc_660 ( N_noxref_3_c_616_n N_noxref_6_c_1263_n ) capacitor c=0.0260398f \
 //x=8.765 //y=3.33 //x2=4.07 //y2=3.7
cc_661 ( N_noxref_3_c_620_n N_noxref_6_c_1263_n ) capacitor c=0.00179385f \
 //x=3.445 //y=3.33 //x2=4.07 //y2=3.7
cc_662 ( N_noxref_3_c_622_n N_noxref_6_c_1263_n ) capacitor c=0.0831612f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_663 ( N_noxref_3_c_700_p N_noxref_6_c_1263_n ) capacitor c=0.00877984f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_664 ( N_noxref_3_c_710_p N_noxref_6_c_1263_n ) capacitor c=0.00283672f \
 //x=3.33 //y=1.915 //x2=4.07 //y2=3.7
cc_665 ( N_noxref_3_c_695_p N_noxref_6_c_1263_n ) capacitor c=0.013693f \
 //x=3.33 //y=4.7 //x2=4.07 //y2=3.7
cc_666 ( N_noxref_3_c_616_n N_noxref_6_c_1226_n ) capacitor c=0.0268062f \
 //x=8.765 //y=3.33 //x2=5.92 //y2=2.08
cc_667 ( N_noxref_3_c_622_n N_noxref_6_c_1226_n ) capacitor c=9.66956e-19 \
 //x=3.33 //y=2.08 //x2=5.92 //y2=2.08
cc_668 ( N_noxref_3_c_622_n N_noxref_6_c_1321_n ) capacitor c=0.0171303f \
 //x=3.33 //y=2.08 //x2=3.29 //y2=5.155
cc_669 ( N_noxref_3_c_695_p N_noxref_6_c_1321_n ) capacitor c=0.00475601f \
 //x=3.33 //y=4.7 //x2=3.29 //y2=5.155
cc_670 ( N_noxref_3_c_641_n N_noxref_6_M22_noxref_g ) capacitor c=0.0213876f \
 //x=6.425 //y=5.155 //x2=6.12 //y2=6.02
cc_671 ( N_noxref_3_c_637_n N_noxref_6_M23_noxref_g ) capacitor c=0.0168349f \
 //x=7.135 //y=5.155 //x2=6.56 //y2=6.02
cc_672 ( N_noxref_3_M22_noxref_d N_noxref_6_M23_noxref_g ) capacitor \
 c=0.0180032f //x=6.195 //y=5.02 //x2=6.56 //y2=6.02
cc_673 ( N_noxref_3_c_641_n N_noxref_6_c_1326_n ) capacitor c=0.00428486f \
 //x=6.425 //y=5.155 //x2=6.485 //y2=4.79
cc_674 ( N_noxref_3_c_705_p N_noxref_6_M2_noxref_d ) capacitor c=0.00217566f \
 //x=3.32 //y=0.915 //x2=3.395 //y2=0.915
cc_675 ( N_noxref_3_c_706_p N_noxref_6_M2_noxref_d ) capacitor c=0.0034598f \
 //x=3.32 //y=1.26 //x2=3.395 //y2=0.915
cc_676 ( N_noxref_3_c_707_p N_noxref_6_M2_noxref_d ) capacitor c=0.00544291f \
 //x=3.32 //y=1.57 //x2=3.395 //y2=0.915
cc_677 ( N_noxref_3_c_747_p N_noxref_6_M2_noxref_d ) capacitor c=0.00241102f \
 //x=3.695 //y=0.76 //x2=3.395 //y2=0.915
cc_678 ( N_noxref_3_c_727_p N_noxref_6_M2_noxref_d ) capacitor c=0.0140297f \
 //x=3.695 //y=1.415 //x2=3.395 //y2=0.915
cc_679 ( N_noxref_3_c_749_p N_noxref_6_M2_noxref_d ) capacitor c=0.00219619f \
 //x=3.85 //y=0.915 //x2=3.395 //y2=0.915
cc_680 ( N_noxref_3_c_728_p N_noxref_6_M2_noxref_d ) capacitor c=0.00603828f \
 //x=3.85 //y=1.26 //x2=3.395 //y2=0.915
cc_681 ( N_noxref_3_c_710_p N_noxref_6_M2_noxref_d ) capacitor c=0.00661782f \
 //x=3.33 //y=1.915 //x2=3.395 //y2=0.915
cc_682 ( N_noxref_3_M20_noxref_g N_noxref_6_M20_noxref_d ) capacitor \
 c=0.0180032f //x=3.07 //y=6.02 //x2=3.145 //y2=5.02
cc_683 ( N_noxref_3_M21_noxref_g N_noxref_6_M20_noxref_d ) capacitor \
 c=0.0194246f //x=3.51 //y=6.02 //x2=3.145 //y2=5.02
cc_684 ( N_noxref_3_c_616_n N_RN_c_1470_n ) capacitor c=0.0140941f //x=8.765 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_685 ( N_noxref_3_c_621_n N_RN_c_1470_n ) capacitor c=0.0541047f //x=10.615 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_686 ( N_noxref_3_c_719_p N_RN_c_1470_n ) capacitor c=0.00680007f //x=8.995 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_687 ( N_noxref_3_c_757_p N_RN_c_1470_n ) capacitor c=0.016327f //x=8.48 \
 //y=1.665 //x2=16.165 //y2=2.22
cc_688 ( N_noxref_3_c_651_n N_RN_c_1470_n ) capacitor c=0.0236835f //x=8.88 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_689 ( N_noxref_3_c_624_n N_RN_c_1470_n ) capacitor c=0.022454f //x=10.73 \
 //y=2.08 //x2=16.165 //y2=2.22
cc_690 ( N_noxref_3_c_629_n N_RN_c_1470_n ) capacitor c=0.00814985f //x=10.535 \
 //y=1.915 //x2=16.165 //y2=2.22
cc_691 ( N_noxref_3_c_616_n N_RN_c_1478_n ) capacitor c=0.00756268f //x=8.765 \
 //y=3.33 //x2=8.255 //y2=2.22
cc_692 ( N_noxref_3_c_651_n N_RN_c_1478_n ) capacitor c=0.00184436f //x=8.88 \
 //y=3.33 //x2=8.255 //y2=2.22
cc_693 ( N_noxref_3_c_616_n N_RN_c_1485_n ) capacitor c=0.0219712f //x=8.765 \
 //y=3.33 //x2=8.14 //y2=2.08
cc_694 ( N_noxref_3_c_719_p N_RN_c_1485_n ) capacitor c=0.00131333f //x=8.995 \
 //y=3.33 //x2=8.14 //y2=2.08
cc_695 ( N_noxref_3_c_651_n N_RN_c_1485_n ) capacitor c=0.0804535f //x=8.88 \
 //y=3.33 //x2=8.14 //y2=2.08
cc_696 ( N_noxref_3_c_624_n N_RN_c_1485_n ) capacitor c=7.44267e-19 //x=10.73 \
 //y=2.08 //x2=8.14 //y2=2.08
cc_697 ( N_noxref_3_c_767_p N_RN_c_1485_n ) capacitor c=0.0166016f //x=8.1 \
 //y=5.155 //x2=8.14 //y2=2.08
cc_698 ( N_noxref_3_c_643_n N_RN_M26_noxref_g ) capacitor c=0.01736f //x=8.015 \
 //y=5.155 //x2=7.88 //y2=6.02
cc_699 ( N_noxref_3_M26_noxref_d N_RN_M26_noxref_g ) capacitor c=0.0180032f \
 //x=7.955 //y=5.02 //x2=7.88 //y2=6.02
cc_700 ( N_noxref_3_c_647_n N_RN_M27_noxref_g ) capacitor c=0.0194981f \
 //x=8.795 //y=5.155 //x2=8.32 //y2=6.02
cc_701 ( N_noxref_3_M26_noxref_d N_RN_M27_noxref_g ) capacitor c=0.0194246f \
 //x=7.955 //y=5.02 //x2=8.32 //y2=6.02
cc_702 ( N_noxref_3_M5_noxref_d N_RN_c_1522_n ) capacitor c=0.00217566f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=0.915
cc_703 ( N_noxref_3_M5_noxref_d N_RN_c_1523_n ) capacitor c=0.0034598f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=1.26
cc_704 ( N_noxref_3_M5_noxref_d N_RN_c_1524_n ) capacitor c=0.00546784f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=1.57
cc_705 ( N_noxref_3_M5_noxref_d N_RN_c_1525_n ) capacitor c=0.00241102f \
 //x=8.205 //y=0.915 //x2=8.505 //y2=0.76
cc_706 ( N_noxref_3_c_623_n N_RN_c_1526_n ) capacitor c=0.00371277f //x=8.795 \
 //y=1.665 //x2=8.505 //y2=1.415
cc_707 ( N_noxref_3_M5_noxref_d N_RN_c_1526_n ) capacitor c=0.0138621f \
 //x=8.205 //y=0.915 //x2=8.505 //y2=1.415
cc_708 ( N_noxref_3_M5_noxref_d N_RN_c_1528_n ) capacitor c=0.00219619f \
 //x=8.205 //y=0.915 //x2=8.66 //y2=0.915
cc_709 ( N_noxref_3_c_623_n N_RN_c_1529_n ) capacitor c=0.00457401f //x=8.795 \
 //y=1.665 //x2=8.66 //y2=1.26
cc_710 ( N_noxref_3_M5_noxref_d N_RN_c_1529_n ) capacitor c=0.00603828f \
 //x=8.205 //y=0.915 //x2=8.66 //y2=1.26
cc_711 ( N_noxref_3_c_651_n N_RN_c_1531_n ) capacitor c=0.00709342f //x=8.88 \
 //y=3.33 //x2=8.14 //y2=2.08
cc_712 ( N_noxref_3_c_651_n N_RN_c_1532_n ) capacitor c=0.00283672f //x=8.88 \
 //y=3.33 //x2=8.14 //y2=1.915
cc_713 ( N_noxref_3_M5_noxref_d N_RN_c_1532_n ) capacitor c=0.00661782f \
 //x=8.205 //y=0.915 //x2=8.14 //y2=1.915
cc_714 ( N_noxref_3_c_647_n N_RN_c_1534_n ) capacitor c=0.00201851f //x=8.795 \
 //y=5.155 //x2=8.14 //y2=4.7
cc_715 ( N_noxref_3_c_651_n N_RN_c_1534_n ) capacitor c=0.013844f //x=8.88 \
 //y=3.33 //x2=8.14 //y2=4.7
cc_716 ( N_noxref_3_c_767_p N_RN_c_1534_n ) capacitor c=0.00475601f //x=8.1 \
 //y=5.155 //x2=8.14 //y2=4.7
cc_717 ( N_noxref_3_c_616_n N_noxref_9_c_1895_n ) capacitor c=0.0558554f \
 //x=8.765 //y=3.33 //x2=11.355 //y2=4.07
cc_718 ( N_noxref_3_c_620_n N_noxref_9_c_1895_n ) capacitor c=0.0135672f \
 //x=3.445 //y=3.33 //x2=11.355 //y2=4.07
cc_719 ( N_noxref_3_c_621_n N_noxref_9_c_1895_n ) capacitor c=0.010979f \
 //x=10.615 //y=3.33 //x2=11.355 //y2=4.07
cc_720 ( N_noxref_3_c_719_p N_noxref_9_c_1895_n ) capacitor c=4.80262e-19 \
 //x=8.995 //y=3.33 //x2=11.355 //y2=4.07
cc_721 ( N_noxref_3_c_622_n N_noxref_9_c_1895_n ) capacitor c=0.0206302f \
 //x=3.33 //y=2.08 //x2=11.355 //y2=4.07
cc_722 ( N_noxref_3_c_651_n N_noxref_9_c_1895_n ) capacitor c=0.0181982f \
 //x=8.88 //y=3.33 //x2=11.355 //y2=4.07
cc_723 ( N_noxref_3_c_624_n N_noxref_9_c_1895_n ) capacitor c=0.0184765f \
 //x=10.73 //y=2.08 //x2=11.355 //y2=4.07
cc_724 ( N_noxref_3_c_624_n N_noxref_9_c_1998_n ) capacitor c=0.00179385f \
 //x=10.73 //y=2.08 //x2=11.585 //y2=4.07
cc_725 ( N_noxref_3_c_622_n N_noxref_9_c_1898_n ) capacitor c=0.00175117f \
 //x=3.33 //y=2.08 //x2=1.11 //y2=2.08
cc_726 ( N_noxref_3_c_624_n N_noxref_9_c_2000_n ) capacitor c=0.00400249f \
 //x=10.73 //y=2.08 //x2=11.47 //y2=4.535
cc_727 ( N_noxref_3_c_663_n N_noxref_9_c_2000_n ) capacitor c=0.00417994f \
 //x=10.73 //y=4.7 //x2=11.47 //y2=4.535
cc_728 ( N_noxref_3_c_621_n N_noxref_9_c_1899_n ) capacitor c=0.00318578f \
 //x=10.615 //y=3.33 //x2=11.47 //y2=2.08
cc_729 ( N_noxref_3_c_651_n N_noxref_9_c_1899_n ) capacitor c=9.69022e-19 \
 //x=8.88 //y=3.33 //x2=11.47 //y2=2.08
cc_730 ( N_noxref_3_c_624_n N_noxref_9_c_1899_n ) capacitor c=0.0771626f \
 //x=10.73 //y=2.08 //x2=11.47 //y2=2.08
cc_731 ( N_noxref_3_c_629_n N_noxref_9_c_1899_n ) capacitor c=0.00284029f \
 //x=10.535 //y=1.915 //x2=11.47 //y2=2.08
cc_732 ( N_noxref_3_M28_noxref_g N_noxref_9_M30_noxref_g ) capacitor \
 c=0.0104611f //x=10.63 //y=6.02 //x2=11.51 //y2=6.02
cc_733 ( N_noxref_3_M29_noxref_g N_noxref_9_M30_noxref_g ) capacitor \
 c=0.106811f //x=11.07 //y=6.02 //x2=11.51 //y2=6.02
cc_734 ( N_noxref_3_M29_noxref_g N_noxref_9_M31_noxref_g ) capacitor \
 c=0.0100341f //x=11.07 //y=6.02 //x2=11.95 //y2=6.02
cc_735 ( N_noxref_3_c_625_n N_noxref_9_c_2009_n ) capacitor c=4.86506e-19 \
 //x=10.535 //y=0.865 //x2=11.505 //y2=0.905
cc_736 ( N_noxref_3_c_627_n N_noxref_9_c_2009_n ) capacitor c=0.00152104f \
 //x=10.535 //y=1.21 //x2=11.505 //y2=0.905
cc_737 ( N_noxref_3_c_632_n N_noxref_9_c_2009_n ) capacitor c=0.0151475f \
 //x=11.065 //y=0.865 //x2=11.505 //y2=0.905
cc_738 ( N_noxref_3_c_628_n N_noxref_9_c_2012_n ) capacitor c=0.00109982f \
 //x=10.535 //y=1.52 //x2=11.505 //y2=1.25
cc_739 ( N_noxref_3_c_634_n N_noxref_9_c_2012_n ) capacitor c=0.0111064f \
 //x=11.065 //y=1.21 //x2=11.505 //y2=1.25
cc_740 ( N_noxref_3_c_628_n N_noxref_9_c_2014_n ) capacitor c=9.57794e-19 \
 //x=10.535 //y=1.52 //x2=11.505 //y2=1.56
cc_741 ( N_noxref_3_c_629_n N_noxref_9_c_2014_n ) capacitor c=0.00662747f \
 //x=10.535 //y=1.915 //x2=11.505 //y2=1.56
cc_742 ( N_noxref_3_c_634_n N_noxref_9_c_2014_n ) capacitor c=0.00862358f \
 //x=11.065 //y=1.21 //x2=11.505 //y2=1.56
cc_743 ( N_noxref_3_c_632_n N_noxref_9_c_2017_n ) capacitor c=0.00124821f \
 //x=11.065 //y=0.865 //x2=12.035 //y2=0.905
cc_744 ( N_noxref_3_c_634_n N_noxref_9_c_2018_n ) capacitor c=0.00200715f \
 //x=11.065 //y=1.21 //x2=12.035 //y2=1.25
cc_745 ( N_noxref_3_c_624_n N_noxref_9_c_2019_n ) capacitor c=0.00282278f \
 //x=10.73 //y=2.08 //x2=11.47 //y2=2.08
cc_746 ( N_noxref_3_c_629_n N_noxref_9_c_2019_n ) capacitor c=0.0172771f \
 //x=10.535 //y=1.915 //x2=11.47 //y2=2.08
cc_747 ( N_noxref_3_c_624_n N_noxref_9_c_2021_n ) capacitor c=0.00344981f \
 //x=10.73 //y=2.08 //x2=11.5 //y2=4.7
cc_748 ( N_noxref_3_c_663_n N_noxref_9_c_2021_n ) capacitor c=0.0293367f \
 //x=10.73 //y=4.7 //x2=11.5 //y2=4.7
cc_749 ( N_noxref_3_c_616_n N_noxref_12_c_2475_n ) capacitor c=2.45218e-19 \
 //x=8.765 //y=3.33 //x2=3.985 //y2=0.54
cc_750 ( N_noxref_3_c_622_n N_noxref_12_c_2475_n ) capacitor c=0.00208521f \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_751 ( N_noxref_3_c_705_p N_noxref_12_c_2475_n ) capacitor c=0.0194423f \
 //x=3.32 //y=0.915 //x2=3.985 //y2=0.54
cc_752 ( N_noxref_3_c_749_p N_noxref_12_c_2475_n ) capacitor c=0.00656458f \
 //x=3.85 //y=0.915 //x2=3.985 //y2=0.54
cc_753 ( N_noxref_3_c_700_p N_noxref_12_c_2475_n ) capacitor c=2.20712e-19 \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_754 ( N_noxref_3_c_706_p N_noxref_12_c_2489_n ) capacitor c=0.00538829f \
 //x=3.32 //y=1.26 //x2=3.1 //y2=0.995
cc_755 ( N_noxref_3_c_705_p N_noxref_12_M2_noxref_s ) capacitor c=0.00538829f \
 //x=3.32 //y=0.915 //x2=2.965 //y2=0.375
cc_756 ( N_noxref_3_c_707_p N_noxref_12_M2_noxref_s ) capacitor c=0.00538829f \
 //x=3.32 //y=1.57 //x2=2.965 //y2=0.375
cc_757 ( N_noxref_3_c_749_p N_noxref_12_M2_noxref_s ) capacitor c=0.0143002f \
 //x=3.85 //y=0.915 //x2=2.965 //y2=0.375
cc_758 ( N_noxref_3_c_728_p N_noxref_12_M2_noxref_s ) capacitor c=0.00290153f \
 //x=3.85 //y=1.26 //x2=2.965 //y2=0.375
cc_759 ( N_noxref_3_c_616_n N_D_c_2523_n ) capacitor c=0.0242474f //x=8.765 \
 //y=3.33 //x2=7.03 //y2=2.08
cc_760 ( N_noxref_3_c_637_n N_D_c_2523_n ) capacitor c=0.0144268f //x=7.135 \
 //y=5.155 //x2=7.03 //y2=2.08
cc_761 ( N_noxref_3_c_651_n N_D_c_2523_n ) capacitor c=0.00254853f //x=8.88 \
 //y=3.33 //x2=7.03 //y2=2.08
cc_762 ( N_noxref_3_c_637_n N_D_M24_noxref_g ) capacitor c=0.0165266f \
 //x=7.135 //y=5.155 //x2=7 //y2=6.02
cc_763 ( N_noxref_3_M24_noxref_d N_D_M24_noxref_g ) capacitor c=0.0180032f \
 //x=7.075 //y=5.02 //x2=7 //y2=6.02
cc_764 ( N_noxref_3_c_643_n N_D_M25_noxref_g ) capacitor c=0.01736f //x=8.015 \
 //y=5.155 //x2=7.44 //y2=6.02
cc_765 ( N_noxref_3_M24_noxref_d N_D_M25_noxref_g ) capacitor c=0.0180032f \
 //x=7.075 //y=5.02 //x2=7.44 //y2=6.02
cc_766 ( N_noxref_3_c_836_p N_D_c_2537_n ) capacitor c=0.00426767f //x=7.22 \
 //y=5.155 //x2=7.365 //y2=4.79
cc_767 ( N_noxref_3_c_637_n N_D_c_2538_n ) capacitor c=0.00322054f //x=7.135 \
 //y=5.155 //x2=7.03 //y2=4.7
cc_768 ( N_noxref_3_c_616_n N_noxref_14_c_2619_n ) capacitor c=0.00243521f \
 //x=8.765 //y=3.33 //x2=5.4 //y2=1.505
cc_769 ( N_noxref_3_c_616_n N_noxref_14_c_2603_n ) capacitor c=0.0103731f \
 //x=8.765 //y=3.33 //x2=6.285 //y2=1.59
cc_770 ( N_noxref_3_c_616_n N_noxref_14_c_2621_n ) capacitor c=0.00864153f \
 //x=8.765 //y=3.33 //x2=7.255 //y2=1.59
cc_771 ( N_noxref_3_c_616_n N_noxref_14_M3_noxref_s ) capacitor c=0.00470578f \
 //x=8.765 //y=3.33 //x2=5.265 //y2=0.375
cc_772 ( N_noxref_3_M5_noxref_d N_noxref_14_M3_noxref_s ) capacitor \
 c=0.00309936f //x=8.205 //y=0.915 //x2=5.265 //y2=0.375
cc_773 ( N_noxref_3_c_616_n N_noxref_15_c_2653_n ) capacitor c=0.00306157f \
 //x=8.765 //y=3.33 //x2=7.825 //y2=0.995
cc_774 ( N_noxref_3_c_623_n N_noxref_15_c_2658_n ) capacitor c=0.00457167f \
 //x=8.795 //y=1.665 //x2=8.795 //y2=0.54
cc_775 ( N_noxref_3_M5_noxref_d N_noxref_15_c_2658_n ) capacitor c=0.0115903f \
 //x=8.205 //y=0.915 //x2=8.795 //y2=0.54
cc_776 ( N_noxref_3_c_757_p N_noxref_15_c_2670_n ) capacitor c=0.020048f \
 //x=8.48 //y=1.665 //x2=7.91 //y2=0.995
cc_777 ( N_noxref_3_M5_noxref_d N_noxref_15_M4_noxref_d ) capacitor \
 c=5.27807e-19 //x=8.205 //y=0.915 //x2=6.67 //y2=0.91
cc_778 ( N_noxref_3_c_616_n N_noxref_15_M5_noxref_s ) capacitor c=0.00243521f \
 //x=8.765 //y=3.33 //x2=7.775 //y2=0.375
cc_779 ( N_noxref_3_c_623_n N_noxref_15_M5_noxref_s ) capacitor c=0.0196084f \
 //x=8.795 //y=1.665 //x2=7.775 //y2=0.375
cc_780 ( N_noxref_3_M5_noxref_d N_noxref_15_M5_noxref_s ) capacitor \
 c=0.0426444f //x=8.205 //y=0.915 //x2=7.775 //y2=0.375
cc_781 ( N_noxref_3_c_623_n N_noxref_16_c_2726_n ) capacitor c=3.04182e-19 \
 //x=8.795 //y=1.665 //x2=10.315 //y2=1.495
cc_782 ( N_noxref_3_c_629_n N_noxref_16_c_2726_n ) capacitor c=0.0034165f \
 //x=10.535 //y=1.915 //x2=10.315 //y2=1.495
cc_783 ( N_noxref_3_c_624_n N_noxref_16_c_2707_n ) capacitor c=0.011618f \
 //x=10.73 //y=2.08 //x2=11.2 //y2=1.58
cc_784 ( N_noxref_3_c_628_n N_noxref_16_c_2707_n ) capacitor c=0.00696403f \
 //x=10.535 //y=1.52 //x2=11.2 //y2=1.58
cc_785 ( N_noxref_3_c_629_n N_noxref_16_c_2707_n ) capacitor c=0.0174694f \
 //x=10.535 //y=1.915 //x2=11.2 //y2=1.58
cc_786 ( N_noxref_3_c_631_n N_noxref_16_c_2707_n ) capacitor c=0.00776811f \
 //x=10.91 //y=1.365 //x2=11.2 //y2=1.58
cc_787 ( N_noxref_3_c_634_n N_noxref_16_c_2707_n ) capacitor c=0.00339872f \
 //x=11.065 //y=1.21 //x2=11.2 //y2=1.58
cc_788 ( N_noxref_3_c_629_n N_noxref_16_c_2714_n ) capacitor c=6.71402e-19 \
 //x=10.535 //y=1.915 //x2=11.285 //y2=1.495
cc_789 ( N_noxref_3_c_625_n N_noxref_16_M6_noxref_s ) capacitor c=0.0327502f \
 //x=10.535 //y=0.865 //x2=10.18 //y2=0.365
cc_790 ( N_noxref_3_c_628_n N_noxref_16_M6_noxref_s ) capacitor c=3.48408e-19 \
 //x=10.535 //y=1.52 //x2=10.18 //y2=0.365
cc_791 ( N_noxref_3_c_632_n N_noxref_16_M6_noxref_s ) capacitor c=0.0120759f \
 //x=11.065 //y=0.865 //x2=10.18 //y2=0.365
cc_792 ( N_noxref_4_c_879_n N_CLK_c_1011_n ) capacitor c=0.0185297f //x=11.645 \
 //y=5.2 //x2=15.055 //y2=4.44
cc_793 ( N_noxref_4_c_883_n N_CLK_c_1011_n ) capacitor c=0.018142f //x=10.935 \
 //y=5.2 //x2=15.055 //y2=4.44
cc_794 ( N_noxref_4_c_864_n N_CLK_c_1011_n ) capacitor c=0.0208321f //x=12.21 \
 //y=3.33 //x2=15.055 //y2=4.44
cc_795 ( N_noxref_4_c_865_n N_CLK_c_1011_n ) capacitor c=0.0224037f //x=14.06 \
 //y=2.08 //x2=15.055 //y2=4.44
cc_796 ( N_noxref_4_c_897_n N_CLK_c_1011_n ) capacitor c=0.0168539f //x=14.335 \
 //y=4.79 //x2=15.055 //y2=4.44
cc_797 ( N_noxref_4_c_862_n N_CLK_c_1010_n ) capacitor c=0.00520283f \
 //x=13.945 //y=3.33 //x2=15.17 //y2=2.08
cc_798 ( N_noxref_4_c_864_n N_CLK_c_1010_n ) capacitor c=5.77178e-19 //x=12.21 \
 //y=3.33 //x2=15.17 //y2=2.08
cc_799 ( N_noxref_4_c_865_n N_CLK_c_1010_n ) capacitor c=0.0469865f //x=14.06 \
 //y=2.08 //x2=15.17 //y2=2.08
cc_800 ( N_noxref_4_c_870_n N_CLK_c_1010_n ) capacitor c=0.00210802f //x=13.76 \
 //y=1.915 //x2=15.17 //y2=2.08
cc_801 ( N_noxref_4_c_927_p N_CLK_c_1010_n ) capacitor c=0.00147352f \
 //x=14.625 //y=4.79 //x2=15.17 //y2=2.08
cc_802 ( N_noxref_4_c_897_n N_CLK_c_1010_n ) capacitor c=0.00141297f \
 //x=14.335 //y=4.79 //x2=15.17 //y2=2.08
cc_803 ( N_noxref_4_M32_noxref_g N_CLK_M34_noxref_g ) capacitor c=0.0105869f \
 //x=14.26 //y=6.02 //x2=15.14 //y2=6.02
cc_804 ( N_noxref_4_M33_noxref_g N_CLK_M34_noxref_g ) capacitor c=0.10632f \
 //x=14.7 //y=6.02 //x2=15.14 //y2=6.02
cc_805 ( N_noxref_4_M33_noxref_g N_CLK_M35_noxref_g ) capacitor c=0.0101598f \
 //x=14.7 //y=6.02 //x2=15.58 //y2=6.02
cc_806 ( N_noxref_4_c_866_n N_CLK_c_1082_n ) capacitor c=5.72482e-19 //x=13.76 \
 //y=0.875 //x2=14.735 //y2=0.91
cc_807 ( N_noxref_4_c_868_n N_CLK_c_1082_n ) capacitor c=0.00149976f //x=13.76 \
 //y=1.22 //x2=14.735 //y2=0.91
cc_808 ( N_noxref_4_c_873_n N_CLK_c_1082_n ) capacitor c=0.0160123f //x=14.29 \
 //y=0.875 //x2=14.735 //y2=0.91
cc_809 ( N_noxref_4_c_869_n N_CLK_c_1085_n ) capacitor c=0.00111227f //x=13.76 \
 //y=1.53 //x2=14.735 //y2=1.22
cc_810 ( N_noxref_4_c_875_n N_CLK_c_1085_n ) capacitor c=0.0124075f //x=14.29 \
 //y=1.22 //x2=14.735 //y2=1.22
cc_811 ( N_noxref_4_c_873_n N_CLK_c_1087_n ) capacitor c=0.00103227f //x=14.29 \
 //y=0.875 //x2=15.26 //y2=0.91
cc_812 ( N_noxref_4_c_875_n N_CLK_c_1088_n ) capacitor c=0.0010154f //x=14.29 \
 //y=1.22 //x2=15.26 //y2=1.22
cc_813 ( N_noxref_4_c_875_n N_CLK_c_1089_n ) capacitor c=9.23422e-19 //x=14.29 \
 //y=1.22 //x2=15.26 //y2=1.45
cc_814 ( N_noxref_4_c_865_n N_CLK_c_1090_n ) capacitor c=0.00203769f //x=14.06 \
 //y=2.08 //x2=15.26 //y2=1.915
cc_815 ( N_noxref_4_c_870_n N_CLK_c_1090_n ) capacitor c=0.00834532f //x=13.76 \
 //y=1.915 //x2=15.26 //y2=1.915
cc_816 ( N_noxref_4_c_865_n N_CLK_c_1092_n ) capacitor c=0.00183762f //x=14.06 \
 //y=2.08 //x2=15.17 //y2=4.7
cc_817 ( N_noxref_4_c_927_p N_CLK_c_1092_n ) capacitor c=0.0168581f //x=14.625 \
 //y=4.79 //x2=15.17 //y2=4.7
cc_818 ( N_noxref_4_c_897_n N_CLK_c_1092_n ) capacitor c=0.00484466f \
 //x=14.335 //y=4.79 //x2=15.17 //y2=4.7
cc_819 ( N_noxref_4_c_862_n N_noxref_6_c_1224_n ) capacitor c=0.176049f \
 //x=13.945 //y=3.33 //x2=18.755 //y2=3.7
cc_820 ( N_noxref_4_c_910_n N_noxref_6_c_1224_n ) capacitor c=0.0293967f \
 //x=12.325 //y=3.33 //x2=18.755 //y2=3.7
cc_821 ( N_noxref_4_c_864_n N_noxref_6_c_1224_n ) capacitor c=0.0206034f \
 //x=12.21 //y=3.33 //x2=18.755 //y2=3.7
cc_822 ( N_noxref_4_c_865_n N_noxref_6_c_1224_n ) capacitor c=0.0216236f \
 //x=14.06 //y=2.08 //x2=18.755 //y2=3.7
cc_823 ( N_noxref_4_c_862_n N_RN_c_1470_n ) capacitor c=0.0546488f //x=13.945 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_824 ( N_noxref_4_c_910_n N_RN_c_1470_n ) capacitor c=0.00761783f //x=12.325 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_825 ( N_noxref_4_c_951_p N_RN_c_1470_n ) capacitor c=0.0146822f //x=11.855 \
 //y=1.655 //x2=16.165 //y2=2.22
cc_826 ( N_noxref_4_c_864_n N_RN_c_1470_n ) capacitor c=0.0238578f //x=12.21 \
 //y=3.33 //x2=16.165 //y2=2.22
cc_827 ( N_noxref_4_c_865_n N_RN_c_1470_n ) capacitor c=0.0232222f //x=14.06 \
 //y=2.08 //x2=16.165 //y2=2.22
cc_828 ( N_noxref_4_c_870_n N_RN_c_1470_n ) capacitor c=0.0104117f //x=13.76 \
 //y=1.915 //x2=16.165 //y2=2.22
cc_829 ( N_noxref_4_c_865_n N_RN_c_1486_n ) capacitor c=0.0014519f //x=14.06 \
 //y=2.08 //x2=16.28 //y2=2.08
cc_830 ( N_noxref_4_c_862_n N_noxref_9_c_1922_n ) capacitor c=0.0107156f \
 //x=13.945 //y=3.33 //x2=16.905 //y2=4.07
cc_831 ( N_noxref_4_c_910_n N_noxref_9_c_1922_n ) capacitor c=8.88358e-19 \
 //x=12.325 //y=3.33 //x2=16.905 //y2=4.07
cc_832 ( N_noxref_4_c_864_n N_noxref_9_c_1922_n ) capacitor c=0.0181936f \
 //x=12.21 //y=3.33 //x2=16.905 //y2=4.07
cc_833 ( N_noxref_4_c_865_n N_noxref_9_c_1922_n ) capacitor c=0.019517f \
 //x=14.06 //y=2.08 //x2=16.905 //y2=4.07
cc_834 ( N_noxref_4_c_864_n N_noxref_9_c_1998_n ) capacitor c=0.00179385f \
 //x=12.21 //y=3.33 //x2=11.585 //y2=4.07
cc_835 ( N_noxref_4_c_879_n N_noxref_9_c_2000_n ) capacitor c=0.0127164f \
 //x=11.645 //y=5.2 //x2=11.47 //y2=4.535
cc_836 ( N_noxref_4_c_864_n N_noxref_9_c_2000_n ) capacitor c=0.0101115f \
 //x=12.21 //y=3.33 //x2=11.47 //y2=4.535
cc_837 ( N_noxref_4_c_910_n N_noxref_9_c_1899_n ) capacitor c=0.00329059f \
 //x=12.325 //y=3.33 //x2=11.47 //y2=2.08
cc_838 ( N_noxref_4_c_864_n N_noxref_9_c_1899_n ) capacitor c=0.0721848f \
 //x=12.21 //y=3.33 //x2=11.47 //y2=2.08
cc_839 ( N_noxref_4_c_865_n N_noxref_9_c_1899_n ) capacitor c=9.69022e-19 \
 //x=14.06 //y=2.08 //x2=11.47 //y2=2.08
cc_840 ( N_noxref_4_M33_noxref_g N_noxref_9_c_1943_n ) capacitor c=0.0168349f \
 //x=14.7 //y=6.02 //x2=15.275 //y2=5.155
cc_841 ( N_noxref_4_c_864_n N_noxref_9_c_1947_n ) capacitor c=2.97874e-19 \
 //x=12.21 //y=3.33 //x2=14.565 //y2=5.155
cc_842 ( N_noxref_4_M32_noxref_g N_noxref_9_c_1947_n ) capacitor c=0.0213876f \
 //x=14.26 //y=6.02 //x2=14.565 //y2=5.155
cc_843 ( N_noxref_4_c_927_p N_noxref_9_c_1947_n ) capacitor c=0.00428486f \
 //x=14.625 //y=4.79 //x2=14.565 //y2=5.155
cc_844 ( N_noxref_4_c_879_n N_noxref_9_M30_noxref_g ) capacitor c=0.0166421f \
 //x=11.645 //y=5.2 //x2=11.51 //y2=6.02
cc_845 ( N_noxref_4_M30_noxref_d N_noxref_9_M30_noxref_g ) capacitor \
 c=0.0173476f //x=11.585 //y=5.02 //x2=11.51 //y2=6.02
cc_846 ( N_noxref_4_c_885_n N_noxref_9_M31_noxref_g ) capacitor c=0.018922f \
 //x=12.125 //y=5.2 //x2=11.95 //y2=6.02
cc_847 ( N_noxref_4_M30_noxref_d N_noxref_9_M31_noxref_g ) capacitor \
 c=0.0179769f //x=11.585 //y=5.02 //x2=11.95 //y2=6.02
cc_848 ( N_noxref_4_M7_noxref_d N_noxref_9_c_2009_n ) capacitor c=0.00217566f \
 //x=11.58 //y=0.905 //x2=11.505 //y2=0.905
cc_849 ( N_noxref_4_M7_noxref_d N_noxref_9_c_2012_n ) capacitor c=0.0034598f \
 //x=11.58 //y=0.905 //x2=11.505 //y2=1.25
cc_850 ( N_noxref_4_M7_noxref_d N_noxref_9_c_2014_n ) capacitor c=0.00669531f \
 //x=11.58 //y=0.905 //x2=11.505 //y2=1.56
cc_851 ( N_noxref_4_c_864_n N_noxref_9_c_2044_n ) capacitor c=0.0142673f \
 //x=12.21 //y=3.33 //x2=11.875 //y2=4.79
cc_852 ( N_noxref_4_c_978_p N_noxref_9_c_2044_n ) capacitor c=0.00407665f \
 //x=11.73 //y=5.2 //x2=11.875 //y2=4.79
cc_853 ( N_noxref_4_M7_noxref_d N_noxref_9_c_2046_n ) capacitor c=0.00241102f \
 //x=11.58 //y=0.905 //x2=11.88 //y2=0.75
cc_854 ( N_noxref_4_c_863_n N_noxref_9_c_2047_n ) capacitor c=0.00371277f \
 //x=12.125 //y=1.655 //x2=11.88 //y2=1.405
cc_855 ( N_noxref_4_M7_noxref_d N_noxref_9_c_2047_n ) capacitor c=0.0137169f \
 //x=11.58 //y=0.905 //x2=11.88 //y2=1.405
cc_856 ( N_noxref_4_M7_noxref_d N_noxref_9_c_2017_n ) capacitor c=0.00132245f \
 //x=11.58 //y=0.905 //x2=12.035 //y2=0.905
cc_857 ( N_noxref_4_c_863_n N_noxref_9_c_2018_n ) capacitor c=0.00457401f \
 //x=12.125 //y=1.655 //x2=12.035 //y2=1.25
cc_858 ( N_noxref_4_M7_noxref_d N_noxref_9_c_2018_n ) capacitor c=0.00566463f \
 //x=11.58 //y=0.905 //x2=12.035 //y2=1.25
cc_859 ( N_noxref_4_c_864_n N_noxref_9_c_2019_n ) capacitor c=0.00731987f \
 //x=12.21 //y=3.33 //x2=11.47 //y2=2.08
cc_860 ( N_noxref_4_c_864_n N_noxref_9_c_2053_n ) capacitor c=0.00306024f \
 //x=12.21 //y=3.33 //x2=11.47 //y2=1.915
cc_861 ( N_noxref_4_M7_noxref_d N_noxref_9_c_2053_n ) capacitor c=0.00660593f \
 //x=11.58 //y=0.905 //x2=11.47 //y2=1.915
cc_862 ( N_noxref_4_c_879_n N_noxref_9_c_2021_n ) capacitor c=0.00346527f \
 //x=11.645 //y=5.2 //x2=11.5 //y2=4.7
cc_863 ( N_noxref_4_c_864_n N_noxref_9_c_2021_n ) capacitor c=0.00517969f \
 //x=12.21 //y=3.33 //x2=11.5 //y2=4.7
cc_864 ( N_noxref_4_M33_noxref_g N_noxref_9_M32_noxref_d ) capacitor \
 c=0.0180032f //x=14.7 //y=6.02 //x2=14.335 //y2=5.02
cc_865 ( N_noxref_4_c_951_p N_noxref_16_c_2726_n ) capacitor c=3.15806e-19 \
 //x=11.855 //y=1.655 //x2=10.315 //y2=1.495
cc_866 ( N_noxref_4_c_951_p N_noxref_16_c_2714_n ) capacitor c=0.020324f \
 //x=11.855 //y=1.655 //x2=11.285 //y2=1.495
cc_867 ( N_noxref_4_c_863_n N_noxref_16_c_2715_n ) capacitor c=0.00457164f \
 //x=12.125 //y=1.655 //x2=12.17 //y2=0.53
cc_868 ( N_noxref_4_M7_noxref_d N_noxref_16_c_2715_n ) capacitor c=0.0115831f \
 //x=11.58 //y=0.905 //x2=12.17 //y2=0.53
cc_869 ( N_noxref_4_c_863_n N_noxref_16_M6_noxref_s ) capacitor c=0.013435f \
 //x=12.125 //y=1.655 //x2=10.18 //y2=0.365
cc_870 ( N_noxref_4_M7_noxref_d N_noxref_16_M6_noxref_s ) capacitor \
 c=0.0439476f //x=11.58 //y=0.905 //x2=10.18 //y2=0.365
cc_871 ( N_noxref_4_c_863_n N_noxref_17_c_2775_n ) capacitor c=4.08644e-19 \
 //x=12.125 //y=1.655 //x2=13.54 //y2=1.505
cc_872 ( N_noxref_4_c_870_n N_noxref_17_c_2775_n ) capacitor c=0.0034165f \
 //x=13.76 //y=1.915 //x2=13.54 //y2=1.505
cc_873 ( N_noxref_4_c_865_n N_noxref_17_c_2759_n ) capacitor c=0.0115578f \
 //x=14.06 //y=2.08 //x2=14.425 //y2=1.59
cc_874 ( N_noxref_4_c_869_n N_noxref_17_c_2759_n ) capacitor c=0.00697148f \
 //x=13.76 //y=1.53 //x2=14.425 //y2=1.59
cc_875 ( N_noxref_4_c_870_n N_noxref_17_c_2759_n ) capacitor c=0.0204849f \
 //x=13.76 //y=1.915 //x2=14.425 //y2=1.59
cc_876 ( N_noxref_4_c_872_n N_noxref_17_c_2759_n ) capacitor c=0.00610316f \
 //x=14.135 //y=1.375 //x2=14.425 //y2=1.59
cc_877 ( N_noxref_4_c_875_n N_noxref_17_c_2759_n ) capacitor c=0.00698822f \
 //x=14.29 //y=1.22 //x2=14.425 //y2=1.59
cc_878 ( N_noxref_4_c_866_n N_noxref_17_M8_noxref_s ) capacitor c=0.0327271f \
 //x=13.76 //y=0.875 //x2=13.405 //y2=0.375
cc_879 ( N_noxref_4_c_869_n N_noxref_17_M8_noxref_s ) capacitor c=7.99997e-19 \
 //x=13.76 //y=1.53 //x2=13.405 //y2=0.375
cc_880 ( N_noxref_4_c_870_n N_noxref_17_M8_noxref_s ) capacitor c=0.00122123f \
 //x=13.76 //y=1.915 //x2=13.405 //y2=0.375
cc_881 ( N_noxref_4_c_873_n N_noxref_17_M8_noxref_s ) capacitor c=0.0121427f \
 //x=14.29 //y=0.875 //x2=13.405 //y2=0.375
cc_882 ( N_noxref_4_M7_noxref_d N_noxref_17_M8_noxref_s ) capacitor \
 c=2.53688e-19 //x=11.58 //y=0.905 //x2=13.405 //y2=0.375
cc_883 ( N_CLK_c_1011_n N_noxref_6_c_1297_n ) capacitor c=0.00910993f \
 //x=15.055 //y=4.44 //x2=5.805 //y2=3.7
cc_884 ( N_CLK_c_1011_n N_noxref_6_c_1298_n ) capacitor c=7.95009e-19 \
 //x=15.055 //y=4.44 //x2=4.185 //y2=3.7
cc_885 ( N_CLK_c_1011_n N_noxref_6_c_1224_n ) capacitor c=0.06678f //x=15.055 \
 //y=4.44 //x2=18.755 //y2=3.7
cc_886 ( N_CLK_c_1010_n N_noxref_6_c_1224_n ) capacitor c=0.0238781f //x=15.17 \
 //y=2.08 //x2=18.755 //y2=3.7
cc_887 ( N_CLK_c_1011_n N_noxref_6_c_1305_n ) capacitor c=6.59178e-19 \
 //x=15.055 //y=4.44 //x2=6.035 //y2=3.7
cc_888 ( N_CLK_c_1028_n N_noxref_6_c_1249_n ) capacitor c=0.00330099f \
 //x=2.335 //y=4.44 //x2=2.325 //y2=5.155
cc_889 ( N_CLK_c_1009_n N_noxref_6_c_1249_n ) capacitor c=0.014564f //x=2.22 \
 //y=2.08 //x2=2.325 //y2=5.155
cc_890 ( N_CLK_M18_noxref_g N_noxref_6_c_1249_n ) capacitor c=0.016514f \
 //x=2.19 //y=6.02 //x2=2.325 //y2=5.155
cc_891 ( N_CLK_c_1066_n N_noxref_6_c_1249_n ) capacitor c=0.00322046f //x=2.22 \
 //y=4.7 //x2=2.325 //y2=5.155
cc_892 ( N_CLK_M19_noxref_g N_noxref_6_c_1255_n ) capacitor c=0.01736f \
 //x=2.63 //y=6.02 //x2=3.205 //y2=5.155
cc_893 ( N_CLK_c_1011_n N_noxref_6_c_1259_n ) capacitor c=0.0183122f \
 //x=15.055 //y=4.44 //x2=3.985 //y2=5.155
cc_894 ( N_CLK_c_1011_n N_noxref_6_c_1263_n ) capacitor c=0.0210274f \
 //x=15.055 //y=4.44 //x2=4.07 //y2=3.7
cc_895 ( N_CLK_c_1009_n N_noxref_6_c_1263_n ) capacitor c=0.00319363f //x=2.22 \
 //y=2.08 //x2=4.07 //y2=3.7
cc_896 ( N_CLK_c_1011_n N_noxref_6_c_1226_n ) capacitor c=0.0208709f \
 //x=15.055 //y=4.44 //x2=5.92 //y2=2.08
cc_897 ( N_CLK_c_1011_n N_noxref_6_c_1355_n ) capacitor c=0.0311227f \
 //x=15.055 //y=4.44 //x2=2.41 //y2=5.155
cc_898 ( N_CLK_c_1065_n N_noxref_6_c_1355_n ) capacitor c=0.00426767f \
 //x=2.555 //y=4.79 //x2=2.41 //y2=5.155
cc_899 ( N_CLK_c_1011_n N_noxref_6_c_1278_n ) capacitor c=0.0166984f \
 //x=15.055 //y=4.44 //x2=6.195 //y2=4.79
cc_900 ( N_CLK_M18_noxref_g N_noxref_6_M18_noxref_d ) capacitor c=0.0180032f \
 //x=2.19 //y=6.02 //x2=2.265 //y2=5.02
cc_901 ( N_CLK_M19_noxref_g N_noxref_6_M18_noxref_d ) capacitor c=0.0180032f \
 //x=2.63 //y=6.02 //x2=2.265 //y2=5.02
cc_902 ( N_CLK_c_1010_n N_RN_c_1470_n ) capacitor c=0.0242349f //x=15.17 \
 //y=2.08 //x2=16.165 //y2=2.22
cc_903 ( N_CLK_c_1090_n N_RN_c_1470_n ) capacitor c=0.00615803f //x=15.26 \
 //y=1.915 //x2=16.165 //y2=2.22
cc_904 ( N_CLK_c_1010_n N_RN_c_1484_n ) capacitor c=0.00165648f //x=15.17 \
 //y=2.08 //x2=16.395 //y2=2.22
cc_905 ( N_CLK_c_1090_n N_RN_c_1484_n ) capacitor c=2.3323e-19 //x=15.26 \
 //y=1.915 //x2=16.395 //y2=2.22
cc_906 ( N_CLK_c_1011_n N_RN_c_1485_n ) capacitor c=0.0200057f //x=15.055 \
 //y=4.44 //x2=8.14 //y2=2.08
cc_907 ( N_CLK_c_1011_n N_RN_c_1486_n ) capacitor c=0.00551083f //x=15.055 \
 //y=4.44 //x2=16.28 //y2=2.08
cc_908 ( N_CLK_c_1010_n N_RN_c_1486_n ) capacitor c=0.0492003f //x=15.17 \
 //y=2.08 //x2=16.28 //y2=2.08
cc_909 ( N_CLK_c_1090_n N_RN_c_1486_n ) capacitor c=0.00203728f //x=15.26 \
 //y=1.915 //x2=16.28 //y2=2.08
cc_910 ( N_CLK_c_1092_n N_RN_c_1486_n ) capacitor c=0.00142741f //x=15.17 \
 //y=4.7 //x2=16.28 //y2=2.08
cc_911 ( N_CLK_M34_noxref_g N_RN_M36_noxref_g ) capacitor c=0.0101598f \
 //x=15.14 //y=6.02 //x2=16.02 //y2=6.02
cc_912 ( N_CLK_M35_noxref_g N_RN_M36_noxref_g ) capacitor c=0.0602553f \
 //x=15.58 //y=6.02 //x2=16.02 //y2=6.02
cc_913 ( N_CLK_M35_noxref_g N_RN_M37_noxref_g ) capacitor c=0.0101598f \
 //x=15.58 //y=6.02 //x2=16.46 //y2=6.02
cc_914 ( N_CLK_c_1087_n N_RN_c_1556_n ) capacitor c=0.00456962f //x=15.26 \
 //y=0.91 //x2=16.27 //y2=0.915
cc_915 ( N_CLK_c_1088_n N_RN_c_1557_n ) capacitor c=0.00438372f //x=15.26 \
 //y=1.22 //x2=16.27 //y2=1.26
cc_916 ( N_CLK_c_1089_n N_RN_c_1558_n ) capacitor c=0.00438372f //x=15.26 \
 //y=1.45 //x2=16.27 //y2=1.57
cc_917 ( N_CLK_c_1011_n N_RN_c_1534_n ) capacitor c=0.0111881f //x=15.055 \
 //y=4.44 //x2=8.14 //y2=4.7
cc_918 ( N_CLK_c_1010_n N_RN_c_1560_n ) capacitor c=0.00201097f //x=15.17 \
 //y=2.08 //x2=16.28 //y2=2.08
cc_919 ( N_CLK_c_1090_n N_RN_c_1560_n ) capacitor c=0.00828003f //x=15.26 \
 //y=1.915 //x2=16.28 //y2=2.08
cc_920 ( N_CLK_c_1090_n N_RN_c_1562_n ) capacitor c=0.00438372f //x=15.26 \
 //y=1.915 //x2=16.28 //y2=1.915
cc_921 ( N_CLK_c_1010_n N_RN_c_1563_n ) capacitor c=0.00218014f //x=15.17 \
 //y=2.08 //x2=16.28 //y2=4.7
cc_922 ( N_CLK_c_1134_p N_RN_c_1563_n ) capacitor c=0.0611812f //x=15.505 \
 //y=4.79 //x2=16.28 //y2=4.7
cc_923 ( N_CLK_c_1092_n N_RN_c_1563_n ) capacitor c=0.00487508f //x=15.17 \
 //y=4.7 //x2=16.28 //y2=4.7
cc_924 ( N_CLK_c_1011_n N_noxref_9_c_1895_n ) capacitor c=0.784553f //x=15.055 \
 //y=4.44 //x2=11.355 //y2=4.07
cc_925 ( N_CLK_c_1028_n N_noxref_9_c_1895_n ) capacitor c=0.0291328f //x=2.335 \
 //y=4.44 //x2=11.355 //y2=4.07
cc_926 ( N_CLK_c_1009_n N_noxref_9_c_1895_n ) capacitor c=0.0265867f //x=2.22 \
 //y=2.08 //x2=11.355 //y2=4.07
cc_927 ( N_CLK_c_1066_n N_noxref_9_c_1895_n ) capacitor c=6.38735e-19 //x=2.22 \
 //y=4.7 //x2=11.355 //y2=4.07
cc_928 ( N_CLK_c_1009_n N_noxref_9_c_1896_n ) capacitor c=0.00128547f //x=2.22 \
 //y=2.08 //x2=1.225 //y2=4.07
cc_929 ( N_CLK_c_1011_n N_noxref_9_c_1922_n ) capacitor c=0.331988f //x=15.055 \
 //y=4.44 //x2=16.905 //y2=4.07
cc_930 ( N_CLK_c_1010_n N_noxref_9_c_1922_n ) capacitor c=0.0208526f //x=15.17 \
 //y=2.08 //x2=16.905 //y2=4.07
cc_931 ( N_CLK_c_1134_p N_noxref_9_c_1922_n ) capacitor c=0.00660387f \
 //x=15.505 //y=4.79 //x2=16.905 //y2=4.07
cc_932 ( N_CLK_c_1011_n N_noxref_9_c_1998_n ) capacitor c=0.0263375f \
 //x=15.055 //y=4.44 //x2=11.585 //y2=4.07
cc_933 ( N_CLK_c_1028_n N_noxref_9_c_1898_n ) capacitor c=0.00551083f \
 //x=2.335 //y=4.44 //x2=1.11 //y2=2.08
cc_934 ( N_CLK_c_1009_n N_noxref_9_c_1898_n ) capacitor c=0.0535714f //x=2.22 \
 //y=2.08 //x2=1.11 //y2=2.08
cc_935 ( N_CLK_c_1062_n N_noxref_9_c_1898_n ) capacitor c=0.00231304f //x=2.31 \
 //y=1.915 //x2=1.11 //y2=2.08
cc_936 ( N_CLK_c_1066_n N_noxref_9_c_1898_n ) capacitor c=0.00183762f //x=2.22 \
 //y=4.7 //x2=1.11 //y2=2.08
cc_937 ( N_CLK_c_1011_n N_noxref_9_c_2000_n ) capacitor c=0.0016972f \
 //x=15.055 //y=4.44 //x2=11.47 //y2=4.535
cc_938 ( N_CLK_c_1011_n N_noxref_9_c_1899_n ) capacitor c=0.0207534f \
 //x=15.055 //y=4.44 //x2=11.47 //y2=2.08
cc_939 ( N_CLK_c_1011_n N_noxref_9_c_1943_n ) capacitor c=0.00241768f \
 //x=15.055 //y=4.44 //x2=15.275 //y2=5.155
cc_940 ( N_CLK_c_1010_n N_noxref_9_c_1943_n ) capacitor c=0.0143918f //x=15.17 \
 //y=2.08 //x2=15.275 //y2=5.155
cc_941 ( N_CLK_M34_noxref_g N_noxref_9_c_1943_n ) capacitor c=0.016514f \
 //x=15.14 //y=6.02 //x2=15.275 //y2=5.155
cc_942 ( N_CLK_c_1092_n N_noxref_9_c_1943_n ) capacitor c=0.00322046f \
 //x=15.17 //y=4.7 //x2=15.275 //y2=5.155
cc_943 ( N_CLK_c_1011_n N_noxref_9_c_1947_n ) capacitor c=0.0219114f \
 //x=15.055 //y=4.44 //x2=14.565 //y2=5.155
cc_944 ( N_CLK_M35_noxref_g N_noxref_9_c_1949_n ) capacitor c=0.0184045f \
 //x=15.58 //y=6.02 //x2=16.155 //y2=5.155
cc_945 ( N_CLK_c_1010_n N_noxref_9_c_1957_n ) capacitor c=0.00317726f \
 //x=15.17 //y=2.08 //x2=17.02 //y2=4.07
cc_946 ( N_CLK_c_1011_n N_noxref_9_c_2080_n ) capacitor c=0.00101864f \
 //x=15.055 //y=4.44 //x2=15.36 //y2=5.155
cc_947 ( N_CLK_c_1134_p N_noxref_9_c_2080_n ) capacitor c=0.00427771f \
 //x=15.505 //y=4.79 //x2=15.36 //y2=5.155
cc_948 ( N_CLK_M18_noxref_g N_noxref_9_M16_noxref_g ) capacitor c=0.0105869f \
 //x=2.19 //y=6.02 //x2=1.31 //y2=6.02
cc_949 ( N_CLK_M18_noxref_g N_noxref_9_M17_noxref_g ) capacitor c=0.10632f \
 //x=2.19 //y=6.02 //x2=1.75 //y2=6.02
cc_950 ( N_CLK_M19_noxref_g N_noxref_9_M17_noxref_g ) capacitor c=0.0101598f \
 //x=2.63 //y=6.02 //x2=1.75 //y2=6.02
cc_951 ( N_CLK_c_1163_p N_noxref_9_c_1904_n ) capacitor c=5.72482e-19 \
 //x=1.785 //y=0.91 //x2=0.81 //y2=0.875
cc_952 ( N_CLK_c_1163_p N_noxref_9_c_1906_n ) capacitor c=0.00149976f \
 //x=1.785 //y=0.91 //x2=0.81 //y2=1.22
cc_953 ( N_CLK_c_1165_p N_noxref_9_c_1907_n ) capacitor c=0.00111227f \
 //x=1.785 //y=1.22 //x2=0.81 //y2=1.53
cc_954 ( N_CLK_c_1009_n N_noxref_9_c_1908_n ) capacitor c=0.00238338f //x=2.22 \
 //y=2.08 //x2=0.81 //y2=1.915
cc_955 ( N_CLK_c_1062_n N_noxref_9_c_1908_n ) capacitor c=0.00964411f //x=2.31 \
 //y=1.915 //x2=0.81 //y2=1.915
cc_956 ( N_CLK_c_1163_p N_noxref_9_c_1911_n ) capacitor c=0.0160123f //x=1.785 \
 //y=0.91 //x2=1.34 //y2=0.875
cc_957 ( N_CLK_c_1059_n N_noxref_9_c_1911_n ) capacitor c=0.00103227f //x=2.31 \
 //y=0.91 //x2=1.34 //y2=0.875
cc_958 ( N_CLK_c_1165_p N_noxref_9_c_1913_n ) capacitor c=0.0124075f //x=1.785 \
 //y=1.22 //x2=1.34 //y2=1.22
cc_959 ( N_CLK_c_1060_n N_noxref_9_c_1913_n ) capacitor c=0.0010154f //x=2.31 \
 //y=1.22 //x2=1.34 //y2=1.22
cc_960 ( N_CLK_c_1061_n N_noxref_9_c_1913_n ) capacitor c=9.23422e-19 //x=2.31 \
 //y=1.45 //x2=1.34 //y2=1.22
cc_961 ( N_CLK_c_1009_n N_noxref_9_c_2095_n ) capacitor c=0.00147352f //x=2.22 \
 //y=2.08 //x2=1.675 //y2=4.79
cc_962 ( N_CLK_c_1066_n N_noxref_9_c_2095_n ) capacitor c=0.0168581f //x=2.22 \
 //y=4.7 //x2=1.675 //y2=4.79
cc_963 ( N_CLK_c_1009_n N_noxref_9_c_1974_n ) capacitor c=0.00141297f //x=2.22 \
 //y=2.08 //x2=1.385 //y2=4.79
cc_964 ( N_CLK_c_1066_n N_noxref_9_c_1974_n ) capacitor c=0.00484466f //x=2.22 \
 //y=4.7 //x2=1.385 //y2=4.79
cc_965 ( N_CLK_c_1011_n N_noxref_9_c_2044_n ) capacitor c=0.00960248f \
 //x=15.055 //y=4.44 //x2=11.875 //y2=4.79
cc_966 ( N_CLK_c_1011_n N_noxref_9_c_2021_n ) capacitor c=0.00203982f \
 //x=15.055 //y=4.44 //x2=11.5 //y2=4.7
cc_967 ( N_CLK_M34_noxref_g N_noxref_9_M34_noxref_d ) capacitor c=0.0180032f \
 //x=15.14 //y=6.02 //x2=15.215 //y2=5.02
cc_968 ( N_CLK_M35_noxref_g N_noxref_9_M34_noxref_d ) capacitor c=0.0180032f \
 //x=15.58 //y=6.02 //x2=15.215 //y2=5.02
cc_969 ( N_CLK_c_1163_p N_noxref_11_c_2430_n ) capacitor c=0.0167228f \
 //x=1.785 //y=0.91 //x2=2.445 //y2=0.54
cc_970 ( N_CLK_c_1059_n N_noxref_11_c_2430_n ) capacitor c=0.00534519f \
 //x=2.31 //y=0.91 //x2=2.445 //y2=0.54
cc_971 ( N_CLK_c_1009_n N_noxref_11_c_2441_n ) capacitor c=0.012357f //x=2.22 \
 //y=2.08 //x2=2.445 //y2=1.59
cc_972 ( N_CLK_c_1165_p N_noxref_11_c_2441_n ) capacitor c=0.0153476f \
 //x=1.785 //y=1.22 //x2=2.445 //y2=1.59
cc_973 ( N_CLK_c_1062_n N_noxref_11_c_2441_n ) capacitor c=0.0230663f //x=2.31 \
 //y=1.915 //x2=2.445 //y2=1.59
cc_974 ( N_CLK_c_1163_p N_noxref_11_M0_noxref_s ) capacitor c=0.00798959f \
 //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_975 ( N_CLK_c_1061_n N_noxref_11_M0_noxref_s ) capacitor c=0.00212176f \
 //x=2.31 //y=1.45 //x2=0.455 //y2=0.375
cc_976 ( N_CLK_c_1062_n N_noxref_11_M0_noxref_s ) capacitor c=0.00298115f \
 //x=2.31 //y=1.915 //x2=0.455 //y2=0.375
cc_977 ( N_CLK_c_1189_p N_noxref_12_c_2470_n ) capacitor c=2.14837e-19 \
 //x=2.155 //y=0.755 //x2=3.015 //y2=0.995
cc_978 ( N_CLK_c_1059_n N_noxref_12_c_2470_n ) capacitor c=0.00123426f \
 //x=2.31 //y=0.91 //x2=3.015 //y2=0.995
cc_979 ( N_CLK_c_1060_n N_noxref_12_c_2470_n ) capacitor c=0.0129288f //x=2.31 \
 //y=1.22 //x2=3.015 //y2=0.995
cc_980 ( N_CLK_c_1061_n N_noxref_12_c_2470_n ) capacitor c=0.00142359f \
 //x=2.31 //y=1.45 //x2=3.015 //y2=0.995
cc_981 ( N_CLK_c_1163_p N_noxref_12_M1_noxref_d ) capacitor c=0.00223875f \
 //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_982 ( N_CLK_c_1165_p N_noxref_12_M1_noxref_d ) capacitor c=0.00262485f \
 //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_983 ( N_CLK_c_1189_p N_noxref_12_M1_noxref_d ) capacitor c=0.00220746f \
 //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_984 ( N_CLK_c_1196_p N_noxref_12_M1_noxref_d ) capacitor c=0.00194798f \
 //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_985 ( N_CLK_c_1059_n N_noxref_12_M1_noxref_d ) capacitor c=0.00198465f \
 //x=2.31 //y=0.91 //x2=1.86 //y2=0.91
cc_986 ( N_CLK_c_1060_n N_noxref_12_M1_noxref_d ) capacitor c=0.00128384f \
 //x=2.31 //y=1.22 //x2=1.86 //y2=0.91
cc_987 ( N_CLK_c_1059_n N_noxref_12_M2_noxref_s ) capacitor c=7.21316e-19 \
 //x=2.31 //y=0.91 //x2=2.965 //y2=0.375
cc_988 ( N_CLK_c_1060_n N_noxref_12_M2_noxref_s ) capacitor c=0.00348171f \
 //x=2.31 //y=1.22 //x2=2.965 //y2=0.375
cc_989 ( N_CLK_c_1011_n N_D_c_2523_n ) capacitor c=0.0210462f //x=15.055 \
 //y=4.44 //x2=7.03 //y2=2.08
cc_990 ( N_CLK_c_1011_n N_D_c_2537_n ) capacitor c=0.0085986f //x=15.055 \
 //y=4.44 //x2=7.365 //y2=4.79
cc_991 ( N_CLK_c_1011_n N_D_c_2538_n ) capacitor c=0.00293313f //x=15.055 \
 //y=4.44 //x2=7.03 //y2=4.7
cc_992 ( N_CLK_c_1082_n N_noxref_17_c_2766_n ) capacitor c=0.0167228f \
 //x=14.735 //y=0.91 //x2=15.395 //y2=0.54
cc_993 ( N_CLK_c_1087_n N_noxref_17_c_2766_n ) capacitor c=0.00534519f \
 //x=15.26 //y=0.91 //x2=15.395 //y2=0.54
cc_994 ( N_CLK_c_1010_n N_noxref_17_c_2789_n ) capacitor c=0.0120267f \
 //x=15.17 //y=2.08 //x2=15.395 //y2=1.59
cc_995 ( N_CLK_c_1085_n N_noxref_17_c_2789_n ) capacitor c=0.0157358f \
 //x=14.735 //y=1.22 //x2=15.395 //y2=1.59
cc_996 ( N_CLK_c_1090_n N_noxref_17_c_2789_n ) capacitor c=0.021347f //x=15.26 \
 //y=1.915 //x2=15.395 //y2=1.59
cc_997 ( N_CLK_c_1082_n N_noxref_17_M8_noxref_s ) capacitor c=0.00798959f \
 //x=14.735 //y=0.91 //x2=13.405 //y2=0.375
cc_998 ( N_CLK_c_1089_n N_noxref_17_M8_noxref_s ) capacitor c=0.00212176f \
 //x=15.26 //y=1.45 //x2=13.405 //y2=0.375
cc_999 ( N_CLK_c_1090_n N_noxref_17_M8_noxref_s ) capacitor c=0.00298115f \
 //x=15.26 //y=1.915 //x2=13.405 //y2=0.375
cc_1000 ( N_CLK_c_1212_p N_noxref_18_c_2809_n ) capacitor c=2.14837e-19 \
 //x=15.105 //y=0.755 //x2=15.965 //y2=0.995
cc_1001 ( N_CLK_c_1087_n N_noxref_18_c_2809_n ) capacitor c=0.00123426f \
 //x=15.26 //y=0.91 //x2=15.965 //y2=0.995
cc_1002 ( N_CLK_c_1088_n N_noxref_18_c_2809_n ) capacitor c=0.0129288f \
 //x=15.26 //y=1.22 //x2=15.965 //y2=0.995
cc_1003 ( N_CLK_c_1089_n N_noxref_18_c_2809_n ) capacitor c=0.00142359f \
 //x=15.26 //y=1.45 //x2=15.965 //y2=0.995
cc_1004 ( N_CLK_c_1082_n N_noxref_18_M9_noxref_d ) capacitor c=0.00223875f \
 //x=14.735 //y=0.91 //x2=14.81 //y2=0.91
cc_1005 ( N_CLK_c_1085_n N_noxref_18_M9_noxref_d ) capacitor c=0.00262485f \
 //x=14.735 //y=1.22 //x2=14.81 //y2=0.91
cc_1006 ( N_CLK_c_1212_p N_noxref_18_M9_noxref_d ) capacitor c=0.00220746f \
 //x=15.105 //y=0.755 //x2=14.81 //y2=0.91
cc_1007 ( N_CLK_c_1219_p N_noxref_18_M9_noxref_d ) capacitor c=0.00194798f \
 //x=15.105 //y=1.375 //x2=14.81 //y2=0.91
cc_1008 ( N_CLK_c_1087_n N_noxref_18_M9_noxref_d ) capacitor c=0.00198465f \
 //x=15.26 //y=0.91 //x2=14.81 //y2=0.91
cc_1009 ( N_CLK_c_1088_n N_noxref_18_M9_noxref_d ) capacitor c=0.00128384f \
 //x=15.26 //y=1.22 //x2=14.81 //y2=0.91
cc_1010 ( N_CLK_c_1087_n N_noxref_18_M10_noxref_s ) capacitor c=7.21316e-19 \
 //x=15.26 //y=0.91 //x2=15.915 //y2=0.375
cc_1011 ( N_CLK_c_1088_n N_noxref_18_M10_noxref_s ) capacitor c=0.00348171f \
 //x=15.26 //y=1.22 //x2=15.915 //y2=0.375
cc_1012 ( N_noxref_6_c_1224_n N_RN_c_1470_n ) capacitor c=0.0824003f \
 //x=18.755 //y=3.7 //x2=16.165 //y2=2.22
cc_1013 ( N_noxref_6_c_1224_n N_RN_c_1478_n ) capacitor c=4.865e-19 //x=18.755 \
 //y=3.7 //x2=8.255 //y2=2.22
cc_1014 ( N_noxref_6_c_1224_n N_RN_c_1480_n ) capacitor c=0.055674f //x=18.755 \
 //y=3.7 //x2=19.865 //y2=2.22
cc_1015 ( N_noxref_6_c_1227_n N_RN_c_1480_n ) capacitor c=0.0251492f //x=18.87 \
 //y=2.08 //x2=19.865 //y2=2.22
cc_1016 ( N_noxref_6_c_1242_n N_RN_c_1480_n ) capacitor c=0.0106236f //x=18.57 \
 //y=1.915 //x2=19.865 //y2=2.22
cc_1017 ( N_noxref_6_c_1224_n N_RN_c_1484_n ) capacitor c=0.00444609f \
 //x=18.755 //y=3.7 //x2=16.395 //y2=2.22
cc_1018 ( N_noxref_6_c_1224_n N_RN_c_1485_n ) capacitor c=0.0179999f \
 //x=18.755 //y=3.7 //x2=8.14 //y2=2.08
cc_1019 ( N_noxref_6_c_1226_n N_RN_c_1485_n ) capacitor c=0.00108603f //x=5.92 \
 //y=2.08 //x2=8.14 //y2=2.08
cc_1020 ( N_noxref_6_c_1224_n N_RN_c_1486_n ) capacitor c=0.022876f //x=18.755 \
 //y=3.7 //x2=16.28 //y2=2.08
cc_1021 ( N_noxref_6_c_1227_n N_RN_c_1486_n ) capacitor c=8.87185e-19 \
 //x=18.87 //y=2.08 //x2=16.28 //y2=2.08
cc_1022 ( N_noxref_6_c_1224_n N_RN_c_1487_n ) capacitor c=0.0027353f \
 //x=18.755 //y=3.7 //x2=19.98 //y2=2.08
cc_1023 ( N_noxref_6_c_1227_n N_RN_c_1487_n ) capacitor c=0.0521309f //x=18.87 \
 //y=2.08 //x2=19.98 //y2=2.08
cc_1024 ( N_noxref_6_c_1242_n N_RN_c_1487_n ) capacitor c=0.00208635f \
 //x=18.57 //y=1.915 //x2=19.98 //y2=2.08
cc_1025 ( N_noxref_6_c_1373_p N_RN_c_1487_n ) capacitor c=0.00147352f \
 //x=19.435 //y=4.79 //x2=19.98 //y2=2.08
cc_1026 ( N_noxref_6_c_1280_n N_RN_c_1487_n ) capacitor c=0.00142741f \
 //x=19.145 //y=4.79 //x2=19.98 //y2=2.08
cc_1027 ( N_noxref_6_M38_noxref_g N_RN_M40_noxref_g ) capacitor c=0.0105869f \
 //x=19.07 //y=6.02 //x2=19.95 //y2=6.02
cc_1028 ( N_noxref_6_M39_noxref_g N_RN_M40_noxref_g ) capacitor c=0.10632f \
 //x=19.51 //y=6.02 //x2=19.95 //y2=6.02
cc_1029 ( N_noxref_6_M39_noxref_g N_RN_M41_noxref_g ) capacitor c=0.0101598f \
 //x=19.51 //y=6.02 //x2=20.39 //y2=6.02
cc_1030 ( N_noxref_6_c_1238_n N_RN_c_1584_n ) capacitor c=5.72482e-19 \
 //x=18.57 //y=0.875 //x2=19.545 //y2=0.91
cc_1031 ( N_noxref_6_c_1240_n N_RN_c_1584_n ) capacitor c=0.00149976f \
 //x=18.57 //y=1.22 //x2=19.545 //y2=0.91
cc_1032 ( N_noxref_6_c_1245_n N_RN_c_1584_n ) capacitor c=0.0160123f //x=19.1 \
 //y=0.875 //x2=19.545 //y2=0.91
cc_1033 ( N_noxref_6_c_1241_n N_RN_c_1587_n ) capacitor c=0.00111227f \
 //x=18.57 //y=1.53 //x2=19.545 //y2=1.22
cc_1034 ( N_noxref_6_c_1247_n N_RN_c_1587_n ) capacitor c=0.0124075f //x=19.1 \
 //y=1.22 //x2=19.545 //y2=1.22
cc_1035 ( N_noxref_6_c_1245_n N_RN_c_1589_n ) capacitor c=0.00103227f //x=19.1 \
 //y=0.875 //x2=20.07 //y2=0.91
cc_1036 ( N_noxref_6_c_1247_n N_RN_c_1590_n ) capacitor c=0.0010154f //x=19.1 \
 //y=1.22 //x2=20.07 //y2=1.22
cc_1037 ( N_noxref_6_c_1247_n N_RN_c_1591_n ) capacitor c=9.23422e-19 //x=19.1 \
 //y=1.22 //x2=20.07 //y2=1.45
cc_1038 ( N_noxref_6_c_1227_n N_RN_c_1592_n ) capacitor c=0.00203769f \
 //x=18.87 //y=2.08 //x2=20.07 //y2=1.915
cc_1039 ( N_noxref_6_c_1242_n N_RN_c_1592_n ) capacitor c=0.00834532f \
 //x=18.57 //y=1.915 //x2=20.07 //y2=1.915
cc_1040 ( N_noxref_6_c_1227_n N_RN_c_1594_n ) capacitor c=0.00183762f \
 //x=18.87 //y=2.08 //x2=19.98 //y2=4.7
cc_1041 ( N_noxref_6_c_1373_p N_RN_c_1594_n ) capacitor c=0.0168581f \
 //x=19.435 //y=4.79 //x2=19.98 //y2=4.7
cc_1042 ( N_noxref_6_c_1280_n N_RN_c_1594_n ) capacitor c=0.00484466f \
 //x=19.145 //y=4.79 //x2=19.98 //y2=4.7
cc_1043 ( N_noxref_6_M39_noxref_g N_QN_c_1758_n ) capacitor c=0.0178794f \
 //x=19.51 //y=6.02 //x2=20.085 //y2=5.155
cc_1044 ( N_noxref_6_M38_noxref_g N_QN_c_1762_n ) capacitor c=0.0213876f \
 //x=19.07 //y=6.02 //x2=19.375 //y2=5.155
cc_1045 ( N_noxref_6_c_1373_p N_QN_c_1762_n ) capacitor c=0.00429591f \
 //x=19.435 //y=4.79 //x2=19.375 //y2=5.155
cc_1046 ( N_noxref_6_M39_noxref_g N_QN_M38_noxref_d ) capacitor c=0.0180032f \
 //x=19.51 //y=6.02 //x2=19.145 //y2=5.02
cc_1047 ( N_noxref_6_c_1297_n N_noxref_9_c_1895_n ) capacitor c=0.147447f \
 //x=5.805 //y=3.7 //x2=11.355 //y2=4.07
cc_1048 ( N_noxref_6_c_1298_n N_noxref_9_c_1895_n ) capacitor c=0.0294294f \
 //x=4.185 //y=3.7 //x2=11.355 //y2=4.07
cc_1049 ( N_noxref_6_c_1224_n N_noxref_9_c_1895_n ) capacitor c=0.467539f \
 //x=18.755 //y=3.7 //x2=11.355 //y2=4.07
cc_1050 ( N_noxref_6_c_1305_n N_noxref_9_c_1895_n ) capacitor c=0.0264476f \
 //x=6.035 //y=3.7 //x2=11.355 //y2=4.07
cc_1051 ( N_noxref_6_c_1253_n N_noxref_9_c_1895_n ) capacitor c=0.0154449f \
 //x=1.615 //y=5.155 //x2=11.355 //y2=4.07
cc_1052 ( N_noxref_6_c_1263_n N_noxref_9_c_1895_n ) capacitor c=0.0200328f \
 //x=4.07 //y=3.7 //x2=11.355 //y2=4.07
cc_1053 ( N_noxref_6_c_1226_n N_noxref_9_c_1895_n ) capacitor c=0.0213516f \
 //x=5.92 //y=2.08 //x2=11.355 //y2=4.07
cc_1054 ( N_noxref_6_c_1224_n N_noxref_9_c_1922_n ) capacitor c=0.468066f \
 //x=18.755 //y=3.7 //x2=16.905 //y2=4.07
cc_1055 ( N_noxref_6_c_1224_n N_noxref_9_c_1998_n ) capacitor c=0.0267832f \
 //x=18.755 //y=3.7 //x2=11.585 //y2=4.07
cc_1056 ( N_noxref_6_c_1224_n N_noxref_9_c_1897_n ) capacitor c=0.176507f \
 //x=18.755 //y=3.7 //x2=24.305 //y2=4.07
cc_1057 ( N_noxref_6_c_1227_n N_noxref_9_c_1897_n ) capacitor c=0.0252746f \
 //x=18.87 //y=2.08 //x2=24.305 //y2=4.07
cc_1058 ( N_noxref_6_c_1280_n N_noxref_9_c_1897_n ) capacitor c=0.0115418f \
 //x=19.145 //y=4.79 //x2=24.305 //y2=4.07
cc_1059 ( N_noxref_6_c_1224_n N_noxref_9_c_1935_n ) capacitor c=0.0268461f \
 //x=18.755 //y=3.7 //x2=17.135 //y2=4.07
cc_1060 ( N_noxref_6_c_1227_n N_noxref_9_c_1935_n ) capacitor c=3.50683e-19 \
 //x=18.87 //y=2.08 //x2=17.135 //y2=4.07
cc_1061 ( N_noxref_6_c_1224_n N_noxref_9_c_1899_n ) capacitor c=0.0236433f \
 //x=18.755 //y=3.7 //x2=11.47 //y2=2.08
cc_1062 ( N_noxref_6_c_1224_n N_noxref_9_c_1957_n ) capacitor c=0.0261231f \
 //x=18.755 //y=3.7 //x2=17.02 //y2=4.07
cc_1063 ( N_noxref_6_c_1227_n N_noxref_9_c_1957_n ) capacitor c=0.0144739f \
 //x=18.87 //y=2.08 //x2=17.02 //y2=4.07
cc_1064 ( N_noxref_6_c_1253_n N_noxref_9_M16_noxref_g ) capacitor c=0.0213876f \
 //x=1.615 //y=5.155 //x2=1.31 //y2=6.02
cc_1065 ( N_noxref_6_c_1249_n N_noxref_9_M17_noxref_g ) capacitor c=0.0178794f \
 //x=2.325 //y=5.155 //x2=1.75 //y2=6.02
cc_1066 ( N_noxref_6_M16_noxref_d N_noxref_9_M17_noxref_g ) capacitor \
 c=0.0180032f //x=1.385 //y=5.02 //x2=1.75 //y2=6.02
cc_1067 ( N_noxref_6_c_1253_n N_noxref_9_c_2095_n ) capacitor c=0.00429591f \
 //x=1.615 //y=5.155 //x2=1.675 //y2=4.79
cc_1068 ( N_noxref_6_c_1224_n N_noxref_10_c_2280_n ) capacitor c=0.00740361f \
 //x=18.755 //y=3.7 //x2=21.205 //y2=3.7
cc_1069 ( N_noxref_6_c_1227_n N_noxref_10_c_2281_n ) capacitor c=0.00138947f \
 //x=18.87 //y=2.08 //x2=21.09 //y2=2.08
cc_1070 ( N_noxref_6_M2_noxref_d N_noxref_11_M0_noxref_s ) capacitor \
 c=0.00309936f //x=3.395 //y=0.915 //x2=0.455 //y2=0.375
cc_1071 ( N_noxref_6_c_1225_n N_noxref_12_c_2475_n ) capacitor c=0.00466084f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_1072 ( N_noxref_6_M2_noxref_d N_noxref_12_c_2475_n ) capacitor c=0.0117786f \
 //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_1073 ( N_noxref_6_c_1312_n N_noxref_12_c_2489_n ) capacitor c=0.0200405f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_1074 ( N_noxref_6_M2_noxref_d N_noxref_12_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_1075 ( N_noxref_6_c_1225_n N_noxref_12_M2_noxref_s ) capacitor c=0.0207678f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_1076 ( N_noxref_6_M2_noxref_d N_noxref_12_M2_noxref_s ) capacitor \
 c=0.0426368f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
cc_1077 ( N_noxref_6_c_1224_n N_D_c_2523_n ) capacitor c=0.0190398f //x=18.755 \
 //y=3.7 //x2=7.03 //y2=2.08
cc_1078 ( N_noxref_6_c_1305_n N_D_c_2523_n ) capacitor c=9.95819e-19 //x=6.035 \
 //y=3.7 //x2=7.03 //y2=2.08
cc_1079 ( N_noxref_6_c_1263_n N_D_c_2523_n ) capacitor c=4.0219e-19 //x=4.07 \
 //y=3.7 //x2=7.03 //y2=2.08
cc_1080 ( N_noxref_6_c_1226_n N_D_c_2523_n ) capacitor c=0.048337f //x=5.92 \
 //y=2.08 //x2=7.03 //y2=2.08
cc_1081 ( N_noxref_6_c_1232_n N_D_c_2523_n ) capacitor c=0.00238338f //x=5.62 \
 //y=1.915 //x2=7.03 //y2=2.08
cc_1082 ( N_noxref_6_c_1326_n N_D_c_2523_n ) capacitor c=0.00147352f //x=6.485 \
 //y=4.79 //x2=7.03 //y2=2.08
cc_1083 ( N_noxref_6_c_1278_n N_D_c_2523_n ) capacitor c=0.00142741f //x=6.195 \
 //y=4.79 //x2=7.03 //y2=2.08
cc_1084 ( N_noxref_6_M22_noxref_g N_D_M24_noxref_g ) capacitor c=0.0105869f \
 //x=6.12 //y=6.02 //x2=7 //y2=6.02
cc_1085 ( N_noxref_6_M23_noxref_g N_D_M24_noxref_g ) capacitor c=0.10632f \
 //x=6.56 //y=6.02 //x2=7 //y2=6.02
cc_1086 ( N_noxref_6_M23_noxref_g N_D_M25_noxref_g ) capacitor c=0.0101598f \
 //x=6.56 //y=6.02 //x2=7.44 //y2=6.02
cc_1087 ( N_noxref_6_c_1228_n N_D_c_2552_n ) capacitor c=5.72482e-19 //x=5.62 \
 //y=0.875 //x2=6.595 //y2=0.91
cc_1088 ( N_noxref_6_c_1230_n N_D_c_2552_n ) capacitor c=0.00149976f //x=5.62 \
 //y=1.22 //x2=6.595 //y2=0.91
cc_1089 ( N_noxref_6_c_1235_n N_D_c_2552_n ) capacitor c=0.0160123f //x=6.15 \
 //y=0.875 //x2=6.595 //y2=0.91
cc_1090 ( N_noxref_6_c_1231_n N_D_c_2555_n ) capacitor c=0.00111227f //x=5.62 \
 //y=1.53 //x2=6.595 //y2=1.22
cc_1091 ( N_noxref_6_c_1237_n N_D_c_2555_n ) capacitor c=0.0124075f //x=6.15 \
 //y=1.22 //x2=6.595 //y2=1.22
cc_1092 ( N_noxref_6_c_1235_n N_D_c_2557_n ) capacitor c=0.00103227f //x=6.15 \
 //y=0.875 //x2=7.12 //y2=0.91
cc_1093 ( N_noxref_6_c_1237_n N_D_c_2558_n ) capacitor c=0.0010154f //x=6.15 \
 //y=1.22 //x2=7.12 //y2=1.22
cc_1094 ( N_noxref_6_c_1237_n N_D_c_2559_n ) capacitor c=9.23422e-19 //x=6.15 \
 //y=1.22 //x2=7.12 //y2=1.45
cc_1095 ( N_noxref_6_c_1226_n N_D_c_2560_n ) capacitor c=0.00231304f //x=5.92 \
 //y=2.08 //x2=7.12 //y2=1.915
cc_1096 ( N_noxref_6_c_1232_n N_D_c_2560_n ) capacitor c=0.00964411f //x=5.62 \
 //y=1.915 //x2=7.12 //y2=1.915
cc_1097 ( N_noxref_6_c_1226_n N_D_c_2538_n ) capacitor c=0.00183762f //x=5.92 \
 //y=2.08 //x2=7.03 //y2=4.7
cc_1098 ( N_noxref_6_c_1326_n N_D_c_2538_n ) capacitor c=0.0168581f //x=6.485 \
 //y=4.79 //x2=7.03 //y2=4.7
cc_1099 ( N_noxref_6_c_1278_n N_D_c_2538_n ) capacitor c=0.00484466f //x=6.195 \
 //y=4.79 //x2=7.03 //y2=4.7
cc_1100 ( N_noxref_6_c_1225_n N_noxref_14_c_2619_n ) capacitor c=3.84569e-19 \
 //x=3.985 //y=1.665 //x2=5.4 //y2=1.505
cc_1101 ( N_noxref_6_c_1232_n N_noxref_14_c_2619_n ) capacitor c=0.0034165f \
 //x=5.62 //y=1.915 //x2=5.4 //y2=1.505
cc_1102 ( N_noxref_6_c_1226_n N_noxref_14_c_2603_n ) capacitor c=0.0125801f \
 //x=5.92 //y=2.08 //x2=6.285 //y2=1.59
cc_1103 ( N_noxref_6_c_1231_n N_noxref_14_c_2603_n ) capacitor c=0.00703864f \
 //x=5.62 //y=1.53 //x2=6.285 //y2=1.59
cc_1104 ( N_noxref_6_c_1232_n N_noxref_14_c_2603_n ) capacitor c=0.0245895f \
 //x=5.62 //y=1.915 //x2=6.285 //y2=1.59
cc_1105 ( N_noxref_6_c_1234_n N_noxref_14_c_2603_n ) capacitor c=0.00708583f \
 //x=5.995 //y=1.375 //x2=6.285 //y2=1.59
cc_1106 ( N_noxref_6_c_1237_n N_noxref_14_c_2603_n ) capacitor c=0.00698822f \
 //x=6.15 //y=1.22 //x2=6.285 //y2=1.59
cc_1107 ( N_noxref_6_c_1228_n N_noxref_14_M3_noxref_s ) capacitor c=0.0327271f \
 //x=5.62 //y=0.875 //x2=5.265 //y2=0.375
cc_1108 ( N_noxref_6_c_1231_n N_noxref_14_M3_noxref_s ) capacitor \
 c=7.99997e-19 //x=5.62 //y=1.53 //x2=5.265 //y2=0.375
cc_1109 ( N_noxref_6_c_1232_n N_noxref_14_M3_noxref_s ) capacitor \
 c=0.00122123f //x=5.62 //y=1.915 //x2=5.265 //y2=0.375
cc_1110 ( N_noxref_6_c_1235_n N_noxref_14_M3_noxref_s ) capacitor c=0.0121427f \
 //x=6.15 //y=0.875 //x2=5.265 //y2=0.375
cc_1111 ( N_noxref_6_M2_noxref_d N_noxref_14_M3_noxref_s ) capacitor \
 c=2.55333e-19 //x=3.395 //y=0.915 //x2=5.265 //y2=0.375
cc_1112 ( N_noxref_6_c_1242_n N_noxref_19_c_2879_n ) capacitor c=0.0034165f \
 //x=18.57 //y=1.915 //x2=18.35 //y2=1.505
cc_1113 ( N_noxref_6_c_1227_n N_noxref_19_c_2863_n ) capacitor c=0.0119952f \
 //x=18.87 //y=2.08 //x2=19.235 //y2=1.59
cc_1114 ( N_noxref_6_c_1241_n N_noxref_19_c_2863_n ) capacitor c=0.00697148f \
 //x=18.57 //y=1.53 //x2=19.235 //y2=1.59
cc_1115 ( N_noxref_6_c_1242_n N_noxref_19_c_2863_n ) capacitor c=0.0204849f \
 //x=18.57 //y=1.915 //x2=19.235 //y2=1.59
cc_1116 ( N_noxref_6_c_1244_n N_noxref_19_c_2863_n ) capacitor c=0.00610316f \
 //x=18.945 //y=1.375 //x2=19.235 //y2=1.59
cc_1117 ( N_noxref_6_c_1247_n N_noxref_19_c_2863_n ) capacitor c=0.00698822f \
 //x=19.1 //y=1.22 //x2=19.235 //y2=1.59
cc_1118 ( N_noxref_6_c_1238_n N_noxref_19_M11_noxref_s ) capacitor \
 c=0.0327271f //x=18.57 //y=0.875 //x2=18.215 //y2=0.375
cc_1119 ( N_noxref_6_c_1241_n N_noxref_19_M11_noxref_s ) capacitor \
 c=7.99997e-19 //x=18.57 //y=1.53 //x2=18.215 //y2=0.375
cc_1120 ( N_noxref_6_c_1242_n N_noxref_19_M11_noxref_s ) capacitor \
 c=0.00122123f //x=18.57 //y=1.915 //x2=18.215 //y2=0.375
cc_1121 ( N_noxref_6_c_1245_n N_noxref_19_M11_noxref_s ) capacitor \
 c=0.0121427f //x=19.1 //y=0.875 //x2=18.215 //y2=0.375
cc_1122 ( N_RN_c_1487_n QN ) capacitor c=0.00330955f //x=19.98 //y=2.08 \
 //x2=21.83 //y2=2.22
cc_1123 ( N_RN_c_1487_n N_QN_c_1758_n ) capacitor c=0.0148665f //x=19.98 \
 //y=2.08 //x2=20.085 //y2=5.155
cc_1124 ( N_RN_M40_noxref_g N_QN_c_1758_n ) capacitor c=0.0166659f //x=19.95 \
 //y=6.02 //x2=20.085 //y2=5.155
cc_1125 ( N_RN_c_1594_n N_QN_c_1758_n ) capacitor c=0.00322396f //x=19.98 \
 //y=4.7 //x2=20.085 //y2=5.155
cc_1126 ( N_RN_M41_noxref_g N_QN_c_1764_n ) capacitor c=0.0184045f //x=20.39 \
 //y=6.02 //x2=20.965 //y2=5.155
cc_1127 ( N_RN_c_1602_p N_QN_c_1804_n ) capacitor c=0.00427862f //x=20.315 \
 //y=4.79 //x2=20.17 //y2=5.155
cc_1128 ( N_RN_M40_noxref_g N_QN_M40_noxref_d ) capacitor c=0.0180032f \
 //x=19.95 //y=6.02 //x2=20.025 //y2=5.02
cc_1129 ( N_RN_M41_noxref_g N_QN_M40_noxref_d ) capacitor c=0.0180032f \
 //x=20.39 //y=6.02 //x2=20.025 //y2=5.02
cc_1130 ( N_RN_c_1470_n N_noxref_9_c_1895_n ) capacitor c=0.00314955f \
 //x=16.165 //y=2.22 //x2=11.355 //y2=4.07
cc_1131 ( N_RN_c_1485_n N_noxref_9_c_1895_n ) capacitor c=0.0179722f //x=8.14 \
 //y=2.08 //x2=11.355 //y2=4.07
cc_1132 ( N_RN_c_1470_n N_noxref_9_c_1922_n ) capacitor c=0.014344f //x=16.165 \
 //y=2.22 //x2=16.905 //y2=4.07
cc_1133 ( N_RN_c_1480_n N_noxref_9_c_1922_n ) capacitor c=0.0031797f \
 //x=19.865 //y=2.22 //x2=16.905 //y2=4.07
cc_1134 ( N_RN_c_1484_n N_noxref_9_c_1922_n ) capacitor c=2.19189e-19 \
 //x=16.395 //y=2.22 //x2=16.905 //y2=4.07
cc_1135 ( N_RN_c_1486_n N_noxref_9_c_1922_n ) capacitor c=0.0219145f //x=16.28 \
 //y=2.08 //x2=16.905 //y2=4.07
cc_1136 ( N_RN_c_1563_n N_noxref_9_c_1922_n ) capacitor c=0.00881004f \
 //x=16.28 //y=4.7 //x2=16.905 //y2=4.07
cc_1137 ( N_RN_c_1470_n N_noxref_9_c_1998_n ) capacitor c=2.80052e-19 \
 //x=16.165 //y=2.22 //x2=11.585 //y2=4.07
cc_1138 ( N_RN_c_1480_n N_noxref_9_c_1897_n ) capacitor c=0.0254729f \
 //x=19.865 //y=2.22 //x2=24.305 //y2=4.07
cc_1139 ( N_RN_c_1487_n N_noxref_9_c_1897_n ) capacitor c=0.0283962f //x=19.98 \
 //y=2.08 //x2=24.305 //y2=4.07
cc_1140 ( N_RN_c_1602_p N_noxref_9_c_1897_n ) capacitor c=0.00495688f \
 //x=20.315 //y=4.79 //x2=24.305 //y2=4.07
cc_1141 ( N_RN_c_1594_n N_noxref_9_c_1897_n ) capacitor c=0.0018068f //x=19.98 \
 //y=4.7 //x2=24.305 //y2=4.07
cc_1142 ( N_RN_c_1480_n N_noxref_9_c_1935_n ) capacitor c=2.98411e-19 \
 //x=19.865 //y=2.22 //x2=17.135 //y2=4.07
cc_1143 ( N_RN_c_1486_n N_noxref_9_c_1935_n ) capacitor c=0.00179385f \
 //x=16.28 //y=2.08 //x2=17.135 //y2=4.07
cc_1144 ( N_RN_c_1470_n N_noxref_9_c_1899_n ) capacitor c=0.0226984f \
 //x=16.165 //y=2.22 //x2=11.47 //y2=2.08
cc_1145 ( N_RN_M36_noxref_g N_noxref_9_c_1949_n ) capacitor c=0.0184045f \
 //x=16.02 //y=6.02 //x2=16.155 //y2=5.155
cc_1146 ( N_RN_M37_noxref_g N_noxref_9_c_1953_n ) capacitor c=0.0205426f \
 //x=16.46 //y=6.02 //x2=16.935 //y2=5.155
cc_1147 ( N_RN_c_1563_n N_noxref_9_c_1953_n ) capacitor c=0.00201851f \
 //x=16.28 //y=4.7 //x2=16.935 //y2=5.155
cc_1148 ( N_RN_c_1623_p N_noxref_9_c_1901_n ) capacitor c=0.00371277f \
 //x=16.645 //y=1.415 //x2=16.935 //y2=1.665
cc_1149 ( N_RN_c_1624_p N_noxref_9_c_1901_n ) capacitor c=0.00457401f //x=16.8 \
 //y=1.26 //x2=16.935 //y2=1.665
cc_1150 ( N_RN_c_1480_n N_noxref_9_c_2144_n ) capacitor c=0.016327f //x=19.865 \
 //y=2.22 //x2=16.62 //y2=1.665
cc_1151 ( N_RN_c_1480_n N_noxref_9_c_1957_n ) capacitor c=0.0245777f \
 //x=19.865 //y=2.22 //x2=17.02 //y2=4.07
cc_1152 ( N_RN_c_1484_n N_noxref_9_c_1957_n ) capacitor c=0.0012045f \
 //x=16.395 //y=2.22 //x2=17.02 //y2=4.07
cc_1153 ( N_RN_c_1486_n N_noxref_9_c_1957_n ) capacitor c=0.0847926f //x=16.28 \
 //y=2.08 //x2=17.02 //y2=4.07
cc_1154 ( N_RN_c_1487_n N_noxref_9_c_1957_n ) capacitor c=7.03136e-19 \
 //x=19.98 //y=2.08 //x2=17.02 //y2=4.07
cc_1155 ( N_RN_c_1560_n N_noxref_9_c_1957_n ) capacitor c=0.00709342f \
 //x=16.28 //y=2.08 //x2=17.02 //y2=4.07
cc_1156 ( N_RN_c_1562_n N_noxref_9_c_1957_n ) capacitor c=0.00283672f \
 //x=16.28 //y=1.915 //x2=17.02 //y2=4.07
cc_1157 ( N_RN_c_1563_n N_noxref_9_c_1957_n ) capacitor c=0.013693f //x=16.28 \
 //y=4.7 //x2=17.02 //y2=4.07
cc_1158 ( N_RN_c_1486_n N_noxref_9_c_2152_n ) capacitor c=0.0174995f //x=16.28 \
 //y=2.08 //x2=16.24 //y2=5.155
cc_1159 ( N_RN_c_1563_n N_noxref_9_c_2152_n ) capacitor c=0.00475729f \
 //x=16.28 //y=4.7 //x2=16.24 //y2=5.155
cc_1160 ( N_RN_c_1470_n N_noxref_9_c_2047_n ) capacitor c=3.11115e-19 \
 //x=16.165 //y=2.22 //x2=11.88 //y2=1.405
cc_1161 ( N_RN_c_1470_n N_noxref_9_c_2019_n ) capacitor c=0.00571486f \
 //x=16.165 //y=2.22 //x2=11.47 //y2=2.08
cc_1162 ( N_RN_c_1556_n N_noxref_9_M10_noxref_d ) capacitor c=0.00217566f \
 //x=16.27 //y=0.915 //x2=16.345 //y2=0.915
cc_1163 ( N_RN_c_1557_n N_noxref_9_M10_noxref_d ) capacitor c=0.0034598f \
 //x=16.27 //y=1.26 //x2=16.345 //y2=0.915
cc_1164 ( N_RN_c_1558_n N_noxref_9_M10_noxref_d ) capacitor c=0.00546784f \
 //x=16.27 //y=1.57 //x2=16.345 //y2=0.915
cc_1165 ( N_RN_c_1640_p N_noxref_9_M10_noxref_d ) capacitor c=0.00241102f \
 //x=16.645 //y=0.76 //x2=16.345 //y2=0.915
cc_1166 ( N_RN_c_1623_p N_noxref_9_M10_noxref_d ) capacitor c=0.0138621f \
 //x=16.645 //y=1.415 //x2=16.345 //y2=0.915
cc_1167 ( N_RN_c_1642_p N_noxref_9_M10_noxref_d ) capacitor c=0.00219619f \
 //x=16.8 //y=0.915 //x2=16.345 //y2=0.915
cc_1168 ( N_RN_c_1624_p N_noxref_9_M10_noxref_d ) capacitor c=0.00603828f \
 //x=16.8 //y=1.26 //x2=16.345 //y2=0.915
cc_1169 ( N_RN_c_1562_n N_noxref_9_M10_noxref_d ) capacitor c=0.00661782f \
 //x=16.28 //y=1.915 //x2=16.345 //y2=0.915
cc_1170 ( N_RN_M36_noxref_g N_noxref_9_M36_noxref_d ) capacitor c=0.0180032f \
 //x=16.02 //y=6.02 //x2=16.095 //y2=5.02
cc_1171 ( N_RN_M37_noxref_g N_noxref_9_M36_noxref_d ) capacitor c=0.0194246f \
 //x=16.46 //y=6.02 //x2=16.095 //y2=5.02
cc_1172 ( N_RN_c_1487_n N_noxref_10_c_2280_n ) capacitor c=0.00273375f \
 //x=19.98 //y=2.08 //x2=21.205 //y2=3.7
cc_1173 ( N_RN_c_1480_n N_noxref_10_c_2281_n ) capacitor c=0.00558344f \
 //x=19.865 //y=2.22 //x2=21.09 //y2=2.08
cc_1174 ( N_RN_c_1487_n N_noxref_10_c_2281_n ) capacitor c=0.0527626f \
 //x=19.98 //y=2.08 //x2=21.09 //y2=2.08
cc_1175 ( N_RN_c_1592_n N_noxref_10_c_2281_n ) capacitor c=0.00213841f \
 //x=20.07 //y=1.915 //x2=21.09 //y2=2.08
cc_1176 ( N_RN_c_1594_n N_noxref_10_c_2281_n ) capacitor c=0.00142741f \
 //x=19.98 //y=4.7 //x2=21.09 //y2=2.08
cc_1177 ( N_RN_M40_noxref_g N_noxref_10_M42_noxref_g ) capacitor c=0.0101598f \
 //x=19.95 //y=6.02 //x2=20.83 //y2=6.02
cc_1178 ( N_RN_M41_noxref_g N_noxref_10_M42_noxref_g ) capacitor c=0.0602553f \
 //x=20.39 //y=6.02 //x2=20.83 //y2=6.02
cc_1179 ( N_RN_M41_noxref_g N_noxref_10_M43_noxref_g ) capacitor c=0.0101598f \
 //x=20.39 //y=6.02 //x2=21.27 //y2=6.02
cc_1180 ( N_RN_c_1589_n N_noxref_10_c_2325_n ) capacitor c=0.00456962f \
 //x=20.07 //y=0.91 //x2=21.08 //y2=0.915
cc_1181 ( N_RN_c_1590_n N_noxref_10_c_2326_n ) capacitor c=0.00438372f \
 //x=20.07 //y=1.22 //x2=21.08 //y2=1.26
cc_1182 ( N_RN_c_1591_n N_noxref_10_c_2327_n ) capacitor c=0.00438372f \
 //x=20.07 //y=1.45 //x2=21.08 //y2=1.57
cc_1183 ( N_RN_c_1480_n N_noxref_10_c_2328_n ) capacitor c=0.00341397f \
 //x=19.865 //y=2.22 //x2=21.09 //y2=2.08
cc_1184 ( N_RN_c_1487_n N_noxref_10_c_2328_n ) capacitor c=0.0021852f \
 //x=19.98 //y=2.08 //x2=21.09 //y2=2.08
cc_1185 ( N_RN_c_1592_n N_noxref_10_c_2328_n ) capacitor c=0.00896806f \
 //x=20.07 //y=1.915 //x2=21.09 //y2=2.08
cc_1186 ( N_RN_c_1592_n N_noxref_10_c_2331_n ) capacitor c=0.00438372f \
 //x=20.07 //y=1.915 //x2=21.09 //y2=1.915
cc_1187 ( N_RN_c_1487_n N_noxref_10_c_2332_n ) capacitor c=0.00219458f \
 //x=19.98 //y=2.08 //x2=21.09 //y2=4.7
cc_1188 ( N_RN_c_1602_p N_noxref_10_c_2332_n ) capacitor c=0.0611812f \
 //x=20.315 //y=4.79 //x2=21.09 //y2=4.7
cc_1189 ( N_RN_c_1594_n N_noxref_10_c_2332_n ) capacitor c=0.00487508f \
 //x=19.98 //y=4.7 //x2=21.09 //y2=4.7
cc_1190 ( N_RN_c_1478_n N_D_c_2523_n ) capacitor c=0.00558344f //x=8.255 \
 //y=2.22 //x2=7.03 //y2=2.08
cc_1191 ( N_RN_c_1485_n N_D_c_2523_n ) capacitor c=0.0471413f //x=8.14 \
 //y=2.08 //x2=7.03 //y2=2.08
cc_1192 ( N_RN_c_1531_n N_D_c_2523_n ) capacitor c=0.00209043f //x=8.14 \
 //y=2.08 //x2=7.03 //y2=2.08
cc_1193 ( N_RN_c_1534_n N_D_c_2523_n ) capacitor c=0.00219458f //x=8.14 \
 //y=4.7 //x2=7.03 //y2=2.08
cc_1194 ( N_RN_M26_noxref_g N_D_M24_noxref_g ) capacitor c=0.0101598f //x=7.88 \
 //y=6.02 //x2=7 //y2=6.02
cc_1195 ( N_RN_M26_noxref_g N_D_M25_noxref_g ) capacitor c=0.0602553f //x=7.88 \
 //y=6.02 //x2=7.44 //y2=6.02
cc_1196 ( N_RN_M27_noxref_g N_D_M25_noxref_g ) capacitor c=0.0101598f //x=8.32 \
 //y=6.02 //x2=7.44 //y2=6.02
cc_1197 ( N_RN_c_1522_n N_D_c_2557_n ) capacitor c=0.00456962f //x=8.13 \
 //y=0.915 //x2=7.12 //y2=0.91
cc_1198 ( N_RN_c_1523_n N_D_c_2558_n ) capacitor c=0.00438372f //x=8.13 \
 //y=1.26 //x2=7.12 //y2=1.22
cc_1199 ( N_RN_c_1524_n N_D_c_2559_n ) capacitor c=0.00438372f //x=8.13 \
 //y=1.57 //x2=7.12 //y2=1.45
cc_1200 ( N_RN_c_1478_n N_D_c_2560_n ) capacitor c=0.00341397f //x=8.255 \
 //y=2.22 //x2=7.12 //y2=1.915
cc_1201 ( N_RN_c_1485_n N_D_c_2560_n ) capacitor c=0.00223318f //x=8.14 \
 //y=2.08 //x2=7.12 //y2=1.915
cc_1202 ( N_RN_c_1531_n N_D_c_2560_n ) capacitor c=0.00881982f //x=8.14 \
 //y=2.08 //x2=7.12 //y2=1.915
cc_1203 ( N_RN_c_1532_n N_D_c_2560_n ) capacitor c=0.00438372f //x=8.14 \
 //y=1.915 //x2=7.12 //y2=1.915
cc_1204 ( N_RN_c_1534_n N_D_c_2537_n ) capacitor c=0.0611812f //x=8.14 //y=4.7 \
 //x2=7.365 //y2=4.79
cc_1205 ( N_RN_c_1485_n N_D_c_2538_n ) capacitor c=0.00142741f //x=8.14 \
 //y=2.08 //x2=7.03 //y2=4.7
cc_1206 ( N_RN_c_1534_n N_D_c_2538_n ) capacitor c=0.00487508f //x=8.14 \
 //y=4.7 //x2=7.03 //y2=4.7
cc_1207 ( N_RN_c_1470_n N_noxref_15_c_2658_n ) capacitor c=7.41833e-19 \
 //x=16.165 //y=2.22 //x2=8.795 //y2=0.54
cc_1208 ( N_RN_c_1478_n N_noxref_15_c_2658_n ) capacitor c=7.4531e-19 \
 //x=8.255 //y=2.22 //x2=8.795 //y2=0.54
cc_1209 ( N_RN_c_1485_n N_noxref_15_c_2658_n ) capacitor c=0.00204178f \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_1210 ( N_RN_c_1522_n N_noxref_15_c_2658_n ) capacitor c=0.0194423f //x=8.13 \
 //y=0.915 //x2=8.795 //y2=0.54
cc_1211 ( N_RN_c_1528_n N_noxref_15_c_2658_n ) capacitor c=0.00656458f \
 //x=8.66 //y=0.915 //x2=8.795 //y2=0.54
cc_1212 ( N_RN_c_1531_n N_noxref_15_c_2658_n ) capacitor c=2.20712e-19 \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_1213 ( N_RN_c_1523_n N_noxref_15_c_2670_n ) capacitor c=0.00538829f \
 //x=8.13 //y=1.26 //x2=7.91 //y2=0.995
cc_1214 ( N_RN_c_1522_n N_noxref_15_M5_noxref_s ) capacitor c=0.00538829f \
 //x=8.13 //y=0.915 //x2=7.775 //y2=0.375
cc_1215 ( N_RN_c_1524_n N_noxref_15_M5_noxref_s ) capacitor c=0.00538829f \
 //x=8.13 //y=1.57 //x2=7.775 //y2=0.375
cc_1216 ( N_RN_c_1528_n N_noxref_15_M5_noxref_s ) capacitor c=0.0143002f \
 //x=8.66 //y=0.915 //x2=7.775 //y2=0.375
cc_1217 ( N_RN_c_1529_n N_noxref_15_M5_noxref_s ) capacitor c=0.00290153f \
 //x=8.66 //y=1.26 //x2=7.775 //y2=0.375
cc_1218 ( N_RN_c_1470_n N_noxref_16_c_2726_n ) capacitor c=0.00635755f \
 //x=16.165 //y=2.22 //x2=10.315 //y2=1.495
cc_1219 ( N_RN_c_1470_n N_noxref_16_c_2707_n ) capacitor c=0.0223494f \
 //x=16.165 //y=2.22 //x2=11.2 //y2=1.58
cc_1220 ( N_RN_c_1470_n N_noxref_16_c_2714_n ) capacitor c=0.00649228f \
 //x=16.165 //y=2.22 //x2=11.285 //y2=1.495
cc_1221 ( N_RN_c_1470_n N_noxref_16_c_2715_n ) capacitor c=0.00178534f \
 //x=16.165 //y=2.22 //x2=12.17 //y2=0.53
cc_1222 ( N_RN_c_1470_n N_noxref_16_M6_noxref_s ) capacitor c=0.00113237f \
 //x=16.165 //y=2.22 //x2=10.18 //y2=0.365
cc_1223 ( N_RN_c_1470_n N_noxref_17_c_2775_n ) capacitor c=0.00642985f \
 //x=16.165 //y=2.22 //x2=13.54 //y2=1.505
cc_1224 ( N_RN_c_1470_n N_noxref_17_c_2759_n ) capacitor c=0.0225733f \
 //x=16.165 //y=2.22 //x2=14.425 //y2=1.59
cc_1225 ( N_RN_c_1470_n N_noxref_17_c_2789_n ) capacitor c=0.0203655f \
 //x=16.165 //y=2.22 //x2=15.395 //y2=1.59
cc_1226 ( N_RN_c_1470_n N_noxref_17_M8_noxref_s ) capacitor c=0.012425f \
 //x=16.165 //y=2.22 //x2=13.405 //y2=0.375
cc_1227 ( N_RN_c_1470_n N_noxref_18_c_2809_n ) capacitor c=0.00657782f \
 //x=16.165 //y=2.22 //x2=15.965 //y2=0.995
cc_1228 ( N_RN_c_1480_n N_noxref_18_c_2814_n ) capacitor c=7.41833e-19 \
 //x=19.865 //y=2.22 //x2=16.935 //y2=0.54
cc_1229 ( N_RN_c_1484_n N_noxref_18_c_2814_n ) capacitor c=7.4531e-19 \
 //x=16.395 //y=2.22 //x2=16.935 //y2=0.54
cc_1230 ( N_RN_c_1486_n N_noxref_18_c_2814_n ) capacitor c=0.00204178f \
 //x=16.28 //y=2.08 //x2=16.935 //y2=0.54
cc_1231 ( N_RN_c_1556_n N_noxref_18_c_2814_n ) capacitor c=0.0194423f \
 //x=16.27 //y=0.915 //x2=16.935 //y2=0.54
cc_1232 ( N_RN_c_1642_p N_noxref_18_c_2814_n ) capacitor c=0.00656458f \
 //x=16.8 //y=0.915 //x2=16.935 //y2=0.54
cc_1233 ( N_RN_c_1560_n N_noxref_18_c_2814_n ) capacitor c=2.20712e-19 \
 //x=16.28 //y=2.08 //x2=16.935 //y2=0.54
cc_1234 ( N_RN_c_1557_n N_noxref_18_c_2842_n ) capacitor c=0.00538829f \
 //x=16.27 //y=1.26 //x2=16.05 //y2=0.995
cc_1235 ( N_RN_c_1470_n N_noxref_18_M10_noxref_s ) capacitor c=0.00642985f \
 //x=16.165 //y=2.22 //x2=15.915 //y2=0.375
cc_1236 ( N_RN_c_1556_n N_noxref_18_M10_noxref_s ) capacitor c=0.00538829f \
 //x=16.27 //y=0.915 //x2=15.915 //y2=0.375
cc_1237 ( N_RN_c_1558_n N_noxref_18_M10_noxref_s ) capacitor c=0.00538829f \
 //x=16.27 //y=1.57 //x2=15.915 //y2=0.375
cc_1238 ( N_RN_c_1642_p N_noxref_18_M10_noxref_s ) capacitor c=0.0143002f \
 //x=16.8 //y=0.915 //x2=15.915 //y2=0.375
cc_1239 ( N_RN_c_1624_p N_noxref_18_M10_noxref_s ) capacitor c=0.00290153f \
 //x=16.8 //y=1.26 //x2=15.915 //y2=0.375
cc_1240 ( N_RN_c_1480_n N_noxref_19_c_2879_n ) capacitor c=0.00642985f \
 //x=19.865 //y=2.22 //x2=18.35 //y2=1.505
cc_1241 ( N_RN_c_1480_n N_noxref_19_c_2863_n ) capacitor c=0.0225733f \
 //x=19.865 //y=2.22 //x2=19.235 //y2=1.59
cc_1242 ( N_RN_c_1584_n N_noxref_19_c_2870_n ) capacitor c=0.0167228f \
 //x=19.545 //y=0.91 //x2=20.205 //y2=0.54
cc_1243 ( N_RN_c_1589_n N_noxref_19_c_2870_n ) capacitor c=0.00534519f \
 //x=20.07 //y=0.91 //x2=20.205 //y2=0.54
cc_1244 ( N_RN_c_1480_n N_noxref_19_c_2893_n ) capacitor c=0.0178105f \
 //x=19.865 //y=2.22 //x2=20.205 //y2=1.59
cc_1245 ( N_RN_c_1487_n N_noxref_19_c_2893_n ) capacitor c=0.0119919f \
 //x=19.98 //y=2.08 //x2=20.205 //y2=1.59
cc_1246 ( N_RN_c_1587_n N_noxref_19_c_2893_n ) capacitor c=0.0157358f \
 //x=19.545 //y=1.22 //x2=20.205 //y2=1.59
cc_1247 ( N_RN_c_1592_n N_noxref_19_c_2893_n ) capacitor c=0.0217576f \
 //x=20.07 //y=1.915 //x2=20.205 //y2=1.59
cc_1248 ( N_RN_c_1480_n N_noxref_19_M11_noxref_s ) capacitor c=0.00642985f \
 //x=19.865 //y=2.22 //x2=18.215 //y2=0.375
cc_1249 ( N_RN_c_1584_n N_noxref_19_M11_noxref_s ) capacitor c=0.00798959f \
 //x=19.545 //y=0.91 //x2=18.215 //y2=0.375
cc_1250 ( N_RN_c_1591_n N_noxref_19_M11_noxref_s ) capacitor c=0.00212176f \
 //x=20.07 //y=1.45 //x2=18.215 //y2=0.375
cc_1251 ( N_RN_c_1592_n N_noxref_19_M11_noxref_s ) capacitor c=0.00298115f \
 //x=20.07 //y=1.915 //x2=18.215 //y2=0.375
cc_1252 ( N_RN_c_1727_p N_noxref_20_c_2915_n ) capacitor c=2.14837e-19 \
 //x=19.915 //y=0.755 //x2=20.775 //y2=0.995
cc_1253 ( N_RN_c_1589_n N_noxref_20_c_2915_n ) capacitor c=0.00123426f \
 //x=20.07 //y=0.91 //x2=20.775 //y2=0.995
cc_1254 ( N_RN_c_1590_n N_noxref_20_c_2915_n ) capacitor c=0.0129288f \
 //x=20.07 //y=1.22 //x2=20.775 //y2=0.995
cc_1255 ( N_RN_c_1591_n N_noxref_20_c_2915_n ) capacitor c=0.00142359f \
 //x=20.07 //y=1.45 //x2=20.775 //y2=0.995
cc_1256 ( N_RN_c_1584_n N_noxref_20_M12_noxref_d ) capacitor c=0.00223875f \
 //x=19.545 //y=0.91 //x2=19.62 //y2=0.91
cc_1257 ( N_RN_c_1587_n N_noxref_20_M12_noxref_d ) capacitor c=0.00262485f \
 //x=19.545 //y=1.22 //x2=19.62 //y2=0.91
cc_1258 ( N_RN_c_1727_p N_noxref_20_M12_noxref_d ) capacitor c=0.00220746f \
 //x=19.915 //y=0.755 //x2=19.62 //y2=0.91
cc_1259 ( N_RN_c_1734_p N_noxref_20_M12_noxref_d ) capacitor c=0.00194798f \
 //x=19.915 //y=1.375 //x2=19.62 //y2=0.91
cc_1260 ( N_RN_c_1589_n N_noxref_20_M12_noxref_d ) capacitor c=0.00198465f \
 //x=20.07 //y=0.91 //x2=19.62 //y2=0.91
cc_1261 ( N_RN_c_1590_n N_noxref_20_M12_noxref_d ) capacitor c=0.00128384f \
 //x=20.07 //y=1.22 //x2=19.62 //y2=0.91
cc_1262 ( N_RN_c_1589_n N_noxref_20_M13_noxref_s ) capacitor c=7.21316e-19 \
 //x=20.07 //y=0.91 //x2=20.725 //y2=0.375
cc_1263 ( N_RN_c_1590_n N_noxref_20_M13_noxref_s ) capacitor c=0.00348171f \
 //x=20.07 //y=1.22 //x2=20.725 //y2=0.375
cc_1264 ( N_QN_c_1739_n N_noxref_9_c_1897_n ) capacitor c=0.010979f //x=23.565 \
 //y=3.33 //x2=24.305 //y2=4.07
cc_1265 ( N_QN_c_1743_n N_noxref_9_c_1897_n ) capacitor c=7.97799e-19 \
 //x=21.945 //y=3.33 //x2=24.305 //y2=4.07
cc_1266 ( QN N_noxref_9_c_1897_n ) capacitor c=0.0232727f //x=21.83 //y=2.22 \
 //x2=24.305 //y2=4.07
cc_1267 ( N_QN_c_1758_n N_noxref_9_c_1897_n ) capacitor c=0.0239852f \
 //x=20.085 //y=5.155 //x2=24.305 //y2=4.07
cc_1268 ( N_QN_c_1762_n N_noxref_9_c_1897_n ) capacitor c=0.0173f //x=19.375 \
 //y=5.155 //x2=24.305 //y2=4.07
cc_1269 ( N_QN_c_1768_n N_noxref_9_c_1897_n ) capacitor c=0.0138556f \
 //x=21.745 //y=5.155 //x2=24.305 //y2=4.07
cc_1270 ( N_QN_c_1745_n N_noxref_9_c_1897_n ) capacitor c=0.0242126f //x=23.68 \
 //y=2.08 //x2=24.305 //y2=4.07
cc_1271 ( N_QN_c_1779_n N_noxref_9_c_1897_n ) capacitor c=0.00844647f \
 //x=23.68 //y=4.7 //x2=24.305 //y2=4.07
cc_1272 ( N_QN_c_1762_n N_noxref_9_c_1953_n ) capacitor c=3.10026e-19 \
 //x=19.375 //y=5.155 //x2=16.935 //y2=5.155
cc_1273 ( N_QN_c_1745_n N_noxref_9_c_2175_n ) capacitor c=0.00400249f \
 //x=23.68 //y=2.08 //x2=24.42 //y2=4.535
cc_1274 ( N_QN_c_1779_n N_noxref_9_c_2175_n ) capacitor c=0.00417994f \
 //x=23.68 //y=4.7 //x2=24.42 //y2=4.535
cc_1275 ( N_QN_c_1739_n N_noxref_9_c_1902_n ) capacitor c=0.00720056f \
 //x=23.565 //y=3.33 //x2=24.42 //y2=2.08
cc_1276 ( QN N_noxref_9_c_1902_n ) capacitor c=0.00107361f //x=21.83 //y=2.22 \
 //x2=24.42 //y2=2.08
cc_1277 ( N_QN_c_1745_n N_noxref_9_c_1902_n ) capacitor c=0.0810987f //x=23.68 \
 //y=2.08 //x2=24.42 //y2=2.08
cc_1278 ( N_QN_c_1750_n N_noxref_9_c_1902_n ) capacitor c=0.00308814f \
 //x=23.485 //y=1.915 //x2=24.42 //y2=2.08
cc_1279 ( N_QN_M44_noxref_g N_noxref_9_M46_noxref_g ) capacitor c=0.0104611f \
 //x=23.58 //y=6.02 //x2=24.46 //y2=6.02
cc_1280 ( N_QN_M45_noxref_g N_noxref_9_M46_noxref_g ) capacitor c=0.106811f \
 //x=24.02 //y=6.02 //x2=24.46 //y2=6.02
cc_1281 ( N_QN_M45_noxref_g N_noxref_9_M47_noxref_g ) capacitor c=0.0100341f \
 //x=24.02 //y=6.02 //x2=24.9 //y2=6.02
cc_1282 ( N_QN_c_1746_n N_noxref_9_c_2184_n ) capacitor c=4.86506e-19 \
 //x=23.485 //y=0.865 //x2=24.455 //y2=0.905
cc_1283 ( N_QN_c_1748_n N_noxref_9_c_2184_n ) capacitor c=0.00152104f \
 //x=23.485 //y=1.21 //x2=24.455 //y2=0.905
cc_1284 ( N_QN_c_1753_n N_noxref_9_c_2184_n ) capacitor c=0.0151475f \
 //x=24.015 //y=0.865 //x2=24.455 //y2=0.905
cc_1285 ( N_QN_c_1749_n N_noxref_9_c_2187_n ) capacitor c=0.00109982f \
 //x=23.485 //y=1.52 //x2=24.455 //y2=1.25
cc_1286 ( N_QN_c_1755_n N_noxref_9_c_2187_n ) capacitor c=0.0111064f \
 //x=24.015 //y=1.21 //x2=24.455 //y2=1.25
cc_1287 ( N_QN_c_1749_n N_noxref_9_c_2189_n ) capacitor c=9.57794e-19 \
 //x=23.485 //y=1.52 //x2=24.455 //y2=1.56
cc_1288 ( N_QN_c_1750_n N_noxref_9_c_2189_n ) capacitor c=0.00662747f \
 //x=23.485 //y=1.915 //x2=24.455 //y2=1.56
cc_1289 ( N_QN_c_1755_n N_noxref_9_c_2189_n ) capacitor c=0.00862358f \
 //x=24.015 //y=1.21 //x2=24.455 //y2=1.56
cc_1290 ( N_QN_c_1753_n N_noxref_9_c_2192_n ) capacitor c=0.00124821f \
 //x=24.015 //y=0.865 //x2=24.985 //y2=0.905
cc_1291 ( N_QN_c_1755_n N_noxref_9_c_2193_n ) capacitor c=0.00200715f \
 //x=24.015 //y=1.21 //x2=24.985 //y2=1.25
cc_1292 ( N_QN_c_1745_n N_noxref_9_c_2194_n ) capacitor c=0.00307062f \
 //x=23.68 //y=2.08 //x2=24.42 //y2=2.08
cc_1293 ( N_QN_c_1750_n N_noxref_9_c_2194_n ) capacitor c=0.0179092f \
 //x=23.485 //y=1.915 //x2=24.42 //y2=2.08
cc_1294 ( N_QN_c_1745_n N_noxref_9_c_2196_n ) capacitor c=0.00344981f \
 //x=23.68 //y=2.08 //x2=24.45 //y2=4.7
cc_1295 ( N_QN_c_1779_n N_noxref_9_c_2196_n ) capacitor c=0.0293367f //x=23.68 \
 //y=4.7 //x2=24.45 //y2=4.7
cc_1296 ( N_QN_c_1739_n N_noxref_10_c_2279_n ) capacitor c=0.175734f \
 //x=23.565 //y=3.33 //x2=25.045 //y2=3.7
cc_1297 ( N_QN_c_1743_n N_noxref_10_c_2279_n ) capacitor c=0.029467f \
 //x=21.945 //y=3.33 //x2=25.045 //y2=3.7
cc_1298 ( QN N_noxref_10_c_2279_n ) capacitor c=0.0206044f //x=21.83 //y=2.22 \
 //x2=25.045 //y2=3.7
cc_1299 ( N_QN_c_1842_p N_noxref_10_c_2279_n ) capacitor c=0.0042996f \
 //x=21.43 //y=1.665 //x2=25.045 //y2=3.7
cc_1300 ( N_QN_c_1745_n N_noxref_10_c_2279_n ) capacitor c=0.0205569f \
 //x=23.68 //y=2.08 //x2=25.045 //y2=3.7
cc_1301 ( QN N_noxref_10_c_2280_n ) capacitor c=0.00117715f //x=21.83 //y=2.22 \
 //x2=21.205 //y2=3.7
cc_1302 ( N_QN_c_1743_n N_noxref_10_c_2281_n ) capacitor c=0.00720056f \
 //x=21.945 //y=3.33 //x2=21.09 //y2=2.08
cc_1303 ( QN N_noxref_10_c_2281_n ) capacitor c=0.0854964f //x=21.83 //y=2.22 \
 //x2=21.09 //y2=2.08
cc_1304 ( N_QN_c_1745_n N_noxref_10_c_2281_n ) capacitor c=0.001003f //x=23.68 \
 //y=2.08 //x2=21.09 //y2=2.08
cc_1305 ( N_QN_c_1848_p N_noxref_10_c_2281_n ) capacitor c=0.0168082f \
 //x=21.05 //y=5.155 //x2=21.09 //y2=2.08
cc_1306 ( N_QN_M45_noxref_g N_noxref_10_c_2290_n ) capacitor c=0.017965f \
 //x=24.02 //y=6.02 //x2=24.595 //y2=5.2
cc_1307 ( N_QN_c_1745_n N_noxref_10_c_2294_n ) capacitor c=0.00549854f \
 //x=23.68 //y=2.08 //x2=23.885 //y2=5.2
cc_1308 ( N_QN_M44_noxref_g N_noxref_10_c_2294_n ) capacitor c=0.0177326f \
 //x=23.58 //y=6.02 //x2=23.885 //y2=5.2
cc_1309 ( N_QN_c_1779_n N_noxref_10_c_2294_n ) capacitor c=0.00582246f \
 //x=23.68 //y=4.7 //x2=23.885 //y2=5.2
cc_1310 ( QN N_noxref_10_c_2283_n ) capacitor c=3.52729e-19 //x=21.83 //y=2.22 \
 //x2=25.16 //y2=3.7
cc_1311 ( N_QN_c_1745_n N_noxref_10_c_2283_n ) capacitor c=0.00407494f \
 //x=23.68 //y=2.08 //x2=25.16 //y2=3.7
cc_1312 ( N_QN_c_1764_n N_noxref_10_M42_noxref_g ) capacitor c=0.0184045f \
 //x=20.965 //y=5.155 //x2=20.83 //y2=6.02
cc_1313 ( N_QN_M42_noxref_d N_noxref_10_M42_noxref_g ) capacitor c=0.0180032f \
 //x=20.905 //y=5.02 //x2=20.83 //y2=6.02
cc_1314 ( N_QN_c_1768_n N_noxref_10_M43_noxref_g ) capacitor c=0.0205426f \
 //x=21.745 //y=5.155 //x2=21.27 //y2=6.02
cc_1315 ( N_QN_M42_noxref_d N_noxref_10_M43_noxref_g ) capacitor c=0.0194246f \
 //x=20.905 //y=5.02 //x2=21.27 //y2=6.02
cc_1316 ( N_QN_M13_noxref_d N_noxref_10_c_2325_n ) capacitor c=0.00217566f \
 //x=21.155 //y=0.915 //x2=21.08 //y2=0.915
cc_1317 ( N_QN_M13_noxref_d N_noxref_10_c_2326_n ) capacitor c=0.0034598f \
 //x=21.155 //y=0.915 //x2=21.08 //y2=1.26
cc_1318 ( N_QN_M13_noxref_d N_noxref_10_c_2327_n ) capacitor c=0.00544291f \
 //x=21.155 //y=0.915 //x2=21.08 //y2=1.57
cc_1319 ( N_QN_M13_noxref_d N_noxref_10_c_2358_n ) capacitor c=0.00241102f \
 //x=21.155 //y=0.915 //x2=21.455 //y2=0.76
cc_1320 ( N_QN_c_1744_n N_noxref_10_c_2359_n ) capacitor c=0.00359704f \
 //x=21.745 //y=1.665 //x2=21.455 //y2=1.415
cc_1321 ( N_QN_M13_noxref_d N_noxref_10_c_2359_n ) capacitor c=0.0140297f \
 //x=21.155 //y=0.915 //x2=21.455 //y2=1.415
cc_1322 ( N_QN_M13_noxref_d N_noxref_10_c_2361_n ) capacitor c=0.00219619f \
 //x=21.155 //y=0.915 //x2=21.61 //y2=0.915
cc_1323 ( N_QN_c_1744_n N_noxref_10_c_2362_n ) capacitor c=0.00457401f \
 //x=21.745 //y=1.665 //x2=21.61 //y2=1.26
cc_1324 ( N_QN_M13_noxref_d N_noxref_10_c_2362_n ) capacitor c=0.00603828f \
 //x=21.155 //y=0.915 //x2=21.61 //y2=1.26
cc_1325 ( QN N_noxref_10_c_2328_n ) capacitor c=0.00772308f //x=21.83 //y=2.22 \
 //x2=21.09 //y2=2.08
cc_1326 ( QN N_noxref_10_c_2331_n ) capacitor c=0.00283672f //x=21.83 //y=2.22 \
 //x2=21.09 //y2=1.915
cc_1327 ( N_QN_M13_noxref_d N_noxref_10_c_2331_n ) capacitor c=0.00661782f \
 //x=21.155 //y=0.915 //x2=21.09 //y2=1.915
cc_1328 ( QN N_noxref_10_c_2332_n ) capacitor c=0.013844f //x=21.83 //y=2.22 \
 //x2=21.09 //y2=4.7
cc_1329 ( N_QN_c_1768_n N_noxref_10_c_2332_n ) capacitor c=0.00201851f \
 //x=21.745 //y=5.155 //x2=21.09 //y2=4.7
cc_1330 ( N_QN_c_1848_p N_noxref_10_c_2332_n ) capacitor c=0.00475729f \
 //x=21.05 //y=5.155 //x2=21.09 //y2=4.7
cc_1331 ( N_QN_M45_noxref_g N_noxref_10_M44_noxref_d ) capacitor c=0.0173476f \
 //x=24.02 //y=6.02 //x2=23.655 //y2=5.02
cc_1332 ( N_QN_M13_noxref_d N_noxref_19_M11_noxref_s ) capacitor c=0.00309936f \
 //x=21.155 //y=0.915 //x2=18.215 //y2=0.375
cc_1333 ( N_QN_c_1744_n N_noxref_20_c_2920_n ) capacitor c=0.00467185f \
 //x=21.745 //y=1.665 //x2=21.745 //y2=0.54
cc_1334 ( N_QN_M13_noxref_d N_noxref_20_c_2920_n ) capacitor c=0.0118029f \
 //x=21.155 //y=0.915 //x2=21.745 //y2=0.54
cc_1335 ( N_QN_c_1842_p N_noxref_20_c_2943_n ) capacitor c=0.020048f //x=21.43 \
 //y=1.665 //x2=20.86 //y2=0.995
cc_1336 ( N_QN_M13_noxref_d N_noxref_20_M12_noxref_d ) capacitor c=5.27807e-19 \
 //x=21.155 //y=0.915 //x2=19.62 //y2=0.91
cc_1337 ( N_QN_c_1744_n N_noxref_20_M13_noxref_s ) capacitor c=0.020752f \
 //x=21.745 //y=1.665 //x2=20.725 //y2=0.375
cc_1338 ( N_QN_M13_noxref_d N_noxref_20_M13_noxref_s ) capacitor c=0.0426444f \
 //x=21.155 //y=0.915 //x2=20.725 //y2=0.375
cc_1339 ( N_QN_c_1739_n N_noxref_21_c_2984_n ) capacitor c=0.00241565f \
 //x=23.565 //y=3.33 //x2=23.265 //y2=1.495
cc_1340 ( N_QN_c_1744_n N_noxref_21_c_2984_n ) capacitor c=3.04182e-19 \
 //x=21.745 //y=1.665 //x2=23.265 //y2=1.495
cc_1341 ( N_QN_c_1750_n N_noxref_21_c_2984_n ) capacitor c=0.0034165f \
 //x=23.485 //y=1.915 //x2=23.265 //y2=1.495
cc_1342 ( N_QN_c_1739_n N_noxref_21_c_2967_n ) capacitor c=0.00649414f \
 //x=23.565 //y=3.33 //x2=24.15 //y2=1.58
cc_1343 ( N_QN_c_1745_n N_noxref_21_c_2967_n ) capacitor c=0.011692f //x=23.68 \
 //y=2.08 //x2=24.15 //y2=1.58
cc_1344 ( N_QN_c_1749_n N_noxref_21_c_2967_n ) capacitor c=0.00703567f \
 //x=23.485 //y=1.52 //x2=24.15 //y2=1.58
cc_1345 ( N_QN_c_1750_n N_noxref_21_c_2967_n ) capacitor c=0.0203514f \
 //x=23.485 //y=1.915 //x2=24.15 //y2=1.58
cc_1346 ( N_QN_c_1752_n N_noxref_21_c_2967_n ) capacitor c=0.00780629f \
 //x=23.86 //y=1.365 //x2=24.15 //y2=1.58
cc_1347 ( N_QN_c_1755_n N_noxref_21_c_2967_n ) capacitor c=0.00339872f \
 //x=24.015 //y=1.21 //x2=24.15 //y2=1.58
cc_1348 ( N_QN_c_1750_n N_noxref_21_c_2974_n ) capacitor c=6.71402e-19 \
 //x=23.485 //y=1.915 //x2=24.235 //y2=1.495
cc_1349 ( N_QN_c_1746_n N_noxref_21_M14_noxref_s ) capacitor c=0.0327502f \
 //x=23.485 //y=0.865 //x2=23.13 //y2=0.365
cc_1350 ( N_QN_c_1749_n N_noxref_21_M14_noxref_s ) capacitor c=3.48408e-19 \
 //x=23.485 //y=1.52 //x2=23.13 //y2=0.365
cc_1351 ( N_QN_c_1753_n N_noxref_21_M14_noxref_s ) capacitor c=0.0120759f \
 //x=24.015 //y=0.865 //x2=23.13 //y2=0.365
cc_1352 ( N_noxref_9_c_1897_n N_noxref_10_c_2279_n ) capacitor c=0.3045f \
 //x=24.305 //y=4.07 //x2=25.045 //y2=3.7
cc_1353 ( N_noxref_9_c_1902_n N_noxref_10_c_2279_n ) capacitor c=0.0255669f \
 //x=24.42 //y=2.08 //x2=25.045 //y2=3.7
cc_1354 ( N_noxref_9_c_2200_p N_noxref_10_c_2279_n ) capacitor c=0.00624857f \
 //x=24.825 //y=4.79 //x2=25.045 //y2=3.7
cc_1355 ( N_noxref_9_c_2196_n N_noxref_10_c_2279_n ) capacitor c=3.27069e-19 \
 //x=24.45 //y=4.7 //x2=25.045 //y2=3.7
cc_1356 ( N_noxref_9_c_1897_n N_noxref_10_c_2280_n ) capacitor c=0.0292842f \
 //x=24.305 //y=4.07 //x2=21.205 //y2=3.7
cc_1357 ( N_noxref_9_c_1897_n N_noxref_10_c_2281_n ) capacitor c=0.0237491f \
 //x=24.305 //y=4.07 //x2=21.09 //y2=2.08
cc_1358 ( N_noxref_9_c_1897_n N_noxref_10_c_2290_n ) capacitor c=0.00208151f \
 //x=24.305 //y=4.07 //x2=24.595 //y2=5.2
cc_1359 ( N_noxref_9_c_2175_n N_noxref_10_c_2290_n ) capacitor c=0.0129205f \
 //x=24.42 //y=4.535 //x2=24.595 //y2=5.2
cc_1360 ( N_noxref_9_M46_noxref_g N_noxref_10_c_2290_n ) capacitor \
 c=0.0166421f //x=24.46 //y=6.02 //x2=24.595 //y2=5.2
cc_1361 ( N_noxref_9_c_2196_n N_noxref_10_c_2290_n ) capacitor c=0.00346627f \
 //x=24.45 //y=4.7 //x2=24.595 //y2=5.2
cc_1362 ( N_noxref_9_c_1897_n N_noxref_10_c_2294_n ) capacitor c=0.01319f \
 //x=24.305 //y=4.07 //x2=23.885 //y2=5.2
cc_1363 ( N_noxref_9_M47_noxref_g N_noxref_10_c_2296_n ) capacitor \
 c=0.0206783f //x=24.9 //y=6.02 //x2=25.075 //y2=5.2
cc_1364 ( N_noxref_9_c_2210_p N_noxref_10_c_2282_n ) capacitor c=0.00359704f \
 //x=24.83 //y=1.405 //x2=25.075 //y2=1.655
cc_1365 ( N_noxref_9_c_2193_n N_noxref_10_c_2282_n ) capacitor c=0.00457401f \
 //x=24.985 //y=1.25 //x2=25.075 //y2=1.655
cc_1366 ( N_noxref_9_c_1897_n N_noxref_10_c_2283_n ) capacitor c=0.00642908f \
 //x=24.305 //y=4.07 //x2=25.16 //y2=3.7
cc_1367 ( N_noxref_9_c_2175_n N_noxref_10_c_2283_n ) capacitor c=0.0101115f \
 //x=24.42 //y=4.535 //x2=25.16 //y2=3.7
cc_1368 ( N_noxref_9_c_1902_n N_noxref_10_c_2283_n ) capacitor c=0.0786723f \
 //x=24.42 //y=2.08 //x2=25.16 //y2=3.7
cc_1369 ( N_noxref_9_c_2200_p N_noxref_10_c_2283_n ) capacitor c=0.0142673f \
 //x=24.825 //y=4.79 //x2=25.16 //y2=3.7
cc_1370 ( N_noxref_9_c_2194_n N_noxref_10_c_2283_n ) capacitor c=0.00877984f \
 //x=24.42 //y=2.08 //x2=25.16 //y2=3.7
cc_1371 ( N_noxref_9_c_2217_p N_noxref_10_c_2283_n ) capacitor c=0.00306024f \
 //x=24.42 //y=1.915 //x2=25.16 //y2=3.7
cc_1372 ( N_noxref_9_c_2196_n N_noxref_10_c_2283_n ) capacitor c=0.00533692f \
 //x=24.45 //y=4.7 //x2=25.16 //y2=3.7
cc_1373 ( N_noxref_9_c_2200_p N_noxref_10_c_2392_n ) capacitor c=0.00421574f \
 //x=24.825 //y=4.79 //x2=24.68 //y2=5.2
cc_1374 ( N_noxref_9_c_1897_n N_noxref_10_c_2332_n ) capacitor c=0.00775263f \
 //x=24.305 //y=4.07 //x2=21.09 //y2=4.7
cc_1375 ( N_noxref_9_c_2184_n N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00217566f //x=24.455 //y=0.905 //x2=24.53 //y2=0.905
cc_1376 ( N_noxref_9_c_2187_n N_noxref_10_M15_noxref_d ) capacitor \
 c=0.0034598f //x=24.455 //y=1.25 //x2=24.53 //y2=0.905
cc_1377 ( N_noxref_9_c_2189_n N_noxref_10_M15_noxref_d ) capacitor \
 c=0.0065582f //x=24.455 //y=1.56 //x2=24.53 //y2=0.905
cc_1378 ( N_noxref_9_c_2224_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00241102f //x=24.83 //y=0.75 //x2=24.53 //y2=0.905
cc_1379 ( N_noxref_9_c_2210_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.0138845f //x=24.83 //y=1.405 //x2=24.53 //y2=0.905
cc_1380 ( N_noxref_9_c_2192_n N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00132245f //x=24.985 //y=0.905 //x2=24.53 //y2=0.905
cc_1381 ( N_noxref_9_c_2193_n N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00566463f //x=24.985 //y=1.25 //x2=24.53 //y2=0.905
cc_1382 ( N_noxref_9_c_2217_p N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00660593f //x=24.42 //y=1.915 //x2=24.53 //y2=0.905
cc_1383 ( N_noxref_9_M46_noxref_g N_noxref_10_M46_noxref_d ) capacitor \
 c=0.0173476f //x=24.46 //y=6.02 //x2=24.535 //y2=5.02
cc_1384 ( N_noxref_9_M47_noxref_g N_noxref_10_M46_noxref_d ) capacitor \
 c=0.0179769f //x=24.9 //y=6.02 //x2=24.535 //y2=5.02
cc_1385 ( N_noxref_9_c_1908_n N_noxref_11_c_2448_n ) capacitor c=0.0034165f \
 //x=0.81 //y=1.915 //x2=0.59 //y2=1.505
cc_1386 ( N_noxref_9_c_1895_n N_noxref_11_c_2423_n ) capacitor c=0.00179505f \
 //x=11.355 //y=4.07 //x2=1.475 //y2=1.59
cc_1387 ( N_noxref_9_c_1896_n N_noxref_11_c_2423_n ) capacitor c=0.00102628f \
 //x=1.225 //y=4.07 //x2=1.475 //y2=1.59
cc_1388 ( N_noxref_9_c_1898_n N_noxref_11_c_2423_n ) capacitor c=0.0122033f \
 //x=1.11 //y=2.08 //x2=1.475 //y2=1.59
cc_1389 ( N_noxref_9_c_1907_n N_noxref_11_c_2423_n ) capacitor c=0.00703864f \
 //x=0.81 //y=1.53 //x2=1.475 //y2=1.59
cc_1390 ( N_noxref_9_c_1908_n N_noxref_11_c_2423_n ) capacitor c=0.0259045f \
 //x=0.81 //y=1.915 //x2=1.475 //y2=1.59
cc_1391 ( N_noxref_9_c_1910_n N_noxref_11_c_2423_n ) capacitor c=0.00708583f \
 //x=1.185 //y=1.375 //x2=1.475 //y2=1.59
cc_1392 ( N_noxref_9_c_1913_n N_noxref_11_c_2423_n ) capacitor c=0.00698822f \
 //x=1.34 //y=1.22 //x2=1.475 //y2=1.59
cc_1393 ( N_noxref_9_c_1895_n N_noxref_11_c_2441_n ) capacitor c=0.0058169f \
 //x=11.355 //y=4.07 //x2=2.445 //y2=1.59
cc_1394 ( N_noxref_9_c_1895_n N_noxref_11_M0_noxref_s ) capacitor \
 c=0.00262629f //x=11.355 //y=4.07 //x2=0.455 //y2=0.375
cc_1395 ( N_noxref_9_c_1904_n N_noxref_11_M0_noxref_s ) capacitor c=0.0327271f \
 //x=0.81 //y=0.875 //x2=0.455 //y2=0.375
cc_1396 ( N_noxref_9_c_1907_n N_noxref_11_M0_noxref_s ) capacitor \
 c=7.99997e-19 //x=0.81 //y=1.53 //x2=0.455 //y2=0.375
cc_1397 ( N_noxref_9_c_1908_n N_noxref_11_M0_noxref_s ) capacitor \
 c=0.00122123f //x=0.81 //y=1.915 //x2=0.455 //y2=0.375
cc_1398 ( N_noxref_9_c_1911_n N_noxref_11_M0_noxref_s ) capacitor c=0.0121427f \
 //x=1.34 //y=0.875 //x2=0.455 //y2=0.375
cc_1399 ( N_noxref_9_c_1895_n N_noxref_12_c_2470_n ) capacitor c=0.0020922f \
 //x=11.355 //y=4.07 //x2=3.015 //y2=0.995
cc_1400 ( N_noxref_9_c_1895_n N_noxref_12_M2_noxref_s ) capacitor \
 c=0.00143334f //x=11.355 //y=4.07 //x2=2.965 //y2=0.375
cc_1401 ( N_noxref_9_c_1895_n N_D_c_2523_n ) capacitor c=0.0190126f //x=11.355 \
 //y=4.07 //x2=7.03 //y2=2.08
cc_1402 ( N_noxref_9_c_2014_n N_noxref_16_c_2714_n ) capacitor c=0.00623646f \
 //x=11.505 //y=1.56 //x2=11.285 //y2=1.495
cc_1403 ( N_noxref_9_c_2019_n N_noxref_16_c_2714_n ) capacitor c=0.00173579f \
 //x=11.47 //y=2.08 //x2=11.285 //y2=1.495
cc_1404 ( N_noxref_9_c_1899_n N_noxref_16_c_2715_n ) capacitor c=0.00156605f \
 //x=11.47 //y=2.08 //x2=12.17 //y2=0.53
cc_1405 ( N_noxref_9_c_2009_n N_noxref_16_c_2715_n ) capacitor c=0.0188655f \
 //x=11.505 //y=0.905 //x2=12.17 //y2=0.53
cc_1406 ( N_noxref_9_c_2017_n N_noxref_16_c_2715_n ) capacitor c=0.00656458f \
 //x=12.035 //y=0.905 //x2=12.17 //y2=0.53
cc_1407 ( N_noxref_9_c_2019_n N_noxref_16_c_2715_n ) capacitor c=2.1838e-19 \
 //x=11.47 //y=2.08 //x2=12.17 //y2=0.53
cc_1408 ( N_noxref_9_c_2009_n N_noxref_16_M6_noxref_s ) capacitor \
 c=0.00623646f //x=11.505 //y=0.905 //x2=10.18 //y2=0.365
cc_1409 ( N_noxref_9_c_2017_n N_noxref_16_M6_noxref_s ) capacitor c=0.0143002f \
 //x=12.035 //y=0.905 //x2=10.18 //y2=0.365
cc_1410 ( N_noxref_9_c_2018_n N_noxref_16_M6_noxref_s ) capacitor \
 c=0.00290153f //x=12.035 //y=1.25 //x2=10.18 //y2=0.365
cc_1411 ( N_noxref_9_M10_noxref_d N_noxref_17_M8_noxref_s ) capacitor \
 c=0.00309936f //x=16.345 //y=0.915 //x2=13.405 //y2=0.375
cc_1412 ( N_noxref_9_c_1901_n N_noxref_18_c_2814_n ) capacitor c=0.00457167f \
 //x=16.935 //y=1.665 //x2=16.935 //y2=0.54
cc_1413 ( N_noxref_9_M10_noxref_d N_noxref_18_c_2814_n ) capacitor \
 c=0.0115903f //x=16.345 //y=0.915 //x2=16.935 //y2=0.54
cc_1414 ( N_noxref_9_c_2144_n N_noxref_18_c_2842_n ) capacitor c=0.0200405f \
 //x=16.62 //y=1.665 //x2=16.05 //y2=0.995
cc_1415 ( N_noxref_9_M10_noxref_d N_noxref_18_M9_noxref_d ) capacitor \
 c=5.27807e-19 //x=16.345 //y=0.915 //x2=14.81 //y2=0.91
cc_1416 ( N_noxref_9_c_1901_n N_noxref_18_M10_noxref_s ) capacitor \
 c=0.0196084f //x=16.935 //y=1.665 //x2=15.915 //y2=0.375
cc_1417 ( N_noxref_9_M10_noxref_d N_noxref_18_M10_noxref_s ) capacitor \
 c=0.0426368f //x=16.345 //y=0.915 //x2=15.915 //y2=0.375
cc_1418 ( N_noxref_9_c_1901_n N_noxref_19_c_2879_n ) capacitor c=3.84569e-19 \
 //x=16.935 //y=1.665 //x2=18.35 //y2=1.505
cc_1419 ( N_noxref_9_c_1897_n N_noxref_19_c_2893_n ) capacitor c=9.18225e-19 \
 //x=24.305 //y=4.07 //x2=20.205 //y2=1.59
cc_1420 ( N_noxref_9_c_1897_n N_noxref_19_M11_noxref_s ) capacitor \
 c=0.00119468f //x=24.305 //y=4.07 //x2=18.215 //y2=0.375
cc_1421 ( N_noxref_9_M10_noxref_d N_noxref_19_M11_noxref_s ) capacitor \
 c=2.55333e-19 //x=16.345 //y=0.915 //x2=18.215 //y2=0.375
cc_1422 ( N_noxref_9_c_1897_n N_noxref_20_c_2915_n ) capacitor c=0.00161795f \
 //x=24.305 //y=4.07 //x2=20.775 //y2=0.995
cc_1423 ( N_noxref_9_c_1897_n N_noxref_20_M13_noxref_s ) capacitor \
 c=0.00122424f //x=24.305 //y=4.07 //x2=20.725 //y2=0.375
cc_1424 ( N_noxref_9_c_2189_n N_noxref_21_c_2974_n ) capacitor c=0.00623646f \
 //x=24.455 //y=1.56 //x2=24.235 //y2=1.495
cc_1425 ( N_noxref_9_c_2194_n N_noxref_21_c_2974_n ) capacitor c=0.00176439f \
 //x=24.42 //y=2.08 //x2=24.235 //y2=1.495
cc_1426 ( N_noxref_9_c_1902_n N_noxref_21_c_2975_n ) capacitor c=0.0016032f \
 //x=24.42 //y=2.08 //x2=25.12 //y2=0.53
cc_1427 ( N_noxref_9_c_2184_n N_noxref_21_c_2975_n ) capacitor c=0.0188655f \
 //x=24.455 //y=0.905 //x2=25.12 //y2=0.53
cc_1428 ( N_noxref_9_c_2192_n N_noxref_21_c_2975_n ) capacitor c=0.00656458f \
 //x=24.985 //y=0.905 //x2=25.12 //y2=0.53
cc_1429 ( N_noxref_9_c_2194_n N_noxref_21_c_2975_n ) capacitor c=2.1838e-19 \
 //x=24.42 //y=2.08 //x2=25.12 //y2=0.53
cc_1430 ( N_noxref_9_c_2184_n N_noxref_21_M14_noxref_s ) capacitor \
 c=0.00623646f //x=24.455 //y=0.905 //x2=23.13 //y2=0.365
cc_1431 ( N_noxref_9_c_2192_n N_noxref_21_M14_noxref_s ) capacitor \
 c=0.0143002f //x=24.985 //y=0.905 //x2=23.13 //y2=0.365
cc_1432 ( N_noxref_9_c_2193_n N_noxref_21_M14_noxref_s ) capacitor \
 c=0.00290153f //x=24.985 //y=1.25 //x2=23.13 //y2=0.365
cc_1433 ( N_noxref_10_c_2281_n N_noxref_20_c_2920_n ) capacitor c=0.00209081f \
 //x=21.09 //y=2.08 //x2=21.745 //y2=0.54
cc_1434 ( N_noxref_10_c_2325_n N_noxref_20_c_2920_n ) capacitor c=0.0194423f \
 //x=21.08 //y=0.915 //x2=21.745 //y2=0.54
cc_1435 ( N_noxref_10_c_2361_n N_noxref_20_c_2920_n ) capacitor c=0.00656458f \
 //x=21.61 //y=0.915 //x2=21.745 //y2=0.54
cc_1436 ( N_noxref_10_c_2328_n N_noxref_20_c_2920_n ) capacitor c=2.20712e-19 \
 //x=21.09 //y=2.08 //x2=21.745 //y2=0.54
cc_1437 ( N_noxref_10_c_2326_n N_noxref_20_c_2943_n ) capacitor c=0.00538829f \
 //x=21.08 //y=1.26 //x2=20.86 //y2=0.995
cc_1438 ( N_noxref_10_c_2325_n N_noxref_20_M13_noxref_s ) capacitor \
 c=0.00538829f //x=21.08 //y=0.915 //x2=20.725 //y2=0.375
cc_1439 ( N_noxref_10_c_2327_n N_noxref_20_M13_noxref_s ) capacitor \
 c=0.00538829f //x=21.08 //y=1.57 //x2=20.725 //y2=0.375
cc_1440 ( N_noxref_10_c_2361_n N_noxref_20_M13_noxref_s ) capacitor \
 c=0.0143002f //x=21.61 //y=0.915 //x2=20.725 //y2=0.375
cc_1441 ( N_noxref_10_c_2362_n N_noxref_20_M13_noxref_s ) capacitor \
 c=0.00290153f //x=21.61 //y=1.26 //x2=20.725 //y2=0.375
cc_1442 ( N_noxref_10_c_2413_p N_noxref_21_c_2984_n ) capacitor c=3.15806e-19 \
 //x=24.805 //y=1.655 //x2=23.265 //y2=1.495
cc_1443 ( N_noxref_10_c_2279_n N_noxref_21_c_2967_n ) capacitor c=0.00299723f \
 //x=25.045 //y=3.7 //x2=24.15 //y2=1.58
cc_1444 ( N_noxref_10_c_2279_n N_noxref_21_c_2974_n ) capacitor c=0.00187232f \
 //x=25.045 //y=3.7 //x2=24.235 //y2=1.495
cc_1445 ( N_noxref_10_c_2413_p N_noxref_21_c_2974_n ) capacitor c=0.020324f \
 //x=24.805 //y=1.655 //x2=24.235 //y2=1.495
cc_1446 ( N_noxref_10_c_2279_n N_noxref_21_c_2975_n ) capacitor c=4.7198e-19 \
 //x=25.045 //y=3.7 //x2=25.12 //y2=0.53
cc_1447 ( N_noxref_10_c_2282_n N_noxref_21_c_2975_n ) capacitor c=0.00467104f \
 //x=25.075 //y=1.655 //x2=25.12 //y2=0.53
cc_1448 ( N_noxref_10_M15_noxref_d N_noxref_21_c_2975_n ) capacitor \
 c=0.0117932f //x=24.53 //y=0.905 //x2=25.12 //y2=0.53
cc_1449 ( N_noxref_10_c_2279_n N_noxref_21_M14_noxref_s ) capacitor \
 c=3.61944e-19 //x=25.045 //y=3.7 //x2=23.13 //y2=0.365
cc_1450 ( N_noxref_10_c_2282_n N_noxref_21_M14_noxref_s ) capacitor \
 c=0.0142774f //x=25.075 //y=1.655 //x2=23.13 //y2=0.365
cc_1451 ( N_noxref_10_M15_noxref_d N_noxref_21_M14_noxref_s ) capacitor \
 c=0.0439476f //x=24.53 //y=0.905 //x2=23.13 //y2=0.365
cc_1452 ( N_noxref_11_c_2430_n N_noxref_12_c_2470_n ) capacitor c=0.0136048f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_1453 ( N_noxref_11_c_2441_n N_noxref_12_c_2470_n ) capacitor c=0.0102225f \
 //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_1454 ( N_noxref_11_M0_noxref_s N_noxref_12_c_2470_n ) capacitor \
 c=0.0228676f //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_1455 ( N_noxref_11_M0_noxref_s N_noxref_12_c_2472_n ) capacitor \
 c=0.0180035f //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_1456 ( N_noxref_11_c_2430_n N_noxref_12_M1_noxref_d ) capacitor \
 c=0.0129526f //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_1457 ( N_noxref_11_c_2441_n N_noxref_12_M1_noxref_d ) capacitor \
 c=0.00908243f //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_1458 ( N_noxref_11_M0_noxref_s N_noxref_12_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_1459 ( N_noxref_11_M0_noxref_s N_noxref_12_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_1460 ( N_noxref_12_c_2478_n N_noxref_14_M3_noxref_s ) capacitor \
 c=0.00191848f //x=4.07 //y=0.625 //x2=5.265 //y2=0.375
cc_1461 ( N_D_c_2552_n N_noxref_14_c_2610_n ) capacitor c=0.0167228f //x=6.595 \
 //y=0.91 //x2=7.255 //y2=0.54
cc_1462 ( N_D_c_2557_n N_noxref_14_c_2610_n ) capacitor c=0.00534519f //x=7.12 \
 //y=0.91 //x2=7.255 //y2=0.54
cc_1463 ( N_D_c_2523_n N_noxref_14_c_2621_n ) capacitor c=0.0125737f //x=7.03 \
 //y=2.08 //x2=7.255 //y2=1.59
cc_1464 ( N_D_c_2555_n N_noxref_14_c_2621_n ) capacitor c=0.0153476f //x=6.595 \
 //y=1.22 //x2=7.255 //y2=1.59
cc_1465 ( N_D_c_2560_n N_noxref_14_c_2621_n ) capacitor c=0.0226946f //x=7.12 \
 //y=1.915 //x2=7.255 //y2=1.59
cc_1466 ( N_D_c_2552_n N_noxref_14_M3_noxref_s ) capacitor c=0.00798959f \
 //x=6.595 //y=0.91 //x2=5.265 //y2=0.375
cc_1467 ( N_D_c_2559_n N_noxref_14_M3_noxref_s ) capacitor c=0.00212176f \
 //x=7.12 //y=1.45 //x2=5.265 //y2=0.375
cc_1468 ( N_D_c_2560_n N_noxref_14_M3_noxref_s ) capacitor c=0.00298115f \
 //x=7.12 //y=1.915 //x2=5.265 //y2=0.375
cc_1469 ( N_D_c_2591_p N_noxref_15_c_2653_n ) capacitor c=2.14837e-19 \
 //x=6.965 //y=0.755 //x2=7.825 //y2=0.995
cc_1470 ( N_D_c_2557_n N_noxref_15_c_2653_n ) capacitor c=0.00123426f //x=7.12 \
 //y=0.91 //x2=7.825 //y2=0.995
cc_1471 ( N_D_c_2558_n N_noxref_15_c_2653_n ) capacitor c=0.0129288f //x=7.12 \
 //y=1.22 //x2=7.825 //y2=0.995
cc_1472 ( N_D_c_2559_n N_noxref_15_c_2653_n ) capacitor c=0.00142359f //x=7.12 \
 //y=1.45 //x2=7.825 //y2=0.995
cc_1473 ( N_D_c_2552_n N_noxref_15_M4_noxref_d ) capacitor c=0.00223875f \
 //x=6.595 //y=0.91 //x2=6.67 //y2=0.91
cc_1474 ( N_D_c_2555_n N_noxref_15_M4_noxref_d ) capacitor c=0.00262485f \
 //x=6.595 //y=1.22 //x2=6.67 //y2=0.91
cc_1475 ( N_D_c_2591_p N_noxref_15_M4_noxref_d ) capacitor c=0.00220746f \
 //x=6.965 //y=0.755 //x2=6.67 //y2=0.91
cc_1476 ( N_D_c_2598_p N_noxref_15_M4_noxref_d ) capacitor c=0.00194798f \
 //x=6.965 //y=1.375 //x2=6.67 //y2=0.91
cc_1477 ( N_D_c_2557_n N_noxref_15_M4_noxref_d ) capacitor c=0.00198465f \
 //x=7.12 //y=0.91 //x2=6.67 //y2=0.91
cc_1478 ( N_D_c_2558_n N_noxref_15_M4_noxref_d ) capacitor c=0.00128384f \
 //x=7.12 //y=1.22 //x2=6.67 //y2=0.91
cc_1479 ( N_D_c_2557_n N_noxref_15_M5_noxref_s ) capacitor c=7.21316e-19 \
 //x=7.12 //y=0.91 //x2=7.775 //y2=0.375
cc_1480 ( N_D_c_2558_n N_noxref_15_M5_noxref_s ) capacitor c=0.00348171f \
 //x=7.12 //y=1.22 //x2=7.775 //y2=0.375
cc_1481 ( N_noxref_14_c_2610_n N_noxref_15_c_2653_n ) capacitor c=0.0134311f \
 //x=7.255 //y=0.54 //x2=7.825 //y2=0.995
cc_1482 ( N_noxref_14_c_2621_n N_noxref_15_c_2653_n ) capacitor c=0.0101712f \
 //x=7.255 //y=1.59 //x2=7.825 //y2=0.995
cc_1483 ( N_noxref_14_M3_noxref_s N_noxref_15_c_2653_n ) capacitor \
 c=0.0227445f //x=5.265 //y=0.375 //x2=7.825 //y2=0.995
cc_1484 ( N_noxref_14_M3_noxref_s N_noxref_15_c_2655_n ) capacitor \
 c=0.0180035f //x=5.265 //y=0.375 //x2=7.91 //y2=0.625
cc_1485 ( N_noxref_14_c_2610_n N_noxref_15_M4_noxref_d ) capacitor \
 c=0.0128913f //x=7.255 //y=0.54 //x2=6.67 //y2=0.91
cc_1486 ( N_noxref_14_c_2621_n N_noxref_15_M4_noxref_d ) capacitor \
 c=0.00899889f //x=7.255 //y=1.59 //x2=6.67 //y2=0.91
cc_1487 ( N_noxref_14_M3_noxref_s N_noxref_15_M4_noxref_d ) capacitor \
 c=0.0159202f //x=5.265 //y=0.375 //x2=6.67 //y2=0.91
cc_1488 ( N_noxref_14_M3_noxref_s N_noxref_15_M5_noxref_s ) capacitor \
 c=0.0213553f //x=5.265 //y=0.375 //x2=7.775 //y2=0.375
cc_1489 ( N_noxref_15_c_2661_n N_noxref_16_M6_noxref_s ) capacitor \
 c=0.00164795f //x=8.88 //y=0.625 //x2=10.18 //y2=0.365
cc_1490 ( N_noxref_16_c_2718_n N_noxref_17_M8_noxref_s ) capacitor \
 c=0.00199452f //x=12.255 //y=0.615 //x2=13.405 //y2=0.375
cc_1491 ( N_noxref_17_c_2766_n N_noxref_18_c_2809_n ) capacitor c=0.0131877f \
 //x=15.395 //y=0.54 //x2=15.965 //y2=0.995
cc_1492 ( N_noxref_17_c_2789_n N_noxref_18_c_2809_n ) capacitor c=0.00981707f \
 //x=15.395 //y=1.59 //x2=15.965 //y2=0.995
cc_1493 ( N_noxref_17_M8_noxref_s N_noxref_18_c_2809_n ) capacitor \
 c=0.0221661f //x=13.405 //y=0.375 //x2=15.965 //y2=0.995
cc_1494 ( N_noxref_17_M8_noxref_s N_noxref_18_c_2811_n ) capacitor \
 c=0.0180035f //x=13.405 //y=0.375 //x2=16.05 //y2=0.625
cc_1495 ( N_noxref_17_c_2766_n N_noxref_18_M9_noxref_d ) capacitor \
 c=0.0127191f //x=15.395 //y=0.54 //x2=14.81 //y2=0.91
cc_1496 ( N_noxref_17_c_2789_n N_noxref_18_M9_noxref_d ) capacitor \
 c=0.00861161f //x=15.395 //y=1.59 //x2=14.81 //y2=0.91
cc_1497 ( N_noxref_17_M8_noxref_s N_noxref_18_M9_noxref_d ) capacitor \
 c=0.0159202f //x=13.405 //y=0.375 //x2=14.81 //y2=0.91
cc_1498 ( N_noxref_17_M8_noxref_s N_noxref_18_M10_noxref_s ) capacitor \
 c=0.0213553f //x=13.405 //y=0.375 //x2=15.915 //y2=0.375
cc_1499 ( N_noxref_18_c_2817_n N_noxref_19_M11_noxref_s ) capacitor \
 c=0.00191848f //x=17.02 //y=0.625 //x2=18.215 //y2=0.375
cc_1500 ( N_noxref_19_c_2870_n N_noxref_20_c_2915_n ) capacitor c=0.0133566f \
 //x=20.205 //y=0.54 //x2=20.775 //y2=0.995
cc_1501 ( N_noxref_19_c_2893_n N_noxref_20_c_2915_n ) capacitor c=0.00992008f \
 //x=20.205 //y=1.59 //x2=20.775 //y2=0.995
cc_1502 ( N_noxref_19_M11_noxref_s N_noxref_20_c_2915_n ) capacitor \
 c=0.0228676f //x=18.215 //y=0.375 //x2=20.775 //y2=0.995
cc_1503 ( N_noxref_19_M11_noxref_s N_noxref_20_c_2917_n ) capacitor \
 c=0.0180035f //x=18.215 //y=0.375 //x2=20.86 //y2=0.625
cc_1504 ( N_noxref_19_c_2870_n N_noxref_20_M12_noxref_d ) capacitor \
 c=0.0127176f //x=20.205 //y=0.54 //x2=19.62 //y2=0.91
cc_1505 ( N_noxref_19_c_2893_n N_noxref_20_M12_noxref_d ) capacitor \
 c=0.0086073f //x=20.205 //y=1.59 //x2=19.62 //y2=0.91
cc_1506 ( N_noxref_19_M11_noxref_s N_noxref_20_M12_noxref_d ) capacitor \
 c=0.0159202f //x=18.215 //y=0.375 //x2=19.62 //y2=0.91
cc_1507 ( N_noxref_19_M11_noxref_s N_noxref_20_M13_noxref_s ) capacitor \
 c=0.0213553f //x=18.215 //y=0.375 //x2=20.725 //y2=0.375
cc_1508 ( N_noxref_20_c_2923_n N_noxref_21_M14_noxref_s ) capacitor \
 c=0.00164795f //x=21.83 //y=0.625 //x2=23.13 //y2=0.365
