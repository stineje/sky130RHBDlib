* SPICE3 file created from DLATCHN.ext - technology: sky130A

.subckt DLATCHN Q D GATE_N VPB VNB
M1000 VPB.t19 a_1105_1004.t5 a_1739_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 Q a_3451_383.t6 VNB.t7 nshort w=-1.83u l=2.06u
+  ad=0.3582p pd=3.15u as=0p ps=0u
M1002 VPB.t12 a_185_182.t3 a_2215_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_3905_1005.t2 Q VPB.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1105_1004.t1 a_629_182.t3 VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t4 a_1739_182.t3 a_3239_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_3905_1005.t0 a_2849_182.t3 a_3451_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_1105_1004.t4 a_185_182.t4 VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t14 D a_629_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VNB a_629_182.t4 a_1000_73.t0 nshort w=-1.605u l=1.765u
+  ad=8.7946p pd=61.42u as=0p ps=0u
M1010 Q a_3451_383.t4 a_3239_1005.t0 pshort w=2u l=0.15u
+  ad=0.58p pd=4.58u as=0p ps=0u
M1011 VPB.t8 a_2215_1004.t5 a_2849_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t9 Q a_3905_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_629_182.t1 D VPB.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1739_182.t0 a_1105_1004.t7 VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPB.t0 a_121_384# a_185_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VNB a_185_182.t5 a_2110_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_2215_1004.t0 a_185_182.t6 VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPB.t7 a_185_182.t8 a_1105_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_2215_1004.t4 D VPB.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_3451_383.t0 a_2849_182.t4 a_3905_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_3239_1005.t3 a_3451_383.t5 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t2 a_629_182.t5 a_1105_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_1739_182.t4 VNB.t1 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_3239_1005.t1 a_1739_182.t5 VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2849_182.t1 a_2215_1004.t7 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_185_182.t1 a_121_384# VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPB.t13 D a_2215_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB Q 0.34fF
C1 D a_121_384# 0.01fF
C2 VPB a_121_384# 0.12fF
C3 VPB D 0.62fF
R0 a_1105_1004.n4 a_1105_1004.t5 512.525
R1 a_1105_1004.n4 a_1105_1004.t7 371.139
R2 a_1105_1004.n5 a_1105_1004.t6 220.263
R3 a_1105_1004.n8 a_1105_1004.n6 194.086
R4 a_1105_1004.n6 a_1105_1004.n3 162.547
R5 a_1105_1004.n5 a_1105_1004.n4 158.3
R6 a_1105_1004.n6 a_1105_1004.n5 153.043
R7 a_1105_1004.n3 a_1105_1004.n2 76.002
R8 a_1105_1004.n9 a_1105_1004.n0 55.263
R9 a_1105_1004.n8 a_1105_1004.n7 30
R10 a_1105_1004.n9 a_1105_1004.n8 23.684
R11 a_1105_1004.n1 a_1105_1004.t2 14.282
R12 a_1105_1004.n1 a_1105_1004.t4 14.282
R13 a_1105_1004.n2 a_1105_1004.t0 14.282
R14 a_1105_1004.n2 a_1105_1004.t1 14.282
R15 a_1105_1004.n3 a_1105_1004.n1 12.85
R16 a_1739_182.n2 a_1739_182.t5 486.819
R17 a_1739_182.n2 a_1739_182.t3 384.527
R18 a_1739_182.n3 a_1739_182.t4 287.101
R19 a_1739_182.n6 a_1739_182.n4 215.257
R20 a_1739_182.n4 a_1739_182.n3 157.396
R21 a_1739_182.n4 a_1739_182.n1 140.59
R22 a_1739_182.n3 a_1739_182.n2 90.041
R23 a_1739_182.n6 a_1739_182.n5 30
R24 a_1739_182.n7 a_1739_182.n0 24.383
R25 a_1739_182.n7 a_1739_182.n6 23.684
R26 a_1739_182.n1 a_1739_182.t2 14.282
R27 a_1739_182.n1 a_1739_182.t0 14.282
R28 VPB VPB.n447 126.832
R29 VPB.n80 VPB.n78 94.117
R30 VPB.n59 VPB.n57 94.117
R31 VPB.n391 VPB.n389 94.117
R32 VPB.n344 VPB.n342 94.117
R33 VPB.n163 VPB.n161 94.117
R34 VPB.n142 VPB.n140 94.117
R35 VPB.n258 VPB.n256 94.117
R36 VPB.n218 VPB.n217 76
R37 VPB.n225 VPB.n224 76
R38 VPB.n229 VPB.n228 76
R39 VPB.n233 VPB.n232 76
R40 VPB.n260 VPB.n259 76
R41 VPB.n264 VPB.n263 76
R42 VPB.n268 VPB.n267 76
R43 VPB.n272 VPB.n271 76
R44 VPB.n277 VPB.n276 76
R45 VPB.n284 VPB.n283 76
R46 VPB.n288 VPB.n287 76
R47 VPB.n292 VPB.n291 76
R48 VPB.n306 VPB.n302 76
R49 VPB.n310 VPB.n95 76
R50 VPB.n315 VPB.n314 76
R51 VPB.n319 VPB.n318 76
R52 VPB.n346 VPB.n345 76
R53 VPB.n352 VPB.n351 76
R54 VPB.n356 VPB.n355 76
R55 VPB.n362 VPB.n361 76
R56 VPB.n366 VPB.n365 76
R57 VPB.n393 VPB.n392 76
R58 VPB.n398 VPB.n397 76
R59 VPB.n403 VPB.n402 76
R60 VPB.n410 VPB.n409 76
R61 VPB.n415 VPB.n414 76
R62 VPB.n420 VPB.n419 76
R63 VPB.n425 VPB.n424 76
R64 VPB.n429 VPB.n428 76
R65 VPB.n440 VPB.n439 76
R66 VPB.n153 VPB.n152 68.979
R67 VPB.n359 VPB.n358 68.979
R68 VPB.n70 VPB.n69 68.979
R69 VPB.n91 VPB.n90 68.979
R70 VPB.n146 VPB.n145 64.528
R71 VPB.n349 VPB.n348 64.528
R72 VPB.n63 VPB.n62 64.528
R73 VPB.n84 VPB.n83 64.528
R74 VPB.n20 VPB.n19 61.764
R75 VPB.n41 VPB.n40 61.764
R76 VPB.n373 VPB.n372 61.764
R77 VPB.n326 VPB.n325 61.764
R78 VPB.n103 VPB.n102 61.764
R79 VPB.n124 VPB.n123 61.764
R80 VPB.n240 VPB.n239 61.764
R81 VPB.n94 VPB.t1 55.106
R82 VPB.n82 VPB.t0 55.106
R83 VPB.n73 VPB.t15 55.106
R84 VPB.n61 VPB.t14 55.106
R85 VPB.n421 VPB.t3 55.106
R86 VPB.n357 VPB.t18 55.106
R87 VPB.n347 VPB.t19 55.106
R88 VPB.n311 VPB.t17 55.106
R89 VPB.n156 VPB.t6 55.106
R90 VPB.n144 VPB.t8 55.106
R91 VPB.n394 VPB.t7 55.106
R92 VPB.n168 VPB.t13 55.106
R93 VPB.n170 VPB.n169 48.952
R94 VPB.n400 VPB.n399 48.952
R95 VPB.n222 VPB.n221 44.502
R96 VPB.n281 VPB.n280 44.502
R97 VPB.n308 VPB.n307 44.502
R98 VPB.n417 VPB.n416 44.502
R99 VPB.n279 VPB.n278 41.183
R100 VPB.n220 VPB.n219 41.183
R101 VPB.n405 VPB.n404 40.824
R102 VPB.n177 VPB.n96 40.824
R103 VPB.n212 VPB.n211 35.118
R104 VPB.n444 VPB.n440 20.452
R105 VPB.n201 VPB.n198 20.452
R106 VPB.n174 VPB.n173 17.801
R107 VPB.n407 VPB.n406 17.801
R108 VPB.n404 VPB.t11 14.282
R109 VPB.n404 VPB.t2 14.282
R110 VPB.n96 VPB.t16 14.282
R111 VPB.n96 VPB.t12 14.282
R112 VPB.n278 VPB.t5 14.282
R113 VPB.n278 VPB.t4 14.282
R114 VPB.n219 VPB.t10 14.282
R115 VPB.n219 VPB.t9 14.282
R116 VPB.n201 VPB.n200 13.653
R117 VPB.n200 VPB.n199 13.653
R118 VPB.n210 VPB.n209 13.653
R119 VPB.n209 VPB.n208 13.653
R120 VPB.n207 VPB.n206 13.653
R121 VPB.n206 VPB.n205 13.653
R122 VPB.n204 VPB.n203 13.653
R123 VPB.n203 VPB.n202 13.653
R124 VPB.n217 VPB.n216 13.653
R125 VPB.n216 VPB.n215 13.653
R126 VPB.n224 VPB.n223 13.653
R127 VPB.n223 VPB.n222 13.653
R128 VPB.n228 VPB.n227 13.653
R129 VPB.n227 VPB.n226 13.653
R130 VPB.n232 VPB.n231 13.653
R131 VPB.n231 VPB.n230 13.653
R132 VPB.n259 VPB.n258 13.653
R133 VPB.n258 VPB.n257 13.653
R134 VPB.n263 VPB.n262 13.653
R135 VPB.n262 VPB.n261 13.653
R136 VPB.n267 VPB.n266 13.653
R137 VPB.n266 VPB.n265 13.653
R138 VPB.n271 VPB.n270 13.653
R139 VPB.n270 VPB.n269 13.653
R140 VPB.n276 VPB.n275 13.653
R141 VPB.n275 VPB.n274 13.653
R142 VPB.n283 VPB.n282 13.653
R143 VPB.n282 VPB.n281 13.653
R144 VPB.n287 VPB.n286 13.653
R145 VPB.n286 VPB.n285 13.653
R146 VPB.n291 VPB.n290 13.653
R147 VPB.n290 VPB.n289 13.653
R148 VPB.n143 VPB.n142 13.653
R149 VPB.n142 VPB.n141 13.653
R150 VPB.n148 VPB.n147 13.653
R151 VPB.n147 VPB.n146 13.653
R152 VPB.n151 VPB.n150 13.653
R153 VPB.n150 VPB.n149 13.653
R154 VPB.n155 VPB.n154 13.653
R155 VPB.n154 VPB.n153 13.653
R156 VPB.n159 VPB.n158 13.653
R157 VPB.n158 VPB.n157 13.653
R158 VPB.n164 VPB.n163 13.653
R159 VPB.n163 VPB.n162 13.653
R160 VPB.n167 VPB.n166 13.653
R161 VPB.n166 VPB.n165 13.653
R162 VPB.n172 VPB.n171 13.653
R163 VPB.n171 VPB.n170 13.653
R164 VPB.n176 VPB.n175 13.653
R165 VPB.n175 VPB.n174 13.653
R166 VPB.n306 VPB.n305 13.653
R167 VPB.n305 VPB.n304 13.653
R168 VPB.n310 VPB.n309 13.653
R169 VPB.n309 VPB.n308 13.653
R170 VPB.n314 VPB.n313 13.653
R171 VPB.n313 VPB.n312 13.653
R172 VPB.n318 VPB.n317 13.653
R173 VPB.n317 VPB.n316 13.653
R174 VPB.n345 VPB.n344 13.653
R175 VPB.n344 VPB.n343 13.653
R176 VPB.n351 VPB.n350 13.653
R177 VPB.n350 VPB.n349 13.653
R178 VPB.n355 VPB.n354 13.653
R179 VPB.n354 VPB.n353 13.653
R180 VPB.n361 VPB.n360 13.653
R181 VPB.n360 VPB.n359 13.653
R182 VPB.n365 VPB.n364 13.653
R183 VPB.n364 VPB.n363 13.653
R184 VPB.n392 VPB.n391 13.653
R185 VPB.n391 VPB.n390 13.653
R186 VPB.n397 VPB.n396 13.653
R187 VPB.n396 VPB.n395 13.653
R188 VPB.n402 VPB.n401 13.653
R189 VPB.n401 VPB.n400 13.653
R190 VPB.n409 VPB.n408 13.653
R191 VPB.n408 VPB.n407 13.653
R192 VPB.n414 VPB.n413 13.653
R193 VPB.n413 VPB.n412 13.653
R194 VPB.n419 VPB.n418 13.653
R195 VPB.n418 VPB.n417 13.653
R196 VPB.n424 VPB.n423 13.653
R197 VPB.n423 VPB.n422 13.653
R198 VPB.n428 VPB.n427 13.653
R199 VPB.n427 VPB.n426 13.653
R200 VPB.n60 VPB.n59 13.653
R201 VPB.n59 VPB.n58 13.653
R202 VPB.n65 VPB.n64 13.653
R203 VPB.n64 VPB.n63 13.653
R204 VPB.n68 VPB.n67 13.653
R205 VPB.n67 VPB.n66 13.653
R206 VPB.n72 VPB.n71 13.653
R207 VPB.n71 VPB.n70 13.653
R208 VPB.n76 VPB.n75 13.653
R209 VPB.n75 VPB.n74 13.653
R210 VPB.n81 VPB.n80 13.653
R211 VPB.n80 VPB.n79 13.653
R212 VPB.n86 VPB.n85 13.653
R213 VPB.n85 VPB.n84 13.653
R214 VPB.n89 VPB.n88 13.653
R215 VPB.n88 VPB.n87 13.653
R216 VPB.n93 VPB.n92 13.653
R217 VPB.n92 VPB.n91 13.653
R218 VPB.n440 VPB.n0 13.653
R219 VPB VPB.n0 13.653
R220 VPB.n215 VPB.n214 13.35
R221 VPB.n274 VPB.n273 13.35
R222 VPB.n304 VPB.n303 13.35
R223 VPB.n412 VPB.n411 13.35
R224 VPB.n444 VPB.n443 13.276
R225 VPB.n443 VPB.n441 13.276
R226 VPB.n34 VPB.n16 13.276
R227 VPB.n16 VPB.n14 13.276
R228 VPB.n55 VPB.n37 13.276
R229 VPB.n37 VPB.n35 13.276
R230 VPB.n387 VPB.n369 13.276
R231 VPB.n369 VPB.n367 13.276
R232 VPB.n340 VPB.n322 13.276
R233 VPB.n322 VPB.n320 13.276
R234 VPB.n117 VPB.n99 13.276
R235 VPB.n99 VPB.n97 13.276
R236 VPB.n138 VPB.n120 13.276
R237 VPB.n120 VPB.n118 13.276
R238 VPB.n254 VPB.n236 13.276
R239 VPB.n236 VPB.n234 13.276
R240 VPB.n210 VPB.n207 13.276
R241 VPB.n207 VPB.n204 13.276
R242 VPB.n259 VPB.n255 13.276
R243 VPB.n143 VPB.n139 13.276
R244 VPB.n151 VPB.n148 13.276
R245 VPB.n155 VPB.n151 13.276
R246 VPB.n160 VPB.n159 13.276
R247 VPB.n164 VPB.n160 13.276
R248 VPB.n167 VPB.n164 13.276
R249 VPB.n176 VPB.n172 13.276
R250 VPB.n310 VPB.n306 13.276
R251 VPB.n345 VPB.n341 13.276
R252 VPB.n392 VPB.n388 13.276
R253 VPB.n60 VPB.n56 13.276
R254 VPB.n68 VPB.n65 13.276
R255 VPB.n72 VPB.n68 13.276
R256 VPB.n77 VPB.n76 13.276
R257 VPB.n81 VPB.n77 13.276
R258 VPB.n89 VPB.n86 13.276
R259 VPB.n93 VPB.n89 13.276
R260 VPB.n198 VPB.n180 13.276
R261 VPB.n180 VPB.n178 13.276
R262 VPB.n185 VPB.n183 12.796
R263 VPB.n185 VPB.n184 12.564
R264 VPB.n194 VPB.n193 12.198
R265 VPB.n192 VPB.n191 12.198
R266 VPB.n188 VPB.n187 12.198
R267 VPB.n172 VPB.n168 11.841
R268 VPB.n311 VPB.n310 11.482
R269 VPB.n159 VPB.n156 10.944
R270 VPB.n76 VPB.n73 10.944
R271 VPB.n440 VPB.n94 10.944
R272 VPB.n144 VPB.n143 10.585
R273 VPB.n61 VPB.n60 10.585
R274 VPB.n82 VPB.n81 10.585
R275 VPB.n198 VPB.n197 7.5
R276 VPB.n183 VPB.n182 7.5
R277 VPB.n187 VPB.n186 7.5
R278 VPB.n191 VPB.n190 7.5
R279 VPB.n180 VPB.n179 7.5
R280 VPB.n195 VPB.n181 7.5
R281 VPB.n236 VPB.n235 7.5
R282 VPB.n249 VPB.n248 7.5
R283 VPB.n243 VPB.n242 7.5
R284 VPB.n245 VPB.n244 7.5
R285 VPB.n238 VPB.n237 7.5
R286 VPB.n254 VPB.n253 7.5
R287 VPB.n120 VPB.n119 7.5
R288 VPB.n133 VPB.n132 7.5
R289 VPB.n127 VPB.n126 7.5
R290 VPB.n129 VPB.n128 7.5
R291 VPB.n122 VPB.n121 7.5
R292 VPB.n138 VPB.n137 7.5
R293 VPB.n99 VPB.n98 7.5
R294 VPB.n112 VPB.n111 7.5
R295 VPB.n106 VPB.n105 7.5
R296 VPB.n108 VPB.n107 7.5
R297 VPB.n101 VPB.n100 7.5
R298 VPB.n117 VPB.n116 7.5
R299 VPB.n322 VPB.n321 7.5
R300 VPB.n335 VPB.n334 7.5
R301 VPB.n329 VPB.n328 7.5
R302 VPB.n331 VPB.n330 7.5
R303 VPB.n324 VPB.n323 7.5
R304 VPB.n340 VPB.n339 7.5
R305 VPB.n369 VPB.n368 7.5
R306 VPB.n382 VPB.n381 7.5
R307 VPB.n376 VPB.n375 7.5
R308 VPB.n378 VPB.n377 7.5
R309 VPB.n371 VPB.n370 7.5
R310 VPB.n387 VPB.n386 7.5
R311 VPB.n37 VPB.n36 7.5
R312 VPB.n50 VPB.n49 7.5
R313 VPB.n44 VPB.n43 7.5
R314 VPB.n46 VPB.n45 7.5
R315 VPB.n39 VPB.n38 7.5
R316 VPB.n55 VPB.n54 7.5
R317 VPB.n16 VPB.n15 7.5
R318 VPB.n29 VPB.n28 7.5
R319 VPB.n23 VPB.n22 7.5
R320 VPB.n25 VPB.n24 7.5
R321 VPB.n18 VPB.n17 7.5
R322 VPB.n34 VPB.n33 7.5
R323 VPB.n443 VPB.n442 7.5
R324 VPB.n12 VPB.n11 7.5
R325 VPB.n6 VPB.n5 7.5
R326 VPB.n8 VPB.n7 7.5
R327 VPB.n2 VPB.n1 7.5
R328 VPB.n445 VPB.n444 7.5
R329 VPB.n77 VPB.n34 7.176
R330 VPB.n56 VPB.n55 7.176
R331 VPB.n388 VPB.n387 7.176
R332 VPB.n341 VPB.n340 7.176
R333 VPB.n160 VPB.n117 7.176
R334 VPB.n139 VPB.n138 7.176
R335 VPB.n255 VPB.n254 7.176
R336 VPB.n306 VPB.n177 6.817
R337 VPB.n250 VPB.n247 6.729
R338 VPB.n246 VPB.n243 6.729
R339 VPB.n241 VPB.n238 6.729
R340 VPB.n134 VPB.n131 6.729
R341 VPB.n130 VPB.n127 6.729
R342 VPB.n125 VPB.n122 6.729
R343 VPB.n113 VPB.n110 6.729
R344 VPB.n109 VPB.n106 6.729
R345 VPB.n104 VPB.n101 6.729
R346 VPB.n336 VPB.n333 6.729
R347 VPB.n332 VPB.n329 6.729
R348 VPB.n327 VPB.n324 6.729
R349 VPB.n383 VPB.n380 6.729
R350 VPB.n379 VPB.n376 6.729
R351 VPB.n374 VPB.n371 6.729
R352 VPB.n51 VPB.n48 6.729
R353 VPB.n47 VPB.n44 6.729
R354 VPB.n42 VPB.n39 6.729
R355 VPB.n30 VPB.n27 6.729
R356 VPB.n26 VPB.n23 6.729
R357 VPB.n21 VPB.n18 6.729
R358 VPB.n13 VPB.n10 6.729
R359 VPB.n9 VPB.n6 6.729
R360 VPB.n4 VPB.n2 6.729
R361 VPB.n241 VPB.n240 6.728
R362 VPB.n246 VPB.n245 6.728
R363 VPB.n250 VPB.n249 6.728
R364 VPB.n253 VPB.n252 6.728
R365 VPB.n125 VPB.n124 6.728
R366 VPB.n130 VPB.n129 6.728
R367 VPB.n134 VPB.n133 6.728
R368 VPB.n137 VPB.n136 6.728
R369 VPB.n104 VPB.n103 6.728
R370 VPB.n109 VPB.n108 6.728
R371 VPB.n113 VPB.n112 6.728
R372 VPB.n116 VPB.n115 6.728
R373 VPB.n327 VPB.n326 6.728
R374 VPB.n332 VPB.n331 6.728
R375 VPB.n336 VPB.n335 6.728
R376 VPB.n339 VPB.n338 6.728
R377 VPB.n374 VPB.n373 6.728
R378 VPB.n379 VPB.n378 6.728
R379 VPB.n383 VPB.n382 6.728
R380 VPB.n386 VPB.n385 6.728
R381 VPB.n42 VPB.n41 6.728
R382 VPB.n47 VPB.n46 6.728
R383 VPB.n51 VPB.n50 6.728
R384 VPB.n54 VPB.n53 6.728
R385 VPB.n21 VPB.n20 6.728
R386 VPB.n26 VPB.n25 6.728
R387 VPB.n30 VPB.n29 6.728
R388 VPB.n33 VPB.n32 6.728
R389 VPB.n4 VPB.n3 6.728
R390 VPB.n9 VPB.n8 6.728
R391 VPB.n13 VPB.n12 6.728
R392 VPB.n446 VPB.n445 6.728
R393 VPB.n177 VPB.n176 6.458
R394 VPB.n409 VPB.n405 6.458
R395 VPB.n197 VPB.n196 6.398
R396 VPB.n211 VPB.n201 6.112
R397 VPB.n211 VPB.n210 6.101
R398 VPB.n224 VPB.n220 4.305
R399 VPB.n283 VPB.n279 4.305
R400 VPB.n148 VPB.n144 2.691
R401 VPB.n351 VPB.n347 2.691
R402 VPB.n65 VPB.n61 2.691
R403 VPB.n86 VPB.n82 2.691
R404 VPB.n156 VPB.n155 2.332
R405 VPB.n361 VPB.n357 2.332
R406 VPB.n73 VPB.n72 2.332
R407 VPB.n94 VPB.n93 2.332
R408 VPB.n314 VPB.n311 1.794
R409 VPB.n424 VPB.n421 1.794
R410 VPB.n168 VPB.n167 1.435
R411 VPB.n397 VPB.n394 1.435
R412 VPB.n195 VPB.n188 1.402
R413 VPB.n195 VPB.n189 1.402
R414 VPB.n195 VPB.n192 1.402
R415 VPB.n195 VPB.n194 1.402
R416 VPB.n196 VPB.n195 0.735
R417 VPB.n195 VPB.n185 0.735
R418 VPB.n251 VPB.n250 0.387
R419 VPB.n251 VPB.n246 0.387
R420 VPB.n251 VPB.n241 0.387
R421 VPB.n252 VPB.n251 0.387
R422 VPB.n135 VPB.n134 0.387
R423 VPB.n135 VPB.n130 0.387
R424 VPB.n135 VPB.n125 0.387
R425 VPB.n136 VPB.n135 0.387
R426 VPB.n114 VPB.n113 0.387
R427 VPB.n114 VPB.n109 0.387
R428 VPB.n114 VPB.n104 0.387
R429 VPB.n115 VPB.n114 0.387
R430 VPB.n337 VPB.n336 0.387
R431 VPB.n337 VPB.n332 0.387
R432 VPB.n337 VPB.n327 0.387
R433 VPB.n338 VPB.n337 0.387
R434 VPB.n384 VPB.n383 0.387
R435 VPB.n384 VPB.n379 0.387
R436 VPB.n384 VPB.n374 0.387
R437 VPB.n385 VPB.n384 0.387
R438 VPB.n52 VPB.n51 0.387
R439 VPB.n52 VPB.n47 0.387
R440 VPB.n52 VPB.n42 0.387
R441 VPB.n53 VPB.n52 0.387
R442 VPB.n31 VPB.n30 0.387
R443 VPB.n31 VPB.n26 0.387
R444 VPB.n31 VPB.n21 0.387
R445 VPB.n32 VPB.n31 0.387
R446 VPB.n447 VPB.n13 0.387
R447 VPB.n447 VPB.n9 0.387
R448 VPB.n447 VPB.n4 0.387
R449 VPB.n447 VPB.n446 0.387
R450 VPB.n260 VPB.n233 0.272
R451 VPB.n293 VPB.n292 0.272
R452 VPB.n298 VPB.n297 0.272
R453 VPB.n346 VPB.n319 0.272
R454 VPB.n393 VPB.n366 0.272
R455 VPB.n430 VPB.n429 0.272
R456 VPB.n435 VPB.n434 0.272
R457 VPB.n439 VPB 0.198
R458 VPB.n213 VPB.n212 0.136
R459 VPB.n218 VPB.n213 0.136
R460 VPB.n225 VPB.n218 0.136
R461 VPB.n229 VPB.n225 0.136
R462 VPB.n233 VPB.n229 0.136
R463 VPB.n264 VPB.n260 0.136
R464 VPB.n268 VPB.n264 0.136
R465 VPB.n272 VPB.n268 0.136
R466 VPB.n277 VPB.n272 0.136
R467 VPB.n284 VPB.n277 0.136
R468 VPB.n288 VPB.n284 0.136
R469 VPB.n292 VPB.n288 0.136
R470 VPB.n294 VPB.n293 0.136
R471 VPB.n295 VPB.n294 0.136
R472 VPB.n296 VPB.n295 0.136
R473 VPB.n297 VPB.n296 0.136
R474 VPB.n299 VPB.n298 0.136
R475 VPB.n300 VPB.n299 0.136
R476 VPB.n301 VPB.n300 0.136
R477 VPB.n302 VPB.n301 0.136
R478 VPB.n302 VPB.n95 0.136
R479 VPB.n315 VPB.n95 0.136
R480 VPB.n319 VPB.n315 0.136
R481 VPB.n352 VPB.n346 0.136
R482 VPB.n356 VPB.n352 0.136
R483 VPB.n362 VPB.n356 0.136
R484 VPB.n366 VPB.n362 0.136
R485 VPB.n398 VPB.n393 0.136
R486 VPB.n403 VPB.n398 0.136
R487 VPB.n410 VPB.n403 0.136
R488 VPB.n415 VPB.n410 0.136
R489 VPB.n420 VPB.n415 0.136
R490 VPB.n425 VPB.n420 0.136
R491 VPB.n429 VPB.n425 0.136
R492 VPB.n431 VPB.n430 0.136
R493 VPB.n432 VPB.n431 0.136
R494 VPB.n433 VPB.n432 0.136
R495 VPB.n434 VPB.n433 0.136
R496 VPB.n436 VPB.n435 0.136
R497 VPB.n437 VPB.n436 0.136
R498 VPB.n438 VPB.n437 0.136
R499 VPB.n439 VPB.n438 0.136
R500 a_185_182.n2 a_185_182.t3 480.392
R501 a_185_182.n4 a_185_182.t8 472.359
R502 a_185_182.n2 a_185_182.t6 403.272
R503 a_185_182.n4 a_185_182.t4 384.527
R504 a_185_182.n3 a_185_182.t5 240.421
R505 a_185_182.n5 a_185_182.t7 198.113
R506 a_185_182.n7 a_185_182.n1 193.696
R507 a_185_182.n9 a_185_182.n7 162.151
R508 a_185_182.n5 a_185_182.n4 146.66
R509 a_185_182.n3 a_185_182.n2 135.047
R510 a_185_182.n6 a_185_182.n3 79.491
R511 a_185_182.n7 a_185_182.n6 79.491
R512 a_185_182.n6 a_185_182.n5 76
R513 a_185_182.n9 a_185_182.n8 30
R514 a_185_182.n10 a_185_182.n0 24.383
R515 a_185_182.n10 a_185_182.n9 23.684
R516 a_185_182.n1 a_185_182.t2 14.282
R517 a_185_182.n1 a_185_182.t1 14.282
R518 a_2215_1004.n4 a_2215_1004.t5 512.525
R519 a_2215_1004.n4 a_2215_1004.t7 371.139
R520 a_2215_1004.n5 a_2215_1004.t6 220.263
R521 a_2215_1004.n8 a_2215_1004.n6 194.086
R522 a_2215_1004.n6 a_2215_1004.n3 162.547
R523 a_2215_1004.n5 a_2215_1004.n4 158.3
R524 a_2215_1004.n6 a_2215_1004.n5 153.043
R525 a_2215_1004.n3 a_2215_1004.n2 76.002
R526 a_2215_1004.n8 a_2215_1004.n7 30
R527 a_2215_1004.n9 a_2215_1004.n0 24.383
R528 a_2215_1004.n9 a_2215_1004.n8 23.684
R529 a_2215_1004.n1 a_2215_1004.t3 14.282
R530 a_2215_1004.n1 a_2215_1004.t4 14.282
R531 a_2215_1004.n2 a_2215_1004.t1 14.282
R532 a_2215_1004.n2 a_2215_1004.t0 14.282
R533 a_2215_1004.n3 a_2215_1004.n1 12.85
R534 a_3905_1005.n0 a_3905_1005.t0 101.66
R535 a_3905_1005.n0 a_3905_1005.t1 101.66
R536 a_3905_1005.n0 a_3905_1005.t3 14.294
R537 a_3905_1005.t2 a_3905_1005.n0 14.282
R538 a_629_182.n2 a_629_182.t5 480.392
R539 a_629_182.n2 a_629_182.t3 403.272
R540 a_629_182.n3 a_629_182.t4 293.527
R541 a_629_182.n6 a_629_182.n4 215.257
R542 a_629_182.n4 a_629_182.n3 153.315
R543 a_629_182.n4 a_629_182.n1 140.59
R544 a_629_182.n3 a_629_182.n2 81.941
R545 a_629_182.n6 a_629_182.n5 30
R546 a_629_182.n7 a_629_182.n0 24.383
R547 a_629_182.n7 a_629_182.n6 23.684
R548 a_629_182.n1 a_629_182.t2 14.282
R549 a_629_182.n1 a_629_182.t1 14.282
R550 a_3239_1005.t2 a_3239_1005.n0 101.66
R551 a_3239_1005.n0 a_3239_1005.t3 101.659
R552 a_3239_1005.n0 a_3239_1005.t0 14.294
R553 a_3239_1005.n0 a_3239_1005.t1 14.282
R554 a_2849_182.n2 a_2849_182.t3 470.752
R555 a_2849_182.n2 a_2849_182.t4 384.527
R556 a_2849_182.n3 a_2849_182.t5 277.772
R557 a_2849_182.n6 a_2849_182.n4 241.81
R558 a_2849_182.n4 a_2849_182.n3 156.307
R559 a_2849_182.n4 a_2849_182.n1 114.038
R560 a_2849_182.n3 a_2849_182.n2 67.114
R561 a_2849_182.n6 a_2849_182.n5 30
R562 a_2849_182.n7 a_2849_182.n0 24.383
R563 a_2849_182.n7 a_2849_182.n6 23.684
R564 a_2849_182.n1 a_2849_182.t2 14.282
R565 a_2849_182.n1 a_2849_182.t1 14.282
R566 a_3451_383.n2 a_3451_383.t5 470.752
R567 a_3451_383.n2 a_3451_383.t4 384.527
R568 a_3451_383.n3 a_3451_383.t6 251.219
R569 a_3451_383.n9 a_3451_383.n4 172.234
R570 a_3451_383.n4 a_3451_383.n3 154.947
R571 a_3451_383.n4 a_3451_383.n1 148.83
R572 a_3451_383.n9 a_3451_383.n8 118.016
R573 a_3451_383.n3 a_3451_383.n2 93.667
R574 a_3451_383.n12 a_3451_383.n0 55.263
R575 a_3451_383.n11 a_3451_383.n9 48.405
R576 a_3451_383.n8 a_3451_383.n7 30
R577 a_3451_383.n11 a_3451_383.n10 30
R578 a_3451_383.n12 a_3451_383.n11 25.263
R579 a_3451_383.n6 a_3451_383.n5 24.383
R580 a_3451_383.n8 a_3451_383.n6 23.684
R581 a_3451_383.n1 a_3451_383.t1 14.282
R582 a_3451_383.n1 a_3451_383.t0 14.282
R583 a_1000_73.n10 a_1000_73.n9 93.333
R584 a_1000_73.n2 a_1000_73.n1 41.622
R585 a_1000_73.n13 a_1000_73.n12 26.667
R586 a_1000_73.n6 a_1000_73.n5 24.977
R587 a_1000_73.t0 a_1000_73.n2 21.209
R588 a_1000_73.t0 a_1000_73.n3 11.595
R589 a_1000_73.t1 a_1000_73.n8 8.137
R590 a_1000_73.t0 a_1000_73.n0 6.109
R591 a_1000_73.t1 a_1000_73.n7 4.864
R592 a_1000_73.t0 a_1000_73.n4 3.871
R593 a_1000_73.t0 a_1000_73.n13 2.535
R594 a_1000_73.n13 a_1000_73.t1 1.145
R595 a_1000_73.n7 a_1000_73.n6 1.13
R596 a_1000_73.t1 a_1000_73.n11 0.804
R597 a_1000_73.n11 a_1000_73.n10 0.136
R598 VNB VNB.n461 300.778
R599 VNB.n249 VNB.n248 199.897
R600 VNB.n137 VNB.n136 199.897
R601 VNB.n110 VNB.n109 199.897
R602 VNB.n344 VNB.n343 199.897
R603 VNB.n396 VNB.n395 199.897
R604 VNB.n52 VNB.n51 199.897
R605 VNB.n25 VNB.n24 199.897
R606 VNB.n146 VNB.n144 154.509
R607 VNB.n258 VNB.n256 154.509
R608 VNB.n353 VNB.n351 154.509
R609 VNB.n166 VNB.n164 154.509
R610 VNB.n61 VNB.n59 154.509
R611 VNB.n405 VNB.n403 154.509
R612 VNB.n81 VNB.n79 154.509
R613 VNB.n316 VNB.n315 121.366
R614 VNB.n425 VNB.n424 84.842
R615 VNB.n202 VNB.n194 76.136
R616 VNB.n202 VNB.n201 76
R617 VNB.n325 VNB.n95 76
R618 VNB.n448 VNB.n447 76
R619 VNB.n437 VNB.n436 76
R620 VNB.n433 VNB.n432 76
R621 VNB.n429 VNB.n428 76
R622 VNB.n423 VNB.n422 76
R623 VNB.n419 VNB.n418 76
R624 VNB.n415 VNB.n414 76
R625 VNB.n411 VNB.n410 76
R626 VNB.n407 VNB.n406 76
R627 VNB.n385 VNB.n384 76
R628 VNB.n381 VNB.n380 76
R629 VNB.n373 VNB.n372 76
R630 VNB.n364 VNB.n363 76
R631 VNB.n355 VNB.n354 76
R632 VNB.n333 VNB.n332 76
R633 VNB.n329 VNB.n328 76
R634 VNB.n319 VNB.n314 76
R635 VNB.n304 VNB.n303 76
R636 VNB.n300 VNB.n299 76
R637 VNB.n292 VNB.n291 76
R638 VNB.n287 VNB.n286 76
R639 VNB.n279 VNB.n278 76
R640 VNB.n275 VNB.n274 76
R641 VNB.n268 VNB.n267 76
R642 VNB.n260 VNB.n259 76
R643 VNB.n238 VNB.n237 76
R644 VNB.n234 VNB.n233 76
R645 VNB.n226 VNB.n225 76
R646 VNB.n221 VNB.n220 76
R647 VNB.n213 VNB.n212 76
R648 VNB.n209 VNB.n208 76
R649 VNB.n320 VNB.n99 63.835
R650 VNB.n154 VNB.n153 49.896
R651 VNB.n371 VNB.n370 49.896
R652 VNB.n69 VNB.n68 49.896
R653 VNB.n89 VNB.n88 49.896
R654 VNB.n218 VNB.n217 36.937
R655 VNB.n284 VNB.n283 36.937
R656 VNB.n317 VNB.n316 36.937
R657 VNB.n427 VNB.n426 36.678
R658 VNB.n207 VNB.n206 36.267
R659 VNB.n273 VNB.n272 36.267
R660 VNB.n126 VNB.n125 35.01
R661 VNB.n359 VNB.n358 35.01
R662 VNB.n41 VNB.n40 35.01
R663 VNB.n14 VNB.n13 35.01
R664 VNB.t4 VNB.n118 32.601
R665 VNB.t8 VNB.n33 32.601
R666 VNB.t0 VNB.n6 32.601
R667 VNB.n357 VNB.n356 29.127
R668 VNB.n99 VNB.n98 28.421
R669 VNB.n323 VNB.n322 27.855
R670 VNB.n99 VNB.n97 25.263
R671 VNB.n97 VNB.n96 24.383
R672 VNB.n367 VNB.t9 20.794
R673 VNB.n194 VNB.n191 20.452
R674 VNB.n449 VNB.n448 20.452
R675 VNB.n148 VNB.n126 20.094
R676 VNB.n152 VNB.n123 20.094
R677 VNB.n159 VNB.n121 20.094
R678 VNB.n360 VNB.n359 20.094
R679 VNB.n369 VNB.n368 20.094
R680 VNB.n377 VNB.n376 20.094
R681 VNB.n63 VNB.n41 20.094
R682 VNB.n67 VNB.n38 20.094
R683 VNB.n74 VNB.n36 20.094
R684 VNB.n83 VNB.n14 20.094
R685 VNB.n87 VNB.n11 20.094
R686 VNB.n94 VNB.n9 20.094
R687 VNB.n223 VNB.n222 19.735
R688 VNB.n216 VNB.n215 19.735
R689 VNB.n205 VNB.n204 19.735
R690 VNB.n198 VNB.n197 19.735
R691 VNB.n230 VNB.n229 19.735
R692 VNB.n289 VNB.n288 19.735
R693 VNB.n282 VNB.n281 19.735
R694 VNB.n271 VNB.n270 19.735
R695 VNB.n264 VNB.n263 19.735
R696 VNB.n296 VNB.n295 19.735
R697 VNB.n204 VNB.t3 19.724
R698 VNB.n222 VNB.t6 19.724
R699 VNB.n270 VNB.t7 19.724
R700 VNB.n288 VNB.t1 19.724
R701 VNB.n126 VNB.n124 19.017
R702 VNB.n359 VNB.n357 19.017
R703 VNB.n41 VNB.n39 19.017
R704 VNB.n14 VNB.n12 19.017
R705 VNB.n120 VNB.t4 17.353
R706 VNB.n35 VNB.t8 17.353
R707 VNB.n8 VNB.t0 17.353
R708 VNB.n324 VNB.n323 16.721
R709 VNB.n201 VNB.n200 13.653
R710 VNB.n200 VNB.n199 13.653
R711 VNB.n208 VNB.n207 13.653
R712 VNB.n212 VNB.n211 13.653
R713 VNB.n211 VNB.n210 13.653
R714 VNB.n220 VNB.n219 13.653
R715 VNB.n219 VNB.n218 13.653
R716 VNB.n225 VNB.n224 13.653
R717 VNB.n233 VNB.n232 13.653
R718 VNB.n232 VNB.n231 13.653
R719 VNB.n237 VNB.n236 13.653
R720 VNB.n236 VNB.n235 13.653
R721 VNB.n259 VNB.n258 13.653
R722 VNB.n258 VNB.n257 13.653
R723 VNB.n267 VNB.n266 13.653
R724 VNB.n266 VNB.n265 13.653
R725 VNB.n274 VNB.n273 13.653
R726 VNB.n278 VNB.n277 13.653
R727 VNB.n277 VNB.n276 13.653
R728 VNB.n286 VNB.n285 13.653
R729 VNB.n285 VNB.n284 13.653
R730 VNB.n291 VNB.n290 13.653
R731 VNB.n299 VNB.n298 13.653
R732 VNB.n298 VNB.n297 13.653
R733 VNB.n303 VNB.n302 13.653
R734 VNB.n302 VNB.n301 13.653
R735 VNB.n147 VNB.n146 13.653
R736 VNB.n146 VNB.n145 13.653
R737 VNB.n151 VNB.n150 13.653
R738 VNB.n150 VNB.n149 13.653
R739 VNB.n155 VNB.n154 13.653
R740 VNB.n158 VNB.n157 13.653
R741 VNB.n157 VNB.n156 13.653
R742 VNB.n162 VNB.n161 13.653
R743 VNB.n161 VNB.n160 13.653
R744 VNB.n167 VNB.n166 13.653
R745 VNB.n166 VNB.n165 13.653
R746 VNB.n170 VNB.n169 13.653
R747 VNB.n169 VNB.n168 13.653
R748 VNB.n173 VNB.n172 13.653
R749 VNB.n172 VNB.n171 13.653
R750 VNB.n176 VNB.n175 13.653
R751 VNB.n175 VNB.n174 13.653
R752 VNB.n319 VNB.n318 13.653
R753 VNB.n318 VNB.n317 13.653
R754 VNB.n325 VNB.n324 13.653
R755 VNB.n328 VNB.n327 13.653
R756 VNB.n327 VNB.n326 13.653
R757 VNB.n332 VNB.n331 13.653
R758 VNB.n331 VNB.n330 13.653
R759 VNB.n354 VNB.n353 13.653
R760 VNB.n353 VNB.n352 13.653
R761 VNB.n363 VNB.n362 13.653
R762 VNB.n362 VNB.n361 13.653
R763 VNB.n372 VNB.n371 13.653
R764 VNB.n380 VNB.n379 13.653
R765 VNB.n379 VNB.n378 13.653
R766 VNB.n384 VNB.n383 13.653
R767 VNB.n383 VNB.n382 13.653
R768 VNB.n406 VNB.n405 13.653
R769 VNB.n405 VNB.n404 13.653
R770 VNB.n410 VNB.n409 13.653
R771 VNB.n409 VNB.n408 13.653
R772 VNB.n414 VNB.n413 13.653
R773 VNB.n413 VNB.n412 13.653
R774 VNB.n418 VNB.n417 13.653
R775 VNB.n417 VNB.n416 13.653
R776 VNB.n422 VNB.n421 13.653
R777 VNB.n421 VNB.n420 13.653
R778 VNB.n428 VNB.n427 13.653
R779 VNB.n432 VNB.n431 13.653
R780 VNB.n431 VNB.n430 13.653
R781 VNB.n436 VNB.n435 13.653
R782 VNB.n435 VNB.n434 13.653
R783 VNB.n62 VNB.n61 13.653
R784 VNB.n61 VNB.n60 13.653
R785 VNB.n66 VNB.n65 13.653
R786 VNB.n65 VNB.n64 13.653
R787 VNB.n70 VNB.n69 13.653
R788 VNB.n73 VNB.n72 13.653
R789 VNB.n72 VNB.n71 13.653
R790 VNB.n77 VNB.n76 13.653
R791 VNB.n76 VNB.n75 13.653
R792 VNB.n82 VNB.n81 13.653
R793 VNB.n81 VNB.n80 13.653
R794 VNB.n86 VNB.n85 13.653
R795 VNB.n85 VNB.n84 13.653
R796 VNB.n90 VNB.n89 13.653
R797 VNB.n93 VNB.n92 13.653
R798 VNB.n92 VNB.n91 13.653
R799 VNB.n448 VNB.n0 13.653
R800 VNB VNB.n0 13.653
R801 VNB.n194 VNB.n193 13.653
R802 VNB.n193 VNB.n192 13.653
R803 VNB.n456 VNB.n453 13.577
R804 VNB.n179 VNB.n177 13.276
R805 VNB.n191 VNB.n179 13.276
R806 VNB.n241 VNB.n239 13.276
R807 VNB.n254 VNB.n241 13.276
R808 VNB.n129 VNB.n127 13.276
R809 VNB.n142 VNB.n129 13.276
R810 VNB.n102 VNB.n100 13.276
R811 VNB.n115 VNB.n102 13.276
R812 VNB.n336 VNB.n334 13.276
R813 VNB.n349 VNB.n336 13.276
R814 VNB.n388 VNB.n386 13.276
R815 VNB.n401 VNB.n388 13.276
R816 VNB.n44 VNB.n42 13.276
R817 VNB.n57 VNB.n44 13.276
R818 VNB.n17 VNB.n15 13.276
R819 VNB.n30 VNB.n17 13.276
R820 VNB.n259 VNB.n255 13.276
R821 VNB.n147 VNB.n143 13.276
R822 VNB.n158 VNB.n155 13.276
R823 VNB.n163 VNB.n162 13.276
R824 VNB.n167 VNB.n163 13.276
R825 VNB.n170 VNB.n167 13.276
R826 VNB.n173 VNB.n170 13.276
R827 VNB.n176 VNB.n173 13.276
R828 VNB.n319 VNB.n176 13.276
R829 VNB.n328 VNB.n325 13.276
R830 VNB.n354 VNB.n350 13.276
R831 VNB.n406 VNB.n402 13.276
R832 VNB.n62 VNB.n58 13.276
R833 VNB.n73 VNB.n70 13.276
R834 VNB.n78 VNB.n77 13.276
R835 VNB.n82 VNB.n78 13.276
R836 VNB.n93 VNB.n90 13.276
R837 VNB.n3 VNB.n1 13.276
R838 VNB.n449 VNB.n3 13.276
R839 VNB.n152 VNB.n151 13.097
R840 VNB.n67 VNB.n66 13.097
R841 VNB.n87 VNB.n86 13.097
R842 VNB.n229 VNB.n228 12.837
R843 VNB.n295 VNB.n294 12.837
R844 VNB.n121 VNB.n120 12.837
R845 VNB.n376 VNB.n375 12.837
R846 VNB.n36 VNB.n35 12.837
R847 VNB.n9 VNB.n8 12.837
R848 VNB.n197 VNB.n196 11.605
R849 VNB.n263 VNB.n262 11.605
R850 VNB.n320 VNB.n319 10.764
R851 VNB.n196 VNB.n195 9.809
R852 VNB.n262 VNB.n261 9.809
R853 VNB.n162 VNB.n159 9.329
R854 VNB.n77 VNB.n74 9.329
R855 VNB.n448 VNB.n94 9.329
R856 VNB.n148 VNB.n147 8.97
R857 VNB.n63 VNB.n62 8.97
R858 VNB.n83 VNB.n82 8.97
R859 VNB.n228 VNB.n227 7.566
R860 VNB.n294 VNB.n293 7.566
R861 VNB.n120 VNB.n119 7.566
R862 VNB.n375 VNB.n374 7.566
R863 VNB.n35 VNB.n34 7.566
R864 VNB.n8 VNB.n7 7.566
R865 VNB.n458 VNB.n457 7.5
R866 VNB.n247 VNB.n246 7.5
R867 VNB.n243 VNB.n242 7.5
R868 VNB.n241 VNB.n240 7.5
R869 VNB.n254 VNB.n253 7.5
R870 VNB.n135 VNB.n134 7.5
R871 VNB.n131 VNB.n130 7.5
R872 VNB.n129 VNB.n128 7.5
R873 VNB.n142 VNB.n141 7.5
R874 VNB.n108 VNB.n107 7.5
R875 VNB.n104 VNB.n103 7.5
R876 VNB.n102 VNB.n101 7.5
R877 VNB.n115 VNB.n114 7.5
R878 VNB.n342 VNB.n341 7.5
R879 VNB.n338 VNB.n337 7.5
R880 VNB.n336 VNB.n335 7.5
R881 VNB.n349 VNB.n348 7.5
R882 VNB.n394 VNB.n393 7.5
R883 VNB.n390 VNB.n389 7.5
R884 VNB.n388 VNB.n387 7.5
R885 VNB.n401 VNB.n400 7.5
R886 VNB.n50 VNB.n49 7.5
R887 VNB.n46 VNB.n45 7.5
R888 VNB.n44 VNB.n43 7.5
R889 VNB.n57 VNB.n56 7.5
R890 VNB.n23 VNB.n22 7.5
R891 VNB.n19 VNB.n18 7.5
R892 VNB.n17 VNB.n16 7.5
R893 VNB.n30 VNB.n29 7.5
R894 VNB.n450 VNB.n449 7.5
R895 VNB.n3 VNB.n2 7.5
R896 VNB.n455 VNB.n454 7.5
R897 VNB.n185 VNB.n184 7.5
R898 VNB.n181 VNB.n180 7.5
R899 VNB.n179 VNB.n178 7.5
R900 VNB.n191 VNB.n190 7.5
R901 VNB.n255 VNB.n254 7.176
R902 VNB.n143 VNB.n142 7.176
R903 VNB.n163 VNB.n115 7.176
R904 VNB.n350 VNB.n349 7.176
R905 VNB.n402 VNB.n401 7.176
R906 VNB.n58 VNB.n57 7.176
R907 VNB.n78 VNB.n30 7.176
R908 VNB.t3 VNB.n203 7.04
R909 VNB.t7 VNB.n269 7.04
R910 VNB.n460 VNB.n458 7.011
R911 VNB.n250 VNB.n247 7.011
R912 VNB.n245 VNB.n243 7.011
R913 VNB.n138 VNB.n135 7.011
R914 VNB.n133 VNB.n131 7.011
R915 VNB.n111 VNB.n108 7.011
R916 VNB.n106 VNB.n104 7.011
R917 VNB.n345 VNB.n342 7.011
R918 VNB.n340 VNB.n338 7.011
R919 VNB.n397 VNB.n394 7.011
R920 VNB.n392 VNB.n390 7.011
R921 VNB.n53 VNB.n50 7.011
R922 VNB.n48 VNB.n46 7.011
R923 VNB.n26 VNB.n23 7.011
R924 VNB.n21 VNB.n19 7.011
R925 VNB.n187 VNB.n185 7.011
R926 VNB.n183 VNB.n181 7.011
R927 VNB.n253 VNB.n252 7.01
R928 VNB.n245 VNB.n244 7.01
R929 VNB.n250 VNB.n249 7.01
R930 VNB.n141 VNB.n140 7.01
R931 VNB.n133 VNB.n132 7.01
R932 VNB.n138 VNB.n137 7.01
R933 VNB.n114 VNB.n113 7.01
R934 VNB.n106 VNB.n105 7.01
R935 VNB.n111 VNB.n110 7.01
R936 VNB.n348 VNB.n347 7.01
R937 VNB.n340 VNB.n339 7.01
R938 VNB.n345 VNB.n344 7.01
R939 VNB.n400 VNB.n399 7.01
R940 VNB.n392 VNB.n391 7.01
R941 VNB.n397 VNB.n396 7.01
R942 VNB.n56 VNB.n55 7.01
R943 VNB.n48 VNB.n47 7.01
R944 VNB.n53 VNB.n52 7.01
R945 VNB.n29 VNB.n28 7.01
R946 VNB.n21 VNB.n20 7.01
R947 VNB.n26 VNB.n25 7.01
R948 VNB.n190 VNB.n189 7.01
R949 VNB.n183 VNB.n182 7.01
R950 VNB.n187 VNB.n186 7.01
R951 VNB.n460 VNB.n459 7.01
R952 VNB.n456 VNB.n455 6.788
R953 VNB.n451 VNB.n450 6.788
R954 VNB.n220 VNB.n216 6.638
R955 VNB.n286 VNB.n282 6.638
R956 VNB.n215 VNB.n214 5.774
R957 VNB.n281 VNB.n280 5.774
R958 VNB.n117 VNB.n116 4.551
R959 VNB.n366 VNB.n365 4.551
R960 VNB.n32 VNB.n31 4.551
R961 VNB.n5 VNB.n4 4.551
R962 VNB.n151 VNB.n148 4.305
R963 VNB.n363 VNB.n360 4.305
R964 VNB.n66 VNB.n63 4.305
R965 VNB.n86 VNB.n83 4.305
R966 VNB.n159 VNB.n158 3.947
R967 VNB.n380 VNB.n377 3.947
R968 VNB.n74 VNB.n73 3.947
R969 VNB.n94 VNB.n93 3.947
R970 VNB.n208 VNB.n205 2.511
R971 VNB.n225 VNB.n223 2.511
R972 VNB.n274 VNB.n271 2.511
R973 VNB.n291 VNB.n289 2.511
R974 VNB.n325 VNB.n320 2.511
R975 VNB.n428 VNB.n425 2.511
R976 VNB.t4 VNB.n117 2.238
R977 VNB.t9 VNB.n366 2.238
R978 VNB.t8 VNB.n32 2.238
R979 VNB.t0 VNB.n5 2.238
R980 VNB.n323 VNB.n321 1.99
R981 VNB.n201 VNB.n198 1.614
R982 VNB.n233 VNB.n230 1.614
R983 VNB.n267 VNB.n264 1.614
R984 VNB.n299 VNB.n296 1.614
R985 VNB.n461 VNB.n452 0.921
R986 VNB.n461 VNB.n456 0.476
R987 VNB.n461 VNB.n451 0.475
R988 VNB.n123 VNB.n122 0.358
R989 VNB.n368 VNB.n367 0.358
R990 VNB.n38 VNB.n37 0.358
R991 VNB.n11 VNB.n10 0.358
R992 VNB.n260 VNB.n238 0.272
R993 VNB.n305 VNB.n304 0.272
R994 VNB.n310 VNB.n309 0.272
R995 VNB.n355 VNB.n333 0.272
R996 VNB.n407 VNB.n385 0.272
R997 VNB.n438 VNB.n437 0.272
R998 VNB.n443 VNB.n442 0.272
R999 VNB.n251 VNB.n245 0.246
R1000 VNB.n252 VNB.n251 0.246
R1001 VNB.n251 VNB.n250 0.246
R1002 VNB.n139 VNB.n133 0.246
R1003 VNB.n140 VNB.n139 0.246
R1004 VNB.n139 VNB.n138 0.246
R1005 VNB.n112 VNB.n106 0.246
R1006 VNB.n113 VNB.n112 0.246
R1007 VNB.n112 VNB.n111 0.246
R1008 VNB.n346 VNB.n340 0.246
R1009 VNB.n347 VNB.n346 0.246
R1010 VNB.n346 VNB.n345 0.246
R1011 VNB.n398 VNB.n392 0.246
R1012 VNB.n399 VNB.n398 0.246
R1013 VNB.n398 VNB.n397 0.246
R1014 VNB.n54 VNB.n48 0.246
R1015 VNB.n55 VNB.n54 0.246
R1016 VNB.n54 VNB.n53 0.246
R1017 VNB.n27 VNB.n21 0.246
R1018 VNB.n28 VNB.n27 0.246
R1019 VNB.n27 VNB.n26 0.246
R1020 VNB.n188 VNB.n183 0.246
R1021 VNB.n189 VNB.n188 0.246
R1022 VNB.n188 VNB.n187 0.246
R1023 VNB.n461 VNB.n460 0.246
R1024 VNB.n447 VNB 0.198
R1025 VNB.n155 VNB.n152 0.179
R1026 VNB.n372 VNB.n369 0.179
R1027 VNB.n70 VNB.n67 0.179
R1028 VNB.n90 VNB.n87 0.179
R1029 VNB.n209 VNB.n202 0.136
R1030 VNB.n213 VNB.n209 0.136
R1031 VNB.n221 VNB.n213 0.136
R1032 VNB.n226 VNB.n221 0.136
R1033 VNB.n234 VNB.n226 0.136
R1034 VNB.n238 VNB.n234 0.136
R1035 VNB.n268 VNB.n260 0.136
R1036 VNB.n275 VNB.n268 0.136
R1037 VNB.n279 VNB.n275 0.136
R1038 VNB.n287 VNB.n279 0.136
R1039 VNB.n292 VNB.n287 0.136
R1040 VNB.n300 VNB.n292 0.136
R1041 VNB.n304 VNB.n300 0.136
R1042 VNB.n306 VNB.n305 0.136
R1043 VNB.n307 VNB.n306 0.136
R1044 VNB.n308 VNB.n307 0.136
R1045 VNB.n309 VNB.n308 0.136
R1046 VNB.n311 VNB.n310 0.136
R1047 VNB.n312 VNB.n311 0.136
R1048 VNB.n313 VNB.n312 0.136
R1049 VNB.n314 VNB.n313 0.136
R1050 VNB.n314 VNB.n95 0.136
R1051 VNB.n329 VNB.n95 0.136
R1052 VNB.n333 VNB.n329 0.136
R1053 VNB.n364 VNB.n355 0.136
R1054 VNB.n373 VNB.n364 0.136
R1055 VNB.n381 VNB.n373 0.136
R1056 VNB.n385 VNB.n381 0.136
R1057 VNB.n411 VNB.n407 0.136
R1058 VNB.n415 VNB.n411 0.136
R1059 VNB.n419 VNB.n415 0.136
R1060 VNB.n423 VNB.n419 0.136
R1061 VNB.n429 VNB.n423 0.136
R1062 VNB.n433 VNB.n429 0.136
R1063 VNB.n437 VNB.n433 0.136
R1064 VNB.n439 VNB.n438 0.136
R1065 VNB.n440 VNB.n439 0.136
R1066 VNB.n441 VNB.n440 0.136
R1067 VNB.n442 VNB.n441 0.136
R1068 VNB.n444 VNB.n443 0.136
R1069 VNB.n445 VNB.n444 0.136
R1070 VNB.n446 VNB.n445 0.136
R1071 VNB.n447 VNB.n446 0.136
R1072 a_2110_73.n12 a_2110_73.n11 26.811
R1073 a_2110_73.n6 a_2110_73.n5 24.977
R1074 a_2110_73.n2 a_2110_73.n1 24.877
R1075 a_2110_73.t0 a_2110_73.n2 12.677
R1076 a_2110_73.t0 a_2110_73.n3 11.595
R1077 a_2110_73.t1 a_2110_73.n8 8.137
R1078 a_2110_73.t0 a_2110_73.n4 7.273
R1079 a_2110_73.t0 a_2110_73.n0 6.109
R1080 a_2110_73.t1 a_2110_73.n7 4.864
R1081 a_2110_73.t0 a_2110_73.n12 2.074
R1082 a_2110_73.n7 a_2110_73.n6 1.13
R1083 a_2110_73.n12 a_2110_73.t1 0.937
R1084 a_2110_73.t1 a_2110_73.n10 0.804
R1085 a_2110_73.n10 a_2110_73.n9 0.136
C4 VPB VNB 18.15fF
C5 a_2110_73.n0 VNB 0.02fF
C6 a_2110_73.n1 VNB 0.10fF
C7 a_2110_73.n2 VNB 0.06fF
C8 a_2110_73.n3 VNB 0.06fF
C9 a_2110_73.n4 VNB 0.00fF
C10 a_2110_73.n5 VNB 0.04fF
C11 a_2110_73.n6 VNB 0.05fF
C12 a_2110_73.n7 VNB 0.02fF
C13 a_2110_73.n8 VNB 0.05fF
C14 a_2110_73.n9 VNB 0.08fF
C15 a_2110_73.n10 VNB 0.18fF
C16 a_2110_73.t1 VNB 0.24fF
C17 a_2110_73.n11 VNB 0.09fF
C18 a_2110_73.n12 VNB 0.00fF
C19 a_1000_73.n0 VNB 0.02fF
C20 a_1000_73.n1 VNB 0.10fF
C21 a_1000_73.n2 VNB 0.07fF
C22 a_1000_73.n3 VNB 0.05fF
C23 a_1000_73.n4 VNB 0.00fF
C24 a_1000_73.n5 VNB 0.04fF
C25 a_1000_73.n6 VNB 0.05fF
C26 a_1000_73.n7 VNB 0.02fF
C27 a_1000_73.n8 VNB 0.05fF
C28 a_1000_73.n9 VNB 0.02fF
C29 a_1000_73.n10 VNB 0.08fF
C30 a_1000_73.n11 VNB 0.18fF
C31 a_1000_73.t1 VNB 0.24fF
C32 a_1000_73.n12 VNB 0.09fF
C33 a_1000_73.n13 VNB 0.00fF
C34 a_3451_383.n0 VNB 0.05fF
C35 a_3451_383.n1 VNB 0.74fF
C36 a_3451_383.n2 VNB 0.36fF
C37 a_3451_383.n3 VNB 0.84fF
C38 a_3451_383.n4 VNB 0.84fF
C39 a_3451_383.n5 VNB 0.05fF
C40 a_3451_383.n6 VNB 0.06fF
C41 a_3451_383.n7 VNB 0.04fF
C42 a_3451_383.n8 VNB 0.21fF
C43 a_3451_383.n9 VNB 0.46fF
C44 a_3451_383.n10 VNB 0.04fF
C45 a_3451_383.n11 VNB 0.11fF
C46 a_3451_383.n12 VNB 0.05fF
C47 a_2849_182.n0 VNB 0.05fF
C48 a_2849_182.n1 VNB 0.82fF
C49 a_2849_182.n2 VNB 0.35fF
C50 a_2849_182.t5 VNB 0.70fF
C51 a_2849_182.n3 VNB 1.08fF
C52 a_2849_182.n4 VNB 1.15fF
C53 a_2849_182.n5 VNB 0.04fF
C54 a_2849_182.n6 VNB 0.40fF
C55 a_2849_182.n7 VNB 0.07fF
C56 a_3239_1005.n0 VNB 0.55fF
C57 a_629_182.n0 VNB 0.04fF
C58 a_629_182.n1 VNB 0.74fF
C59 a_629_182.n2 VNB 0.37fF
C60 a_629_182.n3 VNB 0.59fF
C61 a_629_182.n4 VNB 0.64fF
C62 a_629_182.n5 VNB 0.04fF
C63 a_629_182.n6 VNB 0.32fF
C64 a_629_182.n7 VNB 0.06fF
C65 a_3905_1005.n0 VNB 0.52fF
C66 a_2215_1004.n0 VNB 0.04fF
C67 a_2215_1004.n1 VNB 0.47fF
C68 a_2215_1004.n2 VNB 0.56fF
C69 a_2215_1004.n3 VNB 0.28fF
C70 a_2215_1004.n4 VNB 0.32fF
C71 a_2215_1004.t6 VNB 0.46fF
C72 a_2215_1004.n5 VNB 0.51fF
C73 a_2215_1004.n6 VNB 0.51fF
C74 a_2215_1004.n7 VNB 0.03fF
C75 a_2215_1004.n8 VNB 0.25fF
C76 a_2215_1004.n9 VNB 0.05fF
C77 a_185_182.n0 VNB 0.04fF
C78 a_185_182.n1 VNB 0.74fF
C79 a_185_182.n2 VNB 0.40fF
C80 a_185_182.n3 VNB 0.38fF
C81 a_185_182.n4 VNB 0.36fF
C82 a_185_182.t7 VNB 0.47fF
C83 a_185_182.n5 VNB 0.35fF
C84 a_185_182.n6 VNB 1.54fF
C85 a_185_182.n7 VNB 0.43fF
C86 a_185_182.n8 VNB 0.03fF
C87 a_185_182.n9 VNB 0.23fF
C88 a_185_182.n10 VNB 0.05fF
C89 VPB.n0 VNB 0.03fF
C90 VPB.n1 VNB 0.04fF
C91 VPB.n2 VNB 0.02fF
C92 VPB.n3 VNB 0.10fF
C93 VPB.n5 VNB 0.02fF
C94 VPB.n6 VNB 0.02fF
C95 VPB.n7 VNB 0.02fF
C96 VPB.n8 VNB 0.02fF
C97 VPB.n10 VNB 0.02fF
C98 VPB.n11 VNB 0.02fF
C99 VPB.n12 VNB 0.02fF
C100 VPB.n14 VNB 0.02fF
C101 VPB.n15 VNB 0.02fF
C102 VPB.n16 VNB 0.02fF
C103 VPB.n17 VNB 0.04fF
C104 VPB.n18 VNB 0.02fF
C105 VPB.n19 VNB 0.13fF
C106 VPB.n20 VNB 0.04fF
C107 VPB.n22 VNB 0.02fF
C108 VPB.n23 VNB 0.02fF
C109 VPB.n24 VNB 0.02fF
C110 VPB.n25 VNB 0.02fF
C111 VPB.n27 VNB 0.02fF
C112 VPB.n28 VNB 0.02fF
C113 VPB.n29 VNB 0.02fF
C114 VPB.n31 VNB 0.27fF
C115 VPB.n33 VNB 0.03fF
C116 VPB.n34 VNB 0.02fF
C117 VPB.n35 VNB 0.02fF
C118 VPB.n36 VNB 0.02fF
C119 VPB.n37 VNB 0.02fF
C120 VPB.n38 VNB 0.04fF
C121 VPB.n39 VNB 0.02fF
C122 VPB.n40 VNB 0.16fF
C123 VPB.n41 VNB 0.04fF
C124 VPB.n43 VNB 0.02fF
C125 VPB.n44 VNB 0.02fF
C126 VPB.n45 VNB 0.02fF
C127 VPB.n46 VNB 0.02fF
C128 VPB.n48 VNB 0.02fF
C129 VPB.n49 VNB 0.02fF
C130 VPB.n50 VNB 0.02fF
C131 VPB.n52 VNB 0.27fF
C132 VPB.n54 VNB 0.03fF
C133 VPB.n55 VNB 0.02fF
C134 VPB.n56 VNB 0.03fF
C135 VPB.n57 VNB 0.03fF
C136 VPB.n58 VNB 0.27fF
C137 VPB.n59 VNB 0.01fF
C138 VPB.n60 VNB 0.02fF
C139 VPB.n61 VNB 0.06fF
C140 VPB.n62 VNB 0.13fF
C141 VPB.n63 VNB 0.19fF
C142 VPB.n64 VNB 0.02fF
C143 VPB.n65 VNB 0.01fF
C144 VPB.n66 VNB 0.16fF
C145 VPB.n67 VNB 0.02fF
C146 VPB.n68 VNB 0.02fF
C147 VPB.n69 VNB 0.13fF
C148 VPB.n70 VNB 0.19fF
C149 VPB.n71 VNB 0.02fF
C150 VPB.n72 VNB 0.01fF
C151 VPB.n73 VNB 0.06fF
C152 VPB.n74 VNB 0.27fF
C153 VPB.n75 VNB 0.01fF
C154 VPB.n76 VNB 0.02fF
C155 VPB.n77 VNB 0.03fF
C156 VPB.n78 VNB 0.03fF
C157 VPB.n79 VNB 0.27fF
C158 VPB.n80 VNB 0.01fF
C159 VPB.n81 VNB 0.02fF
C160 VPB.n82 VNB 0.06fF
C161 VPB.n83 VNB 0.13fF
C162 VPB.n84 VNB 0.19fF
C163 VPB.n85 VNB 0.02fF
C164 VPB.n86 VNB 0.01fF
C165 VPB.n87 VNB 0.16fF
C166 VPB.n88 VNB 0.02fF
C167 VPB.n89 VNB 0.02fF
C168 VPB.n90 VNB 0.13fF
C169 VPB.n91 VNB 0.19fF
C170 VPB.n92 VNB 0.02fF
C171 VPB.n93 VNB 0.01fF
C172 VPB.n94 VNB 0.06fF
C173 VPB.n95 VNB 0.02fF
C174 VPB.n96 VNB 0.10fF
C175 VPB.n97 VNB 0.02fF
C176 VPB.n98 VNB 0.02fF
C177 VPB.n99 VNB 0.02fF
C178 VPB.n100 VNB 0.04fF
C179 VPB.n101 VNB 0.02fF
C180 VPB.n102 VNB 0.16fF
C181 VPB.n103 VNB 0.04fF
C182 VPB.n105 VNB 0.02fF
C183 VPB.n106 VNB 0.02fF
C184 VPB.n107 VNB 0.02fF
C185 VPB.n108 VNB 0.02fF
C186 VPB.n110 VNB 0.02fF
C187 VPB.n111 VNB 0.02fF
C188 VPB.n112 VNB 0.02fF
C189 VPB.n114 VNB 0.27fF
C190 VPB.n116 VNB 0.03fF
C191 VPB.n117 VNB 0.02fF
C192 VPB.n118 VNB 0.02fF
C193 VPB.n119 VNB 0.02fF
C194 VPB.n120 VNB 0.02fF
C195 VPB.n121 VNB 0.04fF
C196 VPB.n122 VNB 0.02fF
C197 VPB.n123 VNB 0.16fF
C198 VPB.n124 VNB 0.04fF
C199 VPB.n126 VNB 0.02fF
C200 VPB.n127 VNB 0.02fF
C201 VPB.n128 VNB 0.02fF
C202 VPB.n129 VNB 0.02fF
C203 VPB.n131 VNB 0.02fF
C204 VPB.n132 VNB 0.02fF
C205 VPB.n133 VNB 0.02fF
C206 VPB.n135 VNB 0.27fF
C207 VPB.n137 VNB 0.03fF
C208 VPB.n138 VNB 0.02fF
C209 VPB.n139 VNB 0.03fF
C210 VPB.n140 VNB 0.03fF
C211 VPB.n141 VNB 0.27fF
C212 VPB.n142 VNB 0.01fF
C213 VPB.n143 VNB 0.02fF
C214 VPB.n144 VNB 0.06fF
C215 VPB.n145 VNB 0.13fF
C216 VPB.n146 VNB 0.19fF
C217 VPB.n147 VNB 0.02fF
C218 VPB.n148 VNB 0.01fF
C219 VPB.n149 VNB 0.16fF
C220 VPB.n150 VNB 0.02fF
C221 VPB.n151 VNB 0.02fF
C222 VPB.n152 VNB 0.13fF
C223 VPB.n153 VNB 0.19fF
C224 VPB.n154 VNB 0.02fF
C225 VPB.n155 VNB 0.01fF
C226 VPB.n156 VNB 0.06fF
C227 VPB.n157 VNB 0.27fF
C228 VPB.n158 VNB 0.01fF
C229 VPB.n159 VNB 0.02fF
C230 VPB.n160 VNB 0.03fF
C231 VPB.n161 VNB 0.03fF
C232 VPB.n162 VNB 0.27fF
C233 VPB.n163 VNB 0.01fF
C234 VPB.n164 VNB 0.02fF
C235 VPB.n165 VNB 0.23fF
C236 VPB.n166 VNB 0.02fF
C237 VPB.n167 VNB 0.01fF
C238 VPB.n168 VNB 0.05fF
C239 VPB.n169 VNB 0.13fF
C240 VPB.n170 VNB 0.16fF
C241 VPB.n171 VNB 0.02fF
C242 VPB.n172 VNB 0.02fF
C243 VPB.n173 VNB 0.13fF
C244 VPB.n174 VNB 0.15fF
C245 VPB.n175 VNB 0.02fF
C246 VPB.n176 VNB 0.02fF
C247 VPB.n177 VNB 0.02fF
C248 VPB.n178 VNB 0.02fF
C249 VPB.n179 VNB 0.02fF
C250 VPB.n180 VNB 0.02fF
C251 VPB.n181 VNB 0.14fF
C252 VPB.n182 VNB 0.03fF
C253 VPB.n183 VNB 0.02fF
C254 VPB.n184 VNB 0.05fF
C255 VPB.n185 VNB 0.01fF
C256 VPB.n186 VNB 0.02fF
C257 VPB.n187 VNB 0.02fF
C258 VPB.n190 VNB 0.02fF
C259 VPB.n191 VNB 0.02fF
C260 VPB.n193 VNB 0.02fF
C261 VPB.n195 VNB 0.45fF
C262 VPB.n197 VNB 0.04fF
C263 VPB.n198 VNB 0.04fF
C264 VPB.n199 VNB 0.27fF
C265 VPB.n200 VNB 0.03fF
C266 VPB.n201 VNB 0.03fF
C267 VPB.n202 VNB 0.27fF
C268 VPB.n203 VNB 0.02fF
C269 VPB.n204 VNB 0.02fF
C270 VPB.n205 VNB 0.27fF
C271 VPB.n206 VNB 0.02fF
C272 VPB.n207 VNB 0.02fF
C273 VPB.n208 VNB 0.27fF
C274 VPB.n209 VNB 0.02fF
C275 VPB.n210 VNB 0.02fF
C276 VPB.n211 VNB 0.00fF
C277 VPB.n212 VNB 0.09fF
C278 VPB.n213 VNB 0.02fF
C279 VPB.n214 VNB 0.13fF
C280 VPB.n215 VNB 0.14fF
C281 VPB.n216 VNB 0.02fF
C282 VPB.n217 VNB 0.02fF
C283 VPB.n218 VNB 0.02fF
C284 VPB.n219 VNB 0.10fF
C285 VPB.n220 VNB 0.02fF
C286 VPB.n221 VNB 0.13fF
C287 VPB.n222 VNB 0.16fF
C288 VPB.n223 VNB 0.02fF
C289 VPB.n224 VNB 0.02fF
C290 VPB.n225 VNB 0.02fF
C291 VPB.n226 VNB 0.23fF
C292 VPB.n227 VNB 0.02fF
C293 VPB.n228 VNB 0.02fF
C294 VPB.n229 VNB 0.02fF
C295 VPB.n230 VNB 0.27fF
C296 VPB.n231 VNB 0.01fF
C297 VPB.n232 VNB 0.02fF
C298 VPB.n233 VNB 0.04fF
C299 VPB.n234 VNB 0.02fF
C300 VPB.n235 VNB 0.02fF
C301 VPB.n236 VNB 0.02fF
C302 VPB.n237 VNB 0.04fF
C303 VPB.n238 VNB 0.02fF
C304 VPB.n239 VNB 0.20fF
C305 VPB.n240 VNB 0.04fF
C306 VPB.n242 VNB 0.02fF
C307 VPB.n243 VNB 0.02fF
C308 VPB.n244 VNB 0.02fF
C309 VPB.n245 VNB 0.02fF
C310 VPB.n247 VNB 0.02fF
C311 VPB.n248 VNB 0.02fF
C312 VPB.n249 VNB 0.02fF
C313 VPB.n251 VNB 0.27fF
C314 VPB.n253 VNB 0.03fF
C315 VPB.n254 VNB 0.02fF
C316 VPB.n255 VNB 0.03fF
C317 VPB.n256 VNB 0.03fF
C318 VPB.n257 VNB 0.27fF
C319 VPB.n258 VNB 0.01fF
C320 VPB.n259 VNB 0.02fF
C321 VPB.n260 VNB 0.04fF
C322 VPB.n261 VNB 0.27fF
C323 VPB.n262 VNB 0.02fF
C324 VPB.n263 VNB 0.02fF
C325 VPB.n264 VNB 0.02fF
C326 VPB.n265 VNB 0.27fF
C327 VPB.n266 VNB 0.02fF
C328 VPB.n267 VNB 0.02fF
C329 VPB.n268 VNB 0.02fF
C330 VPB.n269 VNB 0.27fF
C331 VPB.n270 VNB 0.02fF
C332 VPB.n271 VNB 0.02fF
C333 VPB.n272 VNB 0.02fF
C334 VPB.n273 VNB 0.13fF
C335 VPB.n274 VNB 0.14fF
C336 VPB.n275 VNB 0.02fF
C337 VPB.n276 VNB 0.02fF
C338 VPB.n277 VNB 0.02fF
C339 VPB.n278 VNB 0.10fF
C340 VPB.n279 VNB 0.02fF
C341 VPB.n280 VNB 0.13fF
C342 VPB.n281 VNB 0.16fF
C343 VPB.n282 VNB 0.02fF
C344 VPB.n283 VNB 0.02fF
C345 VPB.n284 VNB 0.02fF
C346 VPB.n285 VNB 0.23fF
C347 VPB.n286 VNB 0.02fF
C348 VPB.n287 VNB 0.02fF
C349 VPB.n288 VNB 0.02fF
C350 VPB.n289 VNB 0.27fF
C351 VPB.n290 VNB 0.01fF
C352 VPB.n291 VNB 0.02fF
C353 VPB.n292 VNB 0.04fF
C354 VPB.n293 VNB 0.04fF
C355 VPB.n294 VNB 0.02fF
C356 VPB.n295 VNB 0.02fF
C357 VPB.n296 VNB 0.02fF
C358 VPB.n297 VNB 0.04fF
C359 VPB.n298 VNB 0.04fF
C360 VPB.n299 VNB 0.02fF
C361 VPB.n300 VNB 0.02fF
C362 VPB.n301 VNB 0.02fF
C363 VPB.n302 VNB 0.02fF
C364 VPB.n303 VNB 0.13fF
C365 VPB.n304 VNB 0.14fF
C366 VPB.n305 VNB 0.02fF
C367 VPB.n306 VNB 0.02fF
C368 VPB.n307 VNB 0.13fF
C369 VPB.n308 VNB 0.16fF
C370 VPB.n309 VNB 0.02fF
C371 VPB.n310 VNB 0.02fF
C372 VPB.n311 VNB 0.06fF
C373 VPB.n312 VNB 0.23fF
C374 VPB.n313 VNB 0.02fF
C375 VPB.n314 VNB 0.01fF
C376 VPB.n315 VNB 0.02fF
C377 VPB.n316 VNB 0.27fF
C378 VPB.n317 VNB 0.01fF
C379 VPB.n318 VNB 0.02fF
C380 VPB.n319 VNB 0.04fF
C381 VPB.n320 VNB 0.02fF
C382 VPB.n321 VNB 0.02fF
C383 VPB.n322 VNB 0.02fF
C384 VPB.n323 VNB 0.04fF
C385 VPB.n324 VNB 0.02fF
C386 VPB.n325 VNB 0.16fF
C387 VPB.n326 VNB 0.04fF
C388 VPB.n328 VNB 0.02fF
C389 VPB.n329 VNB 0.02fF
C390 VPB.n330 VNB 0.02fF
C391 VPB.n331 VNB 0.02fF
C392 VPB.n333 VNB 0.02fF
C393 VPB.n334 VNB 0.02fF
C394 VPB.n335 VNB 0.02fF
C395 VPB.n337 VNB 0.27fF
C396 VPB.n339 VNB 0.03fF
C397 VPB.n340 VNB 0.02fF
C398 VPB.n341 VNB 0.03fF
C399 VPB.n342 VNB 0.03fF
C400 VPB.n343 VNB 0.27fF
C401 VPB.n344 VNB 0.01fF
C402 VPB.n345 VNB 0.02fF
C403 VPB.n346 VNB 0.04fF
C404 VPB.n347 VNB 0.06fF
C405 VPB.n348 VNB 0.13fF
C406 VPB.n349 VNB 0.19fF
C407 VPB.n350 VNB 0.02fF
C408 VPB.n351 VNB 0.01fF
C409 VPB.n352 VNB 0.02fF
C410 VPB.n353 VNB 0.16fF
C411 VPB.n354 VNB 0.02fF
C412 VPB.n355 VNB 0.02fF
C413 VPB.n356 VNB 0.02fF
C414 VPB.n357 VNB 0.06fF
C415 VPB.n358 VNB 0.13fF
C416 VPB.n359 VNB 0.19fF
C417 VPB.n360 VNB 0.02fF
C418 VPB.n361 VNB 0.01fF
C419 VPB.n362 VNB 0.02fF
C420 VPB.n363 VNB 0.27fF
C421 VPB.n364 VNB 0.01fF
C422 VPB.n365 VNB 0.02fF
C423 VPB.n366 VNB 0.04fF
C424 VPB.n367 VNB 0.02fF
C425 VPB.n368 VNB 0.02fF
C426 VPB.n369 VNB 0.02fF
C427 VPB.n370 VNB 0.04fF
C428 VPB.n371 VNB 0.02fF
C429 VPB.n372 VNB 0.16fF
C430 VPB.n373 VNB 0.04fF
C431 VPB.n375 VNB 0.02fF
C432 VPB.n376 VNB 0.02fF
C433 VPB.n377 VNB 0.02fF
C434 VPB.n378 VNB 0.02fF
C435 VPB.n380 VNB 0.02fF
C436 VPB.n381 VNB 0.02fF
C437 VPB.n382 VNB 0.02fF
C438 VPB.n384 VNB 0.27fF
C439 VPB.n386 VNB 0.03fF
C440 VPB.n387 VNB 0.02fF
C441 VPB.n388 VNB 0.03fF
C442 VPB.n389 VNB 0.03fF
C443 VPB.n390 VNB 0.27fF
C444 VPB.n391 VNB 0.01fF
C445 VPB.n392 VNB 0.02fF
C446 VPB.n393 VNB 0.04fF
C447 VPB.n394 VNB 0.05fF
C448 VPB.n395 VNB 0.23fF
C449 VPB.n396 VNB 0.02fF
C450 VPB.n397 VNB 0.01fF
C451 VPB.n398 VNB 0.02fF
C452 VPB.n399 VNB 0.13fF
C453 VPB.n400 VNB 0.16fF
C454 VPB.n401 VNB 0.02fF
C455 VPB.n402 VNB 0.02fF
C456 VPB.n403 VNB 0.02fF
C457 VPB.n404 VNB 0.10fF
C458 VPB.n405 VNB 0.02fF
C459 VPB.n406 VNB 0.13fF
C460 VPB.n407 VNB 0.15fF
C461 VPB.n408 VNB 0.02fF
C462 VPB.n409 VNB 0.02fF
C463 VPB.n410 VNB 0.02fF
C464 VPB.n411 VNB 0.13fF
C465 VPB.n412 VNB 0.14fF
C466 VPB.n413 VNB 0.02fF
C467 VPB.n414 VNB 0.02fF
C468 VPB.n415 VNB 0.02fF
C469 VPB.n416 VNB 0.13fF
C470 VPB.n417 VNB 0.16fF
C471 VPB.n418 VNB 0.02fF
C472 VPB.n419 VNB 0.02fF
C473 VPB.n420 VNB 0.02fF
C474 VPB.n421 VNB 0.06fF
C475 VPB.n422 VNB 0.23fF
C476 VPB.n423 VNB 0.02fF
C477 VPB.n424 VNB 0.01fF
C478 VPB.n425 VNB 0.02fF
C479 VPB.n426 VNB 0.27fF
C480 VPB.n427 VNB 0.01fF
C481 VPB.n428 VNB 0.02fF
C482 VPB.n429 VNB 0.04fF
C483 VPB.n430 VNB 0.04fF
C484 VPB.n431 VNB 0.02fF
C485 VPB.n432 VNB 0.02fF
C486 VPB.n433 VNB 0.02fF
C487 VPB.n434 VNB 0.04fF
C488 VPB.n435 VNB 0.04fF
C489 VPB.n436 VNB 0.02fF
C490 VPB.n437 VNB 0.02fF
C491 VPB.n438 VNB 0.02fF
C492 VPB.n439 VNB 0.03fF
C493 VPB.n440 VNB 0.03fF
C494 VPB.n441 VNB 0.02fF
C495 VPB.n442 VNB 0.02fF
C496 VPB.n443 VNB 0.02fF
C497 VPB.n444 VNB 0.04fF
C498 VPB.n445 VNB 0.04fF
C499 VPB.n447 VNB 0.42fF
C500 a_1739_182.n0 VNB 0.05fF
C501 a_1739_182.n1 VNB 0.87fF
C502 a_1739_182.n2 VNB 0.41fF
C503 a_1739_182.n3 VNB 1.27fF
C504 a_1739_182.n4 VNB 1.31fF
C505 a_1739_182.n5 VNB 0.04fF
C506 a_1739_182.n6 VNB 0.37fF
C507 a_1739_182.n7 VNB 0.07fF
C508 a_1105_1004.n0 VNB 0.05fF
C509 a_1105_1004.n1 VNB 0.50fF
C510 a_1105_1004.n2 VNB 0.59fF
C511 a_1105_1004.n3 VNB 0.30fF
C512 a_1105_1004.n4 VNB 0.33fF
C513 a_1105_1004.t6 VNB 0.49fF
C514 a_1105_1004.n5 VNB 0.54fF
C515 a_1105_1004.n6 VNB 0.53fF
C516 a_1105_1004.n7 VNB 0.02fF
C517 a_1105_1004.n8 VNB 0.26fF
C518 a_1105_1004.n9 VNB 0.04fF
.ends
