// File: DLATCH.spi.pex
// Created: Tue Oct 15 15:48:26 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_DLATCH\%GND ( 1 35 47 51 54 65 71 77 82 87 91 94 99 103 111 119 122 \
 127 131 153 157 165 169 177 181 189 193 201 205 217 228 231 243 245 257 277 \
 288 299 300 301 302 303 304 305 )
c278 ( 305 0 ) capacitor c=0.0706776f //x=17.21 //y=0.365
c279 ( 304 0 ) capacitor c=0.0706539f //x=13.88 //y=0.365
c280 ( 303 0 ) capacitor c=0.0578714f //x=11.595 //y=0.37
c281 ( 302 0 ) capacitor c=0.0207878f //x=8.76 //y=0.865
c282 ( 301 0 ) capacitor c=0.0572693f //x=6.045 //y=0.37
c283 ( 300 0 ) capacitor c=0.0208124f //x=3.21 //y=0.865
c284 ( 299 0 ) capacitor c=0.0589275f //x=0.495 //y=0.37
c285 ( 288 0 ) capacitor c=0.270488f //x=19.285 //y=0
c286 ( 277 0 ) capacitor c=0.10534f //x=16.65 //y=0
c287 ( 257 0 ) capacitor c=0.103812f //x=13.32 //y=0
c288 ( 245 0 ) capacitor c=0.10149f //x=11.1 //y=0
c289 ( 244 0 ) capacitor c=0.00440095f //x=8.95 //y=0
c290 ( 243 0 ) capacitor c=0.102231f //x=7.77 //y=0
c291 ( 231 0 ) capacitor c=0.10097f //x=5.55 //y=0
c292 ( 230 0 ) capacitor c=0.00440095f //x=3.33 //y=0
c293 ( 228 0 ) capacitor c=0.103282f //x=2.22 //y=0
c294 ( 217 0 ) capacitor c=0.192978f //x=0.63 //y=0
c295 ( 208 0 ) capacitor c=0.00609805f //x=19.285 //y=0.445
c296 ( 205 0 ) capacitor c=0.00505637f //x=19.2 //y=0.53
c297 ( 204 0 ) capacitor c=0.00468234f //x=18.8 //y=0.445
c298 ( 201 0 ) capacitor c=0.00537084f //x=18.715 //y=0.53
c299 ( 196 0 ) capacitor c=0.00468234f //x=18.315 //y=0.445
c300 ( 193 0 ) capacitor c=0.00537084f //x=18.23 //y=0.53
c301 ( 192 0 ) capacitor c=0.00468234f //x=17.83 //y=0.445
c302 ( 189 0 ) capacitor c=0.00634502f //x=17.745 //y=0.53
c303 ( 184 0 ) capacitor c=0.00609805f //x=17.345 //y=0.445
c304 ( 181 0 ) capacitor c=0.0195795f //x=17.26 //y=0
c305 ( 178 0 ) capacitor c=0.0659516f //x=16.04 //y=0
c306 ( 177 0 ) capacitor c=0.0195795f //x=16.48 //y=0
c307 ( 172 0 ) capacitor c=0.00609805f //x=15.955 //y=0.445
c308 ( 169 0 ) capacitor c=0.00505127f //x=15.87 //y=0.53
c309 ( 168 0 ) capacitor c=0.00468234f //x=15.47 //y=0.445
c310 ( 165 0 ) capacitor c=0.00537002f //x=15.385 //y=0.53
c311 ( 160 0 ) capacitor c=0.00468234f //x=14.985 //y=0.445
c312 ( 157 0 ) capacitor c=0.00556167f //x=14.9 //y=0.53
c313 ( 156 0 ) capacitor c=0.00468234f //x=14.5 //y=0.445
c314 ( 153 0 ) capacitor c=0.00642891f //x=14.415 //y=0.53
c315 ( 148 0 ) capacitor c=0.00609805f //x=14.015 //y=0.445
c316 ( 143 0 ) capacitor c=0.0227441f //x=13.93 //y=0
c317 ( 140 0 ) capacitor c=0.0360689f //x=12.785 //y=0
c318 ( 139 0 ) capacitor c=0.0184787f //x=13.15 //y=0
c319 ( 134 0 ) capacitor c=0.00583665f //x=12.7 //y=0.45
c320 ( 131 0 ) capacitor c=0.00536917f //x=12.615 //y=0.535
c321 ( 130 0 ) capacitor c=0.00479856f //x=12.215 //y=0.45
c322 ( 127 0 ) capacitor c=0.00640467f //x=12.13 //y=0.535
c323 ( 122 0 ) capacitor c=0.00588377f //x=11.73 //y=0.45
c324 ( 119 0 ) capacitor c=0.0164879f //x=11.645 //y=0
c325 ( 111 0 ) capacitor c=0.0720403f //x=10.93 //y=0
c326 ( 103 0 ) capacitor c=0.0389171f //x=8.865 //y=0
c327 ( 100 0 ) capacitor c=0.0360881f //x=7.235 //y=0
c328 ( 99 0 ) capacitor c=0.0160123f //x=7.6 //y=0
c329 ( 94 0 ) capacitor c=0.00583665f //x=7.15 //y=0.45
c330 ( 91 0 ) capacitor c=0.00531808f //x=7.065 //y=0.535
c331 ( 90 0 ) capacitor c=0.00479856f //x=6.665 //y=0.45
c332 ( 87 0 ) capacitor c=0.006266f //x=6.58 //y=0.535
c333 ( 82 0 ) capacitor c=0.00588377f //x=6.18 //y=0.45
c334 ( 77 0 ) capacitor c=0.0164879f //x=6.095 //y=0
c335 ( 71 0 ) capacitor c=0.0722769f //x=5.38 //y=0
c336 ( 65 0 ) capacitor c=0.0426751f //x=3.315 //y=0
c337 ( 60 0 ) capacitor c=0.0360484f //x=1.685 //y=0
c338 ( 59 0 ) capacitor c=0.0184787f //x=2.05 //y=0
c339 ( 54 0 ) capacitor c=0.00583665f //x=1.6 //y=0.45
c340 ( 51 0 ) capacitor c=0.00539433f //x=1.515 //y=0.535
c341 ( 50 0 ) capacitor c=0.00479856f //x=1.115 //y=0.45
c342 ( 47 0 ) capacitor c=0.00707849f //x=1.03 //y=0.535
c343 ( 42 0 ) capacitor c=0.00592191f //x=0.63 //y=0.45
c344 ( 35 0 ) capacitor c=0.67826f //x=19.24 //y=0
r345 (  287 288 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=19.24 //y=0 //x2=19.285 //y2=0
r346 (  285 287 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=18.8 //y=0 //x2=19.24 //y2=0
r347 (  284 285 ) resistor r=10.7563 //w=0.357 //l=0.3 //layer=li \
 //thickness=0.1 //x=18.5 //y=0 //x2=18.8 //y2=0
r348 (  282 284 ) resistor r=6.63305 //w=0.357 //l=0.185 //layer=li \
 //thickness=0.1 //x=18.315 //y=0 //x2=18.5 //y2=0
r349 (  281 282 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.83 //y=0 //x2=18.315 //y2=0
r350 (  280 281 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=17.39 //y=0 //x2=17.83 //y2=0
r351 (  278 280 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=17.345 //y=0 //x2=17.39 //y2=0
r352 (  265 266 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=15.91 //y=0 //x2=15.955 //y2=0
r353 (  263 265 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=15.47 //y=0 //x2=15.91 //y2=0
r354 (  262 263 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.985 //y=0 //x2=15.47 //y2=0
r355 (  261 262 ) resistor r=6.63305 //w=0.357 //l=0.185 //layer=li \
 //thickness=0.1 //x=14.8 //y=0 //x2=14.985 //y2=0
r356 (  259 261 ) resistor r=10.7563 //w=0.357 //l=0.3 //layer=li \
 //thickness=0.1 //x=14.5 //y=0 //x2=14.8 //y2=0
r357 (  258 259 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.015 //y=0 //x2=14.5 //y2=0
r358 (  249 250 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.215 //y=0 //x2=12.7 //y2=0
r359 (  248 249 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=12.21 //y=0 //x2=12.215 //y2=0
r360 (  246 248 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=11.73 //y=0 //x2=12.21 //y2=0
r361 (  235 236 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=7.03 //y=0 //x2=7.15 //y2=0
r362 (  233 235 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=6.665 //y=0 //x2=7.03 //y2=0
r363 (  232 233 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.18 //y=0 //x2=6.665 //y2=0
r364 (  220 221 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.115 //y=0 //x2=1.6 //y2=0
r365 (  219 220 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.115 //y2=0
r366 (  217 219 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=0.63 //y=0 //x2=0.74 //y2=0
r367 (  209 305 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.285 //y=0.615 //x2=19.285 //y2=0.53
r368 (  209 305 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=19.285 //y=0.615 //x2=19.285 //y2=0.88
r369 (  208 305 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.285 //y=0.445 //x2=19.285 //y2=0.53
r370 (  207 288 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.285 //y=0.17 //x2=19.285 //y2=0
r371 (  207 208 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=19.285 //y=0.17 //x2=19.285 //y2=0.445
r372 (  206 305 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.885 //y=0.53 //x2=18.8 //y2=0.53
r373 (  205 305 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.2 //y=0.53 //x2=19.285 //y2=0.53
r374 (  205 206 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=19.2 //y=0.53 //x2=18.885 //y2=0.53
r375 (  204 305 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.8 //y=0.445 //x2=18.8 //y2=0.53
r376 (  203 285 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.8 //y=0.17 //x2=18.8 //y2=0
r377 (  203 204 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=18.8 //y=0.17 //x2=18.8 //y2=0.445
r378 (  202 305 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=18.4 //y=0.53 //x2=18.315 //y2=0.53
r379 (  201 305 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.715 //y=0.53 //x2=18.8 //y2=0.53
r380 (  201 202 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=18.715 //y=0.53 //x2=18.4 //y2=0.53
r381 (  197 305 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=18.315 //y=0.615 //x2=18.315 //y2=0.53
r382 (  197 305 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.315 //y=0.615 //x2=18.315 //y2=0.88
r383 (  196 305 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=18.315 //y=0.445 //x2=18.315 //y2=0.53
r384 (  195 282 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.315 //y=0.17 //x2=18.315 //y2=0
r385 (  195 196 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=18.315 //y=0.17 //x2=18.315 //y2=0.445
r386 (  194 305 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.915 //y=0.53 //x2=17.83 //y2=0.53
r387 (  193 305 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=18.23 //y=0.53 //x2=18.315 //y2=0.53
r388 (  193 194 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=18.23 //y=0.53 //x2=17.915 //y2=0.53
r389 (  192 305 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.83 //y=0.445 //x2=17.83 //y2=0.53
r390 (  191 281 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.83 //y=0.17 //x2=17.83 //y2=0
r391 (  191 192 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=17.83 //y=0.17 //x2=17.83 //y2=0.445
r392 (  190 305 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.43 //y=0.53 //x2=17.345 //y2=0.53
r393 (  189 305 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.745 //y=0.53 //x2=17.83 //y2=0.53
r394 (  189 190 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=17.745 //y=0.53 //x2=17.43 //y2=0.53
r395 (  185 305 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.345 //y=0.615 //x2=17.345 //y2=0.53
r396 (  185 305 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=17.345 //y=0.615 //x2=17.345 //y2=1.22
r397 (  184 305 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.345 //y=0.445 //x2=17.345 //y2=0.53
r398 (  183 278 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.345 //y=0.17 //x2=17.345 //y2=0
r399 (  183 184 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=17.345 //y=0.17 //x2=17.345 //y2=0.445
r400 (  182 277 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.82 //y=0 //x2=16.65 //y2=0
r401 (  181 278 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.26 //y=0 //x2=17.345 //y2=0
r402 (  181 182 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=17.26 //y=0 //x2=16.82 //y2=0
r403 (  178 266 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.04 //y=0 //x2=15.955 //y2=0
r404 (  177 277 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.48 //y=0 //x2=16.65 //y2=0
r405 (  177 178 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=16.48 //y=0 //x2=16.04 //y2=0
r406 (  173 304 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.955 //y=0.615 //x2=15.955 //y2=0.53
r407 (  173 304 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.955 //y=0.615 //x2=15.955 //y2=0.88
r408 (  172 304 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.955 //y=0.445 //x2=15.955 //y2=0.53
r409 (  171 266 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.955 //y=0.17 //x2=15.955 //y2=0
r410 (  171 172 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=15.955 //y=0.17 //x2=15.955 //y2=0.445
r411 (  170 304 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.555 //y=0.53 //x2=15.47 //y2=0.53
r412 (  169 304 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.87 //y=0.53 //x2=15.955 //y2=0.53
r413 (  169 170 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=15.87 //y=0.53 //x2=15.555 //y2=0.53
r414 (  168 304 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.47 //y=0.445 //x2=15.47 //y2=0.53
r415 (  167 263 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.47 //y=0.17 //x2=15.47 //y2=0
r416 (  167 168 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=15.47 //y=0.17 //x2=15.47 //y2=0.445
r417 (  166 304 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=15.07 //y=0.53 //x2=14.985 //y2=0.53
r418 (  165 304 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.385 //y=0.53 //x2=15.47 //y2=0.53
r419 (  165 166 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=15.385 //y=0.53 //x2=15.07 //y2=0.53
r420 (  161 304 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=14.985 //y=0.615 //x2=14.985 //y2=0.53
r421 (  161 304 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=14.985 //y=0.615 //x2=14.985 //y2=0.88
r422 (  160 304 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=14.985 //y=0.445 //x2=14.985 //y2=0.53
r423 (  159 262 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.985 //y=0.17 //x2=14.985 //y2=0
r424 (  159 160 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=14.985 //y=0.17 //x2=14.985 //y2=0.445
r425 (  158 304 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.585 //y=0.53 //x2=14.5 //y2=0.53
r426 (  157 304 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=14.9 //y=0.53 //x2=14.985 //y2=0.53
r427 (  157 158 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=14.9 //y=0.53 //x2=14.585 //y2=0.53
r428 (  156 304 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.5 //y=0.445 //x2=14.5 //y2=0.53
r429 (  155 259 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.5 //y=0.17 //x2=14.5 //y2=0
r430 (  155 156 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=14.5 //y=0.17 //x2=14.5 //y2=0.445
r431 (  154 304 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.1 //y=0.53 //x2=14.015 //y2=0.53
r432 (  153 304 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.415 //y=0.53 //x2=14.5 //y2=0.53
r433 (  153 154 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=14.415 //y=0.53 //x2=14.1 //y2=0.53
r434 (  149 304 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.015 //y=0.615 //x2=14.015 //y2=0.53
r435 (  149 304 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=14.015 //y=0.615 //x2=14.015 //y2=1.22
r436 (  148 304 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.015 //y=0.445 //x2=14.015 //y2=0.53
r437 (  147 258 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.015 //y=0.17 //x2=14.015 //y2=0
r438 (  147 148 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=14.015 //y=0.17 //x2=14.015 //y2=0.445
r439 (  144 257 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.49 //y=0 //x2=13.32 //y2=0
r440 (  144 146 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=13.49 //y=0 //x2=13.69 //y2=0
r441 (  143 258 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.93 //y=0 //x2=14.015 //y2=0
r442 (  143 146 ) resistor r=8.60504 //w=0.357 //l=0.24 //layer=li \
 //thickness=0.1 //x=13.93 //y=0 //x2=13.69 //y2=0
r443 (  140 250 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.785 //y=0 //x2=12.7 //y2=0
r444 (  139 257 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.15 //y=0 //x2=13.32 //y2=0
r445 (  139 140 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=13.15 //y=0 //x2=12.785 //y2=0
r446 (  135 303 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.62 //x2=12.7 //y2=0.535
r447 (  135 303 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.62 //x2=12.7 //y2=1.225
r448 (  134 303 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.45 //x2=12.7 //y2=0.535
r449 (  133 250 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.17 //x2=12.7 //y2=0
r450 (  133 134 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.17 //x2=12.7 //y2=0.45
r451 (  132 303 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.3 //y=0.535 //x2=12.215 //y2=0.535
r452 (  131 303 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.615 //y=0.535 //x2=12.7 //y2=0.535
r453 (  131 132 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=12.615 //y=0.535 //x2=12.3 //y2=0.535
r454 (  130 303 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.215 //y=0.45 //x2=12.215 //y2=0.535
r455 (  129 249 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.215 //y=0.17 //x2=12.215 //y2=0
r456 (  129 130 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=12.215 //y=0.17 //x2=12.215 //y2=0.45
r457 (  128 303 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.815 //y=0.535 //x2=11.73 //y2=0.535
r458 (  127 303 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.13 //y=0.535 //x2=12.215 //y2=0.535
r459 (  127 128 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=12.13 //y=0.535 //x2=11.815 //y2=0.535
r460 (  123 303 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.62 //x2=11.73 //y2=0.535
r461 (  123 303 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.62 //x2=11.73 //y2=1.225
r462 (  122 303 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.45 //x2=11.73 //y2=0.535
r463 (  121 246 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.17 //x2=11.73 //y2=0
r464 (  121 122 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.17 //x2=11.73 //y2=0.45
r465 (  120 245 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.27 //y=0 //x2=11.1 //y2=0
r466 (  119 246 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.645 //y=0 //x2=11.73 //y2=0
r467 (  119 120 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=11.645 //y=0 //x2=11.27 //y2=0
r468 (  114 116 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=9.62 //y=0 //x2=10.73 //y2=0
r469 (  112 244 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.035 //y=0 //x2=8.95 //y2=0
r470 (  112 114 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=9.035 //y=0 //x2=9.62 //y2=0
r471 (  111 245 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.93 //y=0 //x2=11.1 //y2=0
r472 (  111 116 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=10.93 //y=0 //x2=10.73 //y2=0
r473 (  107 244 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.95 //y=0.17 //x2=8.95 //y2=0
r474 (  107 302 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=8.95 //y=0.17 //x2=8.95 //y2=0.955
r475 (  104 243 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.94 //y=0 //x2=7.77 //y2=0
r476 (  104 106 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=7.94 //y=0 //x2=8.51 //y2=0
r477 (  103 244 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.865 //y=0 //x2=8.95 //y2=0
r478 (  103 106 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=8.865 //y=0 //x2=8.51 //y2=0
r479 (  100 236 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.235 //y=0 //x2=7.15 //y2=0
r480 (  99 243 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.6 //y=0 //x2=7.77 //y2=0
r481 (  99 100 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=7.6 //y=0 //x2=7.235 //y2=0
r482 (  95 301 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.62 //x2=7.15 //y2=0.535
r483 (  95 301 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.62 //x2=7.15 //y2=1.225
r484 (  94 301 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.45 //x2=7.15 //y2=0.535
r485 (  93 236 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.17 //x2=7.15 //y2=0
r486 (  93 94 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.17 //x2=7.15 //y2=0.45
r487 (  92 301 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.75 //y=0.535 //x2=6.665 //y2=0.535
r488 (  91 301 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.065 //y=0.535 //x2=7.15 //y2=0.535
r489 (  91 92 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=7.065 //y=0.535 //x2=6.75 //y2=0.535
r490 (  90 301 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.665 //y=0.45 //x2=6.665 //y2=0.535
r491 (  89 233 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.665 //y=0.17 //x2=6.665 //y2=0
r492 (  89 90 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=6.665 //y=0.17 //x2=6.665 //y2=0.45
r493 (  88 301 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.265 //y=0.535 //x2=6.18 //y2=0.535
r494 (  87 301 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.58 //y=0.535 //x2=6.665 //y2=0.535
r495 (  87 88 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=6.58 //y=0.535 //x2=6.265 //y2=0.535
r496 (  83 301 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.62 //x2=6.18 //y2=0.535
r497 (  83 301 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.62 //x2=6.18 //y2=1.225
r498 (  82 301 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.45 //x2=6.18 //y2=0.535
r499 (  81 232 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.17 //x2=6.18 //y2=0
r500 (  81 82 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.17 //x2=6.18 //y2=0.45
r501 (  78 231 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.55 //y2=0
r502 (  78 80 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.92 //y2=0
r503 (  77 232 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.095 //y=0 //x2=6.18 //y2=0
r504 (  77 80 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=6.095 //y=0 //x2=5.92 //y2=0
r505 (  72 230 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.485 //y=0 //x2=3.4 //y2=0
r506 (  72 74 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=3.485 //y=0 //x2=4.44 //y2=0
r507 (  71 231 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=5.55 //y2=0
r508 (  71 74 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=4.44 //y2=0
r509 (  67 230 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.4 //y=0.17 //x2=3.4 //y2=0
r510 (  67 300 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=3.4 //y=0.17 //x2=3.4 //y2=0.955
r511 (  66 228 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.39 //y=0 //x2=2.22 //y2=0
r512 (  65 230 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.315 //y=0 //x2=3.4 //y2=0
r513 (  65 66 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=3.315 //y=0 //x2=2.39 //y2=0
r514 (  60 221 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.6 //y2=0
r515 (  60 62 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.85 //y2=0
r516 (  59 228 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=2.22 //y2=0
r517 (  59 62 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=1.85 //y2=0
r518 (  55 299 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=0.535
r519 (  55 299 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=1.225
r520 (  54 299 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.45 //x2=1.6 //y2=0.535
r521 (  53 221 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0
r522 (  53 54 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0.45
r523 (  52 299 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.2 //y=0.535 //x2=1.115 //y2=0.535
r524 (  51 299 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.6 //y2=0.535
r525 (  51 52 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.2 //y2=0.535
r526 (  50 299 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.45 //x2=1.115 //y2=0.535
r527 (  49 220 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0
r528 (  49 50 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0.45
r529 (  48 299 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.715 //y=0.535 //x2=0.63 //y2=0.535
r530 (  47 299 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=1.115 //y2=0.535
r531 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=0.715 //y2=0.535
r532 (  43 299 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=0.535
r533 (  43 299 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=1.225
r534 (  42 299 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.45 //x2=0.63 //y2=0.535
r535 (  41 217 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0
r536 (  41 42 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0.45
r537 (  35 287 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=19.24 //y=0 //x2=19.24 //y2=0
r538 (  33 284 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=0 //x2=18.5 //y2=0
r539 (  33 35 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=0 //x2=19.24 //y2=0
r540 (  31 280 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=0 //x2=17.39 //y2=0
r541 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=0 //x2=18.5 //y2=0
r542 (  29 265 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.91 //y=0 //x2=15.91 //y2=0
r543 (  29 31 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.91 //y=0 //x2=17.39 //y2=0
r544 (  27 261 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.8 //y=0 //x2=14.8 //y2=0
r545 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.8 //y=0 //x2=15.91 //y2=0
r546 (  25 146 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=0 //x2=13.69 //y2=0
r547 (  25 27 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=0 //x2=14.8 //y2=0
r548 (  23 248 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.21 //y=0 //x2=12.21 //y2=0
r549 (  23 25 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=0 //x2=13.69 //y2=0
r550 (  21 116 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=0 //x2=10.73 //y2=0
r551 (  21 23 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=0 //x2=12.21 //y2=0
r552 (  18 114 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=0 //x2=9.62 //y2=0
r553 (  16 106 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.51 //y=0 //x2=8.51 //y2=0
r554 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.51 //y=0 //x2=9.62 //y2=0
r555 (  14 235 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=0 //x2=7.03 //y2=0
r556 (  14 16 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=0 //x2=8.51 //y2=0
r557 (  12 80 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=0 //x2=5.92 //y2=0
r558 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=0 //x2=7.03 //y2=0
r559 (  10 74 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r560 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.92 //y2=0
r561 (  8 230 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=0 //x2=3.33 //y2=0
r562 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=0 //x2=4.44 //y2=0
r563 (  6 62 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r564 (  6 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=3.33 //y2=0
r565 (  3 219 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r566 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r567 (  1 21 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=9.99 //y=0 //x2=10.73 //y2=0
r568 (  1 18 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=9.99 //y=0 //x2=9.62 //y2=0
ends PM_DLATCH\%GND

subckt PM_DLATCH\%VDD ( 1 35 47 55 61 69 79 89 93 103 111 115 123 131 155 165 \
 169 179 187 202 206 208 212 216 221 224 226 228 229 230 231 232 233 234 235 \
 236 237 238 239 240 241 )
c267 ( 241 0 ) capacitor c=0.0255388f //x=17.735 //y=5.025
c268 ( 240 0 ) capacitor c=0.0255739f //x=14.405 //y=5.025
c269 ( 239 0 ) capacitor c=0.0433929f //x=12.51 //y=5.02
c270 ( 238 0 ) capacitor c=0.0422979f //x=11.64 //y=5.02
c271 ( 237 0 ) capacitor c=0.0382117f //x=10.175 //y=5.02
c272 ( 236 0 ) capacitor c=0.0240874f //x=9.295 //y=5.02
c273 ( 235 0 ) capacitor c=0.0494569f //x=8.425 //y=5.02
c274 ( 234 0 ) capacitor c=0.0432963f //x=6.96 //y=5.02
c275 ( 233 0 ) capacitor c=0.0422219f //x=6.09 //y=5.02
c276 ( 232 0 ) capacitor c=0.0381505f //x=4.625 //y=5.02
c277 ( 231 0 ) capacitor c=0.0240879f //x=3.745 //y=5.02
c278 ( 230 0 ) capacitor c=0.0494569f //x=2.875 //y=5.02
c279 ( 229 0 ) capacitor c=0.0432963f //x=1.41 //y=5.02
c280 ( 228 0 ) capacitor c=0.0421443f //x=0.54 //y=5.02
c281 ( 227 0 ) capacitor c=0.00591168f //x=17.88 //y=7.4
c282 ( 226 0 ) capacitor c=0.111374f //x=16.65 //y=7.4
c283 ( 225 0 ) capacitor c=0.00591168f //x=14.55 //y=7.4
c284 ( 224 0 ) capacitor c=0.109883f //x=13.32 //y=7.4
c285 ( 223 0 ) capacitor c=0.00591168f //x=12.655 //y=7.4
c286 ( 222 0 ) capacitor c=0.00591168f //x=11.775 //y=7.4
c287 ( 221 0 ) capacitor c=0.109921f //x=11.1 //y=7.4
c288 ( 220 0 ) capacitor c=0.00591168f //x=10.32 //y=7.4
c289 ( 219 0 ) capacitor c=0.00591168f //x=9.44 //y=7.4
c290 ( 218 0 ) capacitor c=0.00591168f //x=8.51 //y=7.4
c291 ( 216 0 ) capacitor c=0.114228f //x=7.77 //y=7.4
c292 ( 215 0 ) capacitor c=0.00591168f //x=7.03 //y=7.4
c293 ( 213 0 ) capacitor c=0.00591168f //x=6.225 //y=7.4
c294 ( 212 0 ) capacitor c=0.108342f //x=5.55 //y=7.4
c295 ( 211 0 ) capacitor c=0.00591168f //x=4.77 //y=7.4
c296 ( 210 0 ) capacitor c=0.00591168f //x=3.89 //y=7.4
c297 ( 209 0 ) capacitor c=0.00591168f //x=3.01 //y=7.4
c298 ( 208 0 ) capacitor c=0.114226f //x=2.22 //y=7.4
c299 ( 207 0 ) capacitor c=0.00591168f //x=1.555 //y=7.4
c300 ( 206 0 ) capacitor c=0.232987f //x=0.74 //y=7.4
c301 ( 202 0 ) capacitor c=0.287249f //x=19.24 //y=7.4
c302 ( 187 0 ) capacitor c=0.0427882f //x=17.795 //y=7.4
c303 ( 179 0 ) capacitor c=0.074729f //x=16.48 //y=7.4
c304 ( 169 0 ) capacitor c=0.0427882f //x=14.465 //y=7.4
c305 ( 165 0 ) capacitor c=0.0181526f //x=13.15 //y=7.4
c306 ( 155 0 ) capacitor c=0.0288426f //x=12.57 //y=7.4
c307 ( 147 0 ) capacitor c=0.0216067f //x=11.69 //y=7.4
c308 ( 141 0 ) capacitor c=0.0275781f //x=10.93 //y=7.4
c309 ( 131 0 ) capacitor c=0.0284327f //x=10.235 //y=7.4
c310 ( 123 0 ) capacitor c=0.0288633f //x=9.355 //y=7.4
c311 ( 115 0 ) capacitor c=0.0240981f //x=8.475 //y=7.4
c312 ( 111 0 ) capacitor c=0.0181526f //x=7.6 //y=7.4
c313 ( 103 0 ) capacitor c=0.0289624f //x=7.02 //y=7.4
c314 ( 93 0 ) capacitor c=0.0186283f //x=6.14 //y=7.4
c315 ( 89 0 ) capacitor c=0.0236224f //x=5.38 //y=7.4
c316 ( 79 0 ) capacitor c=0.0288639f //x=4.685 //y=7.4
c317 ( 69 0 ) capacitor c=0.0288633f //x=3.805 //y=7.4
c318 ( 61 0 ) capacitor c=0.0240981f //x=2.925 //y=7.4
c319 ( 55 0 ) capacitor c=0.0181526f //x=2.05 //y=7.4
c320 ( 47 0 ) capacitor c=0.0291066f //x=1.47 //y=7.4
c321 ( 35 0 ) capacitor c=0.691865f //x=19.24 //y=7.4
r322 (  200 202 ) resistor r=26.5322 //w=0.357 //l=0.74 //layer=li \
 //thickness=0.1 //x=18.5 //y=7.4 //x2=19.24 //y2=7.4
r323 (  198 227 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.965 //y=7.4 //x2=17.88 //y2=7.4
r324 (  198 200 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=17.965 //y=7.4 //x2=18.5 //y2=7.4
r325 (  191 227 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.88 //y=7.23 //x2=17.88 //y2=7.4
r326 (  191 241 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=17.88 //y=7.23 //x2=17.88 //y2=6.74
r327 (  188 226 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.82 //y=7.4 //x2=16.65 //y2=7.4
r328 (  188 190 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.82 //y=7.4 //x2=17.39 //y2=7.4
r329 (  187 227 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.795 //y=7.4 //x2=17.88 //y2=7.4
r330 (  187 190 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=17.795 //y=7.4 //x2=17.39 //y2=7.4
r331 (  182 184 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=14.8 //y=7.4 //x2=15.91 //y2=7.4
r332 (  180 225 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.635 //y=7.4 //x2=14.55 //y2=7.4
r333 (  180 182 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=14.635 //y=7.4 //x2=14.8 //y2=7.4
r334 (  179 226 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.48 //y=7.4 //x2=16.65 //y2=7.4
r335 (  179 184 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.48 //y=7.4 //x2=15.91 //y2=7.4
r336 (  173 225 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.55 //y=7.23 //x2=14.55 //y2=7.4
r337 (  173 240 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=14.55 //y=7.23 //x2=14.55 //y2=6.74
r338 (  170 224 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.49 //y=7.4 //x2=13.32 //y2=7.4
r339 (  170 172 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=13.49 //y=7.4 //x2=13.69 //y2=7.4
r340 (  169 225 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.465 //y=7.4 //x2=14.55 //y2=7.4
r341 (  169 172 ) resistor r=27.7871 //w=0.357 //l=0.775 //layer=li \
 //thickness=0.1 //x=14.465 //y=7.4 //x2=13.69 //y2=7.4
r342 (  166 223 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.74 //y=7.4 //x2=12.655 //y2=7.4
r343 (  165 224 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.15 //y=7.4 //x2=13.32 //y2=7.4
r344 (  165 166 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=13.15 //y=7.4 //x2=12.74 //y2=7.4
r345 (  159 223 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.655 //y=7.23 //x2=12.655 //y2=7.4
r346 (  159 239 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=12.655 //y=7.23 //x2=12.655 //y2=6.405
r347 (  156 222 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.86 //y=7.4 //x2=11.775 //y2=7.4
r348 (  156 158 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li \
 //thickness=0.1 //x=11.86 //y=7.4 //x2=12.21 //y2=7.4
r349 (  155 223 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.57 //y=7.4 //x2=12.655 //y2=7.4
r350 (  155 158 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=12.57 //y=7.4 //x2=12.21 //y2=7.4
r351 (  149 222 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.775 //y=7.23 //x2=11.775 //y2=7.4
r352 (  149 238 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=11.775 //y=7.23 //x2=11.775 //y2=6.405
r353 (  148 221 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.27 //y=7.4 //x2=11.1 //y2=7.4
r354 (  147 222 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.69 //y=7.4 //x2=11.775 //y2=7.4
r355 (  147 148 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=11.69 //y=7.4 //x2=11.27 //y2=7.4
r356 (  142 220 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.405 //y=7.4 //x2=10.32 //y2=7.4
r357 (  142 144 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=10.405 //y=7.4 //x2=10.73 //y2=7.4
r358 (  141 221 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.93 //y=7.4 //x2=11.1 //y2=7.4
r359 (  141 144 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=10.93 //y=7.4 //x2=10.73 //y2=7.4
r360 (  135 220 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.32 //y=7.23 //x2=10.32 //y2=7.4
r361 (  135 237 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.32 //y=7.23 //x2=10.32 //y2=6.745
r362 (  132 219 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.525 //y=7.4 //x2=9.44 //y2=7.4
r363 (  132 134 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=9.525 //y=7.4 //x2=9.62 //y2=7.4
r364 (  131 220 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.235 //y=7.4 //x2=10.32 //y2=7.4
r365 (  131 134 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.235 //y=7.4 //x2=9.62 //y2=7.4
r366 (  125 219 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.44 //y=7.23 //x2=9.44 //y2=7.4
r367 (  125 236 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.44 //y=7.23 //x2=9.44 //y2=6.745
r368 (  124 218 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.645 //y=7.4 //x2=8.56 //y2=7.4
r369 (  123 219 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.355 //y=7.4 //x2=9.44 //y2=7.4
r370 (  123 124 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=9.355 //y=7.4 //x2=8.645 //y2=7.4
r371 (  117 218 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.56 //y=7.23 //x2=8.56 //y2=7.4
r372 (  117 235 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=8.56 //y=7.23 //x2=8.56 //y2=6.405
r373 (  116 216 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.94 //y=7.4 //x2=7.77 //y2=7.4
r374 (  115 218 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.475 //y=7.4 //x2=8.56 //y2=7.4
r375 (  115 116 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=8.475 //y=7.4 //x2=7.94 //y2=7.4
r376 (  112 215 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.19 //y=7.4 //x2=7.105 //y2=7.4
r377 (  111 216 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.6 //y=7.4 //x2=7.77 //y2=7.4
r378 (  111 112 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=7.6 //y=7.4 //x2=7.19 //y2=7.4
r379 (  105 215 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.105 //y=7.23 //x2=7.105 //y2=7.4
r380 (  105 234 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=7.105 //y=7.23 //x2=7.105 //y2=6.405
r381 (  104 213 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.31 //y=7.4 //x2=6.225 //y2=7.4
r382 (  103 215 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.02 //y=7.4 //x2=7.105 //y2=7.4
r383 (  103 104 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.02 //y=7.4 //x2=6.31 //y2=7.4
r384 (  97 213 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.225 //y=7.23 //x2=6.225 //y2=7.4
r385 (  97 233 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=6.225 //y=7.23 //x2=6.225 //y2=6.405
r386 (  94 212 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.55 //y2=7.4
r387 (  94 96 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.92 //y2=7.4
r388 (  93 213 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.14 //y=7.4 //x2=6.225 //y2=7.4
r389 (  93 96 ) resistor r=7.88796 //w=0.357 //l=0.22 //layer=li \
 //thickness=0.1 //x=6.14 //y=7.4 //x2=5.92 //y2=7.4
r390 (  90 211 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.855 //y=7.4 //x2=4.77 //y2=7.4
r391 (  89 212 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=5.55 //y2=7.4
r392 (  89 90 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=4.855 //y2=7.4
r393 (  83 211 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.77 //y=7.23 //x2=4.77 //y2=7.4
r394 (  83 232 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.77 //y=7.23 //x2=4.77 //y2=6.745
r395 (  80 210 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.975 //y=7.4 //x2=3.89 //y2=7.4
r396 (  80 82 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=3.975 //y=7.4 //x2=4.44 //y2=7.4
r397 (  79 211 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.685 //y=7.4 //x2=4.77 //y2=7.4
r398 (  79 82 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=4.685 //y=7.4 //x2=4.44 //y2=7.4
r399 (  73 210 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.89 //y=7.23 //x2=3.89 //y2=7.4
r400 (  73 231 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.89 //y=7.23 //x2=3.89 //y2=6.745
r401 (  70 209 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.095 //y=7.4 //x2=3.01 //y2=7.4
r402 (  70 72 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=3.095 //y=7.4 //x2=3.33 //y2=7.4
r403 (  69 210 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.805 //y=7.4 //x2=3.89 //y2=7.4
r404 (  69 72 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=3.805 //y=7.4 //x2=3.33 //y2=7.4
r405 (  63 209 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.01 //y=7.23 //x2=3.01 //y2=7.4
r406 (  63 230 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=3.01 //y=7.23 //x2=3.01 //y2=6.405
r407 (  62 208 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.39 //y=7.4 //x2=2.22 //y2=7.4
r408 (  61 209 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.925 //y=7.4 //x2=3.01 //y2=7.4
r409 (  61 62 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=2.925 //y=7.4 //x2=2.39 //y2=7.4
r410 (  56 207 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.555 //y2=7.4
r411 (  56 58 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.85 //y2=7.4
r412 (  55 208 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.05 //y=7.4 //x2=2.22 //y2=7.4
r413 (  55 58 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=7.4 //x2=1.85 //y2=7.4
r414 (  49 207 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=7.4
r415 (  49 229 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=6.405
r416 (  48 206 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.76 //y=7.4 //x2=0.675 //y2=7.4
r417 (  47 207 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=1.555 //y2=7.4
r418 (  47 48 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=0.76 //y2=7.4
r419 (  41 206 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=7.4
r420 (  41 228 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=6.405
r421 (  35 202 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=19.24 //y=7.4 //x2=19.24 //y2=7.4
r422 (  33 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=7.4 //x2=18.5 //y2=7.4
r423 (  33 35 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=7.4 //x2=19.24 //y2=7.4
r424 (  31 190 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r425 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.4 //x2=18.5 //y2=7.4
r426 (  29 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.91 //y=7.4 //x2=15.91 //y2=7.4
r427 (  29 31 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.91 //y=7.4 //x2=17.39 //y2=7.4
r428 (  27 182 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.8 //y=7.4 //x2=14.8 //y2=7.4
r429 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.8 //y=7.4 //x2=15.91 //y2=7.4
r430 (  25 172 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=7.4 //x2=13.69 //y2=7.4
r431 (  25 27 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=7.4 //x2=14.8 //y2=7.4
r432 (  23 158 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.21 //y=7.4 //x2=12.21 //y2=7.4
r433 (  23 25 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=7.4 //x2=13.69 //y2=7.4
r434 (  21 144 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=7.4 //x2=10.73 //y2=7.4
r435 (  21 23 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=7.4 //x2=12.21 //y2=7.4
r436 (  18 134 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=7.4 //x2=9.62 //y2=7.4
r437 (  16 218 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.51 //y=7.4 //x2=8.51 //y2=7.4
r438 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.51 //y=7.4 //x2=9.62 //y2=7.4
r439 (  14 215 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=7.4 //x2=7.03 //y2=7.4
r440 (  14 16 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=7.4 //x2=8.51 //y2=7.4
r441 (  12 96 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=7.4 //x2=5.92 //y2=7.4
r442 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=7.4 //x2=7.03 //y2=7.4
r443 (  10 82 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r444 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.92 //y2=7.4
r445 (  8 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=7.4 //x2=3.33 //y2=7.4
r446 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=7.4 //x2=4.44 //y2=7.4
r447 (  6 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r448 (  6 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=3.33 //y2=7.4
r449 (  3 206 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r450 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r451 (  1 21 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=9.99 //y=7.4 //x2=10.73 //y2=7.4
r452 (  1 18 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=9.99 //y=7.4 //x2=9.62 //y2=7.4
ends PM_DLATCH\%VDD

subckt PM_DLATCH\%noxref_3 ( 1 2 17 18 19 20 24 26 33 34 35 36 37 38 39 43 45 \
 48 49 59 62 64 )
c117 ( 64 0 ) capacitor c=0.0288745f //x=0.97 //y=5.02
c118 ( 62 0 ) capacitor c=0.0173218f //x=0.925 //y=0.91
c119 ( 59 0 ) capacitor c=0.0593152f //x=3.33 //y=4.7
c120 ( 49 0 ) capacitor c=0.0318948f //x=3.665 //y=1.21
c121 ( 48 0 ) capacitor c=0.0187384f //x=3.665 //y=0.865
c122 ( 45 0 ) capacitor c=0.0141798f //x=3.51 //y=1.365
c123 ( 43 0 ) capacitor c=0.0149844f //x=3.51 //y=0.71
c124 ( 39 0 ) capacitor c=0.0860049f //x=3.135 //y=1.915
c125 ( 38 0 ) capacitor c=0.0229722f //x=3.135 //y=1.52
c126 ( 37 0 ) capacitor c=0.0234352f //x=3.135 //y=1.21
c127 ( 36 0 ) capacitor c=0.0199343f //x=3.135 //y=0.865
c128 ( 35 0 ) capacitor c=0.110275f //x=3.67 //y=6.02
c129 ( 34 0 ) capacitor c=0.154305f //x=3.23 //y=6.02
c130 ( 26 0 ) capacitor c=0.0954186f //x=3.33 //y=2.08
c131 ( 24 0 ) capacitor c=0.0861298f //x=1.48 //y=3.7
c132 ( 20 0 ) capacitor c=0.00417404f //x=1.2 //y=4.58
c133 ( 19 0 ) capacitor c=0.0118896f //x=1.395 //y=4.58
c134 ( 18 0 ) capacitor c=0.00621372f //x=1.195 //y=2.08
c135 ( 17 0 ) capacitor c=0.0139616f //x=1.395 //y=2.08
c136 ( 2 0 ) capacitor c=0.0139226f //x=1.595 //y=3.7
c137 ( 1 0 ) capacitor c=0.0681917f //x=3.215 //y=3.7
r138 (  57 59 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=3.23 //y=4.7 //x2=3.33 //y2=4.7
r139 (  50 59 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=3.67 //y=4.865 //x2=3.33 //y2=4.7
r140 (  49 61 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.665 //y=1.21 //x2=3.625 //y2=1.365
r141 (  48 60 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.665 //y=0.865 //x2=3.625 //y2=0.71
r142 (  48 49 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.665 //y=0.865 //x2=3.665 //y2=1.21
r143 (  46 56 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.29 //y=1.365 //x2=3.175 //y2=1.365
r144 (  45 61 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.51 //y=1.365 //x2=3.625 //y2=1.365
r145 (  44 55 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.29 //y=0.71 //x2=3.175 //y2=0.71
r146 (  43 60 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.51 //y=0.71 //x2=3.625 //y2=0.71
r147 (  43 44 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.51 //y=0.71 //x2=3.29 //y2=0.71
r148 (  40 57 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.23 //y=4.865 //x2=3.23 //y2=4.7
r149 (  39 54 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.915 //x2=3.33 //y2=2.08
r150 (  38 56 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.52 //x2=3.175 //y2=1.365
r151 (  38 39 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.52 //x2=3.135 //y2=1.915
r152 (  37 56 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.21 //x2=3.175 //y2=1.365
r153 (  36 55 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=0.865 //x2=3.175 //y2=0.71
r154 (  36 37 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.135 //y=0.865 //x2=3.135 //y2=1.21
r155 (  35 50 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.67 //y=6.02 //x2=3.67 //y2=4.865
r156 (  34 40 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.23 //y=6.02 //x2=3.23 //y2=4.865
r157 (  33 45 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.4 //y=1.365 //x2=3.51 //y2=1.365
r158 (  33 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.4 //y=1.365 //x2=3.29 //y2=1.365
r159 (  31 59 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r160 (  29 31 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=3.33 //y=3.7 //x2=3.33 //y2=4.7
r161 (  26 54 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r162 (  26 29 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.7
r163 (  22 24 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.48 //y=4.495 //x2=1.48 //y2=3.7
r164 (  21 24 ) resistor r=105.07 //w=0.187 //l=1.535 //layer=li \
 //thickness=0.1 //x=1.48 //y=2.165 //x2=1.48 //y2=3.7
r165 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.48 //y2=4.495
r166 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.2 //y2=4.58
r167 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.48 //y2=2.165
r168 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.195 //y2=2.08
r169 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.2 //y2=4.58
r170 (  11 64 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.115 //y2=5.725
r171 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.195 //y2=2.08
r172 (  7 62 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.11 //y2=1.005
r173 (  6 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.7 //x2=3.33 //y2=3.7
r174 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.48 //y=3.7 //x2=1.48 //y2=3.7
r175 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.595 //y=3.7 //x2=1.48 //y2=3.7
r176 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.215 //y=3.7 //x2=3.33 //y2=3.7
r177 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=3.215 //y=3.7 //x2=1.595 //y2=3.7
ends PM_DLATCH\%noxref_3

subckt PM_DLATCH\%noxref_4 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 \
 52 53 54 56 62 63 65 73 75 76 )
c134 ( 76 0 ) capacitor c=0.0220291f //x=4.185 //y=5.02
c135 ( 75 0 ) capacitor c=0.0217503f //x=3.305 //y=5.02
c136 ( 73 0 ) capacitor c=0.0084702f //x=4.18 //y=0.905
c137 ( 65 0 ) capacitor c=0.0511458f //x=6.29 //y=2.085
c138 ( 63 0 ) capacitor c=0.0435629f //x=6.93 //y=1.255
c139 ( 62 0 ) capacitor c=0.0200386f //x=6.93 //y=0.91
c140 ( 56 0 ) capacitor c=0.0152946f //x=6.775 //y=1.41
c141 ( 54 0 ) capacitor c=0.0157804f //x=6.775 //y=0.755
c142 ( 53 0 ) capacitor c=0.0490829f //x=6.52 //y=4.79
c143 ( 52 0 ) capacitor c=0.0303096f //x=6.81 //y=4.79
c144 ( 48 0 ) capacitor c=0.0290017f //x=6.4 //y=1.92
c145 ( 47 0 ) capacitor c=0.0250027f //x=6.4 //y=1.565
c146 ( 46 0 ) capacitor c=0.0234316f //x=6.4 //y=1.255
c147 ( 45 0 ) capacitor c=0.0200596f //x=6.4 //y=0.91
c148 ( 44 0 ) capacitor c=0.154218f //x=6.885 //y=6.02
c149 ( 43 0 ) capacitor c=0.154243f //x=6.445 //y=6.02
c150 ( 41 0 ) capacitor c=0.0023043f //x=4.33 //y=5.2
c151 ( 34 0 ) capacitor c=0.0884603f //x=6.29 //y=2.085
c152 ( 32 0 ) capacitor c=0.10682f //x=4.81 //y=3.33
c153 ( 28 0 ) capacitor c=0.00468667f //x=4.455 //y=1.655
c154 ( 27 0 ) capacitor c=0.0131863f //x=4.725 //y=1.655
c155 ( 25 0 ) capacitor c=0.0141863f //x=4.725 //y=5.2
c156 ( 14 0 ) capacitor c=0.00265825f //x=3.535 //y=5.2
c157 ( 13 0 ) capacitor c=0.0149089f //x=4.245 //y=5.2
c158 ( 2 0 ) capacitor c=0.0120846f //x=4.925 //y=3.33
c159 ( 1 0 ) capacitor c=0.0361557f //x=6.175 //y=3.33
r160 (  65 66 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.29 //y=2.085 //x2=6.4 //y2=2.085
r161 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.93 //y=1.255 //x2=6.89 //y2=1.41
r162 (  62 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.93 //y=0.91 //x2=6.89 //y2=0.755
r163 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.93 //y=0.91 //x2=6.93 //y2=1.255
r164 (  57 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.555 //y=1.41 //x2=6.44 //y2=1.41
r165 (  56 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.775 //y=1.41 //x2=6.89 //y2=1.41
r166 (  55 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.555 //y=0.755 //x2=6.44 //y2=0.755
r167 (  54 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.775 //y=0.755 //x2=6.89 //y2=0.755
r168 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.775 //y=0.755 //x2=6.555 //y2=0.755
r169 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.81 //y=4.79 //x2=6.885 //y2=4.865
r170 (  52 53 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=6.81 //y=4.79 //x2=6.52 //y2=4.79
r171 (  49 53 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.445 //y=4.865 //x2=6.52 //y2=4.79
r172 (  49 68 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=6.445 //y=4.865 //x2=6.29 //y2=4.7
r173 (  48 66 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.4 //y=1.92 //x2=6.4 //y2=2.085
r174 (  47 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.4 //y=1.565 //x2=6.44 //y2=1.41
r175 (  47 48 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=6.4 //y=1.565 //x2=6.4 //y2=1.92
r176 (  46 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.4 //y=1.255 //x2=6.44 //y2=1.41
r177 (  45 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.4 //y=0.91 //x2=6.44 //y2=0.755
r178 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.4 //y=0.91 //x2=6.4 //y2=1.255
r179 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.885 //y=6.02 //x2=6.885 //y2=4.865
r180 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.445 //y=6.02 //x2=6.445 //y2=4.865
r181 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.665 //y=1.41 //x2=6.775 //y2=1.41
r182 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.665 //y=1.41 //x2=6.555 //y2=1.41
r183 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.29 //y=4.7 //x2=6.29 //y2=4.7
r184 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=6.29 //y=3.33 //x2=6.29 //y2=4.7
r185 (  34 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.29 //y=2.085 //x2=6.29 //y2=2.085
r186 (  34 37 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=6.29 //y=2.085 //x2=6.29 //y2=3.33
r187 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=4.81 //y=5.115 //x2=4.81 //y2=3.33
r188 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=4.81 //y=1.74 //x2=4.81 //y2=3.33
r189 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=1.655 //x2=4.81 //y2=1.74
r190 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=4.725 //y=1.655 //x2=4.455 //y2=1.655
r191 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.415 //y=5.2 //x2=4.33 //y2=5.2
r192 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=5.2 //x2=4.81 //y2=5.115
r193 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=4.725 //y=5.2 //x2=4.415 //y2=5.2
r194 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.37 //y=1.57 //x2=4.455 //y2=1.655
r195 (  21 73 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.37 //y=1.57 //x2=4.37 //y2=1
r196 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.33 //y=5.285 //x2=4.33 //y2=5.2
r197 (  15 76 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=4.33 //y=5.285 //x2=4.33 //y2=5.725
r198 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.245 //y=5.2 //x2=4.33 //y2=5.2
r199 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=4.245 //y=5.2 //x2=3.535 //y2=5.2
r200 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.45 //y=5.285 //x2=3.535 //y2=5.2
r201 (  7 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=3.45 //y=5.285 //x2=3.45 //y2=5.725
r202 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.29 //y=3.33 //x2=6.29 //y2=3.33
r203 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.81 //y=3.33 //x2=4.81 //y2=3.33
r204 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.925 //y=3.33 //x2=4.81 //y2=3.33
r205 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.175 //y=3.33 //x2=6.29 //y2=3.33
r206 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=6.175 //y=3.33 //x2=4.925 //y2=3.33
ends PM_DLATCH\%noxref_4

subckt PM_DLATCH\%GATE ( 1 2 7 8 9 10 11 12 13 14 15 16 18 27 39 40 41 42 43 \
 44 45 46 47 52 54 56 62 63 64 65 66 67 71 73 76 77 82 83 86 100 )
c161 ( 100 0 ) capacitor c=0.0593152f //x=8.88 //y=4.7
c162 ( 86 0 ) capacitor c=0.0331552f //x=4.1 //y=4.7
c163 ( 83 0 ) capacitor c=0.0279499f //x=4.07 //y=1.915
c164 ( 82 0 ) capacitor c=0.0422509f //x=4.07 //y=2.08
c165 ( 77 0 ) capacitor c=0.0318948f //x=9.215 //y=1.21
c166 ( 76 0 ) capacitor c=0.0187384f //x=9.215 //y=0.865
c167 ( 73 0 ) capacitor c=0.0141798f //x=9.06 //y=1.365
c168 ( 71 0 ) capacitor c=0.0149844f //x=9.06 //y=0.71
c169 ( 67 0 ) capacitor c=0.0819722f //x=8.685 //y=1.915
c170 ( 66 0 ) capacitor c=0.0229722f //x=8.685 //y=1.52
c171 ( 65 0 ) capacitor c=0.0234352f //x=8.685 //y=1.21
c172 ( 64 0 ) capacitor c=0.0199343f //x=8.685 //y=0.865
c173 ( 63 0 ) capacitor c=0.0429696f //x=4.635 //y=1.25
c174 ( 62 0 ) capacitor c=0.0192208f //x=4.635 //y=0.905
c175 ( 56 0 ) capacitor c=0.0158629f //x=4.48 //y=1.405
c176 ( 54 0 ) capacitor c=0.0157803f //x=4.48 //y=0.75
c177 ( 52 0 ) capacitor c=0.0300505f //x=4.475 //y=4.79
c178 ( 47 0 ) capacitor c=0.0205163f //x=4.105 //y=1.56
c179 ( 46 0 ) capacitor c=0.0168481f //x=4.105 //y=1.25
c180 ( 45 0 ) capacitor c=0.0174783f //x=4.105 //y=0.905
c181 ( 44 0 ) capacitor c=0.110275f //x=9.22 //y=6.02
c182 ( 43 0 ) capacitor c=0.154305f //x=8.78 //y=6.02
c183 ( 42 0 ) capacitor c=0.15358f //x=4.55 //y=6.02
c184 ( 41 0 ) capacitor c=0.110281f //x=4.11 //y=6.02
c185 ( 27 0 ) capacitor c=0.0925986f //x=8.88 //y=2.08
c186 ( 18 0 ) capacitor c=0.0756836f //x=4.07 //y=2.08
c187 ( 16 0 ) capacitor c=0.00453889f //x=4.07 //y=4.535
c188 ( 2 0 ) capacitor c=0.0165749f //x=4.185 //y=2.96
c189 ( 1 0 ) capacitor c=0.14924f //x=8.765 //y=2.96
r190 (  98 100 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=8.78 //y=4.7 //x2=8.88 //y2=4.7
r191 (  88 89 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=4.1 //y=4.79 //x2=4.1 //y2=4.865
r192 (  86 88 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=4.1 //y=4.7 //x2=4.1 //y2=4.79
r193 (  82 83 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=4.07 //y=2.08 //x2=4.07 //y2=1.915
r194 (  78 100 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=9.22 //y=4.865 //x2=8.88 //y2=4.7
r195 (  77 102 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.21 //x2=9.175 //y2=1.365
r196 (  76 101 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.215 //y=0.865 //x2=9.175 //y2=0.71
r197 (  76 77 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.215 //y=0.865 //x2=9.215 //y2=1.21
r198 (  74 97 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.84 //y=1.365 //x2=8.725 //y2=1.365
r199 (  73 102 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.06 //y=1.365 //x2=9.175 //y2=1.365
r200 (  72 96 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.84 //y=0.71 //x2=8.725 //y2=0.71
r201 (  71 101 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.06 //y=0.71 //x2=9.175 //y2=0.71
r202 (  71 72 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=9.06 //y=0.71 //x2=8.84 //y2=0.71
r203 (  68 98 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.78 //y=4.865 //x2=8.78 //y2=4.7
r204 (  67 95 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=8.685 //y=1.915 //x2=8.88 //y2=2.08
r205 (  66 97 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.685 //y=1.52 //x2=8.725 //y2=1.365
r206 (  66 67 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=8.685 //y=1.52 //x2=8.685 //y2=1.915
r207 (  65 97 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.685 //y=1.21 //x2=8.725 //y2=1.365
r208 (  64 96 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.685 //y=0.865 //x2=8.725 //y2=0.71
r209 (  64 65 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.685 //y=0.865 //x2=8.685 //y2=1.21
r210 (  63 93 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.635 //y=1.25 //x2=4.595 //y2=1.405
r211 (  62 92 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.635 //y=0.905 //x2=4.595 //y2=0.75
r212 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.635 //y=0.905 //x2=4.635 //y2=1.25
r213 (  57 91 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.26 //y=1.405 //x2=4.145 //y2=1.405
r214 (  56 93 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.48 //y=1.405 //x2=4.595 //y2=1.405
r215 (  55 90 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.26 //y=0.75 //x2=4.145 //y2=0.75
r216 (  54 92 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.48 //y=0.75 //x2=4.595 //y2=0.75
r217 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.48 //y=0.75 //x2=4.26 //y2=0.75
r218 (  53 88 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=4.235 //y=4.79 //x2=4.1 //y2=4.79
r219 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.475 //y=4.79 //x2=4.55 //y2=4.865
r220 (  52 53 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=4.475 //y=4.79 //x2=4.235 //y2=4.79
r221 (  47 91 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.56 //x2=4.145 //y2=1.405
r222 (  47 83 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.56 //x2=4.105 //y2=1.915
r223 (  46 91 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.25 //x2=4.145 //y2=1.405
r224 (  45 90 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=0.905 //x2=4.145 //y2=0.75
r225 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.105 //y=0.905 //x2=4.105 //y2=1.25
r226 (  44 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.22 //y=6.02 //x2=9.22 //y2=4.865
r227 (  43 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.78 //y=6.02 //x2=8.78 //y2=4.865
r228 (  42 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.55 //y=6.02 //x2=4.55 //y2=4.865
r229 (  41 89 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.11 //y=6.02 //x2=4.11 //y2=4.865
r230 (  40 73 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.365 //x2=9.06 //y2=1.365
r231 (  40 74 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.365 //x2=8.84 //y2=1.365
r232 (  39 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.37 //y=1.405 //x2=4.48 //y2=1.405
r233 (  39 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.37 //y=1.405 //x2=4.26 //y2=1.405
r234 (  38 86 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.1 //y=4.7 //x2=4.1 //y2=4.7
r235 (  35 100 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.88 //y=4.7 //x2=8.88 //y2=4.7
r236 (  27 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.88 //y=2.08 //x2=8.88 //y2=2.08
r237 (  18 82 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=2.08 //x2=4.07 //y2=2.08
r238 (  16 38 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=4.07 //y=4.535 //x2=4.085 //y2=4.7
r239 (  15 35 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=8.88 //y=4.44 //x2=8.88 //y2=4.7
r240 (  14 15 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=8.88 //y=3.33 //x2=8.88 //y2=4.44
r241 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=8.88 //y=2.96 //x2=8.88 //y2=3.33
r242 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=8.88 //y=2.59 //x2=8.88 //y2=2.96
r243 (  12 27 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=8.88 //y=2.59 //x2=8.88 //y2=2.08
r244 (  11 16 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=4.07 //y=4.44 //x2=4.07 //y2=4.535
r245 (  10 11 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=4.07 //y=3.7 //x2=4.07 //y2=4.44
r246 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=3.33 //x2=4.07 //y2=3.7
r247 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.07 //y=2.96 //x2=4.07 //y2=3.33
r248 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.07 //y=2.59 //x2=4.07 //y2=2.96
r249 (  7 18 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=4.07 //y=2.59 //x2=4.07 //y2=2.08
r250 (  6 13 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.88 //y=2.96 //x2=8.88 //y2=2.96
r251 (  4 8 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=4.07 \
 //y=2.96 //x2=4.07 //y2=2.96
r252 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=2.96 //x2=4.07 //y2=2.96
r253 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=2.96 //x2=8.88 //y2=2.96
r254 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=2.96 //x2=4.185 //y2=2.96
ends PM_DLATCH\%GATE

subckt PM_DLATCH\%D ( 1 2 7 8 9 10 11 12 13 14 15 16 17 18 19 21 34 36 47 48 \
 49 50 51 52 53 54 55 56 60 61 62 64 70 71 72 73 74 79 81 83 89 90 92 101 102 \
 105 )
c177 ( 105 0 ) capacitor c=0.0331844f //x=9.65 //y=4.7
c178 ( 102 0 ) capacitor c=0.0279499f //x=9.62 //y=1.915
c179 ( 101 0 ) capacitor c=0.0437302f //x=9.62 //y=2.08
c180 ( 92 0 ) capacitor c=0.0537799f //x=0.74 //y=2.085
c181 ( 90 0 ) capacitor c=0.0429696f //x=10.185 //y=1.25
c182 ( 89 0 ) capacitor c=0.0192208f //x=10.185 //y=0.905
c183 ( 83 0 ) capacitor c=0.0158629f //x=10.03 //y=1.405
c184 ( 81 0 ) capacitor c=0.0157803f //x=10.03 //y=0.75
c185 ( 79 0 ) capacitor c=0.0307199f //x=10.025 //y=4.79
c186 ( 74 0 ) capacitor c=0.0205163f //x=9.655 //y=1.56
c187 ( 73 0 ) capacitor c=0.0168481f //x=9.655 //y=1.25
c188 ( 72 0 ) capacitor c=0.0174783f //x=9.655 //y=0.905
c189 ( 71 0 ) capacitor c=0.0435629f //x=1.38 //y=1.255
c190 ( 70 0 ) capacitor c=0.0200386f //x=1.38 //y=0.91
c191 ( 64 0 ) capacitor c=0.0152946f //x=1.225 //y=1.41
c192 ( 62 0 ) capacitor c=0.0157804f //x=1.225 //y=0.755
c193 ( 61 0 ) capacitor c=0.048995f //x=0.97 //y=4.79
c194 ( 60 0 ) capacitor c=0.0303096f //x=1.26 //y=4.79
c195 ( 56 0 ) capacitor c=0.0290017f //x=0.85 //y=1.92
c196 ( 55 0 ) capacitor c=0.0250027f //x=0.85 //y=1.565
c197 ( 54 0 ) capacitor c=0.0234316f //x=0.85 //y=1.255
c198 ( 53 0 ) capacitor c=0.0200596f //x=0.85 //y=0.91
c199 ( 52 0 ) capacitor c=0.15358f //x=10.1 //y=6.02
c200 ( 51 0 ) capacitor c=0.110281f //x=9.66 //y=6.02
c201 ( 50 0 ) capacitor c=0.154218f //x=1.335 //y=6.02
c202 ( 49 0 ) capacitor c=0.154243f //x=0.895 //y=6.02
c203 ( 36 0 ) capacitor c=0.0762219f //x=9.62 //y=2.08
c204 ( 34 0 ) capacitor c=0.00453889f //x=9.62 //y=4.535
c205 ( 21 0 ) capacitor c=0.110709f //x=0.74 //y=2.085
c206 ( 2 0 ) capacitor c=0.0162171f //x=0.855 //y=4.07
c207 ( 1 0 ) capacitor c=0.257694f //x=9.505 //y=4.07
r208 (  107 108 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=9.65 //y=4.79 //x2=9.65 //y2=4.865
r209 (  105 107 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=9.65 //y=4.7 //x2=9.65 //y2=4.79
r210 (  101 102 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=9.62 //y=2.08 //x2=9.62 //y2=1.915
r211 (  92 93 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=0.74 //y=2.085 //x2=0.85 //y2=2.085
r212 (  90 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.185 //y=1.25 //x2=10.145 //y2=1.405
r213 (  89 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.185 //y=0.905 //x2=10.145 //y2=0.75
r214 (  89 90 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.185 //y=0.905 //x2=10.185 //y2=1.25
r215 (  84 110 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.81 //y=1.405 //x2=9.695 //y2=1.405
r216 (  83 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.03 //y=1.405 //x2=10.145 //y2=1.405
r217 (  82 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.81 //y=0.75 //x2=9.695 //y2=0.75
r218 (  81 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.03 //y=0.75 //x2=10.145 //y2=0.75
r219 (  81 82 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.03 //y=0.75 //x2=9.81 //y2=0.75
r220 (  80 107 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=9.785 //y=4.79 //x2=9.65 //y2=4.79
r221 (  79 86 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.025 //y=4.79 //x2=10.1 //y2=4.865
r222 (  79 80 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=10.025 //y=4.79 //x2=9.785 //y2=4.79
r223 (  74 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.655 //y=1.56 //x2=9.695 //y2=1.405
r224 (  74 102 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=9.655 //y=1.56 //x2=9.655 //y2=1.915
r225 (  73 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.655 //y=1.25 //x2=9.695 //y2=1.405
r226 (  72 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.655 //y=0.905 //x2=9.695 //y2=0.75
r227 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.655 //y=0.905 //x2=9.655 //y2=1.25
r228 (  71 99 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=1.255 //x2=1.34 //y2=1.41
r229 (  70 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.34 //y2=0.755
r230 (  70 71 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.38 //y2=1.255
r231 (  65 97 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=1.41 //x2=0.89 //y2=1.41
r232 (  64 99 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=1.41 //x2=1.34 //y2=1.41
r233 (  63 96 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=0.755 //x2=0.89 //y2=0.755
r234 (  62 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.34 //y2=0.755
r235 (  62 63 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.005 //y2=0.755
r236 (  60 67 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=1.335 //y2=4.865
r237 (  60 61 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=0.97 //y2=4.79
r238 (  57 61 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.97 //y2=4.79
r239 (  57 95 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.74 //y2=4.7
r240 (  56 93 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.92 //x2=0.85 //y2=2.085
r241 (  55 97 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.89 //y2=1.41
r242 (  55 56 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.85 //y2=1.92
r243 (  54 97 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.255 //x2=0.89 //y2=1.41
r244 (  53 96 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.89 //y2=0.755
r245 (  53 54 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.85 //y2=1.255
r246 (  52 86 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.1 //y=6.02 //x2=10.1 //y2=4.865
r247 (  51 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.66 //y=6.02 //x2=9.66 //y2=4.865
r248 (  50 67 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.335 //y=6.02 //x2=1.335 //y2=4.865
r249 (  49 57 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.895 //y=6.02 //x2=0.895 //y2=4.865
r250 (  48 83 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.92 //y=1.405 //x2=10.03 //y2=1.405
r251 (  48 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.92 //y=1.405 //x2=9.81 //y2=1.405
r252 (  47 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.225 //y2=1.41
r253 (  47 65 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.005 //y2=1.41
r254 (  46 105 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.65 //y=4.7 //x2=9.65 //y2=4.7
r255 (  36 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.62 //y=2.08 //x2=9.62 //y2=2.08
r256 (  34 46 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=9.62 //y=4.535 //x2=9.635 //y2=4.7
r257 (  32 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.7 //x2=0.74 //y2=4.7
r258 (  21 92 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=2.085
r259 (  19 34 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=9.62 //y=4.44 //x2=9.62 //y2=4.535
r260 (  18 19 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=9.62 //y=4.07 //x2=9.62 //y2=4.44
r261 (  17 18 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=9.62 //y=3.33 //x2=9.62 //y2=4.07
r262 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=9.62 //y=2.96 //x2=9.62 //y2=3.33
r263 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=9.62 //y=2.59 //x2=9.62 //y2=2.96
r264 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=9.62 //y=2.22 //x2=9.62 //y2=2.59
r265 (  14 36 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=9.62 //y=2.22 //x2=9.62 //y2=2.08
r266 (  13 32 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=0.74 //y=4.44 //x2=0.74 //y2=4.7
r267 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=4.07 //x2=0.74 //y2=4.44
r268 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=3.7 //x2=0.74 //y2=4.07
r269 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=3.33 //x2=0.74 //y2=3.7
r270 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=2.96 //x2=0.74 //y2=3.33
r271 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.59 //x2=0.74 //y2=2.96
r272 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.22 //x2=0.74 //y2=2.59
r273 (  7 21 ) resistor r=9.24064 //w=0.187 //l=0.135 //layer=li \
 //thickness=0.1 //x=0.74 //y=2.22 //x2=0.74 //y2=2.085
r274 (  6 18 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.62 //y=4.07 //x2=9.62 //y2=4.07
r275 (  4 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=0.74 //y=4.07 //x2=0.74 //y2=4.07
r276 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=0.855 //y=4.07 //x2=0.74 //y2=4.07
r277 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=4.07 //x2=9.62 //y2=4.07
r278 (  1 2 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=4.07 //x2=0.855 //y2=4.07
ends PM_DLATCH\%D

subckt PM_DLATCH\%noxref_7 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 \
 52 53 54 56 62 63 65 73 75 76 )
c139 ( 76 0 ) capacitor c=0.0220291f //x=9.735 //y=5.02
c140 ( 75 0 ) capacitor c=0.0217503f //x=8.855 //y=5.02
c141 ( 73 0 ) capacitor c=0.0084702f //x=9.73 //y=0.905
c142 ( 65 0 ) capacitor c=0.0528806f //x=11.84 //y=2.085
c143 ( 63 0 ) capacitor c=0.0435629f //x=12.48 //y=1.255
c144 ( 62 0 ) capacitor c=0.0200386f //x=12.48 //y=0.91
c145 ( 56 0 ) capacitor c=0.0152946f //x=12.325 //y=1.41
c146 ( 54 0 ) capacitor c=0.0157804f //x=12.325 //y=0.755
c147 ( 53 0 ) capacitor c=0.0493989f //x=12.07 //y=4.79
c148 ( 52 0 ) capacitor c=0.0304843f //x=12.36 //y=4.79
c149 ( 48 0 ) capacitor c=0.0290017f //x=11.95 //y=1.92
c150 ( 47 0 ) capacitor c=0.0250027f //x=11.95 //y=1.565
c151 ( 46 0 ) capacitor c=0.0234316f //x=11.95 //y=1.255
c152 ( 45 0 ) capacitor c=0.0200596f //x=11.95 //y=0.91
c153 ( 44 0 ) capacitor c=0.154218f //x=12.435 //y=6.02
c154 ( 43 0 ) capacitor c=0.154243f //x=11.995 //y=6.02
c155 ( 41 0 ) capacitor c=0.0024826f //x=9.88 //y=5.2
c156 ( 34 0 ) capacitor c=0.0908493f //x=11.84 //y=2.085
c157 ( 32 0 ) capacitor c=0.108527f //x=10.36 //y=3.33
c158 ( 28 0 ) capacitor c=0.00525782f //x=10.005 //y=1.655
c159 ( 27 0 ) capacitor c=0.0139525f //x=10.275 //y=1.655
c160 ( 25 0 ) capacitor c=0.0144648f //x=10.275 //y=5.2
c161 ( 14 0 ) capacitor c=0.00265825f //x=9.085 //y=5.2
c162 ( 13 0 ) capacitor c=0.0150834f //x=9.795 //y=5.2
c163 ( 2 0 ) capacitor c=0.0111324f //x=10.475 //y=3.33
c164 ( 1 0 ) capacitor c=0.0522233f //x=11.725 //y=3.33
r165 (  65 66 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.84 //y=2.085 //x2=11.95 //y2=2.085
r166 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.48 //y=1.255 //x2=12.44 //y2=1.41
r167 (  62 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.48 //y=0.91 //x2=12.44 //y2=0.755
r168 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.48 //y=0.91 //x2=12.48 //y2=1.255
r169 (  57 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.105 //y=1.41 //x2=11.99 //y2=1.41
r170 (  56 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.325 //y=1.41 //x2=12.44 //y2=1.41
r171 (  55 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.105 //y=0.755 //x2=11.99 //y2=0.755
r172 (  54 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.325 //y=0.755 //x2=12.44 //y2=0.755
r173 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=12.325 //y=0.755 //x2=12.105 //y2=0.755
r174 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=12.36 //y=4.79 //x2=12.435 //y2=4.865
r175 (  52 53 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=12.36 //y=4.79 //x2=12.07 //y2=4.79
r176 (  49 53 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.995 //y=4.865 //x2=12.07 //y2=4.79
r177 (  49 68 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=11.995 //y=4.865 //x2=11.84 //y2=4.7
r178 (  48 66 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11.95 //y=1.92 //x2=11.95 //y2=2.085
r179 (  47 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.95 //y=1.565 //x2=11.99 //y2=1.41
r180 (  47 48 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=11.95 //y=1.565 //x2=11.95 //y2=1.92
r181 (  46 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.95 //y=1.255 //x2=11.99 //y2=1.41
r182 (  45 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.95 //y=0.91 //x2=11.99 //y2=0.755
r183 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.95 //y=0.91 //x2=11.95 //y2=1.255
r184 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.435 //y=6.02 //x2=12.435 //y2=4.865
r185 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.995 //y=6.02 //x2=11.995 //y2=4.865
r186 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.215 //y=1.41 //x2=12.325 //y2=1.41
r187 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.215 //y=1.41 //x2=12.105 //y2=1.41
r188 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=4.7 //x2=11.84 //y2=4.7
r189 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=11.84 //y=3.33 //x2=11.84 //y2=4.7
r190 (  34 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=2.085 //x2=11.84 //y2=2.085
r191 (  34 37 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.085 //x2=11.84 //y2=3.33
r192 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=10.36 //y=5.115 //x2=10.36 //y2=3.33
r193 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=10.36 //y=1.74 //x2=10.36 //y2=3.33
r194 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.275 //y=1.655 //x2=10.36 //y2=1.74
r195 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=10.275 //y=1.655 //x2=10.005 //y2=1.655
r196 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.965 //y=5.2 //x2=9.88 //y2=5.2
r197 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.275 //y=5.2 //x2=10.36 //y2=5.115
r198 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=10.275 //y=5.2 //x2=9.965 //y2=5.2
r199 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.92 //y=1.57 //x2=10.005 //y2=1.655
r200 (  21 73 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.92 //y=1.57 //x2=9.92 //y2=1
r201 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.88 //y=5.285 //x2=9.88 //y2=5.2
r202 (  15 76 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=9.88 //y=5.285 //x2=9.88 //y2=5.725
r203 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.795 //y=5.2 //x2=9.88 //y2=5.2
r204 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=9.795 //y=5.2 //x2=9.085 //y2=5.2
r205 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9 //y=5.285 //x2=9.085 //y2=5.2
r206 (  7 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=9 //y=5.285 //x2=9 //y2=5.725
r207 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.84 //y=3.33 //x2=11.84 //y2=3.33
r208 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=3.33 //x2=10.36 //y2=3.33
r209 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.475 //y=3.33 //x2=10.36 //y2=3.33
r210 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.725 //y=3.33 //x2=11.84 //y2=3.33
r211 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=11.725 //y=3.33 //x2=10.475 //y2=3.33
ends PM_DLATCH\%noxref_7

subckt PM_DLATCH\%noxref_8 ( 1 2 17 18 19 20 24 27 32 34 35 36 37 38 39 40 44 \
 46 49 51 52 57 67 69 )
c164 ( 69 0 ) capacitor c=0.0288745f //x=6.52 //y=5.02
c165 ( 67 0 ) capacitor c=0.0173218f //x=6.475 //y=0.91
c166 ( 57 0 ) capacitor c=0.0403405f //x=14.275 //y=4.705
c167 ( 52 0 ) capacitor c=0.0321911f //x=14.765 //y=1.25
c168 ( 51 0 ) capacitor c=0.0185201f //x=14.765 //y=0.905
c169 ( 49 0 ) capacitor c=0.0288104f //x=14.695 //y=4.795
c170 ( 46 0 ) capacitor c=0.0133656f //x=14.61 //y=1.405
c171 ( 44 0 ) capacitor c=0.0157804f //x=14.61 //y=0.75
c172 ( 40 0 ) capacitor c=0.0828832f //x=14.235 //y=1.915
c173 ( 39 0 ) capacitor c=0.022867f //x=14.235 //y=1.56
c174 ( 38 0 ) capacitor c=0.0234318f //x=14.235 //y=1.25
c175 ( 37 0 ) capacitor c=0.0192004f //x=14.235 //y=0.905
c176 ( 36 0 ) capacitor c=0.110795f //x=14.77 //y=6.025
c177 ( 35 0 ) capacitor c=0.153847f //x=14.33 //y=6.025
c178 ( 32 0 ) capacitor c=0.00993392f //x=14.275 //y=4.705
c179 ( 27 0 ) capacitor c=0.0921227f //x=14.43 //y=2.08
c180 ( 24 0 ) capacitor c=0.0820607f //x=7.03 //y=3.7
c181 ( 20 0 ) capacitor c=0.00417404f //x=6.75 //y=4.58
c182 ( 19 0 ) capacitor c=0.0118896f //x=6.945 //y=4.58
c183 ( 18 0 ) capacitor c=0.00549299f //x=6.745 //y=2.08
c184 ( 17 0 ) capacitor c=0.013178f //x=6.945 //y=2.08
c185 ( 2 0 ) capacitor c=0.0108199f //x=7.145 //y=3.7
c186 ( 1 0 ) capacitor c=0.214055f //x=14.315 //y=3.7
r187 (  59 60 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=14.275 //y=4.795 //x2=14.275 //y2=4.87
r188 (  57 59 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=14.275 //y=4.705 //x2=14.275 //y2=4.795
r189 (  52 66 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.765 //y=1.25 //x2=14.725 //y2=1.405
r190 (  51 65 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.765 //y=0.905 //x2=14.725 //y2=0.75
r191 (  51 52 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.765 //y=0.905 //x2=14.765 //y2=1.25
r192 (  50 59 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=14.41 //y=4.795 //x2=14.275 //y2=4.795
r193 (  49 53 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=14.695 //y=4.795 //x2=14.77 //y2=4.87
r194 (  49 50 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=14.695 //y=4.795 //x2=14.41 //y2=4.795
r195 (  47 64 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.39 //y=1.405 //x2=14.275 //y2=1.405
r196 (  46 66 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.61 //y=1.405 //x2=14.725 //y2=1.405
r197 (  45 63 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.39 //y=0.75 //x2=14.275 //y2=0.75
r198 (  44 65 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.61 //y=0.75 //x2=14.725 //y2=0.75
r199 (  44 45 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=14.61 //y=0.75 //x2=14.39 //y2=0.75
r200 (  40 62 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=14.235 //y=1.915 //x2=14.43 //y2=2.08
r201 (  39 64 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.235 //y=1.56 //x2=14.275 //y2=1.405
r202 (  39 40 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=14.235 //y=1.56 //x2=14.235 //y2=1.915
r203 (  38 64 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.235 //y=1.25 //x2=14.275 //y2=1.405
r204 (  37 63 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.235 //y=0.905 //x2=14.275 //y2=0.75
r205 (  37 38 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.235 //y=0.905 //x2=14.235 //y2=1.25
r206 (  36 53 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.77 //y=6.025 //x2=14.77 //y2=4.87
r207 (  35 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.33 //y=6.025 //x2=14.33 //y2=4.87
r208 (  34 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.5 //y=1.405 //x2=14.61 //y2=1.405
r209 (  34 47 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.5 //y=1.405 //x2=14.39 //y2=1.405
r210 (  32 57 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.275 //y=4.705 //x2=14.275 //y2=4.705
r211 (  32 33 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=14.275 //y=4.705 //x2=14.43 //y2=4.705
r212 (  27 62 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.43 //y=2.08 //x2=14.43 //y2=2.08
r213 (  27 30 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=14.43 //y=2.08 //x2=14.43 //y2=3.7
r214 (  25 33 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=14.43 //y=4.54 //x2=14.43 //y2=4.705
r215 (  25 30 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=14.43 //y=4.54 //x2=14.43 //y2=3.7
r216 (  22 24 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=7.03 //y=4.495 //x2=7.03 //y2=3.7
r217 (  21 24 ) resistor r=105.07 //w=0.187 //l=1.535 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.165 //x2=7.03 //y2=3.7
r218 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.945 //y=4.58 //x2=7.03 //y2=4.495
r219 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=6.945 //y=4.58 //x2=6.75 //y2=4.58
r220 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.945 //y=2.08 //x2=7.03 //y2=2.165
r221 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=6.945 //y=2.08 //x2=6.745 //y2=2.08
r222 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.665 //y=4.665 //x2=6.75 //y2=4.58
r223 (  11 69 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=6.665 //y=4.665 //x2=6.665 //y2=5.725
r224 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.66 //y=1.995 //x2=6.745 //y2=2.08
r225 (  7 67 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=6.66 //y=1.995 //x2=6.66 //y2=1.005
r226 (  6 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.43 //y=3.7 //x2=14.43 //y2=3.7
r227 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.03 //y=3.7 //x2=7.03 //y2=3.7
r228 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.145 //y=3.7 //x2=7.03 //y2=3.7
r229 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.315 //y=3.7 //x2=14.43 //y2=3.7
r230 (  1 2 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=14.315 //y=3.7 //x2=7.145 //y2=3.7
ends PM_DLATCH\%noxref_8

subckt PM_DLATCH\%Q ( 1 2 7 8 9 10 11 12 13 14 15 16 21 22 33 34 35 47 57 59 \
 60 61 62 63 64 65 69 71 74 76 77 82 92 93 96 )
c167 ( 96 0 ) capacitor c=0.0159573f //x=15.285 //y=5.025
c168 ( 93 0 ) capacitor c=0.00923651f //x=15.28 //y=0.905
c169 ( 92 0 ) capacitor c=0.007684f //x=14.31 //y=0.905
c170 ( 82 0 ) capacitor c=0.0402699f //x=17.605 //y=4.705
c171 ( 77 0 ) capacitor c=0.0321911f //x=18.095 //y=1.25
c172 ( 76 0 ) capacitor c=0.0185201f //x=18.095 //y=0.905
c173 ( 74 0 ) capacitor c=0.0288104f //x=18.025 //y=4.795
c174 ( 71 0 ) capacitor c=0.0133656f //x=17.94 //y=1.405
c175 ( 69 0 ) capacitor c=0.0157804f //x=17.94 //y=0.75
c176 ( 65 0 ) capacitor c=0.0822075f //x=17.565 //y=1.915
c177 ( 64 0 ) capacitor c=0.022867f //x=17.565 //y=1.56
c178 ( 63 0 ) capacitor c=0.0234318f //x=17.565 //y=1.25
c179 ( 62 0 ) capacitor c=0.0192004f //x=17.565 //y=0.905
c180 ( 61 0 ) capacitor c=0.110795f //x=18.1 //y=6.025
c181 ( 60 0 ) capacitor c=0.153847f //x=17.66 //y=6.025
c182 ( 57 0 ) capacitor c=0.00993392f //x=17.605 //y=4.705
c183 ( 55 0 ) capacitor c=0.00454201f //x=15.47 //y=1.655
c184 ( 47 0 ) capacitor c=0.0893171f //x=17.76 //y=2.08
c185 ( 35 0 ) capacitor c=0.0140918f //x=15.825 //y=1.655
c186 ( 34 0 ) capacitor c=0.00308317f //x=15.515 //y=5.21
c187 ( 33 0 ) capacitor c=0.0137261f //x=15.825 //y=5.21
c188 ( 22 0 ) capacitor c=0.00224268f //x=14.585 //y=1.655
c189 ( 21 0 ) capacitor c=0.0218623f //x=15.385 //y=1.655
c190 ( 7 0 ) capacitor c=0.110461f //x=15.91 //y=2.22
c191 ( 2 0 ) capacitor c=0.0112178f //x=16.025 //y=3.33
c192 ( 1 0 ) capacitor c=0.0678125f //x=17.645 //y=3.33
r193 (  84 85 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=17.605 //y=4.795 //x2=17.605 //y2=4.87
r194 (  82 84 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=17.605 //y=4.705 //x2=17.605 //y2=4.795
r195 (  77 91 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.095 //y=1.25 //x2=18.055 //y2=1.405
r196 (  76 90 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.095 //y=0.905 //x2=18.055 //y2=0.75
r197 (  76 77 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.095 //y=0.905 //x2=18.095 //y2=1.25
r198 (  75 84 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=17.74 //y=4.795 //x2=17.605 //y2=4.795
r199 (  74 78 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=18.025 //y=4.795 //x2=18.1 //y2=4.87
r200 (  74 75 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=18.025 //y=4.795 //x2=17.74 //y2=4.795
r201 (  72 89 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.72 //y=1.405 //x2=17.605 //y2=1.405
r202 (  71 91 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.94 //y=1.405 //x2=18.055 //y2=1.405
r203 (  70 88 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.72 //y=0.75 //x2=17.605 //y2=0.75
r204 (  69 90 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.94 //y=0.75 //x2=18.055 //y2=0.75
r205 (  69 70 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.94 //y=0.75 //x2=17.72 //y2=0.75
r206 (  65 87 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=17.565 //y=1.915 //x2=17.76 //y2=2.08
r207 (  64 89 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.565 //y=1.56 //x2=17.605 //y2=1.405
r208 (  64 65 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=17.565 //y=1.56 //x2=17.565 //y2=1.915
r209 (  63 89 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.565 //y=1.25 //x2=17.605 //y2=1.405
r210 (  62 88 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.565 //y=0.905 //x2=17.605 //y2=0.75
r211 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.565 //y=0.905 //x2=17.565 //y2=1.25
r212 (  61 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.1 //y=6.025 //x2=18.1 //y2=4.87
r213 (  60 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.66 //y=6.025 //x2=17.66 //y2=4.87
r214 (  59 71 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.83 //y=1.405 //x2=17.94 //y2=1.405
r215 (  59 72 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.83 //y=1.405 //x2=17.72 //y2=1.405
r216 (  57 82 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.605 //y=4.705 //x2=17.605 //y2=4.705
r217 (  57 58 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=17.605 //y=4.705 //x2=17.76 //y2=4.705
r218 (  47 87 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=2.08 //x2=17.76 //y2=2.08
r219 (  45 58 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=17.76 //y=4.54 //x2=17.76 //y2=4.705
r220 (  36 55 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.555 //y=1.655 //x2=15.47 //y2=1.655
r221 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.825 //y=1.655 //x2=15.91 //y2=1.74
r222 (  35 36 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=15.825 //y=1.655 //x2=15.555 //y2=1.655
r223 (  33 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.825 //y=5.21 //x2=15.91 //y2=5.125
r224 (  33 34 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=15.825 //y=5.21 //x2=15.515 //y2=5.21
r225 (  29 55 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.47 //y=1.57 //x2=15.47 //y2=1.655
r226 (  29 93 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=15.47 //y=1.57 //x2=15.47 //y2=1
r227 (  23 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.43 //y=5.295 //x2=15.515 //y2=5.21
r228 (  23 96 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=15.43 //y=5.295 //x2=15.43 //y2=5.72
r229 (  21 55 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.385 //y=1.655 //x2=15.47 //y2=1.655
r230 (  21 22 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=15.385 //y=1.655 //x2=14.585 //y2=1.655
r231 (  17 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.5 //y=1.57 //x2=14.585 //y2=1.655
r232 (  17 92 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.5 //y=1.57 //x2=14.5 //y2=1
r233 (  16 45 ) resistor r=6.84492 //w=0.187 //l=0.1 //layer=li \
 //thickness=0.1 //x=17.76 //y=4.44 //x2=17.76 //y2=4.54
r234 (  15 16 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.76 //y=3.33 //x2=17.76 //y2=4.44
r235 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.96 //x2=17.76 //y2=3.33
r236 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.59 //x2=17.76 //y2=2.96
r237 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.22 //x2=17.76 //y2=2.59
r238 (  12 47 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.22 //x2=17.76 //y2=2.08
r239 (  11 38 ) resistor r=46.8877 //w=0.187 //l=0.685 //layer=li \
 //thickness=0.1 //x=15.91 //y=4.44 //x2=15.91 //y2=5.125
r240 (  10 11 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=15.91 //y=3.33 //x2=15.91 //y2=4.44
r241 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.91 //y=2.96 //x2=15.91 //y2=3.33
r242 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=15.91 //y=2.59 //x2=15.91 //y2=2.96
r243 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=15.91 //y=2.22 //x2=15.91 //y2=2.59
r244 (  7 37 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li \
 //thickness=0.1 //x=15.91 //y=2.22 //x2=15.91 //y2=1.74
r245 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.76 //y=3.33 //x2=17.76 //y2=3.33
r246 (  4 10 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.91 //y=3.33 //x2=15.91 //y2=3.33
r247 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.025 //y=3.33 //x2=15.91 //y2=3.33
r248 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.645 //y=3.33 //x2=17.76 //y2=3.33
r249 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=17.645 //y=3.33 //x2=16.025 //y2=3.33
ends PM_DLATCH\%Q

subckt PM_DLATCH\%noxref_10 ( 1 2 17 18 19 20 24 25 27 33 34 35 36 37 38 43 45 \
 47 53 54 56 57 60 68 70 )
c162 ( 70 0 ) capacitor c=0.028853f //x=12.07 //y=5.02
c163 ( 68 0 ) capacitor c=0.0173218f //x=12.025 //y=0.91
c164 ( 60 0 ) capacitor c=0.0354945f //x=18.535 //y=4.705
c165 ( 57 0 ) capacitor c=0.0279572f //x=18.5 //y=1.915
c166 ( 56 0 ) capacitor c=0.0422144f //x=18.5 //y=2.08
c167 ( 54 0 ) capacitor c=0.0237734f //x=19.065 //y=1.255
c168 ( 53 0 ) capacitor c=0.0191782f //x=19.065 //y=0.905
c169 ( 47 0 ) capacitor c=0.0346941f //x=18.91 //y=1.405
c170 ( 45 0 ) capacitor c=0.0157803f //x=18.91 //y=0.75
c171 ( 43 0 ) capacitor c=0.030194f //x=18.905 //y=4.795
c172 ( 38 0 ) capacitor c=0.0199921f //x=18.535 //y=1.56
c173 ( 37 0 ) capacitor c=0.0169608f //x=18.535 //y=1.255
c174 ( 36 0 ) capacitor c=0.0185462f //x=18.535 //y=0.905
c175 ( 35 0 ) capacitor c=0.15325f //x=18.98 //y=6.025
c176 ( 34 0 ) capacitor c=0.110232f //x=18.54 //y=6.025
c177 ( 27 0 ) capacitor c=0.0760752f //x=18.5 //y=2.08
c178 ( 25 0 ) capacitor c=0.00514985f //x=18.5 //y=4.54
c179 ( 24 0 ) capacitor c=0.0855616f //x=12.58 //y=4.07
c180 ( 20 0 ) capacitor c=0.00497659f //x=12.3 //y=4.58
c181 ( 19 0 ) capacitor c=0.012509f //x=12.495 //y=4.58
c182 ( 18 0 ) capacitor c=0.00612032f //x=12.295 //y=2.08
c183 ( 17 0 ) capacitor c=0.0138937f //x=12.495 //y=2.08
c184 ( 2 0 ) capacitor c=0.0119148f //x=12.695 //y=4.07
c185 ( 1 0 ) capacitor c=0.169542f //x=18.385 //y=4.07
r186 (  62 63 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.795 //x2=18.535 //y2=4.87
r187 (  60 62 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.705 //x2=18.535 //y2=4.795
r188 (  56 57 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=18.5 //y=2.08 //x2=18.5 //y2=1.915
r189 (  54 67 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=19.065 //y=1.255 //x2=19.065 //y2=1.367
r190 (  53 66 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.065 //y=0.905 //x2=19.025 //y2=0.75
r191 (  53 54 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=19.065 //y=0.905 //x2=19.065 //y2=1.255
r192 (  48 65 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.69 //y=1.405 //x2=18.575 //y2=1.405
r193 (  47 67 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=18.91 //y=1.405 //x2=19.065 //y2=1.367
r194 (  46 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.69 //y=0.75 //x2=18.575 //y2=0.75
r195 (  45 66 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.91 //y=0.75 //x2=19.025 //y2=0.75
r196 (  45 46 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.91 //y=0.75 //x2=18.69 //y2=0.75
r197 (  44 62 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=18.67 //y=4.795 //x2=18.535 //y2=4.795
r198 (  43 50 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=18.905 //y=4.795 //x2=18.98 //y2=4.87
r199 (  43 44 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=18.905 //y=4.795 //x2=18.67 //y2=4.795
r200 (  38 65 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.535 //y=1.56 //x2=18.575 //y2=1.405
r201 (  38 57 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=18.535 //y=1.56 //x2=18.535 //y2=1.915
r202 (  37 65 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=18.535 //y=1.255 //x2=18.575 //y2=1.405
r203 (  36 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.535 //y=0.905 //x2=18.575 //y2=0.75
r204 (  36 37 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=18.535 //y=0.905 //x2=18.535 //y2=1.255
r205 (  35 50 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.98 //y=6.025 //x2=18.98 //y2=4.87
r206 (  34 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.54 //y=6.025 //x2=18.54 //y2=4.87
r207 (  33 47 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.8 //y=1.405 //x2=18.91 //y2=1.405
r208 (  33 48 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.8 //y=1.405 //x2=18.69 //y2=1.405
r209 (  32 60 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.535 //y=4.705 //x2=18.535 //y2=4.705
r210 (  27 56 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.5 //y=2.08 //x2=18.5 //y2=2.08
r211 (  27 30 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=18.5 //y=2.08 //x2=18.5 //y2=4.07
r212 (  25 32 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=18.5 //y=4.54 //x2=18.517 //y2=4.705
r213 (  25 30 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=18.5 //y=4.54 //x2=18.5 //y2=4.07
r214 (  22 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=12.58 //y=4.495 //x2=12.58 //y2=4.07
r215 (  21 24 ) resistor r=130.396 //w=0.187 //l=1.905 //layer=li \
 //thickness=0.1 //x=12.58 //y=2.165 //x2=12.58 //y2=4.07
r216 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.495 //y=4.58 //x2=12.58 //y2=4.495
r217 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=12.495 //y=4.58 //x2=12.3 //y2=4.58
r218 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.495 //y=2.08 //x2=12.58 //y2=2.165
r219 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.495 //y=2.08 //x2=12.295 //y2=2.08
r220 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.215 //y=4.665 //x2=12.3 //y2=4.58
r221 (  11 70 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=12.215 //y=4.665 //x2=12.215 //y2=5.725
r222 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.995 //x2=12.295 //y2=2.08
r223 (  7 68 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.995 //x2=12.21 //y2=1.005
r224 (  6 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.5 //y=4.07 //x2=18.5 //y2=4.07
r225 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.58 //y=4.07 //x2=12.58 //y2=4.07
r226 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.695 //y=4.07 //x2=12.58 //y2=4.07
r227 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=4.07 //x2=18.5 //y2=4.07
r228 (  1 2 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=4.07 //x2=12.695 //y2=4.07
ends PM_DLATCH\%noxref_10

subckt PM_DLATCH\%noxref_11 ( 1 2 7 9 17 18 29 30 31 36 40 41 42 43 44 45 50 \
 52 54 60 61 63 64 67 75 76 79 )
c162 ( 79 0 ) capacitor c=0.0159573f //x=18.615 //y=5.025
c163 ( 76 0 ) capacitor c=0.00905936f //x=18.61 //y=0.905
c164 ( 75 0 ) capacitor c=0.007684f //x=17.64 //y=0.905
c165 ( 67 0 ) capacitor c=0.0354569f //x=15.205 //y=4.705
c166 ( 64 0 ) capacitor c=0.0279572f //x=15.17 //y=1.915
c167 ( 63 0 ) capacitor c=0.0422144f //x=15.17 //y=2.08
c168 ( 61 0 ) capacitor c=0.0237734f //x=15.735 //y=1.255
c169 ( 60 0 ) capacitor c=0.0191782f //x=15.735 //y=0.905
c170 ( 54 0 ) capacitor c=0.0346941f //x=15.58 //y=1.405
c171 ( 52 0 ) capacitor c=0.0157803f //x=15.58 //y=0.75
c172 ( 50 0 ) capacitor c=0.0295389f //x=15.575 //y=4.795
c173 ( 45 0 ) capacitor c=0.0199921f //x=15.205 //y=1.56
c174 ( 44 0 ) capacitor c=0.0169608f //x=15.205 //y=1.255
c175 ( 43 0 ) capacitor c=0.0185462f //x=15.205 //y=0.905
c176 ( 42 0 ) capacitor c=0.15325f //x=15.65 //y=6.025
c177 ( 41 0 ) capacitor c=0.110232f //x=15.21 //y=6.025
c178 ( 39 0 ) capacitor c=0.00454201f //x=18.8 //y=1.655
c179 ( 36 0 ) capacitor c=0.128643f //x=19.24 //y=3.7
c180 ( 31 0 ) capacitor c=0.0141769f //x=19.155 //y=1.655
c181 ( 30 0 ) capacitor c=0.00326058f //x=18.845 //y=5.21
c182 ( 29 0 ) capacitor c=0.014f //x=19.155 //y=5.21
c183 ( 18 0 ) capacitor c=0.00217843f //x=17.915 //y=1.655
c184 ( 17 0 ) capacitor c=0.0212471f //x=18.715 //y=1.655
c185 ( 9 0 ) capacitor c=0.0762833f //x=15.17 //y=2.08
c186 ( 7 0 ) capacitor c=0.00514991f //x=15.17 //y=4.54
c187 ( 2 0 ) capacitor c=0.00669602f //x=15.285 //y=3.7
c188 ( 1 0 ) capacitor c=0.100901f //x=19.125 //y=3.7
r189 (  69 70 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.795 //x2=15.205 //y2=4.87
r190 (  67 69 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.705 //x2=15.205 //y2=4.795
r191 (  63 64 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=15.17 //y=2.08 //x2=15.17 //y2=1.915
r192 (  61 74 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=15.735 //y=1.255 //x2=15.735 //y2=1.367
r193 (  60 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.735 //y=0.905 //x2=15.695 //y2=0.75
r194 (  60 61 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=15.735 //y=0.905 //x2=15.735 //y2=1.255
r195 (  55 72 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.36 //y=1.405 //x2=15.245 //y2=1.405
r196 (  54 74 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=15.58 //y=1.405 //x2=15.735 //y2=1.367
r197 (  53 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.36 //y=0.75 //x2=15.245 //y2=0.75
r198 (  52 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.58 //y=0.75 //x2=15.695 //y2=0.75
r199 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.58 //y=0.75 //x2=15.36 //y2=0.75
r200 (  51 69 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=15.34 //y=4.795 //x2=15.205 //y2=4.795
r201 (  50 57 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.575 //y=4.795 //x2=15.65 //y2=4.87
r202 (  50 51 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=15.575 //y=4.795 //x2=15.34 //y2=4.795
r203 (  45 72 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.205 //y=1.56 //x2=15.245 //y2=1.405
r204 (  45 64 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=15.205 //y=1.56 //x2=15.205 //y2=1.915
r205 (  44 72 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=15.205 //y=1.255 //x2=15.245 //y2=1.405
r206 (  43 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.205 //y=0.905 //x2=15.245 //y2=0.75
r207 (  43 44 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=15.205 //y=0.905 //x2=15.205 //y2=1.255
r208 (  42 57 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.65 //y=6.025 //x2=15.65 //y2=4.87
r209 (  41 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.21 //y=6.025 //x2=15.21 //y2=4.87
r210 (  40 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.47 //y=1.405 //x2=15.58 //y2=1.405
r211 (  40 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.47 //y=1.405 //x2=15.36 //y2=1.405
r212 (  38 67 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.205 //y=4.705 //x2=15.205 //y2=4.705
r213 (  34 36 ) resistor r=97.5401 //w=0.187 //l=1.425 //layer=li \
 //thickness=0.1 //x=19.24 //y=5.125 //x2=19.24 //y2=3.7
r214 (  33 36 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=19.24 //y=1.74 //x2=19.24 //y2=3.7
r215 (  32 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.885 //y=1.655 //x2=18.8 //y2=1.655
r216 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.155 //y=1.655 //x2=19.24 //y2=1.74
r217 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=19.155 //y=1.655 //x2=18.885 //y2=1.655
r218 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.155 //y=5.21 //x2=19.24 //y2=5.125
r219 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=19.155 //y=5.21 //x2=18.845 //y2=5.21
r220 (  25 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.8 //y=1.57 //x2=18.8 //y2=1.655
r221 (  25 76 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=18.8 //y=1.57 //x2=18.8 //y2=1
r222 (  19 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.76 //y=5.295 //x2=18.845 //y2=5.21
r223 (  19 79 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=18.76 //y=5.295 //x2=18.76 //y2=5.72
r224 (  17 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.715 //y=1.655 //x2=18.8 //y2=1.655
r225 (  17 18 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=18.715 //y=1.655 //x2=17.915 //y2=1.655
r226 (  13 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.83 //y=1.57 //x2=17.915 //y2=1.655
r227 (  13 75 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=17.83 //y=1.57 //x2=17.83 //y2=1
r228 (  9 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.17 //y=2.08 //x2=15.17 //y2=2.08
r229 (  9 12 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=15.17 //y=2.08 //x2=15.17 //y2=3.7
r230 (  7 38 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=15.17 //y=4.54 //x2=15.187 //y2=4.705
r231 (  7 12 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=15.17 //y=4.54 //x2=15.17 //y2=3.7
r232 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.24 //y=3.7 //x2=19.24 //y2=3.7
r233 (  4 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.17 //y=3.7 //x2=15.17 //y2=3.7
r234 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.285 //y=3.7 //x2=15.17 //y2=3.7
r235 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.125 //y=3.7 //x2=19.24 //y2=3.7
r236 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=19.125 //y=3.7 //x2=15.285 //y2=3.7
ends PM_DLATCH\%noxref_11

subckt PM_DLATCH\%noxref_12 ( 1 5 9 10 13 17 29 )
c55 ( 29 0 ) capacitor c=0.0631306f //x=2.78 //y=0.365
c56 ( 17 0 ) capacitor c=0.00722223f //x=4.855 //y=0.615
c57 ( 13 0 ) capacitor c=0.0149611f //x=4.77 //y=0.53
c58 ( 10 0 ) capacitor c=0.00698743f //x=3.885 //y=1.495
c59 ( 9 0 ) capacitor c=0.006761f //x=3.885 //y=0.615
c60 ( 5 0 ) capacitor c=0.0207245f //x=3.8 //y=1.58
c61 ( 1 0 ) capacitor c=0.00856252f //x=2.915 //y=1.495
r62 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.855 //y=0.615 //x2=4.855 //y2=0.49
r63 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.855 //y=0.615 //x2=4.855 //y2=0.88
r64 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.97 //y=0.53 //x2=3.885 //y2=0.49
r65 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.97 //y=0.53 //x2=4.37 //y2=0.53
r66 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.77 //y=0.53 //x2=4.855 //y2=0.49
r67 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.77 //y=0.53 //x2=4.37 //y2=0.53
r68 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=3.885 //y=1.495 //x2=3.885 //y2=1.62
r69 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=3.885 //y=1.495 //x2=3.885 //y2=0.88
r70 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.885 //y=0.615 //x2=3.885 //y2=0.49
r71 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.885 //y=0.615 //x2=3.885 //y2=0.88
r72 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3 //y=1.58 //x2=2.915 //y2=1.62
r73 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3 //y=1.58 //x2=3.4 //y2=1.58
r74 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.8 //y=1.58 //x2=3.885 //y2=1.62
r75 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.8 //y=1.58 //x2=3.4 //y2=1.58
r76 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=2.915 //y=1.495 //x2=2.915 //y2=1.62
r77 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.915 //y=1.495 //x2=2.915 //y2=0.88
ends PM_DLATCH\%noxref_12

subckt PM_DLATCH\%noxref_13 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0633899f //x=8.33 //y=0.365
c55 ( 17 0 ) capacitor c=0.00722223f //x=10.405 //y=0.615
c56 ( 13 0 ) capacitor c=0.0149613f //x=10.32 //y=0.53
c57 ( 10 0 ) capacitor c=0.00687696f //x=9.435 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=9.435 //y=0.615
c59 ( 5 0 ) capacitor c=0.0199444f //x=9.35 //y=1.58
c60 ( 1 0 ) capacitor c=0.00798521f //x=8.465 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=10.405 //y=0.615 //x2=10.405 //y2=0.49
r62 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=10.405 //y=0.615 //x2=10.405 //y2=0.88
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.52 //y=0.53 //x2=9.435 //y2=0.49
r64 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.52 //y=0.53 //x2=9.92 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.32 //y=0.53 //x2=10.405 //y2=0.49
r66 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.32 //y=0.53 //x2=9.92 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.435 //y=1.495 //x2=9.435 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.435 //y=1.495 //x2=9.435 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.435 //y=0.615 //x2=9.435 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=9.435 //y=0.615 //x2=9.435 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.55 //y=1.58 //x2=8.465 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.55 //y=1.58 //x2=8.95 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.35 //y=1.58 //x2=9.435 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.35 //y=1.58 //x2=8.95 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.465 //y=1.495 //x2=8.465 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.465 //y=1.495 //x2=8.465 //y2=0.88
ends PM_DLATCH\%noxref_13

subckt PM_DLATCH\%noxref_14 ( 7 8 15 16 23 24 25 )
c43 ( 25 0 ) capacitor c=0.0306628f //x=15.725 //y=5.025
c44 ( 24 0 ) capacitor c=0.0185379f //x=14.845 //y=5.025
c45 ( 23 0 ) capacitor c=0.0409962f //x=13.975 //y=5.025
c46 ( 16 0 ) capacitor c=0.00193672f //x=15.075 //y=6.91
c47 ( 15 0 ) capacitor c=0.0129692f //x=15.785 //y=6.91
c48 ( 8 0 ) capacitor c=0.00576007f //x=14.195 //y=5.21
c49 ( 7 0 ) capacitor c=0.0170172f //x=14.905 //y=5.21
r50 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.87 //y=6.825 //x2=15.87 //y2=6.74
r51 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.785 //y=6.91 //x2=15.87 //y2=6.825
r52 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=15.785 //y=6.91 //x2=15.075 //y2=6.91
r53 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.99 //y=6.825 //x2=15.075 //y2=6.91
r54 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=14.99 //y=6.825 //x2=14.99 //y2=6.4
r55 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=14.99 //y=5.295 //x2=14.99 //y2=5.72
r56 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.905 //y=5.21 //x2=14.99 //y2=5.295
r57 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=14.905 //y=5.21 //x2=14.195 //y2=5.21
r58 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.11 //y=5.295 //x2=14.195 //y2=5.21
r59 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=14.11 //y=5.295 //x2=14.11 //y2=5.72
ends PM_DLATCH\%noxref_14

subckt PM_DLATCH\%noxref_15 ( 7 8 15 16 23 24 25 )
c42 ( 25 0 ) capacitor c=0.0307189f //x=19.055 //y=5.025
c43 ( 24 0 ) capacitor c=0.0185379f //x=18.175 //y=5.025
c44 ( 23 0 ) capacitor c=0.0410313f //x=17.305 //y=5.025
c45 ( 16 0 ) capacitor c=0.00193672f //x=18.405 //y=6.91
c46 ( 15 0 ) capacitor c=0.0132919f //x=19.115 //y=6.91
c47 ( 8 0 ) capacitor c=0.0056411f //x=17.525 //y=5.21
c48 ( 7 0 ) capacitor c=0.0169676f //x=18.235 //y=5.21
r49 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.2 //y=6.825 //x2=19.2 //y2=6.74
r50 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.115 //y=6.91 //x2=19.2 //y2=6.825
r51 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=19.115 //y=6.91 //x2=18.405 //y2=6.91
r52 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.32 //y=6.825 //x2=18.405 //y2=6.91
r53 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=18.32 //y=6.825 //x2=18.32 //y2=6.4
r54 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=18.32 //y=5.295 //x2=18.32 //y2=5.72
r55 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.235 //y=5.21 //x2=18.32 //y2=5.295
r56 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=18.235 //y=5.21 //x2=17.525 //y2=5.21
r57 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.44 //y=5.295 //x2=17.525 //y2=5.21
r58 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=17.44 //y=5.295 //x2=17.44 //y2=5.72
ends PM_DLATCH\%noxref_15

