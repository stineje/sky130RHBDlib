* SPICE3 file created from AND3X1.ext - technology: sky130A

.subckt AND3X1 Y A B C VPB VNB
X0 VPB a_342_166# a_277_1004# VPB sky130_fd_pr__pfet_01v8 ad=3.36e+12p pd=2.736e+07u as=0p ps=0u w=2e+06u l=150000u M=2
X1 VNB a_147_159# a_91_75# VNB sky130_fd_pr__nfet_01v8 ad=1.3199e+12p pd=9.67e+06u as=0p ps=0u w=3e+06u l=150000u
X2 VPB a_599_943# a_277_1004# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X3 a_372_182# a_342_166# a_91_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4 a_277_1004# a_147_159# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X5 VPB a_277_1004# a_1147_182# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X6 a_1147_182# a_277_1004# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X7 a_277_1004# a_599_943# a_372_182# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends
