magic
tech sky130A
magscale 1 2
timestamp 1652332182
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 1611 945 1645 979
rect 131 871 165 905
rect 649 871 683 905
rect 871 871 905 905
rect 945 871 979 905
rect 2055 871 2089 905
rect 131 797 165 831
rect 649 797 683 831
rect 871 797 905 831
rect 2055 797 2089 831
rect 131 723 165 757
rect 649 723 683 757
rect 945 723 979 757
rect 1611 723 1645 757
rect 2055 723 2089 757
rect 131 649 165 683
rect 649 649 683 683
rect 945 649 979 683
rect 1315 649 1349 683
rect 2055 649 2089 683
rect 131 575 165 609
rect 649 575 683 609
rect 2055 575 2089 609
rect 131 501 165 535
rect 649 501 683 535
rect 1611 501 1645 535
rect 2055 501 2089 535
rect 945 427 979 461
rect 1315 427 1349 461
rect 1611 427 1645 461
<< metal1 >>
rect -34 1446 2254 1514
rect -34 -34 2254 34
use xnor2x1_pcell  xnor2x1_pcell_0 pcells
timestamp 1652332156
transform 1 0 0 0 1 0
box -87 -34 2307 1550
<< labels >>
rlabel locali 1611 723 1645 757 1 Y
port 1 nsew signal output
rlabel locali 1611 501 1645 535 1 Y
port 1 nsew signal output
rlabel locali 1611 427 1645 461 1 Y
port 1 nsew signal output
rlabel locali 1611 945 1645 979 1 Y
port 1 nsew signal output
rlabel locali 945 723 979 757 1 Y
port 1 nsew signal output
rlabel locali 945 649 979 683 1 Y
port 1 nsew signal output
rlabel locali 945 427 979 461 1 Y
port 1 nsew signal output
rlabel locali 945 871 979 905 1 Y
port 1 nsew signal output
rlabel locali 131 871 165 905 1 A
port 2 nsew signal input
rlabel locali 131 797 165 831 1 A
port 2 nsew signal input
rlabel locali 131 723 165 757 1 A
port 2 nsew signal input
rlabel locali 131 649 165 683 1 A
port 2 nsew signal input
rlabel locali 131 575 165 609 1 A
port 2 nsew signal input
rlabel locali 131 501 165 535 1 A
port 2 nsew signal input
rlabel locali 649 501 683 535 1 A
port 2 nsew signal input
rlabel locali 649 575 683 609 1 A
port 2 nsew signal input
rlabel locali 649 649 683 683 1 A
port 2 nsew signal input
rlabel locali 649 723 683 757 1 A
port 2 nsew signal input
rlabel locali 649 797 683 831 1 A
port 2 nsew signal input
rlabel locali 649 871 683 905 1 A
port 2 nsew signal input
rlabel locali 2055 649 2089 683 1 B
port 3 nsew signal input
rlabel locali 2055 575 2089 609 1 B
port 3 nsew signal input
rlabel locali 2055 723 2089 757 1 B
port 3 nsew signal input
rlabel locali 2055 501 2089 535 1 B
port 3 nsew signal input
rlabel locali 2055 797 2089 831 1 B
port 3 nsew signal input
rlabel locali 2055 871 2089 905 1 B
port 3 nsew signal input
rlabel locali 871 797 905 831 1 B
port 3 nsew signal input
rlabel locali 1315 649 1349 683 1 B
port 3 nsew signal input
rlabel locali 1315 427 1349 461 1 B
port 3 nsew signal input
rlabel locali 871 871 905 905 1 B
port 3 nsew signal input
rlabel metal1 -34 1446 2254 1514 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 -34 -34 2254 34 1 GND
port 5 nsew ground bidirectional abutment


<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 2220 1480
string LEFsymmetry X Y R90
<< end >>
