magic
tech sky130A
magscale 1 2
timestamp 1651250933
<< nwell >>
rect -84 832 1416 1575
<< nmos >>
rect 168 316 198 377
tri 198 316 214 332 sw
rect 362 324 392 377
tri 392 324 408 340 sw
rect 168 286 274 316
tri 274 286 304 316 sw
rect 362 294 468 324
tri 468 294 498 324 sw
rect 168 185 198 286
tri 198 270 214 286 nw
tri 258 270 274 286 ne
tri 198 185 214 201 sw
tri 258 185 274 201 se
rect 274 185 304 286
rect 362 193 392 294
tri 392 278 408 294 nw
tri 452 278 468 294 ne
tri 392 193 408 209 sw
tri 452 193 468 209 se
rect 468 193 498 294
tri 168 155 198 185 ne
rect 198 155 274 185
tri 274 155 304 185 nw
tri 362 163 392 193 ne
rect 392 163 468 193
tri 468 163 498 193 nw
rect 834 324 864 377
tri 864 324 880 340 sw
rect 1028 324 1058 377
tri 1058 324 1074 340 sw
rect 834 294 940 324
tri 940 294 970 324 sw
rect 834 193 864 294
tri 864 278 880 294 nw
tri 924 278 940 294 ne
tri 864 193 880 209 sw
tri 924 193 940 209 se
rect 940 193 970 294
rect 1028 294 1134 324
tri 1134 294 1164 324 sw
rect 1028 279 1059 294
tri 1059 279 1074 294 nw
tri 1118 279 1133 294 ne
rect 1133 279 1164 294
tri 834 163 864 193 ne
rect 864 163 940 193
tri 940 163 970 193 nw
rect 1028 193 1058 279
tri 1058 193 1074 209 sw
tri 1118 193 1134 209 se
rect 1134 193 1164 279
tri 1028 163 1058 193 ne
rect 1058 163 1134 193
tri 1134 163 1164 193 nw
<< pmos >>
rect 187 1050 217 1450
rect 275 1050 305 1450
rect 363 1050 393 1450
rect 451 1050 481 1450
rect 853 1051 883 1451
rect 941 1051 971 1451
rect 1029 1051 1059 1451
rect 1117 1051 1147 1451
<< ndiff >>
rect 112 361 168 377
rect 112 327 122 361
rect 156 327 168 361
rect 112 289 168 327
rect 198 361 362 377
rect 198 332 219 361
tri 198 316 214 332 ne
rect 214 327 219 332
rect 253 327 316 361
rect 350 327 362 361
rect 214 316 362 327
rect 392 340 554 377
tri 392 324 408 340 ne
rect 408 324 554 340
rect 112 255 122 289
rect 156 255 168 289
tri 274 286 304 316 ne
rect 304 289 362 316
tri 468 294 498 324 ne
rect 112 221 168 255
rect 112 187 122 221
rect 156 187 168 221
rect 112 155 168 187
tri 198 270 214 286 se
rect 214 270 258 286
tri 258 270 274 286 sw
rect 198 236 274 270
rect 198 202 219 236
rect 253 202 274 236
rect 198 201 274 202
tri 198 185 214 201 ne
rect 214 185 258 201
tri 258 185 274 201 nw
rect 304 255 316 289
rect 350 255 362 289
rect 304 221 362 255
rect 304 187 316 221
rect 350 187 362 221
tri 392 278 408 294 se
rect 408 278 452 294
tri 452 278 468 294 sw
rect 392 245 468 278
rect 392 211 413 245
rect 447 211 468 245
rect 392 209 468 211
tri 392 193 408 209 ne
rect 408 193 452 209
tri 452 193 468 209 nw
rect 498 289 554 324
rect 498 255 510 289
rect 544 255 554 289
rect 498 221 554 255
tri 168 155 198 185 sw
tri 274 155 304 185 se
rect 304 163 362 187
tri 362 163 392 193 sw
tri 468 163 498 193 se
rect 498 187 510 221
rect 544 187 554 221
rect 498 163 554 187
rect 304 155 554 163
rect 112 151 554 155
rect 112 117 122 151
rect 156 117 316 151
rect 350 117 413 151
rect 447 117 510 151
rect 544 117 554 151
rect 112 101 554 117
rect 778 361 834 377
rect 778 327 788 361
rect 822 327 834 361
rect 778 289 834 327
rect 864 340 1028 377
tri 864 324 880 340 ne
rect 880 324 1028 340
rect 1058 340 1220 377
tri 1058 324 1074 340 ne
rect 1074 324 1220 340
tri 940 294 970 324 ne
rect 778 255 788 289
rect 822 255 834 289
rect 778 221 834 255
rect 778 187 788 221
rect 822 187 834 221
tri 864 278 880 294 se
rect 880 278 924 294
tri 924 278 940 294 sw
rect 864 245 940 278
rect 864 211 885 245
rect 919 211 940 245
rect 864 209 940 211
tri 864 193 880 209 ne
rect 880 193 924 209
tri 924 193 940 209 nw
rect 970 289 1028 324
tri 1134 294 1164 324 ne
rect 970 255 982 289
rect 1016 255 1028 289
tri 1059 279 1074 294 se
rect 1074 279 1118 294
tri 1118 279 1133 294 sw
rect 1164 289 1220 324
rect 970 221 1028 255
rect 778 163 834 187
tri 834 163 864 193 sw
tri 940 163 970 193 se
rect 970 187 982 221
rect 1016 187 1028 221
rect 1058 245 1134 279
rect 1058 211 1079 245
rect 1113 211 1134 245
rect 1058 209 1134 211
tri 1058 193 1074 209 ne
rect 1074 193 1118 209
tri 1118 193 1134 209 nw
rect 1164 255 1176 289
rect 1210 255 1220 289
rect 1164 221 1220 255
rect 970 163 1028 187
tri 1028 163 1058 193 sw
tri 1134 163 1164 193 se
rect 1164 187 1176 221
rect 1210 187 1220 221
rect 1164 163 1220 187
rect 778 151 1220 163
rect 778 117 788 151
rect 822 117 885 151
rect 919 117 982 151
rect 1016 117 1079 151
rect 1113 117 1176 151
rect 1210 117 1220 151
rect 778 101 1220 117
<< pdiff >>
rect 131 1412 187 1450
rect 131 1378 141 1412
rect 175 1378 187 1412
rect 131 1344 187 1378
rect 131 1310 141 1344
rect 175 1310 187 1344
rect 131 1276 187 1310
rect 131 1242 141 1276
rect 175 1242 187 1276
rect 131 1208 187 1242
rect 131 1174 141 1208
rect 175 1174 187 1208
rect 131 1139 187 1174
rect 131 1105 141 1139
rect 175 1105 187 1139
rect 131 1050 187 1105
rect 217 1412 275 1450
rect 217 1378 229 1412
rect 263 1378 275 1412
rect 217 1344 275 1378
rect 217 1310 229 1344
rect 263 1310 275 1344
rect 217 1276 275 1310
rect 217 1242 229 1276
rect 263 1242 275 1276
rect 217 1208 275 1242
rect 217 1174 229 1208
rect 263 1174 275 1208
rect 217 1139 275 1174
rect 217 1105 229 1139
rect 263 1105 275 1139
rect 217 1050 275 1105
rect 305 1412 363 1450
rect 305 1378 317 1412
rect 351 1378 363 1412
rect 305 1344 363 1378
rect 305 1310 317 1344
rect 351 1310 363 1344
rect 305 1276 363 1310
rect 305 1242 317 1276
rect 351 1242 363 1276
rect 305 1208 363 1242
rect 305 1174 317 1208
rect 351 1174 363 1208
rect 305 1050 363 1174
rect 393 1412 451 1450
rect 393 1378 405 1412
rect 439 1378 451 1412
rect 393 1344 451 1378
rect 393 1310 405 1344
rect 439 1310 451 1344
rect 393 1276 451 1310
rect 393 1242 405 1276
rect 439 1242 451 1276
rect 393 1208 451 1242
rect 393 1174 405 1208
rect 439 1174 451 1208
rect 393 1139 451 1174
rect 393 1105 405 1139
rect 439 1105 451 1139
rect 393 1050 451 1105
rect 481 1412 535 1450
rect 481 1378 493 1412
rect 527 1378 535 1412
rect 481 1344 535 1378
rect 481 1310 493 1344
rect 527 1310 535 1344
rect 481 1276 535 1310
rect 481 1242 493 1276
rect 527 1242 535 1276
rect 481 1208 535 1242
rect 481 1174 493 1208
rect 527 1174 535 1208
rect 481 1050 535 1174
rect 797 1411 853 1451
rect 797 1377 807 1411
rect 841 1377 853 1411
rect 797 1343 853 1377
rect 797 1309 807 1343
rect 841 1309 853 1343
rect 797 1275 853 1309
rect 797 1241 807 1275
rect 841 1241 853 1275
rect 797 1207 853 1241
rect 797 1173 807 1207
rect 841 1173 853 1207
rect 797 1139 853 1173
rect 797 1105 807 1139
rect 841 1105 853 1139
rect 797 1051 853 1105
rect 883 1411 941 1451
rect 883 1377 895 1411
rect 929 1377 941 1411
rect 883 1343 941 1377
rect 883 1309 895 1343
rect 929 1309 941 1343
rect 883 1275 941 1309
rect 883 1241 895 1275
rect 929 1241 941 1275
rect 883 1207 941 1241
rect 883 1173 895 1207
rect 929 1173 941 1207
rect 883 1051 941 1173
rect 971 1411 1029 1451
rect 971 1377 983 1411
rect 1017 1377 1029 1411
rect 971 1343 1029 1377
rect 971 1309 983 1343
rect 1017 1309 1029 1343
rect 971 1275 1029 1309
rect 971 1241 983 1275
rect 1017 1241 1029 1275
rect 971 1207 1029 1241
rect 971 1173 983 1207
rect 1017 1173 1029 1207
rect 971 1139 1029 1173
rect 971 1105 983 1139
rect 1017 1105 1029 1139
rect 971 1051 1029 1105
rect 1059 1343 1117 1451
rect 1059 1309 1071 1343
rect 1105 1309 1117 1343
rect 1059 1275 1117 1309
rect 1059 1241 1071 1275
rect 1105 1241 1117 1275
rect 1059 1207 1117 1241
rect 1059 1173 1071 1207
rect 1105 1173 1117 1207
rect 1059 1139 1117 1173
rect 1059 1105 1071 1139
rect 1105 1105 1117 1139
rect 1059 1051 1117 1105
rect 1147 1411 1201 1451
rect 1147 1377 1159 1411
rect 1193 1377 1201 1411
rect 1147 1343 1201 1377
rect 1147 1309 1159 1343
rect 1193 1309 1201 1343
rect 1147 1275 1201 1309
rect 1147 1241 1159 1275
rect 1193 1241 1201 1275
rect 1147 1207 1201 1241
rect 1147 1173 1159 1207
rect 1193 1173 1201 1207
rect 1147 1051 1201 1173
<< ndiffc >>
rect 122 327 156 361
rect 219 327 253 361
rect 316 327 350 361
rect 122 255 156 289
rect 122 187 156 221
rect 219 202 253 236
rect 316 255 350 289
rect 316 187 350 221
rect 413 211 447 245
rect 510 255 544 289
rect 510 187 544 221
rect 122 117 156 151
rect 316 117 350 151
rect 413 117 447 151
rect 510 117 544 151
rect 788 327 822 361
rect 788 255 822 289
rect 788 187 822 221
rect 885 211 919 245
rect 982 255 1016 289
rect 982 187 1016 221
rect 1079 211 1113 245
rect 1176 255 1210 289
rect 1176 187 1210 221
rect 788 117 822 151
rect 885 117 919 151
rect 982 117 1016 151
rect 1079 117 1113 151
rect 1176 117 1210 151
<< pdiffc >>
rect 141 1378 175 1412
rect 141 1310 175 1344
rect 141 1242 175 1276
rect 141 1174 175 1208
rect 141 1105 175 1139
rect 229 1378 263 1412
rect 229 1310 263 1344
rect 229 1242 263 1276
rect 229 1174 263 1208
rect 229 1105 263 1139
rect 317 1378 351 1412
rect 317 1310 351 1344
rect 317 1242 351 1276
rect 317 1174 351 1208
rect 405 1378 439 1412
rect 405 1310 439 1344
rect 405 1242 439 1276
rect 405 1174 439 1208
rect 405 1105 439 1139
rect 493 1378 527 1412
rect 493 1310 527 1344
rect 493 1242 527 1276
rect 493 1174 527 1208
rect 807 1377 841 1411
rect 807 1309 841 1343
rect 807 1241 841 1275
rect 807 1173 841 1207
rect 807 1105 841 1139
rect 895 1377 929 1411
rect 895 1309 929 1343
rect 895 1241 929 1275
rect 895 1173 929 1207
rect 983 1377 1017 1411
rect 983 1309 1017 1343
rect 983 1241 1017 1275
rect 983 1173 1017 1207
rect 983 1105 1017 1139
rect 1071 1309 1105 1343
rect 1071 1241 1105 1275
rect 1071 1173 1105 1207
rect 1071 1105 1105 1139
rect 1159 1377 1193 1411
rect 1159 1309 1193 1343
rect 1159 1241 1193 1275
rect 1159 1173 1193 1207
<< psubdiff >>
rect -31 546 1363 572
rect -31 512 -17 546
rect 17 512 649 546
rect 683 512 1315 546
rect 1349 512 1363 546
rect -31 510 1363 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 635 474 697 510
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 635 368 649 402
rect 683 368 697 402
rect 1301 474 1363 510
rect 1301 440 1315 474
rect 1349 440 1363 474
rect 1301 402 1363 440
rect 635 330 697 368
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect -31 47 31 80
rect 635 80 649 114
rect 683 80 697 114
rect 1301 368 1315 402
rect 1349 368 1363 402
rect 1301 330 1363 368
rect 1301 296 1315 330
rect 1349 296 1363 330
rect 1301 258 1363 296
rect 1301 224 1315 258
rect 1349 224 1363 258
rect 1301 186 1363 224
rect 1301 152 1315 186
rect 1349 152 1363 186
rect 1301 114 1363 152
rect 635 47 697 80
rect 1301 80 1315 114
rect 1349 80 1363 114
rect 1301 47 1363 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1027 47
rect 1061 13 1099 47
rect 1133 13 1171 47
rect 1205 13 1243 47
rect 1277 13 1363 47
rect -31 11 31 13
rect 635 11 697 13
rect 1301 11 1363 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1027 1539
rect 1061 1505 1099 1539
rect 1133 1505 1171 1539
rect 1205 1505 1243 1539
rect 1277 1505 1363 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 635 1470 697 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 1301 1470 1363 1505
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 635 1076 649 1110
rect 683 1076 697 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 635 1038 697 1076
rect 1301 1436 1315 1470
rect 1349 1436 1363 1470
rect 1301 1398 1363 1436
rect 1301 1364 1315 1398
rect 1349 1364 1363 1398
rect 1301 1326 1363 1364
rect 1301 1292 1315 1326
rect 1349 1292 1363 1326
rect 1301 1254 1363 1292
rect 1301 1220 1315 1254
rect 1349 1220 1363 1254
rect 1301 1182 1363 1220
rect 1301 1148 1315 1182
rect 1349 1148 1363 1182
rect 1301 1110 1363 1148
rect 1301 1076 1315 1110
rect 1349 1076 1363 1110
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect -31 930 31 932
rect 635 932 649 966
rect 683 932 697 966
rect 1301 1038 1363 1076
rect 1301 1004 1315 1038
rect 1349 1004 1363 1038
rect 1301 966 1363 1004
rect 635 930 697 932
rect 1301 932 1315 966
rect 1349 932 1363 966
rect 1301 930 1363 932
rect -31 868 1363 930
<< psubdiffcont >>
rect -17 512 17 546
rect 649 512 683 546
rect 1315 512 1349 546
rect -17 440 17 474
rect -17 368 17 402
rect 649 440 683 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 649 368 683 402
rect 1315 440 1349 474
rect 649 296 683 330
rect 649 224 683 258
rect 649 152 683 186
rect 649 80 683 114
rect 1315 368 1349 402
rect 1315 296 1349 330
rect 1315 224 1349 258
rect 1315 152 1349 186
rect 1315 80 1349 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1027 13 1061 47
rect 1099 13 1133 47
rect 1171 13 1205 47
rect 1243 13 1277 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1027 1505 1061 1539
rect 1099 1505 1133 1539
rect 1171 1505 1205 1539
rect 1243 1505 1277 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 649 1436 683 1470
rect 649 1364 683 1398
rect 649 1292 683 1326
rect 649 1220 683 1254
rect 649 1148 683 1182
rect 649 1076 683 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1315 1436 1349 1470
rect 1315 1364 1349 1398
rect 1315 1292 1349 1326
rect 1315 1220 1349 1254
rect 1315 1148 1349 1182
rect 1315 1076 1349 1110
rect 649 1004 683 1038
rect 649 932 683 966
rect 1315 1004 1349 1038
rect 1315 932 1349 966
<< poly >>
rect 187 1450 217 1476
rect 275 1450 305 1476
rect 363 1450 393 1476
rect 451 1450 481 1476
rect 853 1451 883 1477
rect 941 1451 971 1477
rect 1029 1451 1059 1477
rect 1117 1451 1147 1477
rect 187 1019 217 1050
rect 275 1019 305 1050
rect 363 1019 393 1050
rect 451 1019 481 1050
rect 187 1003 305 1019
rect 187 989 205 1003
rect 195 969 205 989
rect 239 989 305 1003
rect 349 1003 481 1019
rect 239 969 249 989
rect 195 953 249 969
rect 349 969 359 1003
rect 393 989 481 1003
rect 853 1020 883 1051
rect 941 1020 971 1051
rect 1029 1020 1059 1051
rect 1117 1020 1147 1051
rect 393 969 403 989
rect 349 953 403 969
rect 830 1004 971 1020
rect 830 970 840 1004
rect 874 990 971 1004
rect 1016 1004 1147 1020
rect 874 970 884 990
rect 830 954 884 970
rect 1016 970 1026 1004
rect 1060 990 1147 1004
rect 1060 970 1070 990
rect 1016 954 1070 970
rect 195 461 249 477
rect 195 441 205 461
rect 168 427 205 441
rect 239 427 249 461
rect 168 411 249 427
rect 343 461 397 477
rect 343 427 353 461
rect 387 427 397 461
rect 343 411 397 427
rect 861 461 915 477
rect 861 441 871 461
rect 168 377 198 411
rect 362 377 392 411
rect 834 427 871 441
rect 905 427 915 461
rect 834 411 915 427
rect 1009 461 1063 477
rect 1009 427 1019 461
rect 1053 427 1063 461
rect 1009 411 1063 427
rect 834 377 864 411
rect 1028 377 1058 411
<< polycont >>
rect 205 969 239 1003
rect 359 969 393 1003
rect 840 970 874 1004
rect 1026 970 1060 1004
rect 205 427 239 461
rect 353 427 387 461
rect 871 427 905 461
rect 1019 427 1053 461
<< locali >>
rect -31 1539 1363 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1027 1539
rect 1061 1505 1099 1539
rect 1133 1505 1171 1539
rect 1205 1505 1243 1539
rect 1277 1505 1363 1539
rect -31 1492 1363 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 141 1412 175 1492
rect 141 1344 175 1378
rect 141 1276 175 1310
rect 141 1208 175 1242
rect 141 1139 175 1174
rect 141 1073 175 1105
rect 229 1412 263 1450
rect 229 1344 263 1378
rect 229 1276 263 1310
rect 229 1208 263 1242
rect 229 1139 263 1174
rect 317 1412 351 1492
rect 317 1344 351 1378
rect 317 1276 351 1310
rect 317 1208 351 1242
rect 317 1157 351 1174
rect 405 1412 439 1450
rect 405 1344 439 1378
rect 405 1276 439 1310
rect 405 1208 439 1242
rect 229 1103 263 1105
rect 405 1139 439 1174
rect 493 1412 527 1492
rect 493 1344 527 1378
rect 493 1276 527 1310
rect 493 1208 527 1242
rect 493 1157 527 1174
rect 635 1470 697 1492
rect 635 1436 649 1470
rect 683 1436 697 1470
rect 635 1398 697 1436
rect 635 1364 649 1398
rect 683 1364 697 1398
rect 635 1326 697 1364
rect 635 1292 649 1326
rect 683 1292 697 1326
rect 635 1254 697 1292
rect 635 1220 649 1254
rect 683 1220 697 1254
rect 635 1182 697 1220
rect 405 1103 439 1105
rect 635 1148 649 1182
rect 683 1148 697 1182
rect 635 1110 697 1148
rect 229 1069 535 1103
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 359 1003 393 1019
rect 205 609 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 575
rect 205 411 239 427
rect 353 969 359 988
rect 353 953 393 969
rect 353 683 387 953
rect 353 461 387 649
rect 353 411 387 427
rect 501 535 535 1069
rect 635 1076 649 1110
rect 683 1076 697 1110
rect 635 1038 697 1076
rect 807 1411 841 1451
rect 807 1343 841 1377
rect 807 1275 841 1309
rect 807 1207 841 1241
rect 807 1139 841 1173
rect 895 1411 929 1492
rect 1301 1470 1363 1492
rect 895 1343 929 1377
rect 895 1275 929 1309
rect 895 1207 929 1241
rect 895 1157 929 1173
rect 983 1411 1193 1445
rect 983 1343 1017 1377
rect 983 1275 1017 1309
rect 983 1207 1017 1241
rect 983 1139 1017 1173
rect 807 1071 1017 1105
rect 1071 1343 1105 1359
rect 1071 1275 1105 1309
rect 1071 1207 1105 1241
rect 1071 1139 1105 1173
rect 1159 1343 1193 1377
rect 1159 1275 1193 1309
rect 1159 1207 1193 1241
rect 1159 1157 1193 1173
rect 1301 1436 1315 1470
rect 1349 1436 1363 1470
rect 1301 1398 1363 1436
rect 1301 1364 1315 1398
rect 1349 1364 1363 1398
rect 1301 1326 1363 1364
rect 1301 1292 1315 1326
rect 1349 1292 1363 1326
rect 1301 1254 1363 1292
rect 1301 1220 1315 1254
rect 1349 1220 1363 1254
rect 1301 1182 1363 1220
rect 1301 1148 1315 1182
rect 1349 1148 1363 1182
rect 1301 1110 1363 1148
rect 1071 1071 1201 1105
rect 635 1004 649 1038
rect 683 1004 697 1038
rect 635 966 697 1004
rect 635 932 649 966
rect 683 932 697 966
rect 840 1004 874 1020
rect 1026 1004 1060 1020
rect 874 970 905 988
rect 840 954 905 970
rect 635 868 697 932
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 122 361 156 377
rect 316 361 350 377
rect 501 376 535 501
rect 156 327 219 361
rect 253 327 316 361
rect 122 289 156 327
rect 122 221 156 255
rect 316 289 350 327
rect 122 151 156 187
rect 122 101 156 117
rect 219 236 253 252
rect -31 62 31 80
rect 219 62 253 202
rect 316 221 350 255
rect 413 342 535 376
rect 635 546 697 572
rect 635 512 649 546
rect 683 512 697 546
rect 635 474 697 512
rect 635 440 649 474
rect 683 440 697 474
rect 635 402 697 440
rect 871 535 905 954
rect 871 461 905 501
rect 871 411 905 427
rect 1019 970 1026 988
rect 1019 954 1060 970
rect 1019 757 1053 954
rect 1019 461 1053 723
rect 1019 411 1053 427
rect 1167 831 1201 1071
rect 1301 1076 1315 1110
rect 1349 1076 1363 1110
rect 1301 1038 1363 1076
rect 1301 1004 1315 1038
rect 1349 1004 1363 1038
rect 1301 966 1363 1004
rect 1301 932 1315 966
rect 1349 932 1363 966
rect 1301 868 1363 932
rect 635 368 649 402
rect 683 368 697 402
rect 413 245 447 342
rect 635 330 697 368
rect 413 195 447 211
rect 510 289 544 305
rect 510 221 544 255
rect 316 151 350 187
rect 510 151 544 187
rect 350 117 413 151
rect 447 117 510 151
rect 316 101 350 117
rect 510 101 544 117
rect 635 296 649 330
rect 683 296 697 330
rect 635 258 697 296
rect 635 224 649 258
rect 683 224 697 258
rect 635 186 697 224
rect 635 152 649 186
rect 683 152 697 186
rect 635 114 697 152
rect 635 80 649 114
rect 683 80 697 114
rect 635 62 697 80
rect 788 361 822 377
rect 1167 376 1201 797
rect 788 289 822 327
rect 788 221 822 255
rect 885 342 1201 376
rect 1301 546 1363 572
rect 1301 512 1315 546
rect 1349 512 1363 546
rect 1301 474 1363 512
rect 1301 440 1315 474
rect 1349 440 1363 474
rect 1301 402 1363 440
rect 1301 368 1315 402
rect 1349 368 1363 402
rect 885 245 919 342
rect 885 195 919 211
rect 982 289 1016 306
rect 982 221 1016 255
rect 788 151 822 187
rect 1079 245 1113 342
rect 1301 330 1363 368
rect 1079 195 1113 211
rect 1176 289 1210 306
rect 1176 221 1210 255
rect 982 151 1016 187
rect 1176 151 1210 187
rect 822 117 885 151
rect 919 117 982 151
rect 1016 117 1079 151
rect 1113 117 1176 151
rect 788 62 822 117
rect 885 62 919 117
rect 982 62 1016 117
rect 1079 62 1113 117
rect 1176 62 1210 117
rect 1301 296 1315 330
rect 1349 296 1363 330
rect 1301 258 1363 296
rect 1301 224 1315 258
rect 1349 224 1363 258
rect 1301 186 1363 224
rect 1301 152 1315 186
rect 1349 152 1363 186
rect 1301 114 1363 152
rect 1301 80 1315 114
rect 1349 80 1363 114
rect 1301 62 1363 80
rect -31 47 1363 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1027 47
rect 1061 13 1099 47
rect 1133 13 1171 47
rect 1205 13 1243 47
rect 1277 13 1363 47
rect -31 0 1363 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 721 1505 755 1539
rect 793 1505 827 1539
rect 865 1505 899 1539
rect 937 1505 971 1539
rect 1027 1505 1061 1539
rect 1099 1505 1133 1539
rect 1171 1505 1205 1539
rect 1243 1505 1277 1539
rect 205 575 239 609
rect 353 649 387 683
rect 501 501 535 535
rect 871 501 905 535
rect 1019 723 1053 757
rect 1167 797 1201 831
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
rect 721 13 755 47
rect 793 13 827 47
rect 865 13 899 47
rect 937 13 971 47
rect 1027 13 1061 47
rect 1099 13 1133 47
rect 1171 13 1205 47
rect 1243 13 1277 47
<< metal1 >>
rect -31 1539 1363 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 721 1539
rect 755 1505 793 1539
rect 827 1505 865 1539
rect 899 1505 937 1539
rect 971 1505 1027 1539
rect 1061 1505 1099 1539
rect 1133 1505 1171 1539
rect 1205 1505 1243 1539
rect 1277 1505 1363 1539
rect -31 1492 1363 1505
rect 1161 831 1207 837
rect 1155 797 1167 831
rect 1201 797 1237 831
rect 1161 791 1207 797
rect 1013 757 1059 763
rect 983 723 1019 757
rect 1053 723 1065 757
rect 1013 717 1059 723
rect 347 683 393 689
rect 317 649 353 683
rect 387 649 399 683
rect 347 643 393 649
rect 199 609 245 615
rect 169 575 205 609
rect 239 575 251 609
rect 199 569 245 575
rect 495 535 541 541
rect 865 535 911 541
rect 489 501 501 535
rect 535 501 871 535
rect 905 501 917 535
rect 495 495 541 501
rect 865 495 911 501
rect -31 47 1363 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 721 47
rect 755 13 793 47
rect 827 13 865 47
rect 899 13 937 47
rect 971 13 1027 47
rect 1061 13 1099 47
rect 1133 13 1171 47
rect 1205 13 1243 47
rect 1277 13 1363 47
rect -31 0 1363 13
<< labels >>
rlabel metal1 1167 797 1201 831 1 YN
port 1 n
rlabel metal1 205 575 239 609 1 A
port 2 n
rlabel metal1 353 649 387 683 1 B
port 3 n
rlabel metal1 1019 723 1053 757 1 C
port 4 n
rlabel metal1 -31 1492 1363 1554 1 VDD
port 5 n
rlabel metal1 -31 0 1363 62 1 GND
port 6 n
<< end >>
