magic
tech sky130A
magscale 1 2
timestamp 1652367648
<< metal1 >>
rect 1201 501 1443 535
use invx1_pcell  invx1_pcell_0
timestamp 1652329846
transform 1 0 1332 0 1 0
box -87 -34 531 1550
use aoi3x1_pcell  aoi3x1_pcell_0
timestamp 1652367586
transform 1 0 0 0 1 0
box -87 -34 1419 1550
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 1480 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 1184 0 -1 518
box -53 -33 29 33
<< end >>
