// File: xor2X1_pcell.spi.pex
// Created: Tue Oct 15 16:01:28 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_XOR2X1_PCELL\%noxref_1 ( 19 31 35 38 43 49 55 61 69 77 80 85 89 101 \
 112 115 117 124 131 132 133 134 )
c165 ( 134 0 ) capacitor c=0.0583152f //x=9.375 //y=0.37
c166 ( 133 0 ) capacitor c=0.0210151f //x=6.54 //y=0.87
c167 ( 132 0 ) capacitor c=0.0210151f //x=3.21 //y=0.87
c168 ( 131 0 ) capacitor c=0.0582156f //x=0.495 //y=0.37
c169 ( 124 0 ) capacitor c=0.229233f //x=10.47 //y=0
c170 ( 117 0 ) capacitor c=0.103612f //x=8.88 //y=0
c171 ( 116 0 ) capacitor c=0.0044012f //x=6.73 //y=0
c172 ( 115 0 ) capacitor c=0.104587f //x=5.55 //y=0
c173 ( 114 0 ) capacitor c=0.0044012f //x=3.33 //y=0
c174 ( 112 0 ) capacitor c=0.102385f //x=2.22 //y=0
c175 ( 101 0 ) capacitor c=0.192508f //x=0.63 //y=0
c176 ( 92 0 ) capacitor c=0.00592191f //x=10.47 //y=0.45
c177 ( 89 0 ) capacitor c=0.00644318f //x=10.385 //y=0.535
c178 ( 88 0 ) capacitor c=0.00479856f //x=9.985 //y=0.45
c179 ( 85 0 ) capacitor c=0.00531808f //x=9.9 //y=0.535
c180 ( 80 0 ) capacitor c=0.00587411f //x=9.5 //y=0.45
c181 ( 77 0 ) capacitor c=0.0160123f //x=9.415 //y=0
c182 ( 69 0 ) capacitor c=0.0720515f //x=8.71 //y=0
c183 ( 61 0 ) capacitor c=0.0389232f //x=6.645 //y=0
c184 ( 55 0 ) capacitor c=0.072035f //x=5.38 //y=0
c185 ( 49 0 ) capacitor c=0.0389232f //x=3.315 //y=0
c186 ( 44 0 ) capacitor c=0.0360673f //x=1.685 //y=0
c187 ( 43 0 ) capacitor c=0.0160123f //x=2.05 //y=0
c188 ( 38 0 ) capacitor c=0.00587411f //x=1.6 //y=0.45
c189 ( 35 0 ) capacitor c=0.00534353f //x=1.515 //y=0.535
c190 ( 34 0 ) capacitor c=0.00479856f //x=1.115 //y=0.45
c191 ( 31 0 ) capacitor c=0.00707849f //x=1.03 //y=0.535
c192 ( 26 0 ) capacitor c=0.00592191f //x=0.63 //y=0.45
c193 ( 19 0 ) capacitor c=0.388313f //x=10.36 //y=0
r194 (  123 124 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=10.36 //y=0 //x2=10.47 //y2=0
r195 (  121 123 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=9.985 //y=0 //x2=10.36 //y2=0
r196 (  120 121 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=9.62 //y=0 //x2=9.985 //y2=0
r197 (  118 120 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=9.5 //y=0 //x2=9.62 //y2=0
r198 (  104 105 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.115 //y=0 //x2=1.6 //y2=0
r199 (  103 104 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.115 //y2=0
r200 (  101 103 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=0.63 //y=0 //x2=0.74 //y2=0
r201 (  93 134 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.62 //x2=10.47 //y2=0.535
r202 (  93 134 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.62 //x2=10.47 //y2=1.225
r203 (  92 134 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.45 //x2=10.47 //y2=0.535
r204 (  91 124 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.17 //x2=10.47 //y2=0
r205 (  91 92 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.17 //x2=10.47 //y2=0.45
r206 (  90 134 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.07 //y=0.535 //x2=9.985 //y2=0.535
r207 (  89 134 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.385 //y=0.535 //x2=10.47 //y2=0.535
r208 (  89 90 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=10.385 //y=0.535 //x2=10.07 //y2=0.535
r209 (  88 134 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.985 //y=0.45 //x2=9.985 //y2=0.535
r210 (  87 121 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.985 //y=0.17 //x2=9.985 //y2=0
r211 (  87 88 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=9.985 //y=0.17 //x2=9.985 //y2=0.45
r212 (  86 134 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.585 //y=0.535 //x2=9.5 //y2=0.535
r213 (  85 134 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.9 //y=0.535 //x2=9.985 //y2=0.535
r214 (  85 86 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=9.9 //y=0.535 //x2=9.585 //y2=0.535
r215 (  81 134 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.62 //x2=9.5 //y2=0.535
r216 (  81 134 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.62 //x2=9.5 //y2=1.225
r217 (  80 134 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.45 //x2=9.5 //y2=0.535
r218 (  79 118 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.17 //x2=9.5 //y2=0
r219 (  79 80 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.17 //x2=9.5 //y2=0.45
r220 (  78 117 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.05 //y=0 //x2=8.88 //y2=0
r221 (  77 118 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.415 //y=0 //x2=9.5 //y2=0
r222 (  77 78 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=9.415 //y=0 //x2=9.05 //y2=0
r223 (  72 74 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.03 //y=0 //x2=8.14 //y2=0
r224 (  70 116 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.815 //y=0 //x2=6.73 //y2=0
r225 (  70 72 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=6.815 //y=0 //x2=7.03 //y2=0
r226 (  69 117 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.71 //y=0 //x2=8.88 //y2=0
r227 (  69 74 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.71 //y=0 //x2=8.14 //y2=0
r228 (  65 116 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.73 //y=0.17 //x2=6.73 //y2=0
r229 (  65 133 ) resistor r=54.0749 //w=0.187 //l=0.79 //layer=li \
 //thickness=0.1 //x=6.73 //y=0.17 //x2=6.73 //y2=0.96
r230 (  62 115 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.55 //y2=0
r231 (  62 64 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.92 //y2=0
r232 (  61 116 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.645 //y=0 //x2=6.73 //y2=0
r233 (  61 64 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=6.645 //y=0 //x2=5.92 //y2=0
r234 (  56 114 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.485 //y=0 //x2=3.4 //y2=0
r235 (  56 58 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=3.485 //y=0 //x2=4.44 //y2=0
r236 (  55 115 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=5.55 //y2=0
r237 (  55 58 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=4.44 //y2=0
r238 (  51 114 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.4 //y=0.17 //x2=3.4 //y2=0
r239 (  51 132 ) resistor r=54.0749 //w=0.187 //l=0.79 //layer=li \
 //thickness=0.1 //x=3.4 //y=0.17 //x2=3.4 //y2=0.96
r240 (  50 112 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.39 //y=0 //x2=2.22 //y2=0
r241 (  49 114 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.315 //y=0 //x2=3.4 //y2=0
r242 (  49 50 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=3.315 //y=0 //x2=2.39 //y2=0
r243 (  44 105 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.6 //y2=0
r244 (  44 46 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.85 //y2=0
r245 (  43 112 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=2.22 //y2=0
r246 (  43 46 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=1.85 //y2=0
r247 (  39 131 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=0.535
r248 (  39 131 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=1.225
r249 (  38 131 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.45 //x2=1.6 //y2=0.535
r250 (  37 105 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0
r251 (  37 38 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0.45
r252 (  36 131 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.2 //y=0.535 //x2=1.115 //y2=0.535
r253 (  35 131 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.6 //y2=0.535
r254 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.2 //y2=0.535
r255 (  34 131 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.45 //x2=1.115 //y2=0.535
r256 (  33 104 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0
r257 (  33 34 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0.45
r258 (  32 131 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.715 //y=0.535 //x2=0.63 //y2=0.535
r259 (  31 131 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=1.115 //y2=0.535
r260 (  31 32 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=0.715 //y2=0.535
r261 (  27 131 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=0.535
r262 (  27 131 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=1.225
r263 (  26 131 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.45 //x2=0.63 //y2=0.535
r264 (  25 101 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0
r265 (  25 26 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0.45
r266 (  19 123 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r267 (  17 120 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=0 //x2=9.62 //y2=0
r268 (  17 19 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=9.62 //y=0 //x2=10.36 //y2=0
r269 (  15 74 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=0 //x2=8.14 //y2=0
r270 (  15 17 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=0 //x2=9.62 //y2=0
r271 (  13 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=0 //x2=7.03 //y2=0
r272 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=0 //x2=8.14 //y2=0
r273 (  11 64 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=0 //x2=5.92 //y2=0
r274 (  11 13 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=0 //x2=7.03 //y2=0
r275 (  9 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r276 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.92 //y2=0
r277 (  7 114 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=0 //x2=3.33 //y2=0
r278 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=0 //x2=4.44 //y2=0
r279 (  5 46 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r280 (  5 7 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=3.33 //y2=0
r281 (  2 103 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r282 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_XOR2X1_PCELL\%noxref_1

subckt PM_XOR2X1_PCELL\%noxref_2 ( 19 31 39 45 53 59 67 75 83 96 98 100 102 \
 106 107 108 109 110 111 112 )
c156 ( 112 0 ) capacitor c=0.0420685f //x=10.28 //y=5.02
c157 ( 111 0 ) capacitor c=0.0433633f //x=9.42 //y=5.02
c158 ( 110 0 ) capacitor c=0.0266033f //x=6.635 //y=5.02
c159 ( 109 0 ) capacitor c=0.0265296f //x=3.305 //y=5.02
c160 ( 108 0 ) capacitor c=0.0432963f //x=1.41 //y=5.02
c161 ( 107 0 ) capacitor c=0.0421443f //x=0.54 //y=5.02
c162 ( 106 0 ) capacitor c=0.232571f //x=10.36 //y=7.4
c163 ( 104 0 ) capacitor c=0.00591168f //x=9.62 //y=7.4
c164 ( 102 0 ) capacitor c=0.105702f //x=8.88 //y=7.4
c165 ( 101 0 ) capacitor c=0.00591168f //x=6.78 //y=7.4
c166 ( 100 0 ) capacitor c=0.111763f //x=5.55 //y=7.4
c167 ( 99 0 ) capacitor c=0.00591168f //x=3.45 //y=7.4
c168 ( 98 0 ) capacitor c=0.111559f //x=2.22 //y=7.4
c169 ( 97 0 ) capacitor c=0.00591168f //x=1.555 //y=7.4
c170 ( 96 0 ) capacitor c=0.232987f //x=0.74 //y=7.4
c171 ( 83 0 ) capacitor c=0.0289356f //x=10.34 //y=7.4
c172 ( 75 0 ) capacitor c=0.0181526f //x=9.46 //y=7.4
c173 ( 67 0 ) capacitor c=0.0747638f //x=8.71 //y=7.4
c174 ( 59 0 ) capacitor c=0.042882f //x=6.695 //y=7.4
c175 ( 53 0 ) capacitor c=0.074629f //x=5.38 //y=7.4
c176 ( 45 0 ) capacitor c=0.042884f //x=3.365 //y=7.4
c177 ( 39 0 ) capacitor c=0.0181526f //x=2.05 //y=7.4
c178 ( 31 0 ) capacitor c=0.0291066f //x=1.47 //y=7.4
c179 ( 19 0 ) capacitor c=0.40033f //x=10.36 //y=7.4
r180 (  85 106 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.425 //y=7.23 //x2=10.425 //y2=7.4
r181 (  85 112 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.425 //y=7.23 //x2=10.425 //y2=6.405
r182 (  84 104 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.63 //y=7.4 //x2=9.545 //y2=7.4
r183 (  83 106 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.34 //y=7.4 //x2=10.425 //y2=7.4
r184 (  83 84 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.34 //y=7.4 //x2=9.63 //y2=7.4
r185 (  77 104 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.545 //y=7.23 //x2=9.545 //y2=7.4
r186 (  77 111 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=9.545 //y=7.23 //x2=9.545 //y2=6.405
r187 (  76 102 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.05 //y=7.4 //x2=8.88 //y2=7.4
r188 (  75 104 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.46 //y=7.4 //x2=9.545 //y2=7.4
r189 (  75 76 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=9.46 //y=7.4 //x2=9.05 //y2=7.4
r190 (  70 72 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.03 //y=7.4 //x2=8.14 //y2=7.4
r191 (  68 101 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=6.78 //y2=7.4
r192 (  68 70 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=7.03 //y2=7.4
r193 (  67 102 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.71 //y=7.4 //x2=8.88 //y2=7.4
r194 (  67 72 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.71 //y=7.4 //x2=8.14 //y2=7.4
r195 (  63 101 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=7.4
r196 (  63 110 ) resistor r=80.4278 //w=0.187 //l=1.175 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=6.055
r197 (  60 100 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.55 //y2=7.4
r198 (  60 62 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.92 //y2=7.4
r199 (  59 101 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.78 //y2=7.4
r200 (  59 62 ) resistor r=27.7871 //w=0.357 //l=0.775 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=5.92 //y2=7.4
r201 (  54 99 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.535 //y=7.4 //x2=3.45 //y2=7.4
r202 (  54 56 ) resistor r=32.4482 //w=0.357 //l=0.905 //layer=li \
 //thickness=0.1 //x=3.535 //y=7.4 //x2=4.44 //y2=7.4
r203 (  53 100 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=5.55 //y2=7.4
r204 (  53 56 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=4.44 //y2=7.4
r205 (  49 99 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.45 //y=7.23 //x2=3.45 //y2=7.4
r206 (  49 109 ) resistor r=80.4278 //w=0.187 //l=1.175 //layer=li \
 //thickness=0.1 //x=3.45 //y=7.23 //x2=3.45 //y2=6.055
r207 (  46 98 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.39 //y=7.4 //x2=2.22 //y2=7.4
r208 (  46 48 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=2.39 //y=7.4 //x2=3.33 //y2=7.4
r209 (  45 99 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.365 //y=7.4 //x2=3.45 //y2=7.4
r210 (  45 48 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=3.365 //y=7.4 //x2=3.33 //y2=7.4
r211 (  40 97 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.555 //y2=7.4
r212 (  40 42 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.85 //y2=7.4
r213 (  39 98 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.05 //y=7.4 //x2=2.22 //y2=7.4
r214 (  39 42 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=7.4 //x2=1.85 //y2=7.4
r215 (  33 97 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=7.4
r216 (  33 108 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=6.405
r217 (  32 96 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.76 //y=7.4 //x2=0.675 //y2=7.4
r218 (  31 97 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=1.555 //y2=7.4
r219 (  31 32 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=0.76 //y2=7.4
r220 (  25 96 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=7.4
r221 (  25 107 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=6.405
r222 (  19 106 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r223 (  17 104 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=7.4 //x2=9.62 //y2=7.4
r224 (  17 19 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=9.62 //y=7.4 //x2=10.36 //y2=7.4
r225 (  15 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=7.4 //x2=8.14 //y2=7.4
r226 (  15 17 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=7.4 //x2=9.62 //y2=7.4
r227 (  13 70 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=7.4 //x2=7.03 //y2=7.4
r228 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=7.4 //x2=8.14 //y2=7.4
r229 (  11 62 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=7.4 //x2=5.92 //y2=7.4
r230 (  11 13 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=7.4 //x2=7.03 //y2=7.4
r231 (  9 56 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r232 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.92 //y2=7.4
r233 (  7 48 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=7.4 //x2=3.33 //y2=7.4
r234 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=7.4 //x2=4.44 //y2=7.4
r235 (  5 42 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r236 (  5 7 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=3.33 //y2=7.4
r237 (  2 96 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r238 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_XOR2X1_PCELL\%noxref_2

subckt PM_XOR2X1_PCELL\%noxref_3 ( 1 2 8 16 23 24 25 26 27 28 29 30 31 32 36 \
 37 38 40 46 47 48 49 50 51 55 57 60 61 66 80 )
c133 ( 80 0 ) capacitor c=0.0661295f //x=3.33 //y=4.7
c134 ( 66 0 ) capacitor c=0.0537799f //x=0.74 //y=2.085
c135 ( 61 0 ) capacitor c=0.0318948f //x=3.665 //y=1.215
c136 ( 60 0 ) capacitor c=0.0187407f //x=3.665 //y=0.87
c137 ( 57 0 ) capacitor c=0.0141798f //x=3.51 //y=1.37
c138 ( 55 0 ) capacitor c=0.0149852f //x=3.51 //y=0.715
c139 ( 51 0 ) capacitor c=0.0836807f //x=3.135 //y=1.92
c140 ( 50 0 ) capacitor c=0.0229722f //x=3.135 //y=1.525
c141 ( 49 0 ) capacitor c=0.0234352f //x=3.135 //y=1.215
c142 ( 48 0 ) capacitor c=0.0199366f //x=3.135 //y=0.87
c143 ( 47 0 ) capacitor c=0.0435629f //x=1.38 //y=1.255
c144 ( 46 0 ) capacitor c=0.0200386f //x=1.38 //y=0.91
c145 ( 40 0 ) capacitor c=0.0152946f //x=1.225 //y=1.41
c146 ( 38 0 ) capacitor c=0.0157804f //x=1.225 //y=0.755
c147 ( 37 0 ) capacitor c=0.048995f //x=0.97 //y=4.79
c148 ( 36 0 ) capacitor c=0.0303096f //x=1.26 //y=4.79
c149 ( 32 0 ) capacitor c=0.0290017f //x=0.85 //y=1.92
c150 ( 31 0 ) capacitor c=0.0250027f //x=0.85 //y=1.565
c151 ( 30 0 ) capacitor c=0.0234316f //x=0.85 //y=1.255
c152 ( 29 0 ) capacitor c=0.0200596f //x=0.85 //y=0.91
c153 ( 28 0 ) capacitor c=0.110797f //x=3.67 //y=6.02
c154 ( 27 0 ) capacitor c=0.154322f //x=3.23 //y=6.02
c155 ( 26 0 ) capacitor c=0.154218f //x=1.335 //y=6.02
c156 ( 25 0 ) capacitor c=0.154243f //x=0.895 //y=6.02
c157 ( 16 0 ) capacitor c=0.109612f //x=3.33 //y=2.085
c158 ( 8 0 ) capacitor c=0.11095f //x=0.74 //y=2.085
c159 ( 2 0 ) capacitor c=0.0144527f //x=0.855 //y=4.07
c160 ( 1 0 ) capacitor c=0.0971867f //x=3.215 //y=4.07
r161 (  78 80 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=3.23 //y=4.7 //x2=3.33 //y2=4.7
r162 (  66 67 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=0.74 //y=2.085 //x2=0.85 //y2=2.085
r163 (  62 80 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=3.67 //y=4.865 //x2=3.33 //y2=4.7
r164 (  61 82 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.665 //y=1.215 //x2=3.625 //y2=1.37
r165 (  60 81 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.665 //y=0.87 //x2=3.625 //y2=0.715
r166 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.665 //y=0.87 //x2=3.665 //y2=1.215
r167 (  58 77 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.29 //y=1.37 //x2=3.175 //y2=1.37
r168 (  57 82 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.51 //y=1.37 //x2=3.625 //y2=1.37
r169 (  56 76 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.29 //y=0.715 //x2=3.175 //y2=0.715
r170 (  55 81 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.51 //y=0.715 //x2=3.625 //y2=0.715
r171 (  55 56 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.51 //y=0.715 //x2=3.29 //y2=0.715
r172 (  52 78 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.23 //y=4.865 //x2=3.23 //y2=4.7
r173 (  51 75 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.92 //x2=3.33 //y2=2.085
r174 (  50 77 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.525 //x2=3.175 //y2=1.37
r175 (  50 51 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.525 //x2=3.135 //y2=1.92
r176 (  49 77 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.215 //x2=3.175 //y2=1.37
r177 (  48 76 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=0.87 //x2=3.175 //y2=0.715
r178 (  48 49 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.135 //y=0.87 //x2=3.135 //y2=1.215
r179 (  47 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=1.255 //x2=1.34 //y2=1.41
r180 (  46 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.34 //y2=0.755
r181 (  46 47 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.38 //y2=1.255
r182 (  41 71 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=1.41 //x2=0.89 //y2=1.41
r183 (  40 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=1.41 //x2=1.34 //y2=1.41
r184 (  39 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=0.755 //x2=0.89 //y2=0.755
r185 (  38 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.34 //y2=0.755
r186 (  38 39 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.005 //y2=0.755
r187 (  36 43 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=1.335 //y2=4.865
r188 (  36 37 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=0.97 //y2=4.79
r189 (  33 37 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.97 //y2=4.79
r190 (  33 69 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.74 //y2=4.7
r191 (  32 67 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.92 //x2=0.85 //y2=2.085
r192 (  31 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.89 //y2=1.41
r193 (  31 32 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.85 //y2=1.92
r194 (  30 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.255 //x2=0.89 //y2=1.41
r195 (  29 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.89 //y2=0.755
r196 (  29 30 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.85 //y2=1.255
r197 (  28 62 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.67 //y=6.02 //x2=3.67 //y2=4.865
r198 (  27 52 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.23 //y=6.02 //x2=3.23 //y2=4.865
r199 (  26 43 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.335 //y=6.02 //x2=1.335 //y2=4.865
r200 (  25 33 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.895 //y=6.02 //x2=0.895 //y2=4.865
r201 (  24 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.4 //y=1.37 //x2=3.51 //y2=1.37
r202 (  24 58 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.4 //y=1.37 //x2=3.29 //y2=1.37
r203 (  23 40 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.225 //y2=1.41
r204 (  23 41 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.005 //y2=1.41
r205 (  21 80 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r206 (  19 21 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=3.33 //y=4.07 //x2=3.33 //y2=4.7
r207 (  16 75 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.085 //x2=3.33 //y2=2.085
r208 (  16 19 ) resistor r=135.872 //w=0.187 //l=1.985 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.085 //x2=3.33 //y2=4.07
r209 (  13 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.7 //x2=0.74 //y2=4.7
r210 (  11 13 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=0.74 //y=4.07 //x2=0.74 //y2=4.7
r211 (  8 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=2.085
r212 (  8 11 ) resistor r=135.872 //w=0.187 //l=1.985 //layer=li \
 //thickness=0.1 //x=0.74 //y=2.085 //x2=0.74 //y2=4.07
r213 (  6 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=4.07 //x2=3.33 //y2=4.07
r214 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=0.74 //y=4.07 //x2=0.74 //y2=4.07
r215 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=0.855 //y=4.07 //x2=0.74 //y2=4.07
r216 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.215 //y=4.07 //x2=3.33 //y2=4.07
r217 (  1 2 ) resistor r=2.25191 //w=0.131 //l=2.36 //layer=m1 \
 //thickness=0.36 //x=3.215 //y=4.07 //x2=0.855 //y2=4.07
ends PM_XOR2X1_PCELL\%noxref_3

subckt PM_XOR2X1_PCELL\%noxref_4 ( 1 2 17 18 19 20 24 26 33 34 35 36 37 38 39 \
 43 45 51 52 60 62 64 )
c169 ( 64 0 ) capacitor c=0.0288629f //x=0.97 //y=5.02
c170 ( 62 0 ) capacitor c=0.0173218f //x=0.925 //y=0.91
c171 ( 60 0 ) capacitor c=0.058481f //x=7.77 //y=4.7
c172 ( 52 0 ) capacitor c=0.0417768f //x=7.965 //y=1.255
c173 ( 51 0 ) capacitor c=0.0192208f //x=7.965 //y=0.91
c174 ( 45 0 ) capacitor c=0.0124204f //x=7.81 //y=1.41
c175 ( 43 0 ) capacitor c=0.0157803f //x=7.81 //y=0.755
c176 ( 39 0 ) capacitor c=0.0903287f //x=7.435 //y=1.92
c177 ( 38 0 ) capacitor c=0.0194674f //x=7.435 //y=1.565
c178 ( 37 0 ) capacitor c=0.0168481f //x=7.435 //y=1.255
c179 ( 36 0 ) capacitor c=0.0174345f //x=7.435 //y=0.91
c180 ( 35 0 ) capacitor c=0.153255f //x=7.88 //y=6.02
c181 ( 34 0 ) capacitor c=0.110227f //x=7.44 //y=6.02
c182 ( 26 0 ) capacitor c=0.0737449f //x=7.77 //y=2.085
c183 ( 24 0 ) capacitor c=0.0868472f //x=1.48 //y=2.59
c184 ( 20 0 ) capacitor c=0.00417404f //x=1.2 //y=4.58
c185 ( 19 0 ) capacitor c=0.0118896f //x=1.395 //y=4.58
c186 ( 18 0 ) capacitor c=0.00621372f //x=1.195 //y=2.08
c187 ( 17 0 ) capacitor c=0.013454f //x=1.395 //y=2.08
c188 ( 2 0 ) capacitor c=0.0163395f //x=1.595 //y=2.59
c189 ( 1 0 ) capacitor c=0.188407f //x=7.655 //y=2.59
r190 (  60 61 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.77 //y=4.7 //x2=7.88 //y2=4.7
r191 (  52 58 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.965 //y=1.255 //x2=7.925 //y2=1.41
r192 (  51 57 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.965 //y=0.91 //x2=7.925 //y2=0.755
r193 (  51 52 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.965 //y=0.91 //x2=7.965 //y2=1.255
r194 (  48 61 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=7.88 //y=4.865 //x2=7.88 //y2=4.7
r195 (  46 54 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.59 //y=1.41 //x2=7.475 //y2=1.41
r196 (  45 58 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.81 //y=1.41 //x2=7.925 //y2=1.41
r197 (  44 53 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.59 //y=0.755 //x2=7.475 //y2=0.755
r198 (  43 57 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.81 //y=0.755 //x2=7.925 //y2=0.755
r199 (  43 44 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.81 //y=0.755 //x2=7.59 //y2=0.755
r200 (  40 60 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=7.44 //y=4.865 //x2=7.77 //y2=4.7
r201 (  39 56 ) resistor r=67.2792 //w=0.24 //l=0.438891 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.92 //x2=7.77 //y2=2.16
r202 (  38 54 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.565 //x2=7.475 //y2=1.41
r203 (  38 39 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.565 //x2=7.435 //y2=1.92
r204 (  37 54 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.255 //x2=7.475 //y2=1.41
r205 (  36 53 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.435 //y=0.91 //x2=7.475 //y2=0.755
r206 (  36 37 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.435 //y=0.91 //x2=7.435 //y2=1.255
r207 (  35 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.88 //y=6.02 //x2=7.88 //y2=4.865
r208 (  34 40 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.44 //y=6.02 //x2=7.44 //y2=4.865
r209 (  33 45 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.7 //y=1.41 //x2=7.81 //y2=1.41
r210 (  33 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.7 //y=1.41 //x2=7.59 //y2=1.41
r211 (  31 60 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.77 //y=4.7 //x2=7.77 //y2=4.7
r212 (  29 31 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=7.77 //y=2.59 //x2=7.77 //y2=4.7
r213 (  26 56 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.77 //y=2.085 //x2=7.77 //y2=2.085
r214 (  26 29 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=7.77 //y=2.085 //x2=7.77 //y2=2.59
r215 (  22 24 ) resistor r=130.396 //w=0.187 //l=1.905 //layer=li \
 //thickness=0.1 //x=1.48 //y=4.495 //x2=1.48 //y2=2.59
r216 (  21 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.48 //y=2.165 //x2=1.48 //y2=2.59
r217 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.48 //y2=4.495
r218 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.2 //y2=4.58
r219 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.48 //y2=2.165
r220 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.195 //y2=2.08
r221 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.2 //y2=4.58
r222 (  11 64 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.115 //y2=5.725
r223 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.195 //y2=2.08
r224 (  7 62 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.11 //y2=1.005
r225 (  6 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.77 //y=2.59 //x2=7.77 //y2=2.59
r226 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.48 //y=2.59 //x2=1.48 //y2=2.59
r227 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.595 //y=2.59 //x2=1.48 //y2=2.59
r228 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.655 //y=2.59 //x2=7.77 //y2=2.59
r229 (  1 2 ) resistor r=5.78244 //w=0.131 //l=6.06 //layer=m1 \
 //thickness=0.36 //x=7.655 //y=2.59 //x2=1.595 //y2=2.59
ends PM_XOR2X1_PCELL\%noxref_4

subckt PM_XOR2X1_PCELL\%noxref_5 ( 1 2 17 18 19 20 24 35 36 37 38 42 43 44 47 \
 48 )
c149 ( 48 0 ) capacitor c=0.0159588f //x=7.515 //y=5.02
c150 ( 47 0 ) capacitor c=0.0159588f //x=4.185 //y=5.02
c151 ( 44 0 ) capacitor c=0.00827922f //x=7.51 //y=0.91
c152 ( 43 0 ) capacitor c=0.00846882f //x=4.18 //y=0.91
c153 ( 42 0 ) capacitor c=0.0892717f //x=8.14 //y=3.7
c154 ( 38 0 ) capacitor c=0.00178322f //x=7.785 //y=1.655
c155 ( 37 0 ) capacitor c=0.0112025f //x=8.055 //y=1.655
c156 ( 36 0 ) capacitor c=0.00235465f //x=7.745 //y=5.205
c157 ( 35 0 ) capacitor c=0.0121398f //x=8.055 //y=5.205
c158 ( 24 0 ) capacitor c=0.10559f //x=4.81 //y=3.7
c159 ( 20 0 ) capacitor c=0.00178606f //x=4.455 //y=1.655
c160 ( 19 0 ) capacitor c=0.0109582f //x=4.725 //y=1.655
c161 ( 18 0 ) capacitor c=0.0027221f //x=4.415 //y=5.205
c162 ( 17 0 ) capacitor c=0.0121701f //x=4.725 //y=5.205
c163 ( 2 0 ) capacitor c=0.0132457f //x=4.925 //y=3.7
c164 ( 1 0 ) capacitor c=0.0664267f //x=8.025 //y=3.7
r165 (  40 42 ) resistor r=97.1979 //w=0.187 //l=1.42 //layer=li \
 //thickness=0.1 //x=8.14 //y=5.12 //x2=8.14 //y2=3.7
r166 (  39 42 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=8.14 //y=1.74 //x2=8.14 //y2=3.7
r167 (  37 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.055 //y=1.655 //x2=8.14 //y2=1.74
r168 (  37 38 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=8.055 //y=1.655 //x2=7.785 //y2=1.655
r169 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.055 //y=5.205 //x2=8.14 //y2=5.12
r170 (  35 36 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=8.055 //y=5.205 //x2=7.745 //y2=5.205
r171 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.7 //y=1.57 //x2=7.785 //y2=1.655
r172 (  31 44 ) resistor r=38.6738 //w=0.187 //l=0.565 //layer=li \
 //thickness=0.1 //x=7.7 //y=1.57 //x2=7.7 //y2=1.005
r173 (  25 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.66 //y=5.29 //x2=7.745 //y2=5.205
r174 (  25 48 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=7.66 //y=5.29 //x2=7.66 //y2=5.715
r175 (  22 24 ) resistor r=97.1979 //w=0.187 //l=1.42 //layer=li \
 //thickness=0.1 //x=4.81 //y=5.12 //x2=4.81 //y2=3.7
r176 (  21 24 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=4.81 //y=1.74 //x2=4.81 //y2=3.7
r177 (  19 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=1.655 //x2=4.81 //y2=1.74
r178 (  19 20 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=4.725 //y=1.655 //x2=4.455 //y2=1.655
r179 (  17 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=5.205 //x2=4.81 //y2=5.12
r180 (  17 18 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=4.725 //y=5.205 //x2=4.415 //y2=5.205
r181 (  13 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.37 //y=1.57 //x2=4.455 //y2=1.655
r182 (  13 43 ) resistor r=38.6738 //w=0.187 //l=0.565 //layer=li \
 //thickness=0.1 //x=4.37 //y=1.57 //x2=4.37 //y2=1.005
r183 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.33 //y=5.29 //x2=4.415 //y2=5.205
r184 (  7 47 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=4.33 //y=5.29 //x2=4.33 //y2=5.715
r185 (  6 42 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.14 //y=3.7 //x2=8.14 //y2=3.7
r186 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.81 //y=3.7 //x2=4.81 //y2=3.7
r187 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.925 //y=3.7 //x2=4.81 //y2=3.7
r188 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.025 //y=3.7 //x2=8.14 //y2=3.7
r189 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=8.025 //y=3.7 //x2=4.925 //y2=3.7
ends PM_XOR2X1_PCELL\%noxref_5

subckt PM_XOR2X1_PCELL\%noxref_6 ( 1 2 3 4 14 20 28 31 32 33 34 45 46 47 54 55 \
 56 57 58 60 63 64 66 74 76 )
c165 ( 76 0 ) capacitor c=0.028734f //x=9.84 //y=5.02
c166 ( 74 0 ) capacitor c=0.0173218f //x=9.795 //y=0.91
c167 ( 66 0 ) capacitor c=0.0636249f //x=4.44 //y=4.7
c168 ( 64 0 ) capacitor c=0.0318948f //x=6.995 //y=1.215
c169 ( 63 0 ) capacitor c=0.0187407f //x=6.995 //y=0.87
c170 ( 60 0 ) capacitor c=0.0141798f //x=6.84 //y=1.37
c171 ( 58 0 ) capacitor c=0.0149852f //x=6.84 //y=0.715
c172 ( 57 0 ) capacitor c=0.0836807f //x=6.465 //y=1.92
c173 ( 56 0 ) capacitor c=0.0229722f //x=6.465 //y=1.525
c174 ( 55 0 ) capacitor c=0.0234352f //x=6.465 //y=1.215
c175 ( 54 0 ) capacitor c=0.0199366f //x=6.465 //y=0.87
c176 ( 47 0 ) capacitor c=0.153255f //x=4.55 //y=6.02
c177 ( 46 0 ) capacitor c=0.110227f //x=4.11 //y=6.02
c178 ( 34 0 ) capacitor c=0.00670488f //x=9.705 //y=4.58
c179 ( 33 0 ) capacitor c=0.0137356f //x=9.9 //y=4.58
c180 ( 32 0 ) capacitor c=0.00580686f //x=9.705 //y=2.08
c181 ( 31 0 ) capacitor c=0.0128831f //x=9.905 //y=2.08
c182 ( 28 0 ) capacitor c=0.0775792f //x=9.62 //y=3.33
c183 ( 20 0 ) capacitor c=0.0551449f //x=6.66 //y=2.085
c184 ( 14 0 ) capacitor c=0.024985f //x=4.44 //y=4.07
c185 ( 4 0 ) capacitor c=0.0126928f //x=6.775 //y=3.33
c186 ( 3 0 ) capacitor c=0.0544915f //x=9.505 //y=3.33
c187 ( 2 0 ) capacitor c=0.01091f //x=4.555 //y=4.07
c188 ( 1 0 ) capacitor c=0.109416f //x=9.505 //y=4.07
r189 (  66 67 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.44 //y=4.7 //x2=4.55 //y2=4.7
r190 (  64 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.995 //y=1.215 //x2=6.955 //y2=1.37
r191 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.995 //y=0.87 //x2=6.955 //y2=0.715
r192 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.995 //y=0.87 //x2=6.995 //y2=1.215
r193 (  61 71 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.62 //y=1.37 //x2=6.505 //y2=1.37
r194 (  60 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.84 //y=1.37 //x2=6.955 //y2=1.37
r195 (  59 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.62 //y=0.715 //x2=6.505 //y2=0.715
r196 (  58 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.84 //y=0.715 //x2=6.955 //y2=0.715
r197 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.84 //y=0.715 //x2=6.62 //y2=0.715
r198 (  57 69 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.92 //x2=6.66 //y2=2.085
r199 (  56 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.525 //x2=6.505 //y2=1.37
r200 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.525 //x2=6.465 //y2=1.92
r201 (  55 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.215 //x2=6.505 //y2=1.37
r202 (  54 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.465 //y=0.87 //x2=6.505 //y2=0.715
r203 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.465 //y=0.87 //x2=6.465 //y2=1.215
r204 (  51 67 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=4.55 //y=4.865 //x2=4.55 //y2=4.7
r205 (  48 66 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=4.11 //y=4.865 //x2=4.44 //y2=4.7
r206 (  47 51 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.55 //y=6.02 //x2=4.55 //y2=4.865
r207 (  46 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.11 //y=6.02 //x2=4.11 //y2=4.865
r208 (  45 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.73 //y=1.37 //x2=6.84 //y2=1.37
r209 (  45 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.73 //y=1.37 //x2=6.62 //y2=1.37
r210 (  41 74 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=9.99 //y=1.995 //x2=9.99 //y2=1.005
r211 (  35 76 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=9.985 //y=4.665 //x2=9.985 //y2=5.725
r212 (  33 35 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.9 //y=4.58 //x2=9.985 //y2=4.665
r213 (  33 34 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=9.9 //y=4.58 //x2=9.705 //y2=4.58
r214 (  31 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.905 //y=2.08 //x2=9.99 //y2=1.995
r215 (  31 32 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=9.905 //y=2.08 //x2=9.705 //y2=2.08
r216 (  28 30 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=9.62 //y=3.33 //x2=9.62 //y2=4.07
r217 (  26 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.62 //y=4.495 //x2=9.705 //y2=4.58
r218 (  26 30 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=9.62 //y=4.495 //x2=9.62 //y2=4.07
r219 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.62 //y=2.165 //x2=9.705 //y2=2.08
r220 (  25 28 ) resistor r=79.7433 //w=0.187 //l=1.165 //layer=li \
 //thickness=0.1 //x=9.62 //y=2.165 //x2=9.62 //y2=3.33
r221 (  20 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.085 //x2=6.66 //y2=2.085
r222 (  20 23 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.085 //x2=6.66 //y2=3.33
r223 (  17 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=4.7 //x2=4.44 //y2=4.7
r224 (  14 17 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=4.44 //y=4.07 //x2=4.44 //y2=4.7
r225 (  12 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.62 //y=4.07 //x2=9.62 //y2=4.07
r226 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.62 //y=3.33 //x2=9.62 //y2=3.33
r227 (  8 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=3.33 //x2=6.66 //y2=3.33
r228 (  6 14 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=4.07 //x2=4.44 //y2=4.07
r229 (  4 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.775 //y=3.33 //x2=6.66 //y2=3.33
r230 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=3.33 //x2=9.62 //y2=3.33
r231 (  3 4 ) resistor r=2.60496 //w=0.131 //l=2.73 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=3.33 //x2=6.775 //y2=3.33
r232 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.555 //y=4.07 //x2=4.44 //y2=4.07
r233 (  1 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=4.07 //x2=9.62 //y2=4.07
r234 (  1 2 ) resistor r=4.72328 //w=0.131 //l=4.95 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=4.07 //x2=4.555 //y2=4.07
ends PM_XOR2X1_PCELL\%noxref_6

subckt PM_XOR2X1_PCELL\%noxref_7 ( 1 2 3 4 14 20 26 35 36 37 38 39 40 41 42 43 \
 44 45 47 50 51 58 59 63 64 65 67 70 73 74 75 76 85 90 )
c173 ( 90 0 ) capacitor c=0.051138f //x=10.25 //y=2.085
c174 ( 85 0 ) capacitor c=0.0606915f //x=6.66 //y=4.7
c175 ( 76 0 ) capacitor c=0.0290017f //x=10.25 //y=1.92
c176 ( 75 0 ) capacitor c=0.0250171f //x=10.25 //y=1.565
c177 ( 74 0 ) capacitor c=0.0234316f //x=10.25 //y=1.255
c178 ( 73 0 ) capacitor c=0.0200712f //x=10.25 //y=0.91
c179 ( 70 0 ) capacitor c=0.0488625f //x=10.205 //y=4.865
c180 ( 67 0 ) capacitor c=0.0152946f //x=10.095 //y=1.41
c181 ( 65 0 ) capacitor c=0.0157804f //x=10.095 //y=0.755
c182 ( 64 0 ) capacitor c=0.0129718f //x=9.84 //y=4.79
c183 ( 63 0 ) capacitor c=0.0172687f //x=10.13 //y=4.79
c184 ( 59 0 ) capacitor c=0.0435512f //x=9.72 //y=1.255
c185 ( 58 0 ) capacitor c=0.0200269f //x=9.72 //y=0.91
c186 ( 51 0 ) capacitor c=0.0417768f //x=4.635 //y=1.255
c187 ( 50 0 ) capacitor c=0.0192208f //x=4.635 //y=0.91
c188 ( 47 0 ) capacitor c=0.0124204f //x=4.48 //y=1.41
c189 ( 45 0 ) capacitor c=0.0157803f //x=4.48 //y=0.755
c190 ( 44 0 ) capacitor c=0.0903325f //x=4.105 //y=1.92
c191 ( 43 0 ) capacitor c=0.0194674f //x=4.105 //y=1.565
c192 ( 42 0 ) capacitor c=0.0168481f //x=4.105 //y=1.255
c193 ( 41 0 ) capacitor c=0.0174345f //x=4.105 //y=0.91
c194 ( 40 0 ) capacitor c=0.154243f //x=10.205 //y=6.02
c195 ( 39 0 ) capacitor c=0.154218f //x=9.765 //y=6.02
c196 ( 38 0 ) capacitor c=0.110797f //x=7 //y=6.02
c197 ( 37 0 ) capacitor c=0.154322f //x=6.56 //y=6.02
c198 ( 26 0 ) capacitor c=0.106666f //x=10.36 //y=2.085
c199 ( 20 0 ) capacitor c=0.0150587f //x=6.66 //y=4.44
c200 ( 14 0 ) capacitor c=0.0306114f //x=4.44 //y=2.085
c201 ( 4 0 ) capacitor c=0.015004f //x=6.775 //y=4.44
c202 ( 3 0 ) capacitor c=0.0929962f //x=10.245 //y=4.44
c203 ( 2 0 ) capacitor c=0.0154186f //x=4.555 //y=2.96
c204 ( 1 0 ) capacitor c=0.130205f //x=10.245 //y=2.96
r205 (  90 92 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.25 //y=2.085 //x2=10.36 //y2=2.085
r206 (  83 85 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=6.56 //y=4.7 //x2=6.66 //y2=4.7
r207 (  76 90 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=10.25 //y=1.92 //x2=10.25 //y2=2.085
r208 (  75 89 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.25 //y=1.565 //x2=10.21 //y2=1.41
r209 (  75 76 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=10.25 //y=1.565 //x2=10.25 //y2=1.92
r210 (  74 89 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.25 //y=1.255 //x2=10.21 //y2=1.41
r211 (  73 88 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.25 //y=0.91 //x2=10.21 //y2=0.755
r212 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.25 //y=0.91 //x2=10.25 //y2=1.255
r213 (  70 94 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=10.205 //y=4.865 //x2=10.36 //y2=4.7
r214 (  68 87 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.875 //y=1.41 //x2=9.76 //y2=1.41
r215 (  67 89 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.095 //y=1.41 //x2=10.21 //y2=1.41
r216 (  66 86 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.875 //y=0.755 //x2=9.76 //y2=0.755
r217 (  65 88 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.095 //y=0.755 //x2=10.21 //y2=0.755
r218 (  65 66 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.095 //y=0.755 //x2=9.875 //y2=0.755
r219 (  63 70 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.13 //y=4.79 //x2=10.205 //y2=4.865
r220 (  63 64 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=10.13 //y=4.79 //x2=9.84 //y2=4.79
r221 (  60 64 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.765 //y=4.865 //x2=9.84 //y2=4.79
r222 (  59 87 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.72 //y=1.255 //x2=9.76 //y2=1.41
r223 (  58 86 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.72 //y=0.91 //x2=9.76 //y2=0.755
r224 (  58 59 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.72 //y=0.91 //x2=9.72 //y2=1.255
r225 (  55 85 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=7 //y=4.865 //x2=6.66 //y2=4.7
r226 (  52 83 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.56 //y=4.865 //x2=6.56 //y2=4.7
r227 (  51 82 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.635 //y=1.255 //x2=4.595 //y2=1.41
r228 (  50 81 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.635 //y=0.91 //x2=4.595 //y2=0.755
r229 (  50 51 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.635 //y=0.91 //x2=4.635 //y2=1.255
r230 (  48 78 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.26 //y=1.41 //x2=4.145 //y2=1.41
r231 (  47 82 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.48 //y=1.41 //x2=4.595 //y2=1.41
r232 (  46 77 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.26 //y=0.755 //x2=4.145 //y2=0.755
r233 (  45 81 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.48 //y=0.755 //x2=4.595 //y2=0.755
r234 (  45 46 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.48 //y=0.755 //x2=4.26 //y2=0.755
r235 (  44 80 ) resistor r=67.2792 //w=0.24 //l=0.438891 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.92 //x2=4.44 //y2=2.16
r236 (  43 78 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.565 //x2=4.145 //y2=1.41
r237 (  43 44 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.565 //x2=4.105 //y2=1.92
r238 (  42 78 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.255 //x2=4.145 //y2=1.41
r239 (  41 77 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=0.91 //x2=4.145 //y2=0.755
r240 (  41 42 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.105 //y=0.91 //x2=4.105 //y2=1.255
r241 (  40 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.205 //y=6.02 //x2=10.205 //y2=4.865
r242 (  39 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.765 //y=6.02 //x2=9.765 //y2=4.865
r243 (  38 55 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7 //y=6.02 //x2=7 //y2=4.865
r244 (  37 52 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.56 //y=6.02 //x2=6.56 //y2=4.865
r245 (  36 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.985 //y=1.41 //x2=10.095 //y2=1.41
r246 (  36 68 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.985 //y=1.41 //x2=9.875 //y2=1.41
r247 (  35 47 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.37 //y=1.41 //x2=4.48 //y2=1.41
r248 (  35 48 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.37 //y=1.41 //x2=4.26 //y2=1.41
r249 (  33 94 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=4.7 //x2=10.36 //y2=4.7
r250 (  31 33 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=10.36 //y=4.44 //x2=10.36 //y2=4.7
r251 (  29 31 ) resistor r=101.305 //w=0.187 //l=1.48 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.96 //x2=10.36 //y2=4.44
r252 (  26 92 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=2.085 //x2=10.36 //y2=2.085
r253 (  26 29 ) resistor r=59.893 //w=0.187 //l=0.875 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.085 //x2=10.36 //y2=2.96
r254 (  23 85 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=4.7 //x2=6.66 //y2=4.7
r255 (  20 23 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=6.66 //y=4.44 //x2=6.66 //y2=4.7
r256 (  14 80 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=2.085 //x2=4.44 //y2=2.085
r257 (  14 17 ) resistor r=59.893 //w=0.187 //l=0.875 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.085 //x2=4.44 //y2=2.96
r258 (  12 31 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=4.44 //x2=10.36 //y2=4.44
r259 (  10 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=2.96 //x2=10.36 //y2=2.96
r260 (  8 20 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=4.44 //x2=6.66 //y2=4.44
r261 (  6 17 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=2.96 //x2=4.44 //y2=2.96
r262 (  4 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.775 //y=4.44 //x2=6.66 //y2=4.44
r263 (  3 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.245 //y=4.44 //x2=10.36 //y2=4.44
r264 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=10.245 //y=4.44 //x2=6.775 //y2=4.44
r265 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.555 //y=2.96 //x2=4.44 //y2=2.96
r266 (  1 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.245 //y=2.96 //x2=10.36 //y2=2.96
r267 (  1 2 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=10.245 //y=2.96 //x2=4.555 //y2=2.96
ends PM_XOR2X1_PCELL\%noxref_7

subckt PM_XOR2X1_PCELL\%noxref_8 ( 7 8 15 16 23 24 25 )
c40 ( 25 0 ) capacitor c=0.0306618f //x=4.625 //y=5.02
c41 ( 24 0 ) capacitor c=0.0185379f //x=3.745 //y=5.02
c42 ( 23 0 ) capacitor c=0.0384176f //x=2.875 //y=5.02
c43 ( 16 0 ) capacitor c=0.00194711f //x=3.975 //y=6.905
c44 ( 15 0 ) capacitor c=0.014216f //x=4.685 //y=6.905
c45 ( 8 0 ) capacitor c=0.00644339f //x=3.095 //y=5.205
c46 ( 7 0 ) capacitor c=0.0212224f //x=3.805 //y=5.205
r47 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.77 //y=6.82 //x2=4.77 //y2=6.735
r48 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.685 //y=6.905 //x2=4.77 //y2=6.82
r49 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=4.685 //y=6.905 //x2=3.975 //y2=6.905
r50 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.89 //y=6.82 //x2=3.975 //y2=6.905
r51 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=3.89 //y=6.82 //x2=3.89 //y2=6.395
r52 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=3.89 //y=5.29 //x2=3.89 //y2=5.715
r53 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.805 //y=5.205 //x2=3.89 //y2=5.29
r54 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=3.805 //y=5.205 //x2=3.095 //y2=5.205
r55 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.01 //y=5.29 //x2=3.095 //y2=5.205
r56 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=3.01 //y=5.29 //x2=3.01 //y2=5.715
ends PM_XOR2X1_PCELL\%noxref_8

subckt PM_XOR2X1_PCELL\%noxref_9 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632228f //x=2.78 //y=0.37
c53 ( 17 0 ) capacitor c=0.00723243f //x=4.855 //y=0.62
c54 ( 13 0 ) capacitor c=0.0153475f //x=4.77 //y=0.535
c55 ( 10 0 ) capacitor c=0.00656687f //x=3.885 //y=1.5
c56 ( 9 0 ) capacitor c=0.00677124f //x=3.885 //y=0.62
c57 ( 5 0 ) capacitor c=0.0181169f //x=3.8 //y=1.585
c58 ( 1 0 ) capacitor c=0.0076549f //x=2.915 //y=1.5
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.855 //y=0.62 //x2=4.855 //y2=0.495
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.855 //y=0.62 //x2=4.855 //y2=0.885
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.97 //y=0.535 //x2=3.885 //y2=0.495
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.97 //y=0.535 //x2=4.37 //y2=0.535
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.77 //y=0.535 //x2=4.855 //y2=0.495
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.77 //y=0.535 //x2=4.37 //y2=0.535
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=3.885 //y=1.5 //x2=3.885 //y2=1.625
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=3.885 //y=1.5 //x2=3.885 //y2=0.885
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.885 //y=0.62 //x2=3.885 //y2=0.495
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.885 //y=0.62 //x2=3.885 //y2=0.885
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3 //y=1.585 //x2=2.915 //y2=1.625
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3 //y=1.585 //x2=3.4 //y2=1.585
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.8 //y=1.585 //x2=3.885 //y2=1.625
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.8 //y=1.585 //x2=3.4 //y2=1.585
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=2.915 //y=1.5 //x2=2.915 //y2=1.625
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.915 //y=1.5 //x2=2.915 //y2=0.885
ends PM_XOR2X1_PCELL\%noxref_9

subckt PM_XOR2X1_PCELL\%noxref_10 ( 7 8 15 16 23 24 25 )
c43 ( 25 0 ) capacitor c=0.0305804f //x=7.955 //y=5.02
c44 ( 24 0 ) capacitor c=0.0185379f //x=7.075 //y=5.02
c45 ( 23 0 ) capacitor c=0.0384176f //x=6.205 //y=5.02
c46 ( 16 0 ) capacitor c=0.00194711f //x=7.305 //y=6.905
c47 ( 15 0 ) capacitor c=0.0133643f //x=8.015 //y=6.905
c48 ( 8 0 ) capacitor c=0.00631451f //x=6.425 //y=5.205
c49 ( 7 0 ) capacitor c=0.0183784f //x=7.135 //y=5.205
r50 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.1 //y=6.82 //x2=8.1 //y2=6.735
r51 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.015 //y=6.905 //x2=8.1 //y2=6.82
r52 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.015 //y=6.905 //x2=7.305 //y2=6.905
r53 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.22 //y=6.82 //x2=7.305 //y2=6.905
r54 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=7.22 //y=6.82 //x2=7.22 //y2=6.395
r55 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.29 //x2=7.22 //y2=5.715
r56 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.205 //x2=7.22 //y2=5.29
r57 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=7.135 //y=5.205 //x2=6.425 //y2=5.205
r58 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.29 //x2=6.425 //y2=5.205
r59 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.29 //x2=6.34 //y2=5.715
ends PM_XOR2X1_PCELL\%noxref_10

subckt PM_XOR2X1_PCELL\%noxref_11 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.063541f //x=6.11 //y=0.37
c54 ( 17 0 ) capacitor c=0.00723243f //x=8.185 //y=0.62
c55 ( 13 0 ) capacitor c=0.0153645f //x=8.1 //y=0.535
c56 ( 10 0 ) capacitor c=0.00656687f //x=7.215 //y=1.5
c57 ( 9 0 ) capacitor c=0.00677124f //x=7.215 //y=0.62
c58 ( 5 0 ) capacitor c=0.0181169f //x=7.13 //y=1.585
c59 ( 1 0 ) capacitor c=0.0076549f //x=6.245 //y=1.5
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.185 //y=0.62 //x2=8.185 //y2=0.495
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=8.185 //y=0.62 //x2=8.185 //y2=0.885
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.3 //y=0.535 //x2=7.215 //y2=0.495
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.3 //y=0.535 //x2=7.7 //y2=0.535
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.1 //y=0.535 //x2=8.185 //y2=0.495
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.1 //y=0.535 //x2=7.7 //y2=0.535
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.215 //y=1.5 //x2=7.215 //y2=1.625
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=7.215 //y=1.5 //x2=7.215 //y2=0.885
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.215 //y=0.62 //x2=7.215 //y2=0.495
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=7.215 //y=0.62 //x2=7.215 //y2=0.885
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.33 //y=1.585 //x2=6.245 //y2=1.625
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.33 //y=1.585 //x2=6.73 //y2=1.585
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.13 //y=1.585 //x2=7.215 //y2=1.625
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.13 //y=1.585 //x2=6.73 //y2=1.585
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.245 //y=1.5 //x2=6.245 //y2=1.625
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.245 //y=1.5 //x2=6.245 //y2=0.885
ends PM_XOR2X1_PCELL\%noxref_11

