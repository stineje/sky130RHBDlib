* SPICE3 file created from TIELO.ext - technology: sky130A

.subckt TIELO YN VDD VSS
X0 a_121_411 a_121_411 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.0011 ps=9.1 w=2 l=0.15 M=2
X1 YN a_121_411 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0.0011408 ps=8.1 w=3 l=0.15
.ends
