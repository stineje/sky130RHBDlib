* SPICE3 file created from VOTER3X1.ext - technology: sky130A

.subckt VOTER3X1 Y A B C VDD GND
X0 GND B voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X1 GND B voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X2 GND C voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X3 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# B VDD VDD pshort w=2 l=0.15
X4 voter3x1_pcell_0/m1_1867_797# C voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X5 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# A VDD VDD pshort w=2 l=0.15
X6 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# C voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X7 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# B voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X8 voter3x1_pcell_0/m1_1867_797# C voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X9 voter3x1_pcell_0/m1_1867_797# A voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X10 voter3x1_pcell_0/m1_1867_797# A voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X11 voter3x1_pcell_0/m1_1867_797# A voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X12 Y voter3x1_pcell_0/m1_1867_797# GND GND nshort w=3 l=0.15
X13 VDD voter3x1_pcell_0/m1_1867_797# Y VDD pshort w=2 l=0.15
C0 VDD GND 17.75fF
.ends
