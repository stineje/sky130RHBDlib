magic
tech sky130A
magscale 1 2
timestamp 1669564280
<< nwell >>
rect -87 786 4971 1550
<< pwell >>
rect -34 -34 4918 544
<< nmos >>
rect 168 288 198 349
tri 198 288 214 304 sw
rect 362 296 392 349
tri 392 296 408 312 sw
rect 168 258 274 288
tri 274 258 304 288 sw
rect 362 266 468 296
tri 468 266 498 296 sw
rect 168 157 198 258
tri 198 242 214 258 nw
tri 258 242 274 258 ne
tri 198 157 214 173 sw
tri 258 157 274 173 se
rect 274 157 304 258
rect 362 165 392 266
tri 392 250 408 266 nw
tri 452 250 468 266 ne
tri 392 165 408 181 sw
tri 452 165 468 181 se
rect 468 165 498 266
tri 168 127 198 157 ne
rect 198 127 274 157
tri 274 127 304 157 nw
tri 362 135 392 165 ne
rect 392 135 468 165
tri 468 135 498 165 nw
rect 813 290 843 351
tri 843 290 859 306 sw
rect 1113 290 1143 351
rect 813 260 919 290
tri 919 260 949 290 sw
rect 813 159 843 260
tri 843 244 859 260 nw
tri 903 244 919 260 ne
tri 843 159 859 175 sw
tri 903 159 919 175 se
rect 919 159 949 260
tri 1008 260 1038 290 se
rect 1038 260 1143 290
rect 1008 166 1038 260
tri 1038 244 1054 260 nw
tri 1097 244 1113 260 ne
tri 1038 166 1054 182 sw
tri 1097 166 1113 182 se
rect 1113 166 1143 260
tri 813 129 843 159 ne
rect 843 129 919 159
tri 919 129 949 159 nw
tri 1008 136 1038 166 ne
rect 1038 136 1113 166
tri 1113 136 1143 166 nw
rect 1315 298 1345 351
tri 1345 298 1361 314 sw
rect 1315 268 1421 298
tri 1421 268 1451 298 sw
rect 1315 167 1345 268
tri 1345 252 1361 268 nw
tri 1405 252 1421 268 ne
tri 1345 167 1361 183 sw
tri 1405 167 1421 183 se
rect 1421 167 1451 268
tri 1315 137 1345 167 ne
rect 1345 137 1421 167
tri 1421 137 1451 167 nw
rect 1775 290 1805 351
tri 1805 290 1821 306 sw
rect 2075 290 2105 351
rect 1775 260 1881 290
tri 1881 260 1911 290 sw
rect 1775 159 1805 260
tri 1805 244 1821 260 nw
tri 1865 244 1881 260 ne
tri 1805 159 1821 175 sw
tri 1865 159 1881 175 se
rect 1881 159 1911 260
tri 1970 260 2000 290 se
rect 2000 260 2105 290
rect 1970 166 2000 260
tri 2000 244 2016 260 nw
tri 2059 244 2075 260 ne
tri 2000 166 2016 182 sw
tri 2059 166 2075 182 se
rect 2075 166 2105 260
tri 1775 129 1805 159 ne
rect 1805 129 1881 159
tri 1881 129 1911 159 nw
tri 1970 136 2000 166 ne
rect 2000 136 2075 166
tri 2075 136 2105 166 nw
rect 2277 298 2307 351
tri 2307 298 2323 314 sw
rect 2277 268 2383 298
tri 2383 268 2413 298 sw
rect 2277 167 2307 268
tri 2307 252 2323 268 nw
tri 2367 252 2383 268 ne
tri 2307 167 2323 183 sw
tri 2367 167 2383 183 se
rect 2383 167 2413 268
tri 2277 137 2307 167 ne
rect 2307 137 2383 167
tri 2383 137 2413 167 nw
rect 2758 288 2788 349
tri 2788 288 2804 304 sw
rect 2952 296 2982 349
tri 2982 296 2998 312 sw
rect 2758 258 2864 288
tri 2864 258 2894 288 sw
rect 2952 266 3058 296
tri 3058 266 3088 296 sw
rect 2758 157 2788 258
tri 2788 242 2804 258 nw
tri 2848 242 2864 258 ne
tri 2788 157 2804 173 sw
tri 2848 157 2864 173 se
rect 2864 157 2894 258
rect 2952 165 2982 266
tri 2982 250 2998 266 nw
tri 3042 250 3058 266 ne
tri 2982 165 2998 181 sw
tri 3042 165 3058 181 se
rect 3058 165 3088 266
tri 2758 127 2788 157 ne
rect 2788 127 2864 157
tri 2864 127 2894 157 nw
tri 2952 135 2982 165 ne
rect 2982 135 3058 165
tri 3058 135 3088 165 nw
rect 3424 288 3454 349
tri 3454 288 3470 304 sw
rect 3618 296 3648 349
tri 3648 296 3664 312 sw
rect 3424 258 3530 288
tri 3530 258 3560 288 sw
rect 3618 266 3724 296
tri 3724 266 3754 296 sw
rect 3424 157 3454 258
tri 3454 242 3470 258 nw
tri 3514 242 3530 258 ne
tri 3454 157 3470 173 sw
tri 3514 157 3530 173 se
rect 3530 157 3560 258
rect 3618 165 3648 266
tri 3648 250 3664 266 nw
tri 3708 250 3724 266 ne
tri 3648 165 3664 181 sw
tri 3708 165 3724 181 se
rect 3724 165 3754 266
tri 3424 127 3454 157 ne
rect 3454 127 3530 157
tri 3530 127 3560 157 nw
tri 3618 135 3648 165 ne
rect 3648 135 3724 165
tri 3724 135 3754 165 nw
rect 4069 290 4099 351
tri 4099 290 4115 306 sw
rect 4369 290 4399 351
rect 4069 260 4175 290
tri 4175 260 4205 290 sw
rect 4069 159 4099 260
tri 4099 244 4115 260 nw
tri 4159 244 4175 260 ne
tri 4099 159 4115 175 sw
tri 4159 159 4175 175 se
rect 4175 159 4205 260
tri 4264 260 4294 290 se
rect 4294 260 4399 290
rect 4264 166 4294 260
tri 4294 244 4310 260 nw
tri 4353 244 4369 260 ne
tri 4294 166 4310 182 sw
tri 4353 166 4369 182 se
rect 4369 166 4399 260
tri 4069 129 4099 159 ne
rect 4099 129 4175 159
tri 4175 129 4205 159 nw
tri 4264 136 4294 166 ne
rect 4294 136 4369 166
tri 4369 136 4399 166 nw
rect 4571 298 4601 351
tri 4601 298 4617 314 sw
rect 4571 268 4677 298
tri 4677 268 4707 298 sw
rect 4571 167 4601 268
tri 4601 252 4617 268 nw
tri 4661 252 4677 268 ne
tri 4601 167 4617 183 sw
tri 4661 167 4677 183 se
rect 4677 167 4707 268
tri 4571 137 4601 167 ne
rect 4601 137 4677 167
tri 4677 137 4707 167 nw
<< pmos >>
rect 187 1004 217 1404
rect 275 1004 305 1404
rect 363 1004 393 1404
rect 451 1004 481 1404
rect 913 1004 943 1404
rect 1001 1004 1031 1404
rect 1089 1004 1119 1404
rect 1177 1004 1207 1404
rect 1265 1004 1295 1404
rect 1353 1004 1383 1404
rect 1875 1004 1905 1404
rect 1963 1004 1993 1404
rect 2051 1004 2081 1404
rect 2139 1004 2169 1404
rect 2227 1004 2257 1404
rect 2315 1004 2345 1404
rect 2777 1004 2807 1404
rect 2865 1004 2895 1404
rect 2953 1004 2983 1404
rect 3041 1004 3071 1404
rect 3443 1004 3473 1404
rect 3531 1004 3561 1404
rect 3619 1004 3649 1404
rect 3707 1004 3737 1404
rect 4169 1004 4199 1404
rect 4257 1004 4287 1404
rect 4345 1004 4375 1404
rect 4433 1004 4463 1404
rect 4521 1004 4551 1404
rect 4609 1004 4639 1404
<< ndiff >>
rect 112 333 168 349
rect 112 299 122 333
rect 156 299 168 333
rect 112 261 168 299
rect 198 333 362 349
rect 198 304 219 333
tri 198 288 214 304 ne
rect 214 299 219 304
rect 253 299 316 333
rect 350 299 362 333
rect 214 288 362 299
rect 392 312 554 349
tri 392 296 408 312 ne
rect 408 296 554 312
rect 112 227 122 261
rect 156 227 168 261
tri 274 258 304 288 ne
rect 304 261 362 288
tri 468 266 498 296 ne
rect 112 193 168 227
rect 112 159 122 193
rect 156 159 168 193
rect 112 127 168 159
tri 198 242 214 258 se
rect 214 242 258 258
tri 258 242 274 258 sw
rect 198 208 274 242
rect 198 174 219 208
rect 253 174 274 208
rect 198 173 274 174
tri 198 157 214 173 ne
rect 214 157 258 173
tri 258 157 274 173 nw
rect 304 227 316 261
rect 350 227 362 261
rect 304 193 362 227
rect 304 159 316 193
rect 350 159 362 193
tri 392 250 408 266 se
rect 408 250 452 266
tri 452 250 468 266 sw
rect 392 217 468 250
rect 392 183 413 217
rect 447 183 468 217
rect 392 181 468 183
tri 392 165 408 181 ne
rect 408 165 452 181
tri 452 165 468 181 nw
rect 498 261 554 296
rect 498 227 510 261
rect 544 227 554 261
rect 498 193 554 227
tri 168 127 198 157 sw
tri 274 127 304 157 se
rect 304 135 362 159
tri 362 135 392 165 sw
tri 468 135 498 165 se
rect 498 159 510 193
rect 544 159 554 193
rect 498 135 554 159
rect 304 127 554 135
rect 112 123 554 127
rect 112 89 122 123
rect 156 89 316 123
rect 350 89 413 123
rect 447 89 510 123
rect 544 89 554 123
rect 112 73 554 89
rect 757 335 813 351
rect 757 301 767 335
rect 801 301 813 335
rect 757 263 813 301
rect 843 335 1113 351
rect 843 306 864 335
tri 843 290 859 306 ne
rect 859 301 864 306
rect 898 301 961 335
rect 995 301 1058 335
rect 1092 301 1113 335
rect 859 290 1113 301
rect 1143 335 1199 351
rect 1143 301 1155 335
rect 1189 301 1199 335
rect 757 229 767 263
rect 801 229 813 263
tri 919 260 949 290 ne
rect 949 263 1008 290
rect 757 195 813 229
rect 757 161 767 195
rect 801 161 813 195
rect 757 129 813 161
tri 843 244 859 260 se
rect 859 244 903 260
tri 903 244 919 260 sw
rect 843 210 919 244
rect 843 176 864 210
rect 898 176 919 210
rect 843 175 919 176
tri 843 159 859 175 ne
rect 859 159 903 175
tri 903 159 919 175 nw
rect 949 229 961 263
rect 995 229 1008 263
tri 1008 260 1038 290 nw
rect 949 195 1008 229
rect 949 161 961 195
rect 995 161 1008 195
tri 1038 244 1054 260 se
rect 1054 244 1097 260
tri 1097 244 1113 260 sw
rect 1038 216 1113 244
rect 1038 182 1059 216
rect 1093 182 1113 216
tri 1038 166 1054 182 ne
rect 1054 166 1097 182
tri 1097 166 1113 182 nw
tri 813 129 843 159 sw
tri 919 129 949 159 se
rect 949 136 1008 161
tri 1008 136 1038 166 sw
tri 1113 136 1143 166 se
rect 1143 136 1199 301
rect 949 129 1199 136
rect 757 125 1199 129
rect 757 91 767 125
rect 801 91 961 125
rect 995 91 1058 125
rect 1092 91 1155 125
rect 1189 91 1199 125
rect 757 75 1199 91
rect 1259 335 1315 351
rect 1259 301 1269 335
rect 1303 301 1315 335
rect 1259 263 1315 301
rect 1345 314 1507 351
tri 1345 298 1361 314 ne
rect 1361 298 1507 314
tri 1421 268 1451 298 ne
rect 1259 229 1269 263
rect 1303 229 1315 263
rect 1259 195 1315 229
rect 1259 161 1269 195
rect 1303 161 1315 195
tri 1345 252 1361 268 se
rect 1361 252 1405 268
tri 1405 252 1421 268 sw
rect 1345 219 1421 252
rect 1345 185 1366 219
rect 1400 185 1421 219
rect 1345 183 1421 185
tri 1345 167 1361 183 ne
rect 1361 167 1405 183
tri 1405 167 1421 183 nw
rect 1451 263 1507 298
rect 1451 229 1463 263
rect 1497 229 1507 263
rect 1451 195 1507 229
rect 1259 137 1315 161
tri 1315 137 1345 167 sw
tri 1421 137 1451 167 se
rect 1451 161 1463 195
rect 1497 161 1507 195
rect 1451 137 1507 161
rect 1259 125 1507 137
rect 1259 91 1269 125
rect 1303 91 1366 125
rect 1400 91 1463 125
rect 1497 91 1507 125
rect 1259 75 1507 91
rect 1719 335 1775 351
rect 1719 301 1729 335
rect 1763 301 1775 335
rect 1719 263 1775 301
rect 1805 335 2075 351
rect 1805 306 1826 335
tri 1805 290 1821 306 ne
rect 1821 301 1826 306
rect 1860 301 1923 335
rect 1957 301 2020 335
rect 2054 301 2075 335
rect 1821 290 2075 301
rect 2105 335 2161 351
rect 2105 301 2117 335
rect 2151 301 2161 335
rect 1719 229 1729 263
rect 1763 229 1775 263
tri 1881 260 1911 290 ne
rect 1911 263 1970 290
rect 1719 195 1775 229
rect 1719 161 1729 195
rect 1763 161 1775 195
rect 1719 129 1775 161
tri 1805 244 1821 260 se
rect 1821 244 1865 260
tri 1865 244 1881 260 sw
rect 1805 210 1881 244
rect 1805 176 1826 210
rect 1860 176 1881 210
rect 1805 175 1881 176
tri 1805 159 1821 175 ne
rect 1821 159 1865 175
tri 1865 159 1881 175 nw
rect 1911 229 1923 263
rect 1957 229 1970 263
tri 1970 260 2000 290 nw
rect 1911 195 1970 229
rect 1911 161 1923 195
rect 1957 161 1970 195
tri 2000 244 2016 260 se
rect 2016 244 2059 260
tri 2059 244 2075 260 sw
rect 2000 216 2075 244
rect 2000 182 2021 216
rect 2055 182 2075 216
tri 2000 166 2016 182 ne
rect 2016 166 2059 182
tri 2059 166 2075 182 nw
tri 1775 129 1805 159 sw
tri 1881 129 1911 159 se
rect 1911 136 1970 161
tri 1970 136 2000 166 sw
tri 2075 136 2105 166 se
rect 2105 136 2161 301
rect 1911 129 2161 136
rect 1719 125 2161 129
rect 1719 91 1729 125
rect 1763 91 1923 125
rect 1957 91 2020 125
rect 2054 91 2117 125
rect 2151 91 2161 125
rect 1719 75 2161 91
rect 2221 335 2277 351
rect 2221 301 2231 335
rect 2265 301 2277 335
rect 2221 263 2277 301
rect 2307 314 2469 351
tri 2307 298 2323 314 ne
rect 2323 298 2469 314
tri 2383 268 2413 298 ne
rect 2221 229 2231 263
rect 2265 229 2277 263
rect 2221 195 2277 229
rect 2221 161 2231 195
rect 2265 161 2277 195
tri 2307 252 2323 268 se
rect 2323 252 2367 268
tri 2367 252 2383 268 sw
rect 2307 219 2383 252
rect 2307 185 2328 219
rect 2362 185 2383 219
rect 2307 183 2383 185
tri 2307 167 2323 183 ne
rect 2323 167 2367 183
tri 2367 167 2383 183 nw
rect 2413 263 2469 298
rect 2413 229 2425 263
rect 2459 229 2469 263
rect 2413 195 2469 229
rect 2221 137 2277 161
tri 2277 137 2307 167 sw
tri 2383 137 2413 167 se
rect 2413 161 2425 195
rect 2459 161 2469 195
rect 2413 137 2469 161
rect 2221 125 2469 137
rect 2221 91 2231 125
rect 2265 91 2328 125
rect 2362 91 2425 125
rect 2459 91 2469 125
rect 2221 75 2469 91
rect 2702 333 2758 349
rect 2702 299 2712 333
rect 2746 299 2758 333
rect 2702 261 2758 299
rect 2788 333 2952 349
rect 2788 304 2809 333
tri 2788 288 2804 304 ne
rect 2804 299 2809 304
rect 2843 299 2906 333
rect 2940 299 2952 333
rect 2804 288 2952 299
rect 2982 312 3144 349
tri 2982 296 2998 312 ne
rect 2998 296 3144 312
rect 2702 227 2712 261
rect 2746 227 2758 261
tri 2864 258 2894 288 ne
rect 2894 261 2952 288
tri 3058 266 3088 296 ne
rect 2702 193 2758 227
rect 2702 159 2712 193
rect 2746 159 2758 193
rect 2702 127 2758 159
tri 2788 242 2804 258 se
rect 2804 242 2848 258
tri 2848 242 2864 258 sw
rect 2788 208 2864 242
rect 2788 174 2809 208
rect 2843 174 2864 208
rect 2788 173 2864 174
tri 2788 157 2804 173 ne
rect 2804 157 2848 173
tri 2848 157 2864 173 nw
rect 2894 227 2906 261
rect 2940 227 2952 261
rect 2894 193 2952 227
rect 2894 159 2906 193
rect 2940 159 2952 193
tri 2982 250 2998 266 se
rect 2998 250 3042 266
tri 3042 250 3058 266 sw
rect 2982 217 3058 250
rect 2982 183 3003 217
rect 3037 183 3058 217
rect 2982 181 3058 183
tri 2982 165 2998 181 ne
rect 2998 165 3042 181
tri 3042 165 3058 181 nw
rect 3088 261 3144 296
rect 3088 227 3100 261
rect 3134 227 3144 261
rect 3088 193 3144 227
tri 2758 127 2788 157 sw
tri 2864 127 2894 157 se
rect 2894 135 2952 159
tri 2952 135 2982 165 sw
tri 3058 135 3088 165 se
rect 3088 159 3100 193
rect 3134 159 3144 193
rect 3088 135 3144 159
rect 2894 127 3144 135
rect 2702 123 3144 127
rect 2702 89 2712 123
rect 2746 89 2906 123
rect 2940 89 3003 123
rect 3037 89 3100 123
rect 3134 89 3144 123
rect 2702 73 3144 89
rect 3368 333 3424 349
rect 3368 299 3378 333
rect 3412 299 3424 333
rect 3368 261 3424 299
rect 3454 333 3618 349
rect 3454 304 3475 333
tri 3454 288 3470 304 ne
rect 3470 299 3475 304
rect 3509 299 3572 333
rect 3606 299 3618 333
rect 3470 288 3618 299
rect 3648 312 3810 349
tri 3648 296 3664 312 ne
rect 3664 296 3810 312
rect 3368 227 3378 261
rect 3412 227 3424 261
tri 3530 258 3560 288 ne
rect 3560 261 3618 288
tri 3724 266 3754 296 ne
rect 3368 193 3424 227
rect 3368 159 3378 193
rect 3412 159 3424 193
rect 3368 127 3424 159
tri 3454 242 3470 258 se
rect 3470 242 3514 258
tri 3514 242 3530 258 sw
rect 3454 208 3530 242
rect 3454 174 3475 208
rect 3509 174 3530 208
rect 3454 173 3530 174
tri 3454 157 3470 173 ne
rect 3470 157 3514 173
tri 3514 157 3530 173 nw
rect 3560 227 3572 261
rect 3606 227 3618 261
rect 3560 193 3618 227
rect 3560 159 3572 193
rect 3606 159 3618 193
tri 3648 250 3664 266 se
rect 3664 250 3708 266
tri 3708 250 3724 266 sw
rect 3648 217 3724 250
rect 3648 183 3669 217
rect 3703 183 3724 217
rect 3648 181 3724 183
tri 3648 165 3664 181 ne
rect 3664 165 3708 181
tri 3708 165 3724 181 nw
rect 3754 261 3810 296
rect 3754 227 3766 261
rect 3800 227 3810 261
rect 3754 193 3810 227
tri 3424 127 3454 157 sw
tri 3530 127 3560 157 se
rect 3560 135 3618 159
tri 3618 135 3648 165 sw
tri 3724 135 3754 165 se
rect 3754 159 3766 193
rect 3800 159 3810 193
rect 3754 135 3810 159
rect 3560 127 3810 135
rect 3368 123 3810 127
rect 3368 89 3378 123
rect 3412 89 3572 123
rect 3606 89 3669 123
rect 3703 89 3766 123
rect 3800 89 3810 123
rect 3368 73 3810 89
rect 4013 335 4069 351
rect 4013 301 4023 335
rect 4057 301 4069 335
rect 4013 263 4069 301
rect 4099 335 4369 351
rect 4099 306 4120 335
tri 4099 290 4115 306 ne
rect 4115 301 4120 306
rect 4154 301 4217 335
rect 4251 301 4314 335
rect 4348 301 4369 335
rect 4115 290 4369 301
rect 4399 335 4455 351
rect 4399 301 4411 335
rect 4445 301 4455 335
rect 4013 229 4023 263
rect 4057 229 4069 263
tri 4175 260 4205 290 ne
rect 4205 263 4264 290
rect 4013 195 4069 229
rect 4013 161 4023 195
rect 4057 161 4069 195
rect 4013 129 4069 161
tri 4099 244 4115 260 se
rect 4115 244 4159 260
tri 4159 244 4175 260 sw
rect 4099 210 4175 244
rect 4099 176 4120 210
rect 4154 176 4175 210
rect 4099 175 4175 176
tri 4099 159 4115 175 ne
rect 4115 159 4159 175
tri 4159 159 4175 175 nw
rect 4205 229 4217 263
rect 4251 229 4264 263
tri 4264 260 4294 290 nw
rect 4205 195 4264 229
rect 4205 161 4217 195
rect 4251 161 4264 195
tri 4294 244 4310 260 se
rect 4310 244 4353 260
tri 4353 244 4369 260 sw
rect 4294 216 4369 244
rect 4294 182 4315 216
rect 4349 182 4369 216
tri 4294 166 4310 182 ne
rect 4310 166 4353 182
tri 4353 166 4369 182 nw
tri 4069 129 4099 159 sw
tri 4175 129 4205 159 se
rect 4205 136 4264 161
tri 4264 136 4294 166 sw
tri 4369 136 4399 166 se
rect 4399 136 4455 301
rect 4205 129 4455 136
rect 4013 125 4455 129
rect 4013 91 4023 125
rect 4057 91 4217 125
rect 4251 91 4314 125
rect 4348 91 4411 125
rect 4445 91 4455 125
rect 4013 75 4455 91
rect 4515 335 4571 351
rect 4515 301 4525 335
rect 4559 301 4571 335
rect 4515 263 4571 301
rect 4601 314 4763 351
tri 4601 298 4617 314 ne
rect 4617 298 4763 314
tri 4677 268 4707 298 ne
rect 4515 229 4525 263
rect 4559 229 4571 263
rect 4515 195 4571 229
rect 4515 161 4525 195
rect 4559 161 4571 195
tri 4601 252 4617 268 se
rect 4617 252 4661 268
tri 4661 252 4677 268 sw
rect 4601 219 4677 252
rect 4601 185 4622 219
rect 4656 185 4677 219
rect 4601 183 4677 185
tri 4601 167 4617 183 ne
rect 4617 167 4661 183
tri 4661 167 4677 183 nw
rect 4707 263 4763 298
rect 4707 229 4719 263
rect 4753 229 4763 263
rect 4707 195 4763 229
rect 4515 137 4571 161
tri 4571 137 4601 167 sw
tri 4677 137 4707 167 se
rect 4707 161 4719 195
rect 4753 161 4763 195
rect 4707 137 4763 161
rect 4515 125 4763 137
rect 4515 91 4525 125
rect 4559 91 4622 125
rect 4656 91 4719 125
rect 4753 91 4763 125
rect 4515 75 4763 91
<< pdiff >>
rect 131 1366 187 1404
rect 131 1332 141 1366
rect 175 1332 187 1366
rect 131 1298 187 1332
rect 131 1264 141 1298
rect 175 1264 187 1298
rect 131 1230 187 1264
rect 131 1196 141 1230
rect 175 1196 187 1230
rect 131 1162 187 1196
rect 131 1128 141 1162
rect 175 1128 187 1162
rect 131 1093 187 1128
rect 131 1059 141 1093
rect 175 1059 187 1093
rect 131 1004 187 1059
rect 217 1366 275 1404
rect 217 1332 229 1366
rect 263 1332 275 1366
rect 217 1298 275 1332
rect 217 1264 229 1298
rect 263 1264 275 1298
rect 217 1230 275 1264
rect 217 1196 229 1230
rect 263 1196 275 1230
rect 217 1162 275 1196
rect 217 1128 229 1162
rect 263 1128 275 1162
rect 217 1093 275 1128
rect 217 1059 229 1093
rect 263 1059 275 1093
rect 217 1004 275 1059
rect 305 1366 363 1404
rect 305 1332 317 1366
rect 351 1332 363 1366
rect 305 1298 363 1332
rect 305 1264 317 1298
rect 351 1264 363 1298
rect 305 1230 363 1264
rect 305 1196 317 1230
rect 351 1196 363 1230
rect 305 1162 363 1196
rect 305 1128 317 1162
rect 351 1128 363 1162
rect 305 1004 363 1128
rect 393 1366 451 1404
rect 393 1332 405 1366
rect 439 1332 451 1366
rect 393 1298 451 1332
rect 393 1264 405 1298
rect 439 1264 451 1298
rect 393 1230 451 1264
rect 393 1196 405 1230
rect 439 1196 451 1230
rect 393 1162 451 1196
rect 393 1128 405 1162
rect 439 1128 451 1162
rect 393 1093 451 1128
rect 393 1059 405 1093
rect 439 1059 451 1093
rect 393 1004 451 1059
rect 481 1366 535 1404
rect 481 1332 493 1366
rect 527 1332 535 1366
rect 481 1298 535 1332
rect 481 1264 493 1298
rect 527 1264 535 1298
rect 481 1230 535 1264
rect 481 1196 493 1230
rect 527 1196 535 1230
rect 481 1162 535 1196
rect 481 1128 493 1162
rect 527 1128 535 1162
rect 481 1004 535 1128
rect 857 1366 913 1404
rect 857 1332 867 1366
rect 901 1332 913 1366
rect 857 1298 913 1332
rect 857 1264 867 1298
rect 901 1264 913 1298
rect 857 1230 913 1264
rect 857 1196 867 1230
rect 901 1196 913 1230
rect 857 1162 913 1196
rect 857 1128 867 1162
rect 901 1128 913 1162
rect 857 1093 913 1128
rect 857 1059 867 1093
rect 901 1059 913 1093
rect 857 1004 913 1059
rect 943 1366 1001 1404
rect 943 1332 955 1366
rect 989 1332 1001 1366
rect 943 1298 1001 1332
rect 943 1264 955 1298
rect 989 1264 1001 1298
rect 943 1230 1001 1264
rect 943 1196 955 1230
rect 989 1196 1001 1230
rect 943 1162 1001 1196
rect 943 1128 955 1162
rect 989 1128 1001 1162
rect 943 1093 1001 1128
rect 943 1059 955 1093
rect 989 1059 1001 1093
rect 943 1004 1001 1059
rect 1031 1366 1089 1404
rect 1031 1332 1043 1366
rect 1077 1332 1089 1366
rect 1031 1298 1089 1332
rect 1031 1264 1043 1298
rect 1077 1264 1089 1298
rect 1031 1230 1089 1264
rect 1031 1196 1043 1230
rect 1077 1196 1089 1230
rect 1031 1162 1089 1196
rect 1031 1128 1043 1162
rect 1077 1128 1089 1162
rect 1031 1004 1089 1128
rect 1119 1366 1177 1404
rect 1119 1332 1131 1366
rect 1165 1332 1177 1366
rect 1119 1298 1177 1332
rect 1119 1264 1131 1298
rect 1165 1264 1177 1298
rect 1119 1230 1177 1264
rect 1119 1196 1131 1230
rect 1165 1196 1177 1230
rect 1119 1162 1177 1196
rect 1119 1128 1131 1162
rect 1165 1128 1177 1162
rect 1119 1093 1177 1128
rect 1119 1059 1131 1093
rect 1165 1059 1177 1093
rect 1119 1004 1177 1059
rect 1207 1366 1265 1404
rect 1207 1332 1219 1366
rect 1253 1332 1265 1366
rect 1207 1298 1265 1332
rect 1207 1264 1219 1298
rect 1253 1264 1265 1298
rect 1207 1230 1265 1264
rect 1207 1196 1219 1230
rect 1253 1196 1265 1230
rect 1207 1162 1265 1196
rect 1207 1128 1219 1162
rect 1253 1128 1265 1162
rect 1207 1004 1265 1128
rect 1295 1366 1353 1404
rect 1295 1332 1307 1366
rect 1341 1332 1353 1366
rect 1295 1298 1353 1332
rect 1295 1264 1307 1298
rect 1341 1264 1353 1298
rect 1295 1230 1353 1264
rect 1295 1196 1307 1230
rect 1341 1196 1353 1230
rect 1295 1162 1353 1196
rect 1295 1128 1307 1162
rect 1341 1128 1353 1162
rect 1295 1093 1353 1128
rect 1295 1059 1307 1093
rect 1341 1059 1353 1093
rect 1295 1004 1353 1059
rect 1383 1366 1437 1404
rect 1383 1332 1395 1366
rect 1429 1332 1437 1366
rect 1383 1298 1437 1332
rect 1383 1264 1395 1298
rect 1429 1264 1437 1298
rect 1383 1230 1437 1264
rect 1383 1196 1395 1230
rect 1429 1196 1437 1230
rect 1383 1162 1437 1196
rect 1383 1128 1395 1162
rect 1429 1128 1437 1162
rect 1383 1004 1437 1128
rect 1819 1366 1875 1404
rect 1819 1332 1829 1366
rect 1863 1332 1875 1366
rect 1819 1298 1875 1332
rect 1819 1264 1829 1298
rect 1863 1264 1875 1298
rect 1819 1230 1875 1264
rect 1819 1196 1829 1230
rect 1863 1196 1875 1230
rect 1819 1162 1875 1196
rect 1819 1128 1829 1162
rect 1863 1128 1875 1162
rect 1819 1093 1875 1128
rect 1819 1059 1829 1093
rect 1863 1059 1875 1093
rect 1819 1004 1875 1059
rect 1905 1366 1963 1404
rect 1905 1332 1917 1366
rect 1951 1332 1963 1366
rect 1905 1298 1963 1332
rect 1905 1264 1917 1298
rect 1951 1264 1963 1298
rect 1905 1230 1963 1264
rect 1905 1196 1917 1230
rect 1951 1196 1963 1230
rect 1905 1162 1963 1196
rect 1905 1128 1917 1162
rect 1951 1128 1963 1162
rect 1905 1093 1963 1128
rect 1905 1059 1917 1093
rect 1951 1059 1963 1093
rect 1905 1004 1963 1059
rect 1993 1366 2051 1404
rect 1993 1332 2005 1366
rect 2039 1332 2051 1366
rect 1993 1298 2051 1332
rect 1993 1264 2005 1298
rect 2039 1264 2051 1298
rect 1993 1230 2051 1264
rect 1993 1196 2005 1230
rect 2039 1196 2051 1230
rect 1993 1162 2051 1196
rect 1993 1128 2005 1162
rect 2039 1128 2051 1162
rect 1993 1004 2051 1128
rect 2081 1366 2139 1404
rect 2081 1332 2093 1366
rect 2127 1332 2139 1366
rect 2081 1298 2139 1332
rect 2081 1264 2093 1298
rect 2127 1264 2139 1298
rect 2081 1230 2139 1264
rect 2081 1196 2093 1230
rect 2127 1196 2139 1230
rect 2081 1162 2139 1196
rect 2081 1128 2093 1162
rect 2127 1128 2139 1162
rect 2081 1093 2139 1128
rect 2081 1059 2093 1093
rect 2127 1059 2139 1093
rect 2081 1004 2139 1059
rect 2169 1366 2227 1404
rect 2169 1332 2181 1366
rect 2215 1332 2227 1366
rect 2169 1298 2227 1332
rect 2169 1264 2181 1298
rect 2215 1264 2227 1298
rect 2169 1230 2227 1264
rect 2169 1196 2181 1230
rect 2215 1196 2227 1230
rect 2169 1162 2227 1196
rect 2169 1128 2181 1162
rect 2215 1128 2227 1162
rect 2169 1004 2227 1128
rect 2257 1366 2315 1404
rect 2257 1332 2269 1366
rect 2303 1332 2315 1366
rect 2257 1298 2315 1332
rect 2257 1264 2269 1298
rect 2303 1264 2315 1298
rect 2257 1230 2315 1264
rect 2257 1196 2269 1230
rect 2303 1196 2315 1230
rect 2257 1162 2315 1196
rect 2257 1128 2269 1162
rect 2303 1128 2315 1162
rect 2257 1093 2315 1128
rect 2257 1059 2269 1093
rect 2303 1059 2315 1093
rect 2257 1004 2315 1059
rect 2345 1366 2399 1404
rect 2345 1332 2357 1366
rect 2391 1332 2399 1366
rect 2345 1298 2399 1332
rect 2345 1264 2357 1298
rect 2391 1264 2399 1298
rect 2345 1230 2399 1264
rect 2345 1196 2357 1230
rect 2391 1196 2399 1230
rect 2345 1162 2399 1196
rect 2345 1128 2357 1162
rect 2391 1128 2399 1162
rect 2345 1004 2399 1128
rect 2721 1366 2777 1404
rect 2721 1332 2731 1366
rect 2765 1332 2777 1366
rect 2721 1298 2777 1332
rect 2721 1264 2731 1298
rect 2765 1264 2777 1298
rect 2721 1230 2777 1264
rect 2721 1196 2731 1230
rect 2765 1196 2777 1230
rect 2721 1162 2777 1196
rect 2721 1128 2731 1162
rect 2765 1128 2777 1162
rect 2721 1093 2777 1128
rect 2721 1059 2731 1093
rect 2765 1059 2777 1093
rect 2721 1004 2777 1059
rect 2807 1366 2865 1404
rect 2807 1332 2819 1366
rect 2853 1332 2865 1366
rect 2807 1298 2865 1332
rect 2807 1264 2819 1298
rect 2853 1264 2865 1298
rect 2807 1230 2865 1264
rect 2807 1196 2819 1230
rect 2853 1196 2865 1230
rect 2807 1162 2865 1196
rect 2807 1128 2819 1162
rect 2853 1128 2865 1162
rect 2807 1093 2865 1128
rect 2807 1059 2819 1093
rect 2853 1059 2865 1093
rect 2807 1004 2865 1059
rect 2895 1366 2953 1404
rect 2895 1332 2907 1366
rect 2941 1332 2953 1366
rect 2895 1298 2953 1332
rect 2895 1264 2907 1298
rect 2941 1264 2953 1298
rect 2895 1230 2953 1264
rect 2895 1196 2907 1230
rect 2941 1196 2953 1230
rect 2895 1162 2953 1196
rect 2895 1128 2907 1162
rect 2941 1128 2953 1162
rect 2895 1004 2953 1128
rect 2983 1366 3041 1404
rect 2983 1332 2995 1366
rect 3029 1332 3041 1366
rect 2983 1298 3041 1332
rect 2983 1264 2995 1298
rect 3029 1264 3041 1298
rect 2983 1230 3041 1264
rect 2983 1196 2995 1230
rect 3029 1196 3041 1230
rect 2983 1162 3041 1196
rect 2983 1128 2995 1162
rect 3029 1128 3041 1162
rect 2983 1093 3041 1128
rect 2983 1059 2995 1093
rect 3029 1059 3041 1093
rect 2983 1004 3041 1059
rect 3071 1366 3125 1404
rect 3071 1332 3083 1366
rect 3117 1332 3125 1366
rect 3071 1298 3125 1332
rect 3071 1264 3083 1298
rect 3117 1264 3125 1298
rect 3071 1230 3125 1264
rect 3071 1196 3083 1230
rect 3117 1196 3125 1230
rect 3071 1162 3125 1196
rect 3071 1128 3083 1162
rect 3117 1128 3125 1162
rect 3071 1004 3125 1128
rect 3387 1366 3443 1404
rect 3387 1332 3397 1366
rect 3431 1332 3443 1366
rect 3387 1298 3443 1332
rect 3387 1264 3397 1298
rect 3431 1264 3443 1298
rect 3387 1230 3443 1264
rect 3387 1196 3397 1230
rect 3431 1196 3443 1230
rect 3387 1162 3443 1196
rect 3387 1128 3397 1162
rect 3431 1128 3443 1162
rect 3387 1093 3443 1128
rect 3387 1059 3397 1093
rect 3431 1059 3443 1093
rect 3387 1004 3443 1059
rect 3473 1366 3531 1404
rect 3473 1332 3485 1366
rect 3519 1332 3531 1366
rect 3473 1298 3531 1332
rect 3473 1264 3485 1298
rect 3519 1264 3531 1298
rect 3473 1230 3531 1264
rect 3473 1196 3485 1230
rect 3519 1196 3531 1230
rect 3473 1162 3531 1196
rect 3473 1128 3485 1162
rect 3519 1128 3531 1162
rect 3473 1093 3531 1128
rect 3473 1059 3485 1093
rect 3519 1059 3531 1093
rect 3473 1004 3531 1059
rect 3561 1366 3619 1404
rect 3561 1332 3573 1366
rect 3607 1332 3619 1366
rect 3561 1298 3619 1332
rect 3561 1264 3573 1298
rect 3607 1264 3619 1298
rect 3561 1230 3619 1264
rect 3561 1196 3573 1230
rect 3607 1196 3619 1230
rect 3561 1162 3619 1196
rect 3561 1128 3573 1162
rect 3607 1128 3619 1162
rect 3561 1004 3619 1128
rect 3649 1366 3707 1404
rect 3649 1332 3661 1366
rect 3695 1332 3707 1366
rect 3649 1298 3707 1332
rect 3649 1264 3661 1298
rect 3695 1264 3707 1298
rect 3649 1230 3707 1264
rect 3649 1196 3661 1230
rect 3695 1196 3707 1230
rect 3649 1162 3707 1196
rect 3649 1128 3661 1162
rect 3695 1128 3707 1162
rect 3649 1093 3707 1128
rect 3649 1059 3661 1093
rect 3695 1059 3707 1093
rect 3649 1004 3707 1059
rect 3737 1366 3791 1404
rect 3737 1332 3749 1366
rect 3783 1332 3791 1366
rect 3737 1298 3791 1332
rect 3737 1264 3749 1298
rect 3783 1264 3791 1298
rect 3737 1230 3791 1264
rect 3737 1196 3749 1230
rect 3783 1196 3791 1230
rect 3737 1162 3791 1196
rect 3737 1128 3749 1162
rect 3783 1128 3791 1162
rect 3737 1004 3791 1128
rect 4113 1366 4169 1404
rect 4113 1332 4123 1366
rect 4157 1332 4169 1366
rect 4113 1298 4169 1332
rect 4113 1264 4123 1298
rect 4157 1264 4169 1298
rect 4113 1230 4169 1264
rect 4113 1196 4123 1230
rect 4157 1196 4169 1230
rect 4113 1162 4169 1196
rect 4113 1128 4123 1162
rect 4157 1128 4169 1162
rect 4113 1093 4169 1128
rect 4113 1059 4123 1093
rect 4157 1059 4169 1093
rect 4113 1004 4169 1059
rect 4199 1366 4257 1404
rect 4199 1332 4211 1366
rect 4245 1332 4257 1366
rect 4199 1298 4257 1332
rect 4199 1264 4211 1298
rect 4245 1264 4257 1298
rect 4199 1230 4257 1264
rect 4199 1196 4211 1230
rect 4245 1196 4257 1230
rect 4199 1162 4257 1196
rect 4199 1128 4211 1162
rect 4245 1128 4257 1162
rect 4199 1093 4257 1128
rect 4199 1059 4211 1093
rect 4245 1059 4257 1093
rect 4199 1004 4257 1059
rect 4287 1366 4345 1404
rect 4287 1332 4299 1366
rect 4333 1332 4345 1366
rect 4287 1298 4345 1332
rect 4287 1264 4299 1298
rect 4333 1264 4345 1298
rect 4287 1230 4345 1264
rect 4287 1196 4299 1230
rect 4333 1196 4345 1230
rect 4287 1162 4345 1196
rect 4287 1128 4299 1162
rect 4333 1128 4345 1162
rect 4287 1004 4345 1128
rect 4375 1366 4433 1404
rect 4375 1332 4387 1366
rect 4421 1332 4433 1366
rect 4375 1298 4433 1332
rect 4375 1264 4387 1298
rect 4421 1264 4433 1298
rect 4375 1230 4433 1264
rect 4375 1196 4387 1230
rect 4421 1196 4433 1230
rect 4375 1162 4433 1196
rect 4375 1128 4387 1162
rect 4421 1128 4433 1162
rect 4375 1093 4433 1128
rect 4375 1059 4387 1093
rect 4421 1059 4433 1093
rect 4375 1004 4433 1059
rect 4463 1366 4521 1404
rect 4463 1332 4475 1366
rect 4509 1332 4521 1366
rect 4463 1298 4521 1332
rect 4463 1264 4475 1298
rect 4509 1264 4521 1298
rect 4463 1230 4521 1264
rect 4463 1196 4475 1230
rect 4509 1196 4521 1230
rect 4463 1162 4521 1196
rect 4463 1128 4475 1162
rect 4509 1128 4521 1162
rect 4463 1004 4521 1128
rect 4551 1366 4609 1404
rect 4551 1332 4563 1366
rect 4597 1332 4609 1366
rect 4551 1298 4609 1332
rect 4551 1264 4563 1298
rect 4597 1264 4609 1298
rect 4551 1230 4609 1264
rect 4551 1196 4563 1230
rect 4597 1196 4609 1230
rect 4551 1162 4609 1196
rect 4551 1128 4563 1162
rect 4597 1128 4609 1162
rect 4551 1093 4609 1128
rect 4551 1059 4563 1093
rect 4597 1059 4609 1093
rect 4551 1004 4609 1059
rect 4639 1366 4693 1404
rect 4639 1332 4651 1366
rect 4685 1332 4693 1366
rect 4639 1298 4693 1332
rect 4639 1264 4651 1298
rect 4685 1264 4693 1298
rect 4639 1230 4693 1264
rect 4639 1196 4651 1230
rect 4685 1196 4693 1230
rect 4639 1162 4693 1196
rect 4639 1128 4651 1162
rect 4685 1128 4693 1162
rect 4639 1004 4693 1128
<< ndiffc >>
rect 122 299 156 333
rect 219 299 253 333
rect 316 299 350 333
rect 122 227 156 261
rect 122 159 156 193
rect 219 174 253 208
rect 316 227 350 261
rect 316 159 350 193
rect 413 183 447 217
rect 510 227 544 261
rect 510 159 544 193
rect 122 89 156 123
rect 316 89 350 123
rect 413 89 447 123
rect 510 89 544 123
rect 767 301 801 335
rect 864 301 898 335
rect 961 301 995 335
rect 1058 301 1092 335
rect 1155 301 1189 335
rect 767 229 801 263
rect 767 161 801 195
rect 864 176 898 210
rect 961 229 995 263
rect 961 161 995 195
rect 1059 182 1093 216
rect 767 91 801 125
rect 961 91 995 125
rect 1058 91 1092 125
rect 1155 91 1189 125
rect 1269 301 1303 335
rect 1269 229 1303 263
rect 1269 161 1303 195
rect 1366 185 1400 219
rect 1463 229 1497 263
rect 1463 161 1497 195
rect 1269 91 1303 125
rect 1366 91 1400 125
rect 1463 91 1497 125
rect 1729 301 1763 335
rect 1826 301 1860 335
rect 1923 301 1957 335
rect 2020 301 2054 335
rect 2117 301 2151 335
rect 1729 229 1763 263
rect 1729 161 1763 195
rect 1826 176 1860 210
rect 1923 229 1957 263
rect 1923 161 1957 195
rect 2021 182 2055 216
rect 1729 91 1763 125
rect 1923 91 1957 125
rect 2020 91 2054 125
rect 2117 91 2151 125
rect 2231 301 2265 335
rect 2231 229 2265 263
rect 2231 161 2265 195
rect 2328 185 2362 219
rect 2425 229 2459 263
rect 2425 161 2459 195
rect 2231 91 2265 125
rect 2328 91 2362 125
rect 2425 91 2459 125
rect 2712 299 2746 333
rect 2809 299 2843 333
rect 2906 299 2940 333
rect 2712 227 2746 261
rect 2712 159 2746 193
rect 2809 174 2843 208
rect 2906 227 2940 261
rect 2906 159 2940 193
rect 3003 183 3037 217
rect 3100 227 3134 261
rect 3100 159 3134 193
rect 2712 89 2746 123
rect 2906 89 2940 123
rect 3003 89 3037 123
rect 3100 89 3134 123
rect 3378 299 3412 333
rect 3475 299 3509 333
rect 3572 299 3606 333
rect 3378 227 3412 261
rect 3378 159 3412 193
rect 3475 174 3509 208
rect 3572 227 3606 261
rect 3572 159 3606 193
rect 3669 183 3703 217
rect 3766 227 3800 261
rect 3766 159 3800 193
rect 3378 89 3412 123
rect 3572 89 3606 123
rect 3669 89 3703 123
rect 3766 89 3800 123
rect 4023 301 4057 335
rect 4120 301 4154 335
rect 4217 301 4251 335
rect 4314 301 4348 335
rect 4411 301 4445 335
rect 4023 229 4057 263
rect 4023 161 4057 195
rect 4120 176 4154 210
rect 4217 229 4251 263
rect 4217 161 4251 195
rect 4315 182 4349 216
rect 4023 91 4057 125
rect 4217 91 4251 125
rect 4314 91 4348 125
rect 4411 91 4445 125
rect 4525 301 4559 335
rect 4525 229 4559 263
rect 4525 161 4559 195
rect 4622 185 4656 219
rect 4719 229 4753 263
rect 4719 161 4753 195
rect 4525 91 4559 125
rect 4622 91 4656 125
rect 4719 91 4753 125
<< pdiffc >>
rect 141 1332 175 1366
rect 141 1264 175 1298
rect 141 1196 175 1230
rect 141 1128 175 1162
rect 141 1059 175 1093
rect 229 1332 263 1366
rect 229 1264 263 1298
rect 229 1196 263 1230
rect 229 1128 263 1162
rect 229 1059 263 1093
rect 317 1332 351 1366
rect 317 1264 351 1298
rect 317 1196 351 1230
rect 317 1128 351 1162
rect 405 1332 439 1366
rect 405 1264 439 1298
rect 405 1196 439 1230
rect 405 1128 439 1162
rect 405 1059 439 1093
rect 493 1332 527 1366
rect 493 1264 527 1298
rect 493 1196 527 1230
rect 493 1128 527 1162
rect 867 1332 901 1366
rect 867 1264 901 1298
rect 867 1196 901 1230
rect 867 1128 901 1162
rect 867 1059 901 1093
rect 955 1332 989 1366
rect 955 1264 989 1298
rect 955 1196 989 1230
rect 955 1128 989 1162
rect 955 1059 989 1093
rect 1043 1332 1077 1366
rect 1043 1264 1077 1298
rect 1043 1196 1077 1230
rect 1043 1128 1077 1162
rect 1131 1332 1165 1366
rect 1131 1264 1165 1298
rect 1131 1196 1165 1230
rect 1131 1128 1165 1162
rect 1131 1059 1165 1093
rect 1219 1332 1253 1366
rect 1219 1264 1253 1298
rect 1219 1196 1253 1230
rect 1219 1128 1253 1162
rect 1307 1332 1341 1366
rect 1307 1264 1341 1298
rect 1307 1196 1341 1230
rect 1307 1128 1341 1162
rect 1307 1059 1341 1093
rect 1395 1332 1429 1366
rect 1395 1264 1429 1298
rect 1395 1196 1429 1230
rect 1395 1128 1429 1162
rect 1829 1332 1863 1366
rect 1829 1264 1863 1298
rect 1829 1196 1863 1230
rect 1829 1128 1863 1162
rect 1829 1059 1863 1093
rect 1917 1332 1951 1366
rect 1917 1264 1951 1298
rect 1917 1196 1951 1230
rect 1917 1128 1951 1162
rect 1917 1059 1951 1093
rect 2005 1332 2039 1366
rect 2005 1264 2039 1298
rect 2005 1196 2039 1230
rect 2005 1128 2039 1162
rect 2093 1332 2127 1366
rect 2093 1264 2127 1298
rect 2093 1196 2127 1230
rect 2093 1128 2127 1162
rect 2093 1059 2127 1093
rect 2181 1332 2215 1366
rect 2181 1264 2215 1298
rect 2181 1196 2215 1230
rect 2181 1128 2215 1162
rect 2269 1332 2303 1366
rect 2269 1264 2303 1298
rect 2269 1196 2303 1230
rect 2269 1128 2303 1162
rect 2269 1059 2303 1093
rect 2357 1332 2391 1366
rect 2357 1264 2391 1298
rect 2357 1196 2391 1230
rect 2357 1128 2391 1162
rect 2731 1332 2765 1366
rect 2731 1264 2765 1298
rect 2731 1196 2765 1230
rect 2731 1128 2765 1162
rect 2731 1059 2765 1093
rect 2819 1332 2853 1366
rect 2819 1264 2853 1298
rect 2819 1196 2853 1230
rect 2819 1128 2853 1162
rect 2819 1059 2853 1093
rect 2907 1332 2941 1366
rect 2907 1264 2941 1298
rect 2907 1196 2941 1230
rect 2907 1128 2941 1162
rect 2995 1332 3029 1366
rect 2995 1264 3029 1298
rect 2995 1196 3029 1230
rect 2995 1128 3029 1162
rect 2995 1059 3029 1093
rect 3083 1332 3117 1366
rect 3083 1264 3117 1298
rect 3083 1196 3117 1230
rect 3083 1128 3117 1162
rect 3397 1332 3431 1366
rect 3397 1264 3431 1298
rect 3397 1196 3431 1230
rect 3397 1128 3431 1162
rect 3397 1059 3431 1093
rect 3485 1332 3519 1366
rect 3485 1264 3519 1298
rect 3485 1196 3519 1230
rect 3485 1128 3519 1162
rect 3485 1059 3519 1093
rect 3573 1332 3607 1366
rect 3573 1264 3607 1298
rect 3573 1196 3607 1230
rect 3573 1128 3607 1162
rect 3661 1332 3695 1366
rect 3661 1264 3695 1298
rect 3661 1196 3695 1230
rect 3661 1128 3695 1162
rect 3661 1059 3695 1093
rect 3749 1332 3783 1366
rect 3749 1264 3783 1298
rect 3749 1196 3783 1230
rect 3749 1128 3783 1162
rect 4123 1332 4157 1366
rect 4123 1264 4157 1298
rect 4123 1196 4157 1230
rect 4123 1128 4157 1162
rect 4123 1059 4157 1093
rect 4211 1332 4245 1366
rect 4211 1264 4245 1298
rect 4211 1196 4245 1230
rect 4211 1128 4245 1162
rect 4211 1059 4245 1093
rect 4299 1332 4333 1366
rect 4299 1264 4333 1298
rect 4299 1196 4333 1230
rect 4299 1128 4333 1162
rect 4387 1332 4421 1366
rect 4387 1264 4421 1298
rect 4387 1196 4421 1230
rect 4387 1128 4421 1162
rect 4387 1059 4421 1093
rect 4475 1332 4509 1366
rect 4475 1264 4509 1298
rect 4475 1196 4509 1230
rect 4475 1128 4509 1162
rect 4563 1332 4597 1366
rect 4563 1264 4597 1298
rect 4563 1196 4597 1230
rect 4563 1128 4597 1162
rect 4563 1059 4597 1093
rect 4651 1332 4685 1366
rect 4651 1264 4685 1298
rect 4651 1196 4685 1230
rect 4651 1128 4685 1162
<< psubdiff >>
rect -34 482 4918 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 632 461 700 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 632 427 649 461
rect 683 427 700 461
rect 1594 461 1662 482
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 632 313 700 353
rect 1594 427 1611 461
rect 1645 427 1662 461
rect 2556 461 2624 482
rect 1594 387 1662 427
rect 1594 353 1611 387
rect 1645 353 1662 387
rect 632 279 649 313
rect 683 279 700 313
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect -34 17 34 57
rect 632 57 649 91
rect 683 57 700 91
rect 1594 313 1662 353
rect 2556 427 2573 461
rect 2607 427 2624 461
rect 3222 461 3290 482
rect 2556 387 2624 427
rect 2556 353 2573 387
rect 2607 353 2624 387
rect 1594 279 1611 313
rect 1645 279 1662 313
rect 1594 239 1662 279
rect 1594 205 1611 239
rect 1645 205 1662 239
rect 1594 165 1662 205
rect 1594 131 1611 165
rect 1645 131 1662 165
rect 1594 91 1662 131
rect 632 17 700 57
rect 1594 57 1611 91
rect 1645 57 1662 91
rect 2556 313 2624 353
rect 3222 427 3239 461
rect 3273 427 3290 461
rect 3888 461 3956 482
rect 3222 387 3290 427
rect 3222 353 3239 387
rect 3273 353 3290 387
rect 2556 279 2573 313
rect 2607 279 2624 313
rect 2556 239 2624 279
rect 2556 205 2573 239
rect 2607 205 2624 239
rect 2556 165 2624 205
rect 2556 131 2573 165
rect 2607 131 2624 165
rect 2556 91 2624 131
rect 1594 17 1662 57
rect 2556 57 2573 91
rect 2607 57 2624 91
rect 3222 313 3290 353
rect 3888 427 3905 461
rect 3939 427 3956 461
rect 4850 461 4918 482
rect 3888 387 3956 427
rect 3888 353 3905 387
rect 3939 353 3956 387
rect 3222 279 3239 313
rect 3273 279 3290 313
rect 3222 239 3290 279
rect 3222 205 3239 239
rect 3273 205 3290 239
rect 3222 165 3290 205
rect 3222 131 3239 165
rect 3273 131 3290 165
rect 3222 91 3290 131
rect 2556 17 2624 57
rect 3222 57 3239 91
rect 3273 57 3290 91
rect 3888 313 3956 353
rect 4850 427 4867 461
rect 4901 427 4918 461
rect 4850 387 4918 427
rect 4850 353 4867 387
rect 4901 353 4918 387
rect 3888 279 3905 313
rect 3939 279 3956 313
rect 3888 239 3956 279
rect 3888 205 3905 239
rect 3939 205 3956 239
rect 3888 165 3956 205
rect 3888 131 3905 165
rect 3939 131 3956 165
rect 3888 91 3956 131
rect 3222 17 3290 57
rect 3888 57 3905 91
rect 3939 57 3956 91
rect 4850 313 4918 353
rect 4850 279 4867 313
rect 4901 279 4918 313
rect 4850 239 4918 279
rect 4850 205 4867 239
rect 4901 205 4918 239
rect 4850 165 4918 205
rect 4850 131 4867 165
rect 4901 131 4918 165
rect 4850 91 4918 131
rect 3888 17 3956 57
rect 4850 57 4867 91
rect 4901 57 4918 91
rect 4850 17 4918 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4918 17
rect -34 -34 4918 -17
<< nsubdiff >>
rect -34 1497 4918 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4918 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 632 1423 700 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 1594 1423 1662 1463
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 632 979 700 1019
rect 1594 1389 1611 1423
rect 1645 1389 1662 1423
rect 2556 1423 2624 1463
rect 1594 1349 1662 1389
rect 1594 1315 1611 1349
rect 1645 1315 1662 1349
rect 1594 1275 1662 1315
rect 1594 1241 1611 1275
rect 1645 1241 1662 1275
rect 1594 1201 1662 1241
rect 1594 1167 1611 1201
rect 1645 1167 1662 1201
rect 1594 1127 1662 1167
rect 1594 1093 1611 1127
rect 1645 1093 1662 1127
rect 1594 1053 1662 1093
rect 1594 1019 1611 1053
rect 1645 1019 1662 1053
rect 632 945 649 979
rect 683 945 700 979
rect -34 871 -17 905
rect 17 884 34 905
rect 632 905 700 945
rect 1594 979 1662 1019
rect 2556 1389 2573 1423
rect 2607 1389 2624 1423
rect 3222 1423 3290 1463
rect 2556 1349 2624 1389
rect 2556 1315 2573 1349
rect 2607 1315 2624 1349
rect 2556 1275 2624 1315
rect 2556 1241 2573 1275
rect 2607 1241 2624 1275
rect 2556 1201 2624 1241
rect 2556 1167 2573 1201
rect 2607 1167 2624 1201
rect 2556 1127 2624 1167
rect 2556 1093 2573 1127
rect 2607 1093 2624 1127
rect 2556 1053 2624 1093
rect 2556 1019 2573 1053
rect 2607 1019 2624 1053
rect 1594 945 1611 979
rect 1645 945 1662 979
rect 632 884 649 905
rect 17 871 649 884
rect 683 884 700 905
rect 1594 905 1662 945
rect 2556 979 2624 1019
rect 3222 1389 3239 1423
rect 3273 1389 3290 1423
rect 3888 1423 3956 1463
rect 3222 1349 3290 1389
rect 3222 1315 3239 1349
rect 3273 1315 3290 1349
rect 3222 1275 3290 1315
rect 3222 1241 3239 1275
rect 3273 1241 3290 1275
rect 3222 1201 3290 1241
rect 3222 1167 3239 1201
rect 3273 1167 3290 1201
rect 3222 1127 3290 1167
rect 3222 1093 3239 1127
rect 3273 1093 3290 1127
rect 3222 1053 3290 1093
rect 3222 1019 3239 1053
rect 3273 1019 3290 1053
rect 2556 945 2573 979
rect 2607 945 2624 979
rect 1594 884 1611 905
rect 683 871 1611 884
rect 1645 884 1662 905
rect 2556 905 2624 945
rect 3222 979 3290 1019
rect 3888 1389 3905 1423
rect 3939 1389 3956 1423
rect 4850 1423 4918 1463
rect 3888 1349 3956 1389
rect 3888 1315 3905 1349
rect 3939 1315 3956 1349
rect 3888 1275 3956 1315
rect 3888 1241 3905 1275
rect 3939 1241 3956 1275
rect 3888 1201 3956 1241
rect 3888 1167 3905 1201
rect 3939 1167 3956 1201
rect 3888 1127 3956 1167
rect 3888 1093 3905 1127
rect 3939 1093 3956 1127
rect 3888 1053 3956 1093
rect 3888 1019 3905 1053
rect 3939 1019 3956 1053
rect 3222 945 3239 979
rect 3273 945 3290 979
rect 2556 884 2573 905
rect 1645 871 2573 884
rect 2607 884 2624 905
rect 3222 905 3290 945
rect 3888 979 3956 1019
rect 4850 1389 4867 1423
rect 4901 1389 4918 1423
rect 4850 1349 4918 1389
rect 4850 1315 4867 1349
rect 4901 1315 4918 1349
rect 4850 1275 4918 1315
rect 4850 1241 4867 1275
rect 4901 1241 4918 1275
rect 4850 1201 4918 1241
rect 4850 1167 4867 1201
rect 4901 1167 4918 1201
rect 4850 1127 4918 1167
rect 4850 1093 4867 1127
rect 4901 1093 4918 1127
rect 4850 1053 4918 1093
rect 4850 1019 4867 1053
rect 4901 1019 4918 1053
rect 3888 945 3905 979
rect 3939 945 3956 979
rect 3222 884 3239 905
rect 2607 871 3239 884
rect 3273 884 3290 905
rect 3888 905 3956 945
rect 4850 979 4918 1019
rect 4850 945 4867 979
rect 4901 945 4918 979
rect 3888 884 3905 905
rect 3273 871 3905 884
rect 3939 884 3956 905
rect 4850 905 4918 945
rect 4850 884 4867 905
rect 3939 871 4867 884
rect 4901 871 4918 905
rect -34 822 4918 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 649 427 683 461
rect 649 353 683 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1611 427 1645 461
rect 1611 353 1645 387
rect 649 279 683 313
rect 649 205 683 239
rect 649 131 683 165
rect 649 57 683 91
rect 2573 427 2607 461
rect 2573 353 2607 387
rect 1611 279 1645 313
rect 1611 205 1645 239
rect 1611 131 1645 165
rect 1611 57 1645 91
rect 3239 427 3273 461
rect 3239 353 3273 387
rect 2573 279 2607 313
rect 2573 205 2607 239
rect 2573 131 2607 165
rect 2573 57 2607 91
rect 3905 427 3939 461
rect 3905 353 3939 387
rect 3239 279 3273 313
rect 3239 205 3273 239
rect 3239 131 3273 165
rect 3239 57 3273 91
rect 4867 427 4901 461
rect 4867 353 4901 387
rect 3905 279 3939 313
rect 3905 205 3939 239
rect 3905 131 3939 165
rect 3905 57 3939 91
rect 4867 279 4901 313
rect 4867 205 4901 239
rect 4867 131 4901 165
rect 4867 57 4901 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 649 1389 683 1423
rect 649 1315 683 1349
rect 649 1241 683 1275
rect 649 1167 683 1201
rect 649 1093 683 1127
rect 649 1019 683 1053
rect -17 945 17 979
rect 1611 1389 1645 1423
rect 1611 1315 1645 1349
rect 1611 1241 1645 1275
rect 1611 1167 1645 1201
rect 1611 1093 1645 1127
rect 1611 1019 1645 1053
rect 649 945 683 979
rect -17 871 17 905
rect 2573 1389 2607 1423
rect 2573 1315 2607 1349
rect 2573 1241 2607 1275
rect 2573 1167 2607 1201
rect 2573 1093 2607 1127
rect 2573 1019 2607 1053
rect 1611 945 1645 979
rect 649 871 683 905
rect 3239 1389 3273 1423
rect 3239 1315 3273 1349
rect 3239 1241 3273 1275
rect 3239 1167 3273 1201
rect 3239 1093 3273 1127
rect 3239 1019 3273 1053
rect 2573 945 2607 979
rect 1611 871 1645 905
rect 3905 1389 3939 1423
rect 3905 1315 3939 1349
rect 3905 1241 3939 1275
rect 3905 1167 3939 1201
rect 3905 1093 3939 1127
rect 3905 1019 3939 1053
rect 3239 945 3273 979
rect 2573 871 2607 905
rect 4867 1389 4901 1423
rect 4867 1315 4901 1349
rect 4867 1241 4901 1275
rect 4867 1167 4901 1201
rect 4867 1093 4901 1127
rect 4867 1019 4901 1053
rect 3905 945 3939 979
rect 3239 871 3273 905
rect 4867 945 4901 979
rect 3905 871 3939 905
rect 4867 871 4901 905
<< poly >>
rect 187 1404 217 1430
rect 275 1404 305 1430
rect 363 1404 393 1430
rect 451 1404 481 1430
rect 913 1404 943 1430
rect 1001 1404 1031 1430
rect 1089 1404 1119 1430
rect 1177 1404 1207 1430
rect 1265 1404 1295 1430
rect 1353 1404 1383 1430
rect 187 973 217 1004
rect 275 973 305 1004
rect 363 973 393 1004
rect 451 973 481 1004
rect 187 957 305 973
rect 187 943 205 957
rect 195 923 205 943
rect 239 943 305 957
rect 349 957 481 973
rect 239 923 249 943
rect 195 907 249 923
rect 349 923 359 957
rect 393 943 481 957
rect 1875 1404 1905 1430
rect 1963 1404 1993 1430
rect 2051 1404 2081 1430
rect 2139 1404 2169 1430
rect 2227 1404 2257 1430
rect 2315 1404 2345 1430
rect 913 973 943 1004
rect 1001 973 1031 1004
rect 1089 973 1119 1004
rect 1177 973 1207 1004
rect 393 923 403 943
rect 349 907 403 923
rect 861 957 1031 973
rect 861 923 871 957
rect 905 943 1031 957
rect 1083 957 1207 973
rect 905 923 915 943
rect 861 907 915 923
rect 1083 923 1093 957
rect 1127 943 1207 957
rect 1265 973 1295 1004
rect 1353 973 1383 1004
rect 1265 957 1383 973
rect 1265 943 1315 957
rect 1127 923 1137 943
rect 1083 907 1137 923
rect 1305 923 1315 943
rect 1349 943 1383 957
rect 2777 1404 2807 1430
rect 2865 1404 2895 1430
rect 2953 1404 2983 1430
rect 3041 1404 3071 1430
rect 1875 973 1905 1004
rect 1963 973 1993 1004
rect 2051 973 2081 1004
rect 2139 973 2169 1004
rect 1349 923 1359 943
rect 1305 907 1359 923
rect 1823 957 1993 973
rect 1823 923 1833 957
rect 1867 943 1993 957
rect 2045 957 2169 973
rect 1867 923 1877 943
rect 1823 907 1877 923
rect 2045 923 2055 957
rect 2089 943 2169 957
rect 2227 973 2257 1004
rect 2315 973 2345 1004
rect 2227 957 2345 973
rect 2227 943 2277 957
rect 2089 923 2099 943
rect 2045 907 2099 923
rect 2267 923 2277 943
rect 2311 943 2345 957
rect 3443 1404 3473 1430
rect 3531 1404 3561 1430
rect 3619 1404 3649 1430
rect 3707 1404 3737 1430
rect 2311 923 2321 943
rect 2267 907 2321 923
rect 2777 973 2807 1004
rect 2865 973 2895 1004
rect 2953 973 2983 1004
rect 3041 973 3071 1004
rect 2777 957 2895 973
rect 2777 943 2795 957
rect 2785 923 2795 943
rect 2829 943 2895 957
rect 2939 957 3071 973
rect 2829 923 2839 943
rect 2785 907 2839 923
rect 2939 923 2949 957
rect 2983 943 3071 957
rect 4169 1404 4199 1430
rect 4257 1404 4287 1430
rect 4345 1404 4375 1430
rect 4433 1404 4463 1430
rect 4521 1404 4551 1430
rect 4609 1404 4639 1430
rect 2983 923 2993 943
rect 2939 907 2993 923
rect 3443 973 3473 1004
rect 3531 973 3561 1004
rect 3619 973 3649 1004
rect 3707 973 3737 1004
rect 3443 957 3561 973
rect 3443 943 3461 957
rect 3451 923 3461 943
rect 3495 943 3561 957
rect 3605 957 3737 973
rect 3495 923 3505 943
rect 3451 907 3505 923
rect 3605 923 3615 957
rect 3649 943 3737 957
rect 4169 973 4199 1004
rect 4257 973 4287 1004
rect 4345 973 4375 1004
rect 4433 973 4463 1004
rect 3649 923 3659 943
rect 3605 907 3659 923
rect 4117 957 4287 973
rect 4117 923 4127 957
rect 4161 943 4287 957
rect 4339 957 4463 973
rect 4161 923 4171 943
rect 4117 907 4171 923
rect 4339 923 4349 957
rect 4383 943 4463 957
rect 4521 973 4551 1004
rect 4609 973 4639 1004
rect 4521 957 4639 973
rect 4521 943 4571 957
rect 4383 923 4393 943
rect 4339 907 4393 923
rect 4561 923 4571 943
rect 4605 943 4639 957
rect 4605 923 4615 943
rect 4561 907 4615 923
rect 195 433 249 449
rect 195 413 205 433
rect 168 399 205 413
rect 239 399 249 433
rect 168 383 249 399
rect 343 433 397 449
rect 343 399 353 433
rect 387 399 397 433
rect 343 383 397 399
rect 861 433 915 449
rect 861 413 871 433
rect 168 349 198 383
rect 362 349 392 383
rect 813 399 871 413
rect 905 399 915 433
rect 813 383 915 399
rect 1083 433 1137 449
rect 1083 399 1093 433
rect 1127 413 1137 433
rect 1305 433 1359 449
rect 1127 399 1143 413
rect 1083 383 1143 399
rect 1305 399 1315 433
rect 1349 399 1359 433
rect 1305 383 1359 399
rect 1823 433 1877 449
rect 1823 413 1833 433
rect 813 351 843 383
rect 1113 351 1143 383
rect 1315 351 1345 383
rect 1775 399 1833 413
rect 1867 399 1877 433
rect 1775 383 1877 399
rect 2045 433 2099 449
rect 2045 399 2055 433
rect 2089 413 2099 433
rect 2267 433 2321 449
rect 2089 399 2105 413
rect 2045 383 2105 399
rect 2267 399 2277 433
rect 2311 399 2321 433
rect 2267 383 2321 399
rect 2785 433 2839 449
rect 2785 413 2795 433
rect 1775 351 1805 383
rect 2075 351 2105 383
rect 2277 351 2307 383
rect 2758 399 2795 413
rect 2829 399 2839 433
rect 2758 383 2839 399
rect 2933 433 2987 449
rect 2933 399 2943 433
rect 2977 399 2987 433
rect 2933 383 2987 399
rect 3451 433 3505 449
rect 3451 413 3461 433
rect 2758 349 2788 383
rect 2952 349 2982 383
rect 3424 399 3461 413
rect 3495 399 3505 433
rect 3424 383 3505 399
rect 3599 433 3653 449
rect 3599 399 3609 433
rect 3643 399 3653 433
rect 3599 383 3653 399
rect 4117 433 4171 449
rect 4117 413 4127 433
rect 3424 349 3454 383
rect 3618 349 3648 383
rect 4069 399 4127 413
rect 4161 399 4171 433
rect 4069 383 4171 399
rect 4339 433 4393 449
rect 4339 399 4349 433
rect 4383 413 4393 433
rect 4561 433 4615 449
rect 4383 399 4399 413
rect 4339 383 4399 399
rect 4561 399 4571 433
rect 4605 399 4615 433
rect 4561 383 4615 399
rect 4069 351 4099 383
rect 4369 351 4399 383
rect 4571 351 4601 383
<< polycont >>
rect 205 923 239 957
rect 359 923 393 957
rect 871 923 905 957
rect 1093 923 1127 957
rect 1315 923 1349 957
rect 1833 923 1867 957
rect 2055 923 2089 957
rect 2277 923 2311 957
rect 2795 923 2829 957
rect 2949 923 2983 957
rect 3461 923 3495 957
rect 3615 923 3649 957
rect 4127 923 4161 957
rect 4349 923 4383 957
rect 4571 923 4605 957
rect 205 399 239 433
rect 353 399 387 433
rect 871 399 905 433
rect 1093 399 1127 433
rect 1315 399 1349 433
rect 1833 399 1867 433
rect 2055 399 2089 433
rect 2277 399 2311 433
rect 2795 399 2829 433
rect 2943 399 2977 433
rect 3461 399 3495 433
rect 3609 399 3643 433
rect 4127 399 4161 433
rect 4349 399 4383 433
rect 4571 399 4605 433
<< locali >>
rect -34 1497 4918 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4918 1497
rect -34 1446 4918 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 141 1366 175 1446
rect 141 1298 175 1332
rect 141 1230 175 1264
rect 141 1162 175 1196
rect 141 1093 175 1128
rect 141 1027 175 1059
rect 229 1366 263 1404
rect 229 1298 263 1332
rect 229 1230 263 1264
rect 229 1162 263 1196
rect 229 1093 263 1128
rect 317 1366 351 1446
rect 317 1298 351 1332
rect 317 1230 351 1264
rect 317 1162 351 1196
rect 317 1111 351 1128
rect 405 1366 439 1404
rect 405 1298 439 1332
rect 405 1230 439 1264
rect 405 1162 439 1196
rect 229 1057 263 1059
rect 405 1093 439 1128
rect 493 1366 527 1446
rect 493 1298 527 1332
rect 493 1230 527 1264
rect 493 1162 527 1196
rect 493 1111 527 1128
rect 632 1423 700 1446
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 405 1057 439 1059
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 229 1023 535 1057
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 359 957 393 973
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 923
rect 205 383 239 399
rect 353 923 359 942
rect 353 907 393 923
rect 353 831 387 907
rect 353 433 387 797
rect 353 383 387 399
rect 501 535 535 1023
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect 867 1366 901 1446
rect 867 1298 901 1332
rect 867 1230 901 1264
rect 867 1162 901 1196
rect 867 1093 901 1128
rect 867 1043 901 1059
rect 955 1366 989 1404
rect 955 1298 989 1332
rect 955 1230 989 1264
rect 955 1162 989 1196
rect 955 1093 989 1128
rect 1043 1366 1077 1446
rect 1043 1298 1077 1332
rect 1043 1230 1077 1264
rect 1043 1162 1077 1196
rect 1043 1111 1077 1128
rect 1131 1366 1165 1404
rect 1131 1298 1165 1332
rect 1131 1230 1165 1264
rect 1131 1162 1165 1196
rect 955 1048 989 1059
rect 1131 1093 1165 1128
rect 1219 1366 1253 1446
rect 1219 1298 1253 1332
rect 1219 1230 1253 1264
rect 1219 1162 1253 1196
rect 1219 1111 1253 1128
rect 1307 1366 1341 1404
rect 1307 1298 1341 1332
rect 1307 1230 1341 1264
rect 1307 1162 1341 1196
rect 1131 1048 1165 1059
rect 1307 1093 1341 1128
rect 1395 1366 1429 1446
rect 1395 1298 1429 1332
rect 1395 1230 1429 1264
rect 1395 1162 1429 1196
rect 1395 1111 1429 1128
rect 1594 1423 1662 1446
rect 1594 1389 1611 1423
rect 1645 1389 1662 1423
rect 1594 1349 1662 1389
rect 1594 1315 1611 1349
rect 1645 1315 1662 1349
rect 1594 1275 1662 1315
rect 1594 1241 1611 1275
rect 1645 1241 1662 1275
rect 1594 1201 1662 1241
rect 1594 1167 1611 1201
rect 1645 1167 1662 1201
rect 1594 1127 1662 1167
rect 1307 1048 1341 1059
rect 1594 1093 1611 1127
rect 1645 1093 1662 1127
rect 1594 1053 1662 1093
rect 632 979 700 1019
rect 955 1014 1497 1048
rect 632 945 649 979
rect 683 945 700 979
rect 632 905 700 945
rect 632 871 649 905
rect 683 871 700 905
rect 632 822 700 871
rect 871 957 905 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 122 333 156 349
rect 316 333 350 349
rect 501 348 535 501
rect 156 299 219 333
rect 253 299 316 333
rect 122 261 156 299
rect 122 193 156 227
rect 316 261 350 299
rect 122 123 156 159
rect 122 73 156 89
rect 219 208 253 224
rect -34 34 34 57
rect 219 34 253 174
rect 316 193 350 227
rect 413 314 535 348
rect 632 461 700 544
rect 632 427 649 461
rect 683 427 700 461
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect 871 534 905 923
rect 871 433 905 500
rect 871 383 905 399
rect 1093 957 1127 973
rect 1093 905 1127 923
rect 1093 433 1127 871
rect 1093 383 1127 399
rect 1315 957 1349 973
rect 1315 757 1349 923
rect 1463 847 1497 1014
rect 1462 831 1497 847
rect 1496 797 1497 831
rect 1594 1019 1611 1053
rect 1645 1019 1662 1053
rect 1829 1366 1863 1446
rect 1829 1298 1863 1332
rect 1829 1230 1863 1264
rect 1829 1162 1863 1196
rect 1829 1093 1863 1128
rect 1829 1043 1863 1059
rect 1917 1366 1951 1404
rect 1917 1298 1951 1332
rect 1917 1230 1951 1264
rect 1917 1162 1951 1196
rect 1917 1093 1951 1128
rect 2005 1366 2039 1446
rect 2005 1298 2039 1332
rect 2005 1230 2039 1264
rect 2005 1162 2039 1196
rect 2005 1111 2039 1128
rect 2093 1366 2127 1404
rect 2093 1298 2127 1332
rect 2093 1230 2127 1264
rect 2093 1162 2127 1196
rect 1917 1048 1951 1059
rect 2093 1093 2127 1128
rect 2181 1366 2215 1446
rect 2181 1298 2215 1332
rect 2181 1230 2215 1264
rect 2181 1162 2215 1196
rect 2181 1111 2215 1128
rect 2269 1366 2303 1404
rect 2269 1298 2303 1332
rect 2269 1230 2303 1264
rect 2269 1162 2303 1196
rect 2093 1048 2127 1059
rect 2269 1093 2303 1128
rect 2357 1366 2391 1446
rect 2357 1298 2391 1332
rect 2357 1230 2391 1264
rect 2357 1162 2391 1196
rect 2357 1111 2391 1128
rect 2556 1423 2624 1446
rect 2556 1389 2573 1423
rect 2607 1389 2624 1423
rect 2556 1349 2624 1389
rect 2556 1315 2573 1349
rect 2607 1315 2624 1349
rect 2556 1275 2624 1315
rect 2556 1241 2573 1275
rect 2607 1241 2624 1275
rect 2556 1201 2624 1241
rect 2556 1167 2573 1201
rect 2607 1167 2624 1201
rect 2556 1127 2624 1167
rect 2269 1048 2303 1059
rect 2556 1093 2573 1127
rect 2607 1093 2624 1127
rect 2556 1053 2624 1093
rect 1594 979 1662 1019
rect 1917 1014 2459 1048
rect 1594 945 1611 979
rect 1645 945 1662 979
rect 1594 905 1662 945
rect 1594 871 1611 905
rect 1645 871 1662 905
rect 1594 822 1662 871
rect 1833 957 1867 973
rect 1462 781 1497 797
rect 1315 433 1349 723
rect 1315 383 1349 399
rect 413 217 447 314
rect 632 313 700 353
rect 632 279 649 313
rect 683 279 700 313
rect 413 167 447 183
rect 510 261 544 277
rect 510 193 544 227
rect 316 123 350 159
rect 510 123 544 159
rect 350 89 413 123
rect 447 89 510 123
rect 316 73 350 89
rect 510 73 544 89
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect 632 57 649 91
rect 683 57 700 91
rect 767 335 801 351
rect 961 335 995 351
rect 1155 335 1189 351
rect 801 301 864 335
rect 898 301 961 335
rect 995 301 1058 335
rect 1092 301 1155 335
rect 767 263 801 301
rect 767 195 801 229
rect 961 263 995 301
rect 1155 285 1189 301
rect 1269 335 1303 351
rect 1463 350 1497 781
rect 1269 263 1303 301
rect 767 125 801 161
rect 767 75 801 91
rect 864 210 898 226
rect 632 34 700 57
rect 864 34 898 176
rect 961 195 995 229
rect 1059 216 1093 232
rect 1269 216 1303 229
rect 1093 195 1303 216
rect 1093 182 1269 195
rect 1059 166 1093 182
rect 961 125 995 161
rect 1366 316 1497 350
rect 1594 461 1662 544
rect 1594 427 1611 461
rect 1645 427 1662 461
rect 1594 387 1662 427
rect 1594 353 1611 387
rect 1645 353 1662 387
rect 1833 535 1867 923
rect 1833 433 1867 501
rect 1833 383 1867 399
rect 2055 957 2089 973
rect 2055 461 2089 923
rect 2055 383 2089 399
rect 2277 957 2311 973
rect 2277 757 2311 923
rect 2277 433 2311 723
rect 2277 383 2311 399
rect 2425 535 2459 1014
rect 2556 1019 2573 1053
rect 2607 1019 2624 1053
rect 2731 1366 2765 1446
rect 2731 1298 2765 1332
rect 2731 1230 2765 1264
rect 2731 1162 2765 1196
rect 2731 1093 2765 1128
rect 2731 1027 2765 1059
rect 2819 1366 2853 1404
rect 2819 1298 2853 1332
rect 2819 1230 2853 1264
rect 2819 1162 2853 1196
rect 2819 1093 2853 1128
rect 2907 1366 2941 1446
rect 2907 1298 2941 1332
rect 2907 1230 2941 1264
rect 2907 1162 2941 1196
rect 2907 1111 2941 1128
rect 2995 1366 3029 1404
rect 2995 1298 3029 1332
rect 2995 1230 3029 1264
rect 2995 1162 3029 1196
rect 2819 1057 2853 1059
rect 2995 1093 3029 1128
rect 3083 1366 3117 1446
rect 3083 1298 3117 1332
rect 3083 1230 3117 1264
rect 3083 1162 3117 1196
rect 3083 1111 3117 1128
rect 3222 1423 3290 1446
rect 3222 1389 3239 1423
rect 3273 1389 3290 1423
rect 3222 1349 3290 1389
rect 3222 1315 3239 1349
rect 3273 1315 3290 1349
rect 3222 1275 3290 1315
rect 3222 1241 3239 1275
rect 3273 1241 3290 1275
rect 3222 1201 3290 1241
rect 3222 1167 3239 1201
rect 3273 1167 3290 1201
rect 3222 1127 3290 1167
rect 2995 1057 3029 1059
rect 3222 1093 3239 1127
rect 3273 1093 3290 1127
rect 2819 1023 3125 1057
rect 2556 979 2624 1019
rect 2556 945 2573 979
rect 2607 945 2624 979
rect 2556 905 2624 945
rect 2556 871 2573 905
rect 2607 871 2624 905
rect 2556 822 2624 871
rect 2795 957 2829 973
rect 2949 957 2983 973
rect 1366 219 1400 316
rect 1594 313 1662 353
rect 1594 279 1611 313
rect 1645 279 1662 313
rect 1366 169 1400 185
rect 1463 263 1497 279
rect 1463 195 1497 229
rect 1155 125 1189 141
rect 995 91 1058 125
rect 1092 91 1155 125
rect 961 75 995 91
rect 1155 75 1189 91
rect 1269 125 1303 161
rect 1463 125 1497 161
rect 1303 91 1366 125
rect 1400 91 1463 125
rect 1269 75 1303 91
rect 1463 75 1497 91
rect 1594 239 1662 279
rect 1594 205 1611 239
rect 1645 205 1662 239
rect 1594 165 1662 205
rect 1594 131 1611 165
rect 1645 131 1662 165
rect 1594 91 1662 131
rect 1594 57 1611 91
rect 1645 57 1662 91
rect 1729 335 1763 351
rect 1923 335 1957 351
rect 2117 335 2151 351
rect 1763 301 1826 335
rect 1860 301 1923 335
rect 1957 301 2020 335
rect 2054 301 2117 335
rect 1729 263 1763 301
rect 1729 195 1763 229
rect 1923 263 1957 301
rect 2117 285 2151 301
rect 2231 335 2265 351
rect 2425 350 2459 501
rect 2231 263 2265 301
rect 1729 125 1763 161
rect 1729 75 1763 91
rect 1826 210 1860 226
rect 1594 34 1662 57
rect 1826 34 1860 176
rect 1923 195 1957 229
rect 2021 216 2055 232
rect 2231 216 2265 229
rect 2055 195 2265 216
rect 2055 182 2231 195
rect 2021 166 2055 182
rect 1923 125 1957 161
rect 2328 316 2459 350
rect 2556 461 2624 544
rect 2556 427 2573 461
rect 2607 427 2624 461
rect 2556 387 2624 427
rect 2556 353 2573 387
rect 2607 353 2624 387
rect 2795 535 2829 923
rect 2795 433 2829 501
rect 2795 383 2829 399
rect 2943 923 2949 942
rect 2943 907 2983 923
rect 2943 905 2977 907
rect 2943 433 2977 871
rect 2943 383 2977 399
rect 3091 757 3125 1023
rect 3222 1053 3290 1093
rect 3222 1019 3239 1053
rect 3273 1019 3290 1053
rect 3397 1366 3431 1446
rect 3397 1298 3431 1332
rect 3397 1230 3431 1264
rect 3397 1162 3431 1196
rect 3397 1093 3431 1128
rect 3397 1027 3431 1059
rect 3485 1366 3519 1404
rect 3485 1298 3519 1332
rect 3485 1230 3519 1264
rect 3485 1162 3519 1196
rect 3485 1093 3519 1128
rect 3573 1366 3607 1446
rect 3573 1298 3607 1332
rect 3573 1230 3607 1264
rect 3573 1162 3607 1196
rect 3573 1111 3607 1128
rect 3661 1366 3695 1404
rect 3661 1298 3695 1332
rect 3661 1230 3695 1264
rect 3661 1162 3695 1196
rect 3485 1057 3519 1059
rect 3661 1093 3695 1128
rect 3749 1366 3783 1446
rect 3749 1298 3783 1332
rect 3749 1230 3783 1264
rect 3749 1162 3783 1196
rect 3749 1111 3783 1128
rect 3888 1423 3956 1446
rect 3888 1389 3905 1423
rect 3939 1389 3956 1423
rect 3888 1349 3956 1389
rect 3888 1315 3905 1349
rect 3939 1315 3956 1349
rect 3888 1275 3956 1315
rect 3888 1241 3905 1275
rect 3939 1241 3956 1275
rect 3888 1201 3956 1241
rect 3888 1167 3905 1201
rect 3939 1167 3956 1201
rect 3888 1127 3956 1167
rect 3661 1057 3695 1059
rect 3888 1093 3905 1127
rect 3939 1093 3956 1127
rect 3485 1023 3791 1057
rect 3222 979 3290 1019
rect 3222 945 3239 979
rect 3273 945 3290 979
rect 3222 905 3290 945
rect 3222 871 3239 905
rect 3273 871 3290 905
rect 3222 822 3290 871
rect 3461 957 3495 973
rect 3615 957 3649 973
rect 3461 831 3495 923
rect 2328 219 2362 316
rect 2556 313 2624 353
rect 2556 279 2573 313
rect 2607 279 2624 313
rect 2328 169 2362 185
rect 2425 263 2459 279
rect 2425 195 2459 229
rect 2117 125 2151 141
rect 1957 91 2020 125
rect 2054 91 2117 125
rect 1923 75 1957 91
rect 2117 75 2151 91
rect 2231 125 2265 161
rect 2425 125 2459 161
rect 2265 91 2328 125
rect 2362 91 2425 125
rect 2231 75 2265 91
rect 2425 75 2459 91
rect 2556 239 2624 279
rect 2556 205 2573 239
rect 2607 205 2624 239
rect 2556 165 2624 205
rect 2556 131 2573 165
rect 2607 131 2624 165
rect 2556 91 2624 131
rect 2556 57 2573 91
rect 2607 57 2624 91
rect 2712 333 2746 349
rect 2906 333 2940 349
rect 3091 348 3125 723
rect 2746 299 2809 333
rect 2843 299 2906 333
rect 2712 261 2746 299
rect 2712 193 2746 227
rect 2906 261 2940 299
rect 2712 123 2746 159
rect 2712 73 2746 89
rect 2809 208 2843 224
rect 2556 34 2624 57
rect 2809 34 2843 174
rect 2906 193 2940 227
rect 3003 314 3125 348
rect 3222 461 3290 544
rect 3222 427 3239 461
rect 3273 427 3290 461
rect 3222 387 3290 427
rect 3222 353 3239 387
rect 3273 353 3290 387
rect 3461 433 3495 797
rect 3461 383 3495 399
rect 3609 923 3615 942
rect 3609 907 3649 923
rect 3609 683 3643 907
rect 3609 433 3643 649
rect 3609 383 3643 399
rect 3757 609 3791 1023
rect 3888 1053 3956 1093
rect 3888 1019 3905 1053
rect 3939 1019 3956 1053
rect 4123 1366 4157 1446
rect 4123 1298 4157 1332
rect 4123 1230 4157 1264
rect 4123 1162 4157 1196
rect 4123 1093 4157 1128
rect 4123 1043 4157 1059
rect 4211 1366 4245 1404
rect 4211 1298 4245 1332
rect 4211 1230 4245 1264
rect 4211 1162 4245 1196
rect 4211 1093 4245 1128
rect 4299 1366 4333 1446
rect 4299 1298 4333 1332
rect 4299 1230 4333 1264
rect 4299 1162 4333 1196
rect 4299 1111 4333 1128
rect 4387 1366 4421 1404
rect 4387 1298 4421 1332
rect 4387 1230 4421 1264
rect 4387 1162 4421 1196
rect 4211 1048 4245 1059
rect 4387 1093 4421 1128
rect 4475 1366 4509 1446
rect 4475 1298 4509 1332
rect 4475 1230 4509 1264
rect 4475 1162 4509 1196
rect 4475 1111 4509 1128
rect 4563 1366 4597 1404
rect 4563 1298 4597 1332
rect 4563 1230 4597 1264
rect 4563 1162 4597 1196
rect 4387 1048 4421 1059
rect 4563 1093 4597 1128
rect 4651 1366 4685 1446
rect 4651 1298 4685 1332
rect 4651 1230 4685 1264
rect 4651 1162 4685 1196
rect 4651 1111 4685 1128
rect 4850 1423 4918 1446
rect 4850 1389 4867 1423
rect 4901 1389 4918 1423
rect 4850 1349 4918 1389
rect 4850 1315 4867 1349
rect 4901 1315 4918 1349
rect 4850 1275 4918 1315
rect 4850 1241 4867 1275
rect 4901 1241 4918 1275
rect 4850 1201 4918 1241
rect 4850 1167 4867 1201
rect 4901 1167 4918 1201
rect 4850 1127 4918 1167
rect 4563 1048 4597 1059
rect 4850 1093 4867 1127
rect 4901 1093 4918 1127
rect 4850 1053 4918 1093
rect 3888 979 3956 1019
rect 4211 1014 4753 1048
rect 3888 945 3905 979
rect 3939 945 3956 979
rect 3888 905 3956 945
rect 3888 871 3905 905
rect 3939 871 3956 905
rect 3888 822 3956 871
rect 4127 957 4161 973
rect 3003 217 3037 314
rect 3222 313 3290 353
rect 3222 279 3239 313
rect 3273 279 3290 313
rect 3003 167 3037 183
rect 3100 261 3134 277
rect 3100 193 3134 227
rect 2906 123 2940 159
rect 3100 123 3134 159
rect 2940 89 3003 123
rect 3037 89 3100 123
rect 2906 73 2940 89
rect 3100 73 3134 89
rect 3222 239 3290 279
rect 3222 205 3239 239
rect 3273 205 3290 239
rect 3222 165 3290 205
rect 3222 131 3239 165
rect 3273 131 3290 165
rect 3222 91 3290 131
rect 3222 57 3239 91
rect 3273 57 3290 91
rect 3378 333 3412 349
rect 3572 333 3606 349
rect 3757 348 3791 575
rect 4127 609 4161 923
rect 3412 299 3475 333
rect 3509 299 3572 333
rect 3378 261 3412 299
rect 3378 193 3412 227
rect 3572 261 3606 299
rect 3378 123 3412 159
rect 3378 73 3412 89
rect 3475 208 3509 224
rect 3222 34 3290 57
rect 3475 34 3509 174
rect 3572 193 3606 227
rect 3669 314 3791 348
rect 3888 461 3956 544
rect 3888 427 3905 461
rect 3939 427 3956 461
rect 3888 387 3956 427
rect 3888 353 3905 387
rect 3939 353 3956 387
rect 4127 433 4161 575
rect 4127 383 4161 399
rect 4349 957 4383 973
rect 4349 461 4383 923
rect 4349 383 4383 399
rect 4571 957 4605 973
rect 4571 757 4605 923
rect 4571 433 4605 723
rect 4571 383 4605 399
rect 4719 683 4753 1014
rect 4850 1019 4867 1053
rect 4901 1019 4918 1053
rect 4850 979 4918 1019
rect 4850 945 4867 979
rect 4901 945 4918 979
rect 4850 905 4918 945
rect 4850 871 4867 905
rect 4901 871 4918 905
rect 4850 822 4918 871
rect 3669 217 3703 314
rect 3888 313 3956 353
rect 3888 279 3905 313
rect 3939 279 3956 313
rect 3669 167 3703 183
rect 3766 261 3800 277
rect 3766 193 3800 227
rect 3572 123 3606 159
rect 3766 123 3800 159
rect 3606 89 3669 123
rect 3703 89 3766 123
rect 3572 73 3606 89
rect 3766 73 3800 89
rect 3888 239 3956 279
rect 3888 205 3905 239
rect 3939 205 3956 239
rect 3888 165 3956 205
rect 3888 131 3905 165
rect 3939 131 3956 165
rect 3888 91 3956 131
rect 3888 57 3905 91
rect 3939 57 3956 91
rect 4023 335 4057 351
rect 4217 335 4251 351
rect 4411 335 4445 351
rect 4057 301 4120 335
rect 4154 301 4217 335
rect 4251 301 4314 335
rect 4348 301 4411 335
rect 4023 263 4057 301
rect 4023 195 4057 229
rect 4217 263 4251 301
rect 4411 285 4445 301
rect 4525 335 4559 351
rect 4719 350 4753 649
rect 4525 263 4559 301
rect 4023 125 4057 161
rect 4023 75 4057 91
rect 4120 210 4154 226
rect 3888 34 3956 57
rect 4120 34 4154 176
rect 4217 195 4251 229
rect 4315 216 4349 232
rect 4525 216 4559 229
rect 4349 195 4559 216
rect 4349 182 4525 195
rect 4315 166 4349 182
rect 4217 125 4251 161
rect 4622 316 4753 350
rect 4850 461 4918 544
rect 4850 427 4867 461
rect 4901 427 4918 461
rect 4850 387 4918 427
rect 4850 353 4867 387
rect 4901 353 4918 387
rect 4622 219 4656 316
rect 4850 313 4918 353
rect 4850 279 4867 313
rect 4901 279 4918 313
rect 4622 169 4656 185
rect 4719 263 4753 279
rect 4719 195 4753 229
rect 4411 125 4445 141
rect 4251 91 4314 125
rect 4348 91 4411 125
rect 4217 75 4251 91
rect 4411 75 4445 91
rect 4525 125 4559 161
rect 4719 125 4753 161
rect 4559 91 4622 125
rect 4656 91 4719 125
rect 4525 75 4559 91
rect 4719 75 4753 91
rect 4850 239 4918 279
rect 4850 205 4867 239
rect 4901 205 4918 239
rect 4850 165 4918 205
rect 4850 131 4867 165
rect 4901 131 4918 165
rect 4850 91 4918 131
rect 4850 57 4867 91
rect 4901 57 4918 91
rect 4850 34 4918 57
rect -34 17 4918 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4918 17
rect -34 -34 4918 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 353 797 387 831
rect 501 501 535 535
rect 871 500 905 534
rect 1093 871 1127 905
rect 1462 797 1496 831
rect 1315 723 1349 757
rect 1833 501 1867 535
rect 2055 433 2089 461
rect 2055 427 2089 433
rect 2277 723 2311 757
rect 2425 501 2459 535
rect 2795 501 2829 535
rect 2943 871 2977 905
rect 3091 723 3125 757
rect 3461 797 3495 831
rect 3609 649 3643 683
rect 3757 575 3791 609
rect 4127 575 4161 609
rect 4349 433 4383 461
rect 4349 427 4383 433
rect 4571 723 4605 757
rect 4719 649 4753 683
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
<< metal1 >>
rect -34 1497 4918 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4918 1497
rect -34 1446 4918 1463
rect 1087 905 1133 911
rect 2937 905 2983 911
rect 1081 871 1093 905
rect 1127 871 2943 905
rect 2977 871 2989 905
rect 1087 865 1133 871
rect 2937 865 2983 871
rect 347 831 393 837
rect 1456 831 1502 837
rect 3455 831 3501 837
rect 341 797 353 831
rect 387 797 1462 831
rect 1496 797 3461 831
rect 3495 797 3507 831
rect 347 791 393 797
rect 1456 791 1502 797
rect 3455 791 3501 797
rect 1309 757 1355 763
rect 2271 757 2317 763
rect 3085 757 3131 763
rect 4565 757 4611 763
rect 1303 723 1315 757
rect 1349 723 2277 757
rect 2311 723 3091 757
rect 3125 723 4571 757
rect 4605 723 4617 757
rect 1309 717 1355 723
rect 2271 717 2317 723
rect 3085 717 3131 723
rect 4565 717 4611 723
rect 3603 683 3649 689
rect 4713 683 4759 689
rect 3597 649 3609 683
rect 3643 649 4719 683
rect 4753 649 4765 683
rect 3603 643 3649 649
rect 4713 643 4759 649
rect 3751 609 3797 615
rect 4121 609 4167 615
rect 3745 575 3757 609
rect 3791 575 4127 609
rect 4161 575 4173 609
rect 3751 569 3797 575
rect 4121 569 4167 575
rect 495 535 541 541
rect 865 535 911 540
rect 1827 535 1873 541
rect 2419 535 2465 541
rect 2789 535 2835 541
rect 489 501 501 535
rect 535 534 1833 535
rect 535 501 871 534
rect 495 495 541 501
rect 859 500 871 501
rect 905 501 1833 534
rect 1867 501 1879 535
rect 2413 501 2425 535
rect 2459 501 2795 535
rect 2829 501 2841 535
rect 905 500 941 501
rect 865 494 911 500
rect 1827 495 1873 501
rect 2419 495 2465 501
rect 2789 495 2835 501
rect 2049 461 2095 467
rect 4343 461 4389 467
rect 2043 427 2055 461
rect 2089 427 4349 461
rect 4383 427 4395 461
rect 2049 421 2095 427
rect 4343 421 4389 427
rect -34 17 4918 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4918 17
rect -34 -34 4918 -17
<< labels >>
rlabel metal1 4127 575 4161 609 1 QN
port 1 n
rlabel metal1 4127 797 4161 831 1 QN
port 2 n
rlabel metal1 4127 871 4161 905 1 QN
port 3 n
rlabel metal1 4127 501 4161 535 1 QN
port 4 n
rlabel metal1 3757 501 3791 535 1 QN
port 5 n
rlabel metal1 3757 575 3791 609 1 QN
port 6 n
rlabel metal1 3757 797 3791 831 1 QN
port 7 n
rlabel metal1 3757 871 3791 905 1 QN
port 8 n
rlabel metal1 3757 945 3791 979 1 QN
port 9 n
rlabel metal1 205 723 239 757 1 D
port 10 n
rlabel metal1 205 649 239 683 1 D
port 11 n
rlabel metal1 205 575 239 609 1 D
port 12 n
rlabel metal1 205 501 239 535 1 D
port 13 n
rlabel metal1 205 427 239 461 1 D
port 14 n
rlabel metal1 205 797 239 831 1 D
port 15 n
rlabel metal1 205 871 239 905 1 D
port 16 n
rlabel metal1 1093 871 1127 905 1 CLK
port 17 n
rlabel metal1 1093 723 1127 757 1 CLK
port 18 n
rlabel metal1 1093 649 1127 683 1 CLK
port 19 n
rlabel metal1 1093 575 1127 609 1 CLK
port 20 n
rlabel metal1 2943 575 2977 609 1 CLK
port 21 n
rlabel metal1 2943 649 2977 683 1 CLK
port 22 n
rlabel metal1 2943 871 2977 905 1 CLK
port 23 n
rlabel metal1 2943 501 2977 535 1 CLK
port 24 n
rlabel metal1 2055 427 2089 461 1 SN
port 25 n
rlabel metal1 2055 501 2089 535 1 SN
port 26 n
rlabel metal1 2055 575 2089 609 1 SN
port 27 n
rlabel metal1 2055 649 2089 683 1 SN
port 28 n
rlabel metal1 4349 427 4383 461 1 SN
port 29 n
rlabel metal1 4349 501 4383 535 1 SN
port 30 n
rlabel metal1 4349 575 4383 609 1 SN
port 31 n
rlabel metal1 4349 797 4383 831 1 SN
port 32 n
rlabel metal1 4349 871 4383 905 1 SN
port 33 n
rlabel metal1 -34 1446 4918 1514 1 VPWR
port 34 n
rlabel metal1 -34 -34 4918 34 1 VGND
port 35 n
rlabel nwell 57 1463 91 1497 1 VPB
port 36 n
rlabel pwell 57 -17 91 17 1 VNB
port 37 n
<< end >>
