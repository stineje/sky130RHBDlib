* SPICE3 file created from AND2X1.ext - technology: sky130A

.subckt AND2X1 Y A B VDD GND
X0 VDD B a_217_1004 VDD pshort w=2 l=0.15 M=2
X1 GND A a_112_73 GND nshort w=3 l=0.15
X2 Y a_217_1004 GND GND nshort w=3 l=0.15
X3 VDD a_217_1004 Y VDD pshort w=2 l=0.15 M=2
X4 a_217_1004 A VDD VDD pshort w=2 l=0.15 M=2
X5 a_217_1004 B a_112_73 GND nshort w=3 l=0.15
C0 VDD GND 3.02fF
.ends
