* SPICE3 file created from DFFSNRNQX1.ext - technology: sky130A

.subckt DFFSNRNQX1 Q D CLK SN RN VPB VNB
M1000 Q SN VPB.t24 pshort w=2u l=0.15u
+  ad=1.74p pd=13.74u as=0p ps=0u
M1001 VNB a_4125_1004.t8 a_4901_75.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1002 VPB.t28 a_147_159# a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_599_943.t4 CLK VPB.t32 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPB.t33 CLK a_1561_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t7 a_277_1004.t7 a_2201_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t6 RN a_277_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_599_943.t0 a_1561_943.t8 VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t22 SN a_2201_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPB.t5 RN a_1561_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_4125_1004.t6 a_599_943.t7 VPB.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1561_943.t3 CLK VPB.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_4125_1004.t3 Q VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VNB a_147_159# a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPB.t10 a_599_943.t8 a_277_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_1561_943.t10 a_5182_182.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1016 a_4125_1004.t1 RN VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t8 a_1561_943.t11 a_2201_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1561_943.t6 a_2201_1004.t8 VPB.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPB.t11 a_4125_1004.t7 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_277_1004.t5 a_147_159# VPB.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPB.t16 a_277_1004.t10 a_599_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t25 a_1561_943.t12 a_599_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPB.t23 SN Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VNB a_277_1004.t8 a_2015_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_277_1004.t0 RN VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPB.t30 CLK a_599_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_2201_1004.t0 SN VPB.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1561_943.t0 RN VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB.t2 RN a_4125_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPB.t12 a_1561_943.t13 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_599_943.t5 a_277_1004.t11 VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_277_1004.t2 a_599_943.t10 VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 VNB a_2201_1004.t7 a_2977_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1034 VNB a_277_1004.t9 a_1053_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_2201_1004.t5 a_277_1004.t12 VPB.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_2201_1004.t3 a_1561_943.t14 VPB.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPB.t26 a_599_943.t12 a_4125_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPB.t17 Q a_4125_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 Q a_4125_1004.t9 VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 Q a_1561_943.t15 VPB.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VNB a_599_943.t9 a_3939_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPB.t34 a_2201_1004.t9 a_1561_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB a_147_159# 0.08fF
C1 SN Q 0.38fF
C2 SN CLK 0.48fF
C3 RN Q 0.18fF
C4 RN CLK 0.73fF
C5 SN RN 0.37fF
C6 VPB Q 1.83fF
C7 CLK VPB 0.10fF
C8 RN a_147_159# 0.18fF
C9 SN VPB 0.10fF
C10 RN VPB 1.10fF
R0 VPB VPB.n513 126.832
R1 VPB.n40 VPB.n38 94.117
R2 VPB.n435 VPB.n433 94.117
R3 VPB.n352 VPB.n350 94.117
R4 VPB.n129 VPB.n127 94.117
R5 VPB.n275 VPB.n273 94.117
R6 VPB.n199 VPB.n198 84.554
R7 VPB.n288 VPB.n287 80.104
R8 VPB.n139 VPB.n138 80.104
R9 VPB.n365 VPB.n364 80.104
R10 VPB.n448 VPB.n447 80.104
R11 VPB.n50 VPB.n49 80.104
R12 VPB.n215 VPB.n214 76
R13 VPB.n220 VPB.n219 76
R14 VPB.n225 VPB.n224 76
R15 VPB.n232 VPB.n231 76
R16 VPB.n237 VPB.n236 76
R17 VPB.n242 VPB.n241 76
R18 VPB.n246 VPB.n245 76
R19 VPB.n250 VPB.n249 76
R20 VPB.n277 VPB.n276 76
R21 VPB.n281 VPB.n280 76
R22 VPB.n286 VPB.n285 76
R23 VPB.n291 VPB.n290 76
R24 VPB.n298 VPB.n297 76
R25 VPB.n303 VPB.n302 76
R26 VPB.n308 VPB.n307 76
R27 VPB.n315 VPB.n314 76
R28 VPB.n320 VPB.n319 76
R29 VPB.n325 VPB.n324 76
R30 VPB.n329 VPB.n328 76
R31 VPB.n333 VPB.n332 76
R32 VPB.n348 VPB.n345 76
R33 VPB.n354 VPB.n353 76
R34 VPB.n358 VPB.n357 76
R35 VPB.n363 VPB.n362 76
R36 VPB.n368 VPB.n367 76
R37 VPB.n375 VPB.n374 76
R38 VPB.n380 VPB.n379 76
R39 VPB.n385 VPB.n384 76
R40 VPB.n392 VPB.n391 76
R41 VPB.n397 VPB.n396 76
R42 VPB.n402 VPB.n401 76
R43 VPB.n406 VPB.n405 76
R44 VPB.n410 VPB.n409 76
R45 VPB.n437 VPB.n436 76
R46 VPB.n441 VPB.n440 76
R47 VPB.n446 VPB.n445 76
R48 VPB.n451 VPB.n450 76
R49 VPB.n458 VPB.n457 76
R50 VPB.n463 VPB.n462 76
R51 VPB.n468 VPB.n467 76
R52 VPB.n475 VPB.n474 76
R53 VPB.n480 VPB.n479 76
R54 VPB.n485 VPB.n484 76
R55 VPB.n489 VPB.n488 76
R56 VPB.n493 VPB.n492 76
R57 VPB.n506 VPB.n505 76
R58 VPB.n234 VPB.n233 75.654
R59 VPB.n317 VPB.n316 75.654
R60 VPB.n161 VPB.n160 75.654
R61 VPB.n394 VPB.n393 75.654
R62 VPB.n477 VPB.n476 75.654
R63 VPB.n72 VPB.n71 75.654
R64 VPB.n22 VPB.n21 61.764
R65 VPB.n417 VPB.n416 61.764
R66 VPB.n88 VPB.n87 61.764
R67 VPB.n111 VPB.n110 61.764
R68 VPB.n257 VPB.n256 61.764
R69 VPB.n78 VPB.t29 55.106
R70 VPB.n481 VPB.t20 55.106
R71 VPB.n398 VPB.t19 55.106
R72 VPB.n167 VPB.t35 55.106
R73 VPB.n321 VPB.t27 55.106
R74 VPB.n238 VPB.t0 55.106
R75 VPB.n45 VPB.t10 55.106
R76 VPB.n442 VPB.t25 55.106
R77 VPB.n359 VPB.t8 55.106
R78 VPB.n134 VPB.t5 55.106
R79 VPB.n282 VPB.t17 55.106
R80 VPB.n202 VPB.t12 55.106
R81 VPB.n212 VPB.n211 48.952
R82 VPB.n295 VPB.n294 48.952
R83 VPB.n143 VPB.n142 48.952
R84 VPB.n372 VPB.n371 48.952
R85 VPB.n455 VPB.n454 48.952
R86 VPB.n54 VPB.n53 48.952
R87 VPB.n229 VPB.n228 44.502
R88 VPB.n312 VPB.n311 44.502
R89 VPB.n157 VPB.n156 44.502
R90 VPB.n389 VPB.n388 44.502
R91 VPB.n472 VPB.n471 44.502
R92 VPB.n68 VPB.n67 44.502
R93 VPB.n66 VPB.n14 40.824
R94 VPB.n57 VPB.n15 40.824
R95 VPB.n470 VPB.n469 40.824
R96 VPB.n453 VPB.n452 40.824
R97 VPB.n387 VPB.n386 40.824
R98 VPB.n370 VPB.n369 40.824
R99 VPB.n155 VPB.n103 40.824
R100 VPB.n146 VPB.n104 40.824
R101 VPB.n310 VPB.n309 40.824
R102 VPB.n293 VPB.n292 40.824
R103 VPB.n227 VPB.n226 40.824
R104 VPB.n210 VPB.n209 40.824
R105 VPB.n207 VPB.n206 35.118
R106 VPB.n510 VPB.n506 20.452
R107 VPB.n194 VPB.n191 20.452
R108 VPB.n217 VPB.n216 17.801
R109 VPB.n300 VPB.n299 17.801
R110 VPB.n148 VPB.n147 17.801
R111 VPB.n377 VPB.n376 17.801
R112 VPB.n460 VPB.n459 17.801
R113 VPB.n59 VPB.n58 17.801
R114 VPB.n14 VPB.t1 14.282
R115 VPB.n14 VPB.t28 14.282
R116 VPB.n15 VPB.t9 14.282
R117 VPB.n15 VPB.t6 14.282
R118 VPB.n469 VPB.t32 14.282
R119 VPB.n469 VPB.t16 14.282
R120 VPB.n452 VPB.t14 14.282
R121 VPB.n452 VPB.t30 14.282
R122 VPB.n386 VPB.t21 14.282
R123 VPB.n386 VPB.t7 14.282
R124 VPB.n369 VPB.t13 14.282
R125 VPB.n369 VPB.t22 14.282
R126 VPB.n103 VPB.t31 14.282
R127 VPB.n103 VPB.t34 14.282
R128 VPB.n104 VPB.t4 14.282
R129 VPB.n104 VPB.t33 14.282
R130 VPB.n309 VPB.t3 14.282
R131 VPB.n309 VPB.t26 14.282
R132 VPB.n292 VPB.t18 14.282
R133 VPB.n292 VPB.t2 14.282
R134 VPB.n226 VPB.t24 14.282
R135 VPB.n226 VPB.t11 14.282
R136 VPB.n209 VPB.t15 14.282
R137 VPB.n209 VPB.t23 14.282
R138 VPB.n194 VPB.n193 13.653
R139 VPB.n193 VPB.n192 13.653
R140 VPB.n205 VPB.n204 13.653
R141 VPB.n204 VPB.n203 13.653
R142 VPB.n201 VPB.n200 13.653
R143 VPB.n200 VPB.n199 13.653
R144 VPB.n197 VPB.n196 13.653
R145 VPB.n196 VPB.n195 13.653
R146 VPB.n214 VPB.n213 13.653
R147 VPB.n213 VPB.n212 13.653
R148 VPB.n219 VPB.n218 13.653
R149 VPB.n218 VPB.n217 13.653
R150 VPB.n224 VPB.n223 13.653
R151 VPB.n223 VPB.n222 13.653
R152 VPB.n231 VPB.n230 13.653
R153 VPB.n230 VPB.n229 13.653
R154 VPB.n236 VPB.n235 13.653
R155 VPB.n235 VPB.n234 13.653
R156 VPB.n241 VPB.n240 13.653
R157 VPB.n240 VPB.n239 13.653
R158 VPB.n245 VPB.n244 13.653
R159 VPB.n244 VPB.n243 13.653
R160 VPB.n249 VPB.n248 13.653
R161 VPB.n248 VPB.n247 13.653
R162 VPB.n276 VPB.n275 13.653
R163 VPB.n275 VPB.n274 13.653
R164 VPB.n280 VPB.n279 13.653
R165 VPB.n279 VPB.n278 13.653
R166 VPB.n285 VPB.n284 13.653
R167 VPB.n284 VPB.n283 13.653
R168 VPB.n290 VPB.n289 13.653
R169 VPB.n289 VPB.n288 13.653
R170 VPB.n297 VPB.n296 13.653
R171 VPB.n296 VPB.n295 13.653
R172 VPB.n302 VPB.n301 13.653
R173 VPB.n301 VPB.n300 13.653
R174 VPB.n307 VPB.n306 13.653
R175 VPB.n306 VPB.n305 13.653
R176 VPB.n314 VPB.n313 13.653
R177 VPB.n313 VPB.n312 13.653
R178 VPB.n319 VPB.n318 13.653
R179 VPB.n318 VPB.n317 13.653
R180 VPB.n324 VPB.n323 13.653
R181 VPB.n323 VPB.n322 13.653
R182 VPB.n328 VPB.n327 13.653
R183 VPB.n327 VPB.n326 13.653
R184 VPB.n332 VPB.n331 13.653
R185 VPB.n331 VPB.n330 13.653
R186 VPB.n130 VPB.n129 13.653
R187 VPB.n129 VPB.n128 13.653
R188 VPB.n133 VPB.n132 13.653
R189 VPB.n132 VPB.n131 13.653
R190 VPB.n137 VPB.n136 13.653
R191 VPB.n136 VPB.n135 13.653
R192 VPB.n141 VPB.n140 13.653
R193 VPB.n140 VPB.n139 13.653
R194 VPB.n145 VPB.n144 13.653
R195 VPB.n144 VPB.n143 13.653
R196 VPB.n150 VPB.n149 13.653
R197 VPB.n149 VPB.n148 13.653
R198 VPB.n154 VPB.n153 13.653
R199 VPB.n153 VPB.n152 13.653
R200 VPB.n159 VPB.n158 13.653
R201 VPB.n158 VPB.n157 13.653
R202 VPB.n163 VPB.n162 13.653
R203 VPB.n162 VPB.n161 13.653
R204 VPB.n166 VPB.n165 13.653
R205 VPB.n165 VPB.n164 13.653
R206 VPB.n170 VPB.n169 13.653
R207 VPB.n169 VPB.n168 13.653
R208 VPB.n348 VPB.n347 13.653
R209 VPB.n347 VPB.n346 13.653
R210 VPB.n353 VPB.n352 13.653
R211 VPB.n352 VPB.n351 13.653
R212 VPB.n357 VPB.n356 13.653
R213 VPB.n356 VPB.n355 13.653
R214 VPB.n362 VPB.n361 13.653
R215 VPB.n361 VPB.n360 13.653
R216 VPB.n367 VPB.n366 13.653
R217 VPB.n366 VPB.n365 13.653
R218 VPB.n374 VPB.n373 13.653
R219 VPB.n373 VPB.n372 13.653
R220 VPB.n379 VPB.n378 13.653
R221 VPB.n378 VPB.n377 13.653
R222 VPB.n384 VPB.n383 13.653
R223 VPB.n383 VPB.n382 13.653
R224 VPB.n391 VPB.n390 13.653
R225 VPB.n390 VPB.n389 13.653
R226 VPB.n396 VPB.n395 13.653
R227 VPB.n395 VPB.n394 13.653
R228 VPB.n401 VPB.n400 13.653
R229 VPB.n400 VPB.n399 13.653
R230 VPB.n405 VPB.n404 13.653
R231 VPB.n404 VPB.n403 13.653
R232 VPB.n409 VPB.n408 13.653
R233 VPB.n408 VPB.n407 13.653
R234 VPB.n436 VPB.n435 13.653
R235 VPB.n435 VPB.n434 13.653
R236 VPB.n440 VPB.n439 13.653
R237 VPB.n439 VPB.n438 13.653
R238 VPB.n445 VPB.n444 13.653
R239 VPB.n444 VPB.n443 13.653
R240 VPB.n450 VPB.n449 13.653
R241 VPB.n449 VPB.n448 13.653
R242 VPB.n457 VPB.n456 13.653
R243 VPB.n456 VPB.n455 13.653
R244 VPB.n462 VPB.n461 13.653
R245 VPB.n461 VPB.n460 13.653
R246 VPB.n467 VPB.n466 13.653
R247 VPB.n466 VPB.n465 13.653
R248 VPB.n474 VPB.n473 13.653
R249 VPB.n473 VPB.n472 13.653
R250 VPB.n479 VPB.n478 13.653
R251 VPB.n478 VPB.n477 13.653
R252 VPB.n484 VPB.n483 13.653
R253 VPB.n483 VPB.n482 13.653
R254 VPB.n488 VPB.n487 13.653
R255 VPB.n487 VPB.n486 13.653
R256 VPB.n492 VPB.n491 13.653
R257 VPB.n491 VPB.n490 13.653
R258 VPB.n41 VPB.n40 13.653
R259 VPB.n40 VPB.n39 13.653
R260 VPB.n44 VPB.n43 13.653
R261 VPB.n43 VPB.n42 13.653
R262 VPB.n48 VPB.n47 13.653
R263 VPB.n47 VPB.n46 13.653
R264 VPB.n52 VPB.n51 13.653
R265 VPB.n51 VPB.n50 13.653
R266 VPB.n56 VPB.n55 13.653
R267 VPB.n55 VPB.n54 13.653
R268 VPB.n61 VPB.n60 13.653
R269 VPB.n60 VPB.n59 13.653
R270 VPB.n65 VPB.n64 13.653
R271 VPB.n64 VPB.n63 13.653
R272 VPB.n70 VPB.n69 13.653
R273 VPB.n69 VPB.n68 13.653
R274 VPB.n74 VPB.n73 13.653
R275 VPB.n73 VPB.n72 13.653
R276 VPB.n77 VPB.n76 13.653
R277 VPB.n76 VPB.n75 13.653
R278 VPB.n81 VPB.n80 13.653
R279 VPB.n80 VPB.n79 13.653
R280 VPB.n506 VPB.n0 13.653
R281 VPB VPB.n0 13.653
R282 VPB.n222 VPB.n221 13.35
R283 VPB.n305 VPB.n304 13.35
R284 VPB.n152 VPB.n151 13.35
R285 VPB.n382 VPB.n381 13.35
R286 VPB.n465 VPB.n464 13.35
R287 VPB.n63 VPB.n62 13.35
R288 VPB.n510 VPB.n509 13.276
R289 VPB.n509 VPB.n507 13.276
R290 VPB.n36 VPB.n18 13.276
R291 VPB.n18 VPB.n16 13.276
R292 VPB.n431 VPB.n413 13.276
R293 VPB.n413 VPB.n411 13.276
R294 VPB.n102 VPB.n84 13.276
R295 VPB.n84 VPB.n82 13.276
R296 VPB.n125 VPB.n107 13.276
R297 VPB.n107 VPB.n105 13.276
R298 VPB.n271 VPB.n253 13.276
R299 VPB.n253 VPB.n251 13.276
R300 VPB.n201 VPB.n197 13.276
R301 VPB.n276 VPB.n272 13.276
R302 VPB.n130 VPB.n126 13.276
R303 VPB.n133 VPB.n130 13.276
R304 VPB.n141 VPB.n137 13.276
R305 VPB.n145 VPB.n141 13.276
R306 VPB.n154 VPB.n150 13.276
R307 VPB.n163 VPB.n159 13.276
R308 VPB.n166 VPB.n163 13.276
R309 VPB.n348 VPB.n170 13.276
R310 VPB.n349 VPB.n348 13.276
R311 VPB.n353 VPB.n349 13.276
R312 VPB.n436 VPB.n432 13.276
R313 VPB.n41 VPB.n37 13.276
R314 VPB.n44 VPB.n41 13.276
R315 VPB.n52 VPB.n48 13.276
R316 VPB.n56 VPB.n52 13.276
R317 VPB.n65 VPB.n61 13.276
R318 VPB.n74 VPB.n70 13.276
R319 VPB.n77 VPB.n74 13.276
R320 VPB.n506 VPB.n81 13.276
R321 VPB.n191 VPB.n173 13.276
R322 VPB.n173 VPB.n171 13.276
R323 VPB.n178 VPB.n176 12.796
R324 VPB.n178 VPB.n177 12.564
R325 VPB.n170 VPB.n167 12.558
R326 VPB.n81 VPB.n78 12.558
R327 VPB.n205 VPB.n202 12.2
R328 VPB.n134 VPB.n133 12.2
R329 VPB.n45 VPB.n44 12.2
R330 VPB.n186 VPB.n185 12.198
R331 VPB.n184 VPB.n183 12.198
R332 VPB.n181 VPB.n180 12.198
R333 VPB.n150 VPB.n146 9.329
R334 VPB.n61 VPB.n57 9.329
R335 VPB.n155 VPB.n154 8.97
R336 VPB.n66 VPB.n65 8.97
R337 VPB.n191 VPB.n190 7.5
R338 VPB.n176 VPB.n175 7.5
R339 VPB.n180 VPB.n179 7.5
R340 VPB.n183 VPB.n182 7.5
R341 VPB.n173 VPB.n172 7.5
R342 VPB.n188 VPB.n174 7.5
R343 VPB.n253 VPB.n252 7.5
R344 VPB.n266 VPB.n265 7.5
R345 VPB.n260 VPB.n259 7.5
R346 VPB.n262 VPB.n261 7.5
R347 VPB.n255 VPB.n254 7.5
R348 VPB.n271 VPB.n270 7.5
R349 VPB.n107 VPB.n106 7.5
R350 VPB.n120 VPB.n119 7.5
R351 VPB.n114 VPB.n113 7.5
R352 VPB.n116 VPB.n115 7.5
R353 VPB.n109 VPB.n108 7.5
R354 VPB.n125 VPB.n124 7.5
R355 VPB.n84 VPB.n83 7.5
R356 VPB.n97 VPB.n96 7.5
R357 VPB.n91 VPB.n90 7.5
R358 VPB.n93 VPB.n92 7.5
R359 VPB.n86 VPB.n85 7.5
R360 VPB.n102 VPB.n101 7.5
R361 VPB.n413 VPB.n412 7.5
R362 VPB.n426 VPB.n425 7.5
R363 VPB.n420 VPB.n419 7.5
R364 VPB.n422 VPB.n421 7.5
R365 VPB.n415 VPB.n414 7.5
R366 VPB.n431 VPB.n430 7.5
R367 VPB.n18 VPB.n17 7.5
R368 VPB.n31 VPB.n30 7.5
R369 VPB.n25 VPB.n24 7.5
R370 VPB.n27 VPB.n26 7.5
R371 VPB.n20 VPB.n19 7.5
R372 VPB.n36 VPB.n35 7.5
R373 VPB.n509 VPB.n508 7.5
R374 VPB.n12 VPB.n11 7.5
R375 VPB.n6 VPB.n5 7.5
R376 VPB.n8 VPB.n7 7.5
R377 VPB.n2 VPB.n1 7.5
R378 VPB.n511 VPB.n510 7.5
R379 VPB.n37 VPB.n36 7.176
R380 VPB.n432 VPB.n431 7.176
R381 VPB.n349 VPB.n102 7.176
R382 VPB.n126 VPB.n125 7.176
R383 VPB.n272 VPB.n271 7.176
R384 VPB.n267 VPB.n264 6.729
R385 VPB.n263 VPB.n260 6.729
R386 VPB.n258 VPB.n255 6.729
R387 VPB.n121 VPB.n118 6.729
R388 VPB.n117 VPB.n114 6.729
R389 VPB.n112 VPB.n109 6.729
R390 VPB.n98 VPB.n95 6.729
R391 VPB.n94 VPB.n91 6.729
R392 VPB.n89 VPB.n86 6.729
R393 VPB.n427 VPB.n424 6.729
R394 VPB.n423 VPB.n420 6.729
R395 VPB.n418 VPB.n415 6.729
R396 VPB.n32 VPB.n29 6.729
R397 VPB.n28 VPB.n25 6.729
R398 VPB.n23 VPB.n20 6.729
R399 VPB.n13 VPB.n10 6.729
R400 VPB.n9 VPB.n6 6.729
R401 VPB.n4 VPB.n2 6.729
R402 VPB.n258 VPB.n257 6.728
R403 VPB.n263 VPB.n262 6.728
R404 VPB.n267 VPB.n266 6.728
R405 VPB.n270 VPB.n269 6.728
R406 VPB.n112 VPB.n111 6.728
R407 VPB.n117 VPB.n116 6.728
R408 VPB.n121 VPB.n120 6.728
R409 VPB.n124 VPB.n123 6.728
R410 VPB.n89 VPB.n88 6.728
R411 VPB.n94 VPB.n93 6.728
R412 VPB.n98 VPB.n97 6.728
R413 VPB.n101 VPB.n100 6.728
R414 VPB.n418 VPB.n417 6.728
R415 VPB.n423 VPB.n422 6.728
R416 VPB.n427 VPB.n426 6.728
R417 VPB.n430 VPB.n429 6.728
R418 VPB.n23 VPB.n22 6.728
R419 VPB.n28 VPB.n27 6.728
R420 VPB.n32 VPB.n31 6.728
R421 VPB.n35 VPB.n34 6.728
R422 VPB.n4 VPB.n3 6.728
R423 VPB.n9 VPB.n8 6.728
R424 VPB.n13 VPB.n12 6.728
R425 VPB.n512 VPB.n511 6.728
R426 VPB.n190 VPB.n189 6.398
R427 VPB.n206 VPB.n194 6.112
R428 VPB.n206 VPB.n205 6.101
R429 VPB.n231 VPB.n227 4.305
R430 VPB.n314 VPB.n310 4.305
R431 VPB.n159 VPB.n155 4.305
R432 VPB.n391 VPB.n387 4.305
R433 VPB.n474 VPB.n470 4.305
R434 VPB.n70 VPB.n66 4.305
R435 VPB.n214 VPB.n210 3.947
R436 VPB.n297 VPB.n293 3.947
R437 VPB.n146 VPB.n145 3.947
R438 VPB.n374 VPB.n370 3.947
R439 VPB.n457 VPB.n453 3.947
R440 VPB.n57 VPB.n56 3.947
R441 VPB.n188 VPB.n181 1.402
R442 VPB.n188 VPB.n184 1.402
R443 VPB.n188 VPB.n186 1.402
R444 VPB.n188 VPB.n187 1.402
R445 VPB.n202 VPB.n201 1.076
R446 VPB.n285 VPB.n282 1.076
R447 VPB.n137 VPB.n134 1.076
R448 VPB.n362 VPB.n359 1.076
R449 VPB.n445 VPB.n442 1.076
R450 VPB.n48 VPB.n45 1.076
R451 VPB.n189 VPB.n188 0.735
R452 VPB.n188 VPB.n178 0.735
R453 VPB.n241 VPB.n238 0.717
R454 VPB.n324 VPB.n321 0.717
R455 VPB.n167 VPB.n166 0.717
R456 VPB.n401 VPB.n398 0.717
R457 VPB.n484 VPB.n481 0.717
R458 VPB.n78 VPB.n77 0.717
R459 VPB.n268 VPB.n267 0.387
R460 VPB.n268 VPB.n263 0.387
R461 VPB.n268 VPB.n258 0.387
R462 VPB.n269 VPB.n268 0.387
R463 VPB.n122 VPB.n121 0.387
R464 VPB.n122 VPB.n117 0.387
R465 VPB.n122 VPB.n112 0.387
R466 VPB.n123 VPB.n122 0.387
R467 VPB.n99 VPB.n98 0.387
R468 VPB.n99 VPB.n94 0.387
R469 VPB.n99 VPB.n89 0.387
R470 VPB.n100 VPB.n99 0.387
R471 VPB.n428 VPB.n427 0.387
R472 VPB.n428 VPB.n423 0.387
R473 VPB.n428 VPB.n418 0.387
R474 VPB.n429 VPB.n428 0.387
R475 VPB.n33 VPB.n32 0.387
R476 VPB.n33 VPB.n28 0.387
R477 VPB.n33 VPB.n23 0.387
R478 VPB.n34 VPB.n33 0.387
R479 VPB.n513 VPB.n13 0.387
R480 VPB.n513 VPB.n9 0.387
R481 VPB.n513 VPB.n4 0.387
R482 VPB.n513 VPB.n512 0.387
R483 VPB.n277 VPB.n250 0.272
R484 VPB.n334 VPB.n333 0.272
R485 VPB.n437 VPB.n410 0.272
R486 VPB.n494 VPB.n493 0.272
R487 VPB.n505 VPB 0.198
R488 VPB.n208 VPB.n207 0.136
R489 VPB.n215 VPB.n208 0.136
R490 VPB.n220 VPB.n215 0.136
R491 VPB.n225 VPB.n220 0.136
R492 VPB.n232 VPB.n225 0.136
R493 VPB.n237 VPB.n232 0.136
R494 VPB.n242 VPB.n237 0.136
R495 VPB.n246 VPB.n242 0.136
R496 VPB.n250 VPB.n246 0.136
R497 VPB.n281 VPB.n277 0.136
R498 VPB.n286 VPB.n281 0.136
R499 VPB.n291 VPB.n286 0.136
R500 VPB.n298 VPB.n291 0.136
R501 VPB.n303 VPB.n298 0.136
R502 VPB.n308 VPB.n303 0.136
R503 VPB.n315 VPB.n308 0.136
R504 VPB.n320 VPB.n315 0.136
R505 VPB.n325 VPB.n320 0.136
R506 VPB.n329 VPB.n325 0.136
R507 VPB.n333 VPB.n329 0.136
R508 VPB.n335 VPB.n334 0.136
R509 VPB.n336 VPB.n335 0.136
R510 VPB.n337 VPB.n336 0.136
R511 VPB.n338 VPB.n337 0.136
R512 VPB.n339 VPB.n338 0.136
R513 VPB.n340 VPB.n339 0.136
R514 VPB.n341 VPB.n340 0.136
R515 VPB.n342 VPB.n341 0.136
R516 VPB.n343 VPB.n342 0.136
R517 VPB.n344 VPB.n343 0.136
R518 VPB.n345 VPB.n344 0.136
R519 VPB.n345 VPB 0.136
R520 VPB.n354 VPB 0.136
R521 VPB.n358 VPB.n354 0.136
R522 VPB.n363 VPB.n358 0.136
R523 VPB.n368 VPB.n363 0.136
R524 VPB.n375 VPB.n368 0.136
R525 VPB.n380 VPB.n375 0.136
R526 VPB.n385 VPB.n380 0.136
R527 VPB.n392 VPB.n385 0.136
R528 VPB.n397 VPB.n392 0.136
R529 VPB.n402 VPB.n397 0.136
R530 VPB.n406 VPB.n402 0.136
R531 VPB.n410 VPB.n406 0.136
R532 VPB.n441 VPB.n437 0.136
R533 VPB.n446 VPB.n441 0.136
R534 VPB.n451 VPB.n446 0.136
R535 VPB.n458 VPB.n451 0.136
R536 VPB.n463 VPB.n458 0.136
R537 VPB.n468 VPB.n463 0.136
R538 VPB.n475 VPB.n468 0.136
R539 VPB.n480 VPB.n475 0.136
R540 VPB.n485 VPB.n480 0.136
R541 VPB.n489 VPB.n485 0.136
R542 VPB.n493 VPB.n489 0.136
R543 VPB.n495 VPB.n494 0.136
R544 VPB.n496 VPB.n495 0.136
R545 VPB.n497 VPB.n496 0.136
R546 VPB.n498 VPB.n497 0.136
R547 VPB.n499 VPB.n498 0.136
R548 VPB.n500 VPB.n499 0.136
R549 VPB.n501 VPB.n500 0.136
R550 VPB.n502 VPB.n501 0.136
R551 VPB.n503 VPB.n502 0.136
R552 VPB.n504 VPB.n503 0.136
R553 VPB.n505 VPB.n504 0.136
R554 a_277_1004.n7 a_277_1004.t10 512.525
R555 a_277_1004.n5 a_277_1004.t7 512.525
R556 a_277_1004.n7 a_277_1004.t11 371.139
R557 a_277_1004.n5 a_277_1004.t12 371.139
R558 a_277_1004.n8 a_277_1004.t9 244.968
R559 a_277_1004.n6 a_277_1004.t8 244.968
R560 a_277_1004.n10 a_277_1004.n4 207.04
R561 a_277_1004.n8 a_277_1004.n7 198.954
R562 a_277_1004.n6 a_277_1004.n5 198.954
R563 a_277_1004.n12 a_277_1004.n10 176.926
R564 a_277_1004.n9 a_277_1004.n6 79.491
R565 a_277_1004.n3 a_277_1004.n2 79.232
R566 a_277_1004.n10 a_277_1004.n9 77.315
R567 a_277_1004.n9 a_277_1004.n8 76
R568 a_277_1004.n4 a_277_1004.n3 63.152
R569 a_277_1004.n4 a_277_1004.n0 16.08
R570 a_277_1004.n3 a_277_1004.n1 16.08
R571 a_277_1004.n12 a_277_1004.n11 15.218
R572 a_277_1004.n0 a_277_1004.t3 14.282
R573 a_277_1004.n0 a_277_1004.t2 14.282
R574 a_277_1004.n1 a_277_1004.t1 14.282
R575 a_277_1004.n1 a_277_1004.t0 14.282
R576 a_277_1004.n2 a_277_1004.t6 14.282
R577 a_277_1004.n2 a_277_1004.t5 14.282
R578 a_277_1004.n13 a_277_1004.n12 12.014
R579 a_599_943.n5 a_599_943.t12 512.525
R580 a_599_943.n7 a_599_943.t10 454.685
R581 a_599_943.n7 a_599_943.t8 428.979
R582 a_599_943.n5 a_599_943.t7 371.139
R583 a_599_943.n6 a_599_943.t9 297.715
R584 a_599_943.n8 a_599_943.t11 248.006
R585 a_599_943.n12 a_599_943.n10 229.673
R586 a_599_943.n10 a_599_943.n4 154.293
R587 a_599_943.n6 a_599_943.n5 146.207
R588 a_599_943.n9 a_599_943.n6 84.388
R589 a_599_943.n8 a_599_943.n7 81.941
R590 a_599_943.n9 a_599_943.n8 80.035
R591 a_599_943.n3 a_599_943.n2 79.232
R592 a_599_943.n10 a_599_943.n9 76
R593 a_599_943.n4 a_599_943.n3 63.152
R594 a_599_943.n4 a_599_943.n0 16.08
R595 a_599_943.n3 a_599_943.n1 16.08
R596 a_599_943.n12 a_599_943.n11 15.218
R597 a_599_943.n0 a_599_943.t2 14.282
R598 a_599_943.n0 a_599_943.t0 14.282
R599 a_599_943.n1 a_599_943.t3 14.282
R600 a_599_943.n1 a_599_943.t4 14.282
R601 a_599_943.n2 a_599_943.t6 14.282
R602 a_599_943.n2 a_599_943.t5 14.282
R603 a_599_943.n13 a_599_943.n12 12.014
R604 a_1561_943.n8 a_1561_943.t14 454.685
R605 a_1561_943.n10 a_1561_943.t8 454.685
R606 a_1561_943.n6 a_1561_943.t15 454.685
R607 a_1561_943.n8 a_1561_943.t11 428.979
R608 a_1561_943.n10 a_1561_943.t12 428.979
R609 a_1561_943.n6 a_1561_943.t13 428.979
R610 a_1561_943.n9 a_1561_943.t7 274.559
R611 a_1561_943.n7 a_1561_943.t10 274.559
R612 a_1561_943.n11 a_1561_943.t9 274.22
R613 a_1561_943.n16 a_1561_943.n14 249.704
R614 a_1561_943.n14 a_1561_943.n5 127.74
R615 a_1561_943.n13 a_1561_943.n7 82.484
R616 a_1561_943.n12 a_1561_943.n11 79.495
R617 a_1561_943.n4 a_1561_943.n3 79.232
R618 a_1561_943.n12 a_1561_943.n9 76
R619 a_1561_943.n14 a_1561_943.n13 76
R620 a_1561_943.n5 a_1561_943.n4 63.152
R621 a_1561_943.n9 a_1561_943.n8 55.388
R622 a_1561_943.n7 a_1561_943.n6 55.388
R623 a_1561_943.n11 a_1561_943.n10 55.049
R624 a_1561_943.n16 a_1561_943.n15 30
R625 a_1561_943.n17 a_1561_943.n0 24.383
R626 a_1561_943.n17 a_1561_943.n16 23.684
R627 a_1561_943.n5 a_1561_943.n1 16.08
R628 a_1561_943.n4 a_1561_943.n2 16.08
R629 a_1561_943.n1 a_1561_943.t1 14.282
R630 a_1561_943.n1 a_1561_943.t0 14.282
R631 a_1561_943.n2 a_1561_943.t4 14.282
R632 a_1561_943.n2 a_1561_943.t3 14.282
R633 a_1561_943.n3 a_1561_943.t5 14.282
R634 a_1561_943.n3 a_1561_943.t6 14.282
R635 a_1561_943.n13 a_1561_943.n12 4.035
R636 a_91_75.t0 a_91_75.n0 117.777
R637 a_91_75.n2 a_91_75.n1 55.228
R638 a_91_75.n4 a_91_75.n3 9.111
R639 a_91_75.n8 a_91_75.n6 7.859
R640 a_91_75.t0 a_91_75.n2 4.04
R641 a_91_75.t0 a_91_75.n8 3.034
R642 a_91_75.n6 a_91_75.n4 1.964
R643 a_91_75.n6 a_91_75.n5 1.964
R644 a_91_75.n8 a_91_75.n7 0.443
R645 a_372_182.n10 a_372_182.n8 82.852
R646 a_372_182.n11 a_372_182.n0 49.6
R647 a_372_182.n7 a_372_182.n6 32.833
R648 a_372_182.n8 a_372_182.t1 32.416
R649 a_372_182.n10 a_372_182.n9 27.2
R650 a_372_182.n3 a_372_182.n2 23.284
R651 a_372_182.n11 a_372_182.n10 22.4
R652 a_372_182.n7 a_372_182.n4 19.017
R653 a_372_182.n6 a_372_182.n5 13.494
R654 a_372_182.t1 a_372_182.n1 7.04
R655 a_372_182.t1 a_372_182.n3 5.727
R656 a_372_182.n8 a_372_182.n7 1.435
R657 a_2296_182.n12 a_2296_182.n10 82.852
R658 a_2296_182.t1 a_2296_182.n2 46.91
R659 a_2296_182.n7 a_2296_182.n5 34.805
R660 a_2296_182.n7 a_2296_182.n6 32.622
R661 a_2296_182.n10 a_2296_182.t1 32.416
R662 a_2296_182.n12 a_2296_182.n11 27.2
R663 a_2296_182.n13 a_2296_182.n0 23.498
R664 a_2296_182.n13 a_2296_182.n12 22.4
R665 a_2296_182.n9 a_2296_182.n7 19.017
R666 a_2296_182.n2 a_2296_182.n1 17.006
R667 a_2296_182.n5 a_2296_182.n4 7.5
R668 a_2296_182.n9 a_2296_182.n8 7.5
R669 a_2296_182.t1 a_2296_182.n3 7.04
R670 a_2296_182.n10 a_2296_182.n9 1.435
R671 a_2201_1004.n5 a_2201_1004.t9 512.525
R672 a_2201_1004.n5 a_2201_1004.t8 371.139
R673 a_2201_1004.n6 a_2201_1004.t7 244.609
R674 a_2201_1004.n7 a_2201_1004.n4 207.399
R675 a_2201_1004.n6 a_2201_1004.n5 199.313
R676 a_2201_1004.n9 a_2201_1004.n7 176.567
R677 a_2201_1004.n7 a_2201_1004.n6 153.315
R678 a_2201_1004.n3 a_2201_1004.n2 79.232
R679 a_2201_1004.n4 a_2201_1004.n3 63.152
R680 a_2201_1004.n4 a_2201_1004.n0 16.08
R681 a_2201_1004.n3 a_2201_1004.n1 16.08
R682 a_2201_1004.n9 a_2201_1004.n8 15.218
R683 a_2201_1004.n0 a_2201_1004.t4 14.282
R684 a_2201_1004.n0 a_2201_1004.t3 14.282
R685 a_2201_1004.n1 a_2201_1004.t1 14.282
R686 a_2201_1004.n1 a_2201_1004.t0 14.282
R687 a_2201_1004.n2 a_2201_1004.t6 14.282
R688 a_2201_1004.n2 a_2201_1004.t5 14.282
R689 a_2201_1004.n10 a_2201_1004.n9 12.014
R690 a_4220_182.n12 a_4220_182.n10 82.852
R691 a_4220_182.t1 a_4220_182.n2 46.91
R692 a_4220_182.n7 a_4220_182.n5 34.805
R693 a_4220_182.n7 a_4220_182.n6 32.622
R694 a_4220_182.n10 a_4220_182.t1 32.416
R695 a_4220_182.n12 a_4220_182.n11 27.2
R696 a_4220_182.n13 a_4220_182.n0 23.498
R697 a_4220_182.n13 a_4220_182.n12 22.4
R698 a_4220_182.n9 a_4220_182.n7 19.017
R699 a_4220_182.n2 a_4220_182.n1 17.006
R700 a_4220_182.n5 a_4220_182.n4 7.5
R701 a_4220_182.n9 a_4220_182.n8 7.5
R702 a_4220_182.t1 a_4220_182.n3 7.04
R703 a_4220_182.n10 a_4220_182.n9 1.435
R704 a_4125_1004.n5 a_4125_1004.t7 512.525
R705 a_4125_1004.n5 a_4125_1004.t9 371.139
R706 a_4125_1004.n6 a_4125_1004.t8 271.162
R707 a_4125_1004.n9 a_4125_1004.n7 203.12
R708 a_4125_1004.n7 a_4125_1004.n4 180.846
R709 a_4125_1004.n6 a_4125_1004.n5 172.76
R710 a_4125_1004.n7 a_4125_1004.n6 153.315
R711 a_4125_1004.n3 a_4125_1004.n2 79.232
R712 a_4125_1004.n4 a_4125_1004.n3 63.152
R713 a_4125_1004.n4 a_4125_1004.n0 16.08
R714 a_4125_1004.n3 a_4125_1004.n1 16.08
R715 a_4125_1004.n9 a_4125_1004.n8 15.218
R716 a_4125_1004.n0 a_4125_1004.t2 14.282
R717 a_4125_1004.n0 a_4125_1004.t3 14.282
R718 a_4125_1004.n1 a_4125_1004.t0 14.282
R719 a_4125_1004.n1 a_4125_1004.t1 14.282
R720 a_4125_1004.n2 a_4125_1004.t5 14.282
R721 a_4125_1004.n2 a_4125_1004.t6 14.282
R722 a_4125_1004.n10 a_4125_1004.n9 12.014
R723 a_1334_182.n9 a_1334_182.n7 82.852
R724 a_1334_182.n3 a_1334_182.n1 44.628
R725 a_1334_182.t0 a_1334_182.n9 32.417
R726 a_1334_182.n7 a_1334_182.n6 27.2
R727 a_1334_182.n5 a_1334_182.n4 23.498
R728 a_1334_182.n3 a_1334_182.n2 23.284
R729 a_1334_182.n7 a_1334_182.n5 22.4
R730 a_1334_182.t0 a_1334_182.n11 20.241
R731 a_1334_182.n11 a_1334_182.n10 13.494
R732 a_1334_182.t0 a_1334_182.n0 8.137
R733 a_1334_182.t0 a_1334_182.n3 5.727
R734 a_1334_182.n9 a_1334_182.n8 1.435
R735 a_2015_75.t0 a_2015_75.n0 117.777
R736 a_2015_75.n2 a_2015_75.n1 55.228
R737 a_2015_75.n4 a_2015_75.n3 9.111
R738 a_2015_75.t0 a_2015_75.n2 4.04
R739 a_2015_75.n8 a_2015_75.n7 2.455
R740 a_2015_75.n6 a_2015_75.n4 1.964
R741 a_2015_75.n6 a_2015_75.n5 1.964
R742 a_2015_75.n8 a_2015_75.n6 0.636
R743 a_2015_75.t0 a_2015_75.n8 0.246
R744 VNB VNB.n446 300.778
R745 VNB.n214 VNB.n213 199.897
R746 VNB.n87 VNB.n86 199.897
R747 VNB.n67 VNB.n66 199.897
R748 VNB.n356 VNB.n355 199.897
R749 VNB.n15 VNB.n14 199.897
R750 VNB.n96 VNB.n94 154.509
R751 VNB.n223 VNB.n221 154.509
R752 VNB.n365 VNB.n363 154.509
R753 VNB.n297 VNB.n295 154.509
R754 VNB.n24 VNB.n22 154.509
R755 VNB.n180 VNB.n179 147.75
R756 VNB.n255 VNB.n254 147.75
R757 VNB.n120 VNB.n119 147.75
R758 VNB.n397 VNB.n396 147.75
R759 VNB.n192 VNB.n189 121.366
R760 VNB.n267 VNB.n264 121.366
R761 VNB.n125 VNB.n123 121.366
R762 VNB.n409 VNB.n406 121.366
R763 VNB.n333 VNB.n332 85.559
R764 VNB.n53 VNB.n4 85.559
R765 VNB.n433 VNB.n432 76
R766 VNB.n420 VNB.n419 76
R767 VNB.n416 VNB.n415 76
R768 VNB.n412 VNB.n411 76
R769 VNB.n400 VNB.n399 76
R770 VNB.n395 VNB.n394 76
R771 VNB.n391 VNB.n390 76
R772 VNB.n387 VNB.n386 76
R773 VNB.n383 VNB.n382 76
R774 VNB.n379 VNB.n378 76
R775 VNB.n375 VNB.n374 76
R776 VNB.n371 VNB.n370 76
R777 VNB.n367 VNB.n366 76
R778 VNB.n345 VNB.n344 76
R779 VNB.n341 VNB.n340 76
R780 VNB.n337 VNB.n336 76
R781 VNB.n331 VNB.n330 76
R782 VNB.n327 VNB.n326 76
R783 VNB.n323 VNB.n322 76
R784 VNB.n319 VNB.n318 76
R785 VNB.n315 VNB.n314 76
R786 VNB.n311 VNB.n310 76
R787 VNB.n307 VNB.n306 76
R788 VNB.n303 VNB.n302 76
R789 VNB.n299 VNB.n298 76
R790 VNB.n293 VNB.n290 76
R791 VNB.n278 VNB.n277 76
R792 VNB.n274 VNB.n273 76
R793 VNB.n270 VNB.n269 76
R794 VNB.n258 VNB.n257 76
R795 VNB.n253 VNB.n252 76
R796 VNB.n249 VNB.n248 76
R797 VNB.n245 VNB.n244 76
R798 VNB.n241 VNB.n240 76
R799 VNB.n237 VNB.n236 76
R800 VNB.n233 VNB.n232 76
R801 VNB.n229 VNB.n228 76
R802 VNB.n225 VNB.n224 76
R803 VNB.n203 VNB.n202 76
R804 VNB.n199 VNB.n198 76
R805 VNB.n195 VNB.n194 76
R806 VNB.n183 VNB.n182 76
R807 VNB.n178 VNB.n177 76
R808 VNB.n174 VNB.n173 76
R809 VNB.n170 VNB.n169 76
R810 VNB.n166 VNB.n165 76
R811 VNB.n130 VNB.n129 73.875
R812 VNB.n188 VNB.n187 64.552
R813 VNB.n263 VNB.n262 64.552
R814 VNB.n128 VNB.n76 64.552
R815 VNB.n405 VNB.n404 64.552
R816 VNB.n335 VNB.n334 41.971
R817 VNB.n51 VNB.n50 41.971
R818 VNB.n192 VNB.n191 36.937
R819 VNB.n267 VNB.n266 36.937
R820 VNB.n125 VNB.n124 36.937
R821 VNB.n409 VNB.n408 36.937
R822 VNB.n161 VNB.n160 35.118
R823 VNB.n191 VNB.n190 29.844
R824 VNB.n266 VNB.n265 29.844
R825 VNB.n408 VNB.n407 29.844
R826 VNB.n187 VNB.n186 28.421
R827 VNB.n262 VNB.n261 28.421
R828 VNB.n76 VNB.n75 28.421
R829 VNB.n404 VNB.n403 28.421
R830 VNB.n187 VNB.n185 25.263
R831 VNB.n262 VNB.n260 25.263
R832 VNB.n76 VNB.n74 25.263
R833 VNB.n404 VNB.n402 25.263
R834 VNB.n185 VNB.n184 24.383
R835 VNB.n260 VNB.n259 24.383
R836 VNB.n74 VNB.n73 24.383
R837 VNB.n402 VNB.n401 24.383
R838 VNB.n150 VNB.n147 20.452
R839 VNB.n434 VNB.n433 20.452
R840 VNB.n159 VNB.n158 13.653
R841 VNB.n158 VNB.n157 13.653
R842 VNB.n156 VNB.n155 13.653
R843 VNB.n155 VNB.n154 13.653
R844 VNB.n153 VNB.n152 13.653
R845 VNB.n152 VNB.n151 13.653
R846 VNB.n165 VNB.n164 13.653
R847 VNB.n164 VNB.n163 13.653
R848 VNB.n169 VNB.n168 13.653
R849 VNB.n168 VNB.n167 13.653
R850 VNB.n173 VNB.n172 13.653
R851 VNB.n172 VNB.n171 13.653
R852 VNB.n177 VNB.n176 13.653
R853 VNB.n176 VNB.n175 13.653
R854 VNB.n182 VNB.n181 13.653
R855 VNB.n181 VNB.n180 13.653
R856 VNB.n194 VNB.n193 13.653
R857 VNB.n193 VNB.n192 13.653
R858 VNB.n198 VNB.n197 13.653
R859 VNB.n197 VNB.n196 13.653
R860 VNB.n202 VNB.n201 13.653
R861 VNB.n201 VNB.n200 13.653
R862 VNB.n224 VNB.n223 13.653
R863 VNB.n223 VNB.n222 13.653
R864 VNB.n228 VNB.n227 13.653
R865 VNB.n227 VNB.n226 13.653
R866 VNB.n232 VNB.n231 13.653
R867 VNB.n231 VNB.n230 13.653
R868 VNB.n236 VNB.n235 13.653
R869 VNB.n235 VNB.n234 13.653
R870 VNB.n240 VNB.n239 13.653
R871 VNB.n239 VNB.n238 13.653
R872 VNB.n244 VNB.n243 13.653
R873 VNB.n243 VNB.n242 13.653
R874 VNB.n248 VNB.n247 13.653
R875 VNB.n247 VNB.n246 13.653
R876 VNB.n252 VNB.n251 13.653
R877 VNB.n251 VNB.n250 13.653
R878 VNB.n257 VNB.n256 13.653
R879 VNB.n256 VNB.n255 13.653
R880 VNB.n269 VNB.n268 13.653
R881 VNB.n268 VNB.n267 13.653
R882 VNB.n273 VNB.n272 13.653
R883 VNB.n272 VNB.n271 13.653
R884 VNB.n277 VNB.n276 13.653
R885 VNB.n276 VNB.n275 13.653
R886 VNB.n97 VNB.n96 13.653
R887 VNB.n96 VNB.n95 13.653
R888 VNB.n100 VNB.n99 13.653
R889 VNB.n99 VNB.n98 13.653
R890 VNB.n103 VNB.n102 13.653
R891 VNB.n102 VNB.n101 13.653
R892 VNB.n106 VNB.n105 13.653
R893 VNB.n105 VNB.n104 13.653
R894 VNB.n109 VNB.n108 13.653
R895 VNB.n108 VNB.n107 13.653
R896 VNB.n112 VNB.n111 13.653
R897 VNB.n111 VNB.n110 13.653
R898 VNB.n115 VNB.n114 13.653
R899 VNB.n114 VNB.n113 13.653
R900 VNB.n118 VNB.n117 13.653
R901 VNB.n117 VNB.n116 13.653
R902 VNB.n122 VNB.n121 13.653
R903 VNB.n121 VNB.n120 13.653
R904 VNB.n127 VNB.n126 13.653
R905 VNB.n126 VNB.n125 13.653
R906 VNB.n132 VNB.n131 13.653
R907 VNB.n131 VNB.n130 13.653
R908 VNB.n293 VNB.n292 13.653
R909 VNB.n292 VNB.n291 13.653
R910 VNB.n298 VNB.n297 13.653
R911 VNB.n297 VNB.n296 13.653
R912 VNB.n302 VNB.n301 13.653
R913 VNB.n301 VNB.n300 13.653
R914 VNB.n306 VNB.n305 13.653
R915 VNB.n305 VNB.n304 13.653
R916 VNB.n310 VNB.n309 13.653
R917 VNB.n309 VNB.n308 13.653
R918 VNB.n314 VNB.n313 13.653
R919 VNB.n313 VNB.n312 13.653
R920 VNB.n318 VNB.n317 13.653
R921 VNB.n317 VNB.n316 13.653
R922 VNB.n322 VNB.n321 13.653
R923 VNB.n321 VNB.n320 13.653
R924 VNB.n326 VNB.n325 13.653
R925 VNB.n325 VNB.n324 13.653
R926 VNB.n330 VNB.n329 13.653
R927 VNB.n329 VNB.n328 13.653
R928 VNB.n336 VNB.n335 13.653
R929 VNB.n340 VNB.n339 13.653
R930 VNB.n339 VNB.n338 13.653
R931 VNB.n344 VNB.n343 13.653
R932 VNB.n343 VNB.n342 13.653
R933 VNB.n366 VNB.n365 13.653
R934 VNB.n365 VNB.n364 13.653
R935 VNB.n370 VNB.n369 13.653
R936 VNB.n369 VNB.n368 13.653
R937 VNB.n374 VNB.n373 13.653
R938 VNB.n373 VNB.n372 13.653
R939 VNB.n378 VNB.n377 13.653
R940 VNB.n377 VNB.n376 13.653
R941 VNB.n382 VNB.n381 13.653
R942 VNB.n381 VNB.n380 13.653
R943 VNB.n386 VNB.n385 13.653
R944 VNB.n385 VNB.n384 13.653
R945 VNB.n390 VNB.n389 13.653
R946 VNB.n389 VNB.n388 13.653
R947 VNB.n394 VNB.n393 13.653
R948 VNB.n393 VNB.n392 13.653
R949 VNB.n399 VNB.n398 13.653
R950 VNB.n398 VNB.n397 13.653
R951 VNB.n411 VNB.n410 13.653
R952 VNB.n410 VNB.n409 13.653
R953 VNB.n415 VNB.n414 13.653
R954 VNB.n414 VNB.n413 13.653
R955 VNB.n419 VNB.n418 13.653
R956 VNB.n418 VNB.n417 13.653
R957 VNB.n25 VNB.n24 13.653
R958 VNB.n24 VNB.n23 13.653
R959 VNB.n28 VNB.n27 13.653
R960 VNB.n27 VNB.n26 13.653
R961 VNB.n31 VNB.n30 13.653
R962 VNB.n30 VNB.n29 13.653
R963 VNB.n34 VNB.n33 13.653
R964 VNB.n33 VNB.n32 13.653
R965 VNB.n37 VNB.n36 13.653
R966 VNB.n36 VNB.n35 13.653
R967 VNB.n40 VNB.n39 13.653
R968 VNB.n39 VNB.n38 13.653
R969 VNB.n43 VNB.n42 13.653
R970 VNB.n42 VNB.n41 13.653
R971 VNB.n46 VNB.n45 13.653
R972 VNB.n45 VNB.n44 13.653
R973 VNB.n49 VNB.n48 13.653
R974 VNB.n48 VNB.n47 13.653
R975 VNB.n52 VNB.n51 13.653
R976 VNB.n56 VNB.n55 13.653
R977 VNB.n55 VNB.n54 13.653
R978 VNB.n433 VNB.n0 13.653
R979 VNB VNB.n0 13.653
R980 VNB.n150 VNB.n149 13.653
R981 VNB.n149 VNB.n148 13.653
R982 VNB.n441 VNB.n438 13.577
R983 VNB.n135 VNB.n133 13.276
R984 VNB.n147 VNB.n135 13.276
R985 VNB.n206 VNB.n204 13.276
R986 VNB.n219 VNB.n206 13.276
R987 VNB.n79 VNB.n77 13.276
R988 VNB.n92 VNB.n79 13.276
R989 VNB.n59 VNB.n57 13.276
R990 VNB.n72 VNB.n59 13.276
R991 VNB.n348 VNB.n346 13.276
R992 VNB.n361 VNB.n348 13.276
R993 VNB.n7 VNB.n5 13.276
R994 VNB.n20 VNB.n7 13.276
R995 VNB.n159 VNB.n156 13.276
R996 VNB.n156 VNB.n153 13.276
R997 VNB.n224 VNB.n220 13.276
R998 VNB.n97 VNB.n93 13.276
R999 VNB.n100 VNB.n97 13.276
R1000 VNB.n103 VNB.n100 13.276
R1001 VNB.n106 VNB.n103 13.276
R1002 VNB.n109 VNB.n106 13.276
R1003 VNB.n112 VNB.n109 13.276
R1004 VNB.n115 VNB.n112 13.276
R1005 VNB.n118 VNB.n115 13.276
R1006 VNB.n122 VNB.n118 13.276
R1007 VNB.n127 VNB.n122 13.276
R1008 VNB.n293 VNB.n132 13.276
R1009 VNB.n294 VNB.n293 13.276
R1010 VNB.n298 VNB.n294 13.276
R1011 VNB.n366 VNB.n362 13.276
R1012 VNB.n25 VNB.n21 13.276
R1013 VNB.n28 VNB.n25 13.276
R1014 VNB.n31 VNB.n28 13.276
R1015 VNB.n34 VNB.n31 13.276
R1016 VNB.n37 VNB.n34 13.276
R1017 VNB.n40 VNB.n37 13.276
R1018 VNB.n43 VNB.n40 13.276
R1019 VNB.n46 VNB.n43 13.276
R1020 VNB.n49 VNB.n46 13.276
R1021 VNB.n52 VNB.n49 13.276
R1022 VNB.n433 VNB.n56 13.276
R1023 VNB.n3 VNB.n1 13.276
R1024 VNB.n434 VNB.n3 13.276
R1025 VNB.n132 VNB.n128 12.02
R1026 VNB.n56 VNB.n53 12.02
R1027 VNB.n443 VNB.n442 7.5
R1028 VNB.n212 VNB.n211 7.5
R1029 VNB.n208 VNB.n207 7.5
R1030 VNB.n206 VNB.n205 7.5
R1031 VNB.n219 VNB.n218 7.5
R1032 VNB.n85 VNB.n84 7.5
R1033 VNB.n81 VNB.n80 7.5
R1034 VNB.n79 VNB.n78 7.5
R1035 VNB.n92 VNB.n91 7.5
R1036 VNB.n65 VNB.n64 7.5
R1037 VNB.n61 VNB.n60 7.5
R1038 VNB.n59 VNB.n58 7.5
R1039 VNB.n72 VNB.n71 7.5
R1040 VNB.n354 VNB.n353 7.5
R1041 VNB.n350 VNB.n349 7.5
R1042 VNB.n348 VNB.n347 7.5
R1043 VNB.n361 VNB.n360 7.5
R1044 VNB.n13 VNB.n12 7.5
R1045 VNB.n9 VNB.n8 7.5
R1046 VNB.n7 VNB.n6 7.5
R1047 VNB.n20 VNB.n19 7.5
R1048 VNB.n435 VNB.n434 7.5
R1049 VNB.n3 VNB.n2 7.5
R1050 VNB.n440 VNB.n439 7.5
R1051 VNB.n141 VNB.n140 7.5
R1052 VNB.n137 VNB.n136 7.5
R1053 VNB.n135 VNB.n134 7.5
R1054 VNB.n147 VNB.n146 7.5
R1055 VNB.n220 VNB.n219 7.176
R1056 VNB.n93 VNB.n92 7.176
R1057 VNB.n294 VNB.n72 7.176
R1058 VNB.n362 VNB.n361 7.176
R1059 VNB.n21 VNB.n20 7.176
R1060 VNB.n445 VNB.n443 7.011
R1061 VNB.n215 VNB.n212 7.011
R1062 VNB.n210 VNB.n208 7.011
R1063 VNB.n88 VNB.n85 7.011
R1064 VNB.n83 VNB.n81 7.011
R1065 VNB.n68 VNB.n65 7.011
R1066 VNB.n63 VNB.n61 7.011
R1067 VNB.n357 VNB.n354 7.011
R1068 VNB.n352 VNB.n350 7.011
R1069 VNB.n16 VNB.n13 7.011
R1070 VNB.n11 VNB.n9 7.011
R1071 VNB.n143 VNB.n141 7.011
R1072 VNB.n139 VNB.n137 7.011
R1073 VNB.n218 VNB.n217 7.01
R1074 VNB.n210 VNB.n209 7.01
R1075 VNB.n215 VNB.n214 7.01
R1076 VNB.n91 VNB.n90 7.01
R1077 VNB.n83 VNB.n82 7.01
R1078 VNB.n88 VNB.n87 7.01
R1079 VNB.n71 VNB.n70 7.01
R1080 VNB.n63 VNB.n62 7.01
R1081 VNB.n68 VNB.n67 7.01
R1082 VNB.n360 VNB.n359 7.01
R1083 VNB.n352 VNB.n351 7.01
R1084 VNB.n357 VNB.n356 7.01
R1085 VNB.n19 VNB.n18 7.01
R1086 VNB.n11 VNB.n10 7.01
R1087 VNB.n16 VNB.n15 7.01
R1088 VNB.n146 VNB.n145 7.01
R1089 VNB.n139 VNB.n138 7.01
R1090 VNB.n143 VNB.n142 7.01
R1091 VNB.n445 VNB.n444 7.01
R1092 VNB.n441 VNB.n440 6.788
R1093 VNB.n436 VNB.n435 6.788
R1094 VNB.n160 VNB.n150 6.111
R1095 VNB.n160 VNB.n159 6.1
R1096 VNB.n194 VNB.n188 1.255
R1097 VNB.n269 VNB.n263 1.255
R1098 VNB.n128 VNB.n127 1.255
R1099 VNB.n336 VNB.n333 1.255
R1100 VNB.n411 VNB.n405 1.255
R1101 VNB.n53 VNB.n52 1.255
R1102 VNB.n446 VNB.n437 0.921
R1103 VNB.n446 VNB.n441 0.476
R1104 VNB.n446 VNB.n436 0.475
R1105 VNB.n225 VNB.n203 0.272
R1106 VNB.n279 VNB.n278 0.272
R1107 VNB.n367 VNB.n345 0.272
R1108 VNB.n421 VNB.n420 0.272
R1109 VNB.n216 VNB.n210 0.246
R1110 VNB.n217 VNB.n216 0.246
R1111 VNB.n216 VNB.n215 0.246
R1112 VNB.n89 VNB.n83 0.246
R1113 VNB.n90 VNB.n89 0.246
R1114 VNB.n89 VNB.n88 0.246
R1115 VNB.n69 VNB.n63 0.246
R1116 VNB.n70 VNB.n69 0.246
R1117 VNB.n69 VNB.n68 0.246
R1118 VNB.n358 VNB.n352 0.246
R1119 VNB.n359 VNB.n358 0.246
R1120 VNB.n358 VNB.n357 0.246
R1121 VNB.n17 VNB.n11 0.246
R1122 VNB.n18 VNB.n17 0.246
R1123 VNB.n17 VNB.n16 0.246
R1124 VNB.n144 VNB.n139 0.246
R1125 VNB.n145 VNB.n144 0.246
R1126 VNB.n144 VNB.n143 0.246
R1127 VNB.n446 VNB.n445 0.246
R1128 VNB.n432 VNB 0.198
R1129 VNB.n162 VNB.n161 0.136
R1130 VNB.n166 VNB.n162 0.136
R1131 VNB.n170 VNB.n166 0.136
R1132 VNB.n174 VNB.n170 0.136
R1133 VNB.n178 VNB.n174 0.136
R1134 VNB.n183 VNB.n178 0.136
R1135 VNB.n195 VNB.n183 0.136
R1136 VNB.n199 VNB.n195 0.136
R1137 VNB.n203 VNB.n199 0.136
R1138 VNB.n229 VNB.n225 0.136
R1139 VNB.n233 VNB.n229 0.136
R1140 VNB.n237 VNB.n233 0.136
R1141 VNB.n241 VNB.n237 0.136
R1142 VNB.n245 VNB.n241 0.136
R1143 VNB.n249 VNB.n245 0.136
R1144 VNB.n253 VNB.n249 0.136
R1145 VNB.n258 VNB.n253 0.136
R1146 VNB.n270 VNB.n258 0.136
R1147 VNB.n274 VNB.n270 0.136
R1148 VNB.n278 VNB.n274 0.136
R1149 VNB.n280 VNB.n279 0.136
R1150 VNB.n281 VNB.n280 0.136
R1151 VNB.n282 VNB.n281 0.136
R1152 VNB.n283 VNB.n282 0.136
R1153 VNB.n284 VNB.n283 0.136
R1154 VNB.n285 VNB.n284 0.136
R1155 VNB.n286 VNB.n285 0.136
R1156 VNB.n287 VNB.n286 0.136
R1157 VNB.n288 VNB.n287 0.136
R1158 VNB.n289 VNB.n288 0.136
R1159 VNB.n290 VNB.n289 0.136
R1160 VNB.n290 VNB 0.136
R1161 VNB.n299 VNB 0.136
R1162 VNB.n303 VNB.n299 0.136
R1163 VNB.n307 VNB.n303 0.136
R1164 VNB.n311 VNB.n307 0.136
R1165 VNB.n315 VNB.n311 0.136
R1166 VNB.n319 VNB.n315 0.136
R1167 VNB.n323 VNB.n319 0.136
R1168 VNB.n327 VNB.n323 0.136
R1169 VNB.n331 VNB.n327 0.136
R1170 VNB.n337 VNB.n331 0.136
R1171 VNB.n341 VNB.n337 0.136
R1172 VNB.n345 VNB.n341 0.136
R1173 VNB.n371 VNB.n367 0.136
R1174 VNB.n375 VNB.n371 0.136
R1175 VNB.n379 VNB.n375 0.136
R1176 VNB.n383 VNB.n379 0.136
R1177 VNB.n387 VNB.n383 0.136
R1178 VNB.n391 VNB.n387 0.136
R1179 VNB.n395 VNB.n391 0.136
R1180 VNB.n400 VNB.n395 0.136
R1181 VNB.n412 VNB.n400 0.136
R1182 VNB.n416 VNB.n412 0.136
R1183 VNB.n420 VNB.n416 0.136
R1184 VNB.n422 VNB.n421 0.136
R1185 VNB.n423 VNB.n422 0.136
R1186 VNB.n424 VNB.n423 0.136
R1187 VNB.n425 VNB.n424 0.136
R1188 VNB.n426 VNB.n425 0.136
R1189 VNB.n427 VNB.n426 0.136
R1190 VNB.n428 VNB.n427 0.136
R1191 VNB.n429 VNB.n428 0.136
R1192 VNB.n430 VNB.n429 0.136
R1193 VNB.n431 VNB.n430 0.136
R1194 VNB.n432 VNB.n431 0.136
R1195 a_3258_182.n9 a_3258_182.n7 82.852
R1196 a_3258_182.n3 a_3258_182.n1 44.628
R1197 a_3258_182.t0 a_3258_182.n9 32.417
R1198 a_3258_182.n7 a_3258_182.n6 27.2
R1199 a_3258_182.n5 a_3258_182.n4 23.498
R1200 a_3258_182.n3 a_3258_182.n2 23.284
R1201 a_3258_182.n7 a_3258_182.n5 22.4
R1202 a_3258_182.t0 a_3258_182.n11 20.241
R1203 a_3258_182.n11 a_3258_182.n10 13.494
R1204 a_3258_182.t0 a_3258_182.n0 8.137
R1205 a_3258_182.t0 a_3258_182.n3 5.727
R1206 a_3258_182.n9 a_3258_182.n8 1.435
R1207 a_5182_182.n10 a_5182_182.n8 82.852
R1208 a_5182_182.n7 a_5182_182.n6 32.833
R1209 a_5182_182.n8 a_5182_182.t1 32.416
R1210 a_5182_182.n10 a_5182_182.n9 27.2
R1211 a_5182_182.n11 a_5182_182.n0 23.498
R1212 a_5182_182.n3 a_5182_182.n2 23.284
R1213 a_5182_182.n11 a_5182_182.n10 22.4
R1214 a_5182_182.n7 a_5182_182.n4 19.017
R1215 a_5182_182.n6 a_5182_182.n5 13.494
R1216 a_5182_182.t1 a_5182_182.n1 7.04
R1217 a_5182_182.t1 a_5182_182.n3 5.727
R1218 a_5182_182.n8 a_5182_182.n7 1.435
R1219 a_2977_75.n5 a_2977_75.n4 19.724
R1220 a_2977_75.t0 a_2977_75.n3 11.595
R1221 a_2977_75.t0 a_2977_75.n5 9.207
R1222 a_2977_75.n2 a_2977_75.n1 2.455
R1223 a_2977_75.n2 a_2977_75.n0 1.32
R1224 a_2977_75.t0 a_2977_75.n2 0.246
R1225 a_1053_75.n1 a_1053_75.n0 25.576
R1226 a_1053_75.n3 a_1053_75.n2 9.111
R1227 a_1053_75.n7 a_1053_75.n6 2.455
R1228 a_1053_75.n5 a_1053_75.n3 1.964
R1229 a_1053_75.n5 a_1053_75.n4 1.964
R1230 a_1053_75.t0 a_1053_75.n1 1.871
R1231 a_1053_75.n7 a_1053_75.n5 0.636
R1232 a_1053_75.t0 a_1053_75.n7 0.246
R1233 a_3939_75.n1 a_3939_75.n0 25.576
R1234 a_3939_75.n3 a_3939_75.n2 9.111
R1235 a_3939_75.n7 a_3939_75.n6 2.455
R1236 a_3939_75.n5 a_3939_75.n3 1.964
R1237 a_3939_75.n5 a_3939_75.n4 1.964
R1238 a_3939_75.t0 a_3939_75.n1 1.871
R1239 a_3939_75.n7 a_3939_75.n5 0.636
R1240 a_3939_75.t0 a_3939_75.n7 0.246
R1241 a_4901_75.n5 a_4901_75.n4 19.724
R1242 a_4901_75.t0 a_4901_75.n3 11.595
R1243 a_4901_75.t0 a_4901_75.n5 9.207
R1244 a_4901_75.n2 a_4901_75.n1 2.455
R1245 a_4901_75.n2 a_4901_75.n0 1.32
R1246 a_4901_75.t0 a_4901_75.n2 0.246
C11 VPB VNB 21.96fF
C12 a_4901_75.n0 VNB 0.10fF
C13 a_4901_75.n1 VNB 0.04fF
C14 a_4901_75.n2 VNB 0.03fF
C15 a_4901_75.n3 VNB 0.07fF
C16 a_4901_75.n4 VNB 0.08fF
C17 a_4901_75.n5 VNB 0.06fF
C18 a_3939_75.n0 VNB 0.09fF
C19 a_3939_75.n1 VNB 0.10fF
C20 a_3939_75.n2 VNB 0.05fF
C21 a_3939_75.n3 VNB 0.03fF
C22 a_3939_75.n4 VNB 0.04fF
C23 a_3939_75.n5 VNB 0.03fF
C24 a_3939_75.n6 VNB 0.04fF
C25 a_1053_75.n0 VNB 0.09fF
C26 a_1053_75.n1 VNB 0.10fF
C27 a_1053_75.n2 VNB 0.05fF
C28 a_1053_75.n3 VNB 0.03fF
C29 a_1053_75.n4 VNB 0.04fF
C30 a_1053_75.n5 VNB 0.03fF
C31 a_1053_75.n6 VNB 0.04fF
C32 a_2977_75.n0 VNB 0.10fF
C33 a_2977_75.n1 VNB 0.04fF
C34 a_2977_75.n2 VNB 0.03fF
C35 a_2977_75.n3 VNB 0.07fF
C36 a_2977_75.n4 VNB 0.08fF
C37 a_2977_75.n5 VNB 0.06fF
C38 a_5182_182.n0 VNB 0.02fF
C39 a_5182_182.n1 VNB 0.09fF
C40 a_5182_182.n2 VNB 0.13fF
C41 a_5182_182.n3 VNB 0.11fF
C42 a_5182_182.n4 VNB 0.09fF
C43 a_5182_182.n5 VNB 0.05fF
C44 a_5182_182.n6 VNB 0.01fF
C45 a_5182_182.n7 VNB 0.03fF
C46 a_5182_182.n8 VNB 0.11fF
C47 a_5182_182.n9 VNB 0.02fF
C48 a_5182_182.n10 VNB 0.05fF
C49 a_5182_182.n11 VNB 0.03fF
C50 a_3258_182.n0 VNB 0.07fF
C51 a_3258_182.n1 VNB 0.09fF
C52 a_3258_182.n2 VNB 0.13fF
C53 a_3258_182.n3 VNB 0.11fF
C54 a_3258_182.n4 VNB 0.02fF
C55 a_3258_182.n5 VNB 0.03fF
C56 a_3258_182.n6 VNB 0.02fF
C57 a_3258_182.n7 VNB 0.05fF
C58 a_3258_182.n8 VNB 0.03fF
C59 a_3258_182.n9 VNB 0.11fF
C60 a_3258_182.n10 VNB 0.06fF
C61 a_3258_182.n11 VNB 0.01fF
C62 a_3258_182.t0 VNB 0.33fF
C63 a_2015_75.n0 VNB 0.03fF
C64 a_2015_75.n1 VNB 0.10fF
C65 a_2015_75.n2 VNB 0.10fF
C66 a_2015_75.n3 VNB 0.05fF
C67 a_2015_75.n4 VNB 0.03fF
C68 a_2015_75.n5 VNB 0.04fF
C69 a_2015_75.n6 VNB 0.03fF
C70 a_2015_75.n7 VNB 0.04fF
C71 a_1334_182.n0 VNB 0.07fF
C72 a_1334_182.n1 VNB 0.09fF
C73 a_1334_182.n2 VNB 0.13fF
C74 a_1334_182.n3 VNB 0.11fF
C75 a_1334_182.n4 VNB 0.02fF
C76 a_1334_182.n5 VNB 0.03fF
C77 a_1334_182.n6 VNB 0.02fF
C78 a_1334_182.n7 VNB 0.05fF
C79 a_1334_182.n8 VNB 0.03fF
C80 a_1334_182.n9 VNB 0.11fF
C81 a_1334_182.n10 VNB 0.06fF
C82 a_1334_182.n11 VNB 0.01fF
C83 a_1334_182.t0 VNB 0.33fF
C84 a_4125_1004.n0 VNB 0.47fF
C85 a_4125_1004.n1 VNB 0.47fF
C86 a_4125_1004.n2 VNB 0.55fF
C87 a_4125_1004.n3 VNB 0.17fF
C88 a_4125_1004.n4 VNB 0.28fF
C89 a_4125_1004.n5 VNB 0.31fF
C90 a_4125_1004.n6 VNB 0.56fF
C91 a_4125_1004.n7 VNB 0.55fF
C92 a_4125_1004.n8 VNB 0.07fF
C93 a_4125_1004.n9 VNB 0.24fF
C94 a_4125_1004.n10 VNB 0.04fF
C95 a_4220_182.n0 VNB 0.02fF
C96 a_4220_182.n1 VNB 0.07fF
C97 a_4220_182.n2 VNB 0.13fF
C98 a_4220_182.n3 VNB 0.09fF
C99 a_4220_182.t1 VNB 0.25fF
C100 a_4220_182.n4 VNB 0.05fF
C101 a_4220_182.n5 VNB 0.06fF
C102 a_4220_182.n6 VNB 0.07fF
C103 a_4220_182.n7 VNB 0.07fF
C104 a_4220_182.n8 VNB 0.03fF
C105 a_4220_182.n9 VNB 0.01fF
C106 a_4220_182.n10 VNB 0.11fF
C107 a_4220_182.n11 VNB 0.02fF
C108 a_4220_182.n12 VNB 0.05fF
C109 a_4220_182.n13 VNB 0.03fF
C110 a_2201_1004.n0 VNB 0.53fF
C111 a_2201_1004.n1 VNB 0.53fF
C112 a_2201_1004.n2 VNB 0.62fF
C113 a_2201_1004.n3 VNB 0.20fF
C114 a_2201_1004.n4 VNB 0.34fF
C115 a_2201_1004.n5 VNB 0.37fF
C116 a_2201_1004.n6 VNB 0.63fF
C117 a_2201_1004.n7 VNB 0.62fF
C118 a_2201_1004.n8 VNB 0.08fF
C119 a_2201_1004.n9 VNB 0.24fF
C120 a_2201_1004.n10 VNB 0.04fF
C121 a_2296_182.n0 VNB 0.02fF
C122 a_2296_182.n1 VNB 0.07fF
C123 a_2296_182.n2 VNB 0.13fF
C124 a_2296_182.n3 VNB 0.09fF
C125 a_2296_182.t1 VNB 0.25fF
C126 a_2296_182.n4 VNB 0.05fF
C127 a_2296_182.n5 VNB 0.06fF
C128 a_2296_182.n6 VNB 0.07fF
C129 a_2296_182.n7 VNB 0.07fF
C130 a_2296_182.n8 VNB 0.03fF
C131 a_2296_182.n9 VNB 0.01fF
C132 a_2296_182.n10 VNB 0.11fF
C133 a_2296_182.n11 VNB 0.02fF
C134 a_2296_182.n12 VNB 0.05fF
C135 a_2296_182.n13 VNB 0.03fF
C136 a_372_182.n0 VNB 0.02fF
C137 a_372_182.n1 VNB 0.09fF
C138 a_372_182.n2 VNB 0.13fF
C139 a_372_182.n3 VNB 0.11fF
C140 a_372_182.t1 VNB 0.30fF
C141 a_372_182.n4 VNB 0.09fF
C142 a_372_182.n5 VNB 0.06fF
C143 a_372_182.n6 VNB 0.01fF
C144 a_372_182.n7 VNB 0.03fF
C145 a_372_182.n8 VNB 0.11fF
C146 a_372_182.n9 VNB 0.02fF
C147 a_372_182.n10 VNB 0.05fF
C148 a_372_182.n11 VNB 0.02fF
C149 a_91_75.n0 VNB 0.03fF
C150 a_91_75.n1 VNB 0.10fF
C151 a_91_75.n2 VNB 0.10fF
C152 a_91_75.n3 VNB 0.04fF
C153 a_91_75.n4 VNB 0.03fF
C154 a_91_75.n5 VNB 0.03fF
C155 a_91_75.n6 VNB 0.11fF
C156 a_91_75.n7 VNB 0.04fF
C157 a_1561_943.n0 VNB 0.06fF
C158 a_1561_943.n1 VNB 0.77fF
C159 a_1561_943.n2 VNB 0.77fF
C160 a_1561_943.n3 VNB 0.90fF
C161 a_1561_943.n4 VNB 0.28fF
C162 a_1561_943.n5 VNB 0.37fF
C163 a_1561_943.n6 VNB 0.47fF
C164 a_1561_943.n7 VNB 0.61fF
C165 a_1561_943.n8 VNB 0.47fF
C166 a_1561_943.t7 VNB 0.82fF
C167 a_1561_943.n9 VNB 0.52fF
C168 a_1561_943.n10 VNB 0.46fF
C169 a_1561_943.t9 VNB 0.82fF
C170 a_1561_943.n11 VNB 0.55fF
C171 a_1561_943.n12 VNB 1.81fF
C172 a_1561_943.n13 VNB 2.70fF
C173 a_1561_943.n14 VNB 0.64fF
C174 a_1561_943.n15 VNB 0.05fF
C175 a_1561_943.n16 VNB 0.49fF
C176 a_1561_943.n17 VNB 0.08fF
C177 a_599_943.n0 VNB 0.78fF
C178 a_599_943.n1 VNB 0.78fF
C179 a_599_943.n2 VNB 0.92fF
C180 a_599_943.n3 VNB 0.29fF
C181 a_599_943.n4 VNB 0.42fF
C182 a_599_943.n5 VNB 0.46fF
C183 a_599_943.n6 VNB 0.83fF
C184 a_599_943.n7 VNB 0.52fF
C185 a_599_943.t11 VNB 0.79fF
C186 a_599_943.n8 VNB 0.56fF
C187 a_599_943.n9 VNB 3.96fF
C188 a_599_943.n10 VNB 0.66fF
C189 a_599_943.n11 VNB 0.12fF
C190 a_599_943.n12 VNB 0.44fF
C191 a_599_943.n13 VNB 0.07fF
C192 a_277_1004.n0 VNB 0.50fF
C193 a_277_1004.n1 VNB 0.50fF
C194 a_277_1004.n2 VNB 0.58fF
C195 a_277_1004.n3 VNB 0.18fF
C196 a_277_1004.n4 VNB 0.32fF
C197 a_277_1004.n5 VNB 0.35fF
C198 a_277_1004.n6 VNB 0.44fF
C199 a_277_1004.n7 VNB 0.35fF
C200 a_277_1004.n8 VNB 0.43fF
C201 a_277_1004.n9 VNB 1.04fF
C202 a_277_1004.n10 VNB 0.42fF
C203 a_277_1004.n11 VNB 0.08fF
C204 a_277_1004.n12 VNB 0.22fF
C205 a_277_1004.n13 VNB 0.04fF
C206 VPB.n0 VNB 0.03fF
C207 VPB.n1 VNB 0.04fF
C208 VPB.n2 VNB 0.02fF
C209 VPB.n3 VNB 0.18fF
C210 VPB.n5 VNB 0.02fF
C211 VPB.n6 VNB 0.02fF
C212 VPB.n7 VNB 0.02fF
C213 VPB.n8 VNB 0.02fF
C214 VPB.n10 VNB 0.02fF
C215 VPB.n11 VNB 0.02fF
C216 VPB.n12 VNB 0.02fF
C217 VPB.n14 VNB 0.10fF
C218 VPB.n15 VNB 0.10fF
C219 VPB.n16 VNB 0.02fF
C220 VPB.n17 VNB 0.02fF
C221 VPB.n18 VNB 0.02fF
C222 VPB.n19 VNB 0.04fF
C223 VPB.n20 VNB 0.02fF
C224 VPB.n21 VNB 0.28fF
C225 VPB.n22 VNB 0.04fF
C226 VPB.n24 VNB 0.02fF
C227 VPB.n25 VNB 0.02fF
C228 VPB.n26 VNB 0.02fF
C229 VPB.n27 VNB 0.02fF
C230 VPB.n29 VNB 0.02fF
C231 VPB.n30 VNB 0.02fF
C232 VPB.n31 VNB 0.02fF
C233 VPB.n33 VNB 0.27fF
C234 VPB.n35 VNB 0.03fF
C235 VPB.n36 VNB 0.02fF
C236 VPB.n37 VNB 0.03fF
C237 VPB.n38 VNB 0.03fF
C238 VPB.n39 VNB 0.27fF
C239 VPB.n40 VNB 0.01fF
C240 VPB.n41 VNB 0.02fF
C241 VPB.n42 VNB 0.27fF
C242 VPB.n43 VNB 0.02fF
C243 VPB.n44 VNB 0.02fF
C244 VPB.n45 VNB 0.05fF
C245 VPB.n46 VNB 0.20fF
C246 VPB.n47 VNB 0.02fF
C247 VPB.n48 VNB 0.01fF
C248 VPB.n49 VNB 0.13fF
C249 VPB.n50 VNB 0.16fF
C250 VPB.n51 VNB 0.02fF
C251 VPB.n52 VNB 0.02fF
C252 VPB.n53 VNB 0.13fF
C253 VPB.n54 VNB 0.16fF
C254 VPB.n55 VNB 0.02fF
C255 VPB.n56 VNB 0.02fF
C256 VPB.n57 VNB 0.02fF
C257 VPB.n58 VNB 0.13fF
C258 VPB.n59 VNB 0.15fF
C259 VPB.n60 VNB 0.02fF
C260 VPB.n61 VNB 0.02fF
C261 VPB.n62 VNB 0.13fF
C262 VPB.n63 VNB 0.15fF
C263 VPB.n64 VNB 0.02fF
C264 VPB.n65 VNB 0.02fF
C265 VPB.n66 VNB 0.02fF
C266 VPB.n67 VNB 0.13fF
C267 VPB.n68 VNB 0.16fF
C268 VPB.n69 VNB 0.02fF
C269 VPB.n70 VNB 0.02fF
C270 VPB.n71 VNB 0.13fF
C271 VPB.n72 VNB 0.16fF
C272 VPB.n73 VNB 0.02fF
C273 VPB.n74 VNB 0.02fF
C274 VPB.n75 VNB 0.21fF
C275 VPB.n76 VNB 0.02fF
C276 VPB.n77 VNB 0.01fF
C277 VPB.n78 VNB 0.06fF
C278 VPB.n79 VNB 0.27fF
C279 VPB.n80 VNB 0.02fF
C280 VPB.n81 VNB 0.02fF
C281 VPB.n82 VNB 0.02fF
C282 VPB.n83 VNB 0.02fF
C283 VPB.n84 VNB 0.02fF
C284 VPB.n85 VNB 0.04fF
C285 VPB.n86 VNB 0.02fF
C286 VPB.n87 VNB 0.28fF
C287 VPB.n88 VNB 0.04fF
C288 VPB.n90 VNB 0.02fF
C289 VPB.n91 VNB 0.02fF
C290 VPB.n92 VNB 0.02fF
C291 VPB.n93 VNB 0.02fF
C292 VPB.n95 VNB 0.02fF
C293 VPB.n96 VNB 0.02fF
C294 VPB.n97 VNB 0.02fF
C295 VPB.n99 VNB 0.27fF
C296 VPB.n101 VNB 0.03fF
C297 VPB.n102 VNB 0.02fF
C298 VPB.n103 VNB 0.10fF
C299 VPB.n104 VNB 0.10fF
C300 VPB.n105 VNB 0.02fF
C301 VPB.n106 VNB 0.02fF
C302 VPB.n107 VNB 0.02fF
C303 VPB.n108 VNB 0.04fF
C304 VPB.n109 VNB 0.02fF
C305 VPB.n110 VNB 0.28fF
C306 VPB.n111 VNB 0.04fF
C307 VPB.n113 VNB 0.02fF
C308 VPB.n114 VNB 0.02fF
C309 VPB.n115 VNB 0.02fF
C310 VPB.n116 VNB 0.02fF
C311 VPB.n118 VNB 0.02fF
C312 VPB.n119 VNB 0.02fF
C313 VPB.n120 VNB 0.02fF
C314 VPB.n122 VNB 0.27fF
C315 VPB.n124 VNB 0.03fF
C316 VPB.n125 VNB 0.02fF
C317 VPB.n126 VNB 0.03fF
C318 VPB.n127 VNB 0.03fF
C319 VPB.n128 VNB 0.27fF
C320 VPB.n129 VNB 0.01fF
C321 VPB.n130 VNB 0.02fF
C322 VPB.n131 VNB 0.27fF
C323 VPB.n132 VNB 0.02fF
C324 VPB.n133 VNB 0.02fF
C325 VPB.n134 VNB 0.05fF
C326 VPB.n135 VNB 0.20fF
C327 VPB.n136 VNB 0.02fF
C328 VPB.n137 VNB 0.01fF
C329 VPB.n138 VNB 0.13fF
C330 VPB.n139 VNB 0.16fF
C331 VPB.n140 VNB 0.02fF
C332 VPB.n141 VNB 0.02fF
C333 VPB.n142 VNB 0.13fF
C334 VPB.n143 VNB 0.16fF
C335 VPB.n144 VNB 0.02fF
C336 VPB.n145 VNB 0.02fF
C337 VPB.n146 VNB 0.02fF
C338 VPB.n147 VNB 0.13fF
C339 VPB.n148 VNB 0.15fF
C340 VPB.n149 VNB 0.02fF
C341 VPB.n150 VNB 0.02fF
C342 VPB.n151 VNB 0.13fF
C343 VPB.n152 VNB 0.15fF
C344 VPB.n153 VNB 0.02fF
C345 VPB.n154 VNB 0.02fF
C346 VPB.n155 VNB 0.02fF
C347 VPB.n156 VNB 0.13fF
C348 VPB.n157 VNB 0.16fF
C349 VPB.n158 VNB 0.02fF
C350 VPB.n159 VNB 0.02fF
C351 VPB.n160 VNB 0.13fF
C352 VPB.n161 VNB 0.16fF
C353 VPB.n162 VNB 0.02fF
C354 VPB.n163 VNB 0.02fF
C355 VPB.n164 VNB 0.21fF
C356 VPB.n165 VNB 0.02fF
C357 VPB.n166 VNB 0.01fF
C358 VPB.n167 VNB 0.06fF
C359 VPB.n168 VNB 0.27fF
C360 VPB.n169 VNB 0.02fF
C361 VPB.n170 VNB 0.02fF
C362 VPB.n171 VNB 0.02fF
C363 VPB.n172 VNB 0.02fF
C364 VPB.n173 VNB 0.02fF
C365 VPB.n174 VNB 0.18fF
C366 VPB.n175 VNB 0.03fF
C367 VPB.n176 VNB 0.02fF
C368 VPB.n177 VNB 0.05fF
C369 VPB.n178 VNB 0.01fF
C370 VPB.n179 VNB 0.02fF
C371 VPB.n180 VNB 0.02fF
C372 VPB.n182 VNB 0.02fF
C373 VPB.n183 VNB 0.02fF
C374 VPB.n185 VNB 0.02fF
C375 VPB.n188 VNB 0.45fF
C376 VPB.n190 VNB 0.04fF
C377 VPB.n191 VNB 0.04fF
C378 VPB.n192 VNB 0.27fF
C379 VPB.n193 VNB 0.03fF
C380 VPB.n194 VNB 0.03fF
C381 VPB.n195 VNB 0.16fF
C382 VPB.n196 VNB 0.02fF
C383 VPB.n197 VNB 0.02fF
C384 VPB.n198 VNB 0.13fF
C385 VPB.n199 VNB 0.20fF
C386 VPB.n200 VNB 0.02fF
C387 VPB.n201 VNB 0.01fF
C388 VPB.n202 VNB 0.05fF
C389 VPB.n203 VNB 0.27fF
C390 VPB.n204 VNB 0.02fF
C391 VPB.n205 VNB 0.02fF
C392 VPB.n206 VNB 0.00fF
C393 VPB.n207 VNB 0.09fF
C394 VPB.n208 VNB 0.02fF
C395 VPB.n209 VNB 0.10fF
C396 VPB.n210 VNB 0.02fF
C397 VPB.n211 VNB 0.13fF
C398 VPB.n212 VNB 0.16fF
C399 VPB.n213 VNB 0.02fF
C400 VPB.n214 VNB 0.02fF
C401 VPB.n215 VNB 0.02fF
C402 VPB.n216 VNB 0.13fF
C403 VPB.n217 VNB 0.15fF
C404 VPB.n218 VNB 0.02fF
C405 VPB.n219 VNB 0.02fF
C406 VPB.n220 VNB 0.02fF
C407 VPB.n221 VNB 0.13fF
C408 VPB.n222 VNB 0.15fF
C409 VPB.n223 VNB 0.02fF
C410 VPB.n224 VNB 0.02fF
C411 VPB.n225 VNB 0.02fF
C412 VPB.n226 VNB 0.10fF
C413 VPB.n227 VNB 0.02fF
C414 VPB.n228 VNB 0.13fF
C415 VPB.n229 VNB 0.16fF
C416 VPB.n230 VNB 0.02fF
C417 VPB.n231 VNB 0.02fF
C418 VPB.n232 VNB 0.02fF
C419 VPB.n233 VNB 0.13fF
C420 VPB.n234 VNB 0.16fF
C421 VPB.n235 VNB 0.02fF
C422 VPB.n236 VNB 0.02fF
C423 VPB.n237 VNB 0.02fF
C424 VPB.n238 VNB 0.06fF
C425 VPB.n239 VNB 0.21fF
C426 VPB.n240 VNB 0.02fF
C427 VPB.n241 VNB 0.01fF
C428 VPB.n242 VNB 0.02fF
C429 VPB.n243 VNB 0.27fF
C430 VPB.n244 VNB 0.02fF
C431 VPB.n245 VNB 0.02fF
C432 VPB.n246 VNB 0.02fF
C433 VPB.n247 VNB 0.27fF
C434 VPB.n248 VNB 0.01fF
C435 VPB.n249 VNB 0.02fF
C436 VPB.n250 VNB 0.04fF
C437 VPB.n251 VNB 0.02fF
C438 VPB.n252 VNB 0.02fF
C439 VPB.n253 VNB 0.02fF
C440 VPB.n254 VNB 0.04fF
C441 VPB.n255 VNB 0.02fF
C442 VPB.n256 VNB 0.28fF
C443 VPB.n257 VNB 0.04fF
C444 VPB.n259 VNB 0.02fF
C445 VPB.n260 VNB 0.02fF
C446 VPB.n261 VNB 0.02fF
C447 VPB.n262 VNB 0.02fF
C448 VPB.n264 VNB 0.02fF
C449 VPB.n265 VNB 0.02fF
C450 VPB.n266 VNB 0.02fF
C451 VPB.n268 VNB 0.27fF
C452 VPB.n270 VNB 0.03fF
C453 VPB.n271 VNB 0.02fF
C454 VPB.n272 VNB 0.03fF
C455 VPB.n273 VNB 0.03fF
C456 VPB.n274 VNB 0.27fF
C457 VPB.n275 VNB 0.01fF
C458 VPB.n276 VNB 0.02fF
C459 VPB.n277 VNB 0.04fF
C460 VPB.n278 VNB 0.27fF
C461 VPB.n279 VNB 0.02fF
C462 VPB.n280 VNB 0.02fF
C463 VPB.n281 VNB 0.02fF
C464 VPB.n282 VNB 0.05fF
C465 VPB.n283 VNB 0.20fF
C466 VPB.n284 VNB 0.02fF
C467 VPB.n285 VNB 0.01fF
C468 VPB.n286 VNB 0.02fF
C469 VPB.n287 VNB 0.13fF
C470 VPB.n288 VNB 0.16fF
C471 VPB.n289 VNB 0.02fF
C472 VPB.n290 VNB 0.02fF
C473 VPB.n291 VNB 0.02fF
C474 VPB.n292 VNB 0.10fF
C475 VPB.n293 VNB 0.02fF
C476 VPB.n294 VNB 0.13fF
C477 VPB.n295 VNB 0.16fF
C478 VPB.n296 VNB 0.02fF
C479 VPB.n297 VNB 0.02fF
C480 VPB.n298 VNB 0.02fF
C481 VPB.n299 VNB 0.13fF
C482 VPB.n300 VNB 0.15fF
C483 VPB.n301 VNB 0.02fF
C484 VPB.n302 VNB 0.02fF
C485 VPB.n303 VNB 0.02fF
C486 VPB.n304 VNB 0.13fF
C487 VPB.n305 VNB 0.15fF
C488 VPB.n306 VNB 0.02fF
C489 VPB.n307 VNB 0.02fF
C490 VPB.n308 VNB 0.02fF
C491 VPB.n309 VNB 0.10fF
C492 VPB.n310 VNB 0.02fF
C493 VPB.n311 VNB 0.13fF
C494 VPB.n312 VNB 0.16fF
C495 VPB.n313 VNB 0.02fF
C496 VPB.n314 VNB 0.02fF
C497 VPB.n315 VNB 0.02fF
C498 VPB.n316 VNB 0.13fF
C499 VPB.n317 VNB 0.16fF
C500 VPB.n318 VNB 0.02fF
C501 VPB.n319 VNB 0.02fF
C502 VPB.n320 VNB 0.02fF
C503 VPB.n321 VNB 0.06fF
C504 VPB.n322 VNB 0.21fF
C505 VPB.n323 VNB 0.02fF
C506 VPB.n324 VNB 0.01fF
C507 VPB.n325 VNB 0.02fF
C508 VPB.n326 VNB 0.27fF
C509 VPB.n327 VNB 0.02fF
C510 VPB.n328 VNB 0.02fF
C511 VPB.n329 VNB 0.02fF
C512 VPB.n330 VNB 0.27fF
C513 VPB.n331 VNB 0.01fF
C514 VPB.n332 VNB 0.02fF
C515 VPB.n333 VNB 0.04fF
C516 VPB.n334 VNB 0.04fF
C517 VPB.n335 VNB 0.02fF
C518 VPB.n336 VNB 0.02fF
C519 VPB.n337 VNB 0.02fF
C520 VPB.n338 VNB 0.02fF
C521 VPB.n339 VNB 0.02fF
C522 VPB.n340 VNB 0.02fF
C523 VPB.n341 VNB 0.02fF
C524 VPB.n342 VNB 0.02fF
C525 VPB.n343 VNB 0.02fF
C526 VPB.n344 VNB 0.02fF
C527 VPB.n345 VNB 0.02fF
C528 VPB.n346 VNB 0.27fF
C529 VPB.n347 VNB 0.01fF
C530 VPB.n348 VNB 0.02fF
C531 VPB.n349 VNB 0.03fF
C532 VPB.n350 VNB 0.03fF
C533 VPB.n351 VNB 0.27fF
C534 VPB.n352 VNB 0.01fF
C535 VPB.n353 VNB 0.02fF
C536 VPB.n354 VNB 0.02fF
C537 VPB.n355 VNB 0.27fF
C538 VPB.n356 VNB 0.02fF
C539 VPB.n357 VNB 0.02fF
C540 VPB.n358 VNB 0.02fF
C541 VPB.n359 VNB 0.05fF
C542 VPB.n360 VNB 0.20fF
C543 VPB.n361 VNB 0.02fF
C544 VPB.n362 VNB 0.01fF
C545 VPB.n363 VNB 0.02fF
C546 VPB.n364 VNB 0.13fF
C547 VPB.n365 VNB 0.16fF
C548 VPB.n366 VNB 0.02fF
C549 VPB.n367 VNB 0.02fF
C550 VPB.n368 VNB 0.02fF
C551 VPB.n369 VNB 0.10fF
C552 VPB.n370 VNB 0.02fF
C553 VPB.n371 VNB 0.13fF
C554 VPB.n372 VNB 0.16fF
C555 VPB.n373 VNB 0.02fF
C556 VPB.n374 VNB 0.02fF
C557 VPB.n375 VNB 0.02fF
C558 VPB.n376 VNB 0.13fF
C559 VPB.n377 VNB 0.15fF
C560 VPB.n378 VNB 0.02fF
C561 VPB.n379 VNB 0.02fF
C562 VPB.n380 VNB 0.02fF
C563 VPB.n381 VNB 0.13fF
C564 VPB.n382 VNB 0.15fF
C565 VPB.n383 VNB 0.02fF
C566 VPB.n384 VNB 0.02fF
C567 VPB.n385 VNB 0.02fF
C568 VPB.n386 VNB 0.10fF
C569 VPB.n387 VNB 0.02fF
C570 VPB.n388 VNB 0.13fF
C571 VPB.n389 VNB 0.16fF
C572 VPB.n390 VNB 0.02fF
C573 VPB.n391 VNB 0.02fF
C574 VPB.n392 VNB 0.02fF
C575 VPB.n393 VNB 0.13fF
C576 VPB.n394 VNB 0.16fF
C577 VPB.n395 VNB 0.02fF
C578 VPB.n396 VNB 0.02fF
C579 VPB.n397 VNB 0.02fF
C580 VPB.n398 VNB 0.06fF
C581 VPB.n399 VNB 0.21fF
C582 VPB.n400 VNB 0.02fF
C583 VPB.n401 VNB 0.01fF
C584 VPB.n402 VNB 0.02fF
C585 VPB.n403 VNB 0.27fF
C586 VPB.n404 VNB 0.02fF
C587 VPB.n405 VNB 0.02fF
C588 VPB.n406 VNB 0.02fF
C589 VPB.n407 VNB 0.27fF
C590 VPB.n408 VNB 0.01fF
C591 VPB.n409 VNB 0.02fF
C592 VPB.n410 VNB 0.04fF
C593 VPB.n411 VNB 0.02fF
C594 VPB.n412 VNB 0.02fF
C595 VPB.n413 VNB 0.02fF
C596 VPB.n414 VNB 0.04fF
C597 VPB.n415 VNB 0.02fF
C598 VPB.n416 VNB 0.28fF
C599 VPB.n417 VNB 0.04fF
C600 VPB.n419 VNB 0.02fF
C601 VPB.n420 VNB 0.02fF
C602 VPB.n421 VNB 0.02fF
C603 VPB.n422 VNB 0.02fF
C604 VPB.n424 VNB 0.02fF
C605 VPB.n425 VNB 0.02fF
C606 VPB.n426 VNB 0.02fF
C607 VPB.n428 VNB 0.27fF
C608 VPB.n430 VNB 0.03fF
C609 VPB.n431 VNB 0.02fF
C610 VPB.n432 VNB 0.03fF
C611 VPB.n433 VNB 0.03fF
C612 VPB.n434 VNB 0.27fF
C613 VPB.n435 VNB 0.01fF
C614 VPB.n436 VNB 0.02fF
C615 VPB.n437 VNB 0.04fF
C616 VPB.n438 VNB 0.27fF
C617 VPB.n439 VNB 0.02fF
C618 VPB.n440 VNB 0.02fF
C619 VPB.n441 VNB 0.02fF
C620 VPB.n442 VNB 0.05fF
C621 VPB.n443 VNB 0.20fF
C622 VPB.n444 VNB 0.02fF
C623 VPB.n445 VNB 0.01fF
C624 VPB.n446 VNB 0.02fF
C625 VPB.n447 VNB 0.13fF
C626 VPB.n448 VNB 0.16fF
C627 VPB.n449 VNB 0.02fF
C628 VPB.n450 VNB 0.02fF
C629 VPB.n451 VNB 0.02fF
C630 VPB.n452 VNB 0.10fF
C631 VPB.n453 VNB 0.02fF
C632 VPB.n454 VNB 0.13fF
C633 VPB.n455 VNB 0.16fF
C634 VPB.n456 VNB 0.02fF
C635 VPB.n457 VNB 0.02fF
C636 VPB.n458 VNB 0.02fF
C637 VPB.n459 VNB 0.13fF
C638 VPB.n460 VNB 0.15fF
C639 VPB.n461 VNB 0.02fF
C640 VPB.n462 VNB 0.02fF
C641 VPB.n463 VNB 0.02fF
C642 VPB.n464 VNB 0.13fF
C643 VPB.n465 VNB 0.15fF
C644 VPB.n466 VNB 0.02fF
C645 VPB.n467 VNB 0.02fF
C646 VPB.n468 VNB 0.02fF
C647 VPB.n469 VNB 0.10fF
C648 VPB.n470 VNB 0.02fF
C649 VPB.n471 VNB 0.13fF
C650 VPB.n472 VNB 0.16fF
C651 VPB.n473 VNB 0.02fF
C652 VPB.n474 VNB 0.02fF
C653 VPB.n475 VNB 0.02fF
C654 VPB.n476 VNB 0.13fF
C655 VPB.n477 VNB 0.16fF
C656 VPB.n478 VNB 0.02fF
C657 VPB.n479 VNB 0.02fF
C658 VPB.n480 VNB 0.02fF
C659 VPB.n481 VNB 0.06fF
C660 VPB.n482 VNB 0.21fF
C661 VPB.n483 VNB 0.02fF
C662 VPB.n484 VNB 0.01fF
C663 VPB.n485 VNB 0.02fF
C664 VPB.n486 VNB 0.27fF
C665 VPB.n487 VNB 0.02fF
C666 VPB.n488 VNB 0.02fF
C667 VPB.n489 VNB 0.02fF
C668 VPB.n490 VNB 0.27fF
C669 VPB.n491 VNB 0.01fF
C670 VPB.n492 VNB 0.02fF
C671 VPB.n493 VNB 0.04fF
C672 VPB.n494 VNB 0.04fF
C673 VPB.n495 VNB 0.02fF
C674 VPB.n496 VNB 0.02fF
C675 VPB.n497 VNB 0.02fF
C676 VPB.n498 VNB 0.02fF
C677 VPB.n499 VNB 0.02fF
C678 VPB.n500 VNB 0.02fF
C679 VPB.n501 VNB 0.02fF
C680 VPB.n502 VNB 0.02fF
C681 VPB.n503 VNB 0.02fF
C682 VPB.n504 VNB 0.02fF
C683 VPB.n505 VNB 0.03fF
C684 VPB.n506 VNB 0.03fF
C685 VPB.n507 VNB 0.02fF
C686 VPB.n508 VNB 0.02fF
C687 VPB.n509 VNB 0.02fF
C688 VPB.n510 VNB 0.04fF
C689 VPB.n511 VNB 0.04fF
C690 VPB.n513 VNB 0.42fF
.ends
