magic
tech sky130A
magscale 1 2
timestamp 1649525376
<< metal1 >>
rect 315 501 569 535
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 592 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 296 0 -1 518
box -53 -33 29 33
use invx1_pcell  invx1_pcell_1
timestamp 1648064504
transform 1 0 444 0 1 0
box -84 0 528 1575
use invx1_pcell  invx1_pcell_0
timestamp 1648064504
transform 1 0 0 0 1 0
box -84 0 528 1575
<< end >>
