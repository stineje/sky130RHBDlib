magic
tech sky130A
magscale 1 2
timestamp 1669564293
<< nwell >>
rect -87 786 4527 1550
<< pwell >>
rect -34 -34 4474 544
<< nmos >>
rect 155 297 185 350
tri 185 297 201 313 sw
rect 155 267 261 297
tri 261 267 291 297 sw
rect 155 166 185 267
tri 185 251 201 267 nw
tri 245 251 261 267 ne
tri 185 166 201 182 sw
tri 245 166 261 182 se
rect 261 166 291 267
tri 155 136 185 166 ne
rect 185 136 261 166
tri 261 136 291 166 nw
rect 599 297 629 350
tri 629 297 645 313 sw
rect 599 267 705 297
tri 705 267 735 297 sw
rect 599 166 629 267
tri 629 251 645 267 nw
tri 689 251 705 267 ne
tri 629 166 645 182 sw
tri 689 166 705 182 se
rect 705 166 735 267
tri 599 136 629 166 ne
rect 629 136 705 166
tri 705 136 735 166 nw
rect 1056 288 1086 349
tri 1086 288 1102 304 sw
rect 1250 296 1280 349
tri 1280 296 1296 312 sw
rect 1056 258 1162 288
tri 1162 258 1192 288 sw
rect 1250 266 1356 296
tri 1356 266 1386 296 sw
rect 1056 157 1086 258
tri 1086 242 1102 258 nw
tri 1146 242 1162 258 ne
tri 1086 157 1102 173 sw
tri 1146 157 1162 173 se
rect 1162 157 1192 258
rect 1250 165 1280 266
tri 1280 250 1296 266 nw
tri 1340 250 1356 266 ne
tri 1280 165 1296 181 sw
tri 1340 165 1356 181 se
rect 1356 165 1386 266
tri 1056 127 1086 157 ne
rect 1086 127 1162 157
tri 1162 127 1192 157 nw
tri 1250 135 1280 165 ne
rect 1280 135 1356 165
tri 1356 135 1386 165 nw
rect 1709 297 1739 350
tri 1739 297 1755 313 sw
rect 1709 267 1815 297
tri 1815 267 1845 297 sw
rect 1709 166 1739 267
tri 1739 251 1755 267 nw
tri 1799 251 1815 267 ne
tri 1739 166 1755 182 sw
tri 1799 166 1815 182 se
rect 1815 166 1845 267
tri 1709 136 1739 166 ne
rect 1739 136 1815 166
tri 1815 136 1845 166 nw
rect 2166 288 2196 349
tri 2196 288 2212 304 sw
rect 2360 296 2390 349
tri 2390 296 2406 312 sw
rect 2166 258 2272 288
tri 2272 258 2302 288 sw
rect 2360 266 2466 296
tri 2466 266 2496 296 sw
rect 2166 157 2196 258
tri 2196 242 2212 258 nw
tri 2256 242 2272 258 ne
tri 2196 157 2212 173 sw
tri 2256 157 2272 173 se
rect 2272 157 2302 258
rect 2360 165 2390 266
tri 2390 250 2406 266 nw
tri 2450 250 2466 266 ne
tri 2390 165 2406 181 sw
tri 2450 165 2466 181 se
rect 2466 165 2496 266
tri 2166 127 2196 157 ne
rect 2196 127 2272 157
tri 2272 127 2302 157 nw
tri 2360 135 2390 165 ne
rect 2390 135 2466 165
tri 2466 135 2496 165 nw
rect 2819 297 2849 350
tri 2849 297 2865 313 sw
rect 2819 267 2925 297
tri 2925 267 2955 297 sw
rect 2819 166 2849 267
tri 2849 251 2865 267 nw
tri 2909 251 2925 267 ne
tri 2849 166 2865 182 sw
tri 2909 166 2925 182 se
rect 2925 166 2955 267
tri 2819 136 2849 166 ne
rect 2849 136 2925 166
tri 2925 136 2955 166 nw
rect 3276 296 3306 349
tri 3306 296 3322 312 sw
rect 3470 296 3500 349
tri 3500 296 3516 312 sw
rect 3276 266 3382 296
tri 3382 266 3412 296 sw
rect 3276 165 3306 266
tri 3306 250 3322 266 nw
tri 3366 250 3382 266 ne
tri 3306 165 3322 181 sw
tri 3366 165 3382 181 se
rect 3382 165 3412 266
rect 3470 266 3576 296
tri 3576 266 3606 296 sw
rect 3470 251 3501 266
tri 3501 251 3516 266 nw
tri 3560 251 3575 266 ne
rect 3575 251 3606 266
tri 3276 135 3306 165 ne
rect 3306 135 3382 165
tri 3382 135 3412 165 nw
rect 3470 165 3500 251
tri 3500 165 3516 181 sw
tri 3560 165 3576 181 se
rect 3576 165 3606 251
tri 3470 135 3500 165 ne
rect 3500 135 3576 165
tri 3576 135 3606 165 nw
rect 3942 296 3972 349
tri 3972 296 3988 312 sw
rect 4136 296 4166 349
tri 4166 296 4182 312 sw
rect 3942 266 4048 296
tri 4048 266 4078 296 sw
rect 3942 165 3972 266
tri 3972 250 3988 266 nw
tri 4032 250 4048 266 ne
tri 3972 165 3988 181 sw
tri 4032 165 4048 181 se
rect 4048 165 4078 266
rect 4136 266 4242 296
tri 4242 266 4272 296 sw
rect 4136 251 4167 266
tri 4167 251 4182 266 nw
tri 4226 251 4241 266 ne
rect 4241 251 4272 266
tri 3942 135 3972 165 ne
rect 3972 135 4048 165
tri 4048 135 4078 165 nw
rect 4136 165 4166 251
tri 4166 165 4182 181 sw
tri 4226 165 4242 181 se
rect 4242 165 4272 251
tri 4136 135 4166 165 ne
rect 4166 135 4242 165
tri 4242 135 4272 165 nw
<< pmos >>
rect 164 1004 194 1404
rect 252 1004 282 1404
rect 608 1004 638 1404
rect 696 1004 726 1404
rect 1075 1004 1105 1404
rect 1163 1004 1193 1404
rect 1251 1004 1281 1404
rect 1339 1004 1369 1404
rect 1718 1004 1748 1404
rect 1806 1004 1836 1404
rect 2185 1004 2215 1404
rect 2273 1004 2303 1404
rect 2361 1004 2391 1404
rect 2449 1004 2479 1404
rect 2828 1004 2858 1404
rect 2916 1004 2946 1404
rect 3295 1005 3325 1405
rect 3383 1005 3413 1405
rect 3471 1005 3501 1405
rect 3559 1005 3589 1405
rect 3961 1005 3991 1405
rect 4049 1005 4079 1405
rect 4137 1005 4167 1405
rect 4225 1005 4255 1405
<< ndiff >>
rect 99 334 155 350
rect 99 300 109 334
rect 143 300 155 334
rect 99 262 155 300
rect 185 334 345 350
rect 185 313 303 334
tri 185 297 201 313 ne
rect 201 300 303 313
rect 337 300 345 334
rect 201 297 345 300
tri 261 267 291 297 ne
rect 99 228 109 262
rect 143 228 155 262
rect 99 194 155 228
rect 99 160 109 194
rect 143 160 155 194
tri 185 251 201 267 se
rect 201 251 245 267
tri 245 251 261 267 sw
rect 185 218 261 251
rect 185 184 205 218
rect 239 184 261 218
rect 185 182 261 184
tri 185 166 201 182 ne
rect 201 166 245 182
tri 245 166 261 182 nw
rect 291 262 345 297
rect 291 228 303 262
rect 337 228 345 262
rect 291 194 345 228
rect 99 136 155 160
tri 155 136 185 166 sw
tri 261 136 291 166 se
rect 291 160 303 194
rect 337 160 345 194
rect 291 136 345 160
rect 99 124 345 136
rect 99 90 109 124
rect 143 90 205 124
rect 239 90 303 124
rect 337 90 345 124
rect 99 74 345 90
rect 543 334 599 350
rect 543 300 553 334
rect 587 300 599 334
rect 543 262 599 300
rect 629 334 789 350
rect 629 313 747 334
tri 629 297 645 313 ne
rect 645 300 747 313
rect 781 300 789 334
rect 645 297 789 300
tri 705 267 735 297 ne
rect 543 228 553 262
rect 587 228 599 262
rect 543 194 599 228
rect 543 160 553 194
rect 587 160 599 194
tri 629 251 645 267 se
rect 645 251 689 267
tri 689 251 705 267 sw
rect 629 218 705 251
rect 629 184 649 218
rect 683 184 705 218
rect 629 182 705 184
tri 629 166 645 182 ne
rect 645 166 689 182
tri 689 166 705 182 nw
rect 735 262 789 297
rect 735 228 747 262
rect 781 228 789 262
rect 735 194 789 228
rect 543 136 599 160
tri 599 136 629 166 sw
tri 705 136 735 166 se
rect 735 160 747 194
rect 781 160 789 194
rect 735 136 789 160
rect 543 124 789 136
rect 543 90 553 124
rect 587 90 649 124
rect 683 90 747 124
rect 781 90 789 124
rect 543 74 789 90
rect 1000 333 1056 349
rect 1000 299 1010 333
rect 1044 299 1056 333
rect 1000 261 1056 299
rect 1086 333 1250 349
rect 1086 304 1107 333
tri 1086 288 1102 304 ne
rect 1102 299 1107 304
rect 1141 299 1204 333
rect 1238 299 1250 333
rect 1102 288 1250 299
rect 1280 312 1442 349
tri 1280 296 1296 312 ne
rect 1296 296 1442 312
rect 1000 227 1010 261
rect 1044 227 1056 261
tri 1162 258 1192 288 ne
rect 1192 261 1250 288
tri 1356 266 1386 296 ne
rect 1000 193 1056 227
rect 1000 159 1010 193
rect 1044 159 1056 193
rect 1000 127 1056 159
tri 1086 242 1102 258 se
rect 1102 242 1146 258
tri 1146 242 1162 258 sw
rect 1086 208 1162 242
rect 1086 174 1107 208
rect 1141 174 1162 208
rect 1086 173 1162 174
tri 1086 157 1102 173 ne
rect 1102 157 1146 173
tri 1146 157 1162 173 nw
rect 1192 227 1204 261
rect 1238 227 1250 261
rect 1192 193 1250 227
rect 1192 159 1204 193
rect 1238 159 1250 193
tri 1280 250 1296 266 se
rect 1296 250 1340 266
tri 1340 250 1356 266 sw
rect 1280 217 1356 250
rect 1280 183 1301 217
rect 1335 183 1356 217
rect 1280 181 1356 183
tri 1280 165 1296 181 ne
rect 1296 165 1340 181
tri 1340 165 1356 181 nw
rect 1386 261 1442 296
rect 1386 227 1398 261
rect 1432 227 1442 261
rect 1386 193 1442 227
tri 1056 127 1086 157 sw
tri 1162 127 1192 157 se
rect 1192 135 1250 159
tri 1250 135 1280 165 sw
tri 1356 135 1386 165 se
rect 1386 159 1398 193
rect 1432 159 1442 193
rect 1386 135 1442 159
rect 1192 127 1442 135
rect 1000 123 1442 127
rect 1000 89 1010 123
rect 1044 89 1204 123
rect 1238 89 1301 123
rect 1335 89 1398 123
rect 1432 89 1442 123
rect 1000 73 1442 89
rect 1653 334 1709 350
rect 1653 300 1663 334
rect 1697 300 1709 334
rect 1653 262 1709 300
rect 1739 334 1899 350
rect 1739 313 1857 334
tri 1739 297 1755 313 ne
rect 1755 300 1857 313
rect 1891 300 1899 334
rect 1755 297 1899 300
tri 1815 267 1845 297 ne
rect 1653 228 1663 262
rect 1697 228 1709 262
rect 1653 194 1709 228
rect 1653 160 1663 194
rect 1697 160 1709 194
tri 1739 251 1755 267 se
rect 1755 251 1799 267
tri 1799 251 1815 267 sw
rect 1739 218 1815 251
rect 1739 184 1759 218
rect 1793 184 1815 218
rect 1739 182 1815 184
tri 1739 166 1755 182 ne
rect 1755 166 1799 182
tri 1799 166 1815 182 nw
rect 1845 262 1899 297
rect 1845 228 1857 262
rect 1891 228 1899 262
rect 1845 194 1899 228
rect 1653 136 1709 160
tri 1709 136 1739 166 sw
tri 1815 136 1845 166 se
rect 1845 160 1857 194
rect 1891 160 1899 194
rect 1845 136 1899 160
rect 1653 124 1899 136
rect 1653 90 1663 124
rect 1697 90 1759 124
rect 1793 90 1857 124
rect 1891 90 1899 124
rect 1653 74 1899 90
rect 2110 333 2166 349
rect 2110 299 2120 333
rect 2154 299 2166 333
rect 2110 261 2166 299
rect 2196 333 2360 349
rect 2196 304 2217 333
tri 2196 288 2212 304 ne
rect 2212 299 2217 304
rect 2251 299 2314 333
rect 2348 299 2360 333
rect 2212 288 2360 299
rect 2390 312 2552 349
tri 2390 296 2406 312 ne
rect 2406 296 2552 312
rect 2110 227 2120 261
rect 2154 227 2166 261
tri 2272 258 2302 288 ne
rect 2302 261 2360 288
tri 2466 266 2496 296 ne
rect 2110 193 2166 227
rect 2110 159 2120 193
rect 2154 159 2166 193
rect 2110 127 2166 159
tri 2196 242 2212 258 se
rect 2212 242 2256 258
tri 2256 242 2272 258 sw
rect 2196 208 2272 242
rect 2196 174 2217 208
rect 2251 174 2272 208
rect 2196 173 2272 174
tri 2196 157 2212 173 ne
rect 2212 157 2256 173
tri 2256 157 2272 173 nw
rect 2302 227 2314 261
rect 2348 227 2360 261
rect 2302 193 2360 227
rect 2302 159 2314 193
rect 2348 159 2360 193
tri 2390 250 2406 266 se
rect 2406 250 2450 266
tri 2450 250 2466 266 sw
rect 2390 217 2466 250
rect 2390 183 2411 217
rect 2445 183 2466 217
rect 2390 181 2466 183
tri 2390 165 2406 181 ne
rect 2406 165 2450 181
tri 2450 165 2466 181 nw
rect 2496 261 2552 296
rect 2496 227 2508 261
rect 2542 227 2552 261
rect 2496 193 2552 227
tri 2166 127 2196 157 sw
tri 2272 127 2302 157 se
rect 2302 135 2360 159
tri 2360 135 2390 165 sw
tri 2466 135 2496 165 se
rect 2496 159 2508 193
rect 2542 159 2552 193
rect 2496 135 2552 159
rect 2302 127 2552 135
rect 2110 123 2552 127
rect 2110 89 2120 123
rect 2154 89 2314 123
rect 2348 89 2411 123
rect 2445 89 2508 123
rect 2542 89 2552 123
rect 2110 73 2552 89
rect 2763 334 2819 350
rect 2763 300 2773 334
rect 2807 300 2819 334
rect 2763 262 2819 300
rect 2849 334 3009 350
rect 2849 313 2967 334
tri 2849 297 2865 313 ne
rect 2865 300 2967 313
rect 3001 300 3009 334
rect 2865 297 3009 300
tri 2925 267 2955 297 ne
rect 2763 228 2773 262
rect 2807 228 2819 262
rect 2763 194 2819 228
rect 2763 160 2773 194
rect 2807 160 2819 194
tri 2849 251 2865 267 se
rect 2865 251 2909 267
tri 2909 251 2925 267 sw
rect 2849 218 2925 251
rect 2849 184 2869 218
rect 2903 184 2925 218
rect 2849 182 2925 184
tri 2849 166 2865 182 ne
rect 2865 166 2909 182
tri 2909 166 2925 182 nw
rect 2955 262 3009 297
rect 2955 228 2967 262
rect 3001 228 3009 262
rect 2955 194 3009 228
rect 2763 136 2819 160
tri 2819 136 2849 166 sw
tri 2925 136 2955 166 se
rect 2955 160 2967 194
rect 3001 160 3009 194
rect 2955 136 3009 160
rect 2763 124 3009 136
rect 2763 90 2773 124
rect 2807 90 2869 124
rect 2903 90 2967 124
rect 3001 90 3009 124
rect 2763 74 3009 90
rect 3220 333 3276 349
rect 3220 299 3230 333
rect 3264 299 3276 333
rect 3220 261 3276 299
rect 3306 312 3470 349
tri 3306 296 3322 312 ne
rect 3322 296 3470 312
rect 3500 312 3662 349
tri 3500 296 3516 312 ne
rect 3516 296 3662 312
tri 3382 266 3412 296 ne
rect 3220 227 3230 261
rect 3264 227 3276 261
rect 3220 193 3276 227
rect 3220 159 3230 193
rect 3264 159 3276 193
tri 3306 250 3322 266 se
rect 3322 250 3366 266
tri 3366 250 3382 266 sw
rect 3306 217 3382 250
rect 3306 183 3327 217
rect 3361 183 3382 217
rect 3306 181 3382 183
tri 3306 165 3322 181 ne
rect 3322 165 3366 181
tri 3366 165 3382 181 nw
rect 3412 261 3470 296
tri 3576 266 3606 296 ne
rect 3412 227 3424 261
rect 3458 227 3470 261
tri 3501 251 3516 266 se
rect 3516 251 3560 266
tri 3560 251 3575 266 sw
rect 3606 261 3662 296
rect 3412 193 3470 227
rect 3220 135 3276 159
tri 3276 135 3306 165 sw
tri 3382 135 3412 165 se
rect 3412 159 3424 193
rect 3458 159 3470 193
rect 3500 217 3576 251
rect 3500 183 3521 217
rect 3555 183 3576 217
rect 3500 181 3576 183
tri 3500 165 3516 181 ne
rect 3516 165 3560 181
tri 3560 165 3576 181 nw
rect 3606 227 3618 261
rect 3652 227 3662 261
rect 3606 193 3662 227
rect 3412 135 3470 159
tri 3470 135 3500 165 sw
tri 3576 135 3606 165 se
rect 3606 159 3618 193
rect 3652 159 3662 193
rect 3606 135 3662 159
rect 3220 123 3662 135
rect 3220 89 3230 123
rect 3264 89 3327 123
rect 3361 89 3424 123
rect 3458 89 3521 123
rect 3555 89 3618 123
rect 3652 89 3662 123
rect 3220 73 3662 89
rect 3886 333 3942 349
rect 3886 299 3896 333
rect 3930 299 3942 333
rect 3886 261 3942 299
rect 3972 312 4136 349
tri 3972 296 3988 312 ne
rect 3988 296 4136 312
rect 4166 312 4328 349
tri 4166 296 4182 312 ne
rect 4182 296 4328 312
tri 4048 266 4078 296 ne
rect 3886 227 3896 261
rect 3930 227 3942 261
rect 3886 193 3942 227
rect 3886 159 3896 193
rect 3930 159 3942 193
tri 3972 250 3988 266 se
rect 3988 250 4032 266
tri 4032 250 4048 266 sw
rect 3972 217 4048 250
rect 3972 183 3993 217
rect 4027 183 4048 217
rect 3972 181 4048 183
tri 3972 165 3988 181 ne
rect 3988 165 4032 181
tri 4032 165 4048 181 nw
rect 4078 261 4136 296
tri 4242 266 4272 296 ne
rect 4078 227 4090 261
rect 4124 227 4136 261
tri 4167 251 4182 266 se
rect 4182 251 4226 266
tri 4226 251 4241 266 sw
rect 4272 261 4328 296
rect 4078 193 4136 227
rect 3886 135 3942 159
tri 3942 135 3972 165 sw
tri 4048 135 4078 165 se
rect 4078 159 4090 193
rect 4124 159 4136 193
rect 4166 217 4242 251
rect 4166 183 4187 217
rect 4221 183 4242 217
rect 4166 181 4242 183
tri 4166 165 4182 181 ne
rect 4182 165 4226 181
tri 4226 165 4242 181 nw
rect 4272 227 4284 261
rect 4318 227 4328 261
rect 4272 193 4328 227
rect 4078 135 4136 159
tri 4136 135 4166 165 sw
tri 4242 135 4272 165 se
rect 4272 159 4284 193
rect 4318 159 4328 193
rect 4272 135 4328 159
rect 3886 123 4328 135
rect 3886 89 3896 123
rect 3930 89 3993 123
rect 4027 89 4090 123
rect 4124 89 4187 123
rect 4221 89 4284 123
rect 4318 89 4328 123
rect 3886 73 4328 89
<< pdiff >>
rect 108 1366 164 1404
rect 108 1332 118 1366
rect 152 1332 164 1366
rect 108 1298 164 1332
rect 108 1264 118 1298
rect 152 1264 164 1298
rect 108 1230 164 1264
rect 108 1196 118 1230
rect 152 1196 164 1230
rect 108 1162 164 1196
rect 108 1128 118 1162
rect 152 1128 164 1162
rect 108 1093 164 1128
rect 108 1059 118 1093
rect 152 1059 164 1093
rect 108 1004 164 1059
rect 194 1366 252 1404
rect 194 1332 206 1366
rect 240 1332 252 1366
rect 194 1298 252 1332
rect 194 1264 206 1298
rect 240 1264 252 1298
rect 194 1230 252 1264
rect 194 1196 206 1230
rect 240 1196 252 1230
rect 194 1162 252 1196
rect 194 1128 206 1162
rect 240 1128 252 1162
rect 194 1093 252 1128
rect 194 1059 206 1093
rect 240 1059 252 1093
rect 194 1004 252 1059
rect 282 1366 336 1404
rect 282 1332 294 1366
rect 328 1332 336 1366
rect 282 1298 336 1332
rect 282 1264 294 1298
rect 328 1264 336 1298
rect 282 1230 336 1264
rect 282 1196 294 1230
rect 328 1196 336 1230
rect 282 1162 336 1196
rect 282 1128 294 1162
rect 328 1128 336 1162
rect 282 1093 336 1128
rect 282 1059 294 1093
rect 328 1059 336 1093
rect 282 1004 336 1059
rect 552 1366 608 1404
rect 552 1332 562 1366
rect 596 1332 608 1366
rect 552 1298 608 1332
rect 552 1264 562 1298
rect 596 1264 608 1298
rect 552 1230 608 1264
rect 552 1196 562 1230
rect 596 1196 608 1230
rect 552 1162 608 1196
rect 552 1128 562 1162
rect 596 1128 608 1162
rect 552 1093 608 1128
rect 552 1059 562 1093
rect 596 1059 608 1093
rect 552 1004 608 1059
rect 638 1366 696 1404
rect 638 1332 650 1366
rect 684 1332 696 1366
rect 638 1298 696 1332
rect 638 1264 650 1298
rect 684 1264 696 1298
rect 638 1230 696 1264
rect 638 1196 650 1230
rect 684 1196 696 1230
rect 638 1162 696 1196
rect 638 1128 650 1162
rect 684 1128 696 1162
rect 638 1093 696 1128
rect 638 1059 650 1093
rect 684 1059 696 1093
rect 638 1004 696 1059
rect 726 1366 780 1404
rect 726 1332 738 1366
rect 772 1332 780 1366
rect 726 1298 780 1332
rect 726 1264 738 1298
rect 772 1264 780 1298
rect 726 1230 780 1264
rect 726 1196 738 1230
rect 772 1196 780 1230
rect 726 1162 780 1196
rect 726 1128 738 1162
rect 772 1128 780 1162
rect 726 1093 780 1128
rect 726 1059 738 1093
rect 772 1059 780 1093
rect 726 1004 780 1059
rect 1019 1366 1075 1404
rect 1019 1332 1029 1366
rect 1063 1332 1075 1366
rect 1019 1298 1075 1332
rect 1019 1264 1029 1298
rect 1063 1264 1075 1298
rect 1019 1230 1075 1264
rect 1019 1196 1029 1230
rect 1063 1196 1075 1230
rect 1019 1162 1075 1196
rect 1019 1128 1029 1162
rect 1063 1128 1075 1162
rect 1019 1093 1075 1128
rect 1019 1059 1029 1093
rect 1063 1059 1075 1093
rect 1019 1004 1075 1059
rect 1105 1366 1163 1404
rect 1105 1332 1117 1366
rect 1151 1332 1163 1366
rect 1105 1298 1163 1332
rect 1105 1264 1117 1298
rect 1151 1264 1163 1298
rect 1105 1230 1163 1264
rect 1105 1196 1117 1230
rect 1151 1196 1163 1230
rect 1105 1162 1163 1196
rect 1105 1128 1117 1162
rect 1151 1128 1163 1162
rect 1105 1093 1163 1128
rect 1105 1059 1117 1093
rect 1151 1059 1163 1093
rect 1105 1004 1163 1059
rect 1193 1366 1251 1404
rect 1193 1332 1205 1366
rect 1239 1332 1251 1366
rect 1193 1298 1251 1332
rect 1193 1264 1205 1298
rect 1239 1264 1251 1298
rect 1193 1230 1251 1264
rect 1193 1196 1205 1230
rect 1239 1196 1251 1230
rect 1193 1162 1251 1196
rect 1193 1128 1205 1162
rect 1239 1128 1251 1162
rect 1193 1004 1251 1128
rect 1281 1366 1339 1404
rect 1281 1332 1293 1366
rect 1327 1332 1339 1366
rect 1281 1298 1339 1332
rect 1281 1264 1293 1298
rect 1327 1264 1339 1298
rect 1281 1230 1339 1264
rect 1281 1196 1293 1230
rect 1327 1196 1339 1230
rect 1281 1162 1339 1196
rect 1281 1128 1293 1162
rect 1327 1128 1339 1162
rect 1281 1093 1339 1128
rect 1281 1059 1293 1093
rect 1327 1059 1339 1093
rect 1281 1004 1339 1059
rect 1369 1366 1423 1404
rect 1369 1332 1381 1366
rect 1415 1332 1423 1366
rect 1369 1298 1423 1332
rect 1369 1264 1381 1298
rect 1415 1264 1423 1298
rect 1369 1230 1423 1264
rect 1369 1196 1381 1230
rect 1415 1196 1423 1230
rect 1369 1162 1423 1196
rect 1369 1128 1381 1162
rect 1415 1128 1423 1162
rect 1369 1004 1423 1128
rect 1662 1366 1718 1404
rect 1662 1332 1672 1366
rect 1706 1332 1718 1366
rect 1662 1298 1718 1332
rect 1662 1264 1672 1298
rect 1706 1264 1718 1298
rect 1662 1230 1718 1264
rect 1662 1196 1672 1230
rect 1706 1196 1718 1230
rect 1662 1162 1718 1196
rect 1662 1128 1672 1162
rect 1706 1128 1718 1162
rect 1662 1093 1718 1128
rect 1662 1059 1672 1093
rect 1706 1059 1718 1093
rect 1662 1004 1718 1059
rect 1748 1366 1806 1404
rect 1748 1332 1760 1366
rect 1794 1332 1806 1366
rect 1748 1298 1806 1332
rect 1748 1264 1760 1298
rect 1794 1264 1806 1298
rect 1748 1230 1806 1264
rect 1748 1196 1760 1230
rect 1794 1196 1806 1230
rect 1748 1162 1806 1196
rect 1748 1128 1760 1162
rect 1794 1128 1806 1162
rect 1748 1093 1806 1128
rect 1748 1059 1760 1093
rect 1794 1059 1806 1093
rect 1748 1004 1806 1059
rect 1836 1366 1890 1404
rect 1836 1332 1848 1366
rect 1882 1332 1890 1366
rect 1836 1298 1890 1332
rect 1836 1264 1848 1298
rect 1882 1264 1890 1298
rect 1836 1230 1890 1264
rect 1836 1196 1848 1230
rect 1882 1196 1890 1230
rect 1836 1162 1890 1196
rect 1836 1128 1848 1162
rect 1882 1128 1890 1162
rect 1836 1093 1890 1128
rect 1836 1059 1848 1093
rect 1882 1059 1890 1093
rect 1836 1004 1890 1059
rect 2129 1366 2185 1404
rect 2129 1332 2139 1366
rect 2173 1332 2185 1366
rect 2129 1298 2185 1332
rect 2129 1264 2139 1298
rect 2173 1264 2185 1298
rect 2129 1230 2185 1264
rect 2129 1196 2139 1230
rect 2173 1196 2185 1230
rect 2129 1162 2185 1196
rect 2129 1128 2139 1162
rect 2173 1128 2185 1162
rect 2129 1093 2185 1128
rect 2129 1059 2139 1093
rect 2173 1059 2185 1093
rect 2129 1004 2185 1059
rect 2215 1366 2273 1404
rect 2215 1332 2227 1366
rect 2261 1332 2273 1366
rect 2215 1298 2273 1332
rect 2215 1264 2227 1298
rect 2261 1264 2273 1298
rect 2215 1230 2273 1264
rect 2215 1196 2227 1230
rect 2261 1196 2273 1230
rect 2215 1162 2273 1196
rect 2215 1128 2227 1162
rect 2261 1128 2273 1162
rect 2215 1093 2273 1128
rect 2215 1059 2227 1093
rect 2261 1059 2273 1093
rect 2215 1004 2273 1059
rect 2303 1366 2361 1404
rect 2303 1332 2315 1366
rect 2349 1332 2361 1366
rect 2303 1298 2361 1332
rect 2303 1264 2315 1298
rect 2349 1264 2361 1298
rect 2303 1230 2361 1264
rect 2303 1196 2315 1230
rect 2349 1196 2361 1230
rect 2303 1162 2361 1196
rect 2303 1128 2315 1162
rect 2349 1128 2361 1162
rect 2303 1004 2361 1128
rect 2391 1366 2449 1404
rect 2391 1332 2403 1366
rect 2437 1332 2449 1366
rect 2391 1298 2449 1332
rect 2391 1264 2403 1298
rect 2437 1264 2449 1298
rect 2391 1230 2449 1264
rect 2391 1196 2403 1230
rect 2437 1196 2449 1230
rect 2391 1162 2449 1196
rect 2391 1128 2403 1162
rect 2437 1128 2449 1162
rect 2391 1093 2449 1128
rect 2391 1059 2403 1093
rect 2437 1059 2449 1093
rect 2391 1004 2449 1059
rect 2479 1366 2533 1404
rect 2479 1332 2491 1366
rect 2525 1332 2533 1366
rect 2479 1298 2533 1332
rect 2479 1264 2491 1298
rect 2525 1264 2533 1298
rect 2479 1230 2533 1264
rect 2479 1196 2491 1230
rect 2525 1196 2533 1230
rect 2479 1162 2533 1196
rect 2479 1128 2491 1162
rect 2525 1128 2533 1162
rect 2479 1004 2533 1128
rect 2772 1366 2828 1404
rect 2772 1332 2782 1366
rect 2816 1332 2828 1366
rect 2772 1298 2828 1332
rect 2772 1264 2782 1298
rect 2816 1264 2828 1298
rect 2772 1230 2828 1264
rect 2772 1196 2782 1230
rect 2816 1196 2828 1230
rect 2772 1162 2828 1196
rect 2772 1128 2782 1162
rect 2816 1128 2828 1162
rect 2772 1093 2828 1128
rect 2772 1059 2782 1093
rect 2816 1059 2828 1093
rect 2772 1004 2828 1059
rect 2858 1366 2916 1404
rect 2858 1332 2870 1366
rect 2904 1332 2916 1366
rect 2858 1298 2916 1332
rect 2858 1264 2870 1298
rect 2904 1264 2916 1298
rect 2858 1230 2916 1264
rect 2858 1196 2870 1230
rect 2904 1196 2916 1230
rect 2858 1162 2916 1196
rect 2858 1128 2870 1162
rect 2904 1128 2916 1162
rect 2858 1093 2916 1128
rect 2858 1059 2870 1093
rect 2904 1059 2916 1093
rect 2858 1004 2916 1059
rect 2946 1366 3000 1404
rect 2946 1332 2958 1366
rect 2992 1332 3000 1366
rect 2946 1298 3000 1332
rect 2946 1264 2958 1298
rect 2992 1264 3000 1298
rect 2946 1230 3000 1264
rect 2946 1196 2958 1230
rect 2992 1196 3000 1230
rect 2946 1162 3000 1196
rect 2946 1128 2958 1162
rect 2992 1128 3000 1162
rect 2946 1093 3000 1128
rect 2946 1059 2958 1093
rect 2992 1059 3000 1093
rect 2946 1004 3000 1059
rect 3239 1365 3295 1405
rect 3239 1331 3249 1365
rect 3283 1331 3295 1365
rect 3239 1297 3295 1331
rect 3239 1263 3249 1297
rect 3283 1263 3295 1297
rect 3239 1229 3295 1263
rect 3239 1195 3249 1229
rect 3283 1195 3295 1229
rect 3239 1161 3295 1195
rect 3239 1127 3249 1161
rect 3283 1127 3295 1161
rect 3239 1093 3295 1127
rect 3239 1059 3249 1093
rect 3283 1059 3295 1093
rect 3239 1005 3295 1059
rect 3325 1365 3383 1405
rect 3325 1331 3337 1365
rect 3371 1331 3383 1365
rect 3325 1297 3383 1331
rect 3325 1263 3337 1297
rect 3371 1263 3383 1297
rect 3325 1229 3383 1263
rect 3325 1195 3337 1229
rect 3371 1195 3383 1229
rect 3325 1161 3383 1195
rect 3325 1127 3337 1161
rect 3371 1127 3383 1161
rect 3325 1005 3383 1127
rect 3413 1365 3471 1405
rect 3413 1331 3425 1365
rect 3459 1331 3471 1365
rect 3413 1297 3471 1331
rect 3413 1263 3425 1297
rect 3459 1263 3471 1297
rect 3413 1229 3471 1263
rect 3413 1195 3425 1229
rect 3459 1195 3471 1229
rect 3413 1161 3471 1195
rect 3413 1127 3425 1161
rect 3459 1127 3471 1161
rect 3413 1093 3471 1127
rect 3413 1059 3425 1093
rect 3459 1059 3471 1093
rect 3413 1005 3471 1059
rect 3501 1297 3559 1405
rect 3501 1263 3513 1297
rect 3547 1263 3559 1297
rect 3501 1229 3559 1263
rect 3501 1195 3513 1229
rect 3547 1195 3559 1229
rect 3501 1161 3559 1195
rect 3501 1127 3513 1161
rect 3547 1127 3559 1161
rect 3501 1093 3559 1127
rect 3501 1059 3513 1093
rect 3547 1059 3559 1093
rect 3501 1005 3559 1059
rect 3589 1365 3643 1405
rect 3589 1331 3601 1365
rect 3635 1331 3643 1365
rect 3589 1297 3643 1331
rect 3589 1263 3601 1297
rect 3635 1263 3643 1297
rect 3589 1229 3643 1263
rect 3589 1195 3601 1229
rect 3635 1195 3643 1229
rect 3589 1161 3643 1195
rect 3589 1127 3601 1161
rect 3635 1127 3643 1161
rect 3589 1005 3643 1127
rect 3905 1365 3961 1405
rect 3905 1331 3915 1365
rect 3949 1331 3961 1365
rect 3905 1297 3961 1331
rect 3905 1263 3915 1297
rect 3949 1263 3961 1297
rect 3905 1229 3961 1263
rect 3905 1195 3915 1229
rect 3949 1195 3961 1229
rect 3905 1161 3961 1195
rect 3905 1127 3915 1161
rect 3949 1127 3961 1161
rect 3905 1093 3961 1127
rect 3905 1059 3915 1093
rect 3949 1059 3961 1093
rect 3905 1005 3961 1059
rect 3991 1365 4049 1405
rect 3991 1331 4003 1365
rect 4037 1331 4049 1365
rect 3991 1297 4049 1331
rect 3991 1263 4003 1297
rect 4037 1263 4049 1297
rect 3991 1229 4049 1263
rect 3991 1195 4003 1229
rect 4037 1195 4049 1229
rect 3991 1161 4049 1195
rect 3991 1127 4003 1161
rect 4037 1127 4049 1161
rect 3991 1005 4049 1127
rect 4079 1365 4137 1405
rect 4079 1331 4091 1365
rect 4125 1331 4137 1365
rect 4079 1297 4137 1331
rect 4079 1263 4091 1297
rect 4125 1263 4137 1297
rect 4079 1229 4137 1263
rect 4079 1195 4091 1229
rect 4125 1195 4137 1229
rect 4079 1161 4137 1195
rect 4079 1127 4091 1161
rect 4125 1127 4137 1161
rect 4079 1093 4137 1127
rect 4079 1059 4091 1093
rect 4125 1059 4137 1093
rect 4079 1005 4137 1059
rect 4167 1297 4225 1405
rect 4167 1263 4179 1297
rect 4213 1263 4225 1297
rect 4167 1229 4225 1263
rect 4167 1195 4179 1229
rect 4213 1195 4225 1229
rect 4167 1161 4225 1195
rect 4167 1127 4179 1161
rect 4213 1127 4225 1161
rect 4167 1093 4225 1127
rect 4167 1059 4179 1093
rect 4213 1059 4225 1093
rect 4167 1005 4225 1059
rect 4255 1365 4309 1405
rect 4255 1331 4267 1365
rect 4301 1331 4309 1365
rect 4255 1297 4309 1331
rect 4255 1263 4267 1297
rect 4301 1263 4309 1297
rect 4255 1229 4309 1263
rect 4255 1195 4267 1229
rect 4301 1195 4309 1229
rect 4255 1161 4309 1195
rect 4255 1127 4267 1161
rect 4301 1127 4309 1161
rect 4255 1005 4309 1127
<< ndiffc >>
rect 109 300 143 334
rect 303 300 337 334
rect 109 228 143 262
rect 109 160 143 194
rect 205 184 239 218
rect 303 228 337 262
rect 303 160 337 194
rect 109 90 143 124
rect 205 90 239 124
rect 303 90 337 124
rect 553 300 587 334
rect 747 300 781 334
rect 553 228 587 262
rect 553 160 587 194
rect 649 184 683 218
rect 747 228 781 262
rect 747 160 781 194
rect 553 90 587 124
rect 649 90 683 124
rect 747 90 781 124
rect 1010 299 1044 333
rect 1107 299 1141 333
rect 1204 299 1238 333
rect 1010 227 1044 261
rect 1010 159 1044 193
rect 1107 174 1141 208
rect 1204 227 1238 261
rect 1204 159 1238 193
rect 1301 183 1335 217
rect 1398 227 1432 261
rect 1398 159 1432 193
rect 1010 89 1044 123
rect 1204 89 1238 123
rect 1301 89 1335 123
rect 1398 89 1432 123
rect 1663 300 1697 334
rect 1857 300 1891 334
rect 1663 228 1697 262
rect 1663 160 1697 194
rect 1759 184 1793 218
rect 1857 228 1891 262
rect 1857 160 1891 194
rect 1663 90 1697 124
rect 1759 90 1793 124
rect 1857 90 1891 124
rect 2120 299 2154 333
rect 2217 299 2251 333
rect 2314 299 2348 333
rect 2120 227 2154 261
rect 2120 159 2154 193
rect 2217 174 2251 208
rect 2314 227 2348 261
rect 2314 159 2348 193
rect 2411 183 2445 217
rect 2508 227 2542 261
rect 2508 159 2542 193
rect 2120 89 2154 123
rect 2314 89 2348 123
rect 2411 89 2445 123
rect 2508 89 2542 123
rect 2773 300 2807 334
rect 2967 300 3001 334
rect 2773 228 2807 262
rect 2773 160 2807 194
rect 2869 184 2903 218
rect 2967 228 3001 262
rect 2967 160 3001 194
rect 2773 90 2807 124
rect 2869 90 2903 124
rect 2967 90 3001 124
rect 3230 299 3264 333
rect 3230 227 3264 261
rect 3230 159 3264 193
rect 3327 183 3361 217
rect 3424 227 3458 261
rect 3424 159 3458 193
rect 3521 183 3555 217
rect 3618 227 3652 261
rect 3618 159 3652 193
rect 3230 89 3264 123
rect 3327 89 3361 123
rect 3424 89 3458 123
rect 3521 89 3555 123
rect 3618 89 3652 123
rect 3896 299 3930 333
rect 3896 227 3930 261
rect 3896 159 3930 193
rect 3993 183 4027 217
rect 4090 227 4124 261
rect 4090 159 4124 193
rect 4187 183 4221 217
rect 4284 227 4318 261
rect 4284 159 4318 193
rect 3896 89 3930 123
rect 3993 89 4027 123
rect 4090 89 4124 123
rect 4187 89 4221 123
rect 4284 89 4318 123
<< pdiffc >>
rect 118 1332 152 1366
rect 118 1264 152 1298
rect 118 1196 152 1230
rect 118 1128 152 1162
rect 118 1059 152 1093
rect 206 1332 240 1366
rect 206 1264 240 1298
rect 206 1196 240 1230
rect 206 1128 240 1162
rect 206 1059 240 1093
rect 294 1332 328 1366
rect 294 1264 328 1298
rect 294 1196 328 1230
rect 294 1128 328 1162
rect 294 1059 328 1093
rect 562 1332 596 1366
rect 562 1264 596 1298
rect 562 1196 596 1230
rect 562 1128 596 1162
rect 562 1059 596 1093
rect 650 1332 684 1366
rect 650 1264 684 1298
rect 650 1196 684 1230
rect 650 1128 684 1162
rect 650 1059 684 1093
rect 738 1332 772 1366
rect 738 1264 772 1298
rect 738 1196 772 1230
rect 738 1128 772 1162
rect 738 1059 772 1093
rect 1029 1332 1063 1366
rect 1029 1264 1063 1298
rect 1029 1196 1063 1230
rect 1029 1128 1063 1162
rect 1029 1059 1063 1093
rect 1117 1332 1151 1366
rect 1117 1264 1151 1298
rect 1117 1196 1151 1230
rect 1117 1128 1151 1162
rect 1117 1059 1151 1093
rect 1205 1332 1239 1366
rect 1205 1264 1239 1298
rect 1205 1196 1239 1230
rect 1205 1128 1239 1162
rect 1293 1332 1327 1366
rect 1293 1264 1327 1298
rect 1293 1196 1327 1230
rect 1293 1128 1327 1162
rect 1293 1059 1327 1093
rect 1381 1332 1415 1366
rect 1381 1264 1415 1298
rect 1381 1196 1415 1230
rect 1381 1128 1415 1162
rect 1672 1332 1706 1366
rect 1672 1264 1706 1298
rect 1672 1196 1706 1230
rect 1672 1128 1706 1162
rect 1672 1059 1706 1093
rect 1760 1332 1794 1366
rect 1760 1264 1794 1298
rect 1760 1196 1794 1230
rect 1760 1128 1794 1162
rect 1760 1059 1794 1093
rect 1848 1332 1882 1366
rect 1848 1264 1882 1298
rect 1848 1196 1882 1230
rect 1848 1128 1882 1162
rect 1848 1059 1882 1093
rect 2139 1332 2173 1366
rect 2139 1264 2173 1298
rect 2139 1196 2173 1230
rect 2139 1128 2173 1162
rect 2139 1059 2173 1093
rect 2227 1332 2261 1366
rect 2227 1264 2261 1298
rect 2227 1196 2261 1230
rect 2227 1128 2261 1162
rect 2227 1059 2261 1093
rect 2315 1332 2349 1366
rect 2315 1264 2349 1298
rect 2315 1196 2349 1230
rect 2315 1128 2349 1162
rect 2403 1332 2437 1366
rect 2403 1264 2437 1298
rect 2403 1196 2437 1230
rect 2403 1128 2437 1162
rect 2403 1059 2437 1093
rect 2491 1332 2525 1366
rect 2491 1264 2525 1298
rect 2491 1196 2525 1230
rect 2491 1128 2525 1162
rect 2782 1332 2816 1366
rect 2782 1264 2816 1298
rect 2782 1196 2816 1230
rect 2782 1128 2816 1162
rect 2782 1059 2816 1093
rect 2870 1332 2904 1366
rect 2870 1264 2904 1298
rect 2870 1196 2904 1230
rect 2870 1128 2904 1162
rect 2870 1059 2904 1093
rect 2958 1332 2992 1366
rect 2958 1264 2992 1298
rect 2958 1196 2992 1230
rect 2958 1128 2992 1162
rect 2958 1059 2992 1093
rect 3249 1331 3283 1365
rect 3249 1263 3283 1297
rect 3249 1195 3283 1229
rect 3249 1127 3283 1161
rect 3249 1059 3283 1093
rect 3337 1331 3371 1365
rect 3337 1263 3371 1297
rect 3337 1195 3371 1229
rect 3337 1127 3371 1161
rect 3425 1331 3459 1365
rect 3425 1263 3459 1297
rect 3425 1195 3459 1229
rect 3425 1127 3459 1161
rect 3425 1059 3459 1093
rect 3513 1263 3547 1297
rect 3513 1195 3547 1229
rect 3513 1127 3547 1161
rect 3513 1059 3547 1093
rect 3601 1331 3635 1365
rect 3601 1263 3635 1297
rect 3601 1195 3635 1229
rect 3601 1127 3635 1161
rect 3915 1331 3949 1365
rect 3915 1263 3949 1297
rect 3915 1195 3949 1229
rect 3915 1127 3949 1161
rect 3915 1059 3949 1093
rect 4003 1331 4037 1365
rect 4003 1263 4037 1297
rect 4003 1195 4037 1229
rect 4003 1127 4037 1161
rect 4091 1331 4125 1365
rect 4091 1263 4125 1297
rect 4091 1195 4125 1229
rect 4091 1127 4125 1161
rect 4091 1059 4125 1093
rect 4179 1263 4213 1297
rect 4179 1195 4213 1229
rect 4179 1127 4213 1161
rect 4179 1059 4213 1093
rect 4267 1331 4301 1365
rect 4267 1263 4301 1297
rect 4267 1195 4301 1229
rect 4267 1127 4301 1161
<< psubdiff >>
rect -34 482 4474 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 410 461 478 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 410 427 427 461
rect 461 427 478 461
rect 854 461 922 482
rect -34 313 34 353
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect 854 427 871 461
rect 905 427 922 461
rect 1520 461 1588 482
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 410 313 478 353
rect 854 387 922 427
rect 854 353 871 387
rect 905 353 922 387
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect -34 17 34 57
rect 410 57 427 91
rect 461 57 478 91
rect 854 313 922 353
rect 1520 427 1537 461
rect 1571 427 1588 461
rect 1964 461 2032 482
rect 1520 387 1588 427
rect 1520 353 1537 387
rect 1571 353 1588 387
rect 1964 427 1981 461
rect 2015 427 2032 461
rect 2630 461 2698 482
rect 854 279 871 313
rect 905 279 922 313
rect 854 239 922 279
rect 854 205 871 239
rect 905 205 922 239
rect 854 165 922 205
rect 854 131 871 165
rect 905 131 922 165
rect 854 91 922 131
rect 410 17 478 57
rect 854 57 871 91
rect 905 57 922 91
rect 1520 313 1588 353
rect 1964 387 2032 427
rect 1964 353 1981 387
rect 2015 353 2032 387
rect 1520 279 1537 313
rect 1571 279 1588 313
rect 1520 239 1588 279
rect 1520 205 1537 239
rect 1571 205 1588 239
rect 1520 165 1588 205
rect 1520 131 1537 165
rect 1571 131 1588 165
rect 1520 91 1588 131
rect 854 17 922 57
rect 1520 57 1537 91
rect 1571 57 1588 91
rect 1964 313 2032 353
rect 2630 427 2647 461
rect 2681 427 2698 461
rect 3074 461 3142 482
rect 2630 387 2698 427
rect 2630 353 2647 387
rect 2681 353 2698 387
rect 3074 427 3091 461
rect 3125 427 3142 461
rect 3740 461 3808 482
rect 1964 279 1981 313
rect 2015 279 2032 313
rect 1964 239 2032 279
rect 1964 205 1981 239
rect 2015 205 2032 239
rect 1964 165 2032 205
rect 1964 131 1981 165
rect 2015 131 2032 165
rect 1964 91 2032 131
rect 1520 17 1588 57
rect 1964 57 1981 91
rect 2015 57 2032 91
rect 2630 313 2698 353
rect 3074 387 3142 427
rect 3074 353 3091 387
rect 3125 353 3142 387
rect 2630 279 2647 313
rect 2681 279 2698 313
rect 2630 239 2698 279
rect 2630 205 2647 239
rect 2681 205 2698 239
rect 2630 165 2698 205
rect 2630 131 2647 165
rect 2681 131 2698 165
rect 2630 91 2698 131
rect 1964 17 2032 57
rect 2630 57 2647 91
rect 2681 57 2698 91
rect 3074 313 3142 353
rect 3740 427 3757 461
rect 3791 427 3808 461
rect 4406 461 4474 482
rect 3740 387 3808 427
rect 3740 353 3757 387
rect 3791 353 3808 387
rect 3074 279 3091 313
rect 3125 279 3142 313
rect 3074 239 3142 279
rect 3074 205 3091 239
rect 3125 205 3142 239
rect 3074 165 3142 205
rect 3074 131 3091 165
rect 3125 131 3142 165
rect 3074 91 3142 131
rect 2630 17 2698 57
rect 3074 57 3091 91
rect 3125 57 3142 91
rect 3740 313 3808 353
rect 4406 427 4423 461
rect 4457 427 4474 461
rect 4406 387 4474 427
rect 4406 353 4423 387
rect 4457 353 4474 387
rect 3740 279 3757 313
rect 3791 279 3808 313
rect 3740 239 3808 279
rect 3740 205 3757 239
rect 3791 205 3808 239
rect 3740 165 3808 205
rect 3740 131 3757 165
rect 3791 131 3808 165
rect 3740 91 3808 131
rect 3074 17 3142 57
rect 3740 57 3757 91
rect 3791 57 3808 91
rect 4406 313 4474 353
rect 4406 279 4423 313
rect 4457 279 4474 313
rect 4406 239 4474 279
rect 4406 205 4423 239
rect 4457 205 4474 239
rect 4406 165 4474 205
rect 4406 131 4423 165
rect 4457 131 4474 165
rect 4406 91 4474 131
rect 3740 17 3808 57
rect 4406 57 4423 91
rect 4457 57 4474 91
rect 4406 17 4474 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4474 17
rect -34 -34 4474 -17
<< nsubdiff >>
rect -34 1497 4474 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4474 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 410 1423 478 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 854 1423 922 1463
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 410 979 478 1019
rect 854 1389 871 1423
rect 905 1389 922 1423
rect 1520 1423 1588 1463
rect 854 1349 922 1389
rect 854 1315 871 1349
rect 905 1315 922 1349
rect 854 1275 922 1315
rect 854 1241 871 1275
rect 905 1241 922 1275
rect 854 1201 922 1241
rect 854 1167 871 1201
rect 905 1167 922 1201
rect 854 1127 922 1167
rect 854 1093 871 1127
rect 905 1093 922 1127
rect 854 1053 922 1093
rect 854 1019 871 1053
rect 905 1019 922 1053
rect 410 945 427 979
rect 461 945 478 979
rect -34 871 -17 905
rect 17 884 34 905
rect 410 905 478 945
rect 854 979 922 1019
rect 1520 1389 1537 1423
rect 1571 1389 1588 1423
rect 1964 1423 2032 1463
rect 1520 1349 1588 1389
rect 1520 1315 1537 1349
rect 1571 1315 1588 1349
rect 1520 1275 1588 1315
rect 1520 1241 1537 1275
rect 1571 1241 1588 1275
rect 1520 1201 1588 1241
rect 1520 1167 1537 1201
rect 1571 1167 1588 1201
rect 1520 1127 1588 1167
rect 1520 1093 1537 1127
rect 1571 1093 1588 1127
rect 1520 1053 1588 1093
rect 1520 1019 1537 1053
rect 1571 1019 1588 1053
rect 854 945 871 979
rect 905 945 922 979
rect 410 884 427 905
rect 17 871 427 884
rect 461 884 478 905
rect 854 905 922 945
rect 1520 979 1588 1019
rect 1964 1389 1981 1423
rect 2015 1389 2032 1423
rect 2630 1423 2698 1463
rect 1964 1349 2032 1389
rect 1964 1315 1981 1349
rect 2015 1315 2032 1349
rect 1964 1275 2032 1315
rect 1964 1241 1981 1275
rect 2015 1241 2032 1275
rect 1964 1201 2032 1241
rect 1964 1167 1981 1201
rect 2015 1167 2032 1201
rect 1964 1127 2032 1167
rect 1964 1093 1981 1127
rect 2015 1093 2032 1127
rect 1964 1053 2032 1093
rect 1964 1019 1981 1053
rect 2015 1019 2032 1053
rect 1520 945 1537 979
rect 1571 945 1588 979
rect 854 884 871 905
rect 461 871 871 884
rect 905 884 922 905
rect 1520 905 1588 945
rect 1964 979 2032 1019
rect 2630 1389 2647 1423
rect 2681 1389 2698 1423
rect 3074 1423 3142 1463
rect 2630 1349 2698 1389
rect 2630 1315 2647 1349
rect 2681 1315 2698 1349
rect 2630 1275 2698 1315
rect 2630 1241 2647 1275
rect 2681 1241 2698 1275
rect 2630 1201 2698 1241
rect 2630 1167 2647 1201
rect 2681 1167 2698 1201
rect 2630 1127 2698 1167
rect 2630 1093 2647 1127
rect 2681 1093 2698 1127
rect 2630 1053 2698 1093
rect 2630 1019 2647 1053
rect 2681 1019 2698 1053
rect 1964 945 1981 979
rect 2015 945 2032 979
rect 1520 884 1537 905
rect 905 871 1537 884
rect 1571 884 1588 905
rect 1964 905 2032 945
rect 2630 979 2698 1019
rect 3074 1389 3091 1423
rect 3125 1389 3142 1423
rect 3740 1423 3808 1463
rect 3074 1349 3142 1389
rect 3074 1315 3091 1349
rect 3125 1315 3142 1349
rect 3074 1275 3142 1315
rect 3074 1241 3091 1275
rect 3125 1241 3142 1275
rect 3074 1201 3142 1241
rect 3074 1167 3091 1201
rect 3125 1167 3142 1201
rect 3074 1127 3142 1167
rect 3074 1093 3091 1127
rect 3125 1093 3142 1127
rect 3074 1053 3142 1093
rect 3074 1019 3091 1053
rect 3125 1019 3142 1053
rect 2630 945 2647 979
rect 2681 945 2698 979
rect 1964 884 1981 905
rect 1571 871 1981 884
rect 2015 884 2032 905
rect 2630 905 2698 945
rect 3074 979 3142 1019
rect 3740 1389 3757 1423
rect 3791 1389 3808 1423
rect 4406 1423 4474 1463
rect 3740 1349 3808 1389
rect 3740 1315 3757 1349
rect 3791 1315 3808 1349
rect 3740 1275 3808 1315
rect 3740 1241 3757 1275
rect 3791 1241 3808 1275
rect 3740 1201 3808 1241
rect 3740 1167 3757 1201
rect 3791 1167 3808 1201
rect 3740 1127 3808 1167
rect 3740 1093 3757 1127
rect 3791 1093 3808 1127
rect 3740 1053 3808 1093
rect 3740 1019 3757 1053
rect 3791 1019 3808 1053
rect 3074 945 3091 979
rect 3125 945 3142 979
rect 2630 884 2647 905
rect 2015 871 2647 884
rect 2681 884 2698 905
rect 3074 905 3142 945
rect 3740 979 3808 1019
rect 4406 1389 4423 1423
rect 4457 1389 4474 1423
rect 4406 1349 4474 1389
rect 4406 1315 4423 1349
rect 4457 1315 4474 1349
rect 4406 1275 4474 1315
rect 4406 1241 4423 1275
rect 4457 1241 4474 1275
rect 4406 1201 4474 1241
rect 4406 1167 4423 1201
rect 4457 1167 4474 1201
rect 4406 1127 4474 1167
rect 4406 1093 4423 1127
rect 4457 1093 4474 1127
rect 4406 1053 4474 1093
rect 4406 1019 4423 1053
rect 4457 1019 4474 1053
rect 3740 945 3757 979
rect 3791 945 3808 979
rect 3074 884 3091 905
rect 2681 871 3091 884
rect 3125 884 3142 905
rect 3740 905 3808 945
rect 4406 979 4474 1019
rect 4406 945 4423 979
rect 4457 945 4474 979
rect 3740 884 3757 905
rect 3125 871 3757 884
rect 3791 884 3808 905
rect 4406 905 4474 945
rect 4406 884 4423 905
rect 3791 871 4423 884
rect 4457 871 4474 905
rect -34 822 4474 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 427 427 461 461
rect 427 353 461 387
rect 871 427 905 461
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 871 353 905 387
rect 427 279 461 313
rect 427 205 461 239
rect 427 131 461 165
rect 427 57 461 91
rect 1537 427 1571 461
rect 1537 353 1571 387
rect 1981 427 2015 461
rect 871 279 905 313
rect 871 205 905 239
rect 871 131 905 165
rect 871 57 905 91
rect 1981 353 2015 387
rect 1537 279 1571 313
rect 1537 205 1571 239
rect 1537 131 1571 165
rect 1537 57 1571 91
rect 2647 427 2681 461
rect 2647 353 2681 387
rect 3091 427 3125 461
rect 1981 279 2015 313
rect 1981 205 2015 239
rect 1981 131 2015 165
rect 1981 57 2015 91
rect 3091 353 3125 387
rect 2647 279 2681 313
rect 2647 205 2681 239
rect 2647 131 2681 165
rect 2647 57 2681 91
rect 3757 427 3791 461
rect 3757 353 3791 387
rect 3091 279 3125 313
rect 3091 205 3125 239
rect 3091 131 3125 165
rect 3091 57 3125 91
rect 4423 427 4457 461
rect 4423 353 4457 387
rect 3757 279 3791 313
rect 3757 205 3791 239
rect 3757 131 3791 165
rect 3757 57 3791 91
rect 4423 279 4457 313
rect 4423 205 4457 239
rect 4423 131 4457 165
rect 4423 57 4457 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 427 1389 461 1423
rect 427 1315 461 1349
rect 427 1241 461 1275
rect 427 1167 461 1201
rect 427 1093 461 1127
rect 427 1019 461 1053
rect -17 945 17 979
rect 871 1389 905 1423
rect 871 1315 905 1349
rect 871 1241 905 1275
rect 871 1167 905 1201
rect 871 1093 905 1127
rect 871 1019 905 1053
rect 427 945 461 979
rect -17 871 17 905
rect 1537 1389 1571 1423
rect 1537 1315 1571 1349
rect 1537 1241 1571 1275
rect 1537 1167 1571 1201
rect 1537 1093 1571 1127
rect 1537 1019 1571 1053
rect 871 945 905 979
rect 427 871 461 905
rect 1981 1389 2015 1423
rect 1981 1315 2015 1349
rect 1981 1241 2015 1275
rect 1981 1167 2015 1201
rect 1981 1093 2015 1127
rect 1981 1019 2015 1053
rect 1537 945 1571 979
rect 871 871 905 905
rect 2647 1389 2681 1423
rect 2647 1315 2681 1349
rect 2647 1241 2681 1275
rect 2647 1167 2681 1201
rect 2647 1093 2681 1127
rect 2647 1019 2681 1053
rect 1981 945 2015 979
rect 1537 871 1571 905
rect 3091 1389 3125 1423
rect 3091 1315 3125 1349
rect 3091 1241 3125 1275
rect 3091 1167 3125 1201
rect 3091 1093 3125 1127
rect 3091 1019 3125 1053
rect 2647 945 2681 979
rect 1981 871 2015 905
rect 3757 1389 3791 1423
rect 3757 1315 3791 1349
rect 3757 1241 3791 1275
rect 3757 1167 3791 1201
rect 3757 1093 3791 1127
rect 3757 1019 3791 1053
rect 3091 945 3125 979
rect 2647 871 2681 905
rect 4423 1389 4457 1423
rect 4423 1315 4457 1349
rect 4423 1241 4457 1275
rect 4423 1167 4457 1201
rect 4423 1093 4457 1127
rect 4423 1019 4457 1053
rect 3757 945 3791 979
rect 3091 871 3125 905
rect 4423 945 4457 979
rect 3757 871 3791 905
rect 4423 871 4457 905
<< poly >>
rect 164 1404 194 1430
rect 252 1404 282 1430
rect 608 1404 638 1430
rect 696 1404 726 1430
rect 164 973 194 1004
rect 252 973 282 1004
rect 121 957 282 973
rect 121 923 131 957
rect 165 943 282 957
rect 1075 1404 1105 1430
rect 1163 1404 1193 1430
rect 1251 1404 1281 1430
rect 1339 1404 1369 1430
rect 608 973 638 1004
rect 696 973 726 1004
rect 165 923 175 943
rect 121 907 175 923
rect 565 957 726 973
rect 565 923 575 957
rect 609 943 726 957
rect 1718 1404 1748 1430
rect 1806 1404 1836 1430
rect 609 923 619 943
rect 565 907 619 923
rect 1075 973 1105 1004
rect 1163 973 1193 1004
rect 1251 973 1281 1004
rect 1339 973 1369 1004
rect 1075 957 1193 973
rect 1075 943 1093 957
rect 1083 923 1093 943
rect 1127 943 1193 957
rect 1237 957 1369 973
rect 1127 923 1137 943
rect 1083 907 1137 923
rect 1237 923 1247 957
rect 1281 943 1369 957
rect 2185 1404 2215 1430
rect 2273 1404 2303 1430
rect 2361 1404 2391 1430
rect 2449 1404 2479 1430
rect 1718 973 1748 1004
rect 1806 973 1836 1004
rect 1281 923 1291 943
rect 1237 907 1291 923
rect 1675 957 1836 973
rect 1675 923 1685 957
rect 1719 943 1836 957
rect 2828 1404 2858 1430
rect 2916 1404 2946 1430
rect 1719 923 1729 943
rect 1675 907 1729 923
rect 2185 973 2215 1004
rect 2273 973 2303 1004
rect 2361 973 2391 1004
rect 2449 973 2479 1004
rect 2185 957 2303 973
rect 2185 943 2203 957
rect 2193 923 2203 943
rect 2237 943 2303 957
rect 2347 957 2479 973
rect 2237 923 2247 943
rect 2193 907 2247 923
rect 2347 923 2357 957
rect 2391 943 2479 957
rect 3295 1405 3325 1431
rect 3383 1405 3413 1431
rect 3471 1405 3501 1431
rect 3559 1405 3589 1431
rect 2828 973 2858 1004
rect 2916 973 2946 1004
rect 2391 923 2401 943
rect 2347 907 2401 923
rect 2785 957 2946 973
rect 2785 923 2795 957
rect 2829 943 2946 957
rect 3961 1405 3991 1431
rect 4049 1405 4079 1431
rect 4137 1405 4167 1431
rect 4225 1405 4255 1431
rect 3295 974 3325 1005
rect 3383 974 3413 1005
rect 3471 974 3501 1005
rect 3559 974 3589 1005
rect 2829 923 2839 943
rect 2785 907 2839 923
rect 3272 958 3413 974
rect 3272 924 3282 958
rect 3316 944 3413 958
rect 3458 958 3589 974
rect 3316 924 3326 944
rect 3272 908 3326 924
rect 3458 924 3468 958
rect 3502 944 3589 958
rect 3961 974 3991 1005
rect 4049 974 4079 1005
rect 4137 974 4167 1005
rect 4225 974 4255 1005
rect 3502 924 3512 944
rect 3458 908 3512 924
rect 3938 958 4079 974
rect 3938 924 3948 958
rect 3982 944 4079 958
rect 4124 958 4255 974
rect 3982 924 3992 944
rect 3938 908 3992 924
rect 4124 924 4134 958
rect 4168 944 4255 958
rect 4168 924 4178 944
rect 4124 908 4178 924
rect 121 434 175 450
rect 121 400 131 434
rect 165 413 175 434
rect 165 400 185 413
rect 121 384 185 400
rect 155 350 185 384
rect 565 434 619 450
rect 565 400 575 434
rect 609 413 619 434
rect 609 400 629 413
rect 565 384 629 400
rect 599 350 629 384
rect 1083 433 1137 449
rect 1083 413 1093 433
rect 1056 399 1093 413
rect 1127 399 1137 433
rect 1056 383 1137 399
rect 1231 433 1285 449
rect 1231 399 1241 433
rect 1275 399 1285 433
rect 1231 383 1285 399
rect 1056 349 1086 383
rect 1250 349 1280 383
rect 1675 434 1729 450
rect 1675 400 1685 434
rect 1719 413 1729 434
rect 1719 400 1739 413
rect 1675 384 1739 400
rect 1709 350 1739 384
rect 2193 433 2247 449
rect 2193 413 2203 433
rect 2166 399 2203 413
rect 2237 399 2247 433
rect 2166 383 2247 399
rect 2341 433 2395 449
rect 2341 399 2351 433
rect 2385 399 2395 433
rect 2341 383 2395 399
rect 2166 349 2196 383
rect 2360 349 2390 383
rect 2785 434 2839 450
rect 2785 400 2795 434
rect 2829 413 2839 434
rect 2829 400 2849 413
rect 2785 384 2849 400
rect 2819 350 2849 384
rect 3303 433 3357 449
rect 3303 413 3313 433
rect 3276 399 3313 413
rect 3347 399 3357 433
rect 3276 383 3357 399
rect 3451 433 3505 449
rect 3451 399 3461 433
rect 3495 399 3505 433
rect 3451 383 3505 399
rect 3969 433 4023 449
rect 3969 413 3979 433
rect 3276 349 3306 383
rect 3470 349 3500 383
rect 3942 399 3979 413
rect 4013 399 4023 433
rect 3942 383 4023 399
rect 4117 433 4171 449
rect 4117 399 4127 433
rect 4161 399 4171 433
rect 4117 383 4171 399
rect 3942 349 3972 383
rect 4136 349 4166 383
<< polycont >>
rect 131 923 165 957
rect 575 923 609 957
rect 1093 923 1127 957
rect 1247 923 1281 957
rect 1685 923 1719 957
rect 2203 923 2237 957
rect 2357 923 2391 957
rect 2795 923 2829 957
rect 3282 924 3316 958
rect 3468 924 3502 958
rect 3948 924 3982 958
rect 4134 924 4168 958
rect 131 400 165 434
rect 575 400 609 434
rect 1093 399 1127 433
rect 1241 399 1275 433
rect 1685 400 1719 434
rect 2203 399 2237 433
rect 2351 399 2385 433
rect 2795 400 2829 434
rect 3313 399 3347 433
rect 3461 399 3495 433
rect 3979 399 4013 433
rect 4127 399 4161 433
<< locali >>
rect -34 1497 4474 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4474 1497
rect -34 1446 4474 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 118 1366 152 1446
rect 118 1298 152 1332
rect 118 1230 152 1264
rect 118 1162 152 1196
rect 118 1093 152 1128
rect 118 1037 152 1059
rect 206 1366 240 1404
rect 206 1298 240 1332
rect 206 1230 240 1264
rect 206 1162 240 1196
rect 206 1093 240 1128
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 131 957 165 973
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 131 434 165 923
rect 206 933 240 1059
rect 294 1366 328 1446
rect 294 1298 328 1332
rect 294 1230 328 1264
rect 294 1162 328 1196
rect 294 1093 328 1128
rect 294 1037 328 1059
rect 410 1423 478 1446
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect 562 1366 596 1446
rect 562 1298 596 1332
rect 562 1230 596 1264
rect 562 1162 596 1196
rect 562 1093 596 1128
rect 562 1037 596 1059
rect 650 1366 684 1404
rect 650 1298 684 1332
rect 650 1230 684 1264
rect 650 1162 684 1196
rect 650 1093 684 1128
rect 410 979 478 1019
rect 410 945 427 979
rect 461 945 478 979
rect 206 899 313 933
rect 279 609 313 899
rect 410 905 478 945
rect 410 871 427 905
rect 461 871 478 905
rect 410 822 478 871
rect 575 957 609 973
rect 575 831 609 923
rect 650 933 684 1059
rect 738 1366 772 1446
rect 738 1298 772 1332
rect 738 1230 772 1264
rect 738 1162 772 1196
rect 738 1093 772 1128
rect 738 1037 772 1059
rect 854 1423 922 1446
rect 854 1389 871 1423
rect 905 1389 922 1423
rect 854 1349 922 1389
rect 854 1315 871 1349
rect 905 1315 922 1349
rect 854 1275 922 1315
rect 854 1241 871 1275
rect 905 1241 922 1275
rect 854 1201 922 1241
rect 854 1167 871 1201
rect 905 1167 922 1201
rect 854 1127 922 1167
rect 854 1093 871 1127
rect 905 1093 922 1127
rect 854 1053 922 1093
rect 854 1019 871 1053
rect 905 1019 922 1053
rect 1029 1366 1063 1446
rect 1029 1298 1063 1332
rect 1029 1230 1063 1264
rect 1029 1162 1063 1196
rect 1029 1093 1063 1128
rect 1029 1027 1063 1059
rect 1117 1366 1151 1404
rect 1117 1298 1151 1332
rect 1117 1230 1151 1264
rect 1117 1162 1151 1196
rect 1117 1093 1151 1128
rect 1205 1366 1239 1446
rect 1205 1298 1239 1332
rect 1205 1230 1239 1264
rect 1205 1162 1239 1196
rect 1205 1111 1239 1128
rect 1293 1366 1327 1404
rect 1293 1298 1327 1332
rect 1293 1230 1327 1264
rect 1293 1162 1327 1196
rect 1117 1057 1151 1059
rect 1293 1093 1327 1128
rect 1381 1366 1415 1446
rect 1381 1298 1415 1332
rect 1381 1230 1415 1264
rect 1381 1162 1415 1196
rect 1381 1111 1415 1128
rect 1520 1423 1588 1446
rect 1520 1389 1537 1423
rect 1571 1389 1588 1423
rect 1520 1349 1588 1389
rect 1520 1315 1537 1349
rect 1571 1315 1588 1349
rect 1520 1275 1588 1315
rect 1520 1241 1537 1275
rect 1571 1241 1588 1275
rect 1520 1201 1588 1241
rect 1520 1167 1537 1201
rect 1571 1167 1588 1201
rect 1520 1127 1588 1167
rect 1293 1057 1327 1059
rect 1520 1093 1537 1127
rect 1571 1093 1588 1127
rect 1117 1023 1423 1057
rect 854 979 922 1019
rect 854 945 871 979
rect 905 945 922 979
rect 650 899 757 933
rect 279 433 313 575
rect 131 384 165 400
rect 205 399 313 433
rect 410 461 478 544
rect 410 427 427 461
rect 461 427 478 461
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 109 334 143 350
rect 109 262 143 300
rect 109 194 143 228
rect 205 218 239 399
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect 575 434 609 797
rect 723 757 757 899
rect 854 905 922 945
rect 854 871 871 905
rect 905 871 922 905
rect 854 822 922 871
rect 1093 957 1127 973
rect 1247 957 1281 973
rect 723 433 757 723
rect 1093 757 1127 923
rect 575 384 609 400
rect 649 399 757 433
rect 854 461 922 544
rect 854 427 871 461
rect 905 427 922 461
rect 205 168 239 184
rect 303 334 337 350
rect 303 262 337 300
rect 303 194 337 228
rect 109 124 143 160
rect 303 124 337 160
rect 143 90 205 124
rect 239 90 303 124
rect 109 34 143 90
rect 206 34 240 90
rect 303 34 337 90
rect 410 313 478 353
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect 410 57 427 91
rect 461 57 478 91
rect 410 34 478 57
rect 553 334 587 350
rect 553 262 587 300
rect 553 194 587 228
rect 649 218 683 399
rect 854 387 922 427
rect 854 353 871 387
rect 905 353 922 387
rect 1093 433 1127 723
rect 1093 383 1127 399
rect 1241 923 1247 942
rect 1241 907 1281 923
rect 1241 609 1275 907
rect 1241 433 1275 575
rect 1241 383 1275 399
rect 1389 683 1423 1023
rect 1520 1053 1588 1093
rect 1520 1019 1537 1053
rect 1571 1019 1588 1053
rect 1672 1366 1706 1446
rect 1672 1298 1706 1332
rect 1672 1230 1706 1264
rect 1672 1162 1706 1196
rect 1672 1093 1706 1128
rect 1672 1037 1706 1059
rect 1760 1366 1794 1404
rect 1760 1298 1794 1332
rect 1760 1230 1794 1264
rect 1760 1162 1794 1196
rect 1760 1093 1794 1128
rect 1520 979 1588 1019
rect 1520 945 1537 979
rect 1571 945 1588 979
rect 1520 905 1588 945
rect 1520 871 1537 905
rect 1571 871 1588 905
rect 1520 822 1588 871
rect 1685 957 1719 973
rect 649 168 683 184
rect 747 334 781 350
rect 747 262 781 300
rect 747 194 781 228
rect 553 124 587 160
rect 747 124 781 160
rect 587 90 649 124
rect 683 90 747 124
rect 553 34 587 90
rect 650 34 684 90
rect 747 34 781 90
rect 854 313 922 353
rect 854 279 871 313
rect 905 279 922 313
rect 854 239 922 279
rect 854 205 871 239
rect 905 205 922 239
rect 854 165 922 205
rect 854 131 871 165
rect 905 131 922 165
rect 854 91 922 131
rect 854 57 871 91
rect 905 57 922 91
rect 1010 333 1044 349
rect 1204 333 1238 349
rect 1389 348 1423 649
rect 1685 683 1719 923
rect 1760 933 1794 1059
rect 1848 1366 1882 1446
rect 1848 1298 1882 1332
rect 1848 1230 1882 1264
rect 1848 1162 1882 1196
rect 1848 1093 1882 1128
rect 1848 1037 1882 1059
rect 1964 1423 2032 1446
rect 1964 1389 1981 1423
rect 2015 1389 2032 1423
rect 1964 1349 2032 1389
rect 1964 1315 1981 1349
rect 2015 1315 2032 1349
rect 1964 1275 2032 1315
rect 1964 1241 1981 1275
rect 2015 1241 2032 1275
rect 1964 1201 2032 1241
rect 1964 1167 1981 1201
rect 2015 1167 2032 1201
rect 1964 1127 2032 1167
rect 1964 1093 1981 1127
rect 2015 1093 2032 1127
rect 1964 1053 2032 1093
rect 1964 1019 1981 1053
rect 2015 1019 2032 1053
rect 2139 1366 2173 1446
rect 2139 1298 2173 1332
rect 2139 1230 2173 1264
rect 2139 1162 2173 1196
rect 2139 1093 2173 1128
rect 2139 1027 2173 1059
rect 2227 1366 2261 1404
rect 2227 1298 2261 1332
rect 2227 1230 2261 1264
rect 2227 1162 2261 1196
rect 2227 1093 2261 1128
rect 2315 1366 2349 1446
rect 2315 1298 2349 1332
rect 2315 1230 2349 1264
rect 2315 1162 2349 1196
rect 2315 1111 2349 1128
rect 2403 1366 2437 1404
rect 2403 1298 2437 1332
rect 2403 1230 2437 1264
rect 2403 1162 2437 1196
rect 2227 1057 2261 1059
rect 2403 1093 2437 1128
rect 2491 1366 2525 1446
rect 2491 1298 2525 1332
rect 2491 1230 2525 1264
rect 2491 1162 2525 1196
rect 2491 1111 2525 1128
rect 2630 1423 2698 1446
rect 2630 1389 2647 1423
rect 2681 1389 2698 1423
rect 2630 1349 2698 1389
rect 2630 1315 2647 1349
rect 2681 1315 2698 1349
rect 2630 1275 2698 1315
rect 2630 1241 2647 1275
rect 2681 1241 2698 1275
rect 2630 1201 2698 1241
rect 2630 1167 2647 1201
rect 2681 1167 2698 1201
rect 2630 1127 2698 1167
rect 2403 1057 2437 1059
rect 2630 1093 2647 1127
rect 2681 1093 2698 1127
rect 2227 1023 2533 1057
rect 1964 979 2032 1019
rect 1964 945 1981 979
rect 2015 945 2032 979
rect 1760 899 1867 933
rect 1044 299 1107 333
rect 1141 299 1204 333
rect 1010 261 1044 299
rect 1010 193 1044 227
rect 1204 261 1238 299
rect 1010 123 1044 159
rect 1010 73 1044 89
rect 1107 208 1141 224
rect 854 34 922 57
rect 1107 34 1141 174
rect 1204 193 1238 227
rect 1301 314 1423 348
rect 1520 461 1588 544
rect 1520 427 1537 461
rect 1571 427 1588 461
rect 1520 387 1588 427
rect 1520 353 1537 387
rect 1571 353 1588 387
rect 1685 434 1719 649
rect 1833 757 1867 899
rect 1964 905 2032 945
rect 1964 871 1981 905
rect 2015 871 2032 905
rect 1964 822 2032 871
rect 2203 957 2237 973
rect 2357 957 2391 973
rect 1833 433 1867 723
rect 2203 609 2237 923
rect 1685 384 1719 400
rect 1759 399 1867 433
rect 1964 461 2032 544
rect 1964 427 1981 461
rect 2015 427 2032 461
rect 1301 217 1335 314
rect 1520 313 1588 353
rect 1520 279 1537 313
rect 1571 279 1588 313
rect 1301 167 1335 183
rect 1398 261 1432 277
rect 1398 193 1432 227
rect 1204 123 1238 159
rect 1398 123 1432 159
rect 1238 89 1301 123
rect 1335 89 1398 123
rect 1204 73 1238 89
rect 1398 73 1432 89
rect 1520 239 1588 279
rect 1520 205 1537 239
rect 1571 205 1588 239
rect 1520 165 1588 205
rect 1520 131 1537 165
rect 1571 131 1588 165
rect 1520 91 1588 131
rect 1520 57 1537 91
rect 1571 57 1588 91
rect 1520 34 1588 57
rect 1663 334 1697 350
rect 1663 262 1697 300
rect 1663 194 1697 228
rect 1759 218 1793 399
rect 1964 387 2032 427
rect 1964 353 1981 387
rect 2015 353 2032 387
rect 2203 433 2237 575
rect 2203 383 2237 399
rect 2351 923 2357 942
rect 2351 907 2391 923
rect 2351 831 2385 907
rect 2351 433 2385 797
rect 2351 383 2385 399
rect 2499 683 2533 1023
rect 2630 1053 2698 1093
rect 2630 1019 2647 1053
rect 2681 1019 2698 1053
rect 2782 1366 2816 1446
rect 2782 1298 2816 1332
rect 2782 1230 2816 1264
rect 2782 1162 2816 1196
rect 2782 1093 2816 1128
rect 2782 1037 2816 1059
rect 2870 1366 2904 1404
rect 2870 1298 2904 1332
rect 2870 1230 2904 1264
rect 2870 1162 2904 1196
rect 2870 1093 2904 1128
rect 2630 979 2698 1019
rect 2630 945 2647 979
rect 2681 945 2698 979
rect 2630 905 2698 945
rect 2630 871 2647 905
rect 2681 871 2698 905
rect 2630 822 2698 871
rect 2795 957 2829 973
rect 1759 168 1793 184
rect 1857 334 1891 350
rect 1857 262 1891 300
rect 1857 194 1891 228
rect 1663 124 1697 160
rect 1857 124 1891 160
rect 1697 90 1759 124
rect 1793 90 1857 124
rect 1663 34 1697 90
rect 1760 34 1794 90
rect 1857 34 1891 90
rect 1964 313 2032 353
rect 1964 279 1981 313
rect 2015 279 2032 313
rect 1964 239 2032 279
rect 1964 205 1981 239
rect 2015 205 2032 239
rect 1964 165 2032 205
rect 1964 131 1981 165
rect 2015 131 2032 165
rect 1964 91 2032 131
rect 1964 57 1981 91
rect 2015 57 2032 91
rect 2120 333 2154 349
rect 2314 333 2348 349
rect 2499 348 2533 649
rect 2795 683 2829 923
rect 2870 933 2904 1059
rect 2958 1366 2992 1446
rect 2958 1298 2992 1332
rect 2958 1230 2992 1264
rect 2958 1162 2992 1196
rect 2958 1093 2992 1128
rect 2958 1037 2992 1059
rect 3074 1423 3142 1446
rect 3074 1389 3091 1423
rect 3125 1389 3142 1423
rect 3074 1349 3142 1389
rect 3074 1315 3091 1349
rect 3125 1315 3142 1349
rect 3074 1275 3142 1315
rect 3074 1241 3091 1275
rect 3125 1241 3142 1275
rect 3074 1201 3142 1241
rect 3074 1167 3091 1201
rect 3125 1167 3142 1201
rect 3074 1127 3142 1167
rect 3074 1093 3091 1127
rect 3125 1093 3142 1127
rect 3074 1053 3142 1093
rect 3074 1019 3091 1053
rect 3125 1019 3142 1053
rect 3249 1365 3283 1405
rect 3249 1297 3283 1331
rect 3249 1229 3283 1263
rect 3249 1161 3283 1195
rect 3249 1093 3283 1127
rect 3337 1365 3371 1446
rect 3740 1423 3808 1446
rect 3337 1297 3371 1331
rect 3337 1229 3371 1263
rect 3337 1161 3371 1195
rect 3337 1111 3371 1127
rect 3425 1365 3635 1399
rect 3425 1297 3459 1331
rect 3425 1229 3459 1263
rect 3425 1161 3459 1195
rect 3425 1093 3459 1127
rect 3249 1025 3459 1059
rect 3513 1297 3547 1313
rect 3513 1229 3547 1263
rect 3513 1161 3547 1195
rect 3513 1093 3547 1127
rect 3601 1297 3635 1331
rect 3601 1229 3635 1263
rect 3601 1161 3635 1195
rect 3601 1111 3635 1127
rect 3740 1389 3757 1423
rect 3791 1389 3808 1423
rect 3740 1349 3808 1389
rect 3740 1315 3757 1349
rect 3791 1315 3808 1349
rect 3740 1275 3808 1315
rect 3740 1241 3757 1275
rect 3791 1241 3808 1275
rect 3740 1201 3808 1241
rect 3740 1167 3757 1201
rect 3791 1167 3808 1201
rect 3740 1127 3808 1167
rect 3740 1093 3757 1127
rect 3791 1093 3808 1127
rect 3513 1025 3643 1059
rect 3074 979 3142 1019
rect 3074 945 3091 979
rect 3125 945 3142 979
rect 2870 899 2977 933
rect 2154 299 2217 333
rect 2251 299 2314 333
rect 2120 261 2154 299
rect 2120 193 2154 227
rect 2314 261 2348 299
rect 2120 123 2154 159
rect 2120 73 2154 89
rect 2217 208 2251 224
rect 1964 34 2032 57
rect 2217 34 2251 174
rect 2314 193 2348 227
rect 2411 314 2533 348
rect 2630 461 2698 544
rect 2630 427 2647 461
rect 2681 427 2698 461
rect 2630 387 2698 427
rect 2630 353 2647 387
rect 2681 353 2698 387
rect 2795 434 2829 649
rect 2943 831 2977 899
rect 3074 905 3142 945
rect 3282 958 3316 974
rect 3468 958 3502 974
rect 3316 924 3347 942
rect 3282 908 3347 924
rect 3074 871 3091 905
rect 3125 871 3142 905
rect 3074 822 3142 871
rect 2943 433 2977 797
rect 3313 757 3347 908
rect 2795 384 2829 400
rect 2869 399 2977 433
rect 3074 461 3142 544
rect 3074 427 3091 461
rect 3125 427 3142 461
rect 2411 217 2445 314
rect 2630 313 2698 353
rect 2630 279 2647 313
rect 2681 279 2698 313
rect 2411 167 2445 183
rect 2508 261 2542 277
rect 2508 193 2542 227
rect 2314 123 2348 159
rect 2508 123 2542 159
rect 2348 89 2411 123
rect 2445 89 2508 123
rect 2314 73 2348 89
rect 2508 73 2542 89
rect 2630 239 2698 279
rect 2630 205 2647 239
rect 2681 205 2698 239
rect 2630 165 2698 205
rect 2630 131 2647 165
rect 2681 131 2698 165
rect 2630 91 2698 131
rect 2630 57 2647 91
rect 2681 57 2698 91
rect 2630 34 2698 57
rect 2773 334 2807 350
rect 2773 262 2807 300
rect 2773 194 2807 228
rect 2869 218 2903 399
rect 3074 387 3142 427
rect 3074 353 3091 387
rect 3125 353 3142 387
rect 3313 433 3347 723
rect 3313 383 3347 399
rect 3461 924 3468 942
rect 3461 908 3502 924
rect 3461 757 3495 908
rect 3461 433 3495 723
rect 3461 383 3495 399
rect 3609 683 3643 1025
rect 3740 1053 3808 1093
rect 3740 1019 3757 1053
rect 3791 1019 3808 1053
rect 3915 1365 3949 1405
rect 3915 1297 3949 1331
rect 3915 1229 3949 1263
rect 3915 1161 3949 1195
rect 3915 1093 3949 1127
rect 4003 1365 4037 1446
rect 4406 1423 4474 1446
rect 4003 1297 4037 1331
rect 4003 1229 4037 1263
rect 4003 1161 4037 1195
rect 4003 1111 4037 1127
rect 4091 1365 4301 1399
rect 4091 1297 4125 1331
rect 4091 1229 4125 1263
rect 4091 1161 4125 1195
rect 4091 1093 4125 1127
rect 3915 1025 4125 1059
rect 4179 1297 4213 1313
rect 4179 1229 4213 1263
rect 4179 1161 4213 1195
rect 4179 1093 4213 1127
rect 4267 1297 4301 1331
rect 4267 1229 4301 1263
rect 4267 1161 4301 1195
rect 4267 1111 4301 1127
rect 4406 1389 4423 1423
rect 4457 1389 4474 1423
rect 4406 1349 4474 1389
rect 4406 1315 4423 1349
rect 4457 1315 4474 1349
rect 4406 1275 4474 1315
rect 4406 1241 4423 1275
rect 4457 1241 4474 1275
rect 4406 1201 4474 1241
rect 4406 1167 4423 1201
rect 4457 1167 4474 1201
rect 4406 1127 4474 1167
rect 4406 1093 4423 1127
rect 4457 1093 4474 1127
rect 4179 1025 4309 1059
rect 3740 979 3808 1019
rect 3740 945 3757 979
rect 3791 945 3808 979
rect 3740 905 3808 945
rect 3948 958 3982 974
rect 4134 958 4168 974
rect 3982 924 4013 942
rect 3948 908 4013 924
rect 3740 871 3757 905
rect 3791 871 3808 905
rect 3740 822 3808 871
rect 2869 168 2903 184
rect 2967 334 3001 350
rect 2967 262 3001 300
rect 2967 194 3001 228
rect 2773 124 2807 160
rect 2967 124 3001 160
rect 2807 90 2869 124
rect 2903 90 2967 124
rect 2773 34 2807 90
rect 2870 34 2904 90
rect 2967 34 3001 90
rect 3074 313 3142 353
rect 3074 279 3091 313
rect 3125 279 3142 313
rect 3074 239 3142 279
rect 3074 205 3091 239
rect 3125 205 3142 239
rect 3074 165 3142 205
rect 3074 131 3091 165
rect 3125 131 3142 165
rect 3074 91 3142 131
rect 3074 57 3091 91
rect 3125 57 3142 91
rect 3074 34 3142 57
rect 3230 333 3264 349
rect 3609 348 3643 649
rect 3979 683 4013 908
rect 3230 261 3264 299
rect 3230 193 3264 227
rect 3327 314 3643 348
rect 3740 461 3808 544
rect 3740 427 3757 461
rect 3791 427 3808 461
rect 3740 387 3808 427
rect 3740 353 3757 387
rect 3791 353 3808 387
rect 3979 433 4013 649
rect 3979 383 4013 399
rect 4127 924 4134 942
rect 4127 908 4168 924
rect 4127 831 4161 908
rect 4127 433 4161 797
rect 4127 383 4161 399
rect 4275 757 4309 1025
rect 4406 1053 4474 1093
rect 4406 1019 4423 1053
rect 4457 1019 4474 1053
rect 4406 979 4474 1019
rect 4406 945 4423 979
rect 4457 945 4474 979
rect 4406 905 4474 945
rect 4406 871 4423 905
rect 4457 871 4474 905
rect 4406 822 4474 871
rect 3327 217 3361 314
rect 3327 167 3361 183
rect 3424 261 3458 278
rect 3424 193 3458 227
rect 3230 123 3264 159
rect 3521 217 3555 314
rect 3740 313 3808 353
rect 3740 279 3757 313
rect 3791 279 3808 313
rect 3521 167 3555 183
rect 3618 261 3652 278
rect 3618 193 3652 227
rect 3424 123 3458 159
rect 3618 123 3652 159
rect 3264 89 3327 123
rect 3361 89 3424 123
rect 3458 89 3521 123
rect 3555 89 3618 123
rect 3230 34 3264 89
rect 3327 34 3361 89
rect 3424 34 3458 89
rect 3521 34 3555 89
rect 3618 34 3652 89
rect 3740 239 3808 279
rect 3740 205 3757 239
rect 3791 205 3808 239
rect 3740 165 3808 205
rect 3740 131 3757 165
rect 3791 131 3808 165
rect 3740 91 3808 131
rect 3740 57 3757 91
rect 3791 57 3808 91
rect 3740 34 3808 57
rect 3896 333 3930 349
rect 4275 348 4309 723
rect 3896 261 3930 299
rect 3896 193 3930 227
rect 3993 314 4309 348
rect 4406 461 4474 544
rect 4406 427 4423 461
rect 4457 427 4474 461
rect 4406 387 4474 427
rect 4406 353 4423 387
rect 4457 353 4474 387
rect 3993 217 4027 314
rect 3993 167 4027 183
rect 4090 261 4124 278
rect 4090 193 4124 227
rect 3896 123 3930 159
rect 4187 217 4221 314
rect 4406 313 4474 353
rect 4406 279 4423 313
rect 4457 279 4474 313
rect 4187 167 4221 183
rect 4284 261 4318 278
rect 4284 193 4318 227
rect 4090 123 4124 159
rect 4284 123 4318 159
rect 3930 89 3993 123
rect 4027 89 4090 123
rect 4124 89 4187 123
rect 4221 89 4284 123
rect 3896 34 3930 89
rect 3993 34 4027 89
rect 4090 34 4124 89
rect 4187 34 4221 89
rect 4284 34 4318 89
rect 4406 239 4474 279
rect 4406 205 4423 239
rect 4457 205 4474 239
rect 4406 165 4474 205
rect 4406 131 4423 165
rect 4457 131 4474 165
rect 4406 91 4474 131
rect 4406 57 4423 91
rect 4457 57 4474 91
rect 4406 34 4474 57
rect -34 17 4474 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4474 17
rect -34 -34 4474 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 279 575 313 609
rect 575 797 609 831
rect 723 723 757 757
rect 1093 723 1127 757
rect 1241 575 1275 609
rect 1389 649 1423 683
rect 1685 649 1719 683
rect 1833 723 1867 757
rect 2203 575 2237 609
rect 2351 797 2385 831
rect 2499 649 2533 683
rect 2795 649 2829 683
rect 2943 797 2977 831
rect 3313 723 3347 757
rect 3461 723 3495 757
rect 3609 649 3643 683
rect 3979 649 4013 683
rect 4127 797 4161 831
rect 4275 723 4309 757
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
<< metal1 >>
rect -34 1497 4474 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4474 1497
rect -34 1446 4474 1463
rect 569 831 615 837
rect 2345 831 2391 837
rect 2937 831 2983 837
rect 4121 831 4167 837
rect 563 797 575 831
rect 609 797 2351 831
rect 2385 797 2397 831
rect 2931 797 2943 831
rect 2977 797 4127 831
rect 4161 797 4173 831
rect 569 791 615 797
rect 2345 791 2391 797
rect 2937 791 2983 797
rect 4121 791 4167 797
rect 717 757 763 763
rect 1087 757 1133 763
rect 1827 757 1873 763
rect 3307 757 3353 763
rect 3455 757 3501 763
rect 4269 757 4315 763
rect 711 723 723 757
rect 757 723 1093 757
rect 1127 723 1139 757
rect 1821 723 1833 757
rect 1867 723 3313 757
rect 3347 723 3359 757
rect 3449 723 3461 757
rect 3495 723 4275 757
rect 4309 723 4321 757
rect 717 717 763 723
rect 1087 717 1133 723
rect 1827 717 1873 723
rect 3307 717 3353 723
rect 3455 717 3501 723
rect 4269 717 4315 723
rect 1383 683 1429 689
rect 1679 683 1725 689
rect 2493 683 2539 689
rect 2789 683 2835 689
rect 3603 683 3649 689
rect 3973 683 4019 689
rect 1377 649 1389 683
rect 1423 649 1685 683
rect 1719 649 1731 683
rect 2487 649 2499 683
rect 2533 649 2795 683
rect 2829 649 2841 683
rect 3597 649 3609 683
rect 3643 649 3979 683
rect 4013 649 4025 683
rect 1383 643 1429 649
rect 1679 643 1725 649
rect 2493 643 2539 649
rect 2789 643 2835 649
rect 3603 643 3649 649
rect 3973 643 4019 649
rect 273 609 319 615
rect 1235 609 1281 615
rect 2197 609 2243 615
rect 267 575 279 609
rect 313 575 1241 609
rect 1275 575 2203 609
rect 2237 575 2249 609
rect 273 569 319 575
rect 1235 569 1281 575
rect 2197 569 2243 575
rect -34 17 4474 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4474 17
rect -34 -34 4474 -17
<< labels >>
rlabel metal1 3609 649 3643 683 1 Q
port 1 n
rlabel metal1 3609 575 3643 609 1 Q
port 2 n
rlabel metal1 3609 501 3643 535 1 Q
port 3 n
rlabel metal1 3609 427 3643 461 1 Q
port 4 n
rlabel metal1 3609 871 3643 905 1 Q
port 5 n
rlabel metal1 3979 427 4013 461 1 Q
port 6 n
rlabel metal1 3979 501 4013 535 1 Q
port 7 n
rlabel metal1 3979 575 4013 609 1 Q
port 8 n
rlabel metal1 3979 649 4013 683 1 Q
port 9 n
rlabel metal1 3979 871 4013 905 1 Q
port 10 n
rlabel metal1 575 797 609 831 1 D
port 11 n
rlabel metal1 575 871 609 905 1 D
port 12 n
rlabel metal1 575 723 609 757 1 D
port 13 n
rlabel metal1 575 649 609 683 1 D
port 14 n
rlabel metal1 575 501 609 535 1 D
port 15 n
rlabel metal1 2351 649 2385 683 1 D
port 16 n
rlabel metal1 2351 797 2385 831 1 D
port 17 n
rlabel metal1 2351 871 2385 905 1 D
port 18 n
rlabel metal1 2351 575 2385 609 1 D
port 19 n
rlabel metal1 2351 501 2385 535 1 D
port 20 n
rlabel metal1 131 575 165 609 1 GATE_N
port 21 n
rlabel metal1 131 501 165 535 1 GATE_N
port 22 n
rlabel metal1 131 649 165 683 1 GATE_N
port 23 n
rlabel metal1 131 723 165 757 1 GATE_N
port 24 n
rlabel metal1 131 797 165 831 1 GATE_N
port 25 n
rlabel metal1 131 871 165 905 1 GATE_N
port 26 n
rlabel metal1 -34 1446 4474 1514 1 VPWR
port 27 n
rlabel metal1 -34 -34 4474 34 1 VGND
port 28 n
rlabel nwell 57 1463 91 1497 1 VPB
port 29 n
rlabel pwell 57 -17 91 17 1 VNB
port 30 n
<< end >>
