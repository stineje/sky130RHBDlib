magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1 21 1650 203
rect 30 -17 64 21
<< locali >>
rect 17 199 66 323
rect 974 323 1040 425
rect 1142 323 1208 425
rect 1310 323 1376 425
rect 1478 323 1544 425
rect 974 289 1544 323
rect 974 170 1050 289
rect 1084 204 1639 255
rect 974 127 1639 170
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 17 391 69 493
rect 103 425 175 527
rect 17 357 175 391
rect 100 265 175 357
rect 215 345 257 493
rect 291 379 357 527
rect 391 345 425 493
rect 459 379 525 527
rect 559 345 593 493
rect 627 379 693 527
rect 727 345 761 493
rect 795 379 861 527
rect 895 459 1639 493
rect 895 345 940 459
rect 215 311 940 345
rect 1074 357 1108 459
rect 1242 357 1276 459
rect 1410 357 1444 459
rect 1578 289 1639 459
rect 100 199 940 265
rect 100 165 139 199
rect 17 131 139 165
rect 207 131 940 165
rect 17 51 69 131
rect 103 17 169 97
rect 207 51 241 131
rect 275 17 341 97
rect 375 51 409 131
rect 443 17 509 97
rect 543 51 577 131
rect 611 17 677 97
rect 711 51 745 131
rect 779 17 847 97
rect 881 93 940 131
rect 881 51 1639 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
rlabel locali s 1084 204 1639 255 6 A
port 1 nsew signal input
rlabel locali s 17 199 66 323 6 TE
port 2 nsew signal input
rlabel metal1 s 0 -48 1656 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1650 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1694 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1656 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 974 127 1639 170 6 Z
port 7 nsew signal output
rlabel locali s 974 170 1050 289 6 Z
port 7 nsew signal output
rlabel locali s 974 289 1544 323 6 Z
port 7 nsew signal output
rlabel locali s 1478 323 1544 425 6 Z
port 7 nsew signal output
rlabel locali s 1310 323 1376 425 6 Z
port 7 nsew signal output
rlabel locali s 1142 323 1208 425 6 Z
port 7 nsew signal output
rlabel locali s 974 323 1040 425 6 Z
port 7 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1656 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2051578
string GDS_START 2038956
<< end >>
