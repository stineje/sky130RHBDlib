* SPICE3 file created from DFFQX1.ext - technology: sky130A

.subckt DFFQX1 Q D CLK VDD GND
M1000 a_599_989.t4 D.t0 VDD.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 GND a_1845_1050.t5 a_2406_101.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1002 a_1845_1050.t4 a_599_989.t5 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t2 a_147_187.t6 a_1845_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD.t22 a_147_187.t7 a_277_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 GND a_147_187.t8 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_3177_1050.t1 a_277_1050.t7 VDD.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t9 a_1845_1050.t6 a_147_187.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t14 CLK.t0 a_277_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 GND a_599_989.t8 a_1740_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1010 VDD.t15 CLK.t1 a_147_187.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_3177_1050.t3 Q.t6 VDD.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 Q.t4 a_3177_1050.t5 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VDD.t12 a_599_989.t7 a_277_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t16 a_277_1050.t8 a_599_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD.t21 a_147_187.t9 Q.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1845_1050.t0 a_147_187.t10 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 GND a_3177_1050.t6 a_3738_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q.t0 a_147_187.t11 VDD.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VDD.t25 D.t2 a_599_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_277_1050.t0 a_147_187.t12 VDD.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 GND a_277_1050.t10 a_1074_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t10 a_599_989.t9 a_1845_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_277_1050.t6 CLK.t4 VDD.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VDD.t3 a_277_1050.t9 a_3177_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_147_187.t3 CLK.t5 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 GND a_277_1050.t12 a_3072_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_277_1050.t4 a_599_989.t10 VDD.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_599_989.t0 a_277_1050.t11 VDD.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q a_147_187.t5 a_3738_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1030 a_147_187.t0 a_1845_1050.t7 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 VDD.t4 Q.t7 a_3177_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 VDD.t7 a_3177_1050.t7 Q.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 CLK D 0.07fF
C1 VDD D 0.07fF
C2 VDD Q 1.43fF
C3 VDD CLK 0.40fF
R0 D.n0 D.t2 472.359
R1 D.n0 D.t0 384.527
R2 D.n1 D.t1 220.772
R3 D.n1 D.n0 136.613
R4 D.n2 D.n1 76
R5 D.n2 D 0.046
R6 VDD.n315 VDD.n313 144.705
R7 VDD.n205 VDD.n203 144.705
R8 VDD.n376 VDD.n374 144.705
R9 VDD.n144 VDD.n142 144.705
R10 VDD.n83 VDD.n81 144.705
R11 VDD.n44 VDD.n43 76
R12 VDD.n49 VDD.n48 76
R13 VDD.n54 VDD.n53 76
R14 VDD.n58 VDD.n57 76
R15 VDD.n85 VDD.n84 76
R16 VDD.n90 VDD.n89 76
R17 VDD.n95 VDD.n94 76
R18 VDD.n101 VDD.n100 76
R19 VDD.n106 VDD.n105 76
R20 VDD.n111 VDD.n110 76
R21 VDD.n116 VDD.n115 76
R22 VDD.n120 VDD.n119 76
R23 VDD.n146 VDD.n145 76
R24 VDD.n151 VDD.n150 76
R25 VDD.n156 VDD.n155 76
R26 VDD.n162 VDD.n161 76
R27 VDD.n167 VDD.n166 76
R28 VDD.n172 VDD.n171 76
R29 VDD.n177 VDD.n176 76
R30 VDD.n181 VDD.n180 76
R31 VDD.n207 VDD.n206 76
R32 VDD.n212 VDD.n211 76
R33 VDD.n404 VDD.n403 76
R34 VDD.n399 VDD.n398 76
R35 VDD.n393 VDD.n392 76
R36 VDD.n388 VDD.n387 76
R37 VDD.n383 VDD.n382 76
R38 VDD.n378 VDD.n377 76
R39 VDD.n352 VDD.n351 76
R40 VDD.n348 VDD.n347 76
R41 VDD.n343 VDD.n342 76
R42 VDD.n338 VDD.n337 76
R43 VDD.n332 VDD.n331 76
R44 VDD.n327 VDD.n326 76
R45 VDD.n322 VDD.n321 76
R46 VDD.n317 VDD.n316 76
R47 VDD.n290 VDD.n289 76
R48 VDD.n286 VDD.n285 76
R49 VDD.n282 VDD.n281 76
R50 VDD.n278 VDD.n277 76
R51 VDD.n273 VDD.n272 76
R52 VDD.n266 VDD.n265 76
R53 VDD.n261 VDD.n260 76
R54 VDD.n256 VDD.n255 76
R55 VDD.n249 VDD.n248 76
R56 VDD.n244 VDD.n243 76
R57 VDD.n239 VDD.n238 76
R58 VDD.n235 VDD.n234 76
R59 VDD.n275 VDD.n274 64.064
R60 VDD.n246 VDD.n245 59.488
R61 VDD.n240 VDD.t17 55.106
R62 VDD.n318 VDD.t13 55.106
R63 VDD.n379 VDD.t0 55.106
R64 VDD.n173 VDD.t1 55.106
R65 VDD.n112 VDD.t6 55.106
R66 VDD.n50 VDD.t8 55.106
R67 VDD.n281 VDD.t12 55.106
R68 VDD.n344 VDD.t25 55.106
R69 VDD.n208 VDD.t2 55.106
R70 VDD.n147 VDD.t15 55.106
R71 VDD.n86 VDD.t4 55.106
R72 VDD.n33 VDD.t21 55.106
R73 VDD.n251 VDD.n250 40.824
R74 VDD.n271 VDD.n270 40.824
R75 VDD.n334 VDD.n333 40.824
R76 VDD.n395 VDD.n394 40.824
R77 VDD.n158 VDD.n157 40.824
R78 VDD.n97 VDD.n96 40.824
R79 VDD.n28 VDD.n27 40.824
R80 VDD.n357 VDD.n356 36.774
R81 VDD.n186 VDD.n185 36.774
R82 VDD.n125 VDD.n124 36.774
R83 VDD.n63 VDD.n62 36.774
R84 VDD.n306 VDD.n305 36.774
R85 VDD.n25 VDD.n24 36.608
R86 VDD.n92 VDD.n91 36.608
R87 VDD.n153 VDD.n152 36.608
R88 VDD.n401 VDD.n400 36.608
R89 VDD.n340 VDD.n339 36.608
R90 VDD.n38 VDD.n37 34.942
R91 VDD.n46 VDD.n45 32.032
R92 VDD.n108 VDD.n107 32.032
R93 VDD.n169 VDD.n168 32.032
R94 VDD.n385 VDD.n384 32.032
R95 VDD.n324 VDD.n323 32.032
R96 VDD.n268 VDD.n267 27.456
R97 VDD.n253 VDD.n252 22.88
R98 VDD.n234 VDD.n231 21.841
R99 VDD.n23 VDD.n20 21.841
R100 VDD.n250 VDD.t19 14.282
R101 VDD.n250 VDD.t22 14.282
R102 VDD.n270 VDD.t11 14.282
R103 VDD.n270 VDD.t14 14.282
R104 VDD.n333 VDD.t24 14.282
R105 VDD.n333 VDD.t16 14.282
R106 VDD.n394 VDD.t5 14.282
R107 VDD.n394 VDD.t10 14.282
R108 VDD.n157 VDD.t18 14.282
R109 VDD.n157 VDD.t9 14.282
R110 VDD.n96 VDD.t20 14.282
R111 VDD.n96 VDD.t3 14.282
R112 VDD.n27 VDD.t23 14.282
R113 VDD.n27 VDD.t7 14.282
R114 VDD.n231 VDD.n214 14.167
R115 VDD.n214 VDD.n213 14.167
R116 VDD.n372 VDD.n354 14.167
R117 VDD.n354 VDD.n353 14.167
R118 VDD.n201 VDD.n183 14.167
R119 VDD.n183 VDD.n182 14.167
R120 VDD.n140 VDD.n122 14.167
R121 VDD.n122 VDD.n121 14.167
R122 VDD.n79 VDD.n60 14.167
R123 VDD.n60 VDD.n59 14.167
R124 VDD.n311 VDD.n292 14.167
R125 VDD.n292 VDD.n291 14.167
R126 VDD.n20 VDD.n19 14.167
R127 VDD.n19 VDD.n17 14.167
R128 VDD.n32 VDD.n31 14.167
R129 VDD.n84 VDD.n80 14.167
R130 VDD.n145 VDD.n141 14.167
R131 VDD.n206 VDD.n202 14.167
R132 VDD.n377 VDD.n373 14.167
R133 VDD.n316 VDD.n312 14.167
R134 VDD.n258 VDD.n257 13.728
R135 VDD.n23 VDD.n22 13.653
R136 VDD.n22 VDD.n21 13.653
R137 VDD.n36 VDD.n35 13.653
R138 VDD.n35 VDD.n34 13.653
R139 VDD.n32 VDD.n26 13.653
R140 VDD.n26 VDD.n25 13.653
R141 VDD.n31 VDD.n30 13.653
R142 VDD.n30 VDD.n29 13.653
R143 VDD.n43 VDD.n42 13.653
R144 VDD.n42 VDD.n41 13.653
R145 VDD.n48 VDD.n47 13.653
R146 VDD.n47 VDD.n46 13.653
R147 VDD.n53 VDD.n52 13.653
R148 VDD.n52 VDD.n51 13.653
R149 VDD.n57 VDD.n56 13.653
R150 VDD.n56 VDD.n55 13.653
R151 VDD.n84 VDD.n83 13.653
R152 VDD.n83 VDD.n82 13.653
R153 VDD.n89 VDD.n88 13.653
R154 VDD.n88 VDD.n87 13.653
R155 VDD.n94 VDD.n93 13.653
R156 VDD.n93 VDD.n92 13.653
R157 VDD.n100 VDD.n99 13.653
R158 VDD.n99 VDD.n98 13.653
R159 VDD.n105 VDD.n104 13.653
R160 VDD.n104 VDD.n103 13.653
R161 VDD.n110 VDD.n109 13.653
R162 VDD.n109 VDD.n108 13.653
R163 VDD.n115 VDD.n114 13.653
R164 VDD.n114 VDD.n113 13.653
R165 VDD.n119 VDD.n118 13.653
R166 VDD.n118 VDD.n117 13.653
R167 VDD.n145 VDD.n144 13.653
R168 VDD.n144 VDD.n143 13.653
R169 VDD.n150 VDD.n149 13.653
R170 VDD.n149 VDD.n148 13.653
R171 VDD.n155 VDD.n154 13.653
R172 VDD.n154 VDD.n153 13.653
R173 VDD.n161 VDD.n160 13.653
R174 VDD.n160 VDD.n159 13.653
R175 VDD.n166 VDD.n165 13.653
R176 VDD.n165 VDD.n164 13.653
R177 VDD.n171 VDD.n170 13.653
R178 VDD.n170 VDD.n169 13.653
R179 VDD.n176 VDD.n175 13.653
R180 VDD.n175 VDD.n174 13.653
R181 VDD.n180 VDD.n179 13.653
R182 VDD.n179 VDD.n178 13.653
R183 VDD.n206 VDD.n205 13.653
R184 VDD.n205 VDD.n204 13.653
R185 VDD.n211 VDD.n210 13.653
R186 VDD.n210 VDD.n209 13.653
R187 VDD.n403 VDD.n402 13.653
R188 VDD.n402 VDD.n401 13.653
R189 VDD.n398 VDD.n397 13.653
R190 VDD.n397 VDD.n396 13.653
R191 VDD.n392 VDD.n391 13.653
R192 VDD.n391 VDD.n390 13.653
R193 VDD.n387 VDD.n386 13.653
R194 VDD.n386 VDD.n385 13.653
R195 VDD.n382 VDD.n381 13.653
R196 VDD.n381 VDD.n380 13.653
R197 VDD.n377 VDD.n376 13.653
R198 VDD.n376 VDD.n375 13.653
R199 VDD.n351 VDD.n350 13.653
R200 VDD.n350 VDD.n349 13.653
R201 VDD.n347 VDD.n346 13.653
R202 VDD.n346 VDD.n345 13.653
R203 VDD.n342 VDD.n341 13.653
R204 VDD.n341 VDD.n340 13.653
R205 VDD.n337 VDD.n336 13.653
R206 VDD.n336 VDD.n335 13.653
R207 VDD.n331 VDD.n330 13.653
R208 VDD.n330 VDD.n329 13.653
R209 VDD.n326 VDD.n325 13.653
R210 VDD.n325 VDD.n324 13.653
R211 VDD.n321 VDD.n320 13.653
R212 VDD.n320 VDD.n319 13.653
R213 VDD.n316 VDD.n315 13.653
R214 VDD.n315 VDD.n314 13.653
R215 VDD.n289 VDD.n288 13.653
R216 VDD.n288 VDD.n287 13.653
R217 VDD.n285 VDD.n284 13.653
R218 VDD.n284 VDD.n283 13.653
R219 VDD.n281 VDD.n280 13.653
R220 VDD.n280 VDD.n279 13.653
R221 VDD.n277 VDD.n276 13.653
R222 VDD.n276 VDD.n275 13.653
R223 VDD.n272 VDD.n269 13.653
R224 VDD.n269 VDD.n268 13.653
R225 VDD.n265 VDD.n264 13.653
R226 VDD.n264 VDD.n263 13.653
R227 VDD.n260 VDD.n259 13.653
R228 VDD.n259 VDD.n258 13.653
R229 VDD.n255 VDD.n254 13.653
R230 VDD.n254 VDD.n253 13.653
R231 VDD.n248 VDD.n247 13.653
R232 VDD.n247 VDD.n246 13.653
R233 VDD.n243 VDD.n242 13.653
R234 VDD.n242 VDD.n241 13.653
R235 VDD.n238 VDD.n237 13.653
R236 VDD.n237 VDD.n236 13.653
R237 VDD.n234 VDD.n233 13.653
R238 VDD.n233 VDD.n232 13.653
R239 VDD.n4 VDD.n2 12.915
R240 VDD.n4 VDD.n3 12.66
R241 VDD.n12 VDD.n11 12.343
R242 VDD.n8 VDD.n7 12.343
R243 VDD.n12 VDD.n9 12.343
R244 VDD.n33 VDD.n32 11.806
R245 VDD.n263 VDD.n262 9.152
R246 VDD.n31 VDD.n28 8.658
R247 VDD.n100 VDD.n97 8.658
R248 VDD.n161 VDD.n158 8.658
R249 VDD.n398 VDD.n395 8.658
R250 VDD.n337 VDD.n334 8.658
R251 VDD.n373 VDD.n372 7.674
R252 VDD.n202 VDD.n201 7.674
R253 VDD.n141 VDD.n140 7.674
R254 VDD.n80 VDD.n79 7.674
R255 VDD.n312 VDD.n311 7.674
R256 VDD.n74 VDD.n73 7.5
R257 VDD.n68 VDD.n67 7.5
R258 VDD.n70 VDD.n69 7.5
R259 VDD.n65 VDD.n64 7.5
R260 VDD.n79 VDD.n78 7.5
R261 VDD.n135 VDD.n134 7.5
R262 VDD.n129 VDD.n128 7.5
R263 VDD.n131 VDD.n130 7.5
R264 VDD.n137 VDD.n127 7.5
R265 VDD.n137 VDD.n125 7.5
R266 VDD.n140 VDD.n139 7.5
R267 VDD.n196 VDD.n195 7.5
R268 VDD.n190 VDD.n189 7.5
R269 VDD.n192 VDD.n191 7.5
R270 VDD.n198 VDD.n188 7.5
R271 VDD.n198 VDD.n186 7.5
R272 VDD.n201 VDD.n200 7.5
R273 VDD.n367 VDD.n366 7.5
R274 VDD.n361 VDD.n360 7.5
R275 VDD.n363 VDD.n362 7.5
R276 VDD.n369 VDD.n359 7.5
R277 VDD.n369 VDD.n357 7.5
R278 VDD.n372 VDD.n371 7.5
R279 VDD.n296 VDD.n295 7.5
R280 VDD.n299 VDD.n298 7.5
R281 VDD.n301 VDD.n300 7.5
R282 VDD.n304 VDD.n303 7.5
R283 VDD.n311 VDD.n310 7.5
R284 VDD.n226 VDD.n225 7.5
R285 VDD.n220 VDD.n219 7.5
R286 VDD.n222 VDD.n221 7.5
R287 VDD.n228 VDD.n218 7.5
R288 VDD.n228 VDD.n216 7.5
R289 VDD.n231 VDD.n230 7.5
R290 VDD.n20 VDD.n16 7.5
R291 VDD.n2 VDD.n1 7.5
R292 VDD.n7 VDD.n6 7.5
R293 VDD.n11 VDD.n10 7.5
R294 VDD.n19 VDD.n18 7.5
R295 VDD.n14 VDD.n0 7.5
R296 VDD.n66 VDD.n63 6.772
R297 VDD.n77 VDD.n61 6.772
R298 VDD.n75 VDD.n72 6.772
R299 VDD.n71 VDD.n68 6.772
R300 VDD.n138 VDD.n123 6.772
R301 VDD.n136 VDD.n133 6.772
R302 VDD.n132 VDD.n129 6.772
R303 VDD.n199 VDD.n184 6.772
R304 VDD.n197 VDD.n194 6.772
R305 VDD.n193 VDD.n190 6.772
R306 VDD.n370 VDD.n355 6.772
R307 VDD.n368 VDD.n365 6.772
R308 VDD.n364 VDD.n361 6.772
R309 VDD.n229 VDD.n215 6.772
R310 VDD.n227 VDD.n224 6.772
R311 VDD.n223 VDD.n220 6.772
R312 VDD.n66 VDD.n65 6.772
R313 VDD.n71 VDD.n70 6.772
R314 VDD.n75 VDD.n74 6.772
R315 VDD.n78 VDD.n77 6.772
R316 VDD.n132 VDD.n131 6.772
R317 VDD.n136 VDD.n135 6.772
R318 VDD.n139 VDD.n138 6.772
R319 VDD.n193 VDD.n192 6.772
R320 VDD.n197 VDD.n196 6.772
R321 VDD.n200 VDD.n199 6.772
R322 VDD.n364 VDD.n363 6.772
R323 VDD.n368 VDD.n367 6.772
R324 VDD.n371 VDD.n370 6.772
R325 VDD.n223 VDD.n222 6.772
R326 VDD.n227 VDD.n226 6.772
R327 VDD.n230 VDD.n229 6.772
R328 VDD.n310 VDD.n309 6.772
R329 VDD.n297 VDD.n294 6.772
R330 VDD.n302 VDD.n299 6.772
R331 VDD.n307 VDD.n304 6.772
R332 VDD.n307 VDD.n306 6.772
R333 VDD.n302 VDD.n301 6.772
R334 VDD.n297 VDD.n296 6.772
R335 VDD.n309 VDD.n293 6.772
R336 VDD.n255 VDD.n251 6.69
R337 VDD.n37 VDD.n23 6.487
R338 VDD.n37 VDD.n36 6.475
R339 VDD.n16 VDD.n15 6.458
R340 VDD.n272 VDD.n271 6.296
R341 VDD.n127 VDD.n126 6.202
R342 VDD.n188 VDD.n187 6.202
R343 VDD.n359 VDD.n358 6.202
R344 VDD.n218 VDD.n217 6.202
R345 VDD.n41 VDD.n40 4.576
R346 VDD.n103 VDD.n102 4.576
R347 VDD.n164 VDD.n163 4.576
R348 VDD.n390 VDD.n389 4.576
R349 VDD.n329 VDD.n328 4.576
R350 VDD.n53 VDD.n50 2.754
R351 VDD.n115 VDD.n112 2.754
R352 VDD.n176 VDD.n173 2.754
R353 VDD.n382 VDD.n379 2.754
R354 VDD.n321 VDD.n318 2.754
R355 VDD.n36 VDD.n33 2.361
R356 VDD.n89 VDD.n86 2.361
R357 VDD.n150 VDD.n147 2.361
R358 VDD.n211 VDD.n208 2.361
R359 VDD.n347 VDD.n344 2.361
R360 VDD.n14 VDD.n5 1.329
R361 VDD.n14 VDD.n8 1.329
R362 VDD.n14 VDD.n12 1.329
R363 VDD.n14 VDD.n13 1.329
R364 VDD.n15 VDD.n14 0.696
R365 VDD.n14 VDD.n4 0.696
R366 VDD.n243 VDD.n240 0.393
R367 VDD.n76 VDD.n75 0.365
R368 VDD.n76 VDD.n71 0.365
R369 VDD.n76 VDD.n66 0.365
R370 VDD.n77 VDD.n76 0.365
R371 VDD.n137 VDD.n136 0.365
R372 VDD.n137 VDD.n132 0.365
R373 VDD.n138 VDD.n137 0.365
R374 VDD.n198 VDD.n197 0.365
R375 VDD.n198 VDD.n193 0.365
R376 VDD.n199 VDD.n198 0.365
R377 VDD.n369 VDD.n368 0.365
R378 VDD.n369 VDD.n364 0.365
R379 VDD.n370 VDD.n369 0.365
R380 VDD.n228 VDD.n227 0.365
R381 VDD.n228 VDD.n223 0.365
R382 VDD.n229 VDD.n228 0.365
R383 VDD.n308 VDD.n307 0.365
R384 VDD.n308 VDD.n302 0.365
R385 VDD.n308 VDD.n297 0.365
R386 VDD.n309 VDD.n308 0.365
R387 VDD.n85 VDD.n58 0.29
R388 VDD.n146 VDD.n120 0.29
R389 VDD.n207 VDD.n181 0.29
R390 VDD.n378 VDD.n352 0.29
R391 VDD.n317 VDD.n290 0.29
R392 VDD.n235 VDD 0.207
R393 VDD.n266 VDD.n261 0.197
R394 VDD.n44 VDD.n39 0.181
R395 VDD.n106 VDD.n101 0.181
R396 VDD.n167 VDD.n162 0.181
R397 VDD.n399 VDD.n393 0.181
R398 VDD.n338 VDD.n332 0.181
R399 VDD.n39 VDD.n38 0.145
R400 VDD.n49 VDD.n44 0.145
R401 VDD.n54 VDD.n49 0.145
R402 VDD.n58 VDD.n54 0.145
R403 VDD.n90 VDD.n85 0.145
R404 VDD.n95 VDD.n90 0.145
R405 VDD.n101 VDD.n95 0.145
R406 VDD.n111 VDD.n106 0.145
R407 VDD.n116 VDD.n111 0.145
R408 VDD.n120 VDD.n116 0.145
R409 VDD.n151 VDD.n146 0.145
R410 VDD.n156 VDD.n151 0.145
R411 VDD.n162 VDD.n156 0.145
R412 VDD.n172 VDD.n167 0.145
R413 VDD.n177 VDD.n172 0.145
R414 VDD.n181 VDD.n177 0.145
R415 VDD.n212 VDD.n207 0.145
R416 VDD.n404 VDD.n399 0.145
R417 VDD.n393 VDD.n388 0.145
R418 VDD.n388 VDD.n383 0.145
R419 VDD.n383 VDD.n378 0.145
R420 VDD.n352 VDD.n348 0.145
R421 VDD.n348 VDD.n343 0.145
R422 VDD.n343 VDD.n338 0.145
R423 VDD.n332 VDD.n327 0.145
R424 VDD.n327 VDD.n322 0.145
R425 VDD.n322 VDD.n317 0.145
R426 VDD.n290 VDD.n286 0.145
R427 VDD.n286 VDD.n282 0.145
R428 VDD.n282 VDD.n278 0.145
R429 VDD.n278 VDD.n273 0.145
R430 VDD.n273 VDD.n266 0.145
R431 VDD.n261 VDD.n256 0.145
R432 VDD.n256 VDD.n249 0.145
R433 VDD.n249 VDD.n244 0.145
R434 VDD.n244 VDD.n239 0.145
R435 VDD.n239 VDD.n235 0.145
R436 VDD VDD.n404 0.137
R437 VDD VDD.n212 0.008
R438 a_599_989.n0 a_599_989.t9 480.392
R439 a_599_989.n2 a_599_989.t10 454.685
R440 a_599_989.n2 a_599_989.t7 428.979
R441 a_599_989.n0 a_599_989.t5 403.272
R442 a_599_989.n1 a_599_989.t8 283.48
R443 a_599_989.n3 a_599_989.t6 237.959
R444 a_599_989.n9 a_599_989.n8 210.592
R445 a_599_989.n11 a_599_989.n9 152.499
R446 a_599_989.n3 a_599_989.n2 98.447
R447 a_599_989.n1 a_599_989.n0 98.447
R448 a_599_989.n4 a_599_989.n3 78.947
R449 a_599_989.n4 a_599_989.n1 77.315
R450 a_599_989.n11 a_599_989.n10 76.002
R451 a_599_989.n9 a_599_989.n4 76
R452 a_599_989.n8 a_599_989.n7 30
R453 a_599_989.n6 a_599_989.n5 24.383
R454 a_599_989.n8 a_599_989.n6 23.684
R455 a_599_989.n10 a_599_989.t1 14.282
R456 a_599_989.n10 a_599_989.t0 14.282
R457 a_599_989.n12 a_599_989.t3 14.282
R458 a_599_989.t4 a_599_989.n12 14.282
R459 a_599_989.n12 a_599_989.n11 12.848
R460 a_147_187.n8 a_147_187.t7 512.525
R461 a_147_187.n6 a_147_187.t6 472.359
R462 a_147_187.n4 a_147_187.t9 472.359
R463 a_147_187.n6 a_147_187.t10 384.527
R464 a_147_187.n4 a_147_187.t11 384.527
R465 a_147_187.n8 a_147_187.t12 371.139
R466 a_147_187.n9 a_147_187.t8 340.774
R467 a_147_187.n7 a_147_187.t13 294.278
R468 a_147_187.n5 a_147_187.t5 294.278
R469 a_147_187.n14 a_147_187.n12 263.698
R470 a_147_187.n9 a_147_187.n8 109.607
R471 a_147_187.n12 a_147_187.n3 99.394
R472 a_147_187.n10 a_147_187.n9 82.484
R473 a_147_187.n11 a_147_187.n5 80.307
R474 a_147_187.n3 a_147_187.n2 76.002
R475 a_147_187.n10 a_147_187.n7 76
R476 a_147_187.n12 a_147_187.n11 76
R477 a_147_187.n7 a_147_187.n6 56.954
R478 a_147_187.n5 a_147_187.n4 56.954
R479 a_147_187.n14 a_147_187.n13 30
R480 a_147_187.n15 a_147_187.n0 24.383
R481 a_147_187.n15 a_147_187.n14 23.684
R482 a_147_187.n1 a_147_187.t2 14.282
R483 a_147_187.n1 a_147_187.t3 14.282
R484 a_147_187.n2 a_147_187.t1 14.282
R485 a_147_187.n2 a_147_187.t0 14.282
R486 a_147_187.n3 a_147_187.n1 12.85
R487 a_147_187.n11 a_147_187.n10 2.947
R488 a_3738_101.n5 a_3738_101.n4 24.877
R489 a_3738_101.t0 a_3738_101.n5 12.677
R490 a_3738_101.t0 a_3738_101.n3 11.595
R491 a_3738_101.t0 a_3738_101.n6 8.137
R492 a_3738_101.n2 a_3738_101.n0 4.031
R493 a_3738_101.n2 a_3738_101.n1 3.644
R494 a_3738_101.t0 a_3738_101.n2 1.093
R495 Q.n5 Q.t7 472.359
R496 Q.n5 Q.t6 384.527
R497 Q.n6 Q.t5 267.725
R498 Q.n4 Q.n3 258.884
R499 Q.n4 Q.n2 125.947
R500 Q.n6 Q.n5 83.507
R501 Q Q.n6 78.901
R502 Q.n2 Q.n1 76.002
R503 Q.n7 Q.n4 76
R504 Q.n0 Q.t1 14.282
R505 Q.n0 Q.t0 14.282
R506 Q.n1 Q.t3 14.282
R507 Q.n1 Q.t4 14.282
R508 Q.n2 Q.n0 12.85
R509 Q.n7 Q 0.046
R510 a_1845_1050.n0 a_1845_1050.t6 480.392
R511 a_1845_1050.n0 a_1845_1050.t7 403.272
R512 a_1845_1050.n1 a_1845_1050.t5 283.48
R513 a_1845_1050.n6 a_1845_1050.n5 210.592
R514 a_1845_1050.n6 a_1845_1050.n1 153.315
R515 a_1845_1050.n8 a_1845_1050.n6 152.499
R516 a_1845_1050.n1 a_1845_1050.n0 98.447
R517 a_1845_1050.n8 a_1845_1050.n7 76.002
R518 a_1845_1050.n5 a_1845_1050.n4 30
R519 a_1845_1050.n3 a_1845_1050.n2 24.383
R520 a_1845_1050.n5 a_1845_1050.n3 23.684
R521 a_1845_1050.n7 a_1845_1050.t3 14.282
R522 a_1845_1050.n7 a_1845_1050.t4 14.282
R523 a_1845_1050.t1 a_1845_1050.n9 14.282
R524 a_1845_1050.n9 a_1845_1050.t0 14.282
R525 a_1845_1050.n9 a_1845_1050.n8 12.848
R526 a_1074_101.n12 a_1074_101.n11 26.811
R527 a_1074_101.n6 a_1074_101.n5 24.977
R528 a_1074_101.n2 a_1074_101.n1 24.877
R529 a_1074_101.t0 a_1074_101.n2 12.677
R530 a_1074_101.t0 a_1074_101.n3 11.595
R531 a_1074_101.t1 a_1074_101.n8 8.137
R532 a_1074_101.t0 a_1074_101.n4 7.273
R533 a_1074_101.t0 a_1074_101.n0 6.109
R534 a_1074_101.t1 a_1074_101.n7 4.864
R535 a_1074_101.t0 a_1074_101.n12 2.074
R536 a_1074_101.n7 a_1074_101.n6 1.13
R537 a_1074_101.n12 a_1074_101.t1 0.937
R538 a_1074_101.t1 a_1074_101.n10 0.804
R539 a_1074_101.n10 a_1074_101.n9 0.136
R540 a_277_1050.n4 a_277_1050.t8 480.392
R541 a_277_1050.n2 a_277_1050.t9 480.392
R542 a_277_1050.n4 a_277_1050.t11 403.272
R543 a_277_1050.n2 a_277_1050.t7 403.272
R544 a_277_1050.n5 a_277_1050.t10 310.033
R545 a_277_1050.n3 a_277_1050.t12 310.033
R546 a_277_1050.n11 a_277_1050.n10 239.657
R547 a_277_1050.n12 a_277_1050.n11 144.246
R548 a_277_1050.n6 a_277_1050.n3 83.3
R549 a_277_1050.n14 a_277_1050.n13 79.231
R550 a_277_1050.n11 a_277_1050.n6 77.315
R551 a_277_1050.n6 a_277_1050.n5 76
R552 a_277_1050.n5 a_277_1050.n4 71.894
R553 a_277_1050.n3 a_277_1050.n2 71.894
R554 a_277_1050.n13 a_277_1050.n12 63.152
R555 a_277_1050.n10 a_277_1050.n9 30
R556 a_277_1050.n8 a_277_1050.n7 24.383
R557 a_277_1050.n10 a_277_1050.n8 23.684
R558 a_277_1050.n12 a_277_1050.n1 16.08
R559 a_277_1050.n13 a_277_1050.n0 16.08
R560 a_277_1050.n1 a_277_1050.t5 14.282
R561 a_277_1050.n1 a_277_1050.t4 14.282
R562 a_277_1050.n0 a_277_1050.t2 14.282
R563 a_277_1050.n0 a_277_1050.t6 14.282
R564 a_277_1050.t1 a_277_1050.n14 14.282
R565 a_277_1050.n14 a_277_1050.t0 14.282
R566 a_3177_1050.n1 a_3177_1050.t7 480.392
R567 a_3177_1050.n1 a_3177_1050.t5 403.272
R568 a_3177_1050.n2 a_3177_1050.t6 283.48
R569 a_3177_1050.n7 a_3177_1050.n6 210.592
R570 a_3177_1050.n7 a_3177_1050.n2 153.315
R571 a_3177_1050.n8 a_3177_1050.n7 152.499
R572 a_3177_1050.n2 a_3177_1050.n1 98.447
R573 a_3177_1050.n9 a_3177_1050.n8 76.001
R574 a_3177_1050.n6 a_3177_1050.n5 30
R575 a_3177_1050.n4 a_3177_1050.n3 24.383
R576 a_3177_1050.n6 a_3177_1050.n4 23.684
R577 a_3177_1050.n0 a_3177_1050.t2 14.282
R578 a_3177_1050.n0 a_3177_1050.t3 14.282
R579 a_3177_1050.n9 a_3177_1050.t0 14.282
R580 a_3177_1050.t1 a_3177_1050.n9 14.282
R581 a_3177_1050.n8 a_3177_1050.n0 12.85
R582 a_372_210.n10 a_372_210.n8 82.852
R583 a_372_210.n11 a_372_210.n0 49.6
R584 a_372_210.n7 a_372_210.n6 32.833
R585 a_372_210.n8 a_372_210.t1 32.416
R586 a_372_210.n10 a_372_210.n9 27.2
R587 a_372_210.n3 a_372_210.n2 23.284
R588 a_372_210.n11 a_372_210.n10 22.4
R589 a_372_210.n7 a_372_210.n4 19.017
R590 a_372_210.n6 a_372_210.n5 13.494
R591 a_372_210.t1 a_372_210.n1 7.04
R592 a_372_210.t1 a_372_210.n3 5.727
R593 a_372_210.n8 a_372_210.n7 1.435
R594 a_2406_101.n10 a_2406_101.n9 93.333
R595 a_2406_101.n2 a_2406_101.n1 41.622
R596 a_2406_101.n13 a_2406_101.n12 26.667
R597 a_2406_101.n6 a_2406_101.n5 24.977
R598 a_2406_101.t0 a_2406_101.n2 21.209
R599 a_2406_101.t0 a_2406_101.n3 11.595
R600 a_2406_101.t1 a_2406_101.n8 8.137
R601 a_2406_101.t0 a_2406_101.n0 6.109
R602 a_2406_101.t1 a_2406_101.n7 4.864
R603 a_2406_101.t0 a_2406_101.n4 3.871
R604 a_2406_101.t0 a_2406_101.n13 2.535
R605 a_2406_101.n13 a_2406_101.t1 1.145
R606 a_2406_101.n7 a_2406_101.n6 1.13
R607 a_2406_101.t1 a_2406_101.n11 0.804
R608 a_2406_101.n11 a_2406_101.n10 0.136
R609 GND.n26 GND.n24 219.745
R610 GND.n141 GND.n140 219.745
R611 GND.n171 GND.n169 219.745
R612 GND.n89 GND.n87 219.745
R613 GND.n59 GND.n58 219.745
R614 GND.n26 GND.n25 85.529
R615 GND.n141 GND.n139 85.529
R616 GND.n171 GND.n170 85.529
R617 GND.n89 GND.n88 85.529
R618 GND.n59 GND.n57 85.529
R619 GND.n14 GND.n13 84.842
R620 GND.n77 GND.n76 84.842
R621 GND.n149 GND.n148 84.842
R622 GND.n99 GND.n98 76
R623 GND.n12 GND.n11 76
R624 GND.n17 GND.n16 76
R625 GND.n20 GND.n19 76
R626 GND.n23 GND.n22 76
R627 GND.n30 GND.n29 76
R628 GND.n33 GND.n32 76
R629 GND.n36 GND.n35 76
R630 GND.n39 GND.n38 76
R631 GND.n42 GND.n41 76
R632 GND.n50 GND.n49 76
R633 GND.n53 GND.n52 76
R634 GND.n56 GND.n55 76
R635 GND.n63 GND.n62 76
R636 GND.n66 GND.n65 76
R637 GND.n69 GND.n68 76
R638 GND.n72 GND.n71 76
R639 GND.n75 GND.n74 76
R640 GND.n80 GND.n79 76
R641 GND.n83 GND.n82 76
R642 GND.n86 GND.n85 76
R643 GND.n93 GND.n92 76
R644 GND.n96 GND.n95 76
R645 GND.n194 GND.n193 76
R646 GND.n191 GND.n190 76
R647 GND.n188 GND.n187 76
R648 GND.n185 GND.n184 76
R649 GND.n177 GND.n176 76
R650 GND.n174 GND.n173 76
R651 GND.n167 GND.n166 76
R652 GND.n164 GND.n163 76
R653 GND.n161 GND.n160 76
R654 GND.n158 GND.n157 76
R655 GND.n155 GND.n154 76
R656 GND.n152 GND.n151 76
R657 GND.n147 GND.n146 76
R658 GND.n144 GND.n143 76
R659 GND.n137 GND.n136 76
R660 GND.n134 GND.n133 76
R661 GND.n131 GND.n130 76
R662 GND.n128 GND.n127 76
R663 GND.n125 GND.n124 76
R664 GND.n122 GND.n121 76
R665 GND.n119 GND.n118 76
R666 GND.n116 GND.n115 76
R667 GND.n113 GND.n112 76
R668 GND.n110 GND.n109 76
R669 GND.n102 GND.n101 76
R670 GND.n108 GND.n107 64.552
R671 GND.n47 GND.n46 63.835
R672 GND.n182 GND.n181 63.835
R673 GND.n8 GND.n7 34.942
R674 GND.n46 GND.n45 28.421
R675 GND.n181 GND.n180 28.421
R676 GND.n107 GND.n106 28.421
R677 GND.n46 GND.n44 25.263
R678 GND.n181 GND.n179 25.263
R679 GND.n107 GND.n105 25.263
R680 GND.n44 GND.n43 24.383
R681 GND.n179 GND.n178 24.383
R682 GND.n105 GND.n104 24.383
R683 GND.n6 GND.n5 14.167
R684 GND.n5 GND.n4 14.167
R685 GND.n29 GND.n27 14.167
R686 GND.n62 GND.n60 14.167
R687 GND.n92 GND.n90 14.167
R688 GND.n173 GND.n172 14.167
R689 GND.n143 GND.n142 14.167
R690 GND.n101 GND.n100 13.653
R691 GND.n109 GND.n103 13.653
R692 GND.n112 GND.n111 13.653
R693 GND.n115 GND.n114 13.653
R694 GND.n118 GND.n117 13.653
R695 GND.n121 GND.n120 13.653
R696 GND.n124 GND.n123 13.653
R697 GND.n127 GND.n126 13.653
R698 GND.n130 GND.n129 13.653
R699 GND.n133 GND.n132 13.653
R700 GND.n136 GND.n135 13.653
R701 GND.n143 GND.n138 13.653
R702 GND.n146 GND.n145 13.653
R703 GND.n151 GND.n150 13.653
R704 GND.n154 GND.n153 13.653
R705 GND.n157 GND.n156 13.653
R706 GND.n160 GND.n159 13.653
R707 GND.n163 GND.n162 13.653
R708 GND.n166 GND.n165 13.653
R709 GND.n173 GND.n168 13.653
R710 GND.n176 GND.n175 13.653
R711 GND.n184 GND.n183 13.653
R712 GND.n187 GND.n186 13.653
R713 GND.n190 GND.n189 13.653
R714 GND.n193 GND.n192 13.653
R715 GND.n95 GND.n94 13.653
R716 GND.n92 GND.n91 13.653
R717 GND.n85 GND.n84 13.653
R718 GND.n82 GND.n81 13.653
R719 GND.n79 GND.n78 13.653
R720 GND.n74 GND.n73 13.653
R721 GND.n71 GND.n70 13.653
R722 GND.n68 GND.n67 13.653
R723 GND.n65 GND.n64 13.653
R724 GND.n62 GND.n61 13.653
R725 GND.n55 GND.n54 13.653
R726 GND.n52 GND.n51 13.653
R727 GND.n49 GND.n48 13.653
R728 GND.n41 GND.n40 13.653
R729 GND.n38 GND.n37 13.653
R730 GND.n35 GND.n34 13.653
R731 GND.n32 GND.n31 13.653
R732 GND.n29 GND.n28 13.653
R733 GND.n22 GND.n21 13.653
R734 GND.n19 GND.n18 13.653
R735 GND.n16 GND.n15 13.653
R736 GND.n11 GND.n10 13.653
R737 GND.n4 GND.n3 13.653
R738 GND.n5 GND.n2 13.653
R739 GND.n6 GND.n1 13.653
R740 GND.n27 GND.n26 7.312
R741 GND.n142 GND.n141 7.312
R742 GND.n172 GND.n171 7.312
R743 GND.n90 GND.n89 7.312
R744 GND.n60 GND.n59 7.312
R745 GND.n7 GND.n0 7.083
R746 GND.n7 GND.n6 6.474
R747 GND.n16 GND.n14 3.935
R748 GND.n49 GND.n47 3.935
R749 GND.n79 GND.n77 3.935
R750 GND.n184 GND.n182 3.935
R751 GND.n151 GND.n149 3.935
R752 GND.n98 GND.n97 0.596
R753 GND.n30 GND.n23 0.29
R754 GND.n63 GND.n56 0.29
R755 GND.n93 GND.n86 0.29
R756 GND.n174 GND.n167 0.29
R757 GND.n144 GND.n137 0.29
R758 GND.n99 GND 0.207
R759 GND.n122 GND.n119 0.197
R760 GND.n109 GND.n108 0.196
R761 GND.n12 GND.n9 0.181
R762 GND.n42 GND.n39 0.181
R763 GND.n75 GND.n72 0.181
R764 GND.n191 GND.n188 0.181
R765 GND.n158 GND.n155 0.181
R766 GND.n9 GND.n8 0.145
R767 GND.n17 GND.n12 0.145
R768 GND.n20 GND.n17 0.145
R769 GND.n23 GND.n20 0.145
R770 GND.n33 GND.n30 0.145
R771 GND.n36 GND.n33 0.145
R772 GND.n39 GND.n36 0.145
R773 GND.n50 GND.n42 0.145
R774 GND.n53 GND.n50 0.145
R775 GND.n56 GND.n53 0.145
R776 GND.n66 GND.n63 0.145
R777 GND.n69 GND.n66 0.145
R778 GND.n72 GND.n69 0.145
R779 GND.n80 GND.n75 0.145
R780 GND.n83 GND.n80 0.145
R781 GND.n86 GND.n83 0.145
R782 GND.n96 GND.n93 0.145
R783 GND.n194 GND.n191 0.145
R784 GND.n188 GND.n185 0.145
R785 GND.n185 GND.n177 0.145
R786 GND.n177 GND.n174 0.145
R787 GND.n167 GND.n164 0.145
R788 GND.n164 GND.n161 0.145
R789 GND.n161 GND.n158 0.145
R790 GND.n155 GND.n152 0.145
R791 GND.n152 GND.n147 0.145
R792 GND.n147 GND.n144 0.145
R793 GND.n137 GND.n134 0.145
R794 GND.n134 GND.n131 0.145
R795 GND.n131 GND.n128 0.145
R796 GND.n128 GND.n125 0.145
R797 GND.n125 GND.n122 0.145
R798 GND.n119 GND.n116 0.145
R799 GND.n116 GND.n113 0.145
R800 GND.n113 GND.n110 0.145
R801 GND.n110 GND.n102 0.145
R802 GND.n102 GND.n99 0.145
R803 GND GND.n194 0.137
R804 GND GND.n96 0.008
R805 CLK.n0 CLK.t1 472.359
R806 CLK.n2 CLK.t0 459.505
R807 CLK.n2 CLK.t4 384.527
R808 CLK.n0 CLK.t5 384.527
R809 CLK.n3 CLK.t2 322.152
R810 CLK.n1 CLK.t3 321.724
R811 CLK.n4 CLK.n3 49.342
R812 CLK.n4 CLK.n1 44.933
R813 CLK.n3 CLK.n2 27.599
R814 CLK.n1 CLK.n0 23.329
R815 CLK.n4 CLK 0.046
R816 a_3072_101.n12 a_3072_101.n11 26.811
R817 a_3072_101.n6 a_3072_101.n5 24.977
R818 a_3072_101.n2 a_3072_101.n1 24.877
R819 a_3072_101.t0 a_3072_101.n2 12.677
R820 a_3072_101.t0 a_3072_101.n3 11.595
R821 a_3072_101.t1 a_3072_101.n8 8.137
R822 a_3072_101.t0 a_3072_101.n4 7.273
R823 a_3072_101.t0 a_3072_101.n0 6.109
R824 a_3072_101.t1 a_3072_101.n7 4.864
R825 a_3072_101.t0 a_3072_101.n12 2.074
R826 a_3072_101.n7 a_3072_101.n6 1.13
R827 a_3072_101.n12 a_3072_101.t1 0.937
R828 a_3072_101.t1 a_3072_101.n10 0.804
R829 a_3072_101.n10 a_3072_101.n9 0.136
R830 a_91_103.n5 a_91_103.n4 19.724
R831 a_91_103.t0 a_91_103.n3 11.595
R832 a_91_103.t0 a_91_103.n5 9.207
R833 a_91_103.n2 a_91_103.n1 2.455
R834 a_91_103.n2 a_91_103.n0 1.32
R835 a_91_103.t0 a_91_103.n2 0.246
R836 a_1740_101.t0 a_1740_101.n1 34.62
R837 a_1740_101.t0 a_1740_101.n0 8.137
R838 a_1740_101.t0 a_1740_101.n2 4.69
C4 VDD GND 16.41fF
C5 a_1740_101.n0 GND 0.05fF
C6 a_1740_101.n1 GND 0.12fF
C7 a_1740_101.n2 GND 0.04fF
C8 a_91_103.n0 GND 0.10fF
C9 a_91_103.n1 GND 0.04fF
C10 a_91_103.n2 GND 0.03fF
C11 a_91_103.n3 GND 0.06fF
C12 a_91_103.n4 GND 0.08fF
C13 a_91_103.n5 GND 0.06fF
C14 a_3072_101.n0 GND 0.02fF
C15 a_3072_101.n1 GND 0.10fF
C16 a_3072_101.n2 GND 0.06fF
C17 a_3072_101.n3 GND 0.06fF
C18 a_3072_101.n4 GND 0.00fF
C19 a_3072_101.n5 GND 0.04fF
C20 a_3072_101.n6 GND 0.05fF
C21 a_3072_101.n7 GND 0.02fF
C22 a_3072_101.n8 GND 0.05fF
C23 a_3072_101.n9 GND 0.08fF
C24 a_3072_101.n10 GND 0.17fF
C25 a_3072_101.t1 GND 0.23fF
C26 a_3072_101.n11 GND 0.09fF
C27 a_3072_101.n12 GND 0.00fF
C28 a_2406_101.n0 GND 0.02fF
C29 a_2406_101.n1 GND 0.10fF
C30 a_2406_101.n2 GND 0.07fF
C31 a_2406_101.n3 GND 0.05fF
C32 a_2406_101.n4 GND 0.00fF
C33 a_2406_101.n5 GND 0.04fF
C34 a_2406_101.n6 GND 0.05fF
C35 a_2406_101.n7 GND 0.02fF
C36 a_2406_101.n8 GND 0.05fF
C37 a_2406_101.n9 GND 0.02fF
C38 a_2406_101.n10 GND 0.08fF
C39 a_2406_101.n11 GND 0.17fF
C40 a_2406_101.t1 GND 0.23fF
C41 a_2406_101.n12 GND 0.09fF
C42 a_2406_101.n13 GND 0.00fF
C43 a_372_210.n0 GND 0.02fF
C44 a_372_210.n1 GND 0.09fF
C45 a_372_210.n2 GND 0.13fF
C46 a_372_210.n3 GND 0.11fF
C47 a_372_210.t1 GND 0.30fF
C48 a_372_210.n4 GND 0.09fF
C49 a_372_210.n5 GND 0.06fF
C50 a_372_210.n6 GND 0.01fF
C51 a_372_210.n7 GND 0.03fF
C52 a_372_210.n8 GND 0.11fF
C53 a_372_210.n9 GND 0.02fF
C54 a_372_210.n10 GND 0.05fF
C55 a_372_210.n11 GND 0.02fF
C56 a_3177_1050.n0 GND 0.50fF
C57 a_3177_1050.n1 GND 0.36fF
C58 a_3177_1050.n2 GND 0.54fF
C59 a_3177_1050.n3 GND 0.04fF
C60 a_3177_1050.n4 GND 0.05fF
C61 a_3177_1050.n5 GND 0.03fF
C62 a_3177_1050.n6 GND 0.28fF
C63 a_3177_1050.n7 GND 0.57fF
C64 a_3177_1050.n8 GND 0.29fF
C65 a_3177_1050.n9 GND 0.59fF
C66 a_277_1050.n0 GND 0.69fF
C67 a_277_1050.n1 GND 0.69fF
C68 a_277_1050.n2 GND 0.44fF
C69 a_277_1050.n3 GND 0.61fF
C70 a_277_1050.n4 GND 0.44fF
C71 a_277_1050.n5 GND 0.51fF
C72 a_277_1050.n6 GND 2.48fF
C73 a_277_1050.n7 GND 0.05fF
C74 a_277_1050.n8 GND 0.07fF
C75 a_277_1050.n9 GND 0.04fF
C76 a_277_1050.n10 GND 0.43fF
C77 a_277_1050.n11 GND 0.58fF
C78 a_277_1050.n12 GND 0.36fF
C79 a_277_1050.n13 GND 0.26fF
C80 a_277_1050.n14 GND 0.81fF
C81 a_1074_101.n0 GND 0.02fF
C82 a_1074_101.n1 GND 0.10fF
C83 a_1074_101.n2 GND 0.06fF
C84 a_1074_101.n3 GND 0.06fF
C85 a_1074_101.n4 GND 0.00fF
C86 a_1074_101.n5 GND 0.04fF
C87 a_1074_101.n6 GND 0.05fF
C88 a_1074_101.n7 GND 0.02fF
C89 a_1074_101.n8 GND 0.05fF
C90 a_1074_101.n9 GND 0.08fF
C91 a_1074_101.n10 GND 0.17fF
C92 a_1074_101.t1 GND 0.23fF
C93 a_1074_101.n11 GND 0.09fF
C94 a_1074_101.n12 GND 0.00fF
C95 a_1845_1050.n0 GND 0.37fF
C96 a_1845_1050.n1 GND 0.56fF
C97 a_1845_1050.n2 GND 0.04fF
C98 a_1845_1050.n3 GND 0.05fF
C99 a_1845_1050.n4 GND 0.03fF
C100 a_1845_1050.n5 GND 0.29fF
C101 a_1845_1050.n6 GND 0.60fF
C102 a_1845_1050.n7 GND 0.62fF
C103 a_1845_1050.n8 GND 0.30fF
C104 a_1845_1050.n9 GND 0.52fF
C105 Q.n0 GND 0.56fF
C106 Q.n1 GND 0.66fF
C107 Q.n2 GND 0.29fF
C108 Q.n3 GND 0.45fF
C109 Q.n4 GND 0.48fF
C110 Q.n5 GND 0.32fF
C111 Q.t5 GND 0.59fF
C112 Q.n6 GND 0.41fF
C113 Q.n7 GND 0.03fF
C114 a_3738_101.n0 GND 0.07fF
C115 a_3738_101.n1 GND 0.02fF
C116 a_3738_101.n2 GND 0.01fF
C117 a_3738_101.n3 GND 0.06fF
C118 a_3738_101.n4 GND 0.10fF
C119 a_3738_101.n5 GND 0.06fF
C120 a_3738_101.n6 GND 0.05fF
C121 a_147_187.n0 GND 0.05fF
C122 a_147_187.n1 GND 0.72fF
C123 a_147_187.n2 GND 0.85fF
C124 a_147_187.n3 GND 0.33fF
C125 a_147_187.n4 GND 0.38fF
C126 a_147_187.n5 GND 0.56fF
C127 a_147_187.n6 GND 0.38fF
C128 a_147_187.t13 GND 0.80fF
C129 a_147_187.n7 GND 0.52fF
C130 a_147_187.n8 GND 0.37fF
C131 a_147_187.n9 GND 0.74fF
C132 a_147_187.n10 GND 2.40fF
C133 a_147_187.n11 GND 1.79fF
C134 a_147_187.n12 GND 0.58fF
C135 a_147_187.n13 GND 0.05fF
C136 a_147_187.n14 GND 0.49fF
C137 a_147_187.n15 GND 0.07fF
C138 a_599_989.n0 GND 0.40fF
C139 a_599_989.n1 GND 0.42fF
C140 a_599_989.n2 GND 0.40fF
C141 a_599_989.t6 GND 0.56fF
C142 a_599_989.n3 GND 0.40fF
C143 a_599_989.n4 GND 1.08fF
C144 a_599_989.n5 GND 0.04fF
C145 a_599_989.n6 GND 0.06fF
C146 a_599_989.n7 GND 0.04fF
C147 a_599_989.n8 GND 0.32fF
C148 a_599_989.n9 GND 0.45fF
C149 a_599_989.n10 GND 0.67fF
C150 a_599_989.n11 GND 0.33fF
C151 a_599_989.n12 GND 0.56fF
C152 VDD.n0 GND 0.16fF
C153 VDD.n1 GND 0.03fF
C154 VDD.n2 GND 0.02fF
C155 VDD.n3 GND 0.05fF
C156 VDD.n4 GND 0.01fF
C157 VDD.n6 GND 0.02fF
C158 VDD.n7 GND 0.02fF
C159 VDD.n9 GND 0.02fF
C160 VDD.n10 GND 0.02fF
C161 VDD.n11 GND 0.02fF
C162 VDD.n14 GND 0.46fF
C163 VDD.n16 GND 0.03fF
C164 VDD.n17 GND 0.02fF
C165 VDD.n18 GND 0.02fF
C166 VDD.n19 GND 0.02fF
C167 VDD.n20 GND 0.04fF
C168 VDD.n21 GND 0.28fF
C169 VDD.n22 GND 0.02fF
C170 VDD.n23 GND 0.03fF
C171 VDD.n24 GND 0.14fF
C172 VDD.n25 GND 0.17fF
C173 VDD.n26 GND 0.01fF
C174 VDD.n27 GND 0.11fF
C175 VDD.n28 GND 0.03fF
C176 VDD.n29 GND 0.31fF
C177 VDD.n30 GND 0.01fF
C178 VDD.n31 GND 0.02fF
C179 VDD.n32 GND 0.02fF
C180 VDD.n33 GND 0.06fF
C181 VDD.n34 GND 0.25fF
C182 VDD.n35 GND 0.01fF
C183 VDD.n36 GND 0.01fF
C184 VDD.n37 GND 0.00fF
C185 VDD.n38 GND 0.09fF
C186 VDD.n39 GND 0.03fF
C187 VDD.n40 GND 0.17fF
C188 VDD.n41 GND 0.14fF
C189 VDD.n42 GND 0.01fF
C190 VDD.n43 GND 0.02fF
C191 VDD.n44 GND 0.03fF
C192 VDD.n45 GND 0.14fF
C193 VDD.n46 GND 0.17fF
C194 VDD.n47 GND 0.01fF
C195 VDD.n48 GND 0.02fF
C196 VDD.n49 GND 0.02fF
C197 VDD.n50 GND 0.06fF
C198 VDD.n51 GND 0.25fF
C199 VDD.n52 GND 0.01fF
C200 VDD.n53 GND 0.01fF
C201 VDD.n54 GND 0.02fF
C202 VDD.n55 GND 0.28fF
C203 VDD.n56 GND 0.01fF
C204 VDD.n57 GND 0.02fF
C205 VDD.n58 GND 0.03fF
C206 VDD.n59 GND 0.02fF
C207 VDD.n60 GND 0.02fF
C208 VDD.n61 GND 0.02fF
C209 VDD.n62 GND 0.22fF
C210 VDD.n63 GND 0.04fF
C211 VDD.n64 GND 0.04fF
C212 VDD.n65 GND 0.02fF
C213 VDD.n67 GND 0.02fF
C214 VDD.n68 GND 0.02fF
C215 VDD.n69 GND 0.02fF
C216 VDD.n70 GND 0.02fF
C217 VDD.n72 GND 0.02fF
C218 VDD.n73 GND 0.02fF
C219 VDD.n74 GND 0.02fF
C220 VDD.n76 GND 0.28fF
C221 VDD.n78 GND 0.02fF
C222 VDD.n79 GND 0.02fF
C223 VDD.n80 GND 0.03fF
C224 VDD.n81 GND 0.02fF
C225 VDD.n82 GND 0.28fF
C226 VDD.n83 GND 0.01fF
C227 VDD.n84 GND 0.02fF
C228 VDD.n85 GND 0.03fF
C229 VDD.n86 GND 0.06fF
C230 VDD.n87 GND 0.25fF
C231 VDD.n88 GND 0.01fF
C232 VDD.n89 GND 0.01fF
C233 VDD.n90 GND 0.02fF
C234 VDD.n91 GND 0.14fF
C235 VDD.n92 GND 0.17fF
C236 VDD.n93 GND 0.01fF
C237 VDD.n94 GND 0.02fF
C238 VDD.n95 GND 0.02fF
C239 VDD.n96 GND 0.11fF
C240 VDD.n97 GND 0.03fF
C241 VDD.n98 GND 0.31fF
C242 VDD.n99 GND 0.01fF
C243 VDD.n100 GND 0.02fF
C244 VDD.n101 GND 0.03fF
C245 VDD.n102 GND 0.17fF
C246 VDD.n103 GND 0.14fF
C247 VDD.n104 GND 0.01fF
C248 VDD.n105 GND 0.02fF
C249 VDD.n106 GND 0.03fF
C250 VDD.n107 GND 0.14fF
C251 VDD.n108 GND 0.17fF
C252 VDD.n109 GND 0.01fF
C253 VDD.n110 GND 0.02fF
C254 VDD.n111 GND 0.02fF
C255 VDD.n112 GND 0.06fF
C256 VDD.n113 GND 0.25fF
C257 VDD.n114 GND 0.01fF
C258 VDD.n115 GND 0.01fF
C259 VDD.n116 GND 0.02fF
C260 VDD.n117 GND 0.28fF
C261 VDD.n118 GND 0.01fF
C262 VDD.n119 GND 0.02fF
C263 VDD.n120 GND 0.03fF
C264 VDD.n121 GND 0.02fF
C265 VDD.n122 GND 0.02fF
C266 VDD.n123 GND 0.02fF
C267 VDD.n124 GND 0.22fF
C268 VDD.n125 GND 0.04fF
C269 VDD.n126 GND 0.03fF
C270 VDD.n127 GND 0.02fF
C271 VDD.n128 GND 0.02fF
C272 VDD.n129 GND 0.02fF
C273 VDD.n130 GND 0.03fF
C274 VDD.n131 GND 0.02fF
C275 VDD.n133 GND 0.02fF
C276 VDD.n134 GND 0.02fF
C277 VDD.n135 GND 0.02fF
C278 VDD.n137 GND 0.28fF
C279 VDD.n139 GND 0.02fF
C280 VDD.n140 GND 0.02fF
C281 VDD.n141 GND 0.03fF
C282 VDD.n142 GND 0.02fF
C283 VDD.n143 GND 0.28fF
C284 VDD.n144 GND 0.01fF
C285 VDD.n145 GND 0.02fF
C286 VDD.n146 GND 0.03fF
C287 VDD.n147 GND 0.06fF
C288 VDD.n148 GND 0.25fF
C289 VDD.n149 GND 0.01fF
C290 VDD.n150 GND 0.01fF
C291 VDD.n151 GND 0.02fF
C292 VDD.n152 GND 0.14fF
C293 VDD.n153 GND 0.17fF
C294 VDD.n154 GND 0.01fF
C295 VDD.n155 GND 0.02fF
C296 VDD.n156 GND 0.02fF
C297 VDD.n157 GND 0.11fF
C298 VDD.n158 GND 0.03fF
C299 VDD.n159 GND 0.31fF
C300 VDD.n160 GND 0.01fF
C301 VDD.n161 GND 0.02fF
C302 VDD.n162 GND 0.03fF
C303 VDD.n163 GND 0.17fF
C304 VDD.n164 GND 0.14fF
C305 VDD.n165 GND 0.01fF
C306 VDD.n166 GND 0.02fF
C307 VDD.n167 GND 0.03fF
C308 VDD.n168 GND 0.14fF
C309 VDD.n169 GND 0.17fF
C310 VDD.n170 GND 0.01fF
C311 VDD.n171 GND 0.02fF
C312 VDD.n172 GND 0.02fF
C313 VDD.n173 GND 0.06fF
C314 VDD.n174 GND 0.25fF
C315 VDD.n175 GND 0.01fF
C316 VDD.n176 GND 0.01fF
C317 VDD.n177 GND 0.02fF
C318 VDD.n178 GND 0.28fF
C319 VDD.n179 GND 0.01fF
C320 VDD.n180 GND 0.02fF
C321 VDD.n181 GND 0.03fF
C322 VDD.n182 GND 0.02fF
C323 VDD.n183 GND 0.02fF
C324 VDD.n184 GND 0.02fF
C325 VDD.n185 GND 0.22fF
C326 VDD.n186 GND 0.04fF
C327 VDD.n187 GND 0.03fF
C328 VDD.n188 GND 0.02fF
C329 VDD.n189 GND 0.02fF
C330 VDD.n190 GND 0.02fF
C331 VDD.n191 GND 0.03fF
C332 VDD.n192 GND 0.02fF
C333 VDD.n194 GND 0.02fF
C334 VDD.n195 GND 0.02fF
C335 VDD.n196 GND 0.02fF
C336 VDD.n198 GND 0.28fF
C337 VDD.n200 GND 0.02fF
C338 VDD.n201 GND 0.02fF
C339 VDD.n202 GND 0.03fF
C340 VDD.n203 GND 0.02fF
C341 VDD.n204 GND 0.28fF
C342 VDD.n205 GND 0.01fF
C343 VDD.n206 GND 0.02fF
C344 VDD.n207 GND 0.03fF
C345 VDD.n208 GND 0.06fF
C346 VDD.n209 GND 0.25fF
C347 VDD.n210 GND 0.01fF
C348 VDD.n211 GND 0.01fF
C349 VDD.n212 GND 0.01fF
C350 VDD.n213 GND 0.02fF
C351 VDD.n214 GND 0.02fF
C352 VDD.n215 GND 0.02fF
C353 VDD.n216 GND 0.20fF
C354 VDD.n217 GND 0.03fF
C355 VDD.n218 GND 0.02fF
C356 VDD.n219 GND 0.02fF
C357 VDD.n220 GND 0.02fF
C358 VDD.n221 GND 0.03fF
C359 VDD.n222 GND 0.02fF
C360 VDD.n224 GND 0.02fF
C361 VDD.n225 GND 0.02fF
C362 VDD.n226 GND 0.02fF
C363 VDD.n228 GND 0.46fF
C364 VDD.n230 GND 0.03fF
C365 VDD.n231 GND 0.04fF
C366 VDD.n232 GND 0.28fF
C367 VDD.n233 GND 0.02fF
C368 VDD.n234 GND 0.03fF
C369 VDD.n235 GND 0.03fF
C370 VDD.n236 GND 0.28fF
C371 VDD.n237 GND 0.01fF
C372 VDD.n238 GND 0.02fF
C373 VDD.n239 GND 0.02fF
C374 VDD.n240 GND 0.06fF
C375 VDD.n241 GND 0.23fF
C376 VDD.n242 GND 0.01fF
C377 VDD.n243 GND 0.01fF
C378 VDD.n244 GND 0.02fF
C379 VDD.n245 GND 0.14fF
C380 VDD.n246 GND 0.17fF
C381 VDD.n247 GND 0.01fF
C382 VDD.n248 GND 0.02fF
C383 VDD.n249 GND 0.02fF
C384 VDD.n250 GND 0.11fF
C385 VDD.n251 GND 0.02fF
C386 VDD.n252 GND 0.14fF
C387 VDD.n253 GND 0.16fF
C388 VDD.n254 GND 0.01fF
C389 VDD.n255 GND 0.02fF
C390 VDD.n256 GND 0.02fF
C391 VDD.n257 GND 0.18fF
C392 VDD.n258 GND 0.15fF
C393 VDD.n259 GND 0.01fF
C394 VDD.n260 GND 0.02fF
C395 VDD.n261 GND 0.03fF
C396 VDD.n262 GND 0.18fF
C397 VDD.n263 GND 0.15fF
C398 VDD.n264 GND 0.01fF
C399 VDD.n265 GND 0.02fF
C400 VDD.n266 GND 0.03fF
C401 VDD.n267 GND 0.14fF
C402 VDD.n268 GND 0.16fF
C403 VDD.n269 GND 0.01fF
C404 VDD.n270 GND 0.11fF
C405 VDD.n271 GND 0.02fF
C406 VDD.n272 GND 0.02fF
C407 VDD.n273 GND 0.02fF
C408 VDD.n274 GND 0.14fF
C409 VDD.n275 GND 0.17fF
C410 VDD.n276 GND 0.01fF
C411 VDD.n277 GND 0.02fF
C412 VDD.n278 GND 0.02fF
C413 VDD.n279 GND 0.22fF
C414 VDD.n280 GND 0.01fF
C415 VDD.n281 GND 0.07fF
C416 VDD.n282 GND 0.02fF
C417 VDD.n283 GND 0.28fF
C418 VDD.n284 GND 0.01fF
C419 VDD.n285 GND 0.02fF
C420 VDD.n286 GND 0.02fF
C421 VDD.n287 GND 0.28fF
C422 VDD.n288 GND 0.01fF
C423 VDD.n289 GND 0.02fF
C424 VDD.n290 GND 0.03fF
C425 VDD.n291 GND 0.02fF
C426 VDD.n292 GND 0.02fF
C427 VDD.n293 GND 0.02fF
C428 VDD.n294 GND 0.02fF
C429 VDD.n295 GND 0.02fF
C430 VDD.n296 GND 0.02fF
C431 VDD.n298 GND 0.02fF
C432 VDD.n299 GND 0.02fF
C433 VDD.n300 GND 0.02fF
C434 VDD.n301 GND 0.02fF
C435 VDD.n303 GND 0.04fF
C436 VDD.n304 GND 0.02fF
C437 VDD.n305 GND 0.27fF
C438 VDD.n306 GND 0.04fF
C439 VDD.n308 GND 0.28fF
C440 VDD.n310 GND 0.02fF
C441 VDD.n311 GND 0.02fF
C442 VDD.n312 GND 0.03fF
C443 VDD.n313 GND 0.02fF
C444 VDD.n314 GND 0.28fF
C445 VDD.n315 GND 0.01fF
C446 VDD.n316 GND 0.02fF
C447 VDD.n317 GND 0.03fF
C448 VDD.n318 GND 0.06fF
C449 VDD.n319 GND 0.25fF
C450 VDD.n320 GND 0.01fF
C451 VDD.n321 GND 0.01fF
C452 VDD.n322 GND 0.02fF
C453 VDD.n323 GND 0.14fF
C454 VDD.n324 GND 0.17fF
C455 VDD.n325 GND 0.01fF
C456 VDD.n326 GND 0.02fF
C457 VDD.n327 GND 0.02fF
C458 VDD.n328 GND 0.17fF
C459 VDD.n329 GND 0.14fF
C460 VDD.n330 GND 0.01fF
C461 VDD.n331 GND 0.02fF
C462 VDD.n332 GND 0.03fF
C463 VDD.n333 GND 0.11fF
C464 VDD.n334 GND 0.03fF
C465 VDD.n335 GND 0.31fF
C466 VDD.n336 GND 0.01fF
C467 VDD.n337 GND 0.02fF
C468 VDD.n338 GND 0.03fF
C469 VDD.n339 GND 0.14fF
C470 VDD.n340 GND 0.17fF
C471 VDD.n341 GND 0.01fF
C472 VDD.n342 GND 0.02fF
C473 VDD.n343 GND 0.02fF
C474 VDD.n344 GND 0.06fF
C475 VDD.n345 GND 0.25fF
C476 VDD.n346 GND 0.01fF
C477 VDD.n347 GND 0.01fF
C478 VDD.n348 GND 0.02fF
C479 VDD.n349 GND 0.28fF
C480 VDD.n350 GND 0.01fF
C481 VDD.n351 GND 0.02fF
C482 VDD.n352 GND 0.03fF
C483 VDD.n353 GND 0.02fF
C484 VDD.n354 GND 0.02fF
C485 VDD.n355 GND 0.02fF
C486 VDD.n356 GND 0.22fF
C487 VDD.n357 GND 0.04fF
C488 VDD.n358 GND 0.03fF
C489 VDD.n359 GND 0.02fF
C490 VDD.n360 GND 0.02fF
C491 VDD.n361 GND 0.02fF
C492 VDD.n362 GND 0.03fF
C493 VDD.n363 GND 0.02fF
C494 VDD.n365 GND 0.02fF
C495 VDD.n366 GND 0.02fF
C496 VDD.n367 GND 0.02fF
C497 VDD.n369 GND 0.28fF
C498 VDD.n371 GND 0.02fF
C499 VDD.n372 GND 0.02fF
C500 VDD.n373 GND 0.03fF
C501 VDD.n374 GND 0.02fF
C502 VDD.n375 GND 0.28fF
C503 VDD.n376 GND 0.01fF
C504 VDD.n377 GND 0.02fF
C505 VDD.n378 GND 0.03fF
C506 VDD.n379 GND 0.06fF
C507 VDD.n380 GND 0.25fF
C508 VDD.n381 GND 0.01fF
C509 VDD.n382 GND 0.01fF
C510 VDD.n383 GND 0.02fF
C511 VDD.n384 GND 0.14fF
C512 VDD.n385 GND 0.17fF
C513 VDD.n386 GND 0.01fF
C514 VDD.n387 GND 0.02fF
C515 VDD.n388 GND 0.02fF
C516 VDD.n389 GND 0.17fF
C517 VDD.n390 GND 0.14fF
C518 VDD.n391 GND 0.01fF
C519 VDD.n392 GND 0.02fF
C520 VDD.n393 GND 0.03fF
C521 VDD.n394 GND 0.11fF
C522 VDD.n395 GND 0.03fF
C523 VDD.n396 GND 0.31fF
C524 VDD.n397 GND 0.01fF
C525 VDD.n398 GND 0.02fF
C526 VDD.n399 GND 0.03fF
C527 VDD.n400 GND 0.14fF
C528 VDD.n401 GND 0.17fF
C529 VDD.n402 GND 0.01fF
C530 VDD.n403 GND 0.02fF
C531 VDD.n404 GND 0.02fF
.ends
