magic
tech sky130A
magscale 1 2
timestamp 1652455121
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 131 871 165 905
rect 797 871 831 905
rect 1759 871 1793 905
rect 1907 871 1941 905
rect 3165 871 3199 905
rect 3535 871 3569 905
rect 131 797 165 831
rect 1907 797 1941 831
rect 131 723 165 757
rect 797 723 831 757
rect 131 649 165 683
rect 797 649 831 683
rect 1759 649 1793 683
rect 1907 649 1941 683
rect 3165 649 3199 683
rect 3535 649 3569 683
rect 131 575 165 609
rect 797 575 831 609
rect 1759 575 1793 609
rect 1907 575 1941 609
rect 3165 575 3199 609
rect 3535 575 3569 609
rect 131 501 165 535
rect 797 501 831 535
rect 1759 501 1793 535
rect 1907 501 1941 535
rect 3165 501 3199 535
rect 3535 501 3569 535
rect 131 427 165 461
rect 1907 427 1941 461
rect 3165 427 3199 461
rect 3535 427 3569 461
<< metal1 >>
rect -34 1446 4030 1514
rect 201 797 1871 831
rect 2569 797 3647 831
rect 349 723 613 757
rect 1459 723 2833 757
rect 3087 723 3795 757
rect 3235 649 3499 683
rect 867 575 1723 609
rect -34 -34 4030 34
use li1_M1_contact  li1_M1_contact_5 pcells
timestamp 1648061256
transform 1 0 666 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 296 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 814 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 148 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 1406 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 1 0 1924 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 1776 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 3182 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 3552 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 3034 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform -1 0 2516 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 3700 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 2886 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform 1 0 3848 0 1 740
box -53 -33 29 33
use nor2x1_pcell  nor2x1_pcell_0 pcells
timestamp 1652323563
transform 1 0 2664 0 1 0
box -87 -34 753 1550
use nor2x1_pcell  nor2x1_pcell_1
timestamp 1652323563
transform 1 0 3330 0 1 0
box -87 -34 753 1550
use and2x1_pcell  and2x1_pcell_0 pcells
timestamp 1652455121
transform 1 0 444 0 1 0
box -87 -34 1197 1550
use and2x1_pcell  and2x1_pcell_1
timestamp 1652455121
transform 1 0 1554 0 1 0
box -87 -34 1197 1550
use invx1_pcell  invx1_pcell_0 pcells
timestamp 1652329846
transform 1 0 0 0 1 0
box -87 -34 531 1550
<< labels >>
rlabel locali 3165 649 3199 683 1 Q
port 1 nsew signal output
rlabel locali 3165 575 3199 609 1 Q
port 1 nsew signal output
rlabel locali 3165 501 3199 535 1 Q
port 1 nsew signal output
rlabel locali 3165 427 3199 461 1 Q
port 1 nsew signal output
rlabel locali 3165 871 3199 905 1 Q
port 1 nsew signal output
rlabel locali 3535 427 3569 461 1 Q
port 1 nsew signal output
rlabel locali 3535 501 3569 535 1 Q
port 1 nsew signal output
rlabel locali 3535 575 3569 609 1 Q
port 1 nsew signal output
rlabel locali 3535 649 3569 683 1 Q
port 1 nsew signal output
rlabel locali 3535 871 3569 905 1 Q
port 1 nsew signal output
rlabel locali 131 797 165 831 1 D
port 2 nsew signal input
rlabel locali 131 871 165 905 1 D
port 2 nsew signal input
rlabel locali 131 723 165 757 1 D
port 2 nsew signal input
rlabel locali 131 649 165 683 1 D
port 2 nsew signal input
rlabel locali 131 575 165 609 1 D
port 2 nsew signal input
rlabel locali 131 501 165 535 1 D
port 2 nsew signal input
rlabel locali 131 427 165 461 1 D
port 2 nsew signal input
rlabel locali 1907 427 1941 461 1 D
port 2 nsew signal input
rlabel locali 1907 501 1941 535 1 D
port 2 nsew signal input
rlabel locali 1907 575 1941 609 1 D
port 2 nsew signal input
rlabel locali 1907 649 1941 683 1 D
port 2 nsew signal input
rlabel locali 1907 797 1941 831 1 D
port 2 nsew signal input
rlabel locali 1907 871 1941 905 1 D
port 2 nsew signal input
rlabel locali 797 575 831 609 1 GATE
port 3 nsew signal input
rlabel locali 797 501 831 535 1 GATE
port 3 nsew signal input
rlabel locali 797 649 831 683 1 GATE
port 3 nsew signal input
rlabel locali 797 723 831 757 1 GATE
port 3 nsew signal input
rlabel locali 797 871 831 905 1 GATE
port 3 nsew signal input
rlabel locali 1759 501 1793 535 1 GATE
port 3 nsew signal input
rlabel locali 1759 575 1793 609 1 GATE
port 3 nsew signal input
rlabel locali 1759 649 1793 683 1 GATE
port 3 nsew signal input
rlabel locali 1759 871 1793 905 1 GATE
port 3 nsew signal input
rlabel metal1 -34 1446 4030 1514 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 -34 -34 4030 34 1 GND
port 5 nsew ground bidirectional abutment


<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 3996 1480
string LEFsymmetry X Y R90
<< end >>
