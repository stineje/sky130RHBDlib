magic
tech sky130A
magscale 1 2
timestamp 1645210163
use sky130_fd_pr__dfl1sd__example_55959141808123  sky130_fd_pr__dfl1sd__example_55959141808123_0
timestamp 1645210163
transform 1 0 200 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808122  sky130_fd_pr__hvdfl1sd__example_55959141808122_0
timestamp 1645210163
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 228 29 228 29 0 FreeSans 300 0 0 0 D
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 37313126
string GDS_START 37312074
<< end >>
