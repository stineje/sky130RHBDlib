magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 710 203
rect 30 -17 64 21
<< scnmos >>
rect 108 47 138 177
rect 208 47 238 177
rect 316 47 346 177
rect 400 47 430 177
rect 496 47 526 177
rect 592 47 622 177
<< scpmoshvt >>
rect 108 297 138 497
rect 208 297 238 497
rect 316 297 346 497
rect 400 297 430 497
rect 496 297 526 497
rect 611 297 641 497
<< ndiff >>
rect 27 165 108 177
rect 27 131 35 165
rect 69 131 108 165
rect 27 93 108 131
rect 27 59 35 93
rect 69 59 108 93
rect 27 47 108 59
rect 138 157 208 177
rect 138 123 148 157
rect 182 123 208 157
rect 138 89 208 123
rect 138 55 148 89
rect 182 55 208 89
rect 138 47 208 55
rect 238 157 316 177
rect 238 123 260 157
rect 294 123 316 157
rect 238 89 316 123
rect 238 55 260 89
rect 294 55 316 89
rect 238 47 316 55
rect 346 129 400 177
rect 346 95 356 129
rect 390 95 400 129
rect 346 47 400 95
rect 430 89 496 177
rect 430 55 446 89
rect 480 55 496 89
rect 430 47 496 55
rect 526 129 592 177
rect 526 95 542 129
rect 576 95 592 129
rect 526 47 592 95
rect 622 157 684 177
rect 622 123 638 157
rect 672 123 684 157
rect 622 89 684 123
rect 622 55 638 89
rect 672 55 684 89
rect 622 47 684 55
<< pdiff >>
rect 27 485 108 497
rect 27 451 35 485
rect 69 451 108 485
rect 27 414 108 451
rect 27 380 35 414
rect 69 380 108 414
rect 27 343 108 380
rect 27 309 35 343
rect 69 309 108 343
rect 27 297 108 309
rect 138 477 208 497
rect 138 443 148 477
rect 182 443 208 477
rect 138 409 208 443
rect 138 375 148 409
rect 182 375 208 409
rect 138 297 208 375
rect 238 477 316 497
rect 238 443 260 477
rect 294 443 316 477
rect 238 409 316 443
rect 238 375 260 409
rect 294 375 316 409
rect 238 297 316 375
rect 346 297 400 497
rect 430 297 496 497
rect 526 477 611 497
rect 526 443 566 477
rect 600 443 611 477
rect 526 349 611 443
rect 526 315 566 349
rect 600 315 611 349
rect 526 297 611 315
rect 641 477 709 497
rect 641 443 667 477
rect 701 443 709 477
rect 641 409 709 443
rect 641 375 667 409
rect 701 375 709 409
rect 641 297 709 375
<< ndiffc >>
rect 35 131 69 165
rect 35 59 69 93
rect 148 123 182 157
rect 148 55 182 89
rect 260 123 294 157
rect 260 55 294 89
rect 356 95 390 129
rect 446 55 480 89
rect 542 95 576 129
rect 638 123 672 157
rect 638 55 672 89
<< pdiffc >>
rect 35 451 69 485
rect 35 380 69 414
rect 35 309 69 343
rect 148 443 182 477
rect 148 375 182 409
rect 260 443 294 477
rect 260 375 294 409
rect 566 443 600 477
rect 566 315 600 349
rect 667 443 701 477
rect 667 375 701 409
<< poly >>
rect 108 497 138 523
rect 208 497 238 523
rect 316 497 346 523
rect 400 497 430 523
rect 496 497 526 523
rect 611 497 641 523
rect 108 265 138 297
rect 208 265 238 297
rect 316 265 346 297
rect 400 265 430 297
rect 496 265 526 297
rect 611 265 641 297
rect 108 249 250 265
rect 108 215 206 249
rect 240 215 250 249
rect 108 199 250 215
rect 292 249 346 265
rect 292 215 302 249
rect 336 215 346 249
rect 292 199 346 215
rect 388 249 442 265
rect 388 215 398 249
rect 432 215 442 249
rect 388 199 442 215
rect 484 249 538 265
rect 484 215 494 249
rect 528 215 538 249
rect 484 199 538 215
rect 580 249 641 265
rect 580 215 590 249
rect 624 215 641 249
rect 580 199 641 215
rect 108 177 138 199
rect 208 177 238 199
rect 316 177 346 199
rect 400 177 430 199
rect 496 177 526 199
rect 592 177 622 199
rect 108 21 138 47
rect 208 21 238 47
rect 316 21 346 47
rect 400 21 430 47
rect 496 21 526 47
rect 592 21 622 47
<< polycont >>
rect 206 215 240 249
rect 302 215 336 249
rect 398 215 432 249
rect 494 215 528 249
rect 590 215 624 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 485 76 527
rect 17 451 35 485
rect 69 451 76 485
rect 17 414 76 451
rect 17 380 35 414
rect 69 380 76 414
rect 17 343 76 380
rect 17 309 35 343
rect 69 309 76 343
rect 17 293 76 309
rect 110 477 198 493
rect 110 443 148 477
rect 182 443 198 477
rect 110 409 198 443
rect 110 375 148 409
rect 182 375 198 409
rect 110 367 198 375
rect 233 477 296 527
rect 233 443 260 477
rect 294 443 296 477
rect 233 409 296 443
rect 233 375 260 409
rect 294 375 296 409
rect 110 259 172 367
rect 233 357 296 375
rect 330 477 616 493
rect 330 459 566 477
rect 330 323 364 459
rect 600 443 616 477
rect 17 215 172 259
rect 17 165 76 181
rect 17 131 35 165
rect 69 131 76 165
rect 17 93 76 131
rect 17 59 35 93
rect 69 59 76 93
rect 17 17 76 59
rect 110 165 172 215
rect 206 289 364 323
rect 206 249 240 289
rect 398 265 438 425
rect 206 199 240 215
rect 274 249 352 255
rect 274 215 302 249
rect 336 215 352 249
rect 274 199 352 215
rect 389 249 438 265
rect 389 215 398 249
rect 432 215 438 249
rect 389 199 438 215
rect 478 249 528 425
rect 566 349 616 443
rect 651 477 718 527
rect 651 443 667 477
rect 701 443 718 477
rect 651 409 718 443
rect 651 375 667 409
rect 701 375 718 409
rect 651 367 718 375
rect 600 333 616 349
rect 600 315 719 333
rect 566 299 719 315
rect 478 215 494 249
rect 478 199 528 215
rect 571 249 651 265
rect 571 215 590 249
rect 624 215 651 249
rect 571 199 651 215
rect 685 165 719 299
rect 110 157 198 165
rect 110 123 148 157
rect 182 123 198 157
rect 110 89 198 123
rect 110 55 148 89
rect 182 55 198 89
rect 110 53 198 55
rect 232 157 322 165
rect 232 123 260 157
rect 294 123 322 157
rect 232 89 322 123
rect 232 55 260 89
rect 294 55 322 89
rect 232 17 322 55
rect 356 131 588 165
rect 356 129 390 131
rect 542 129 588 131
rect 356 51 390 95
rect 424 89 508 97
rect 424 55 446 89
rect 480 55 508 89
rect 424 17 508 55
rect 576 95 588 129
rect 542 51 588 95
rect 622 157 719 165
rect 622 123 638 157
rect 672 123 719 157
rect 622 89 719 123
rect 622 55 638 89
rect 672 55 719 89
rect 622 51 719 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 122 425 156 459 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 398 289 432 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 357 432 391 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 122 153 156 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 122 85 156 119 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 122 289 156 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 122 357 156 391 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o31a_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 1431166
string GDS_START 1423900
string path 0.000 0.000 3.680 0.000 
<< end >>
