magic
tech sky130A
magscale 1 2
timestamp 1652331711
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 945 945 979 979
rect 1611 945 1645 979
rect 131 871 165 905
rect 649 871 683 905
rect 945 871 979 905
rect 1315 871 1349 905
rect 2055 871 2089 905
rect 131 797 165 831
rect 649 797 683 831
rect 2055 797 2089 831
rect 131 723 165 757
rect 649 723 683 757
rect 945 723 979 757
rect 1611 723 1645 757
rect 2055 723 2089 757
rect 131 649 165 683
rect 649 649 683 683
rect 945 649 979 683
rect 2055 649 2089 683
rect 131 575 165 609
rect 649 575 683 609
rect 871 575 905 609
rect 2055 575 2089 609
rect 131 501 165 535
rect 1611 501 1645 535
rect 2055 501 2089 535
rect 131 427 165 461
rect 649 427 683 461
rect 871 427 905 461
rect 945 427 979 461
rect 1611 427 1645 461
rect 2055 427 2089 461
<< metal1 >>
rect -34 1446 2254 1514
rect -34 -34 2254 34
use xor2X1_pcell  xor2X1_pcell_0 pcells
timestamp 1652331234
transform 1 0 0 0 1 0
box -87 -34 2307 1550
<< labels >>
rlabel metal1 1611 723 1645 757 1 Y
port 1 n
rlabel metal1 1611 945 1645 979 1 Y
port 2 n
rlabel metal1 1611 501 1645 535 1 Y
port 3 n
rlabel metal1 1611 427 1645 461 1 Y
port 4 n
rlabel metal1 945 723 979 757 1 Y
port 5 n
rlabel metal1 945 649 979 683 1 Y
port 6 n
rlabel metal1 945 871 979 905 1 Y
port 7 n
rlabel metal1 945 945 979 979 1 Y
port 8 n
rlabel metal1 945 427 979 461 1 Y
port 9 n
rlabel metal1 131 797 165 831 1 A
port 10 n
rlabel metal1 131 723 165 757 1 A
port 11 n
rlabel metal1 131 649 165 683 1 A
port 12 n
rlabel metal1 131 575 165 609 1 A
port 13 n
rlabel metal1 131 501 165 535 1 A
port 14 n
rlabel metal1 131 427 165 461 1 A
port 15 n
rlabel metal1 131 871 165 905 1 A
port 16 n
rlabel metal1 649 871 683 905 1 A
port 17 n
rlabel metal1 649 797 683 831 1 A
port 18 n
rlabel metal1 649 723 683 757 1 A
port 19 n
rlabel metal1 649 649 683 683 1 A
port 20 n
rlabel metal1 649 575 683 609 1 A
port 21 n
rlabel metal1 649 427 683 461 1 A
port 22 n
rlabel metal1 2055 871 2089 905 1 B
port 23 n
rlabel metal1 2055 797 2089 831 1 B
port 24 n
rlabel metal1 2055 723 2089 757 1 B
port 25 n
rlabel metal1 2055 649 2089 683 1 B
port 26 n
rlabel metal1 2055 575 2089 609 1 B
port 27 n
rlabel metal1 2055 501 2089 535 1 B
port 28 n
rlabel metal1 2055 427 2089 461 1 B
port 29 n
rlabel metal1 1315 871 1349 905 1 B
port 30 n
rlabel metal1 871 575 905 609 1 B
port 31 n
rlabel metal1 871 427 905 461 1 B
port 32 n
rlabel metal1 -34 1446 2254 1514 1 VDD
port 33 n
rlabel metal1 -34 -34 2254 34 1 GND
port 34 n
rlabel nwell 57 1463 91 1497 1 VPB
port 35 n
rlabel pwell 57 -17 91 17 1 VNB
port 36 n
<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 2220 1480
string LEFsymmetry X Y R90
<< end >>
