// File: invx1_pcell.spi.pex
// Created: Tue Oct 15 15:57:06 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_INVX1_PCELL\%noxref_2 ( 5 17 30 32 33 34 )
c23 ( 34 0 ) capacitor c=0.0451925f //x=1.41 //y=5.02
c24 ( 33 0 ) capacitor c=0.0427416f //x=0.54 //y=5.02
c25 ( 32 0 ) capacitor c=0.234796f //x=1.48 //y=7.4
c26 ( 30 0 ) capacitor c=0.233263f //x=0.74 //y=7.4
c27 ( 17 0 ) capacitor c=0.028745f //x=1.47 //y=7.4
c28 ( 5 0 ) capacitor c=0.110692f //x=1.48 //y=7.4
r29 (  19 32 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.555 //y=7.23 //x2=1.555 //y2=7.4
r30 (  19 34 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=6.405
r31 (  18 30 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.76 //y=7.4 //x2=0.675 //y2=7.4
r32 (  17 32 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=1.555 //y2=7.4
r33 (  17 18 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=0.76 //y2=7.4
r34 (  11 30 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=0.675 //y=7.23 //x2=0.675 //y2=7.4
r35 (  11 33 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=6.405
r36 (  5 32 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=1.48 //y=7.4 //x2=1.48 //y2=7.4
r37 (  2 30 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=7.4 //x2=0.74 //y2=7.4
r38 (  2 5 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.48 //y2=7.4
ends PM_INVX1_PCELL\%noxref_2

subckt PM_INVX1_PCELL\%noxref_3 ( 2 7 8 9 10 11 12 13 17 18 19 21 27 28 30 )
c38 ( 30 0 ) capacitor c=0.0537799f //x=0.74 //y=2.085
c39 ( 28 0 ) capacitor c=0.0435629f //x=1.38 //y=1.255
c40 ( 27 0 ) capacitor c=0.0200386f //x=1.38 //y=0.91
c41 ( 21 0 ) capacitor c=0.0152946f //x=1.225 //y=1.41
c42 ( 19 0 ) capacitor c=0.0157804f //x=1.225 //y=0.755
c43 ( 18 0 ) capacitor c=0.0524167f //x=0.97 //y=4.79
c44 ( 17 0 ) capacitor c=0.0322983f //x=1.26 //y=4.79
c45 ( 13 0 ) capacitor c=0.0290017f //x=0.85 //y=1.92
c46 ( 12 0 ) capacitor c=0.0250027f //x=0.85 //y=1.565
c47 ( 11 0 ) capacitor c=0.0234316f //x=0.85 //y=1.255
c48 ( 10 0 ) capacitor c=0.0200596f //x=0.85 //y=0.91
c49 ( 9 0 ) capacitor c=0.154218f //x=1.335 //y=6.02
c50 ( 8 0 ) capacitor c=0.154243f //x=0.895 //y=6.02
c51 ( 2 0 ) capacitor c=0.115492f //x=0.74 //y=2.085
r52 (  30 31 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=0.74 //y=2.085 //x2=0.85 //y2=2.085
r53 (  28 37 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=1.255 //x2=1.34 //y2=1.41
r54 (  27 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.34 //y2=0.755
r55 (  27 28 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.38 //y2=1.255
r56 (  22 35 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=1.41 //x2=0.89 //y2=1.41
r57 (  21 37 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=1.41 //x2=1.34 //y2=1.41
r58 (  20 34 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=0.755 //x2=0.89 //y2=0.755
r59 (  19 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.34 //y2=0.755
r60 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.005 //y2=0.755
r61 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=1.335 //y2=4.865
r62 (  17 18 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=0.97 //y2=4.79
r63 (  14 18 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.97 //y2=4.79
r64 (  14 33 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.74 //y2=4.7
r65 (  13 31 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.92 //x2=0.85 //y2=2.085
r66 (  12 35 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.89 //y2=1.41
r67 (  12 13 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.85 //y2=1.92
r68 (  11 35 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.255 //x2=0.89 //y2=1.41
r69 (  10 34 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.89 //y2=0.755
r70 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.85 //y2=1.255
r71 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.335 //y=6.02 //x2=1.335 //y2=4.865
r72 (  8 14 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.895 //y=6.02 //x2=0.895 //y2=4.865
r73 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.225 //y2=1.41
r74 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.005 //y2=1.41
r75 (  5 33 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.7 //x2=0.74 //y2=4.7
r76 (  2 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=2.085
r77 (  2 5 ) resistor r=178.995 //w=0.187 //l=2.615 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=4.7
ends PM_INVX1_PCELL\%noxref_3

subckt PM_INVX1_PCELL\%noxref_4 ( 11 12 13 14 16 17 19 )
c33 ( 19 0 ) capacitor c=0.028734f //x=0.97 //y=5.02
c34 ( 17 0 ) capacitor c=0.0173218f //x=0.925 //y=0.91
c35 ( 16 0 ) capacitor c=0.10647f //x=1.48 //y=4.495
c36 ( 14 0 ) capacitor c=0.00575887f //x=1.2 //y=4.58
c37 ( 13 0 ) capacitor c=0.0146395f //x=1.395 //y=4.58
c38 ( 12 0 ) capacitor c=0.00636159f //x=1.195 //y=2.08
c39 ( 11 0 ) capacitor c=0.0141837f //x=1.395 //y=2.08
r40 (  15 16 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=1.48 //y=2.165 //x2=1.48 //y2=4.495
r41 (  13 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.48 //y2=4.495
r42 (  13 14 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.2 //y2=4.58
r43 (  11 15 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.48 //y2=2.165
r44 (  11 12 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=1.395 //y=2.08 //x2=1.195 //y2=2.08
r45 (  5 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.2 //y2=4.58
r46 (  5 19 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li //thickness=0.1 \
 //x=1.115 //y=4.665 //x2=1.115 //y2=5.725
r47 (  1 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.195 //y2=2.08
r48 (  1 17 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=1.11 //y=1.995 //x2=1.11 //y2=1.005
ends PM_INVX1_PCELL\%noxref_4

