magic
tech sky130A
magscale 1 2
timestamp 1669201001
<< nwell >>
rect -87 786 235 1550
<< pwell >>
rect -34 -34 182 544
<< psubdiff >>
rect -34 482 182 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 17 34 57
rect 114 461 182 482
rect 114 427 131 461
rect 165 427 182 461
rect 114 387 182 427
rect 114 353 131 387
rect 165 353 182 387
rect 114 313 182 353
rect 114 279 131 313
rect 165 279 182 313
rect 114 239 182 279
rect 114 205 131 239
rect 165 205 182 239
rect 114 165 182 205
rect 114 131 131 165
rect 165 131 182 165
rect 114 91 182 131
rect 114 57 131 91
rect 165 57 182 91
rect 114 17 182 57
rect -34 -17 57 17
rect 91 -17 182 17
rect -34 -34 182 -17
<< nsubdiff >>
rect -34 1497 182 1514
rect -34 1463 57 1497
rect 91 1463 182 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 884 34 905
rect 114 1423 182 1463
rect 114 1389 131 1423
rect 165 1389 182 1423
rect 114 1349 182 1389
rect 114 1315 131 1349
rect 165 1315 182 1349
rect 114 1275 182 1315
rect 114 1241 131 1275
rect 165 1241 182 1275
rect 114 1201 182 1241
rect 114 1167 131 1201
rect 165 1167 182 1201
rect 114 1127 182 1167
rect 114 1093 131 1127
rect 165 1093 182 1127
rect 114 1053 182 1093
rect 114 1019 131 1053
rect 165 1019 182 1053
rect 114 979 182 1019
rect 114 945 131 979
rect 165 945 182 979
rect 114 905 182 945
rect 114 884 131 905
rect 17 871 131 884
rect 165 871 182 905
rect -34 822 182 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 131 427 165 461
rect 131 353 165 387
rect 131 279 165 313
rect 131 205 165 239
rect 131 131 165 165
rect 131 57 165 91
rect 57 -17 91 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect -17 945 17 979
rect -17 871 17 905
rect 131 1389 165 1423
rect 131 1315 165 1349
rect 131 1241 165 1275
rect 131 1167 165 1201
rect 131 1093 165 1127
rect 131 1019 165 1053
rect 131 945 165 979
rect 131 871 165 905
<< locali >>
rect -34 1497 182 1514
rect -34 1463 57 1497
rect 91 1463 182 1497
rect -34 1446 182 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 114 1423 182 1446
rect 114 1389 131 1423
rect 165 1389 182 1423
rect 114 1349 182 1389
rect 114 1315 131 1349
rect 165 1315 182 1349
rect 114 1275 182 1315
rect 114 1241 131 1275
rect 165 1241 182 1275
rect 114 1201 182 1241
rect 114 1167 131 1201
rect 165 1167 182 1201
rect 114 1127 182 1167
rect 114 1093 131 1127
rect 165 1093 182 1127
rect 114 1053 182 1093
rect 114 1019 131 1053
rect 165 1019 182 1053
rect 114 979 182 1019
rect 114 945 131 979
rect 165 945 182 979
rect 114 905 182 945
rect 114 871 131 905
rect 165 871 182 905
rect 114 822 182 871
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 114 461 182 544
rect 114 427 131 461
rect 165 427 182 461
rect 114 387 182 427
rect 114 353 131 387
rect 165 353 182 387
rect 114 313 182 353
rect 114 279 131 313
rect 165 279 182 313
rect 114 239 182 279
rect 114 205 131 239
rect 165 205 182 239
rect 114 165 182 205
rect 114 131 131 165
rect 165 131 182 165
rect 114 91 182 131
rect 114 57 131 91
rect 165 57 182 91
rect 114 34 182 57
rect -34 17 182 34
rect -34 -17 57 17
rect 91 -17 182 17
rect -34 -34 182 -17
<< metal1 >>
rect -34 1446 182 1514
rect -34 -34 182 34
<< labels >>
rlabel metal1 -34 1446 182 1514 1 VPWR
port 1 n
rlabel metal1 -34 -34 182 34 1 VGND
port 2 n
rlabel nwell 57 1463 91 1497 1 VPB
port 3 n
rlabel pwell 57 -17 91 17 1 VNB
port 4 n
<< end >>
