* SPICE3 file created from AND2X1.ext - technology: sky130A

.subckt AND2X1 Y A B VDD VSS
X0 VDD A a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0.00278 pd=2.278 as=0 ps=0 w=2 l=0.15 M=2
X1 Y a_217_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0058 pd=4.58 as=0 ps=0 w=2 l=0.15 M=2
X2 Y a_217_1050 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0.0013199 ps=9.67 w=3 l=0.15
X3 VDD B a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X4 VSS A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X5 a_217_1050 B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 VDD a_217_1050 2.24f
.ends
