* SPICE3 file created from BUFX1.ext - technology: sky130A

.subckt BUFX1 Y A VDD VSS
X0 a_185_209 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.0022 ps=1.82 w=2 l=0.15 M=2
X1 a_185_209 A VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.0022816 ps=1.62 w=3 l=0.15
X2 VDD a_185_209 Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.0058 ps=4.58 w=2 l=0.15 M=2
X3 Y a_185_209 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
.ends
