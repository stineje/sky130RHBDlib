magic
tech sky130A
magscale 1 2
timestamp 1669564298
<< nwell >>
rect -87 786 3417 1550
<< pwell >>
rect -34 -34 3364 544
<< nmos >>
rect 168 288 198 349
tri 198 288 214 304 sw
rect 362 296 392 349
tri 392 296 408 312 sw
rect 168 258 274 288
tri 274 258 304 288 sw
rect 362 266 468 296
tri 468 266 498 296 sw
rect 168 157 198 258
tri 198 242 214 258 nw
tri 258 242 274 258 ne
tri 198 157 214 173 sw
tri 258 157 274 173 se
rect 274 157 304 258
rect 362 165 392 266
tri 392 250 408 266 nw
tri 452 250 468 266 ne
tri 392 165 408 181 sw
tri 452 165 468 181 se
rect 468 165 498 266
tri 168 127 198 157 ne
rect 198 127 274 157
tri 274 127 304 157 nw
tri 362 135 392 165 ne
rect 392 135 468 165
tri 468 135 498 165 nw
rect 821 297 851 350
tri 851 297 867 313 sw
rect 821 267 927 297
tri 927 267 957 297 sw
rect 821 166 851 267
tri 851 251 867 267 nw
tri 911 251 927 267 ne
tri 851 166 867 182 sw
tri 911 166 927 182 se
rect 927 166 957 267
tri 821 136 851 166 ne
rect 851 136 927 166
tri 927 136 957 166 nw
rect 1265 297 1295 350
tri 1295 297 1311 313 sw
rect 1265 267 1371 297
tri 1371 267 1401 297 sw
rect 1265 166 1295 267
tri 1295 251 1311 267 nw
tri 1355 251 1371 267 ne
tri 1295 166 1311 182 sw
tri 1355 166 1371 182 se
rect 1371 166 1401 267
tri 1265 136 1295 166 ne
rect 1295 136 1371 166
tri 1371 136 1401 166 nw
rect 1722 289 1752 350
tri 1752 289 1768 305 sw
rect 1916 297 1946 350
tri 1946 297 1962 313 sw
rect 1722 259 1828 289
tri 1828 259 1858 289 sw
rect 1916 267 2022 297
tri 2022 267 2052 297 sw
rect 1722 158 1752 259
tri 1752 243 1768 259 nw
tri 1812 243 1828 259 ne
tri 1752 158 1768 174 sw
tri 1812 158 1828 174 se
rect 1828 158 1858 259
rect 1916 166 1946 267
tri 1946 251 1962 267 nw
tri 2006 251 2022 267 ne
tri 1946 166 1962 182 sw
tri 2006 166 2022 182 se
rect 2022 166 2052 267
tri 1722 128 1752 158 ne
rect 1752 128 1828 158
tri 1828 128 1858 158 nw
tri 1916 136 1946 166 ne
rect 1946 136 2022 166
tri 2022 136 2052 166 nw
rect 2388 289 2418 350
tri 2418 289 2434 305 sw
rect 2582 297 2612 350
tri 2612 297 2628 313 sw
rect 2388 259 2494 289
tri 2494 259 2524 289 sw
rect 2582 267 2688 297
tri 2688 267 2718 297 sw
rect 2388 158 2418 259
tri 2418 243 2434 259 nw
tri 2478 243 2494 259 ne
tri 2418 158 2434 174 sw
tri 2478 158 2494 174 se
rect 2494 158 2524 259
rect 2582 166 2612 267
tri 2612 251 2628 267 nw
tri 2672 251 2688 267 ne
tri 2612 166 2628 182 sw
tri 2672 166 2688 182 se
rect 2688 166 2718 267
tri 2388 128 2418 158 ne
rect 2418 128 2494 158
tri 2494 128 2524 158 nw
tri 2582 136 2612 166 ne
rect 2612 136 2688 166
tri 2688 136 2718 166 nw
tri 3129 297 3145 313 se
rect 3145 297 3175 350
tri 3039 267 3069 297 se
rect 3069 267 3175 297
rect 3039 166 3069 267
tri 3069 251 3085 267 nw
tri 3129 251 3145 267 ne
tri 3069 166 3085 182 sw
tri 3129 166 3145 182 se
rect 3145 166 3175 267
tri 3039 136 3069 166 ne
rect 3069 136 3145 166
tri 3145 136 3175 166 nw
<< pmos >>
rect 187 1004 217 1404
rect 275 1004 305 1404
rect 363 1004 393 1404
rect 451 1004 481 1404
rect 830 1004 860 1404
rect 918 1004 948 1404
rect 1274 1004 1304 1404
rect 1362 1004 1392 1404
rect 1741 1004 1771 1404
rect 1829 1004 1859 1404
rect 1917 1004 1947 1404
rect 2005 1004 2035 1404
rect 2407 1004 2437 1404
rect 2495 1004 2525 1404
rect 2583 1004 2613 1404
rect 2671 1004 2701 1404
rect 3048 1004 3078 1404
rect 3136 1004 3166 1404
<< ndiff >>
rect 112 333 168 349
rect 112 299 122 333
rect 156 299 168 333
rect 112 261 168 299
rect 198 333 362 349
rect 198 304 219 333
tri 198 288 214 304 ne
rect 214 299 219 304
rect 253 299 316 333
rect 350 299 362 333
rect 214 288 362 299
rect 392 312 554 349
tri 392 296 408 312 ne
rect 408 296 554 312
rect 112 227 122 261
rect 156 227 168 261
tri 274 258 304 288 ne
rect 304 261 362 288
tri 468 266 498 296 ne
rect 112 193 168 227
rect 112 159 122 193
rect 156 159 168 193
rect 112 127 168 159
tri 198 242 214 258 se
rect 214 242 258 258
tri 258 242 274 258 sw
rect 198 208 274 242
rect 198 174 219 208
rect 253 174 274 208
rect 198 173 274 174
tri 198 157 214 173 ne
rect 214 157 258 173
tri 258 157 274 173 nw
rect 304 227 316 261
rect 350 227 362 261
rect 304 193 362 227
rect 304 159 316 193
rect 350 159 362 193
tri 392 250 408 266 se
rect 408 250 452 266
tri 452 250 468 266 sw
rect 392 217 468 250
rect 392 183 413 217
rect 447 183 468 217
rect 392 181 468 183
tri 392 165 408 181 ne
rect 408 165 452 181
tri 452 165 468 181 nw
rect 498 261 554 296
rect 498 227 510 261
rect 544 227 554 261
rect 498 193 554 227
tri 168 127 198 157 sw
tri 274 127 304 157 se
rect 304 135 362 159
tri 362 135 392 165 sw
tri 468 135 498 165 se
rect 498 159 510 193
rect 544 159 554 193
rect 498 135 554 159
rect 304 127 554 135
rect 112 123 554 127
rect 112 89 122 123
rect 156 89 316 123
rect 350 89 413 123
rect 447 89 510 123
rect 544 89 554 123
rect 112 73 554 89
rect 765 334 821 350
rect 765 300 775 334
rect 809 300 821 334
rect 765 262 821 300
rect 851 334 1011 350
rect 851 313 969 334
tri 851 297 867 313 ne
rect 867 300 969 313
rect 1003 300 1011 334
rect 867 297 1011 300
tri 927 267 957 297 ne
rect 765 228 775 262
rect 809 228 821 262
rect 765 194 821 228
rect 765 160 775 194
rect 809 160 821 194
tri 851 251 867 267 se
rect 867 251 911 267
tri 911 251 927 267 sw
rect 851 218 927 251
rect 851 184 871 218
rect 905 184 927 218
rect 851 182 927 184
tri 851 166 867 182 ne
rect 867 166 911 182
tri 911 166 927 182 nw
rect 957 262 1011 297
rect 957 228 969 262
rect 1003 228 1011 262
rect 957 194 1011 228
rect 765 136 821 160
tri 821 136 851 166 sw
tri 927 136 957 166 se
rect 957 160 969 194
rect 1003 160 1011 194
rect 957 136 1011 160
rect 765 124 1011 136
rect 765 90 775 124
rect 809 90 871 124
rect 905 90 969 124
rect 1003 90 1011 124
rect 765 74 1011 90
rect 1209 334 1265 350
rect 1209 300 1219 334
rect 1253 300 1265 334
rect 1209 262 1265 300
rect 1295 334 1455 350
rect 1295 313 1413 334
tri 1295 297 1311 313 ne
rect 1311 300 1413 313
rect 1447 300 1455 334
rect 1311 297 1455 300
tri 1371 267 1401 297 ne
rect 1209 228 1219 262
rect 1253 228 1265 262
rect 1209 194 1265 228
rect 1209 160 1219 194
rect 1253 160 1265 194
tri 1295 251 1311 267 se
rect 1311 251 1355 267
tri 1355 251 1371 267 sw
rect 1295 218 1371 251
rect 1295 184 1315 218
rect 1349 184 1371 218
rect 1295 182 1371 184
tri 1295 166 1311 182 ne
rect 1311 166 1355 182
tri 1355 166 1371 182 nw
rect 1401 262 1455 297
rect 1401 228 1413 262
rect 1447 228 1455 262
rect 1401 194 1455 228
rect 1209 136 1265 160
tri 1265 136 1295 166 sw
tri 1371 136 1401 166 se
rect 1401 160 1413 194
rect 1447 160 1455 194
rect 1401 136 1455 160
rect 1209 124 1455 136
rect 1209 90 1219 124
rect 1253 90 1315 124
rect 1349 90 1413 124
rect 1447 90 1455 124
rect 1209 74 1455 90
rect 1666 334 1722 350
rect 1666 300 1676 334
rect 1710 300 1722 334
rect 1666 262 1722 300
rect 1752 334 1916 350
rect 1752 305 1773 334
tri 1752 289 1768 305 ne
rect 1768 300 1773 305
rect 1807 300 1870 334
rect 1904 300 1916 334
rect 1768 289 1916 300
rect 1946 313 2108 350
tri 1946 297 1962 313 ne
rect 1962 297 2108 313
rect 1666 228 1676 262
rect 1710 228 1722 262
tri 1828 259 1858 289 ne
rect 1858 262 1916 289
tri 2022 267 2052 297 ne
rect 1666 194 1722 228
rect 1666 160 1676 194
rect 1710 160 1722 194
rect 1666 128 1722 160
tri 1752 243 1768 259 se
rect 1768 243 1812 259
tri 1812 243 1828 259 sw
rect 1752 209 1828 243
rect 1752 175 1773 209
rect 1807 175 1828 209
rect 1752 174 1828 175
tri 1752 158 1768 174 ne
rect 1768 158 1812 174
tri 1812 158 1828 174 nw
rect 1858 228 1870 262
rect 1904 228 1916 262
rect 1858 194 1916 228
rect 1858 160 1870 194
rect 1904 160 1916 194
tri 1946 251 1962 267 se
rect 1962 251 2006 267
tri 2006 251 2022 267 sw
rect 1946 218 2022 251
rect 1946 184 1967 218
rect 2001 184 2022 218
rect 1946 182 2022 184
tri 1946 166 1962 182 ne
rect 1962 166 2006 182
tri 2006 166 2022 182 nw
rect 2052 262 2108 297
rect 2052 228 2064 262
rect 2098 228 2108 262
rect 2052 194 2108 228
tri 1722 128 1752 158 sw
tri 1828 128 1858 158 se
rect 1858 136 1916 160
tri 1916 136 1946 166 sw
tri 2022 136 2052 166 se
rect 2052 160 2064 194
rect 2098 160 2108 194
rect 2052 136 2108 160
rect 1858 128 2108 136
rect 1666 124 2108 128
rect 1666 90 1676 124
rect 1710 90 1870 124
rect 1904 90 1967 124
rect 2001 90 2064 124
rect 2098 90 2108 124
rect 1666 74 2108 90
rect 2332 334 2388 350
rect 2332 300 2342 334
rect 2376 300 2388 334
rect 2332 262 2388 300
rect 2418 334 2582 350
rect 2418 305 2439 334
tri 2418 289 2434 305 ne
rect 2434 300 2439 305
rect 2473 300 2536 334
rect 2570 300 2582 334
rect 2434 289 2582 300
rect 2612 313 2774 350
tri 2612 297 2628 313 ne
rect 2628 297 2774 313
rect 2332 228 2342 262
rect 2376 228 2388 262
tri 2494 259 2524 289 ne
rect 2524 262 2582 289
tri 2688 267 2718 297 ne
rect 2332 194 2388 228
rect 2332 160 2342 194
rect 2376 160 2388 194
rect 2332 128 2388 160
tri 2418 243 2434 259 se
rect 2434 243 2478 259
tri 2478 243 2494 259 sw
rect 2418 209 2494 243
rect 2418 175 2439 209
rect 2473 175 2494 209
rect 2418 174 2494 175
tri 2418 158 2434 174 ne
rect 2434 158 2478 174
tri 2478 158 2494 174 nw
rect 2524 228 2536 262
rect 2570 228 2582 262
rect 2524 194 2582 228
rect 2524 160 2536 194
rect 2570 160 2582 194
tri 2612 251 2628 267 se
rect 2628 251 2672 267
tri 2672 251 2688 267 sw
rect 2612 218 2688 251
rect 2612 184 2633 218
rect 2667 184 2688 218
rect 2612 182 2688 184
tri 2612 166 2628 182 ne
rect 2628 166 2672 182
tri 2672 166 2688 182 nw
rect 2718 262 2774 297
rect 2718 228 2730 262
rect 2764 228 2774 262
rect 2718 194 2774 228
tri 2388 128 2418 158 sw
tri 2494 128 2524 158 se
rect 2524 136 2582 160
tri 2582 136 2612 166 sw
tri 2688 136 2718 166 se
rect 2718 160 2730 194
rect 2764 160 2774 194
rect 2718 136 2774 160
rect 2524 128 2774 136
rect 2332 124 2774 128
rect 2332 90 2342 124
rect 2376 90 2536 124
rect 2570 90 2633 124
rect 2667 90 2730 124
rect 2764 90 2774 124
rect 2332 74 2774 90
rect 2985 334 3145 350
rect 2985 300 2993 334
rect 3027 313 3145 334
rect 3027 300 3129 313
rect 2985 297 3129 300
tri 3129 297 3145 313 nw
rect 3175 334 3231 350
rect 3175 300 3187 334
rect 3221 300 3231 334
rect 2985 262 3039 297
tri 3039 267 3069 297 nw
rect 2985 228 2993 262
rect 3027 228 3039 262
rect 2985 194 3039 228
rect 2985 160 2993 194
rect 3027 160 3039 194
tri 3069 251 3085 267 se
rect 3085 251 3129 267
tri 3129 251 3145 267 sw
rect 3069 218 3145 251
rect 3069 184 3091 218
rect 3125 184 3145 218
rect 3069 182 3145 184
tri 3069 166 3085 182 ne
rect 3085 166 3129 182
tri 3129 166 3145 182 nw
rect 3175 262 3231 300
rect 3175 228 3187 262
rect 3221 228 3231 262
rect 3175 194 3231 228
rect 2985 136 3039 160
tri 3039 136 3069 166 sw
tri 3145 136 3175 166 se
rect 3175 160 3187 194
rect 3221 160 3231 194
rect 3175 136 3231 160
rect 2985 124 3231 136
rect 2985 90 2993 124
rect 3027 90 3091 124
rect 3125 90 3187 124
rect 3221 90 3231 124
rect 2985 74 3231 90
<< pdiff >>
rect 131 1366 187 1404
rect 131 1332 141 1366
rect 175 1332 187 1366
rect 131 1298 187 1332
rect 131 1264 141 1298
rect 175 1264 187 1298
rect 131 1230 187 1264
rect 131 1196 141 1230
rect 175 1196 187 1230
rect 131 1162 187 1196
rect 131 1128 141 1162
rect 175 1128 187 1162
rect 131 1093 187 1128
rect 131 1059 141 1093
rect 175 1059 187 1093
rect 131 1004 187 1059
rect 217 1366 275 1404
rect 217 1332 229 1366
rect 263 1332 275 1366
rect 217 1298 275 1332
rect 217 1264 229 1298
rect 263 1264 275 1298
rect 217 1230 275 1264
rect 217 1196 229 1230
rect 263 1196 275 1230
rect 217 1162 275 1196
rect 217 1128 229 1162
rect 263 1128 275 1162
rect 217 1093 275 1128
rect 217 1059 229 1093
rect 263 1059 275 1093
rect 217 1004 275 1059
rect 305 1366 363 1404
rect 305 1332 317 1366
rect 351 1332 363 1366
rect 305 1298 363 1332
rect 305 1264 317 1298
rect 351 1264 363 1298
rect 305 1230 363 1264
rect 305 1196 317 1230
rect 351 1196 363 1230
rect 305 1162 363 1196
rect 305 1128 317 1162
rect 351 1128 363 1162
rect 305 1004 363 1128
rect 393 1366 451 1404
rect 393 1332 405 1366
rect 439 1332 451 1366
rect 393 1298 451 1332
rect 393 1264 405 1298
rect 439 1264 451 1298
rect 393 1230 451 1264
rect 393 1196 405 1230
rect 439 1196 451 1230
rect 393 1162 451 1196
rect 393 1128 405 1162
rect 439 1128 451 1162
rect 393 1093 451 1128
rect 393 1059 405 1093
rect 439 1059 451 1093
rect 393 1004 451 1059
rect 481 1366 535 1404
rect 481 1332 493 1366
rect 527 1332 535 1366
rect 481 1298 535 1332
rect 481 1264 493 1298
rect 527 1264 535 1298
rect 481 1230 535 1264
rect 481 1196 493 1230
rect 527 1196 535 1230
rect 481 1162 535 1196
rect 481 1128 493 1162
rect 527 1128 535 1162
rect 481 1004 535 1128
rect 774 1366 830 1404
rect 774 1332 784 1366
rect 818 1332 830 1366
rect 774 1298 830 1332
rect 774 1264 784 1298
rect 818 1264 830 1298
rect 774 1230 830 1264
rect 774 1196 784 1230
rect 818 1196 830 1230
rect 774 1162 830 1196
rect 774 1128 784 1162
rect 818 1128 830 1162
rect 774 1093 830 1128
rect 774 1059 784 1093
rect 818 1059 830 1093
rect 774 1004 830 1059
rect 860 1366 918 1404
rect 860 1332 872 1366
rect 906 1332 918 1366
rect 860 1298 918 1332
rect 860 1264 872 1298
rect 906 1264 918 1298
rect 860 1230 918 1264
rect 860 1196 872 1230
rect 906 1196 918 1230
rect 860 1162 918 1196
rect 860 1128 872 1162
rect 906 1128 918 1162
rect 860 1093 918 1128
rect 860 1059 872 1093
rect 906 1059 918 1093
rect 860 1004 918 1059
rect 948 1366 1002 1404
rect 948 1332 960 1366
rect 994 1332 1002 1366
rect 948 1298 1002 1332
rect 948 1264 960 1298
rect 994 1264 1002 1298
rect 948 1230 1002 1264
rect 948 1196 960 1230
rect 994 1196 1002 1230
rect 948 1162 1002 1196
rect 948 1128 960 1162
rect 994 1128 1002 1162
rect 948 1093 1002 1128
rect 948 1059 960 1093
rect 994 1059 1002 1093
rect 948 1004 1002 1059
rect 1218 1366 1274 1404
rect 1218 1332 1228 1366
rect 1262 1332 1274 1366
rect 1218 1298 1274 1332
rect 1218 1264 1228 1298
rect 1262 1264 1274 1298
rect 1218 1230 1274 1264
rect 1218 1196 1228 1230
rect 1262 1196 1274 1230
rect 1218 1162 1274 1196
rect 1218 1128 1228 1162
rect 1262 1128 1274 1162
rect 1218 1093 1274 1128
rect 1218 1059 1228 1093
rect 1262 1059 1274 1093
rect 1218 1004 1274 1059
rect 1304 1366 1362 1404
rect 1304 1332 1316 1366
rect 1350 1332 1362 1366
rect 1304 1298 1362 1332
rect 1304 1264 1316 1298
rect 1350 1264 1362 1298
rect 1304 1230 1362 1264
rect 1304 1196 1316 1230
rect 1350 1196 1362 1230
rect 1304 1162 1362 1196
rect 1304 1128 1316 1162
rect 1350 1128 1362 1162
rect 1304 1093 1362 1128
rect 1304 1059 1316 1093
rect 1350 1059 1362 1093
rect 1304 1004 1362 1059
rect 1392 1366 1446 1404
rect 1392 1332 1404 1366
rect 1438 1332 1446 1366
rect 1392 1298 1446 1332
rect 1392 1264 1404 1298
rect 1438 1264 1446 1298
rect 1392 1230 1446 1264
rect 1392 1196 1404 1230
rect 1438 1196 1446 1230
rect 1392 1162 1446 1196
rect 1392 1128 1404 1162
rect 1438 1128 1446 1162
rect 1392 1093 1446 1128
rect 1392 1059 1404 1093
rect 1438 1059 1446 1093
rect 1392 1004 1446 1059
rect 1685 1364 1741 1404
rect 1685 1330 1695 1364
rect 1729 1330 1741 1364
rect 1685 1296 1741 1330
rect 1685 1262 1695 1296
rect 1729 1262 1741 1296
rect 1685 1228 1741 1262
rect 1685 1194 1695 1228
rect 1729 1194 1741 1228
rect 1685 1160 1741 1194
rect 1685 1126 1695 1160
rect 1729 1126 1741 1160
rect 1685 1092 1741 1126
rect 1685 1058 1695 1092
rect 1729 1058 1741 1092
rect 1685 1004 1741 1058
rect 1771 1296 1829 1404
rect 1771 1262 1783 1296
rect 1817 1262 1829 1296
rect 1771 1228 1829 1262
rect 1771 1194 1783 1228
rect 1817 1194 1829 1228
rect 1771 1160 1829 1194
rect 1771 1126 1783 1160
rect 1817 1126 1829 1160
rect 1771 1004 1829 1126
rect 1859 1364 1917 1404
rect 1859 1330 1871 1364
rect 1905 1330 1917 1364
rect 1859 1296 1917 1330
rect 1859 1262 1871 1296
rect 1905 1262 1917 1296
rect 1859 1228 1917 1262
rect 1859 1194 1871 1228
rect 1905 1194 1917 1228
rect 1859 1160 1917 1194
rect 1859 1126 1871 1160
rect 1905 1126 1917 1160
rect 1859 1092 1917 1126
rect 1859 1058 1871 1092
rect 1905 1058 1917 1092
rect 1859 1004 1917 1058
rect 1947 1296 2005 1404
rect 1947 1262 1959 1296
rect 1993 1262 2005 1296
rect 1947 1228 2005 1262
rect 1947 1194 1959 1228
rect 1993 1194 2005 1228
rect 1947 1160 2005 1194
rect 1947 1126 1959 1160
rect 1993 1126 2005 1160
rect 1947 1092 2005 1126
rect 1947 1058 1959 1092
rect 1993 1058 2005 1092
rect 1947 1004 2005 1058
rect 2035 1364 2089 1404
rect 2035 1330 2047 1364
rect 2081 1330 2089 1364
rect 2035 1296 2089 1330
rect 2035 1262 2047 1296
rect 2081 1262 2089 1296
rect 2035 1228 2089 1262
rect 2035 1194 2047 1228
rect 2081 1194 2089 1228
rect 2035 1160 2089 1194
rect 2035 1126 2047 1160
rect 2081 1126 2089 1160
rect 2035 1004 2089 1126
rect 2351 1364 2407 1404
rect 2351 1330 2361 1364
rect 2395 1330 2407 1364
rect 2351 1296 2407 1330
rect 2351 1262 2361 1296
rect 2395 1262 2407 1296
rect 2351 1228 2407 1262
rect 2351 1194 2361 1228
rect 2395 1194 2407 1228
rect 2351 1160 2407 1194
rect 2351 1126 2361 1160
rect 2395 1126 2407 1160
rect 2351 1092 2407 1126
rect 2351 1058 2361 1092
rect 2395 1058 2407 1092
rect 2351 1004 2407 1058
rect 2437 1296 2495 1404
rect 2437 1262 2449 1296
rect 2483 1262 2495 1296
rect 2437 1228 2495 1262
rect 2437 1194 2449 1228
rect 2483 1194 2495 1228
rect 2437 1160 2495 1194
rect 2437 1126 2449 1160
rect 2483 1126 2495 1160
rect 2437 1004 2495 1126
rect 2525 1364 2583 1404
rect 2525 1330 2537 1364
rect 2571 1330 2583 1364
rect 2525 1296 2583 1330
rect 2525 1262 2537 1296
rect 2571 1262 2583 1296
rect 2525 1228 2583 1262
rect 2525 1194 2537 1228
rect 2571 1194 2583 1228
rect 2525 1160 2583 1194
rect 2525 1126 2537 1160
rect 2571 1126 2583 1160
rect 2525 1092 2583 1126
rect 2525 1058 2537 1092
rect 2571 1058 2583 1092
rect 2525 1004 2583 1058
rect 2613 1296 2671 1404
rect 2613 1262 2625 1296
rect 2659 1262 2671 1296
rect 2613 1228 2671 1262
rect 2613 1194 2625 1228
rect 2659 1194 2671 1228
rect 2613 1160 2671 1194
rect 2613 1126 2625 1160
rect 2659 1126 2671 1160
rect 2613 1092 2671 1126
rect 2613 1058 2625 1092
rect 2659 1058 2671 1092
rect 2613 1004 2671 1058
rect 2701 1364 2755 1404
rect 2701 1330 2713 1364
rect 2747 1330 2755 1364
rect 2701 1296 2755 1330
rect 2701 1262 2713 1296
rect 2747 1262 2755 1296
rect 2701 1228 2755 1262
rect 2701 1194 2713 1228
rect 2747 1194 2755 1228
rect 2701 1160 2755 1194
rect 2701 1126 2713 1160
rect 2747 1126 2755 1160
rect 2701 1004 2755 1126
rect 2994 1366 3048 1404
rect 2994 1332 3002 1366
rect 3036 1332 3048 1366
rect 2994 1298 3048 1332
rect 2994 1264 3002 1298
rect 3036 1264 3048 1298
rect 2994 1230 3048 1264
rect 2994 1196 3002 1230
rect 3036 1196 3048 1230
rect 2994 1162 3048 1196
rect 2994 1128 3002 1162
rect 3036 1128 3048 1162
rect 2994 1093 3048 1128
rect 2994 1059 3002 1093
rect 3036 1059 3048 1093
rect 2994 1004 3048 1059
rect 3078 1366 3136 1404
rect 3078 1332 3090 1366
rect 3124 1332 3136 1366
rect 3078 1298 3136 1332
rect 3078 1264 3090 1298
rect 3124 1264 3136 1298
rect 3078 1230 3136 1264
rect 3078 1196 3090 1230
rect 3124 1196 3136 1230
rect 3078 1162 3136 1196
rect 3078 1128 3090 1162
rect 3124 1128 3136 1162
rect 3078 1093 3136 1128
rect 3078 1059 3090 1093
rect 3124 1059 3136 1093
rect 3078 1004 3136 1059
rect 3166 1366 3222 1404
rect 3166 1332 3178 1366
rect 3212 1332 3222 1366
rect 3166 1298 3222 1332
rect 3166 1264 3178 1298
rect 3212 1264 3222 1298
rect 3166 1230 3222 1264
rect 3166 1196 3178 1230
rect 3212 1196 3222 1230
rect 3166 1162 3222 1196
rect 3166 1128 3178 1162
rect 3212 1128 3222 1162
rect 3166 1093 3222 1128
rect 3166 1059 3178 1093
rect 3212 1059 3222 1093
rect 3166 1004 3222 1059
<< ndiffc >>
rect 122 299 156 333
rect 219 299 253 333
rect 316 299 350 333
rect 122 227 156 261
rect 122 159 156 193
rect 219 174 253 208
rect 316 227 350 261
rect 316 159 350 193
rect 413 183 447 217
rect 510 227 544 261
rect 510 159 544 193
rect 122 89 156 123
rect 316 89 350 123
rect 413 89 447 123
rect 510 89 544 123
rect 775 300 809 334
rect 969 300 1003 334
rect 775 228 809 262
rect 775 160 809 194
rect 871 184 905 218
rect 969 228 1003 262
rect 969 160 1003 194
rect 775 90 809 124
rect 871 90 905 124
rect 969 90 1003 124
rect 1219 300 1253 334
rect 1413 300 1447 334
rect 1219 228 1253 262
rect 1219 160 1253 194
rect 1315 184 1349 218
rect 1413 228 1447 262
rect 1413 160 1447 194
rect 1219 90 1253 124
rect 1315 90 1349 124
rect 1413 90 1447 124
rect 1676 300 1710 334
rect 1773 300 1807 334
rect 1870 300 1904 334
rect 1676 228 1710 262
rect 1676 160 1710 194
rect 1773 175 1807 209
rect 1870 228 1904 262
rect 1870 160 1904 194
rect 1967 184 2001 218
rect 2064 228 2098 262
rect 2064 160 2098 194
rect 1676 90 1710 124
rect 1870 90 1904 124
rect 1967 90 2001 124
rect 2064 90 2098 124
rect 2342 300 2376 334
rect 2439 300 2473 334
rect 2536 300 2570 334
rect 2342 228 2376 262
rect 2342 160 2376 194
rect 2439 175 2473 209
rect 2536 228 2570 262
rect 2536 160 2570 194
rect 2633 184 2667 218
rect 2730 228 2764 262
rect 2730 160 2764 194
rect 2342 90 2376 124
rect 2536 90 2570 124
rect 2633 90 2667 124
rect 2730 90 2764 124
rect 2993 300 3027 334
rect 3187 300 3221 334
rect 2993 228 3027 262
rect 2993 160 3027 194
rect 3091 184 3125 218
rect 3187 228 3221 262
rect 3187 160 3221 194
rect 2993 90 3027 124
rect 3091 90 3125 124
rect 3187 90 3221 124
<< pdiffc >>
rect 141 1332 175 1366
rect 141 1264 175 1298
rect 141 1196 175 1230
rect 141 1128 175 1162
rect 141 1059 175 1093
rect 229 1332 263 1366
rect 229 1264 263 1298
rect 229 1196 263 1230
rect 229 1128 263 1162
rect 229 1059 263 1093
rect 317 1332 351 1366
rect 317 1264 351 1298
rect 317 1196 351 1230
rect 317 1128 351 1162
rect 405 1332 439 1366
rect 405 1264 439 1298
rect 405 1196 439 1230
rect 405 1128 439 1162
rect 405 1059 439 1093
rect 493 1332 527 1366
rect 493 1264 527 1298
rect 493 1196 527 1230
rect 493 1128 527 1162
rect 784 1332 818 1366
rect 784 1264 818 1298
rect 784 1196 818 1230
rect 784 1128 818 1162
rect 784 1059 818 1093
rect 872 1332 906 1366
rect 872 1264 906 1298
rect 872 1196 906 1230
rect 872 1128 906 1162
rect 872 1059 906 1093
rect 960 1332 994 1366
rect 960 1264 994 1298
rect 960 1196 994 1230
rect 960 1128 994 1162
rect 960 1059 994 1093
rect 1228 1332 1262 1366
rect 1228 1264 1262 1298
rect 1228 1196 1262 1230
rect 1228 1128 1262 1162
rect 1228 1059 1262 1093
rect 1316 1332 1350 1366
rect 1316 1264 1350 1298
rect 1316 1196 1350 1230
rect 1316 1128 1350 1162
rect 1316 1059 1350 1093
rect 1404 1332 1438 1366
rect 1404 1264 1438 1298
rect 1404 1196 1438 1230
rect 1404 1128 1438 1162
rect 1404 1059 1438 1093
rect 1695 1330 1729 1364
rect 1695 1262 1729 1296
rect 1695 1194 1729 1228
rect 1695 1126 1729 1160
rect 1695 1058 1729 1092
rect 1783 1262 1817 1296
rect 1783 1194 1817 1228
rect 1783 1126 1817 1160
rect 1871 1330 1905 1364
rect 1871 1262 1905 1296
rect 1871 1194 1905 1228
rect 1871 1126 1905 1160
rect 1871 1058 1905 1092
rect 1959 1262 1993 1296
rect 1959 1194 1993 1228
rect 1959 1126 1993 1160
rect 1959 1058 1993 1092
rect 2047 1330 2081 1364
rect 2047 1262 2081 1296
rect 2047 1194 2081 1228
rect 2047 1126 2081 1160
rect 2361 1330 2395 1364
rect 2361 1262 2395 1296
rect 2361 1194 2395 1228
rect 2361 1126 2395 1160
rect 2361 1058 2395 1092
rect 2449 1262 2483 1296
rect 2449 1194 2483 1228
rect 2449 1126 2483 1160
rect 2537 1330 2571 1364
rect 2537 1262 2571 1296
rect 2537 1194 2571 1228
rect 2537 1126 2571 1160
rect 2537 1058 2571 1092
rect 2625 1262 2659 1296
rect 2625 1194 2659 1228
rect 2625 1126 2659 1160
rect 2625 1058 2659 1092
rect 2713 1330 2747 1364
rect 2713 1262 2747 1296
rect 2713 1194 2747 1228
rect 2713 1126 2747 1160
rect 3002 1332 3036 1366
rect 3002 1264 3036 1298
rect 3002 1196 3036 1230
rect 3002 1128 3036 1162
rect 3002 1059 3036 1093
rect 3090 1332 3124 1366
rect 3090 1264 3124 1298
rect 3090 1196 3124 1230
rect 3090 1128 3124 1162
rect 3090 1059 3124 1093
rect 3178 1332 3212 1366
rect 3178 1264 3212 1298
rect 3178 1196 3212 1230
rect 3178 1128 3212 1162
rect 3178 1059 3212 1093
<< psubdiff >>
rect -34 482 3364 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 632 461 700 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 632 427 649 461
rect 683 427 700 461
rect 1076 461 1144 482
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 1520 461 1588 482
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 632 313 700 353
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 1520 427 1537 461
rect 1571 427 1588 461
rect 2186 461 2254 482
rect 632 279 649 313
rect 683 279 700 313
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect -34 17 34 57
rect 632 57 649 91
rect 683 57 700 91
rect 1076 313 1144 353
rect 1520 387 1588 427
rect 1520 353 1537 387
rect 1571 353 1588 387
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 632 17 700 57
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1520 313 1588 353
rect 2186 427 2203 461
rect 2237 427 2254 461
rect 2852 461 2920 482
rect 2186 387 2254 427
rect 2186 353 2203 387
rect 2237 353 2254 387
rect 1520 279 1537 313
rect 1571 279 1588 313
rect 1520 239 1588 279
rect 1520 205 1537 239
rect 1571 205 1588 239
rect 1520 165 1588 205
rect 1520 131 1537 165
rect 1571 131 1588 165
rect 1520 91 1588 131
rect 1076 17 1144 57
rect 1520 57 1537 91
rect 1571 57 1588 91
rect 2186 313 2254 353
rect 2852 427 2869 461
rect 2903 427 2920 461
rect 3296 461 3364 482
rect 2852 387 2920 427
rect 2852 353 2869 387
rect 2903 353 2920 387
rect 2186 279 2203 313
rect 2237 279 2254 313
rect 2186 239 2254 279
rect 2186 205 2203 239
rect 2237 205 2254 239
rect 2186 165 2254 205
rect 2186 131 2203 165
rect 2237 131 2254 165
rect 2186 91 2254 131
rect 1520 17 1588 57
rect 2186 57 2203 91
rect 2237 57 2254 91
rect 2852 313 2920 353
rect 3296 427 3313 461
rect 3347 427 3364 461
rect 3296 387 3364 427
rect 3296 353 3313 387
rect 3347 353 3364 387
rect 2852 279 2869 313
rect 2903 279 2920 313
rect 2852 239 2920 279
rect 2852 205 2869 239
rect 2903 205 2920 239
rect 2852 165 2920 205
rect 2852 131 2869 165
rect 2903 131 2920 165
rect 2852 91 2920 131
rect 2186 17 2254 57
rect 2852 57 2869 91
rect 2903 57 2920 91
rect 3296 313 3364 353
rect 3296 279 3313 313
rect 3347 279 3364 313
rect 3296 239 3364 279
rect 3296 205 3313 239
rect 3347 205 3364 239
rect 3296 165 3364 205
rect 3296 131 3313 165
rect 3347 131 3364 165
rect 3296 91 3364 131
rect 2852 17 2920 57
rect 3296 57 3313 91
rect 3347 57 3364 91
rect 3296 17 3364 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3364 17
rect -34 -34 3364 -17
<< nsubdiff >>
rect -34 1497 3364 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3364 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 632 1423 700 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 1076 1423 1144 1463
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 632 979 700 1019
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1520 1423 1588 1463
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 632 945 649 979
rect 683 945 700 979
rect -34 871 -17 905
rect 17 884 34 905
rect 632 905 700 945
rect 1076 979 1144 1019
rect 1520 1389 1537 1423
rect 1571 1389 1588 1423
rect 2186 1423 2254 1463
rect 1520 1349 1588 1389
rect 1520 1315 1537 1349
rect 1571 1315 1588 1349
rect 1520 1275 1588 1315
rect 1520 1241 1537 1275
rect 1571 1241 1588 1275
rect 1520 1201 1588 1241
rect 1520 1167 1537 1201
rect 1571 1167 1588 1201
rect 1520 1127 1588 1167
rect 1520 1093 1537 1127
rect 1571 1093 1588 1127
rect 1520 1053 1588 1093
rect 1520 1019 1537 1053
rect 1571 1019 1588 1053
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 632 884 649 905
rect 17 871 649 884
rect 683 884 700 905
rect 1076 905 1144 945
rect 1520 979 1588 1019
rect 2186 1389 2203 1423
rect 2237 1389 2254 1423
rect 2852 1423 2920 1463
rect 2186 1349 2254 1389
rect 2186 1315 2203 1349
rect 2237 1315 2254 1349
rect 2186 1275 2254 1315
rect 2186 1241 2203 1275
rect 2237 1241 2254 1275
rect 2186 1201 2254 1241
rect 2186 1167 2203 1201
rect 2237 1167 2254 1201
rect 2186 1127 2254 1167
rect 2186 1093 2203 1127
rect 2237 1093 2254 1127
rect 2186 1053 2254 1093
rect 2186 1019 2203 1053
rect 2237 1019 2254 1053
rect 1520 945 1537 979
rect 1571 945 1588 979
rect 1076 884 1093 905
rect 683 871 1093 884
rect 1127 884 1144 905
rect 1520 905 1588 945
rect 2186 979 2254 1019
rect 2852 1389 2869 1423
rect 2903 1389 2920 1423
rect 3296 1423 3364 1463
rect 2852 1349 2920 1389
rect 2852 1315 2869 1349
rect 2903 1315 2920 1349
rect 2852 1275 2920 1315
rect 2852 1241 2869 1275
rect 2903 1241 2920 1275
rect 2852 1201 2920 1241
rect 2852 1167 2869 1201
rect 2903 1167 2920 1201
rect 2852 1127 2920 1167
rect 2852 1093 2869 1127
rect 2903 1093 2920 1127
rect 2852 1053 2920 1093
rect 2852 1019 2869 1053
rect 2903 1019 2920 1053
rect 2186 945 2203 979
rect 2237 945 2254 979
rect 1520 884 1537 905
rect 1127 871 1537 884
rect 1571 884 1588 905
rect 2186 905 2254 945
rect 2852 979 2920 1019
rect 3296 1389 3313 1423
rect 3347 1389 3364 1423
rect 3296 1349 3364 1389
rect 3296 1315 3313 1349
rect 3347 1315 3364 1349
rect 3296 1275 3364 1315
rect 3296 1241 3313 1275
rect 3347 1241 3364 1275
rect 3296 1201 3364 1241
rect 3296 1167 3313 1201
rect 3347 1167 3364 1201
rect 3296 1127 3364 1167
rect 3296 1093 3313 1127
rect 3347 1093 3364 1127
rect 3296 1053 3364 1093
rect 3296 1019 3313 1053
rect 3347 1019 3364 1053
rect 2852 945 2869 979
rect 2903 945 2920 979
rect 2186 884 2203 905
rect 1571 871 2203 884
rect 2237 884 2254 905
rect 2852 905 2920 945
rect 3296 979 3364 1019
rect 3296 945 3313 979
rect 3347 945 3364 979
rect 2852 884 2869 905
rect 2237 871 2869 884
rect 2903 884 2920 905
rect 3296 905 3364 945
rect 3296 884 3313 905
rect 2903 871 3313 884
rect 3347 871 3364 905
rect -34 822 3364 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 649 427 683 461
rect 649 353 683 387
rect 1093 427 1127 461
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1093 353 1127 387
rect 1537 427 1571 461
rect 649 279 683 313
rect 649 205 683 239
rect 649 131 683 165
rect 649 57 683 91
rect 1537 353 1571 387
rect 1093 279 1127 313
rect 1093 205 1127 239
rect 1093 131 1127 165
rect 1093 57 1127 91
rect 2203 427 2237 461
rect 2203 353 2237 387
rect 1537 279 1571 313
rect 1537 205 1571 239
rect 1537 131 1571 165
rect 1537 57 1571 91
rect 2869 427 2903 461
rect 2869 353 2903 387
rect 2203 279 2237 313
rect 2203 205 2237 239
rect 2203 131 2237 165
rect 2203 57 2237 91
rect 3313 427 3347 461
rect 3313 353 3347 387
rect 2869 279 2903 313
rect 2869 205 2903 239
rect 2869 131 2903 165
rect 2869 57 2903 91
rect 3313 279 3347 313
rect 3313 205 3347 239
rect 3313 131 3347 165
rect 3313 57 3347 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 649 1389 683 1423
rect 649 1315 683 1349
rect 649 1241 683 1275
rect 649 1167 683 1201
rect 649 1093 683 1127
rect 649 1019 683 1053
rect -17 945 17 979
rect 1093 1389 1127 1423
rect 1093 1315 1127 1349
rect 1093 1241 1127 1275
rect 1093 1167 1127 1201
rect 1093 1093 1127 1127
rect 1093 1019 1127 1053
rect 649 945 683 979
rect -17 871 17 905
rect 1537 1389 1571 1423
rect 1537 1315 1571 1349
rect 1537 1241 1571 1275
rect 1537 1167 1571 1201
rect 1537 1093 1571 1127
rect 1537 1019 1571 1053
rect 1093 945 1127 979
rect 649 871 683 905
rect 2203 1389 2237 1423
rect 2203 1315 2237 1349
rect 2203 1241 2237 1275
rect 2203 1167 2237 1201
rect 2203 1093 2237 1127
rect 2203 1019 2237 1053
rect 1537 945 1571 979
rect 1093 871 1127 905
rect 2869 1389 2903 1423
rect 2869 1315 2903 1349
rect 2869 1241 2903 1275
rect 2869 1167 2903 1201
rect 2869 1093 2903 1127
rect 2869 1019 2903 1053
rect 2203 945 2237 979
rect 1537 871 1571 905
rect 3313 1389 3347 1423
rect 3313 1315 3347 1349
rect 3313 1241 3347 1275
rect 3313 1167 3347 1201
rect 3313 1093 3347 1127
rect 3313 1019 3347 1053
rect 2869 945 2903 979
rect 2203 871 2237 905
rect 3313 945 3347 979
rect 2869 871 2903 905
rect 3313 871 3347 905
<< poly >>
rect 187 1404 217 1430
rect 275 1404 305 1430
rect 363 1404 393 1430
rect 451 1404 481 1430
rect 830 1404 860 1430
rect 918 1404 948 1430
rect 187 973 217 1004
rect 275 973 305 1004
rect 363 973 393 1004
rect 451 973 481 1004
rect 187 957 305 973
rect 187 943 205 957
rect 195 923 205 943
rect 239 943 305 957
rect 349 957 481 973
rect 239 923 249 943
rect 195 907 249 923
rect 349 923 359 957
rect 393 943 481 957
rect 1274 1404 1304 1430
rect 1362 1404 1392 1430
rect 830 973 860 1004
rect 918 973 948 1004
rect 393 923 403 943
rect 349 907 403 923
rect 787 957 948 973
rect 787 923 797 957
rect 831 943 948 957
rect 1741 1404 1771 1430
rect 1829 1404 1859 1430
rect 1917 1404 1947 1430
rect 2005 1404 2035 1430
rect 1274 973 1304 1004
rect 1362 973 1392 1004
rect 831 923 841 943
rect 787 907 841 923
rect 1231 957 1392 973
rect 1231 923 1241 957
rect 1275 943 1392 957
rect 2407 1404 2437 1430
rect 2495 1404 2525 1430
rect 2583 1404 2613 1430
rect 2671 1404 2701 1430
rect 1275 923 1285 943
rect 1231 907 1285 923
rect 1741 973 1771 1004
rect 1829 973 1859 1004
rect 1741 957 1859 973
rect 1741 943 1759 957
rect 1749 923 1759 943
rect 1793 943 1859 957
rect 1917 973 1947 1004
rect 2005 973 2035 1004
rect 1917 957 2035 973
rect 1917 943 1981 957
rect 1793 923 1803 943
rect 1749 907 1803 923
rect 1971 923 1981 943
rect 2015 943 2035 957
rect 3048 1404 3078 1430
rect 3136 1404 3166 1430
rect 2015 923 2025 943
rect 1971 907 2025 923
rect 2407 973 2437 1004
rect 2495 973 2525 1004
rect 2407 957 2525 973
rect 2407 943 2425 957
rect 2415 923 2425 943
rect 2459 943 2525 957
rect 2583 973 2613 1004
rect 2671 973 2701 1004
rect 2583 957 2701 973
rect 2583 943 2647 957
rect 2459 923 2469 943
rect 2415 907 2469 923
rect 2637 923 2647 943
rect 2681 943 2701 957
rect 2681 923 2691 943
rect 2637 907 2691 923
rect 3048 973 3078 1004
rect 3136 973 3166 1004
rect 3048 957 3209 973
rect 3048 943 3165 957
rect 3155 923 3165 943
rect 3199 923 3209 957
rect 3155 907 3209 923
rect 195 433 249 449
rect 195 413 205 433
rect 168 399 205 413
rect 239 399 249 433
rect 168 383 249 399
rect 343 433 397 449
rect 343 399 353 433
rect 387 399 397 433
rect 343 383 397 399
rect 168 349 198 383
rect 362 349 392 383
rect 787 434 841 450
rect 787 400 797 434
rect 831 413 841 434
rect 831 400 851 413
rect 787 384 851 400
rect 821 350 851 384
rect 1231 434 1285 450
rect 1231 400 1241 434
rect 1275 413 1285 434
rect 1275 400 1295 413
rect 1231 384 1295 400
rect 1265 350 1295 384
rect 1749 434 1803 450
rect 1749 414 1759 434
rect 1722 400 1759 414
rect 1793 400 1803 434
rect 1971 434 2025 450
rect 1971 414 1981 434
rect 1722 384 1803 400
rect 1916 400 1981 414
rect 2015 400 2025 434
rect 1916 384 2025 400
rect 2415 434 2469 450
rect 2415 414 2425 434
rect 1722 350 1752 384
rect 1916 350 1946 384
rect 2388 400 2425 414
rect 2459 400 2469 434
rect 2637 434 2691 450
rect 2637 414 2647 434
rect 2388 384 2469 400
rect 2582 400 2647 414
rect 2681 400 2691 434
rect 2582 384 2691 400
rect 3155 434 3209 450
rect 3155 413 3165 434
rect 2388 350 2418 384
rect 2582 350 2612 384
rect 3145 400 3165 413
rect 3199 400 3209 434
rect 3145 384 3209 400
rect 3145 350 3175 384
<< polycont >>
rect 205 923 239 957
rect 359 923 393 957
rect 797 923 831 957
rect 1241 923 1275 957
rect 1759 923 1793 957
rect 1981 923 2015 957
rect 2425 923 2459 957
rect 2647 923 2681 957
rect 3165 923 3199 957
rect 205 399 239 433
rect 353 399 387 433
rect 797 400 831 434
rect 1241 400 1275 434
rect 1759 400 1793 434
rect 1981 400 2015 434
rect 2425 400 2459 434
rect 2647 400 2681 434
rect 3165 400 3199 434
<< locali >>
rect -34 1497 3364 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3364 1497
rect -34 1446 3364 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 141 1366 175 1446
rect 141 1298 175 1332
rect 141 1230 175 1264
rect 141 1162 175 1196
rect 141 1093 175 1128
rect 141 1027 175 1059
rect 229 1366 263 1404
rect 229 1298 263 1332
rect 229 1230 263 1264
rect 229 1162 263 1196
rect 229 1093 263 1128
rect 317 1366 351 1446
rect 317 1298 351 1332
rect 317 1230 351 1264
rect 317 1162 351 1196
rect 317 1111 351 1128
rect 405 1366 439 1404
rect 405 1298 439 1332
rect 405 1230 439 1264
rect 405 1162 439 1196
rect 229 1057 263 1059
rect 405 1093 439 1128
rect 493 1366 527 1446
rect 493 1298 527 1332
rect 493 1230 527 1264
rect 493 1162 527 1196
rect 493 1111 527 1128
rect 632 1423 700 1446
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 405 1057 439 1059
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 229 1023 535 1057
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 359 957 393 973
rect 205 831 239 923
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 797
rect 205 383 239 399
rect 353 923 359 942
rect 353 907 393 923
rect 353 757 387 907
rect 353 433 387 723
rect 353 383 387 399
rect 501 683 535 1023
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect 784 1366 818 1446
rect 784 1298 818 1332
rect 784 1230 818 1264
rect 784 1162 818 1196
rect 784 1093 818 1128
rect 784 1037 818 1059
rect 872 1366 906 1404
rect 872 1298 906 1332
rect 872 1230 906 1264
rect 872 1162 906 1196
rect 872 1093 906 1128
rect 632 979 700 1019
rect 632 945 649 979
rect 683 945 700 979
rect 632 905 700 945
rect 632 871 649 905
rect 683 871 700 905
rect 632 822 700 871
rect 797 957 831 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 122 333 156 349
rect 316 333 350 349
rect 501 348 535 649
rect 797 683 831 923
rect 872 933 906 1059
rect 960 1366 994 1446
rect 960 1298 994 1332
rect 960 1230 994 1264
rect 960 1162 994 1196
rect 960 1093 994 1128
rect 960 1037 994 1059
rect 1076 1423 1144 1446
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 1228 1366 1262 1446
rect 1228 1298 1262 1332
rect 1228 1230 1262 1264
rect 1228 1162 1262 1196
rect 1228 1093 1262 1128
rect 1228 1037 1262 1059
rect 1316 1366 1350 1404
rect 1316 1298 1350 1332
rect 1316 1230 1350 1264
rect 1316 1162 1350 1196
rect 1316 1093 1350 1128
rect 1076 979 1144 1019
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 872 899 979 933
rect 156 299 219 333
rect 253 299 316 333
rect 122 261 156 299
rect 122 193 156 227
rect 316 261 350 299
rect 122 123 156 159
rect 122 73 156 89
rect 219 208 253 224
rect -34 34 34 57
rect 219 34 253 174
rect 316 193 350 227
rect 413 314 535 348
rect 632 461 700 544
rect 632 427 649 461
rect 683 427 700 461
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect 797 434 831 649
rect 945 433 979 899
rect 1076 905 1144 945
rect 1076 871 1093 905
rect 1127 871 1144 905
rect 1076 822 1144 871
rect 1241 957 1275 973
rect 1241 831 1275 923
rect 1316 933 1350 1059
rect 1404 1366 1438 1446
rect 1404 1298 1438 1332
rect 1404 1230 1438 1264
rect 1404 1162 1438 1196
rect 1404 1093 1438 1128
rect 1404 1037 1438 1059
rect 1520 1423 1588 1446
rect 1520 1389 1537 1423
rect 1571 1389 1588 1423
rect 1520 1349 1588 1389
rect 1520 1315 1537 1349
rect 1571 1315 1588 1349
rect 1520 1275 1588 1315
rect 1520 1241 1537 1275
rect 1571 1241 1588 1275
rect 1520 1201 1588 1241
rect 1520 1167 1537 1201
rect 1571 1167 1588 1201
rect 1520 1127 1588 1167
rect 1520 1093 1537 1127
rect 1571 1093 1588 1127
rect 1520 1053 1588 1093
rect 1520 1019 1537 1053
rect 1571 1019 1588 1053
rect 1695 1364 1729 1380
rect 1695 1296 1729 1330
rect 1695 1228 1729 1262
rect 1695 1160 1729 1194
rect 1695 1092 1729 1126
rect 1783 1296 1817 1446
rect 2186 1423 2254 1446
rect 1783 1228 1817 1262
rect 1783 1160 1817 1194
rect 1783 1110 1817 1126
rect 1871 1364 2081 1398
rect 1871 1296 1905 1330
rect 1871 1228 1905 1262
rect 1871 1160 1905 1194
rect 1871 1092 1905 1126
rect 1695 1024 1905 1058
rect 1959 1296 1993 1312
rect 1959 1228 1993 1262
rect 1959 1160 1993 1194
rect 1959 1092 1993 1126
rect 2047 1296 2081 1330
rect 2047 1228 2081 1262
rect 2047 1160 2081 1194
rect 2047 1110 2081 1126
rect 2186 1389 2203 1423
rect 2237 1389 2254 1423
rect 2186 1349 2254 1389
rect 2186 1315 2203 1349
rect 2237 1315 2254 1349
rect 2186 1275 2254 1315
rect 2186 1241 2203 1275
rect 2237 1241 2254 1275
rect 2186 1201 2254 1241
rect 2186 1167 2203 1201
rect 2237 1167 2254 1201
rect 2186 1127 2254 1167
rect 2186 1093 2203 1127
rect 2237 1093 2254 1127
rect 1959 1024 2089 1058
rect 1520 979 1588 1019
rect 1520 945 1537 979
rect 1571 945 1588 979
rect 1316 899 1423 933
rect 797 384 831 400
rect 871 399 979 433
rect 1076 461 1144 544
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 413 217 447 314
rect 632 313 700 353
rect 632 279 649 313
rect 683 279 700 313
rect 413 167 447 183
rect 510 261 544 277
rect 510 193 544 227
rect 316 123 350 159
rect 510 123 544 159
rect 350 89 413 123
rect 447 89 510 123
rect 316 73 350 89
rect 510 73 544 89
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect 632 57 649 91
rect 683 57 700 91
rect 632 34 700 57
rect 775 334 809 350
rect 775 262 809 300
rect 775 194 809 228
rect 871 218 905 399
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 1241 434 1275 797
rect 1389 535 1423 899
rect 1520 905 1588 945
rect 1520 871 1537 905
rect 1571 871 1588 905
rect 1520 822 1588 871
rect 1759 957 1793 973
rect 1759 831 1793 923
rect 1981 957 2015 973
rect 1389 433 1423 501
rect 1241 384 1275 400
rect 1315 399 1423 433
rect 1520 461 1588 544
rect 1520 427 1537 461
rect 1571 427 1588 461
rect 871 168 905 184
rect 969 334 1003 350
rect 969 262 1003 300
rect 969 194 1003 228
rect 775 124 809 160
rect 969 124 1003 160
rect 809 90 871 124
rect 905 90 969 124
rect 775 34 809 90
rect 872 34 906 90
rect 969 34 1003 90
rect 1076 313 1144 353
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1076 34 1144 57
rect 1219 334 1253 350
rect 1219 262 1253 300
rect 1219 194 1253 228
rect 1315 218 1349 399
rect 1520 387 1588 427
rect 1520 353 1537 387
rect 1571 353 1588 387
rect 1759 434 1793 797
rect 1907 905 1941 921
rect 1907 757 1941 871
rect 1981 831 2015 923
rect 1981 781 2015 797
rect 1907 707 1941 723
rect 2055 757 2089 1024
rect 2186 1053 2254 1093
rect 2186 1019 2203 1053
rect 2237 1019 2254 1053
rect 2361 1364 2395 1380
rect 2361 1296 2395 1330
rect 2361 1228 2395 1262
rect 2361 1160 2395 1194
rect 2361 1092 2395 1126
rect 2449 1296 2483 1446
rect 2852 1423 2920 1446
rect 2449 1228 2483 1262
rect 2449 1160 2483 1194
rect 2449 1110 2483 1126
rect 2537 1364 2747 1398
rect 2537 1296 2571 1330
rect 2537 1228 2571 1262
rect 2537 1160 2571 1194
rect 2537 1092 2571 1126
rect 2361 1024 2571 1058
rect 2625 1296 2659 1312
rect 2625 1228 2659 1262
rect 2625 1160 2659 1194
rect 2625 1092 2659 1126
rect 2713 1296 2747 1330
rect 2713 1228 2747 1262
rect 2713 1160 2747 1194
rect 2713 1110 2747 1126
rect 2852 1389 2869 1423
rect 2903 1389 2920 1423
rect 2852 1349 2920 1389
rect 2852 1315 2869 1349
rect 2903 1315 2920 1349
rect 2852 1275 2920 1315
rect 2852 1241 2869 1275
rect 2903 1241 2920 1275
rect 2852 1201 2920 1241
rect 2852 1167 2869 1201
rect 2903 1167 2920 1201
rect 2852 1127 2920 1167
rect 2852 1093 2869 1127
rect 2903 1093 2920 1127
rect 2625 1024 2755 1058
rect 2186 979 2254 1019
rect 2186 945 2203 979
rect 2237 945 2254 979
rect 2186 905 2254 945
rect 2186 871 2203 905
rect 2237 871 2254 905
rect 2186 822 2254 871
rect 2425 957 2459 973
rect 2425 905 2459 923
rect 2425 855 2459 871
rect 2647 957 2681 973
rect 1759 384 1793 400
rect 1981 609 2015 625
rect 1981 434 2015 575
rect 1981 384 2015 400
rect 1315 168 1349 184
rect 1413 334 1447 350
rect 1413 262 1447 300
rect 1413 194 1447 228
rect 1219 124 1253 160
rect 1413 124 1447 160
rect 1253 90 1315 124
rect 1349 90 1413 124
rect 1219 34 1253 90
rect 1316 34 1350 90
rect 1413 34 1447 90
rect 1520 313 1588 353
rect 1520 279 1537 313
rect 1571 279 1588 313
rect 1520 239 1588 279
rect 1520 205 1537 239
rect 1571 205 1588 239
rect 1520 165 1588 205
rect 1520 131 1537 165
rect 1571 131 1588 165
rect 1520 91 1588 131
rect 1520 57 1537 91
rect 1571 57 1588 91
rect 1676 334 1710 350
rect 1870 334 1904 350
rect 2055 348 2089 723
rect 2425 683 2459 699
rect 1710 300 1773 334
rect 1807 300 1870 334
rect 1676 262 1710 300
rect 1676 194 1710 228
rect 1870 262 1904 300
rect 1676 124 1710 160
rect 1676 74 1710 90
rect 1773 209 1807 225
rect 1520 34 1588 57
rect 1773 34 1807 175
rect 1870 194 1904 228
rect 1967 314 2089 348
rect 2186 461 2254 544
rect 2186 427 2203 461
rect 2237 427 2254 461
rect 2186 387 2254 427
rect 2186 353 2203 387
rect 2237 353 2254 387
rect 2425 434 2459 649
rect 2425 384 2459 400
rect 2647 535 2681 923
rect 2647 434 2681 501
rect 2647 384 2681 400
rect 2721 757 2755 1024
rect 2852 1053 2920 1093
rect 2852 1019 2869 1053
rect 2903 1019 2920 1053
rect 3002 1366 3036 1446
rect 3002 1298 3036 1332
rect 3002 1230 3036 1264
rect 3002 1162 3036 1196
rect 3002 1093 3036 1128
rect 3002 1037 3036 1059
rect 3090 1366 3124 1404
rect 3090 1298 3124 1332
rect 3090 1230 3124 1264
rect 3090 1162 3124 1196
rect 3090 1093 3124 1128
rect 2852 979 2920 1019
rect 2852 945 2869 979
rect 2903 945 2920 979
rect 2852 905 2920 945
rect 3090 933 3124 1059
rect 3178 1366 3212 1446
rect 3178 1298 3212 1332
rect 3178 1230 3212 1264
rect 3178 1162 3212 1196
rect 3178 1093 3212 1128
rect 3178 1037 3212 1059
rect 3296 1423 3364 1446
rect 3296 1389 3313 1423
rect 3347 1389 3364 1423
rect 3296 1349 3364 1389
rect 3296 1315 3313 1349
rect 3347 1315 3364 1349
rect 3296 1275 3364 1315
rect 3296 1241 3313 1275
rect 3347 1241 3364 1275
rect 3296 1201 3364 1241
rect 3296 1167 3313 1201
rect 3347 1167 3364 1201
rect 3296 1127 3364 1167
rect 3296 1093 3313 1127
rect 3347 1093 3364 1127
rect 3296 1053 3364 1093
rect 3296 1019 3313 1053
rect 3347 1019 3364 1053
rect 3296 979 3364 1019
rect 2852 871 2869 905
rect 2903 871 2920 905
rect 2852 822 2920 871
rect 3017 899 3124 933
rect 3165 957 3199 973
rect 3165 905 3199 923
rect 3017 831 3051 899
rect 1967 218 2001 314
rect 2186 313 2254 353
rect 2186 279 2203 313
rect 2237 279 2254 313
rect 1967 168 2001 184
rect 2064 262 2098 278
rect 2064 194 2098 228
rect 1870 124 1904 160
rect 2064 124 2098 160
rect 1904 90 1967 124
rect 2001 90 2064 124
rect 1870 74 1904 90
rect 2064 74 2098 90
rect 2186 239 2254 279
rect 2186 205 2203 239
rect 2237 205 2254 239
rect 2186 165 2254 205
rect 2186 131 2203 165
rect 2237 131 2254 165
rect 2186 91 2254 131
rect 2186 57 2203 91
rect 2237 57 2254 91
rect 2342 334 2376 350
rect 2536 334 2570 350
rect 2721 348 2755 723
rect 3017 683 3051 797
rect 2376 300 2439 334
rect 2473 300 2536 334
rect 2342 262 2376 300
rect 2342 194 2376 228
rect 2536 262 2570 300
rect 2342 124 2376 160
rect 2342 74 2376 90
rect 2439 209 2473 225
rect 2186 34 2254 57
rect 2439 34 2473 175
rect 2536 194 2570 228
rect 2633 314 2755 348
rect 2852 461 2920 544
rect 2852 427 2869 461
rect 2903 427 2920 461
rect 2852 387 2920 427
rect 3017 433 3051 649
rect 3165 609 3199 871
rect 3296 945 3313 979
rect 3347 945 3364 979
rect 3296 905 3364 945
rect 3296 871 3313 905
rect 3347 871 3364 905
rect 3296 822 3364 871
rect 3165 434 3199 575
rect 3017 399 3125 433
rect 2852 353 2869 387
rect 2903 353 2920 387
rect 2633 218 2667 314
rect 2852 313 2920 353
rect 2852 279 2869 313
rect 2903 279 2920 313
rect 2633 168 2667 184
rect 2730 262 2764 278
rect 2730 194 2764 228
rect 2536 124 2570 160
rect 2730 124 2764 160
rect 2570 90 2633 124
rect 2667 90 2730 124
rect 2536 74 2570 90
rect 2730 74 2764 90
rect 2852 239 2920 279
rect 2852 205 2869 239
rect 2903 205 2920 239
rect 2852 165 2920 205
rect 2852 131 2869 165
rect 2903 131 2920 165
rect 2852 91 2920 131
rect 2852 57 2869 91
rect 2903 57 2920 91
rect 2852 34 2920 57
rect 2993 334 3027 350
rect 2993 262 3027 300
rect 2993 194 3027 228
rect 3091 218 3125 399
rect 3165 384 3199 400
rect 3296 461 3364 544
rect 3296 427 3313 461
rect 3347 427 3364 461
rect 3296 387 3364 427
rect 3296 353 3313 387
rect 3347 353 3364 387
rect 3091 168 3125 184
rect 3187 334 3221 350
rect 3187 262 3221 300
rect 3187 194 3221 228
rect 2993 124 3027 160
rect 3187 124 3221 160
rect 3027 90 3091 124
rect 3125 90 3187 124
rect 2993 34 3027 90
rect 3090 34 3124 90
rect 3187 34 3221 90
rect 3296 313 3364 353
rect 3296 279 3313 313
rect 3347 279 3364 313
rect 3296 239 3364 279
rect 3296 205 3313 239
rect 3347 205 3364 239
rect 3296 165 3364 205
rect 3296 131 3313 165
rect 3347 131 3364 165
rect 3296 91 3364 131
rect 3296 57 3313 91
rect 3347 57 3364 91
rect 3296 34 3364 57
rect -34 17 3364 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3364 17
rect -34 -34 3364 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 205 797 239 831
rect 353 723 387 757
rect 501 649 535 683
rect 797 649 831 683
rect 1241 797 1275 831
rect 1759 797 1793 831
rect 1389 501 1423 535
rect 1907 871 1941 905
rect 1981 797 2015 831
rect 1907 723 1941 757
rect 2425 871 2459 905
rect 2055 723 2089 757
rect 1981 575 2015 609
rect 2425 649 2459 683
rect 2647 501 2681 535
rect 2721 723 2755 757
rect 3017 797 3051 831
rect 3017 649 3051 683
rect 3165 871 3199 905
rect 3165 575 3199 609
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
<< metal1 >>
rect -34 1497 3364 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3364 1497
rect -34 1446 3364 1463
rect 1901 905 1947 911
rect 2419 905 2465 911
rect 3159 905 3205 911
rect 1895 871 1907 905
rect 1941 871 2425 905
rect 2459 871 3165 905
rect 3199 871 3211 905
rect 1901 865 1947 871
rect 2419 865 2465 871
rect 3159 865 3205 871
rect 199 831 245 837
rect 1235 831 1281 837
rect 1753 831 1799 837
rect 1975 831 2021 837
rect 3011 831 3057 837
rect 193 797 205 831
rect 239 797 1241 831
rect 1275 797 1759 831
rect 1793 797 1805 831
rect 1969 797 1981 831
rect 2015 797 3017 831
rect 3051 797 3063 831
rect 199 791 245 797
rect 1235 791 1281 797
rect 1753 791 1799 797
rect 1975 791 2021 797
rect 3011 791 3057 797
rect 347 757 393 763
rect 1901 757 1947 763
rect 2049 757 2095 763
rect 2715 757 2761 763
rect 341 723 353 757
rect 387 723 1907 757
rect 1941 723 1953 757
rect 2043 723 2055 757
rect 2089 723 2721 757
rect 2755 723 2767 757
rect 347 717 393 723
rect 1901 717 1947 723
rect 2049 717 2095 723
rect 2715 717 2761 723
rect 495 683 541 689
rect 791 683 837 689
rect 2419 683 2465 689
rect 3011 683 3057 689
rect 489 649 501 683
rect 535 649 797 683
rect 831 649 843 683
rect 2413 649 2425 683
rect 2459 649 3017 683
rect 3051 649 3063 683
rect 495 643 541 649
rect 791 643 837 649
rect 2419 643 2465 649
rect 3011 643 3057 649
rect 1975 609 2021 615
rect 3159 609 3205 615
rect 1969 575 1981 609
rect 2015 575 3165 609
rect 3199 575 3211 609
rect 1975 569 2021 575
rect 3159 569 3205 575
rect 1383 535 1429 541
rect 2641 535 2687 541
rect 1377 501 1389 535
rect 1423 501 2647 535
rect 2681 501 2693 535
rect 1383 495 1429 501
rect 2641 495 2687 501
rect -34 17 3364 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3364 17
rect -34 -34 3364 -17
<< labels >>
rlabel metal1 2721 723 2755 757 1 SUM
port 1 n
rlabel metal1 2055 723 2089 757 1 SUM
port 2 n
rlabel metal1 2721 427 2755 461 1 SUM
port 3 n
rlabel metal1 2721 501 2755 535 1 SUM
port 4 n
rlabel metal1 2721 945 2755 979 1 SUM
port 5 n
rlabel metal1 2055 649 2089 683 1 SUM
port 6 n
rlabel metal1 2055 427 2089 461 1 SUM
port 7 n
rlabel metal1 2055 945 2089 979 1 SUM
port 8 n
rlabel metal1 945 501 979 535 1 COUT
port 9 n
rlabel metal1 945 427 979 461 1 COUT
port 10 n
rlabel metal1 945 649 979 683 1 COUT
port 11 n
rlabel metal1 945 871 979 905 1 COUT
port 12 n
rlabel metal1 945 575 979 609 1 COUT
port 13 n
rlabel metal1 205 797 239 831 1 A
port 14 n
rlabel metal1 205 871 239 905 1 A
port 15 n
rlabel metal1 205 723 239 757 1 A
port 16 n
rlabel metal1 205 649 239 683 1 A
port 17 n
rlabel metal1 205 575 239 609 1 A
port 18 n
rlabel metal1 205 501 239 535 1 A
port 19 n
rlabel metal1 1241 871 1275 905 1 A
port 20 n
rlabel metal1 1241 797 1275 831 1 A
port 21 n
rlabel metal1 1241 649 1275 683 1 A
port 22 n
rlabel metal1 1241 575 1275 609 1 A
port 23 n
rlabel metal1 1241 501 1275 535 1 A
port 24 n
rlabel metal1 1759 871 1793 905 1 A
port 25 n
rlabel metal1 1759 797 1793 831 1 A
port 26 n
rlabel metal1 1759 649 1793 683 1 A
port 27 n
rlabel metal1 1759 575 1793 609 1 A
port 28 n
rlabel metal1 353 723 387 757 1 B
port 29 n
rlabel metal1 353 649 387 683 1 B
port 30 n
rlabel metal1 353 575 387 609 1 B
port 31 n
rlabel metal1 353 501 387 535 1 B
port 32 n
rlabel metal1 353 871 387 905 1 B
port 33 n
rlabel metal1 1907 723 1941 757 1 B
port 34 n
rlabel metal1 1907 797 1941 831 1 B
port 35 n
rlabel metal1 1907 871 1941 905 1 B
port 36 n
rlabel metal1 3165 723 3199 757 1 B
port 37 n
rlabel metal1 1981 575 2015 609 1 B
port 38 n
rlabel metal1 3165 575 3199 609 1 B
port 39 n
rlabel metal1 3165 649 3199 683 1 B
port 40 n
rlabel metal1 3165 501 3199 535 1 B
port 41 n
rlabel metal1 3165 797 3199 831 1 B
port 42 n
rlabel metal1 3165 871 3199 905 1 B
port 43 n
rlabel metal1 2425 871 2459 905 1 B
port 44 n
rlabel metal1 -34 1446 3364 1514 1 VPWR
port 45 n
rlabel metal1 -34 -34 3364 34 1 VGND
port 46 n
rlabel nwell 57 1463 91 1497 1 VPB
port 47 n
rlabel pwell 57 -17 91 17 1 VNB
port 48 n
<< end >>
