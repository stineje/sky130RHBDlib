* SPICE3 file created from DFFRNX1.ext - technology: sky130A

.subckt DFFRNX1 Q QN D CLK RN VDD GND
X0 VDD CLK a_277_1004 VDD pshort w=2 l=0.15 M=2
X1 VDD a_277_1004 QN VDD pshort w=2 l=0.15 M=2
X2 a_599_943 RN VDD VDD pshort w=2 l=0.15 M=2
X3 QN Q VDD VDD pshort w=2 l=0.15 M=2
X4 GND a_147_159 a_91_75 GND nshort w=3 l=0.15
X5 a_147_159 CLK VDD VDD pshort w=2 l=0.15 M=2
X6 Q QN VDD VDD pshort w=2 l=0.15 M=2
X7 QN Q a_3924_182 GND nshort w=3 l=0.15
X8 VDD a_599_943 a_277_1004 VDD pshort w=2 l=0.15 M=2
X9 VDD a_147_159 a_2141_1004 VDD pshort w=2 l=0.15 M=2
X10 VDD a_2141_1004 a_147_159 VDD pshort w=2 l=0.15 M=2
X11 a_147_159 RN VDD VDD pshort w=2 l=0.15 M=2
X12 Q a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X13 a_372_182 CLK a_91_75 GND nshort w=3 l=0.15
X14 GND a_277_1004 a_3643_75 GND nshort w=3 l=0.15
X15 a_277_1004 a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X16 GND QN a_4626_73 GND nshort w=3 l=0.15
X17 VDD a_277_1004 a_599_943 VDD pshort w=2 l=0.15 M=2
X18 a_599_943 RN a_1334_182 GND nshort w=3 l=0.15
X19 GND a_599_943 a_2036_73 GND nshort w=3 l=0.15
X20 GND a_2141_1004 a_2681_75 GND nshort w=3 l=0.15
X21 a_2141_1004 a_599_943 VDD VDD pshort w=2 l=0.15 M=2
X22 a_3924_182 RN a_3643_75 GND nshort w=3 l=0.15
X23 VDD D a_599_943 VDD pshort w=2 l=0.15 M=2
X24 VDD RN QN VDD pshort w=2 l=0.15 M=2
X25 GND a_277_1004 a_1053_75 GND nshort w=3 l=0.15
X26 a_2962_182 CLK a_2681_75 GND nshort w=3 l=0.15
X27 a_1334_182 D a_1053_75 GND nshort w=3 l=0.15
X28 Q a_147_159 a_4626_73 GND nshort w=3 l=0.15
X29 a_2141_1004 a_147_159 a_2036_73 GND nshort w=3 l=0.15
X30 a_277_1004 a_599_943 a_372_182 GND nshort w=3 l=0.15
X31 a_147_159 RN a_2962_182 GND nshort w=3 l=0.15
C0 a_277_1004 a_147_159 3.63fF
C1 a_277_1004 VDD 2.39fF
C2 a_599_943 VDD 2.34fF
C3 a_147_159 VDD 3.82fF
C4 a_147_159 CLK 3.25fF
C5 a_277_1004 a_599_943 2.06fF
C6 VDD GND 12.57fF
.ends
