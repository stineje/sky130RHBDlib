VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
# Standard Cell LEF generated in Magic




MACRO AND2X1
  CLASS CORE ;
  FOREIGN AND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.550 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 5.985 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 5.720 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 3.920 5.185 4.090 7.230 ;
        RECT 4.800 5.185 4.970 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 5.720 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 5.720 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 3.875 0.620 4.045 1.750 ;
        RECT 4.845 0.620 5.015 1.750 ;
        RECT 3.875 0.450 5.015 0.620 ;
        RECT 3.875 0.170 4.045 0.450 ;
        RECT 4.360 0.170 4.530 0.450 ;
        RECT 4.845 0.170 5.015 0.450 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT -0.170 -0.170 5.720 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 5.720 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 3.985 1.920 4.155 4.865 ;
        RECT 4.360 4.665 4.530 7.020 ;
        RECT 4.360 4.495 4.895 4.665 ;
        RECT 4.725 2.165 4.895 4.495 ;
        RECT 4.355 1.995 4.895 2.165 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 4.355 0.840 4.525 1.995 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
      LAYER mcon ;
        RECT 2.505 3.245 2.675 3.415 ;
        RECT 3.985 3.245 4.155 3.415 ;
      LAYER met1 ;
        RECT 2.475 3.415 2.705 3.445 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 2.445 3.245 4.215 3.415 ;
        RECT 2.475 3.215 2.705 3.245 ;
        RECT 3.955 3.215 4.185 3.245 ;
  END
END AND2X1






MACRO AND3X1
  CLASS CORE ;
  FOREIGN AND3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.810 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 7.465 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 7.200 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.400 5.185 5.570 7.230 ;
        RECT 6.280 5.185 6.450 7.230 ;
        RECT 6.860 4.110 7.200 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 7.200 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 7.200 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.355 0.620 5.525 1.750 ;
        RECT 6.325 0.620 6.495 1.750 ;
        RECT 5.355 0.450 6.495 0.620 ;
        RECT 5.355 0.170 5.525 0.450 ;
        RECT 5.840 0.170 6.010 0.450 ;
        RECT 6.325 0.170 6.495 0.450 ;
        RECT 6.860 0.170 7.200 2.720 ;
        RECT -0.170 -0.170 7.200 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 7.200 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.465 1.920 5.635 4.865 ;
        RECT 5.840 4.665 6.010 7.020 ;
        RECT 5.840 4.495 6.375 4.665 ;
        RECT 6.205 2.165 6.375 4.495 ;
        RECT 5.835 1.995 6.375 2.165 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 5.835 0.840 6.005 1.995 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
      LAYER mcon ;
        RECT 3.985 3.245 4.155 3.415 ;
        RECT 5.465 3.245 5.635 3.415 ;
      LAYER met1 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 5.435 3.415 5.665 3.445 ;
        RECT 3.925 3.245 5.695 3.415 ;
        RECT 3.955 3.215 4.185 3.245 ;
        RECT 5.435 3.215 5.665 3.245 ;
  END
END AND3X1






MACRO AO3X1
  CLASS CORE ;
  FOREIGN AO3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.880 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 9.315 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 9.050 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.475 5.555 4.645 7.230 ;
        RECT 6.490 4.110 6.830 7.230 ;
        RECT 7.250 5.185 7.420 7.230 ;
        RECT 8.130 5.185 8.300 7.230 ;
        RECT 8.710 4.110 9.050 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 9.050 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 9.050 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 3.940 0.615 4.110 1.745 ;
        RECT 4.910 0.615 5.080 1.390 ;
        RECT 5.880 0.615 6.050 1.390 ;
        RECT 3.940 0.445 6.050 0.615 ;
        RECT 3.940 0.170 4.110 0.445 ;
        RECT 4.425 0.170 4.595 0.445 ;
        RECT 4.910 0.170 5.080 0.445 ;
        RECT 5.395 0.170 5.565 0.445 ;
        RECT 5.880 0.170 6.050 0.445 ;
        RECT 6.490 0.170 6.830 2.720 ;
        RECT 7.205 0.620 7.375 1.750 ;
        RECT 8.175 0.620 8.345 1.750 ;
        RECT 7.205 0.450 8.345 0.620 ;
        RECT 7.205 0.170 7.375 0.450 ;
        RECT 7.690 0.170 7.860 0.450 ;
        RECT 8.175 0.170 8.345 0.450 ;
        RECT 8.710 0.170 9.050 2.720 ;
        RECT -0.170 -0.170 9.050 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 9.050 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 4.035 5.295 4.205 7.025 ;
        RECT 4.915 6.825 5.965 6.995 ;
        RECT 4.915 5.295 5.085 6.825 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 4.035 5.125 5.085 5.295 ;
        RECT 5.355 5.295 5.525 6.565 ;
        RECT 5.795 5.555 5.965 6.825 ;
        RECT 5.355 5.125 6.005 5.295 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.200 4.710 4.370 4.870 ;
        RECT 5.130 4.710 5.300 4.870 ;
        RECT 4.200 4.540 4.525 4.710 ;
        RECT 4.355 1.915 4.525 4.540 ;
        RECT 5.095 4.540 5.300 4.710 ;
        RECT 5.095 1.915 5.265 4.540 ;
        RECT 5.835 1.740 6.005 5.125 ;
        RECT 7.315 1.920 7.485 4.865 ;
        RECT 7.690 4.665 7.860 7.020 ;
        RECT 7.690 4.495 8.225 4.665 ;
        RECT 8.055 2.165 8.225 4.495 ;
        RECT 7.685 1.995 8.225 2.165 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 4.425 1.570 6.005 1.740 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 4.425 0.835 4.595 1.570 ;
        RECT 5.395 0.835 5.565 1.570 ;
        RECT 7.685 0.840 7.855 1.995 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 7.315 2.505 7.485 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 7.285 2.675 7.515 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 5.775 2.505 7.545 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 7.285 2.475 7.515 2.505 ;
  END
END AO3X1






MACRO AOA4X1
  CLASS CORE ;
  FOREIGN AOA4X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.210 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 12.645 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 12.380 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.475 5.555 4.645 7.230 ;
        RECT 6.490 4.110 6.830 7.230 ;
        RECT 7.365 5.135 7.535 7.230 ;
        RECT 8.245 5.555 8.415 7.230 ;
        RECT 9.125 5.555 9.295 7.230 ;
        RECT 9.820 4.110 10.160 7.230 ;
        RECT 10.580 5.185 10.750 7.230 ;
        RECT 11.460 5.185 11.630 7.230 ;
        RECT 12.040 4.110 12.380 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 12.380 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 12.380 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 3.940 0.615 4.110 1.745 ;
        RECT 4.910 0.615 5.080 1.390 ;
        RECT 5.880 0.615 6.050 1.390 ;
        RECT 3.940 0.445 6.050 0.615 ;
        RECT 3.940 0.170 4.110 0.445 ;
        RECT 4.425 0.170 4.595 0.445 ;
        RECT 4.910 0.170 5.080 0.445 ;
        RECT 5.395 0.170 5.565 0.445 ;
        RECT 5.880 0.170 6.050 0.445 ;
        RECT 6.490 0.170 6.830 2.720 ;
        RECT 7.755 0.170 7.925 1.120 ;
        RECT 9.820 0.170 10.160 2.720 ;
        RECT 10.535 0.620 10.705 1.750 ;
        RECT 11.505 0.620 11.675 1.750 ;
        RECT 10.535 0.450 11.675 0.620 ;
        RECT 10.535 0.170 10.705 0.450 ;
        RECT 11.020 0.170 11.190 0.450 ;
        RECT 11.505 0.170 11.675 0.450 ;
        RECT 12.040 0.170 12.380 2.720 ;
        RECT -0.170 -0.170 12.380 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 12.380 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 4.035 5.295 4.205 7.025 ;
        RECT 4.915 6.825 5.965 6.995 ;
        RECT 4.915 5.295 5.085 6.825 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 4.035 5.125 5.085 5.295 ;
        RECT 5.355 5.295 5.525 6.565 ;
        RECT 5.795 5.555 5.965 6.825 ;
        RECT 5.355 5.125 6.005 5.295 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.200 4.710 4.370 4.870 ;
        RECT 5.130 4.710 5.300 4.870 ;
        RECT 4.200 4.540 4.525 4.710 ;
        RECT 4.355 1.915 4.525 4.540 ;
        RECT 5.095 4.540 5.300 4.710 ;
        RECT 5.095 1.915 5.265 4.540 ;
        RECT 5.835 1.740 6.005 5.125 ;
        RECT 7.805 5.285 7.975 7.020 ;
        RECT 8.685 5.285 8.855 7.020 ;
        RECT 7.805 5.115 9.335 5.285 ;
        RECT 7.685 1.915 7.855 4.865 ;
        RECT 8.455 4.710 8.625 4.865 ;
        RECT 8.425 4.535 8.625 4.710 ;
        RECT 8.425 1.915 8.595 4.535 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 4.425 1.570 6.005 1.740 ;
        RECT 7.270 1.665 7.440 1.745 ;
        RECT 8.240 1.665 8.410 1.745 ;
        RECT 9.165 1.740 9.335 5.115 ;
        RECT 10.645 1.920 10.815 4.865 ;
        RECT 11.020 4.665 11.190 7.020 ;
        RECT 11.020 4.495 11.555 4.665 ;
        RECT 11.385 2.165 11.555 4.495 ;
        RECT 11.015 1.995 11.555 2.165 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 4.425 0.835 4.595 1.570 ;
        RECT 5.395 0.835 5.565 1.570 ;
        RECT 7.270 1.495 8.410 1.665 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 7.270 0.365 7.440 1.495 ;
        RECT 8.240 0.615 8.410 1.495 ;
        RECT 8.725 1.570 9.335 1.740 ;
        RECT 8.725 0.835 8.895 1.570 ;
        RECT 9.210 0.615 9.380 1.385 ;
        RECT 11.015 0.840 11.185 1.995 ;
        RECT 8.240 0.445 9.380 0.615 ;
        RECT 8.240 0.365 8.410 0.445 ;
        RECT 9.210 0.365 9.380 0.445 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 7.685 2.505 7.855 2.675 ;
        RECT 9.165 2.505 9.335 2.675 ;
        RECT 10.645 2.505 10.815 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 9.135 2.675 9.365 2.705 ;
        RECT 10.615 2.675 10.845 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 5.775 2.505 7.915 2.675 ;
        RECT 9.105 2.505 10.875 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
        RECT 9.135 2.475 9.365 2.505 ;
        RECT 10.615 2.475 10.845 2.505 ;
  END
END AOA4X1






MACRO AOAI4X1
  CLASS CORE ;
  FOREIGN AOAI4X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.990 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 10.425 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 10.160 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.475 5.555 4.645 7.230 ;
        RECT 6.490 4.110 6.830 7.230 ;
        RECT 7.365 5.135 7.535 7.230 ;
        RECT 8.245 5.555 8.415 7.230 ;
        RECT 9.125 5.555 9.295 7.230 ;
        RECT 9.820 4.110 10.160 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 10.160 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 10.160 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 3.940 0.615 4.110 1.745 ;
        RECT 4.910 0.615 5.080 1.390 ;
        RECT 5.880 0.615 6.050 1.390 ;
        RECT 3.940 0.445 6.050 0.615 ;
        RECT 3.940 0.170 4.110 0.445 ;
        RECT 4.425 0.170 4.595 0.445 ;
        RECT 4.910 0.170 5.080 0.445 ;
        RECT 5.395 0.170 5.565 0.445 ;
        RECT 5.880 0.170 6.050 0.445 ;
        RECT 6.490 0.170 6.830 2.720 ;
        RECT 7.755 0.170 7.925 1.120 ;
        RECT 9.820 0.170 10.160 2.720 ;
        RECT -0.170 -0.170 10.160 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 10.160 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 4.035 5.295 4.205 7.025 ;
        RECT 4.915 6.825 5.965 6.995 ;
        RECT 4.915 5.295 5.085 6.825 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 4.035 5.125 5.085 5.295 ;
        RECT 5.355 5.295 5.525 6.565 ;
        RECT 5.795 5.555 5.965 6.825 ;
        RECT 5.355 5.125 6.005 5.295 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.200 4.710 4.370 4.870 ;
        RECT 5.130 4.710 5.300 4.870 ;
        RECT 4.200 4.540 4.525 4.710 ;
        RECT 4.355 1.915 4.525 4.540 ;
        RECT 5.095 4.540 5.300 4.710 ;
        RECT 5.095 1.915 5.265 4.540 ;
        RECT 5.835 1.740 6.005 5.125 ;
        RECT 7.805 5.285 7.975 7.020 ;
        RECT 8.685 5.285 8.855 7.020 ;
        RECT 7.805 5.115 9.335 5.285 ;
        RECT 7.685 1.915 7.855 4.865 ;
        RECT 8.455 4.710 8.625 4.865 ;
        RECT 8.425 4.535 8.625 4.710 ;
        RECT 8.425 1.915 8.595 4.535 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 4.425 1.570 6.005 1.740 ;
        RECT 7.270 1.665 7.440 1.745 ;
        RECT 8.240 1.665 8.410 1.745 ;
        RECT 9.165 1.740 9.335 5.115 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 4.425 0.835 4.595 1.570 ;
        RECT 5.395 0.835 5.565 1.570 ;
        RECT 7.270 1.495 8.410 1.665 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 7.270 0.365 7.440 1.495 ;
        RECT 8.240 0.615 8.410 1.495 ;
        RECT 8.725 1.570 9.335 1.740 ;
        RECT 8.725 0.835 8.895 1.570 ;
        RECT 9.210 0.615 9.380 1.385 ;
        RECT 8.240 0.445 9.380 0.615 ;
        RECT 8.240 0.365 8.410 0.445 ;
        RECT 9.210 0.365 9.380 0.445 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 7.685 2.505 7.855 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 5.775 2.505 7.915 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
  END
END AOAI4X1






MACRO AOI3X1
  CLASS CORE ;
  FOREIGN AOI3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.660 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 7.095 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 6.830 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.475 5.555 4.645 7.230 ;
        RECT 6.490 4.110 6.830 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 6.830 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 6.830 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 3.940 0.615 4.110 1.745 ;
        RECT 4.910 0.615 5.080 1.390 ;
        RECT 5.880 0.615 6.050 1.390 ;
        RECT 3.940 0.445 6.050 0.615 ;
        RECT 3.940 0.170 4.110 0.445 ;
        RECT 4.425 0.170 4.595 0.445 ;
        RECT 4.910 0.170 5.080 0.445 ;
        RECT 5.395 0.170 5.565 0.445 ;
        RECT 5.880 0.170 6.050 0.445 ;
        RECT 6.490 0.170 6.830 2.720 ;
        RECT -0.170 -0.170 6.830 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 6.830 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 4.035 5.295 4.205 7.025 ;
        RECT 4.915 6.825 5.965 6.995 ;
        RECT 4.915 5.295 5.085 6.825 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 4.035 5.125 5.085 5.295 ;
        RECT 5.355 5.295 5.525 6.565 ;
        RECT 5.795 5.555 5.965 6.825 ;
        RECT 5.355 5.125 6.005 5.295 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.200 4.710 4.370 4.870 ;
        RECT 5.130 4.710 5.300 4.870 ;
        RECT 4.200 4.540 4.525 4.710 ;
        RECT 4.355 1.915 4.525 4.540 ;
        RECT 5.095 4.540 5.300 4.710 ;
        RECT 5.095 1.915 5.265 4.540 ;
        RECT 5.835 1.740 6.005 5.125 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 4.425 1.570 6.005 1.740 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 4.425 0.835 4.595 1.570 ;
        RECT 5.395 0.835 5.565 1.570 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
  END
END AOI3X1






MACRO BUFX1
  CLASS CORE ;
  FOREIGN BUFX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.440 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 4.875 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 4.610 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
        RECT 2.810 5.185 2.980 7.230 ;
        RECT 3.690 5.185 3.860 7.230 ;
        RECT 4.270 4.110 4.610 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 4.610 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 4.610 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT 2.765 0.620 2.935 1.750 ;
        RECT 3.735 0.620 3.905 1.750 ;
        RECT 2.765 0.450 3.905 0.620 ;
        RECT 2.765 0.170 2.935 0.450 ;
        RECT 3.250 0.170 3.420 0.450 ;
        RECT 3.735 0.170 3.905 0.450 ;
        RECT 4.270 0.170 4.610 2.720 ;
        RECT -0.170 -0.170 4.610 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 4.610 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
        RECT 2.875 1.920 3.045 4.865 ;
        RECT 3.250 4.665 3.420 7.020 ;
        RECT 3.250 4.495 3.785 4.665 ;
        RECT 3.615 2.165 3.785 4.495 ;
        RECT 3.245 1.995 3.785 2.165 ;
        RECT 3.245 0.840 3.415 1.995 ;
      LAYER mcon ;
        RECT 1.395 2.505 1.565 2.675 ;
        RECT 2.875 2.505 3.045 2.675 ;
      LAYER met1 ;
        RECT 1.365 2.675 1.595 2.705 ;
        RECT 2.845 2.675 3.075 2.705 ;
        RECT 1.335 2.505 3.105 2.675 ;
        RECT 1.365 2.475 1.595 2.505 ;
        RECT 2.845 2.475 3.075 2.505 ;
  END
END BUFX1






MACRO DFFQNX1
  CLASS CORE ;
  FOREIGN DFFQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.460 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 15.945 5.285 16.115 7.020 ;
        RECT 16.825 5.285 16.995 7.020 ;
        RECT 15.945 5.115 17.475 5.285 ;
        RECT 17.305 1.740 17.475 5.115 ;
        RECT 19.155 1.915 19.325 4.865 ;
        RECT 16.865 1.570 17.475 1.740 ;
        RECT 16.865 0.835 17.035 1.570 ;
      LAYER mcon ;
        RECT 17.305 3.245 17.475 3.415 ;
        RECT 19.155 3.245 19.325 3.415 ;
      LAYER met1 ;
        RECT 17.275 3.415 17.505 3.445 ;
        RECT 19.125 3.415 19.355 3.445 ;
        RECT 17.245 3.245 19.385 3.415 ;
        RECT 17.275 3.215 17.505 3.245 ;
        RECT 19.125 3.215 19.355 3.245 ;
    END
  END QN
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 13.265 4.710 13.435 4.865 ;
        RECT 13.235 4.535 13.435 4.710 ;
        RECT 13.235 1.915 13.405 4.535 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 13.235 4.355 13.405 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 13.205 4.525 13.435 4.555 ;
        RECT 2.075 4.355 13.465 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 13.205 4.325 13.435 4.355 ;
    END
  END CLK
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 21.895 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 21.630 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.515 5.135 5.685 7.230 ;
        RECT 6.395 5.555 6.565 7.230 ;
        RECT 7.275 5.555 7.445 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 8.845 5.135 9.015 7.230 ;
        RECT 9.725 5.555 9.895 7.230 ;
        RECT 10.605 5.555 10.775 7.230 ;
        RECT 11.300 4.110 11.640 7.230 ;
        RECT 12.175 5.135 12.345 7.230 ;
        RECT 13.055 5.555 13.225 7.230 ;
        RECT 13.935 5.555 14.105 7.230 ;
        RECT 14.630 4.110 14.970 7.230 ;
        RECT 15.505 5.135 15.675 7.230 ;
        RECT 16.385 5.555 16.555 7.230 ;
        RECT 17.265 5.555 17.435 7.230 ;
        RECT 17.960 4.110 18.300 7.230 ;
        RECT 18.835 5.135 19.005 7.230 ;
        RECT 19.715 5.555 19.885 7.230 ;
        RECT 20.595 5.555 20.765 7.230 ;
        RECT 21.290 4.110 21.630 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 21.630 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 21.630 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.905 0.170 6.075 1.120 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.235 0.170 9.405 1.120 ;
        RECT 11.300 0.170 11.640 2.720 ;
        RECT 12.565 0.170 12.735 1.120 ;
        RECT 14.630 0.170 14.970 2.720 ;
        RECT 15.895 0.170 16.065 1.120 ;
        RECT 17.960 0.170 18.300 2.720 ;
        RECT 19.225 0.170 19.395 1.120 ;
        RECT 21.290 0.170 21.630 2.720 ;
        RECT -0.170 -0.170 21.630 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 21.630 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 5.955 5.285 6.125 7.020 ;
        RECT 6.835 5.285 7.005 7.020 ;
        RECT 9.285 5.285 9.455 7.020 ;
        RECT 10.165 5.285 10.335 7.020 ;
        RECT 12.615 5.285 12.785 7.020 ;
        RECT 13.495 5.285 13.665 7.020 ;
        RECT 19.275 5.285 19.445 7.020 ;
        RECT 20.155 5.285 20.325 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 5.955 5.115 7.485 5.285 ;
        RECT 9.285 5.115 10.815 5.285 ;
        RECT 12.615 5.115 14.145 5.285 ;
        RECT 19.275 5.115 20.805 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 6.605 4.710 6.775 4.865 ;
        RECT 6.575 4.535 6.775 4.710 ;
        RECT 6.575 1.915 6.745 4.535 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.420 1.665 5.590 1.745 ;
        RECT 6.390 1.665 6.560 1.745 ;
        RECT 7.315 1.740 7.485 5.115 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 9.935 4.710 10.105 4.865 ;
        RECT 9.905 4.535 10.105 4.710 ;
        RECT 9.905 1.915 10.075 4.535 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.420 1.495 6.560 1.665 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.420 0.365 5.590 1.495 ;
        RECT 6.390 0.615 6.560 1.495 ;
        RECT 6.875 1.570 7.485 1.740 ;
        RECT 8.750 1.665 8.920 1.745 ;
        RECT 9.720 1.665 9.890 1.745 ;
        RECT 10.645 1.740 10.815 5.115 ;
        RECT 12.495 1.915 12.665 4.865 ;
        RECT 6.875 0.835 7.045 1.570 ;
        RECT 8.750 1.495 9.890 1.665 ;
        RECT 7.360 0.615 7.530 1.385 ;
        RECT 6.390 0.445 7.530 0.615 ;
        RECT 6.390 0.365 6.560 0.445 ;
        RECT 7.360 0.365 7.530 0.445 ;
        RECT 8.750 0.365 8.920 1.495 ;
        RECT 9.720 0.615 9.890 1.495 ;
        RECT 10.205 1.570 10.815 1.740 ;
        RECT 12.080 1.665 12.250 1.745 ;
        RECT 13.050 1.665 13.220 1.745 ;
        RECT 13.975 1.740 14.145 5.115 ;
        RECT 15.825 1.915 15.995 4.865 ;
        RECT 16.595 4.710 16.765 4.865 ;
        RECT 19.925 4.710 20.095 4.865 ;
        RECT 16.565 4.535 16.765 4.710 ;
        RECT 19.895 4.535 20.095 4.710 ;
        RECT 16.565 1.915 16.735 4.535 ;
        RECT 19.895 1.915 20.065 4.535 ;
        RECT 10.205 0.835 10.375 1.570 ;
        RECT 12.080 1.495 13.220 1.665 ;
        RECT 10.690 0.615 10.860 1.385 ;
        RECT 9.720 0.445 10.860 0.615 ;
        RECT 9.720 0.365 9.890 0.445 ;
        RECT 10.690 0.365 10.860 0.445 ;
        RECT 12.080 0.365 12.250 1.495 ;
        RECT 13.050 0.615 13.220 1.495 ;
        RECT 13.535 1.570 14.145 1.740 ;
        RECT 15.410 1.665 15.580 1.745 ;
        RECT 16.380 1.665 16.550 1.745 ;
        RECT 13.535 0.835 13.705 1.570 ;
        RECT 15.410 1.495 16.550 1.665 ;
        RECT 14.020 0.615 14.190 1.385 ;
        RECT 13.050 0.445 14.190 0.615 ;
        RECT 13.050 0.365 13.220 0.445 ;
        RECT 14.020 0.365 14.190 0.445 ;
        RECT 15.410 0.365 15.580 1.495 ;
        RECT 16.380 0.615 16.550 1.495 ;
        RECT 18.740 1.665 18.910 1.745 ;
        RECT 19.710 1.665 19.880 1.745 ;
        RECT 20.635 1.740 20.805 5.115 ;
        RECT 18.740 1.495 19.880 1.665 ;
        RECT 17.350 0.615 17.520 1.385 ;
        RECT 16.380 0.445 17.520 0.615 ;
        RECT 16.380 0.365 16.550 0.445 ;
        RECT 17.350 0.365 17.520 0.445 ;
        RECT 18.740 0.365 18.910 1.495 ;
        RECT 19.710 0.615 19.880 1.495 ;
        RECT 20.195 1.570 20.805 1.740 ;
        RECT 20.195 0.835 20.365 1.570 ;
        RECT 20.680 0.615 20.850 1.385 ;
        RECT 19.710 0.445 20.850 0.615 ;
        RECT 19.710 0.365 19.880 0.445 ;
        RECT 20.680 0.365 20.850 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 7.315 3.245 7.485 3.415 ;
        RECT 9.165 3.245 9.335 3.415 ;
        RECT 9.905 3.985 10.075 4.155 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 12.495 3.245 12.665 3.415 ;
        RECT 13.975 3.985 14.145 4.155 ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 16.565 3.615 16.735 3.785 ;
        RECT 19.895 3.985 20.065 4.155 ;
        RECT 20.635 3.615 20.805 3.785 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 9.875 4.155 10.105 4.185 ;
        RECT 13.945 4.155 14.175 4.185 ;
        RECT 19.865 4.155 20.095 4.185 ;
        RECT 0.965 3.985 20.125 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 9.875 3.955 10.105 3.985 ;
        RECT 13.945 3.955 14.175 3.985 ;
        RECT 19.865 3.955 20.095 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 16.535 3.785 16.765 3.815 ;
        RECT 20.605 3.785 20.835 3.815 ;
        RECT 3.925 3.615 16.055 3.785 ;
        RECT 16.505 3.615 20.865 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 16.535 3.585 16.765 3.615 ;
        RECT 20.605 3.585 20.835 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 7.285 3.415 7.515 3.445 ;
        RECT 9.135 3.415 9.365 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.465 3.415 12.695 3.445 ;
        RECT 3.185 3.245 9.395 3.415 ;
        RECT 10.585 3.245 12.725 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 7.285 3.215 7.515 3.245 ;
        RECT 9.135 3.215 9.365 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.465 3.215 12.695 3.245 ;
  END
END DFFQNX1






MACRO DFFQX1
  CLASS CORE ;
  FOREIGN DFFQX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.460 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 19.275 5.285 19.445 7.020 ;
        RECT 20.155 5.285 20.325 7.020 ;
        RECT 19.275 5.115 20.805 5.285 ;
        RECT 16.595 4.710 16.765 4.865 ;
        RECT 16.565 4.535 16.765 4.710 ;
        RECT 16.565 1.915 16.735 4.535 ;
        RECT 20.635 1.740 20.805 5.115 ;
        RECT 20.195 1.570 20.805 1.740 ;
        RECT 20.195 0.835 20.365 1.570 ;
      LAYER mcon ;
        RECT 16.565 3.615 16.735 3.785 ;
        RECT 20.635 3.615 20.805 3.785 ;
      LAYER met1 ;
        RECT 16.535 3.785 16.765 3.815 ;
        RECT 20.605 3.785 20.835 3.815 ;
        RECT 16.505 3.615 20.865 3.785 ;
        RECT 16.535 3.585 16.765 3.615 ;
        RECT 20.605 3.585 20.835 3.615 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 13.265 4.710 13.435 4.865 ;
        RECT 13.235 4.535 13.435 4.710 ;
        RECT 13.235 1.915 13.405 4.535 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 13.235 4.355 13.405 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 13.205 4.525 13.435 4.555 ;
        RECT 2.075 4.355 13.465 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 13.205 4.325 13.435 4.355 ;
    END
  END CLK
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 21.895 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 21.630 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.515 5.135 5.685 7.230 ;
        RECT 6.395 5.555 6.565 7.230 ;
        RECT 7.275 5.555 7.445 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 8.845 5.135 9.015 7.230 ;
        RECT 9.725 5.555 9.895 7.230 ;
        RECT 10.605 5.555 10.775 7.230 ;
        RECT 11.300 4.110 11.640 7.230 ;
        RECT 12.175 5.135 12.345 7.230 ;
        RECT 13.055 5.555 13.225 7.230 ;
        RECT 13.935 5.555 14.105 7.230 ;
        RECT 14.630 4.110 14.970 7.230 ;
        RECT 15.505 5.135 15.675 7.230 ;
        RECT 16.385 5.555 16.555 7.230 ;
        RECT 17.265 5.555 17.435 7.230 ;
        RECT 17.960 4.110 18.300 7.230 ;
        RECT 18.835 5.135 19.005 7.230 ;
        RECT 19.715 5.555 19.885 7.230 ;
        RECT 20.595 5.555 20.765 7.230 ;
        RECT 21.290 4.110 21.630 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 21.630 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 21.630 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.905 0.170 6.075 1.120 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.235 0.170 9.405 1.120 ;
        RECT 11.300 0.170 11.640 2.720 ;
        RECT 12.565 0.170 12.735 1.120 ;
        RECT 14.630 0.170 14.970 2.720 ;
        RECT 15.895 0.170 16.065 1.120 ;
        RECT 17.960 0.170 18.300 2.720 ;
        RECT 19.225 0.170 19.395 1.120 ;
        RECT 21.290 0.170 21.630 2.720 ;
        RECT -0.170 -0.170 21.630 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 21.630 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 5.955 5.285 6.125 7.020 ;
        RECT 6.835 5.285 7.005 7.020 ;
        RECT 9.285 5.285 9.455 7.020 ;
        RECT 10.165 5.285 10.335 7.020 ;
        RECT 12.615 5.285 12.785 7.020 ;
        RECT 13.495 5.285 13.665 7.020 ;
        RECT 15.945 5.285 16.115 7.020 ;
        RECT 16.825 5.285 16.995 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 5.955 5.115 7.485 5.285 ;
        RECT 9.285 5.115 10.815 5.285 ;
        RECT 12.615 5.115 14.145 5.285 ;
        RECT 15.945 5.115 17.475 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 6.605 4.710 6.775 4.865 ;
        RECT 6.575 4.535 6.775 4.710 ;
        RECT 6.575 1.915 6.745 4.535 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.420 1.665 5.590 1.745 ;
        RECT 6.390 1.665 6.560 1.745 ;
        RECT 7.315 1.740 7.485 5.115 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 9.935 4.710 10.105 4.865 ;
        RECT 9.905 4.535 10.105 4.710 ;
        RECT 9.905 1.915 10.075 4.535 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.420 1.495 6.560 1.665 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.420 0.365 5.590 1.495 ;
        RECT 6.390 0.615 6.560 1.495 ;
        RECT 6.875 1.570 7.485 1.740 ;
        RECT 8.750 1.665 8.920 1.745 ;
        RECT 9.720 1.665 9.890 1.745 ;
        RECT 10.645 1.740 10.815 5.115 ;
        RECT 12.495 1.915 12.665 4.865 ;
        RECT 6.875 0.835 7.045 1.570 ;
        RECT 8.750 1.495 9.890 1.665 ;
        RECT 7.360 0.615 7.530 1.385 ;
        RECT 6.390 0.445 7.530 0.615 ;
        RECT 6.390 0.365 6.560 0.445 ;
        RECT 7.360 0.365 7.530 0.445 ;
        RECT 8.750 0.365 8.920 1.495 ;
        RECT 9.720 0.615 9.890 1.495 ;
        RECT 10.205 1.570 10.815 1.740 ;
        RECT 12.080 1.665 12.250 1.745 ;
        RECT 13.050 1.665 13.220 1.745 ;
        RECT 13.975 1.740 14.145 5.115 ;
        RECT 15.825 1.915 15.995 4.865 ;
        RECT 10.205 0.835 10.375 1.570 ;
        RECT 12.080 1.495 13.220 1.665 ;
        RECT 10.690 0.615 10.860 1.385 ;
        RECT 9.720 0.445 10.860 0.615 ;
        RECT 9.720 0.365 9.890 0.445 ;
        RECT 10.690 0.365 10.860 0.445 ;
        RECT 12.080 0.365 12.250 1.495 ;
        RECT 13.050 0.615 13.220 1.495 ;
        RECT 13.535 1.570 14.145 1.740 ;
        RECT 15.410 1.665 15.580 1.745 ;
        RECT 16.380 1.665 16.550 1.745 ;
        RECT 17.305 1.740 17.475 5.115 ;
        RECT 19.155 1.915 19.325 4.865 ;
        RECT 19.925 4.710 20.095 4.865 ;
        RECT 19.895 4.535 20.095 4.710 ;
        RECT 19.895 1.915 20.065 4.535 ;
        RECT 13.535 0.835 13.705 1.570 ;
        RECT 15.410 1.495 16.550 1.665 ;
        RECT 14.020 0.615 14.190 1.385 ;
        RECT 13.050 0.445 14.190 0.615 ;
        RECT 13.050 0.365 13.220 0.445 ;
        RECT 14.020 0.365 14.190 0.445 ;
        RECT 15.410 0.365 15.580 1.495 ;
        RECT 16.380 0.615 16.550 1.495 ;
        RECT 16.865 1.570 17.475 1.740 ;
        RECT 18.740 1.665 18.910 1.745 ;
        RECT 19.710 1.665 19.880 1.745 ;
        RECT 16.865 0.835 17.035 1.570 ;
        RECT 18.740 1.495 19.880 1.665 ;
        RECT 17.350 0.615 17.520 1.385 ;
        RECT 16.380 0.445 17.520 0.615 ;
        RECT 16.380 0.365 16.550 0.445 ;
        RECT 17.350 0.365 17.520 0.445 ;
        RECT 18.740 0.365 18.910 1.495 ;
        RECT 19.710 0.615 19.880 1.495 ;
        RECT 20.680 0.615 20.850 1.385 ;
        RECT 19.710 0.445 20.850 0.615 ;
        RECT 19.710 0.365 19.880 0.445 ;
        RECT 20.680 0.365 20.850 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 7.315 3.245 7.485 3.415 ;
        RECT 9.165 3.245 9.335 3.415 ;
        RECT 9.905 3.985 10.075 4.155 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 12.495 3.245 12.665 3.415 ;
        RECT 13.975 3.985 14.145 4.155 ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 17.305 3.245 17.475 3.415 ;
        RECT 19.155 3.245 19.325 3.415 ;
        RECT 19.895 3.985 20.065 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 9.875 4.155 10.105 4.185 ;
        RECT 13.945 4.155 14.175 4.185 ;
        RECT 19.865 4.155 20.095 4.185 ;
        RECT 0.965 3.985 20.125 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 9.875 3.955 10.105 3.985 ;
        RECT 13.945 3.955 14.175 3.985 ;
        RECT 19.865 3.955 20.095 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 3.925 3.615 16.055 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 7.285 3.415 7.515 3.445 ;
        RECT 9.135 3.415 9.365 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.465 3.415 12.695 3.445 ;
        RECT 17.275 3.415 17.505 3.445 ;
        RECT 19.125 3.415 19.355 3.445 ;
        RECT 3.185 3.245 9.395 3.415 ;
        RECT 10.585 3.245 12.725 3.415 ;
        RECT 17.245 3.245 19.385 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 7.285 3.215 7.515 3.245 ;
        RECT 9.135 3.215 9.365 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.465 3.215 12.695 3.245 ;
        RECT 17.275 3.215 17.505 3.245 ;
        RECT 19.125 3.215 19.355 3.245 ;
  END
END DFFQX1






MACRO DFFRNQNX1
  CLASS CORE ;
  FOREIGN DFFRNQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.900 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 19.205 5.240 19.375 7.020 ;
        RECT 20.085 5.240 20.255 7.020 ;
        RECT 20.965 5.240 21.135 7.020 ;
        RECT 19.205 5.070 21.915 5.240 ;
        RECT 21.745 1.750 21.915 5.070 ;
        RECT 23.595 1.915 23.765 4.865 ;
        RECT 21.260 1.580 21.915 1.750 ;
        RECT 21.260 0.845 21.430 1.580 ;
      LAYER mcon ;
        RECT 21.745 3.245 21.915 3.415 ;
        RECT 23.595 3.245 23.765 3.415 ;
      LAYER met1 ;
        RECT 21.715 3.415 21.945 3.445 ;
        RECT 23.565 3.415 23.795 3.445 ;
        RECT 21.685 3.245 23.825 3.415 ;
        RECT 21.715 3.215 21.945 3.245 ;
        RECT 23.565 3.215 23.795 3.245 ;
    END
  END QN
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 15.085 1.915 15.255 4.865 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 15.085 4.355 15.255 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 15.055 4.525 15.285 4.555 ;
        RECT 2.075 4.355 15.315 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 15.055 4.325 15.285 4.355 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 3.069350 ;
    PORT
      LAYER li1 ;
        RECT 8.055 1.915 8.225 4.865 ;
        RECT 16.195 1.915 16.365 4.865 ;
        RECT 19.895 1.915 20.065 4.865 ;
      LAYER mcon ;
        RECT 8.055 2.135 8.225 2.305 ;
        RECT 16.195 2.135 16.365 2.305 ;
        RECT 19.895 2.135 20.065 2.305 ;
      LAYER met1 ;
        RECT 8.025 2.305 8.255 2.335 ;
        RECT 16.165 2.305 16.395 2.335 ;
        RECT 19.865 2.305 20.095 2.335 ;
        RECT 7.995 2.135 20.125 2.305 ;
        RECT 8.025 2.105 8.255 2.135 ;
        RECT 16.165 2.105 16.395 2.135 ;
        RECT 19.865 2.105 20.095 2.135 ;
    END
  END RN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 26.335 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 26.070 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.325 5.135 10.495 7.230 ;
        RECT 11.205 5.555 11.375 7.230 ;
        RECT 12.085 5.555 12.255 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.955 5.215 14.125 7.230 ;
        RECT 14.835 5.555 15.005 7.230 ;
        RECT 15.715 5.555 15.885 7.230 ;
        RECT 16.595 5.555 16.765 7.230 ;
        RECT 17.590 4.110 17.930 7.230 ;
        RECT 18.765 5.215 18.935 7.230 ;
        RECT 19.645 5.555 19.815 7.230 ;
        RECT 20.525 5.555 20.695 7.230 ;
        RECT 21.405 5.555 21.575 7.230 ;
        RECT 22.400 4.110 22.740 7.230 ;
        RECT 23.275 5.135 23.445 7.230 ;
        RECT 24.155 5.555 24.325 7.230 ;
        RECT 25.035 5.555 25.205 7.230 ;
        RECT 25.730 4.110 26.070 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 26.070 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 26.070 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.715 0.170 10.885 1.120 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 13.940 0.170 14.110 1.130 ;
        RECT 17.590 0.170 17.930 2.720 ;
        RECT 18.750 0.170 18.920 1.130 ;
        RECT 22.400 0.170 22.740 2.720 ;
        RECT 23.665 0.170 23.835 1.120 ;
        RECT 25.730 0.170 26.070 2.720 ;
        RECT -0.170 -0.170 26.070 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 26.070 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 10.765 5.285 10.935 7.020 ;
        RECT 11.645 5.285 11.815 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 10.765 5.115 12.295 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 11.415 4.710 11.585 4.865 ;
        RECT 11.385 4.535 11.585 4.710 ;
        RECT 11.385 1.915 11.555 4.535 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.230 1.665 10.400 1.745 ;
        RECT 11.200 1.665 11.370 1.745 ;
        RECT 12.125 1.740 12.295 5.115 ;
        RECT 14.395 5.240 14.565 7.020 ;
        RECT 15.275 5.240 15.445 7.020 ;
        RECT 16.155 5.240 16.325 7.020 ;
        RECT 23.715 5.285 23.885 7.020 ;
        RECT 24.595 5.285 24.765 7.020 ;
        RECT 14.395 5.070 17.105 5.240 ;
        RECT 23.715 5.115 25.245 5.285 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.230 1.495 11.370 1.665 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.230 0.365 10.400 1.495 ;
        RECT 11.200 0.615 11.370 1.495 ;
        RECT 11.685 1.570 12.295 1.740 ;
        RECT 13.455 1.675 13.625 1.755 ;
        RECT 14.425 1.675 14.595 1.755 ;
        RECT 15.395 1.675 15.565 1.755 ;
        RECT 11.685 0.835 11.855 1.570 ;
        RECT 13.455 1.505 15.565 1.675 ;
        RECT 12.170 0.615 12.340 1.385 ;
        RECT 11.200 0.445 12.340 0.615 ;
        RECT 11.200 0.365 11.370 0.445 ;
        RECT 12.170 0.365 12.340 0.445 ;
        RECT 13.455 0.375 13.625 1.505 ;
        RECT 14.425 0.625 14.595 1.505 ;
        RECT 15.395 1.425 15.565 1.505 ;
        RECT 14.915 1.080 15.085 1.160 ;
        RECT 15.965 1.080 16.135 1.755 ;
        RECT 16.935 1.750 17.105 5.070 ;
        RECT 18.785 1.915 18.955 4.865 ;
        RECT 21.005 1.915 21.175 4.865 ;
        RECT 24.365 4.710 24.535 4.865 ;
        RECT 24.335 4.535 24.535 4.710 ;
        RECT 24.335 1.915 24.505 4.535 ;
        RECT 14.915 0.910 16.135 1.080 ;
        RECT 14.915 0.830 15.085 0.910 ;
        RECT 15.395 0.625 15.565 0.705 ;
        RECT 14.425 0.455 15.565 0.625 ;
        RECT 14.425 0.375 14.595 0.455 ;
        RECT 15.395 0.375 15.565 0.455 ;
        RECT 15.965 0.625 16.135 0.910 ;
        RECT 16.450 1.580 17.105 1.750 ;
        RECT 18.265 1.675 18.435 1.755 ;
        RECT 19.235 1.675 19.405 1.755 ;
        RECT 20.205 1.675 20.375 1.755 ;
        RECT 16.450 0.845 16.620 1.580 ;
        RECT 18.265 1.505 20.375 1.675 ;
        RECT 16.935 0.625 17.105 1.395 ;
        RECT 15.965 0.455 17.105 0.625 ;
        RECT 15.965 0.375 16.135 0.455 ;
        RECT 16.935 0.375 17.105 0.455 ;
        RECT 18.265 0.375 18.435 1.505 ;
        RECT 19.235 0.625 19.405 1.505 ;
        RECT 20.205 1.425 20.375 1.505 ;
        RECT 19.725 1.080 19.895 1.160 ;
        RECT 20.775 1.080 20.945 1.755 ;
        RECT 23.180 1.665 23.350 1.745 ;
        RECT 24.150 1.665 24.320 1.745 ;
        RECT 25.075 1.740 25.245 5.115 ;
        RECT 23.180 1.495 24.320 1.665 ;
        RECT 19.725 0.910 20.945 1.080 ;
        RECT 19.725 0.830 19.895 0.910 ;
        RECT 20.205 0.625 20.375 0.705 ;
        RECT 19.235 0.455 20.375 0.625 ;
        RECT 19.235 0.375 19.405 0.455 ;
        RECT 20.205 0.375 20.375 0.455 ;
        RECT 20.775 0.625 20.945 0.910 ;
        RECT 21.745 0.625 21.915 1.395 ;
        RECT 20.775 0.455 21.915 0.625 ;
        RECT 20.775 0.375 20.945 0.455 ;
        RECT 21.745 0.375 21.915 0.455 ;
        RECT 23.180 0.365 23.350 1.495 ;
        RECT 24.150 0.615 24.320 1.495 ;
        RECT 24.635 1.570 25.245 1.740 ;
        RECT 24.635 0.835 24.805 1.570 ;
        RECT 25.120 0.615 25.290 1.385 ;
        RECT 24.150 0.445 25.290 0.615 ;
        RECT 24.150 0.365 24.320 0.445 ;
        RECT 25.120 0.365 25.290 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 3.245 12.295 3.415 ;
        RECT 13.975 3.245 14.145 3.415 ;
        RECT 16.935 3.985 17.105 4.155 ;
        RECT 18.785 3.615 18.955 3.785 ;
        RECT 21.005 3.615 21.175 3.785 ;
        RECT 24.335 3.985 24.505 4.155 ;
        RECT 25.075 3.615 25.245 3.785 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 16.905 4.155 17.135 4.185 ;
        RECT 24.305 4.155 24.535 4.185 ;
        RECT 0.965 3.985 24.565 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 16.905 3.955 17.135 3.985 ;
        RECT 24.305 3.955 24.535 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 18.755 3.785 18.985 3.815 ;
        RECT 20.975 3.785 21.205 3.815 ;
        RECT 25.045 3.785 25.275 3.815 ;
        RECT 3.925 3.615 19.015 3.785 ;
        RECT 20.945 3.615 25.305 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 18.755 3.585 18.985 3.615 ;
        RECT 20.975 3.585 21.205 3.615 ;
        RECT 25.045 3.585 25.275 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 8.765 3.415 8.995 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.095 3.415 12.325 3.445 ;
        RECT 13.945 3.415 14.175 3.445 ;
        RECT 3.185 3.245 10.875 3.415 ;
        RECT 12.065 3.245 14.205 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 8.765 3.215 8.995 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.095 3.215 12.325 3.245 ;
        RECT 13.945 3.215 14.175 3.245 ;
  END
END DFFRNQNX1






MACRO DFFRNQX1
  CLASS CORE ;
  FOREIGN DFFRNQX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.900 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 23.715 5.285 23.885 7.020 ;
        RECT 24.595 5.285 24.765 7.020 ;
        RECT 23.715 5.115 25.245 5.285 ;
        RECT 21.005 1.915 21.175 4.865 ;
        RECT 25.075 1.740 25.245 5.115 ;
        RECT 24.635 1.570 25.245 1.740 ;
        RECT 24.635 0.835 24.805 1.570 ;
      LAYER mcon ;
        RECT 21.005 3.615 21.175 3.785 ;
        RECT 25.075 3.615 25.245 3.785 ;
      LAYER met1 ;
        RECT 20.975 3.785 21.205 3.815 ;
        RECT 25.045 3.785 25.275 3.815 ;
        RECT 20.945 3.615 25.305 3.785 ;
        RECT 20.975 3.585 21.205 3.615 ;
        RECT 25.045 3.585 25.275 3.615 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 15.085 1.915 15.255 4.865 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 15.085 4.355 15.255 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 15.055 4.525 15.285 4.555 ;
        RECT 2.075 4.355 15.315 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 15.055 4.325 15.285 4.355 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 3.069350 ;
    PORT
      LAYER li1 ;
        RECT 8.055 1.915 8.225 4.865 ;
        RECT 16.195 1.915 16.365 4.865 ;
        RECT 19.895 1.915 20.065 4.865 ;
      LAYER mcon ;
        RECT 8.055 2.135 8.225 2.305 ;
        RECT 16.195 2.135 16.365 2.305 ;
        RECT 19.895 2.135 20.065 2.305 ;
      LAYER met1 ;
        RECT 8.025 2.305 8.255 2.335 ;
        RECT 16.165 2.305 16.395 2.335 ;
        RECT 19.865 2.305 20.095 2.335 ;
        RECT 7.995 2.135 20.125 2.305 ;
        RECT 8.025 2.105 8.255 2.135 ;
        RECT 16.165 2.105 16.395 2.135 ;
        RECT 19.865 2.105 20.095 2.135 ;
    END
  END RN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 26.335 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 26.070 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.325 5.135 10.495 7.230 ;
        RECT 11.205 5.555 11.375 7.230 ;
        RECT 12.085 5.555 12.255 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.955 5.215 14.125 7.230 ;
        RECT 14.835 5.555 15.005 7.230 ;
        RECT 15.715 5.555 15.885 7.230 ;
        RECT 16.595 5.555 16.765 7.230 ;
        RECT 17.590 4.110 17.930 7.230 ;
        RECT 18.765 5.215 18.935 7.230 ;
        RECT 19.645 5.555 19.815 7.230 ;
        RECT 20.525 5.555 20.695 7.230 ;
        RECT 21.405 5.555 21.575 7.230 ;
        RECT 22.400 4.110 22.740 7.230 ;
        RECT 23.275 5.135 23.445 7.230 ;
        RECT 24.155 5.555 24.325 7.230 ;
        RECT 25.035 5.555 25.205 7.230 ;
        RECT 25.730 4.110 26.070 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 26.070 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 26.070 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.715 0.170 10.885 1.120 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 13.940 0.170 14.110 1.130 ;
        RECT 17.590 0.170 17.930 2.720 ;
        RECT 18.750 0.170 18.920 1.130 ;
        RECT 22.400 0.170 22.740 2.720 ;
        RECT 23.665 0.170 23.835 1.120 ;
        RECT 25.730 0.170 26.070 2.720 ;
        RECT -0.170 -0.170 26.070 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 26.070 0.175 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 10.765 5.285 10.935 7.020 ;
        RECT 11.645 5.285 11.815 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 10.765 5.115 12.295 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 11.415 4.710 11.585 4.865 ;
        RECT 11.385 4.535 11.585 4.710 ;
        RECT 11.385 1.915 11.555 4.535 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.230 1.665 10.400 1.745 ;
        RECT 11.200 1.665 11.370 1.745 ;
        RECT 12.125 1.740 12.295 5.115 ;
        RECT 14.395 5.240 14.565 7.020 ;
        RECT 15.275 5.240 15.445 7.020 ;
        RECT 16.155 5.240 16.325 7.020 ;
        RECT 19.205 5.240 19.375 7.020 ;
        RECT 20.085 5.240 20.255 7.020 ;
        RECT 20.965 5.240 21.135 7.020 ;
        RECT 14.395 5.070 17.105 5.240 ;
        RECT 19.205 5.070 21.915 5.240 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.230 1.495 11.370 1.665 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.230 0.365 10.400 1.495 ;
        RECT 11.200 0.615 11.370 1.495 ;
        RECT 11.685 1.570 12.295 1.740 ;
        RECT 13.455 1.675 13.625 1.755 ;
        RECT 14.425 1.675 14.595 1.755 ;
        RECT 15.395 1.675 15.565 1.755 ;
        RECT 11.685 0.835 11.855 1.570 ;
        RECT 13.455 1.505 15.565 1.675 ;
        RECT 12.170 0.615 12.340 1.385 ;
        RECT 11.200 0.445 12.340 0.615 ;
        RECT 11.200 0.365 11.370 0.445 ;
        RECT 12.170 0.365 12.340 0.445 ;
        RECT 13.455 0.375 13.625 1.505 ;
        RECT 14.425 0.625 14.595 1.505 ;
        RECT 15.395 1.425 15.565 1.505 ;
        RECT 14.915 1.080 15.085 1.160 ;
        RECT 15.965 1.080 16.135 1.755 ;
        RECT 16.935 1.750 17.105 5.070 ;
        RECT 18.785 1.915 18.955 4.865 ;
        RECT 14.915 0.910 16.135 1.080 ;
        RECT 14.915 0.830 15.085 0.910 ;
        RECT 15.395 0.625 15.565 0.705 ;
        RECT 14.425 0.455 15.565 0.625 ;
        RECT 14.425 0.375 14.595 0.455 ;
        RECT 15.395 0.375 15.565 0.455 ;
        RECT 15.965 0.625 16.135 0.910 ;
        RECT 16.450 1.580 17.105 1.750 ;
        RECT 18.265 1.675 18.435 1.755 ;
        RECT 19.235 1.675 19.405 1.755 ;
        RECT 20.205 1.675 20.375 1.755 ;
        RECT 16.450 0.845 16.620 1.580 ;
        RECT 18.265 1.505 20.375 1.675 ;
        RECT 16.935 0.625 17.105 1.395 ;
        RECT 15.965 0.455 17.105 0.625 ;
        RECT 15.965 0.375 16.135 0.455 ;
        RECT 16.935 0.375 17.105 0.455 ;
        RECT 18.265 0.375 18.435 1.505 ;
        RECT 19.235 0.625 19.405 1.505 ;
        RECT 20.205 1.425 20.375 1.505 ;
        RECT 19.725 1.080 19.895 1.160 ;
        RECT 20.775 1.080 20.945 1.755 ;
        RECT 21.745 1.750 21.915 5.070 ;
        RECT 23.595 1.915 23.765 4.865 ;
        RECT 24.365 4.710 24.535 4.865 ;
        RECT 24.335 4.535 24.535 4.710 ;
        RECT 24.335 1.915 24.505 4.535 ;
        RECT 19.725 0.910 20.945 1.080 ;
        RECT 19.725 0.830 19.895 0.910 ;
        RECT 20.205 0.625 20.375 0.705 ;
        RECT 19.235 0.455 20.375 0.625 ;
        RECT 19.235 0.375 19.405 0.455 ;
        RECT 20.205 0.375 20.375 0.455 ;
        RECT 20.775 0.625 20.945 0.910 ;
        RECT 21.260 1.580 21.915 1.750 ;
        RECT 23.180 1.665 23.350 1.745 ;
        RECT 24.150 1.665 24.320 1.745 ;
        RECT 21.260 0.845 21.430 1.580 ;
        RECT 23.180 1.495 24.320 1.665 ;
        RECT 21.745 0.625 21.915 1.395 ;
        RECT 20.775 0.455 21.915 0.625 ;
        RECT 20.775 0.375 20.945 0.455 ;
        RECT 21.745 0.375 21.915 0.455 ;
        RECT 23.180 0.365 23.350 1.495 ;
        RECT 24.150 0.615 24.320 1.495 ;
        RECT 25.120 0.615 25.290 1.385 ;
        RECT 24.150 0.445 25.290 0.615 ;
        RECT 24.150 0.365 24.320 0.445 ;
        RECT 25.120 0.365 25.290 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 3.245 12.295 3.415 ;
        RECT 13.975 3.245 14.145 3.415 ;
        RECT 16.935 3.985 17.105 4.155 ;
        RECT 18.785 3.615 18.955 3.785 ;
        RECT 21.745 3.245 21.915 3.415 ;
        RECT 23.595 3.245 23.765 3.415 ;
        RECT 24.335 3.985 24.505 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 16.905 4.155 17.135 4.185 ;
        RECT 24.305 4.155 24.535 4.185 ;
        RECT 0.965 3.985 24.565 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 16.905 3.955 17.135 3.985 ;
        RECT 24.305 3.955 24.535 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 18.755 3.785 18.985 3.815 ;
        RECT 3.925 3.615 19.015 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 18.755 3.585 18.985 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 8.765 3.415 8.995 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.095 3.415 12.325 3.445 ;
        RECT 13.945 3.415 14.175 3.445 ;
        RECT 21.715 3.415 21.945 3.445 ;
        RECT 23.565 3.415 23.795 3.445 ;
        RECT 3.185 3.245 10.875 3.415 ;
        RECT 12.065 3.245 14.205 3.415 ;
        RECT 21.685 3.245 23.825 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 8.765 3.215 8.995 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.095 3.215 12.325 3.245 ;
        RECT 13.945 3.215 14.175 3.245 ;
        RECT 21.715 3.215 21.945 3.245 ;
        RECT 23.565 3.215 23.795 3.245 ;
  END
END DFFRNQX1






MACRO DFFRNX1
  CLASS CORE ;
  FOREIGN DFFRNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 25.900 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 23.715 5.285 23.885 7.020 ;
        RECT 24.595 5.285 24.765 7.020 ;
        RECT 23.715 5.115 25.245 5.285 ;
        RECT 21.005 1.915 21.175 4.865 ;
        RECT 25.075 1.740 25.245 5.115 ;
        RECT 24.635 1.570 25.245 1.740 ;
        RECT 24.635 0.835 24.805 1.570 ;
      LAYER mcon ;
        RECT 21.005 3.615 21.175 3.785 ;
        RECT 25.075 3.615 25.245 3.785 ;
      LAYER met1 ;
        RECT 20.975 3.785 21.205 3.815 ;
        RECT 25.045 3.785 25.275 3.815 ;
        RECT 20.945 3.615 25.305 3.785 ;
        RECT 20.975 3.585 21.205 3.615 ;
        RECT 25.045 3.585 25.275 3.615 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 19.205 5.240 19.375 7.020 ;
        RECT 20.085 5.240 20.255 7.020 ;
        RECT 20.965 5.240 21.135 7.020 ;
        RECT 19.205 5.070 21.915 5.240 ;
        RECT 21.745 1.750 21.915 5.070 ;
        RECT 23.595 1.915 23.765 4.865 ;
        RECT 21.260 1.580 21.915 1.750 ;
        RECT 21.260 0.845 21.430 1.580 ;
      LAYER mcon ;
        RECT 21.745 3.245 21.915 3.415 ;
        RECT 23.595 3.245 23.765 3.415 ;
      LAYER met1 ;
        RECT 21.715 3.415 21.945 3.445 ;
        RECT 23.565 3.415 23.795 3.445 ;
        RECT 21.685 3.245 23.825 3.415 ;
        RECT 21.715 3.215 21.945 3.245 ;
        RECT 23.565 3.215 23.795 3.245 ;
    END
  END QN
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 15.085 1.915 15.255 4.865 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 15.085 4.355 15.255 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 15.055 4.525 15.285 4.555 ;
        RECT 2.075 4.355 15.315 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 15.055 4.325 15.285 4.355 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 3.069350 ;
    PORT
      LAYER li1 ;
        RECT 8.055 1.915 8.225 4.865 ;
        RECT 16.195 1.915 16.365 4.865 ;
        RECT 19.895 1.915 20.065 4.865 ;
      LAYER mcon ;
        RECT 8.055 2.135 8.225 2.305 ;
        RECT 16.195 2.135 16.365 2.305 ;
        RECT 19.895 2.135 20.065 2.305 ;
      LAYER met1 ;
        RECT 8.025 2.305 8.255 2.335 ;
        RECT 16.165 2.305 16.395 2.335 ;
        RECT 19.865 2.305 20.095 2.335 ;
        RECT 7.995 2.135 20.125 2.305 ;
        RECT 8.025 2.105 8.255 2.135 ;
        RECT 16.165 2.105 16.395 2.135 ;
        RECT 19.865 2.105 20.095 2.135 ;
    END
  END RN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 26.335 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 26.070 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.325 5.135 10.495 7.230 ;
        RECT 11.205 5.555 11.375 7.230 ;
        RECT 12.085 5.555 12.255 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.955 5.215 14.125 7.230 ;
        RECT 14.835 5.555 15.005 7.230 ;
        RECT 15.715 5.555 15.885 7.230 ;
        RECT 16.595 5.555 16.765 7.230 ;
        RECT 17.590 4.110 17.930 7.230 ;
        RECT 18.765 5.215 18.935 7.230 ;
        RECT 19.645 5.555 19.815 7.230 ;
        RECT 20.525 5.555 20.695 7.230 ;
        RECT 21.405 5.555 21.575 7.230 ;
        RECT 22.400 4.110 22.740 7.230 ;
        RECT 23.275 5.135 23.445 7.230 ;
        RECT 24.155 5.555 24.325 7.230 ;
        RECT 25.035 5.555 25.205 7.230 ;
        RECT 25.730 4.110 26.070 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 26.070 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 26.070 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.715 0.170 10.885 1.120 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 13.940 0.170 14.110 1.130 ;
        RECT 17.590 0.170 17.930 2.720 ;
        RECT 18.750 0.170 18.920 1.130 ;
        RECT 22.400 0.170 22.740 2.720 ;
        RECT 23.665 0.170 23.835 1.120 ;
        RECT 25.730 0.170 26.070 2.720 ;
        RECT -0.170 -0.170 26.070 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 26.070 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 10.765 5.285 10.935 7.020 ;
        RECT 11.645 5.285 11.815 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 10.765 5.115 12.295 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 11.415 4.710 11.585 4.865 ;
        RECT 11.385 4.535 11.585 4.710 ;
        RECT 11.385 1.915 11.555 4.535 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.230 1.665 10.400 1.745 ;
        RECT 11.200 1.665 11.370 1.745 ;
        RECT 12.125 1.740 12.295 5.115 ;
        RECT 14.395 5.240 14.565 7.020 ;
        RECT 15.275 5.240 15.445 7.020 ;
        RECT 16.155 5.240 16.325 7.020 ;
        RECT 14.395 5.070 17.105 5.240 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.230 1.495 11.370 1.665 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.230 0.365 10.400 1.495 ;
        RECT 11.200 0.615 11.370 1.495 ;
        RECT 11.685 1.570 12.295 1.740 ;
        RECT 13.455 1.675 13.625 1.755 ;
        RECT 14.425 1.675 14.595 1.755 ;
        RECT 15.395 1.675 15.565 1.755 ;
        RECT 11.685 0.835 11.855 1.570 ;
        RECT 13.455 1.505 15.565 1.675 ;
        RECT 12.170 0.615 12.340 1.385 ;
        RECT 11.200 0.445 12.340 0.615 ;
        RECT 11.200 0.365 11.370 0.445 ;
        RECT 12.170 0.365 12.340 0.445 ;
        RECT 13.455 0.375 13.625 1.505 ;
        RECT 14.425 0.625 14.595 1.505 ;
        RECT 15.395 1.425 15.565 1.505 ;
        RECT 14.915 1.080 15.085 1.160 ;
        RECT 15.965 1.080 16.135 1.755 ;
        RECT 16.935 1.750 17.105 5.070 ;
        RECT 18.785 1.915 18.955 4.865 ;
        RECT 24.365 4.710 24.535 4.865 ;
        RECT 24.335 4.535 24.535 4.710 ;
        RECT 24.335 1.915 24.505 4.535 ;
        RECT 14.915 0.910 16.135 1.080 ;
        RECT 14.915 0.830 15.085 0.910 ;
        RECT 15.395 0.625 15.565 0.705 ;
        RECT 14.425 0.455 15.565 0.625 ;
        RECT 14.425 0.375 14.595 0.455 ;
        RECT 15.395 0.375 15.565 0.455 ;
        RECT 15.965 0.625 16.135 0.910 ;
        RECT 16.450 1.580 17.105 1.750 ;
        RECT 18.265 1.675 18.435 1.755 ;
        RECT 19.235 1.675 19.405 1.755 ;
        RECT 20.205 1.675 20.375 1.755 ;
        RECT 16.450 0.845 16.620 1.580 ;
        RECT 18.265 1.505 20.375 1.675 ;
        RECT 16.935 0.625 17.105 1.395 ;
        RECT 15.965 0.455 17.105 0.625 ;
        RECT 15.965 0.375 16.135 0.455 ;
        RECT 16.935 0.375 17.105 0.455 ;
        RECT 18.265 0.375 18.435 1.505 ;
        RECT 19.235 0.625 19.405 1.505 ;
        RECT 20.205 1.425 20.375 1.505 ;
        RECT 19.725 1.080 19.895 1.160 ;
        RECT 20.775 1.080 20.945 1.755 ;
        RECT 23.180 1.665 23.350 1.745 ;
        RECT 24.150 1.665 24.320 1.745 ;
        RECT 23.180 1.495 24.320 1.665 ;
        RECT 19.725 0.910 20.945 1.080 ;
        RECT 19.725 0.830 19.895 0.910 ;
        RECT 20.205 0.625 20.375 0.705 ;
        RECT 19.235 0.455 20.375 0.625 ;
        RECT 19.235 0.375 19.405 0.455 ;
        RECT 20.205 0.375 20.375 0.455 ;
        RECT 20.775 0.625 20.945 0.910 ;
        RECT 21.745 0.625 21.915 1.395 ;
        RECT 20.775 0.455 21.915 0.625 ;
        RECT 20.775 0.375 20.945 0.455 ;
        RECT 21.745 0.375 21.915 0.455 ;
        RECT 23.180 0.365 23.350 1.495 ;
        RECT 24.150 0.615 24.320 1.495 ;
        RECT 25.120 0.615 25.290 1.385 ;
        RECT 24.150 0.445 25.290 0.615 ;
        RECT 24.150 0.365 24.320 0.445 ;
        RECT 25.120 0.365 25.290 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 3.245 12.295 3.415 ;
        RECT 13.975 3.245 14.145 3.415 ;
        RECT 16.935 3.985 17.105 4.155 ;
        RECT 18.785 3.615 18.955 3.785 ;
        RECT 24.335 3.985 24.505 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 16.905 4.155 17.135 4.185 ;
        RECT 24.305 4.155 24.535 4.185 ;
        RECT 0.965 3.985 24.565 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 16.905 3.955 17.135 3.985 ;
        RECT 24.305 3.955 24.535 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 18.755 3.785 18.985 3.815 ;
        RECT 3.925 3.615 19.015 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 18.755 3.585 18.985 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 8.765 3.415 8.995 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.095 3.415 12.325 3.445 ;
        RECT 13.945 3.415 14.175 3.445 ;
        RECT 3.185 3.245 10.875 3.415 ;
        RECT 12.065 3.245 14.205 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 8.765 3.215 8.995 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.095 3.215 12.325 3.245 ;
        RECT 13.945 3.215 14.175 3.245 ;
  END
END DFFRNX1






MACRO DFFSNQNX1
  CLASS CORE ;
  FOREIGN DFFSNQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.420 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 17.425 5.285 17.595 7.020 ;
        RECT 18.305 5.285 18.475 7.020 ;
        RECT 17.425 5.115 18.955 5.285 ;
        RECT 18.785 1.740 18.955 5.115 ;
        RECT 20.635 1.915 20.805 4.865 ;
        RECT 18.345 1.570 18.955 1.740 ;
        RECT 18.345 0.835 18.515 1.570 ;
      LAYER mcon ;
        RECT 18.785 2.875 18.955 3.045 ;
        RECT 20.635 2.875 20.805 3.045 ;
      LAYER met1 ;
        RECT 18.755 3.045 18.985 3.075 ;
        RECT 20.605 3.045 20.835 3.075 ;
        RECT 18.725 2.875 20.865 3.045 ;
        RECT 18.755 2.845 18.985 2.875 ;
        RECT 20.605 2.845 20.835 2.875 ;
    END
  END QN
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 5.465 1.915 5.635 4.865 ;
        RECT 14.745 4.710 14.915 4.865 ;
        RECT 14.715 4.535 14.915 4.710 ;
        RECT 14.715 1.915 14.885 4.535 ;
      LAYER mcon ;
        RECT 5.465 4.355 5.635 4.525 ;
        RECT 14.715 4.355 14.885 4.525 ;
      LAYER met1 ;
        RECT 5.435 4.525 5.665 4.555 ;
        RECT 14.685 4.525 14.915 4.555 ;
        RECT 5.405 4.355 14.945 4.525 ;
        RECT 5.435 4.325 5.665 4.355 ;
        RECT 14.685 4.325 14.915 4.355 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 10.275 1.915 10.445 4.865 ;
        RECT 21.745 1.915 21.915 4.865 ;
      LAYER mcon ;
        RECT 10.275 2.135 10.445 2.305 ;
        RECT 21.745 2.135 21.915 2.305 ;
      LAYER met1 ;
        RECT 10.245 2.305 10.475 2.335 ;
        RECT 21.715 2.305 21.945 2.335 ;
        RECT 10.215 2.135 21.975 2.305 ;
        RECT 10.245 2.105 10.475 2.135 ;
        RECT 21.715 2.105 21.945 2.135 ;
    END
  END SN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 24.855 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 24.590 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.335 5.215 4.505 7.230 ;
        RECT 5.215 5.555 5.385 7.230 ;
        RECT 6.095 5.555 6.265 7.230 ;
        RECT 6.975 5.555 7.145 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 9.145 5.215 9.315 7.230 ;
        RECT 10.025 5.555 10.195 7.230 ;
        RECT 10.905 5.555 11.075 7.230 ;
        RECT 11.785 5.555 11.955 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.655 5.135 13.825 7.230 ;
        RECT 14.535 5.555 14.705 7.230 ;
        RECT 15.415 5.555 15.585 7.230 ;
        RECT 16.110 4.110 16.450 7.230 ;
        RECT 16.985 5.135 17.155 7.230 ;
        RECT 17.865 5.555 18.035 7.230 ;
        RECT 18.745 5.555 18.915 7.230 ;
        RECT 19.440 4.110 19.780 7.230 ;
        RECT 20.615 5.215 20.785 7.230 ;
        RECT 21.495 5.555 21.665 7.230 ;
        RECT 22.375 5.555 22.545 7.230 ;
        RECT 23.255 5.555 23.425 7.230 ;
        RECT 24.250 4.110 24.590 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 24.590 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 24.590 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 4.320 0.170 4.490 1.130 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.130 0.170 9.300 1.130 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 14.045 0.170 14.215 1.120 ;
        RECT 16.110 0.170 16.450 2.720 ;
        RECT 17.375 0.170 17.545 1.120 ;
        RECT 19.440 0.170 19.780 2.720 ;
        RECT 20.600 0.170 20.770 1.130 ;
        RECT 24.250 0.170 24.590 2.720 ;
        RECT -0.170 -0.170 24.590 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 24.590 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.775 5.240 4.945 7.020 ;
        RECT 5.655 5.240 5.825 7.020 ;
        RECT 6.535 5.240 6.705 7.020 ;
        RECT 9.585 5.240 9.755 7.020 ;
        RECT 10.465 5.240 10.635 7.020 ;
        RECT 11.345 5.240 11.515 7.020 ;
        RECT 14.095 5.285 14.265 7.020 ;
        RECT 14.975 5.285 15.145 7.020 ;
        RECT 4.775 5.070 7.485 5.240 ;
        RECT 9.585 5.070 12.295 5.240 ;
        RECT 14.095 5.115 15.625 5.285 ;
        RECT 4.355 1.915 4.525 4.865 ;
        RECT 6.575 1.915 6.745 4.865 ;
        RECT 7.315 4.235 7.485 5.070 ;
        RECT 7.310 3.905 7.485 4.235 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 3.835 1.675 4.005 1.755 ;
        RECT 4.805 1.675 4.975 1.755 ;
        RECT 5.775 1.675 5.945 1.755 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 3.835 1.505 5.945 1.675 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 3.835 0.375 4.005 1.505 ;
        RECT 4.805 0.625 4.975 1.505 ;
        RECT 5.775 1.425 5.945 1.505 ;
        RECT 5.295 1.080 5.465 1.160 ;
        RECT 6.345 1.080 6.515 1.755 ;
        RECT 7.315 1.750 7.485 3.905 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 11.385 1.915 11.555 4.865 ;
        RECT 5.295 0.910 6.515 1.080 ;
        RECT 5.295 0.830 5.465 0.910 ;
        RECT 5.775 0.625 5.945 0.705 ;
        RECT 4.805 0.455 5.945 0.625 ;
        RECT 4.805 0.375 4.975 0.455 ;
        RECT 5.775 0.375 5.945 0.455 ;
        RECT 6.345 0.625 6.515 0.910 ;
        RECT 6.830 1.580 7.485 1.750 ;
        RECT 8.645 1.675 8.815 1.755 ;
        RECT 9.615 1.675 9.785 1.755 ;
        RECT 10.585 1.675 10.755 1.755 ;
        RECT 6.830 0.845 7.000 1.580 ;
        RECT 8.645 1.505 10.755 1.675 ;
        RECT 7.315 0.625 7.485 1.395 ;
        RECT 6.345 0.455 7.485 0.625 ;
        RECT 6.345 0.375 6.515 0.455 ;
        RECT 7.315 0.375 7.485 0.455 ;
        RECT 8.645 0.375 8.815 1.505 ;
        RECT 9.615 0.625 9.785 1.505 ;
        RECT 10.585 1.425 10.755 1.505 ;
        RECT 10.105 1.080 10.275 1.160 ;
        RECT 11.155 1.080 11.325 1.755 ;
        RECT 12.125 1.750 12.295 5.070 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 10.105 0.910 11.325 1.080 ;
        RECT 10.105 0.830 10.275 0.910 ;
        RECT 10.585 0.625 10.755 0.705 ;
        RECT 9.615 0.455 10.755 0.625 ;
        RECT 9.615 0.375 9.785 0.455 ;
        RECT 10.585 0.375 10.755 0.455 ;
        RECT 11.155 0.625 11.325 0.910 ;
        RECT 11.640 1.580 12.295 1.750 ;
        RECT 13.560 1.665 13.730 1.745 ;
        RECT 14.530 1.665 14.700 1.745 ;
        RECT 15.455 1.740 15.625 5.115 ;
        RECT 21.055 5.240 21.225 7.020 ;
        RECT 21.935 5.240 22.105 7.020 ;
        RECT 22.815 5.240 22.985 7.020 ;
        RECT 21.055 5.070 23.765 5.240 ;
        RECT 17.305 1.915 17.475 4.865 ;
        RECT 18.075 4.710 18.245 4.865 ;
        RECT 18.045 4.535 18.245 4.710 ;
        RECT 18.045 1.915 18.215 4.535 ;
        RECT 22.855 1.915 23.025 4.865 ;
        RECT 11.640 0.845 11.810 1.580 ;
        RECT 13.560 1.495 14.700 1.665 ;
        RECT 12.125 0.625 12.295 1.395 ;
        RECT 11.155 0.455 12.295 0.625 ;
        RECT 11.155 0.375 11.325 0.455 ;
        RECT 12.125 0.375 12.295 0.455 ;
        RECT 13.560 0.365 13.730 1.495 ;
        RECT 14.530 0.615 14.700 1.495 ;
        RECT 15.015 1.570 15.625 1.740 ;
        RECT 16.890 1.665 17.060 1.745 ;
        RECT 17.860 1.665 18.030 1.745 ;
        RECT 15.015 0.835 15.185 1.570 ;
        RECT 16.890 1.495 18.030 1.665 ;
        RECT 15.500 0.615 15.670 1.385 ;
        RECT 14.530 0.445 15.670 0.615 ;
        RECT 14.530 0.365 14.700 0.445 ;
        RECT 15.500 0.365 15.670 0.445 ;
        RECT 16.890 0.365 17.060 1.495 ;
        RECT 17.860 0.615 18.030 1.495 ;
        RECT 20.115 1.675 20.285 1.755 ;
        RECT 21.085 1.675 21.255 1.755 ;
        RECT 22.055 1.675 22.225 1.755 ;
        RECT 20.115 1.505 22.225 1.675 ;
        RECT 18.830 0.615 19.000 1.385 ;
        RECT 17.860 0.445 19.000 0.615 ;
        RECT 17.860 0.365 18.030 0.445 ;
        RECT 18.830 0.365 19.000 0.445 ;
        RECT 20.115 0.375 20.285 1.505 ;
        RECT 21.085 0.625 21.255 1.505 ;
        RECT 22.055 1.425 22.225 1.505 ;
        RECT 21.575 1.080 21.745 1.160 ;
        RECT 22.625 1.080 22.795 1.755 ;
        RECT 23.595 1.750 23.765 5.070 ;
        RECT 21.575 0.910 22.795 1.080 ;
        RECT 21.575 0.830 21.745 0.910 ;
        RECT 22.055 0.625 22.225 0.705 ;
        RECT 21.085 0.455 22.225 0.625 ;
        RECT 21.085 0.375 21.255 0.455 ;
        RECT 22.055 0.375 22.225 0.455 ;
        RECT 22.625 0.625 22.795 0.910 ;
        RECT 23.110 1.580 23.765 1.750 ;
        RECT 23.110 0.845 23.280 1.580 ;
        RECT 23.595 0.625 23.765 1.395 ;
        RECT 22.625 0.455 23.765 0.625 ;
        RECT 22.625 0.375 22.795 0.455 ;
        RECT 23.595 0.375 23.765 0.455 ;
      LAYER mcon ;
        RECT 1.765 3.985 1.935 4.155 ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.500 4.525 2.670 ;
        RECT 7.310 3.985 7.480 4.155 ;
        RECT 6.575 3.615 6.745 3.785 ;
        RECT 9.165 2.505 9.335 2.675 ;
        RECT 11.385 3.615 11.555 3.785 ;
        RECT 12.125 2.505 12.295 2.675 ;
        RECT 13.975 2.505 14.145 2.675 ;
        RECT 15.455 3.615 15.625 3.785 ;
        RECT 17.305 3.985 17.475 4.155 ;
        RECT 18.045 3.245 18.215 3.415 ;
        RECT 22.855 3.615 23.025 3.785 ;
        RECT 23.595 3.245 23.765 3.415 ;
      LAYER met1 ;
        RECT 1.735 4.155 1.965 4.185 ;
        RECT 7.280 4.155 7.510 4.185 ;
        RECT 17.275 4.155 17.505 4.185 ;
        RECT 1.705 3.985 17.535 4.155 ;
        RECT 1.735 3.955 1.965 3.985 ;
        RECT 7.280 3.955 7.510 3.985 ;
        RECT 17.275 3.955 17.505 3.985 ;
        RECT 6.545 3.785 6.775 3.815 ;
        RECT 11.355 3.785 11.585 3.815 ;
        RECT 15.425 3.785 15.655 3.815 ;
        RECT 22.825 3.785 23.055 3.815 ;
        RECT 6.515 3.615 23.085 3.785 ;
        RECT 6.545 3.585 6.775 3.615 ;
        RECT 11.355 3.585 11.585 3.615 ;
        RECT 15.425 3.585 15.655 3.615 ;
        RECT 22.825 3.585 23.055 3.615 ;
        RECT 18.015 3.415 18.245 3.445 ;
        RECT 23.565 3.415 23.795 3.445 ;
        RECT 17.985 3.245 23.825 3.415 ;
        RECT 18.015 3.215 18.245 3.245 ;
        RECT 23.565 3.215 23.795 3.245 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.700 ;
        RECT 9.135 2.675 9.365 2.705 ;
        RECT 12.095 2.675 12.325 2.705 ;
        RECT 13.945 2.675 14.175 2.705 ;
        RECT 2.445 2.505 9.395 2.675 ;
        RECT 12.065 2.505 14.205 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.295 2.500 4.705 2.505 ;
        RECT 4.325 2.470 4.555 2.500 ;
        RECT 9.135 2.475 9.365 2.505 ;
        RECT 12.095 2.475 12.325 2.505 ;
        RECT 13.945 2.475 14.175 2.505 ;
  END
END DFFSNQNX1






MACRO DFFSNQX1
  CLASS CORE ;
  FOREIGN DFFSNQX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.420 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 21.055 5.240 21.225 7.020 ;
        RECT 21.935 5.240 22.105 7.020 ;
        RECT 22.815 5.240 22.985 7.020 ;
        RECT 21.055 5.070 23.765 5.240 ;
        RECT 18.075 4.710 18.245 4.865 ;
        RECT 18.045 4.535 18.245 4.710 ;
        RECT 18.045 1.915 18.215 4.535 ;
        RECT 23.595 1.750 23.765 5.070 ;
        RECT 23.110 1.580 23.765 1.750 ;
        RECT 23.110 0.845 23.280 1.580 ;
      LAYER mcon ;
        RECT 18.045 3.245 18.215 3.415 ;
        RECT 23.595 3.245 23.765 3.415 ;
      LAYER met1 ;
        RECT 18.015 3.415 18.245 3.445 ;
        RECT 23.565 3.415 23.795 3.445 ;
        RECT 17.985 3.245 23.825 3.415 ;
        RECT 18.015 3.215 18.245 3.245 ;
        RECT 23.565 3.215 23.795 3.245 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 5.465 1.915 5.635 4.865 ;
        RECT 14.745 4.710 14.915 4.865 ;
        RECT 14.715 4.535 14.915 4.710 ;
        RECT 14.715 1.915 14.885 4.535 ;
      LAYER mcon ;
        RECT 5.465 4.355 5.635 4.525 ;
        RECT 14.715 4.355 14.885 4.525 ;
      LAYER met1 ;
        RECT 5.435 4.525 5.665 4.555 ;
        RECT 14.685 4.525 14.915 4.555 ;
        RECT 5.405 4.355 14.945 4.525 ;
        RECT 5.435 4.325 5.665 4.355 ;
        RECT 14.685 4.325 14.915 4.355 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 10.275 1.915 10.445 4.865 ;
        RECT 21.745 1.915 21.915 4.865 ;
      LAYER mcon ;
        RECT 10.275 2.135 10.445 2.305 ;
        RECT 21.745 2.135 21.915 2.305 ;
      LAYER met1 ;
        RECT 10.245 2.305 10.475 2.335 ;
        RECT 21.715 2.305 21.945 2.335 ;
        RECT 10.215 2.135 21.975 2.305 ;
        RECT 10.245 2.105 10.475 2.135 ;
        RECT 21.715 2.105 21.945 2.135 ;
    END
  END SN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 24.855 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 24.590 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.335 5.215 4.505 7.230 ;
        RECT 5.215 5.555 5.385 7.230 ;
        RECT 6.095 5.555 6.265 7.230 ;
        RECT 6.975 5.555 7.145 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 9.145 5.215 9.315 7.230 ;
        RECT 10.025 5.555 10.195 7.230 ;
        RECT 10.905 5.555 11.075 7.230 ;
        RECT 11.785 5.555 11.955 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.655 5.135 13.825 7.230 ;
        RECT 14.535 5.555 14.705 7.230 ;
        RECT 15.415 5.555 15.585 7.230 ;
        RECT 16.110 4.110 16.450 7.230 ;
        RECT 16.985 5.135 17.155 7.230 ;
        RECT 17.865 5.555 18.035 7.230 ;
        RECT 18.745 5.555 18.915 7.230 ;
        RECT 19.440 4.110 19.780 7.230 ;
        RECT 20.615 5.215 20.785 7.230 ;
        RECT 21.495 5.555 21.665 7.230 ;
        RECT 22.375 5.555 22.545 7.230 ;
        RECT 23.255 5.555 23.425 7.230 ;
        RECT 24.250 4.110 24.590 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 24.590 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 24.590 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 4.320 0.170 4.490 1.130 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.130 0.170 9.300 1.130 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 14.045 0.170 14.215 1.120 ;
        RECT 16.110 0.170 16.450 2.720 ;
        RECT 17.375 0.170 17.545 1.120 ;
        RECT 19.440 0.170 19.780 2.720 ;
        RECT 20.600 0.170 20.770 1.130 ;
        RECT 24.250 0.170 24.590 2.720 ;
        RECT -0.170 -0.170 24.590 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 24.590 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.775 5.240 4.945 7.020 ;
        RECT 5.655 5.240 5.825 7.020 ;
        RECT 6.535 5.240 6.705 7.020 ;
        RECT 9.585 5.240 9.755 7.020 ;
        RECT 10.465 5.240 10.635 7.020 ;
        RECT 11.345 5.240 11.515 7.020 ;
        RECT 14.095 5.285 14.265 7.020 ;
        RECT 14.975 5.285 15.145 7.020 ;
        RECT 17.425 5.285 17.595 7.020 ;
        RECT 18.305 5.285 18.475 7.020 ;
        RECT 4.775 5.070 7.485 5.240 ;
        RECT 9.585 5.070 12.295 5.240 ;
        RECT 14.095 5.115 15.625 5.285 ;
        RECT 17.425 5.115 18.955 5.285 ;
        RECT 4.355 1.915 4.525 4.865 ;
        RECT 6.575 1.915 6.745 4.865 ;
        RECT 7.315 4.235 7.485 5.070 ;
        RECT 7.310 3.905 7.485 4.235 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 3.835 1.675 4.005 1.755 ;
        RECT 4.805 1.675 4.975 1.755 ;
        RECT 5.775 1.675 5.945 1.755 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 3.835 1.505 5.945 1.675 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 3.835 0.375 4.005 1.505 ;
        RECT 4.805 0.625 4.975 1.505 ;
        RECT 5.775 1.425 5.945 1.505 ;
        RECT 5.295 1.080 5.465 1.160 ;
        RECT 6.345 1.080 6.515 1.755 ;
        RECT 7.315 1.750 7.485 3.905 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 11.385 1.915 11.555 4.865 ;
        RECT 5.295 0.910 6.515 1.080 ;
        RECT 5.295 0.830 5.465 0.910 ;
        RECT 5.775 0.625 5.945 0.705 ;
        RECT 4.805 0.455 5.945 0.625 ;
        RECT 4.805 0.375 4.975 0.455 ;
        RECT 5.775 0.375 5.945 0.455 ;
        RECT 6.345 0.625 6.515 0.910 ;
        RECT 6.830 1.580 7.485 1.750 ;
        RECT 8.645 1.675 8.815 1.755 ;
        RECT 9.615 1.675 9.785 1.755 ;
        RECT 10.585 1.675 10.755 1.755 ;
        RECT 6.830 0.845 7.000 1.580 ;
        RECT 8.645 1.505 10.755 1.675 ;
        RECT 7.315 0.625 7.485 1.395 ;
        RECT 6.345 0.455 7.485 0.625 ;
        RECT 6.345 0.375 6.515 0.455 ;
        RECT 7.315 0.375 7.485 0.455 ;
        RECT 8.645 0.375 8.815 1.505 ;
        RECT 9.615 0.625 9.785 1.505 ;
        RECT 10.585 1.425 10.755 1.505 ;
        RECT 10.105 1.080 10.275 1.160 ;
        RECT 11.155 1.080 11.325 1.755 ;
        RECT 12.125 1.750 12.295 5.070 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 10.105 0.910 11.325 1.080 ;
        RECT 10.105 0.830 10.275 0.910 ;
        RECT 10.585 0.625 10.755 0.705 ;
        RECT 9.615 0.455 10.755 0.625 ;
        RECT 9.615 0.375 9.785 0.455 ;
        RECT 10.585 0.375 10.755 0.455 ;
        RECT 11.155 0.625 11.325 0.910 ;
        RECT 11.640 1.580 12.295 1.750 ;
        RECT 13.560 1.665 13.730 1.745 ;
        RECT 14.530 1.665 14.700 1.745 ;
        RECT 15.455 1.740 15.625 5.115 ;
        RECT 17.305 1.915 17.475 4.865 ;
        RECT 11.640 0.845 11.810 1.580 ;
        RECT 13.560 1.495 14.700 1.665 ;
        RECT 12.125 0.625 12.295 1.395 ;
        RECT 11.155 0.455 12.295 0.625 ;
        RECT 11.155 0.375 11.325 0.455 ;
        RECT 12.125 0.375 12.295 0.455 ;
        RECT 13.560 0.365 13.730 1.495 ;
        RECT 14.530 0.615 14.700 1.495 ;
        RECT 15.015 1.570 15.625 1.740 ;
        RECT 16.890 1.665 17.060 1.745 ;
        RECT 17.860 1.665 18.030 1.745 ;
        RECT 18.785 1.740 18.955 5.115 ;
        RECT 20.635 1.915 20.805 4.865 ;
        RECT 22.855 1.915 23.025 4.865 ;
        RECT 15.015 0.835 15.185 1.570 ;
        RECT 16.890 1.495 18.030 1.665 ;
        RECT 15.500 0.615 15.670 1.385 ;
        RECT 14.530 0.445 15.670 0.615 ;
        RECT 14.530 0.365 14.700 0.445 ;
        RECT 15.500 0.365 15.670 0.445 ;
        RECT 16.890 0.365 17.060 1.495 ;
        RECT 17.860 0.615 18.030 1.495 ;
        RECT 18.345 1.570 18.955 1.740 ;
        RECT 20.115 1.675 20.285 1.755 ;
        RECT 21.085 1.675 21.255 1.755 ;
        RECT 22.055 1.675 22.225 1.755 ;
        RECT 18.345 0.835 18.515 1.570 ;
        RECT 20.115 1.505 22.225 1.675 ;
        RECT 18.830 0.615 19.000 1.385 ;
        RECT 17.860 0.445 19.000 0.615 ;
        RECT 17.860 0.365 18.030 0.445 ;
        RECT 18.830 0.365 19.000 0.445 ;
        RECT 20.115 0.375 20.285 1.505 ;
        RECT 21.085 0.625 21.255 1.505 ;
        RECT 22.055 1.425 22.225 1.505 ;
        RECT 21.575 1.080 21.745 1.160 ;
        RECT 22.625 1.080 22.795 1.755 ;
        RECT 21.575 0.910 22.795 1.080 ;
        RECT 21.575 0.830 21.745 0.910 ;
        RECT 22.055 0.625 22.225 0.705 ;
        RECT 21.085 0.455 22.225 0.625 ;
        RECT 21.085 0.375 21.255 0.455 ;
        RECT 22.055 0.375 22.225 0.455 ;
        RECT 22.625 0.625 22.795 0.910 ;
        RECT 23.595 0.625 23.765 1.395 ;
        RECT 22.625 0.455 23.765 0.625 ;
        RECT 22.625 0.375 22.795 0.455 ;
        RECT 23.595 0.375 23.765 0.455 ;
      LAYER mcon ;
        RECT 1.765 3.985 1.935 4.155 ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.500 4.525 2.670 ;
        RECT 7.310 3.985 7.480 4.155 ;
        RECT 6.575 3.615 6.745 3.785 ;
        RECT 9.165 2.505 9.335 2.675 ;
        RECT 11.385 3.615 11.555 3.785 ;
        RECT 12.125 2.505 12.295 2.675 ;
        RECT 13.975 2.505 14.145 2.675 ;
        RECT 15.455 3.615 15.625 3.785 ;
        RECT 17.305 3.985 17.475 4.155 ;
        RECT 18.785 2.875 18.955 3.045 ;
        RECT 20.635 2.875 20.805 3.045 ;
        RECT 22.855 3.615 23.025 3.785 ;
      LAYER met1 ;
        RECT 1.735 4.155 1.965 4.185 ;
        RECT 7.280 4.155 7.510 4.185 ;
        RECT 17.275 4.155 17.505 4.185 ;
        RECT 1.705 3.985 17.535 4.155 ;
        RECT 1.735 3.955 1.965 3.985 ;
        RECT 7.280 3.955 7.510 3.985 ;
        RECT 17.275 3.955 17.505 3.985 ;
        RECT 6.545 3.785 6.775 3.815 ;
        RECT 11.355 3.785 11.585 3.815 ;
        RECT 15.425 3.785 15.655 3.815 ;
        RECT 22.825 3.785 23.055 3.815 ;
        RECT 6.515 3.615 23.085 3.785 ;
        RECT 6.545 3.585 6.775 3.615 ;
        RECT 11.355 3.585 11.585 3.615 ;
        RECT 15.425 3.585 15.655 3.615 ;
        RECT 22.825 3.585 23.055 3.615 ;
        RECT 18.755 3.045 18.985 3.075 ;
        RECT 20.605 3.045 20.835 3.075 ;
        RECT 18.725 2.875 20.865 3.045 ;
        RECT 18.755 2.845 18.985 2.875 ;
        RECT 20.605 2.845 20.835 2.875 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.700 ;
        RECT 9.135 2.675 9.365 2.705 ;
        RECT 12.095 2.675 12.325 2.705 ;
        RECT 13.945 2.675 14.175 2.705 ;
        RECT 2.445 2.505 9.395 2.675 ;
        RECT 12.065 2.505 14.205 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.295 2.500 4.705 2.505 ;
        RECT 4.325 2.470 4.555 2.500 ;
        RECT 9.135 2.475 9.365 2.505 ;
        RECT 12.095 2.475 12.325 2.505 ;
        RECT 13.945 2.475 14.175 2.505 ;
  END
END DFFSNQX1






MACRO DFFSNRNQNX1
  CLASS CORE ;
  FOREIGN DFFSNRNQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.860 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 20.685 5.240 20.855 7.020 ;
        RECT 21.565 5.240 21.735 7.020 ;
        RECT 22.445 5.240 22.615 7.020 ;
        RECT 20.685 5.070 23.395 5.240 ;
        RECT 23.225 1.750 23.395 5.070 ;
        RECT 25.075 1.915 25.245 4.865 ;
        RECT 22.740 1.580 23.395 1.750 ;
        RECT 22.740 0.845 22.910 1.580 ;
      LAYER mcon ;
        RECT 23.225 3.245 23.395 3.415 ;
        RECT 25.075 3.245 25.245 3.415 ;
      LAYER met1 ;
        RECT 23.195 3.415 23.425 3.445 ;
        RECT 25.045 3.415 25.275 3.445 ;
        RECT 23.165 3.245 25.305 3.415 ;
        RECT 23.195 3.215 23.425 3.245 ;
        RECT 25.045 3.215 25.275 3.245 ;
    END
  END QN
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 16.565 1.915 16.735 4.865 ;
      LAYER mcon ;
        RECT 6.945 3.245 7.115 3.415 ;
        RECT 16.565 3.245 16.735 3.415 ;
      LAYER met1 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 16.535 3.415 16.765 3.445 ;
        RECT 6.885 3.245 16.795 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
        RECT 16.535 3.215 16.765 3.245 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 3.056950 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 17.675 1.915 17.845 4.865 ;
        RECT 21.375 1.915 21.545 4.865 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 17.675 4.355 17.845 4.525 ;
        RECT 21.375 4.355 21.545 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 17.645 4.525 17.875 4.555 ;
        RECT 21.345 4.525 21.575 4.555 ;
        RECT 2.075 4.355 21.605 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 17.645 4.325 17.875 4.355 ;
        RECT 21.345 4.325 21.575 4.355 ;
    END
  END RN
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 11.755 1.915 11.925 4.865 ;
        RECT 26.185 1.915 26.355 4.865 ;
      LAYER mcon ;
        RECT 11.755 2.510 11.925 2.680 ;
        RECT 26.185 2.505 26.355 2.675 ;
      LAYER met1 ;
        RECT 11.725 2.680 11.955 2.710 ;
        RECT 11.695 2.675 12.105 2.680 ;
        RECT 26.155 2.675 26.385 2.705 ;
        RECT 11.695 2.510 26.415 2.675 ;
        RECT 11.725 2.480 11.955 2.510 ;
        RECT 12.105 2.505 26.415 2.510 ;
        RECT 26.155 2.475 26.385 2.505 ;
    END
  END SN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 29.295 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 29.030 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.625 5.215 10.795 7.230 ;
        RECT 11.505 5.555 11.675 7.230 ;
        RECT 12.385 5.555 12.555 7.230 ;
        RECT 13.265 5.555 13.435 7.230 ;
        RECT 14.260 4.110 14.600 7.230 ;
        RECT 15.435 5.215 15.605 7.230 ;
        RECT 16.315 5.555 16.485 7.230 ;
        RECT 17.195 5.555 17.365 7.230 ;
        RECT 18.075 5.555 18.245 7.230 ;
        RECT 19.070 4.110 19.410 7.230 ;
        RECT 20.245 5.215 20.415 7.230 ;
        RECT 21.125 5.555 21.295 7.230 ;
        RECT 22.005 5.555 22.175 7.230 ;
        RECT 22.885 5.555 23.055 7.230 ;
        RECT 23.880 4.110 24.220 7.230 ;
        RECT 25.055 5.215 25.225 7.230 ;
        RECT 25.935 5.555 26.105 7.230 ;
        RECT 26.815 5.555 26.985 7.230 ;
        RECT 27.695 5.555 27.865 7.230 ;
        RECT 28.690 4.110 29.030 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 29.030 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 29.030 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.610 0.170 10.780 1.130 ;
        RECT 14.260 0.170 14.600 2.720 ;
        RECT 15.420 0.170 15.590 1.130 ;
        RECT 19.070 0.170 19.410 2.720 ;
        RECT 20.230 0.170 20.400 1.130 ;
        RECT 23.880 0.170 24.220 2.720 ;
        RECT 25.040 0.170 25.210 1.130 ;
        RECT 28.690 0.170 29.030 2.720 ;
        RECT -0.170 -0.170 29.030 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 29.030 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 11.065 5.240 11.235 7.020 ;
        RECT 11.945 5.240 12.115 7.020 ;
        RECT 12.825 5.240 12.995 7.020 ;
        RECT 15.875 5.240 16.045 7.020 ;
        RECT 16.755 5.240 16.925 7.020 ;
        RECT 17.635 5.240 17.805 7.020 ;
        RECT 25.495 5.240 25.665 7.020 ;
        RECT 26.375 5.240 26.545 7.020 ;
        RECT 27.255 5.240 27.425 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 11.065 5.070 13.775 5.240 ;
        RECT 15.875 5.070 18.585 5.240 ;
        RECT 25.495 5.070 28.205 5.240 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 8.055 4.235 8.225 4.865 ;
        RECT 8.050 3.905 8.225 4.235 ;
        RECT 8.055 1.915 8.225 3.905 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 12.865 1.915 13.035 4.865 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.125 1.675 10.295 1.755 ;
        RECT 11.095 1.675 11.265 1.755 ;
        RECT 12.065 1.675 12.235 1.755 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.125 1.505 12.235 1.675 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.125 0.375 10.295 1.505 ;
        RECT 11.095 0.625 11.265 1.505 ;
        RECT 12.065 1.425 12.235 1.505 ;
        RECT 11.585 1.080 11.755 1.160 ;
        RECT 12.635 1.080 12.805 1.755 ;
        RECT 13.605 1.750 13.775 5.070 ;
        RECT 15.455 1.915 15.625 4.865 ;
        RECT 11.585 0.910 12.805 1.080 ;
        RECT 11.585 0.830 11.755 0.910 ;
        RECT 12.065 0.625 12.235 0.705 ;
        RECT 11.095 0.455 12.235 0.625 ;
        RECT 11.095 0.375 11.265 0.455 ;
        RECT 12.065 0.375 12.235 0.455 ;
        RECT 12.635 0.625 12.805 0.910 ;
        RECT 13.120 1.580 13.775 1.750 ;
        RECT 14.935 1.675 15.105 1.755 ;
        RECT 15.905 1.675 16.075 1.755 ;
        RECT 16.875 1.675 17.045 1.755 ;
        RECT 13.120 0.845 13.290 1.580 ;
        RECT 14.935 1.505 17.045 1.675 ;
        RECT 13.605 0.625 13.775 1.395 ;
        RECT 12.635 0.455 13.775 0.625 ;
        RECT 12.635 0.375 12.805 0.455 ;
        RECT 13.605 0.375 13.775 0.455 ;
        RECT 14.935 0.375 15.105 1.505 ;
        RECT 15.905 0.625 16.075 1.505 ;
        RECT 16.875 1.425 17.045 1.505 ;
        RECT 16.395 1.080 16.565 1.160 ;
        RECT 17.445 1.080 17.615 1.755 ;
        RECT 18.415 1.750 18.585 5.070 ;
        RECT 20.265 1.915 20.435 4.865 ;
        RECT 22.485 1.915 22.655 4.865 ;
        RECT 27.295 1.915 27.465 4.865 ;
        RECT 16.395 0.910 17.615 1.080 ;
        RECT 16.395 0.830 16.565 0.910 ;
        RECT 16.875 0.625 17.045 0.705 ;
        RECT 15.905 0.455 17.045 0.625 ;
        RECT 15.905 0.375 16.075 0.455 ;
        RECT 16.875 0.375 17.045 0.455 ;
        RECT 17.445 0.625 17.615 0.910 ;
        RECT 17.930 1.580 18.585 1.750 ;
        RECT 19.745 1.675 19.915 1.755 ;
        RECT 20.715 1.675 20.885 1.755 ;
        RECT 21.685 1.675 21.855 1.755 ;
        RECT 17.930 0.845 18.100 1.580 ;
        RECT 19.745 1.505 21.855 1.675 ;
        RECT 18.415 0.625 18.585 1.395 ;
        RECT 17.445 0.455 18.585 0.625 ;
        RECT 17.445 0.375 17.615 0.455 ;
        RECT 18.415 0.375 18.585 0.455 ;
        RECT 19.745 0.375 19.915 1.505 ;
        RECT 20.715 0.625 20.885 1.505 ;
        RECT 21.685 1.425 21.855 1.505 ;
        RECT 21.205 1.080 21.375 1.160 ;
        RECT 22.255 1.080 22.425 1.755 ;
        RECT 24.555 1.675 24.725 1.755 ;
        RECT 25.525 1.675 25.695 1.755 ;
        RECT 26.495 1.675 26.665 1.755 ;
        RECT 24.555 1.505 26.665 1.675 ;
        RECT 21.205 0.910 22.425 1.080 ;
        RECT 21.205 0.830 21.375 0.910 ;
        RECT 21.685 0.625 21.855 0.705 ;
        RECT 20.715 0.455 21.855 0.625 ;
        RECT 20.715 0.375 20.885 0.455 ;
        RECT 21.685 0.375 21.855 0.455 ;
        RECT 22.255 0.625 22.425 0.910 ;
        RECT 23.225 0.625 23.395 1.395 ;
        RECT 22.255 0.455 23.395 0.625 ;
        RECT 22.255 0.375 22.425 0.455 ;
        RECT 23.225 0.375 23.395 0.455 ;
        RECT 24.555 0.375 24.725 1.505 ;
        RECT 25.525 0.625 25.695 1.505 ;
        RECT 26.495 1.425 26.665 1.505 ;
        RECT 26.015 1.080 26.185 1.160 ;
        RECT 27.065 1.080 27.235 1.755 ;
        RECT 28.035 1.750 28.205 5.070 ;
        RECT 26.015 0.910 27.235 1.080 ;
        RECT 26.015 0.830 26.185 0.910 ;
        RECT 26.495 0.625 26.665 0.705 ;
        RECT 25.525 0.455 26.665 0.625 ;
        RECT 25.525 0.375 25.695 0.455 ;
        RECT 26.495 0.375 26.665 0.455 ;
        RECT 27.065 0.625 27.235 0.910 ;
        RECT 27.550 1.580 28.205 1.750 ;
        RECT 27.550 0.845 27.720 1.580 ;
        RECT 28.035 0.625 28.205 1.395 ;
        RECT 27.065 0.455 28.205 0.625 ;
        RECT 27.065 0.375 27.235 0.455 ;
        RECT 28.035 0.375 28.205 0.455 ;
      LAYER mcon ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 2.880 4.155 3.050 ;
        RECT 8.050 3.985 8.220 4.155 ;
        RECT 5.835 2.880 6.005 3.050 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 2.880 10.815 3.050 ;
        RECT 12.865 3.985 13.035 4.155 ;
        RECT 13.605 2.875 13.775 3.045 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 20.265 3.615 20.435 3.785 ;
        RECT 22.485 3.615 22.655 3.785 ;
        RECT 27.295 3.985 27.465 4.155 ;
        RECT 28.035 3.615 28.205 3.785 ;
      LAYER met1 ;
        RECT 8.020 4.155 8.250 4.185 ;
        RECT 12.835 4.155 13.065 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 7.990 3.985 27.525 4.155 ;
        RECT 8.020 3.955 8.250 3.985 ;
        RECT 12.835 3.955 13.065 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 20.235 3.785 20.465 3.815 ;
        RECT 22.455 3.785 22.685 3.815 ;
        RECT 28.005 3.785 28.235 3.815 ;
        RECT 3.185 3.615 20.495 3.785 ;
        RECT 22.425 3.615 28.265 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 20.235 3.585 20.465 3.615 ;
        RECT 22.455 3.585 22.685 3.615 ;
        RECT 28.005 3.585 28.235 3.615 ;
        RECT 3.955 3.050 4.185 3.080 ;
        RECT 5.805 3.050 6.035 3.080 ;
        RECT 10.615 3.050 10.845 3.080 ;
        RECT 3.925 2.880 10.875 3.050 ;
        RECT 13.575 3.045 13.805 3.075 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 3.955 2.850 4.185 2.880 ;
        RECT 5.805 2.850 6.035 2.880 ;
        RECT 10.615 2.850 10.845 2.880 ;
        RECT 13.545 2.875 15.685 3.045 ;
        RECT 13.575 2.845 13.805 2.875 ;
        RECT 15.425 2.845 15.655 2.875 ;
  END
END DFFSNRNQNX1






MACRO DFFSNRNQX1
  CLASS CORE ;
  FOREIGN DFFSNRNQX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.860 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 25.495 5.240 25.665 7.020 ;
        RECT 26.375 5.240 26.545 7.020 ;
        RECT 27.255 5.240 27.425 7.020 ;
        RECT 25.495 5.070 28.205 5.240 ;
        RECT 22.485 1.915 22.655 4.865 ;
        RECT 28.035 1.750 28.205 5.070 ;
        RECT 27.550 1.580 28.205 1.750 ;
        RECT 27.550 0.845 27.720 1.580 ;
      LAYER mcon ;
        RECT 22.485 3.615 22.655 3.785 ;
        RECT 28.035 3.615 28.205 3.785 ;
      LAYER met1 ;
        RECT 22.455 3.785 22.685 3.815 ;
        RECT 28.005 3.785 28.235 3.815 ;
        RECT 22.425 3.615 28.265 3.785 ;
        RECT 22.455 3.585 22.685 3.615 ;
        RECT 28.005 3.585 28.235 3.615 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 16.565 1.915 16.735 4.865 ;
      LAYER mcon ;
        RECT 6.945 3.245 7.115 3.415 ;
        RECT 16.565 3.245 16.735 3.415 ;
      LAYER met1 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 16.535 3.415 16.765 3.445 ;
        RECT 6.885 3.245 16.795 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
        RECT 16.535 3.215 16.765 3.245 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 11.755 1.915 11.925 4.865 ;
        RECT 26.185 1.915 26.355 4.865 ;
      LAYER mcon ;
        RECT 11.755 2.505 11.925 2.675 ;
        RECT 26.185 2.505 26.355 2.675 ;
      LAYER met1 ;
        RECT 11.725 2.675 11.955 2.705 ;
        RECT 26.155 2.675 26.385 2.705 ;
        RECT 11.695 2.505 26.415 2.675 ;
        RECT 11.725 2.475 11.955 2.505 ;
        RECT 26.155 2.475 26.385 2.505 ;
    END
  END SN
  PIN RN
    ANTENNAGATEAREA 3.056950 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 17.675 1.915 17.845 4.865 ;
        RECT 21.375 1.915 21.545 4.865 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 17.675 4.355 17.845 4.525 ;
        RECT 21.375 4.355 21.545 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 17.645 4.525 17.875 4.555 ;
        RECT 21.345 4.525 21.575 4.555 ;
        RECT 2.075 4.355 21.605 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 17.645 4.325 17.875 4.355 ;
        RECT 21.345 4.325 21.575 4.355 ;
    END
  END RN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 29.295 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 29.030 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.625 5.215 10.795 7.230 ;
        RECT 11.505 5.555 11.675 7.230 ;
        RECT 12.385 5.555 12.555 7.230 ;
        RECT 13.265 5.555 13.435 7.230 ;
        RECT 14.260 4.110 14.600 7.230 ;
        RECT 15.435 5.215 15.605 7.230 ;
        RECT 16.315 5.555 16.485 7.230 ;
        RECT 17.195 5.555 17.365 7.230 ;
        RECT 18.075 5.555 18.245 7.230 ;
        RECT 19.070 4.110 19.410 7.230 ;
        RECT 20.245 5.215 20.415 7.230 ;
        RECT 21.125 5.555 21.295 7.230 ;
        RECT 22.005 5.555 22.175 7.230 ;
        RECT 22.885 5.555 23.055 7.230 ;
        RECT 23.880 4.110 24.220 7.230 ;
        RECT 25.055 5.215 25.225 7.230 ;
        RECT 25.935 5.555 26.105 7.230 ;
        RECT 26.815 5.555 26.985 7.230 ;
        RECT 27.695 5.555 27.865 7.230 ;
        RECT 28.690 4.110 29.030 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 29.030 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 29.030 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.610 0.170 10.780 1.130 ;
        RECT 14.260 0.170 14.600 2.720 ;
        RECT 15.420 0.170 15.590 1.130 ;
        RECT 19.070 0.170 19.410 2.720 ;
        RECT 20.230 0.170 20.400 1.130 ;
        RECT 23.880 0.170 24.220 2.720 ;
        RECT 25.040 0.170 25.210 1.130 ;
        RECT 28.690 0.170 29.030 2.720 ;
        RECT -0.170 -0.170 29.030 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 29.030 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 11.065 5.240 11.235 7.020 ;
        RECT 11.945 5.240 12.115 7.020 ;
        RECT 12.825 5.240 12.995 7.020 ;
        RECT 15.875 5.240 16.045 7.020 ;
        RECT 16.755 5.240 16.925 7.020 ;
        RECT 17.635 5.240 17.805 7.020 ;
        RECT 20.685 5.240 20.855 7.020 ;
        RECT 21.565 5.240 21.735 7.020 ;
        RECT 22.445 5.240 22.615 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 11.065 5.070 13.775 5.240 ;
        RECT 15.875 5.070 18.585 5.240 ;
        RECT 20.685 5.070 23.395 5.240 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 8.055 4.235 8.225 4.865 ;
        RECT 8.050 3.905 8.225 4.235 ;
        RECT 8.055 1.915 8.225 3.905 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 12.865 1.915 13.035 4.865 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.125 1.675 10.295 1.755 ;
        RECT 11.095 1.675 11.265 1.755 ;
        RECT 12.065 1.675 12.235 1.755 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.125 1.505 12.235 1.675 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.125 0.375 10.295 1.505 ;
        RECT 11.095 0.625 11.265 1.505 ;
        RECT 12.065 1.425 12.235 1.505 ;
        RECT 11.585 1.080 11.755 1.160 ;
        RECT 12.635 1.080 12.805 1.755 ;
        RECT 13.605 1.750 13.775 5.070 ;
        RECT 15.455 1.915 15.625 4.865 ;
        RECT 11.585 0.910 12.805 1.080 ;
        RECT 11.585 0.830 11.755 0.910 ;
        RECT 12.065 0.625 12.235 0.705 ;
        RECT 11.095 0.455 12.235 0.625 ;
        RECT 11.095 0.375 11.265 0.455 ;
        RECT 12.065 0.375 12.235 0.455 ;
        RECT 12.635 0.625 12.805 0.910 ;
        RECT 13.120 1.580 13.775 1.750 ;
        RECT 14.935 1.675 15.105 1.755 ;
        RECT 15.905 1.675 16.075 1.755 ;
        RECT 16.875 1.675 17.045 1.755 ;
        RECT 13.120 0.845 13.290 1.580 ;
        RECT 14.935 1.505 17.045 1.675 ;
        RECT 13.605 0.625 13.775 1.395 ;
        RECT 12.635 0.455 13.775 0.625 ;
        RECT 12.635 0.375 12.805 0.455 ;
        RECT 13.605 0.375 13.775 0.455 ;
        RECT 14.935 0.375 15.105 1.505 ;
        RECT 15.905 0.625 16.075 1.505 ;
        RECT 16.875 1.425 17.045 1.505 ;
        RECT 16.395 1.080 16.565 1.160 ;
        RECT 17.445 1.080 17.615 1.755 ;
        RECT 18.415 1.750 18.585 5.070 ;
        RECT 20.265 1.915 20.435 4.865 ;
        RECT 16.395 0.910 17.615 1.080 ;
        RECT 16.395 0.830 16.565 0.910 ;
        RECT 16.875 0.625 17.045 0.705 ;
        RECT 15.905 0.455 17.045 0.625 ;
        RECT 15.905 0.375 16.075 0.455 ;
        RECT 16.875 0.375 17.045 0.455 ;
        RECT 17.445 0.625 17.615 0.910 ;
        RECT 17.930 1.580 18.585 1.750 ;
        RECT 19.745 1.675 19.915 1.755 ;
        RECT 20.715 1.675 20.885 1.755 ;
        RECT 21.685 1.675 21.855 1.755 ;
        RECT 17.930 0.845 18.100 1.580 ;
        RECT 19.745 1.505 21.855 1.675 ;
        RECT 18.415 0.625 18.585 1.395 ;
        RECT 17.445 0.455 18.585 0.625 ;
        RECT 17.445 0.375 17.615 0.455 ;
        RECT 18.415 0.375 18.585 0.455 ;
        RECT 19.745 0.375 19.915 1.505 ;
        RECT 20.715 0.625 20.885 1.505 ;
        RECT 21.685 1.425 21.855 1.505 ;
        RECT 21.205 1.080 21.375 1.160 ;
        RECT 22.255 1.080 22.425 1.755 ;
        RECT 23.225 1.750 23.395 5.070 ;
        RECT 25.075 1.915 25.245 4.865 ;
        RECT 27.295 1.915 27.465 4.865 ;
        RECT 21.205 0.910 22.425 1.080 ;
        RECT 21.205 0.830 21.375 0.910 ;
        RECT 21.685 0.625 21.855 0.705 ;
        RECT 20.715 0.455 21.855 0.625 ;
        RECT 20.715 0.375 20.885 0.455 ;
        RECT 21.685 0.375 21.855 0.455 ;
        RECT 22.255 0.625 22.425 0.910 ;
        RECT 22.740 1.580 23.395 1.750 ;
        RECT 24.555 1.675 24.725 1.755 ;
        RECT 25.525 1.675 25.695 1.755 ;
        RECT 26.495 1.675 26.665 1.755 ;
        RECT 22.740 0.845 22.910 1.580 ;
        RECT 24.555 1.505 26.665 1.675 ;
        RECT 23.225 0.625 23.395 1.395 ;
        RECT 22.255 0.455 23.395 0.625 ;
        RECT 22.255 0.375 22.425 0.455 ;
        RECT 23.225 0.375 23.395 0.455 ;
        RECT 24.555 0.375 24.725 1.505 ;
        RECT 25.525 0.625 25.695 1.505 ;
        RECT 26.495 1.425 26.665 1.505 ;
        RECT 26.015 1.080 26.185 1.160 ;
        RECT 27.065 1.080 27.235 1.755 ;
        RECT 26.015 0.910 27.235 1.080 ;
        RECT 26.015 0.830 26.185 0.910 ;
        RECT 26.495 0.625 26.665 0.705 ;
        RECT 25.525 0.455 26.665 0.625 ;
        RECT 25.525 0.375 25.695 0.455 ;
        RECT 26.495 0.375 26.665 0.455 ;
        RECT 27.065 0.625 27.235 0.910 ;
        RECT 28.035 0.625 28.205 1.395 ;
        RECT 27.065 0.455 28.205 0.625 ;
        RECT 27.065 0.375 27.235 0.455 ;
        RECT 28.035 0.375 28.205 0.455 ;
      LAYER mcon ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 2.880 4.155 3.050 ;
        RECT 8.050 3.985 8.220 4.155 ;
        RECT 5.835 2.880 6.005 3.050 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 2.880 10.815 3.050 ;
        RECT 12.865 3.985 13.035 4.155 ;
        RECT 13.605 2.875 13.775 3.045 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 20.265 3.615 20.435 3.785 ;
        RECT 23.225 3.245 23.395 3.415 ;
        RECT 25.075 3.245 25.245 3.415 ;
        RECT 27.295 3.985 27.465 4.155 ;
      LAYER met1 ;
        RECT 8.020 4.155 8.250 4.185 ;
        RECT 12.835 4.155 13.065 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 7.990 3.985 27.525 4.155 ;
        RECT 8.020 3.955 8.250 3.985 ;
        RECT 12.835 3.955 13.065 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 20.235 3.785 20.465 3.815 ;
        RECT 3.185 3.615 20.495 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 20.235 3.585 20.465 3.615 ;
        RECT 23.195 3.415 23.425 3.445 ;
        RECT 25.045 3.415 25.275 3.445 ;
        RECT 23.165 3.245 25.305 3.415 ;
        RECT 23.195 3.215 23.425 3.245 ;
        RECT 25.045 3.215 25.275 3.245 ;
        RECT 3.955 3.050 4.185 3.080 ;
        RECT 5.805 3.050 6.035 3.080 ;
        RECT 10.615 3.050 10.845 3.080 ;
        RECT 3.925 2.880 10.875 3.050 ;
        RECT 13.575 3.045 13.805 3.075 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 3.955 2.850 4.185 2.880 ;
        RECT 5.805 2.850 6.035 2.880 ;
        RECT 10.615 2.850 10.845 2.880 ;
        RECT 13.545 2.875 15.685 3.045 ;
        RECT 13.575 2.845 13.805 2.875 ;
        RECT 15.425 2.845 15.655 2.875 ;
  END
END DFFSNRNQX1






MACRO DFFSNRNX1
  CLASS CORE ;
  FOREIGN DFFSNRNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 28.860 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 25.495 5.240 25.665 7.020 ;
        RECT 26.375 5.240 26.545 7.020 ;
        RECT 27.255 5.240 27.425 7.020 ;
        RECT 25.495 5.070 28.205 5.240 ;
        RECT 22.485 1.915 22.655 4.865 ;
        RECT 28.035 1.750 28.205 5.070 ;
        RECT 27.550 1.580 28.205 1.750 ;
        RECT 27.550 0.845 27.720 1.580 ;
      LAYER mcon ;
        RECT 22.485 3.615 22.655 3.785 ;
        RECT 28.035 3.615 28.205 3.785 ;
      LAYER met1 ;
        RECT 22.455 3.785 22.685 3.815 ;
        RECT 28.005 3.785 28.235 3.815 ;
        RECT 22.425 3.615 28.265 3.785 ;
        RECT 22.455 3.585 22.685 3.615 ;
        RECT 28.005 3.585 28.235 3.615 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 20.685 5.240 20.855 7.020 ;
        RECT 21.565 5.240 21.735 7.020 ;
        RECT 22.445 5.240 22.615 7.020 ;
        RECT 20.685 5.070 23.395 5.240 ;
        RECT 23.225 1.750 23.395 5.070 ;
        RECT 25.075 1.915 25.245 4.865 ;
        RECT 22.740 1.580 23.395 1.750 ;
        RECT 22.740 0.845 22.910 1.580 ;
      LAYER mcon ;
        RECT 23.225 3.245 23.395 3.415 ;
        RECT 25.075 3.245 25.245 3.415 ;
      LAYER met1 ;
        RECT 23.195 3.415 23.425 3.445 ;
        RECT 25.045 3.415 25.275 3.445 ;
        RECT 23.165 3.245 25.305 3.415 ;
        RECT 23.195 3.215 23.425 3.245 ;
        RECT 25.045 3.215 25.275 3.245 ;
    END
  END QN
  PIN CLK
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 16.565 1.915 16.735 4.865 ;
      LAYER mcon ;
        RECT 6.945 3.245 7.115 3.415 ;
        RECT 16.565 3.245 16.735 3.415 ;
      LAYER met1 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 16.535 3.415 16.765 3.445 ;
        RECT 6.885 3.245 16.795 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
        RECT 16.535 3.215 16.765 3.245 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 11.755 1.915 11.925 4.865 ;
        RECT 26.185 1.915 26.355 4.865 ;
      LAYER mcon ;
        RECT 11.755 2.505 11.925 2.675 ;
        RECT 26.185 2.505 26.355 2.675 ;
      LAYER met1 ;
        RECT 11.725 2.675 11.955 2.705 ;
        RECT 26.155 2.675 26.385 2.705 ;
        RECT 11.695 2.505 26.415 2.675 ;
        RECT 11.725 2.475 11.955 2.505 ;
        RECT 26.155 2.475 26.385 2.505 ;
    END
  END SN
  PIN RN
    ANTENNAGATEAREA 3.056950 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 17.675 1.915 17.845 4.865 ;
        RECT 21.375 1.915 21.545 4.865 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 17.675 4.355 17.845 4.525 ;
        RECT 21.375 4.355 21.545 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 17.645 4.525 17.875 4.555 ;
        RECT 21.345 4.525 21.575 4.555 ;
        RECT 2.075 4.355 21.605 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 17.645 4.325 17.875 4.355 ;
        RECT 21.345 4.325 21.575 4.355 ;
    END
  END RN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 29.295 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 29.030 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.625 5.215 10.795 7.230 ;
        RECT 11.505 5.555 11.675 7.230 ;
        RECT 12.385 5.555 12.555 7.230 ;
        RECT 13.265 5.555 13.435 7.230 ;
        RECT 14.260 4.110 14.600 7.230 ;
        RECT 15.435 5.215 15.605 7.230 ;
        RECT 16.315 5.555 16.485 7.230 ;
        RECT 17.195 5.555 17.365 7.230 ;
        RECT 18.075 5.555 18.245 7.230 ;
        RECT 19.070 4.110 19.410 7.230 ;
        RECT 20.245 5.215 20.415 7.230 ;
        RECT 21.125 5.555 21.295 7.230 ;
        RECT 22.005 5.555 22.175 7.230 ;
        RECT 22.885 5.555 23.055 7.230 ;
        RECT 23.880 4.110 24.220 7.230 ;
        RECT 25.055 5.215 25.225 7.230 ;
        RECT 25.935 5.555 26.105 7.230 ;
        RECT 26.815 5.555 26.985 7.230 ;
        RECT 27.695 5.555 27.865 7.230 ;
        RECT 28.690 4.110 29.030 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 29.030 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 29.030 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.610 0.170 10.780 1.130 ;
        RECT 14.260 0.170 14.600 2.720 ;
        RECT 15.420 0.170 15.590 1.130 ;
        RECT 19.070 0.170 19.410 2.720 ;
        RECT 20.230 0.170 20.400 1.130 ;
        RECT 23.880 0.170 24.220 2.720 ;
        RECT 25.040 0.170 25.210 1.130 ;
        RECT 28.690 0.170 29.030 2.720 ;
        RECT -0.170 -0.170 29.030 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 29.030 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 11.065 5.240 11.235 7.020 ;
        RECT 11.945 5.240 12.115 7.020 ;
        RECT 12.825 5.240 12.995 7.020 ;
        RECT 15.875 5.240 16.045 7.020 ;
        RECT 16.755 5.240 16.925 7.020 ;
        RECT 17.635 5.240 17.805 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 11.065 5.070 13.775 5.240 ;
        RECT 15.875 5.070 18.585 5.240 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 8.055 4.235 8.225 4.865 ;
        RECT 8.050 3.905 8.225 4.235 ;
        RECT 8.055 1.915 8.225 3.905 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 12.865 1.915 13.035 4.865 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.125 1.675 10.295 1.755 ;
        RECT 11.095 1.675 11.265 1.755 ;
        RECT 12.065 1.675 12.235 1.755 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.125 1.505 12.235 1.675 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.125 0.375 10.295 1.505 ;
        RECT 11.095 0.625 11.265 1.505 ;
        RECT 12.065 1.425 12.235 1.505 ;
        RECT 11.585 1.080 11.755 1.160 ;
        RECT 12.635 1.080 12.805 1.755 ;
        RECT 13.605 1.750 13.775 5.070 ;
        RECT 15.455 1.915 15.625 4.865 ;
        RECT 11.585 0.910 12.805 1.080 ;
        RECT 11.585 0.830 11.755 0.910 ;
        RECT 12.065 0.625 12.235 0.705 ;
        RECT 11.095 0.455 12.235 0.625 ;
        RECT 11.095 0.375 11.265 0.455 ;
        RECT 12.065 0.375 12.235 0.455 ;
        RECT 12.635 0.625 12.805 0.910 ;
        RECT 13.120 1.580 13.775 1.750 ;
        RECT 14.935 1.675 15.105 1.755 ;
        RECT 15.905 1.675 16.075 1.755 ;
        RECT 16.875 1.675 17.045 1.755 ;
        RECT 13.120 0.845 13.290 1.580 ;
        RECT 14.935 1.505 17.045 1.675 ;
        RECT 13.605 0.625 13.775 1.395 ;
        RECT 12.635 0.455 13.775 0.625 ;
        RECT 12.635 0.375 12.805 0.455 ;
        RECT 13.605 0.375 13.775 0.455 ;
        RECT 14.935 0.375 15.105 1.505 ;
        RECT 15.905 0.625 16.075 1.505 ;
        RECT 16.875 1.425 17.045 1.505 ;
        RECT 16.395 1.080 16.565 1.160 ;
        RECT 17.445 1.080 17.615 1.755 ;
        RECT 18.415 1.750 18.585 5.070 ;
        RECT 20.265 1.915 20.435 4.865 ;
        RECT 27.295 1.915 27.465 4.865 ;
        RECT 16.395 0.910 17.615 1.080 ;
        RECT 16.395 0.830 16.565 0.910 ;
        RECT 16.875 0.625 17.045 0.705 ;
        RECT 15.905 0.455 17.045 0.625 ;
        RECT 15.905 0.375 16.075 0.455 ;
        RECT 16.875 0.375 17.045 0.455 ;
        RECT 17.445 0.625 17.615 0.910 ;
        RECT 17.930 1.580 18.585 1.750 ;
        RECT 19.745 1.675 19.915 1.755 ;
        RECT 20.715 1.675 20.885 1.755 ;
        RECT 21.685 1.675 21.855 1.755 ;
        RECT 17.930 0.845 18.100 1.580 ;
        RECT 19.745 1.505 21.855 1.675 ;
        RECT 18.415 0.625 18.585 1.395 ;
        RECT 17.445 0.455 18.585 0.625 ;
        RECT 17.445 0.375 17.615 0.455 ;
        RECT 18.415 0.375 18.585 0.455 ;
        RECT 19.745 0.375 19.915 1.505 ;
        RECT 20.715 0.625 20.885 1.505 ;
        RECT 21.685 1.425 21.855 1.505 ;
        RECT 21.205 1.080 21.375 1.160 ;
        RECT 22.255 1.080 22.425 1.755 ;
        RECT 24.555 1.675 24.725 1.755 ;
        RECT 25.525 1.675 25.695 1.755 ;
        RECT 26.495 1.675 26.665 1.755 ;
        RECT 24.555 1.505 26.665 1.675 ;
        RECT 21.205 0.910 22.425 1.080 ;
        RECT 21.205 0.830 21.375 0.910 ;
        RECT 21.685 0.625 21.855 0.705 ;
        RECT 20.715 0.455 21.855 0.625 ;
        RECT 20.715 0.375 20.885 0.455 ;
        RECT 21.685 0.375 21.855 0.455 ;
        RECT 22.255 0.625 22.425 0.910 ;
        RECT 23.225 0.625 23.395 1.395 ;
        RECT 22.255 0.455 23.395 0.625 ;
        RECT 22.255 0.375 22.425 0.455 ;
        RECT 23.225 0.375 23.395 0.455 ;
        RECT 24.555 0.375 24.725 1.505 ;
        RECT 25.525 0.625 25.695 1.505 ;
        RECT 26.495 1.425 26.665 1.505 ;
        RECT 26.015 1.080 26.185 1.160 ;
        RECT 27.065 1.080 27.235 1.755 ;
        RECT 26.015 0.910 27.235 1.080 ;
        RECT 26.015 0.830 26.185 0.910 ;
        RECT 26.495 0.625 26.665 0.705 ;
        RECT 25.525 0.455 26.665 0.625 ;
        RECT 25.525 0.375 25.695 0.455 ;
        RECT 26.495 0.375 26.665 0.455 ;
        RECT 27.065 0.625 27.235 0.910 ;
        RECT 28.035 0.625 28.205 1.395 ;
        RECT 27.065 0.455 28.205 0.625 ;
        RECT 27.065 0.375 27.235 0.455 ;
        RECT 28.035 0.375 28.205 0.455 ;
      LAYER mcon ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 3.985 2.880 4.155 3.050 ;
        RECT 8.050 3.985 8.220 4.155 ;
        RECT 5.835 2.880 6.005 3.050 ;
        RECT 8.795 3.615 8.965 3.785 ;
        RECT 10.645 2.880 10.815 3.050 ;
        RECT 12.865 3.985 13.035 4.155 ;
        RECT 13.605 2.875 13.775 3.045 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 20.265 3.615 20.435 3.785 ;
        RECT 27.295 3.985 27.465 4.155 ;
      LAYER met1 ;
        RECT 8.020 4.155 8.250 4.185 ;
        RECT 12.835 4.155 13.065 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 27.265 4.155 27.495 4.185 ;
        RECT 7.990 3.985 27.525 4.155 ;
        RECT 8.020 3.955 8.250 3.985 ;
        RECT 12.835 3.955 13.065 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 27.265 3.955 27.495 3.985 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 8.765 3.785 8.995 3.815 ;
        RECT 20.235 3.785 20.465 3.815 ;
        RECT 3.185 3.615 20.495 3.785 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 8.765 3.585 8.995 3.615 ;
        RECT 20.235 3.585 20.465 3.615 ;
        RECT 3.955 3.050 4.185 3.080 ;
        RECT 5.805 3.050 6.035 3.080 ;
        RECT 10.615 3.050 10.845 3.080 ;
        RECT 3.925 2.880 10.875 3.050 ;
        RECT 13.575 3.045 13.805 3.075 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 3.955 2.850 4.185 2.880 ;
        RECT 5.805 2.850 6.035 2.880 ;
        RECT 10.615 2.850 10.845 2.880 ;
        RECT 13.545 2.875 15.685 3.045 ;
        RECT 13.575 2.845 13.805 2.875 ;
        RECT 15.425 2.845 15.655 2.875 ;
  END
END DFFSNRNX1






MACRO DFFSNX1
  CLASS CORE ;
  FOREIGN DFFSNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.420 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.931900 ;
    PORT
      LAYER li1 ;
        RECT 21.055 5.240 21.225 7.020 ;
        RECT 21.935 5.240 22.105 7.020 ;
        RECT 22.815 5.240 22.985 7.020 ;
        RECT 21.055 5.070 23.765 5.240 ;
        RECT 18.075 4.710 18.245 4.865 ;
        RECT 18.045 4.535 18.245 4.710 ;
        RECT 18.045 1.915 18.215 4.535 ;
        RECT 23.595 1.750 23.765 5.070 ;
        RECT 23.110 1.580 23.765 1.750 ;
        RECT 23.110 0.845 23.280 1.580 ;
      LAYER mcon ;
        RECT 18.045 3.985 18.215 4.155 ;
        RECT 23.595 3.985 23.765 4.155 ;
      LAYER met1 ;
        RECT 18.015 4.155 18.245 4.185 ;
        RECT 23.565 4.155 23.795 4.185 ;
        RECT 17.985 3.985 23.825 4.155 ;
        RECT 18.015 3.955 18.245 3.985 ;
        RECT 23.565 3.955 23.795 3.985 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 17.425 5.285 17.595 7.020 ;
        RECT 18.305 5.285 18.475 7.020 ;
        RECT 17.425 5.115 18.955 5.285 ;
        RECT 18.785 1.740 18.955 5.115 ;
        RECT 20.635 1.915 20.805 4.865 ;
        RECT 18.345 1.570 18.955 1.740 ;
        RECT 18.345 0.835 18.515 1.570 ;
      LAYER mcon ;
        RECT 18.785 2.875 18.955 3.045 ;
        RECT 20.635 2.875 20.805 3.045 ;
      LAYER met1 ;
        RECT 18.755 3.045 18.985 3.075 ;
        RECT 20.605 3.045 20.835 3.075 ;
        RECT 18.725 2.875 20.865 3.045 ;
        RECT 18.755 2.845 18.985 2.875 ;
        RECT 20.605 2.845 20.835 2.875 ;
    END
  END QN
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 5.465 1.915 5.635 4.865 ;
        RECT 14.745 4.710 14.915 4.865 ;
        RECT 14.715 4.535 14.915 4.710 ;
        RECT 14.715 1.915 14.885 4.535 ;
      LAYER mcon ;
        RECT 5.465 4.355 5.635 4.525 ;
        RECT 14.715 4.355 14.885 4.525 ;
      LAYER met1 ;
        RECT 5.435 4.525 5.665 4.555 ;
        RECT 14.685 4.525 14.915 4.555 ;
        RECT 5.405 4.355 14.945 4.525 ;
        RECT 5.435 4.325 5.665 4.355 ;
        RECT 14.685 4.325 14.915 4.355 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 2.029700 ;
    PORT
      LAYER li1 ;
        RECT 10.275 1.915 10.445 4.865 ;
        RECT 21.745 1.915 21.915 4.865 ;
      LAYER mcon ;
        RECT 10.275 2.135 10.445 2.305 ;
        RECT 21.745 2.135 21.915 2.305 ;
      LAYER met1 ;
        RECT 10.245 2.305 10.475 2.335 ;
        RECT 21.715 2.305 21.945 2.335 ;
        RECT 10.215 2.135 21.975 2.305 ;
        RECT 10.245 2.105 10.475 2.135 ;
        RECT 21.715 2.105 21.945 2.135 ;
    END
  END SN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 24.855 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 24.590 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.335 5.215 4.505 7.230 ;
        RECT 5.215 5.555 5.385 7.230 ;
        RECT 6.095 5.555 6.265 7.230 ;
        RECT 6.975 5.555 7.145 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 9.145 5.215 9.315 7.230 ;
        RECT 10.025 5.555 10.195 7.230 ;
        RECT 10.905 5.555 11.075 7.230 ;
        RECT 11.785 5.555 11.955 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.655 5.135 13.825 7.230 ;
        RECT 14.535 5.555 14.705 7.230 ;
        RECT 15.415 5.555 15.585 7.230 ;
        RECT 16.110 4.110 16.450 7.230 ;
        RECT 16.985 5.135 17.155 7.230 ;
        RECT 17.865 5.555 18.035 7.230 ;
        RECT 18.745 5.555 18.915 7.230 ;
        RECT 19.440 4.110 19.780 7.230 ;
        RECT 20.615 5.215 20.785 7.230 ;
        RECT 21.495 5.555 21.665 7.230 ;
        RECT 22.375 5.555 22.545 7.230 ;
        RECT 23.255 5.555 23.425 7.230 ;
        RECT 24.250 4.110 24.590 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 24.590 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 24.590 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 4.320 0.170 4.490 1.130 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.130 0.170 9.300 1.130 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 14.045 0.170 14.215 1.120 ;
        RECT 16.110 0.170 16.450 2.720 ;
        RECT 17.375 0.170 17.545 1.120 ;
        RECT 19.440 0.170 19.780 2.720 ;
        RECT 20.600 0.170 20.770 1.130 ;
        RECT 24.250 0.170 24.590 2.720 ;
        RECT -0.170 -0.170 24.590 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 24.590 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.775 5.240 4.945 7.020 ;
        RECT 5.655 5.240 5.825 7.020 ;
        RECT 6.535 5.240 6.705 7.020 ;
        RECT 9.585 5.240 9.755 7.020 ;
        RECT 10.465 5.240 10.635 7.020 ;
        RECT 11.345 5.240 11.515 7.020 ;
        RECT 14.095 5.285 14.265 7.020 ;
        RECT 14.975 5.285 15.145 7.020 ;
        RECT 4.775 5.070 7.485 5.240 ;
        RECT 9.585 5.070 12.295 5.240 ;
        RECT 14.095 5.115 15.625 5.285 ;
        RECT 4.355 1.915 4.525 4.865 ;
        RECT 6.575 1.915 6.745 4.865 ;
        RECT 7.315 4.235 7.485 5.070 ;
        RECT 7.310 3.905 7.485 4.235 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 3.835 1.675 4.005 1.755 ;
        RECT 4.805 1.675 4.975 1.755 ;
        RECT 5.775 1.675 5.945 1.755 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 3.835 1.505 5.945 1.675 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 3.835 0.375 4.005 1.505 ;
        RECT 4.805 0.625 4.975 1.505 ;
        RECT 5.775 1.425 5.945 1.505 ;
        RECT 5.295 1.080 5.465 1.160 ;
        RECT 6.345 1.080 6.515 1.755 ;
        RECT 7.315 1.750 7.485 3.905 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 11.385 1.915 11.555 4.865 ;
        RECT 5.295 0.910 6.515 1.080 ;
        RECT 5.295 0.830 5.465 0.910 ;
        RECT 5.775 0.625 5.945 0.705 ;
        RECT 4.805 0.455 5.945 0.625 ;
        RECT 4.805 0.375 4.975 0.455 ;
        RECT 5.775 0.375 5.945 0.455 ;
        RECT 6.345 0.625 6.515 0.910 ;
        RECT 6.830 1.580 7.485 1.750 ;
        RECT 8.645 1.675 8.815 1.755 ;
        RECT 9.615 1.675 9.785 1.755 ;
        RECT 10.585 1.675 10.755 1.755 ;
        RECT 6.830 0.845 7.000 1.580 ;
        RECT 8.645 1.505 10.755 1.675 ;
        RECT 7.315 0.625 7.485 1.395 ;
        RECT 6.345 0.455 7.485 0.625 ;
        RECT 6.345 0.375 6.515 0.455 ;
        RECT 7.315 0.375 7.485 0.455 ;
        RECT 8.645 0.375 8.815 1.505 ;
        RECT 9.615 0.625 9.785 1.505 ;
        RECT 10.585 1.425 10.755 1.505 ;
        RECT 10.105 1.080 10.275 1.160 ;
        RECT 11.155 1.080 11.325 1.755 ;
        RECT 12.125 1.750 12.295 5.070 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 10.105 0.910 11.325 1.080 ;
        RECT 10.105 0.830 10.275 0.910 ;
        RECT 10.585 0.625 10.755 0.705 ;
        RECT 9.615 0.455 10.755 0.625 ;
        RECT 9.615 0.375 9.785 0.455 ;
        RECT 10.585 0.375 10.755 0.455 ;
        RECT 11.155 0.625 11.325 0.910 ;
        RECT 11.640 1.580 12.295 1.750 ;
        RECT 13.560 1.665 13.730 1.745 ;
        RECT 14.530 1.665 14.700 1.745 ;
        RECT 15.455 1.740 15.625 5.115 ;
        RECT 17.305 1.915 17.475 4.865 ;
        RECT 22.855 1.915 23.025 4.865 ;
        RECT 11.640 0.845 11.810 1.580 ;
        RECT 13.560 1.495 14.700 1.665 ;
        RECT 12.125 0.625 12.295 1.395 ;
        RECT 11.155 0.455 12.295 0.625 ;
        RECT 11.155 0.375 11.325 0.455 ;
        RECT 12.125 0.375 12.295 0.455 ;
        RECT 13.560 0.365 13.730 1.495 ;
        RECT 14.530 0.615 14.700 1.495 ;
        RECT 15.015 1.570 15.625 1.740 ;
        RECT 16.890 1.665 17.060 1.745 ;
        RECT 17.860 1.665 18.030 1.745 ;
        RECT 15.015 0.835 15.185 1.570 ;
        RECT 16.890 1.495 18.030 1.665 ;
        RECT 15.500 0.615 15.670 1.385 ;
        RECT 14.530 0.445 15.670 0.615 ;
        RECT 14.530 0.365 14.700 0.445 ;
        RECT 15.500 0.365 15.670 0.445 ;
        RECT 16.890 0.365 17.060 1.495 ;
        RECT 17.860 0.615 18.030 1.495 ;
        RECT 20.115 1.675 20.285 1.755 ;
        RECT 21.085 1.675 21.255 1.755 ;
        RECT 22.055 1.675 22.225 1.755 ;
        RECT 20.115 1.505 22.225 1.675 ;
        RECT 18.830 0.615 19.000 1.385 ;
        RECT 17.860 0.445 19.000 0.615 ;
        RECT 17.860 0.365 18.030 0.445 ;
        RECT 18.830 0.365 19.000 0.445 ;
        RECT 20.115 0.375 20.285 1.505 ;
        RECT 21.085 0.625 21.255 1.505 ;
        RECT 22.055 1.425 22.225 1.505 ;
        RECT 21.575 1.080 21.745 1.160 ;
        RECT 22.625 1.080 22.795 1.755 ;
        RECT 21.575 0.910 22.795 1.080 ;
        RECT 21.575 0.830 21.745 0.910 ;
        RECT 22.055 0.625 22.225 0.705 ;
        RECT 21.085 0.455 22.225 0.625 ;
        RECT 21.085 0.375 21.255 0.455 ;
        RECT 22.055 0.375 22.225 0.455 ;
        RECT 22.625 0.625 22.795 0.910 ;
        RECT 23.595 0.625 23.765 1.395 ;
        RECT 22.625 0.455 23.765 0.625 ;
        RECT 22.625 0.375 22.795 0.455 ;
        RECT 23.595 0.375 23.765 0.455 ;
      LAYER mcon ;
        RECT 1.765 3.985 1.935 4.155 ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.500 4.525 2.670 ;
        RECT 7.310 3.985 7.480 4.155 ;
        RECT 6.575 3.615 6.745 3.785 ;
        RECT 9.165 2.505 9.335 2.675 ;
        RECT 11.385 3.615 11.555 3.785 ;
        RECT 12.125 2.505 12.295 2.675 ;
        RECT 13.975 2.505 14.145 2.675 ;
        RECT 15.455 3.615 15.625 3.785 ;
        RECT 17.305 3.985 17.475 4.155 ;
        RECT 22.855 3.615 23.025 3.785 ;
      LAYER met1 ;
        RECT 1.735 4.155 1.965 4.185 ;
        RECT 7.280 4.155 7.510 4.185 ;
        RECT 17.275 4.155 17.505 4.185 ;
        RECT 1.705 3.985 17.535 4.155 ;
        RECT 1.735 3.955 1.965 3.985 ;
        RECT 7.280 3.955 7.510 3.985 ;
        RECT 17.275 3.955 17.505 3.985 ;
        RECT 6.545 3.785 6.775 3.815 ;
        RECT 11.355 3.785 11.585 3.815 ;
        RECT 15.425 3.785 15.655 3.815 ;
        RECT 22.825 3.785 23.055 3.815 ;
        RECT 6.515 3.615 23.085 3.785 ;
        RECT 6.545 3.585 6.775 3.615 ;
        RECT 11.355 3.585 11.585 3.615 ;
        RECT 15.425 3.585 15.655 3.615 ;
        RECT 22.825 3.585 23.055 3.615 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.700 ;
        RECT 9.135 2.675 9.365 2.705 ;
        RECT 12.095 2.675 12.325 2.705 ;
        RECT 13.945 2.675 14.175 2.705 ;
        RECT 2.445 2.505 9.395 2.675 ;
        RECT 12.065 2.505 14.205 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.295 2.500 4.705 2.505 ;
        RECT 4.325 2.470 4.555 2.500 ;
        RECT 9.135 2.475 9.365 2.505 ;
        RECT 12.095 2.475 12.325 2.505 ;
        RECT 13.945 2.475 14.175 2.505 ;
  END
END DFFSNX1






MACRO DFFX1
  CLASS CORE ;
  FOREIGN DFFX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.460 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 19.275 5.285 19.445 7.020 ;
        RECT 20.155 5.285 20.325 7.020 ;
        RECT 19.275 5.115 20.805 5.285 ;
        RECT 16.595 4.710 16.765 4.865 ;
        RECT 16.565 4.535 16.765 4.710 ;
        RECT 16.565 1.915 16.735 4.535 ;
        RECT 20.635 1.740 20.805 5.115 ;
        RECT 20.195 1.570 20.805 1.740 ;
        RECT 20.195 0.835 20.365 1.570 ;
      LAYER mcon ;
        RECT 16.565 3.615 16.735 3.785 ;
        RECT 20.635 3.615 20.805 3.785 ;
      LAYER met1 ;
        RECT 16.535 3.785 16.765 3.815 ;
        RECT 20.605 3.785 20.835 3.815 ;
        RECT 16.505 3.615 20.865 3.785 ;
        RECT 16.535 3.585 16.765 3.615 ;
        RECT 20.605 3.585 20.835 3.615 ;
    END
  END Q
  PIN QN
    ANTENNAGATEAREA 1.033250 ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 15.945 5.285 16.115 7.020 ;
        RECT 16.825 5.285 16.995 7.020 ;
        RECT 15.945 5.115 17.475 5.285 ;
        RECT 17.305 1.740 17.475 5.115 ;
        RECT 19.155 1.915 19.325 4.865 ;
        RECT 16.865 1.570 17.475 1.740 ;
        RECT 16.865 0.835 17.035 1.570 ;
      LAYER mcon ;
        RECT 17.305 3.245 17.475 3.415 ;
        RECT 19.155 3.245 19.325 3.415 ;
      LAYER met1 ;
        RECT 17.275 3.415 17.505 3.445 ;
        RECT 19.125 3.415 19.355 3.445 ;
        RECT 17.245 3.245 19.385 3.415 ;
        RECT 17.275 3.215 17.505 3.245 ;
        RECT 19.125 3.215 19.355 3.245 ;
    END
  END QN
  PIN CLK
    ANTENNAGATEAREA 2.042100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 13.265 4.710 13.435 4.865 ;
        RECT 13.235 4.535 13.435 4.710 ;
        RECT 13.235 1.915 13.405 4.535 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 13.235 4.355 13.405 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 13.205 4.525 13.435 4.555 ;
        RECT 2.075 4.355 13.465 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 13.205 4.325 13.435 4.355 ;
    END
  END CLK
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 21.895 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 21.630 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.515 5.135 5.685 7.230 ;
        RECT 6.395 5.555 6.565 7.230 ;
        RECT 7.275 5.555 7.445 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 8.845 5.135 9.015 7.230 ;
        RECT 9.725 5.555 9.895 7.230 ;
        RECT 10.605 5.555 10.775 7.230 ;
        RECT 11.300 4.110 11.640 7.230 ;
        RECT 12.175 5.135 12.345 7.230 ;
        RECT 13.055 5.555 13.225 7.230 ;
        RECT 13.935 5.555 14.105 7.230 ;
        RECT 14.630 4.110 14.970 7.230 ;
        RECT 15.505 5.135 15.675 7.230 ;
        RECT 16.385 5.555 16.555 7.230 ;
        RECT 17.265 5.555 17.435 7.230 ;
        RECT 17.960 4.110 18.300 7.230 ;
        RECT 18.835 5.135 19.005 7.230 ;
        RECT 19.715 5.555 19.885 7.230 ;
        RECT 20.595 5.555 20.765 7.230 ;
        RECT 21.290 4.110 21.630 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.225 21.630 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 21.630 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.905 0.170 6.075 1.120 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.235 0.170 9.405 1.120 ;
        RECT 11.300 0.170 11.640 2.720 ;
        RECT 12.565 0.170 12.735 1.120 ;
        RECT 14.630 0.170 14.970 2.720 ;
        RECT 15.895 0.170 16.065 1.120 ;
        RECT 17.960 0.170 18.300 2.720 ;
        RECT 19.225 0.170 19.395 1.120 ;
        RECT 21.290 0.170 21.630 2.720 ;
        RECT -0.170 -0.170 21.630 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 21.630 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 5.955 5.285 6.125 7.020 ;
        RECT 6.835 5.285 7.005 7.020 ;
        RECT 9.285 5.285 9.455 7.020 ;
        RECT 10.165 5.285 10.335 7.020 ;
        RECT 12.615 5.285 12.785 7.020 ;
        RECT 13.495 5.285 13.665 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 5.955 5.115 7.485 5.285 ;
        RECT 9.285 5.115 10.815 5.285 ;
        RECT 12.615 5.115 14.145 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 6.605 4.710 6.775 4.865 ;
        RECT 6.575 4.535 6.775 4.710 ;
        RECT 6.575 1.915 6.745 4.535 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.420 1.665 5.590 1.745 ;
        RECT 6.390 1.665 6.560 1.745 ;
        RECT 7.315 1.740 7.485 5.115 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 9.935 4.710 10.105 4.865 ;
        RECT 9.905 4.535 10.105 4.710 ;
        RECT 9.905 1.915 10.075 4.535 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.420 1.495 6.560 1.665 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.420 0.365 5.590 1.495 ;
        RECT 6.390 0.615 6.560 1.495 ;
        RECT 6.875 1.570 7.485 1.740 ;
        RECT 8.750 1.665 8.920 1.745 ;
        RECT 9.720 1.665 9.890 1.745 ;
        RECT 10.645 1.740 10.815 5.115 ;
        RECT 12.495 1.915 12.665 4.865 ;
        RECT 6.875 0.835 7.045 1.570 ;
        RECT 8.750 1.495 9.890 1.665 ;
        RECT 7.360 0.615 7.530 1.385 ;
        RECT 6.390 0.445 7.530 0.615 ;
        RECT 6.390 0.365 6.560 0.445 ;
        RECT 7.360 0.365 7.530 0.445 ;
        RECT 8.750 0.365 8.920 1.495 ;
        RECT 9.720 0.615 9.890 1.495 ;
        RECT 10.205 1.570 10.815 1.740 ;
        RECT 12.080 1.665 12.250 1.745 ;
        RECT 13.050 1.665 13.220 1.745 ;
        RECT 13.975 1.740 14.145 5.115 ;
        RECT 15.825 1.915 15.995 4.865 ;
        RECT 19.925 4.710 20.095 4.865 ;
        RECT 19.895 4.535 20.095 4.710 ;
        RECT 19.895 1.915 20.065 4.535 ;
        RECT 10.205 0.835 10.375 1.570 ;
        RECT 12.080 1.495 13.220 1.665 ;
        RECT 10.690 0.615 10.860 1.385 ;
        RECT 9.720 0.445 10.860 0.615 ;
        RECT 9.720 0.365 9.890 0.445 ;
        RECT 10.690 0.365 10.860 0.445 ;
        RECT 12.080 0.365 12.250 1.495 ;
        RECT 13.050 0.615 13.220 1.495 ;
        RECT 13.535 1.570 14.145 1.740 ;
        RECT 15.410 1.665 15.580 1.745 ;
        RECT 16.380 1.665 16.550 1.745 ;
        RECT 13.535 0.835 13.705 1.570 ;
        RECT 15.410 1.495 16.550 1.665 ;
        RECT 14.020 0.615 14.190 1.385 ;
        RECT 13.050 0.445 14.190 0.615 ;
        RECT 13.050 0.365 13.220 0.445 ;
        RECT 14.020 0.365 14.190 0.445 ;
        RECT 15.410 0.365 15.580 1.495 ;
        RECT 16.380 0.615 16.550 1.495 ;
        RECT 18.740 1.665 18.910 1.745 ;
        RECT 19.710 1.665 19.880 1.745 ;
        RECT 18.740 1.495 19.880 1.665 ;
        RECT 17.350 0.615 17.520 1.385 ;
        RECT 16.380 0.445 17.520 0.615 ;
        RECT 16.380 0.365 16.550 0.445 ;
        RECT 17.350 0.365 17.520 0.445 ;
        RECT 18.740 0.365 18.910 1.495 ;
        RECT 19.710 0.615 19.880 1.495 ;
        RECT 20.680 0.615 20.850 1.385 ;
        RECT 19.710 0.445 20.850 0.615 ;
        RECT 19.710 0.365 19.880 0.445 ;
        RECT 20.680 0.365 20.850 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 7.315 3.245 7.485 3.415 ;
        RECT 9.165 3.245 9.335 3.415 ;
        RECT 9.905 3.985 10.075 4.155 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 12.495 3.245 12.665 3.415 ;
        RECT 13.975 3.985 14.145 4.155 ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 19.895 3.985 20.065 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 9.875 4.155 10.105 4.185 ;
        RECT 13.945 4.155 14.175 4.185 ;
        RECT 19.865 4.155 20.095 4.185 ;
        RECT 0.965 3.985 20.125 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 9.875 3.955 10.105 3.985 ;
        RECT 13.945 3.955 14.175 3.985 ;
        RECT 19.865 3.955 20.095 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 3.925 3.615 16.055 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 7.285 3.415 7.515 3.445 ;
        RECT 9.135 3.415 9.365 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.465 3.415 12.695 3.445 ;
        RECT 3.185 3.245 9.395 3.415 ;
        RECT 10.585 3.245 12.725 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 7.285 3.215 7.515 3.245 ;
        RECT 9.135 3.215 9.365 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.465 3.215 12.695 3.245 ;
  END
END DFFX1






MACRO DLATCH
  CLASS CORE ;
  FOREIGN DLATCH ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.980 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 0.963050 ;
    PORT
      LAYER li1 ;
        RECT 15.345 5.295 15.515 6.565 ;
        RECT 15.345 5.125 15.995 5.295 ;
        RECT 15.825 1.740 15.995 5.125 ;
        RECT 17.520 4.710 17.690 4.870 ;
        RECT 17.520 4.540 17.845 4.710 ;
        RECT 17.675 1.915 17.845 4.540 ;
        RECT 14.415 1.570 15.995 1.740 ;
        RECT 14.415 0.835 14.585 1.570 ;
        RECT 15.385 0.835 15.555 1.570 ;
      LAYER mcon ;
        RECT 15.825 3.245 15.995 3.415 ;
        RECT 17.675 3.245 17.845 3.415 ;
      LAYER met1 ;
        RECT 15.795 3.415 16.025 3.445 ;
        RECT 17.645 3.415 17.875 3.445 ;
        RECT 15.765 3.245 17.905 3.415 ;
        RECT 15.795 3.215 16.025 3.245 ;
        RECT 17.645 3.215 17.875 3.245 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 2.054500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 9.565 4.710 9.735 4.865 ;
        RECT 9.535 4.535 9.735 4.710 ;
        RECT 9.535 1.915 9.705 4.535 ;
      LAYER mcon ;
        RECT 0.655 3.985 0.825 4.155 ;
        RECT 9.535 3.985 9.705 4.155 ;
      LAYER met1 ;
        RECT 0.625 4.155 0.855 4.185 ;
        RECT 9.505 4.155 9.735 4.185 ;
        RECT 0.595 3.985 9.765 4.155 ;
        RECT 0.625 3.955 0.855 3.985 ;
        RECT 9.505 3.955 9.735 3.985 ;
    END
  END D
  PIN GATE
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 4.015 4.710 4.185 4.865 ;
        RECT 3.985 4.535 4.185 4.710 ;
        RECT 3.985 1.915 4.155 4.535 ;
        RECT 8.795 1.915 8.965 4.865 ;
      LAYER mcon ;
        RECT 3.985 2.875 4.155 3.045 ;
        RECT 8.795 2.875 8.965 3.045 ;
      LAYER met1 ;
        RECT 3.955 3.045 4.185 3.075 ;
        RECT 8.765 3.045 8.995 3.075 ;
        RECT 3.925 2.875 9.025 3.045 ;
        RECT 3.955 2.845 4.185 2.875 ;
        RECT 8.765 2.845 8.995 2.875 ;
    END
  END GATE
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 20.415 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 20.150 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
        RECT 2.925 5.135 3.095 7.230 ;
        RECT 3.805 5.555 3.975 7.230 ;
        RECT 4.685 5.555 4.855 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
        RECT 6.140 5.185 6.310 7.230 ;
        RECT 7.020 5.185 7.190 7.230 ;
        RECT 7.600 4.110 7.940 7.230 ;
        RECT 8.475 5.135 8.645 7.230 ;
        RECT 9.355 5.555 9.525 7.230 ;
        RECT 10.235 5.555 10.405 7.230 ;
        RECT 10.930 4.110 11.270 7.230 ;
        RECT 11.690 5.185 11.860 7.230 ;
        RECT 12.570 5.185 12.740 7.230 ;
        RECT 13.150 4.110 13.490 7.230 ;
        RECT 14.465 5.555 14.635 7.230 ;
        RECT 16.480 4.110 16.820 7.230 ;
        RECT 17.795 5.555 17.965 7.230 ;
        RECT 19.810 4.110 20.150 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 20.150 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 20.150 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT 3.315 0.170 3.485 1.120 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT 6.095 0.620 6.265 1.750 ;
        RECT 7.065 0.620 7.235 1.750 ;
        RECT 6.095 0.450 7.235 0.620 ;
        RECT 6.095 0.170 6.265 0.450 ;
        RECT 6.580 0.170 6.750 0.450 ;
        RECT 7.065 0.170 7.235 0.450 ;
        RECT 7.600 0.170 7.940 2.720 ;
        RECT 8.865 0.170 9.035 1.120 ;
        RECT 10.930 0.170 11.270 2.720 ;
        RECT 11.645 0.620 11.815 1.750 ;
        RECT 12.615 0.620 12.785 1.750 ;
        RECT 11.645 0.450 12.785 0.620 ;
        RECT 11.645 0.170 11.815 0.450 ;
        RECT 12.130 0.170 12.300 0.450 ;
        RECT 12.615 0.170 12.785 0.450 ;
        RECT 13.150 0.170 13.490 2.720 ;
        RECT 13.930 0.615 14.100 1.745 ;
        RECT 14.900 0.615 15.070 1.390 ;
        RECT 15.870 0.615 16.040 1.390 ;
        RECT 13.930 0.445 16.040 0.615 ;
        RECT 13.930 0.170 14.100 0.445 ;
        RECT 14.415 0.170 14.585 0.445 ;
        RECT 14.900 0.170 15.070 0.445 ;
        RECT 15.385 0.170 15.555 0.445 ;
        RECT 15.870 0.170 16.040 0.445 ;
        RECT 16.480 0.170 16.820 2.720 ;
        RECT 17.260 0.615 17.430 1.745 ;
        RECT 18.230 0.615 18.400 1.390 ;
        RECT 19.200 0.615 19.370 1.390 ;
        RECT 17.260 0.445 19.370 0.615 ;
        RECT 17.260 0.170 17.430 0.445 ;
        RECT 17.745 0.170 17.915 0.445 ;
        RECT 18.230 0.170 18.400 0.445 ;
        RECT 18.715 0.170 18.885 0.445 ;
        RECT 19.200 0.170 19.370 0.445 ;
        RECT 19.810 0.170 20.150 2.720 ;
        RECT -0.170 -0.170 20.150 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 20.150 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 3.365 5.285 3.535 7.020 ;
        RECT 4.245 5.285 4.415 7.020 ;
        RECT 3.365 5.115 4.895 5.285 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 2.830 1.665 3.000 1.745 ;
        RECT 3.800 1.665 3.970 1.745 ;
        RECT 4.725 1.740 4.895 5.115 ;
        RECT 6.205 1.920 6.375 4.865 ;
        RECT 6.580 4.665 6.750 7.020 ;
        RECT 8.915 5.285 9.085 7.020 ;
        RECT 9.795 5.285 9.965 7.020 ;
        RECT 8.915 5.115 10.445 5.285 ;
        RECT 6.580 4.495 7.115 4.665 ;
        RECT 6.945 2.165 7.115 4.495 ;
        RECT 6.575 1.995 7.115 2.165 ;
        RECT 2.830 1.495 3.970 1.665 ;
        RECT 2.830 0.365 3.000 1.495 ;
        RECT 3.800 0.615 3.970 1.495 ;
        RECT 4.285 1.570 4.895 1.740 ;
        RECT 4.285 0.835 4.455 1.570 ;
        RECT 4.770 0.615 4.940 1.385 ;
        RECT 6.575 0.840 6.745 1.995 ;
        RECT 8.380 1.665 8.550 1.745 ;
        RECT 9.350 1.665 9.520 1.745 ;
        RECT 10.275 1.740 10.445 5.115 ;
        RECT 11.755 1.920 11.925 4.865 ;
        RECT 12.130 4.665 12.300 7.020 ;
        RECT 14.025 5.295 14.195 7.025 ;
        RECT 14.905 6.825 15.955 6.995 ;
        RECT 14.905 5.295 15.075 6.825 ;
        RECT 15.785 5.555 15.955 6.825 ;
        RECT 14.025 5.125 15.075 5.295 ;
        RECT 17.355 5.295 17.525 7.025 ;
        RECT 18.235 6.825 19.285 6.995 ;
        RECT 18.235 5.295 18.405 6.825 ;
        RECT 17.355 5.125 18.405 5.295 ;
        RECT 18.675 5.295 18.845 6.565 ;
        RECT 19.115 5.555 19.285 6.825 ;
        RECT 18.675 5.125 19.325 5.295 ;
        RECT 14.190 4.710 14.360 4.870 ;
        RECT 15.120 4.710 15.290 4.870 ;
        RECT 18.450 4.710 18.620 4.870 ;
        RECT 12.130 4.495 12.665 4.665 ;
        RECT 14.190 4.540 14.515 4.710 ;
        RECT 12.495 2.165 12.665 4.495 ;
        RECT 12.125 1.995 12.665 2.165 ;
        RECT 8.380 1.495 9.520 1.665 ;
        RECT 3.800 0.445 4.940 0.615 ;
        RECT 3.800 0.365 3.970 0.445 ;
        RECT 4.770 0.365 4.940 0.445 ;
        RECT 8.380 0.365 8.550 1.495 ;
        RECT 9.350 0.615 9.520 1.495 ;
        RECT 9.835 1.570 10.445 1.740 ;
        RECT 9.835 0.835 10.005 1.570 ;
        RECT 10.320 0.615 10.490 1.385 ;
        RECT 12.125 0.840 12.295 1.995 ;
        RECT 14.345 1.915 14.515 4.540 ;
        RECT 15.085 4.540 15.290 4.710 ;
        RECT 18.415 4.540 18.620 4.710 ;
        RECT 15.085 1.915 15.255 4.540 ;
        RECT 18.415 1.915 18.585 4.540 ;
        RECT 19.155 1.740 19.325 5.125 ;
        RECT 17.745 1.570 19.325 1.740 ;
        RECT 17.745 0.835 17.915 1.570 ;
        RECT 18.715 0.835 18.885 1.570 ;
        RECT 9.350 0.445 10.490 0.615 ;
        RECT 9.350 0.365 9.520 0.445 ;
        RECT 10.320 0.365 10.490 0.445 ;
      LAYER mcon ;
        RECT 1.395 3.615 1.565 3.785 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 4.725 3.245 4.895 3.415 ;
        RECT 6.205 3.245 6.375 3.415 ;
        RECT 6.945 3.615 7.115 3.785 ;
        RECT 10.275 3.245 10.445 3.415 ;
        RECT 11.755 3.245 11.925 3.415 ;
        RECT 12.495 3.985 12.665 4.155 ;
        RECT 14.345 3.615 14.515 3.785 ;
        RECT 15.085 3.615 15.255 3.785 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 19.155 3.615 19.325 3.785 ;
      LAYER met1 ;
        RECT 12.465 4.155 12.695 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 12.435 3.985 18.645 4.155 ;
        RECT 12.465 3.955 12.695 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 1.365 3.785 1.595 3.815 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 6.915 3.785 7.145 3.815 ;
        RECT 14.315 3.785 14.545 3.815 ;
        RECT 15.055 3.785 15.285 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 1.335 3.615 3.475 3.785 ;
        RECT 6.885 3.615 14.575 3.785 ;
        RECT 15.025 3.615 19.385 3.785 ;
        RECT 1.365 3.585 1.595 3.615 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 6.915 3.585 7.145 3.615 ;
        RECT 14.315 3.585 14.545 3.615 ;
        RECT 15.055 3.585 15.285 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
        RECT 4.695 3.415 4.925 3.445 ;
        RECT 6.175 3.415 6.405 3.445 ;
        RECT 10.245 3.415 10.475 3.445 ;
        RECT 11.725 3.415 11.955 3.445 ;
        RECT 4.665 3.245 6.435 3.415 ;
        RECT 10.215 3.245 11.985 3.415 ;
        RECT 4.695 3.215 4.925 3.245 ;
        RECT 6.175 3.215 6.405 3.245 ;
        RECT 10.245 3.215 10.475 3.245 ;
        RECT 11.725 3.215 11.955 3.245 ;
  END
END DLATCH






MACRO DLATCHN
  CLASS CORE ;
  FOREIGN DLATCHN ;
  ORIGIN 0.000 0.000 ;
  SIZE 22.200 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 0.963050 ;
    PORT
      LAYER li1 ;
        RECT 17.565 5.295 17.735 6.565 ;
        RECT 17.565 5.125 18.215 5.295 ;
        RECT 18.045 1.740 18.215 5.125 ;
        RECT 19.740 4.710 19.910 4.870 ;
        RECT 19.740 4.540 20.065 4.710 ;
        RECT 19.895 1.915 20.065 4.540 ;
        RECT 16.635 1.570 18.215 1.740 ;
        RECT 16.635 0.835 16.805 1.570 ;
        RECT 17.605 0.835 17.775 1.570 ;
      LAYER mcon ;
        RECT 18.045 3.245 18.215 3.415 ;
        RECT 19.895 3.245 20.065 3.415 ;
      LAYER met1 ;
        RECT 18.015 3.415 18.245 3.445 ;
        RECT 19.865 3.415 20.095 3.445 ;
        RECT 17.985 3.245 20.125 3.415 ;
        RECT 18.015 3.215 18.245 3.245 ;
        RECT 19.865 3.215 20.095 3.245 ;
    END
  END Q
  PIN D
    ANTENNAGATEAREA 2.054500 ;
    PORT
      LAYER li1 ;
        RECT 2.875 1.920 3.045 4.865 ;
        RECT 11.785 4.710 11.955 4.865 ;
        RECT 11.755 4.535 11.955 4.710 ;
        RECT 11.755 1.915 11.925 4.535 ;
      LAYER mcon ;
        RECT 2.875 3.985 3.045 4.155 ;
        RECT 11.755 3.985 11.925 4.155 ;
      LAYER met1 ;
        RECT 2.845 4.155 3.075 4.185 ;
        RECT 11.725 4.155 11.955 4.185 ;
        RECT 2.815 3.985 11.985 4.155 ;
        RECT 2.845 3.955 3.075 3.985 ;
        RECT 11.725 3.955 11.955 3.985 ;
    END
  END D
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 22.635 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 22.370 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
        RECT 2.810 5.185 2.980 7.230 ;
        RECT 3.690 5.185 3.860 7.230 ;
        RECT 4.270 4.110 4.610 7.230 ;
        RECT 5.145 5.135 5.315 7.230 ;
        RECT 6.025 5.555 6.195 7.230 ;
        RECT 6.905 5.555 7.075 7.230 ;
        RECT 7.600 4.110 7.940 7.230 ;
        RECT 8.360 5.185 8.530 7.230 ;
        RECT 9.240 5.185 9.410 7.230 ;
        RECT 9.820 4.110 10.160 7.230 ;
        RECT 10.695 5.135 10.865 7.230 ;
        RECT 11.575 5.555 11.745 7.230 ;
        RECT 12.455 5.555 12.625 7.230 ;
        RECT 13.150 4.110 13.490 7.230 ;
        RECT 13.910 5.185 14.080 7.230 ;
        RECT 14.790 5.185 14.960 7.230 ;
        RECT 15.370 4.110 15.710 7.230 ;
        RECT 16.685 5.555 16.855 7.230 ;
        RECT 18.700 4.110 19.040 7.230 ;
        RECT 20.015 5.555 20.185 7.230 ;
        RECT 22.030 4.110 22.370 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 22.370 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 22.370 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT 2.765 0.620 2.935 1.750 ;
        RECT 3.735 0.620 3.905 1.750 ;
        RECT 2.765 0.450 3.905 0.620 ;
        RECT 2.765 0.170 2.935 0.450 ;
        RECT 3.250 0.170 3.420 0.450 ;
        RECT 3.735 0.170 3.905 0.450 ;
        RECT 4.270 0.170 4.610 2.720 ;
        RECT 5.535 0.170 5.705 1.120 ;
        RECT 7.600 0.170 7.940 2.720 ;
        RECT 8.315 0.620 8.485 1.750 ;
        RECT 9.285 0.620 9.455 1.750 ;
        RECT 8.315 0.450 9.455 0.620 ;
        RECT 8.315 0.170 8.485 0.450 ;
        RECT 8.800 0.170 8.970 0.450 ;
        RECT 9.285 0.170 9.455 0.450 ;
        RECT 9.820 0.170 10.160 2.720 ;
        RECT 11.085 0.170 11.255 1.120 ;
        RECT 13.150 0.170 13.490 2.720 ;
        RECT 13.865 0.620 14.035 1.750 ;
        RECT 14.835 0.620 15.005 1.750 ;
        RECT 13.865 0.450 15.005 0.620 ;
        RECT 13.865 0.170 14.035 0.450 ;
        RECT 14.350 0.170 14.520 0.450 ;
        RECT 14.835 0.170 15.005 0.450 ;
        RECT 15.370 0.170 15.710 2.720 ;
        RECT 16.150 0.615 16.320 1.745 ;
        RECT 17.120 0.615 17.290 1.390 ;
        RECT 18.090 0.615 18.260 1.390 ;
        RECT 16.150 0.445 18.260 0.615 ;
        RECT 16.150 0.170 16.320 0.445 ;
        RECT 16.635 0.170 16.805 0.445 ;
        RECT 17.120 0.170 17.290 0.445 ;
        RECT 17.605 0.170 17.775 0.445 ;
        RECT 18.090 0.170 18.260 0.445 ;
        RECT 18.700 0.170 19.040 2.720 ;
        RECT 19.480 0.615 19.650 1.745 ;
        RECT 20.450 0.615 20.620 1.390 ;
        RECT 21.420 0.615 21.590 1.390 ;
        RECT 19.480 0.445 21.590 0.615 ;
        RECT 19.480 0.170 19.650 0.445 ;
        RECT 19.965 0.170 20.135 0.445 ;
        RECT 20.450 0.170 20.620 0.445 ;
        RECT 20.935 0.170 21.105 0.445 ;
        RECT 21.420 0.170 21.590 0.445 ;
        RECT 22.030 0.170 22.370 2.720 ;
        RECT -0.170 -0.170 22.370 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 22.370 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 3.250 4.665 3.420 7.020 ;
        RECT 5.585 5.285 5.755 7.020 ;
        RECT 6.465 5.285 6.635 7.020 ;
        RECT 5.585 5.115 7.115 5.285 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 3.250 4.495 3.785 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 3.615 2.165 3.785 4.495 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 3.245 1.995 3.785 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
        RECT 3.245 0.840 3.415 1.995 ;
        RECT 5.465 1.915 5.635 4.865 ;
        RECT 6.235 4.710 6.405 4.865 ;
        RECT 6.205 4.535 6.405 4.710 ;
        RECT 6.205 1.915 6.375 4.535 ;
        RECT 5.050 1.665 5.220 1.745 ;
        RECT 6.020 1.665 6.190 1.745 ;
        RECT 6.945 1.740 7.115 5.115 ;
        RECT 8.425 1.920 8.595 4.865 ;
        RECT 8.800 4.665 8.970 7.020 ;
        RECT 11.135 5.285 11.305 7.020 ;
        RECT 12.015 5.285 12.185 7.020 ;
        RECT 11.135 5.115 12.665 5.285 ;
        RECT 8.800 4.495 9.335 4.665 ;
        RECT 9.165 2.165 9.335 4.495 ;
        RECT 8.795 1.995 9.335 2.165 ;
        RECT 5.050 1.495 6.190 1.665 ;
        RECT 5.050 0.365 5.220 1.495 ;
        RECT 6.020 0.615 6.190 1.495 ;
        RECT 6.505 1.570 7.115 1.740 ;
        RECT 6.505 0.835 6.675 1.570 ;
        RECT 6.990 0.615 7.160 1.385 ;
        RECT 8.795 0.840 8.965 1.995 ;
        RECT 11.015 1.915 11.185 4.865 ;
        RECT 10.600 1.665 10.770 1.745 ;
        RECT 11.570 1.665 11.740 1.745 ;
        RECT 12.495 1.740 12.665 5.115 ;
        RECT 13.975 1.920 14.145 4.865 ;
        RECT 14.350 4.665 14.520 7.020 ;
        RECT 16.245 5.295 16.415 7.025 ;
        RECT 17.125 6.825 18.175 6.995 ;
        RECT 17.125 5.295 17.295 6.825 ;
        RECT 18.005 5.555 18.175 6.825 ;
        RECT 16.245 5.125 17.295 5.295 ;
        RECT 19.575 5.295 19.745 7.025 ;
        RECT 20.455 6.825 21.505 6.995 ;
        RECT 20.455 5.295 20.625 6.825 ;
        RECT 19.575 5.125 20.625 5.295 ;
        RECT 20.895 5.295 21.065 6.565 ;
        RECT 21.335 5.555 21.505 6.825 ;
        RECT 20.895 5.125 21.545 5.295 ;
        RECT 16.410 4.710 16.580 4.870 ;
        RECT 17.340 4.710 17.510 4.870 ;
        RECT 20.670 4.710 20.840 4.870 ;
        RECT 14.350 4.495 14.885 4.665 ;
        RECT 16.410 4.540 16.735 4.710 ;
        RECT 14.715 2.165 14.885 4.495 ;
        RECT 14.345 1.995 14.885 2.165 ;
        RECT 10.600 1.495 11.740 1.665 ;
        RECT 6.020 0.445 7.160 0.615 ;
        RECT 6.020 0.365 6.190 0.445 ;
        RECT 6.990 0.365 7.160 0.445 ;
        RECT 10.600 0.365 10.770 1.495 ;
        RECT 11.570 0.615 11.740 1.495 ;
        RECT 12.055 1.570 12.665 1.740 ;
        RECT 12.055 0.835 12.225 1.570 ;
        RECT 12.540 0.615 12.710 1.385 ;
        RECT 14.345 0.840 14.515 1.995 ;
        RECT 16.565 1.915 16.735 4.540 ;
        RECT 17.305 4.540 17.510 4.710 ;
        RECT 20.635 4.540 20.840 4.710 ;
        RECT 17.305 1.915 17.475 4.540 ;
        RECT 20.635 1.915 20.805 4.540 ;
        RECT 21.375 1.740 21.545 5.125 ;
        RECT 19.965 1.570 21.545 1.740 ;
        RECT 19.965 0.835 20.135 1.570 ;
        RECT 20.935 0.835 21.105 1.570 ;
        RECT 11.570 0.445 12.710 0.615 ;
        RECT 11.570 0.365 11.740 0.445 ;
        RECT 12.540 0.365 12.710 0.445 ;
      LAYER mcon ;
        RECT 1.395 2.875 1.565 3.045 ;
        RECT 3.615 3.615 3.785 3.785 ;
        RECT 5.465 3.615 5.635 3.785 ;
        RECT 6.205 2.875 6.375 3.045 ;
        RECT 6.945 3.245 7.115 3.415 ;
        RECT 8.425 3.245 8.595 3.415 ;
        RECT 9.165 3.615 9.335 3.785 ;
        RECT 11.015 2.875 11.185 3.045 ;
        RECT 12.495 3.245 12.665 3.415 ;
        RECT 13.975 3.245 14.145 3.415 ;
        RECT 14.715 3.985 14.885 4.155 ;
        RECT 16.565 3.615 16.735 3.785 ;
        RECT 17.305 3.615 17.475 3.785 ;
        RECT 20.635 3.985 20.805 4.155 ;
        RECT 21.375 3.615 21.545 3.785 ;
      LAYER met1 ;
        RECT 14.685 4.155 14.915 4.185 ;
        RECT 20.605 4.155 20.835 4.185 ;
        RECT 14.655 3.985 20.865 4.155 ;
        RECT 14.685 3.955 14.915 3.985 ;
        RECT 20.605 3.955 20.835 3.985 ;
        RECT 3.585 3.785 3.815 3.815 ;
        RECT 5.435 3.785 5.665 3.815 ;
        RECT 9.135 3.785 9.365 3.815 ;
        RECT 16.535 3.785 16.765 3.815 ;
        RECT 17.275 3.785 17.505 3.815 ;
        RECT 21.345 3.785 21.575 3.815 ;
        RECT 3.555 3.615 5.695 3.785 ;
        RECT 9.105 3.615 16.795 3.785 ;
        RECT 17.245 3.615 21.605 3.785 ;
        RECT 3.585 3.585 3.815 3.615 ;
        RECT 5.435 3.585 5.665 3.615 ;
        RECT 9.135 3.585 9.365 3.615 ;
        RECT 16.535 3.585 16.765 3.615 ;
        RECT 17.275 3.585 17.505 3.615 ;
        RECT 21.345 3.585 21.575 3.615 ;
        RECT 6.915 3.415 7.145 3.445 ;
        RECT 8.395 3.415 8.625 3.445 ;
        RECT 12.465 3.415 12.695 3.445 ;
        RECT 13.945 3.415 14.175 3.445 ;
        RECT 6.885 3.245 8.655 3.415 ;
        RECT 12.435 3.245 14.205 3.415 ;
        RECT 6.915 3.215 7.145 3.245 ;
        RECT 8.395 3.215 8.625 3.245 ;
        RECT 12.465 3.215 12.695 3.245 ;
        RECT 13.945 3.215 14.175 3.245 ;
        RECT 1.365 3.045 1.595 3.075 ;
        RECT 6.175 3.045 6.405 3.075 ;
        RECT 10.985 3.045 11.215 3.075 ;
        RECT 1.335 2.875 11.245 3.045 ;
        RECT 1.365 2.845 1.595 2.875 ;
        RECT 6.175 2.845 6.405 2.875 ;
        RECT 10.985 2.845 11.215 2.875 ;
  END
END DLATCHN






MACRO FA
  CLASS CORE ;
  FOREIGN FA ;
  ORIGIN 0.000 0.000 ;
  SIZE 38.850 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN SUM
    ANTENNADIFFAREA 1.543800 ;
    PORT
      LAYER li1 ;
        RECT 15.345 5.290 15.515 6.560 ;
        RECT 18.675 5.290 18.845 6.560 ;
        RECT 15.345 5.120 15.995 5.290 ;
        RECT 18.675 5.120 19.325 5.290 ;
        RECT 15.825 1.740 15.995 5.120 ;
        RECT 19.155 1.740 19.325 5.120 ;
        RECT 15.385 1.570 15.995 1.740 ;
        RECT 18.715 1.570 19.325 1.740 ;
        RECT 15.385 0.840 15.555 1.570 ;
        RECT 18.715 0.840 18.885 1.570 ;
      LAYER mcon ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 19.155 3.615 19.325 3.785 ;
      LAYER met1 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 15.765 3.615 19.385 3.785 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
    END
  END SUM
  PIN A
    ANTENNAGATEAREA 3.087750 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 3.245 2.305 3.415 4.865 ;
        RECT 29.545 4.710 29.715 4.865 ;
        RECT 29.515 4.535 29.715 4.710 ;
        RECT 29.515 2.305 29.685 4.535 ;
        RECT 3.165 2.135 3.495 2.305 ;
        RECT 29.435 2.135 29.765 2.305 ;
        RECT 3.245 1.920 3.415 2.135 ;
        RECT 29.515 1.915 29.685 2.135 ;
      LAYER mcon ;
        RECT 0.655 3.985 0.825 4.155 ;
        RECT 3.245 3.985 3.415 4.155 ;
        RECT 3.245 2.135 3.415 2.305 ;
        RECT 29.515 2.135 29.685 2.305 ;
      LAYER met1 ;
        RECT 0.625 4.155 0.855 4.185 ;
        RECT 3.215 4.155 3.445 4.185 ;
        RECT 0.595 3.985 3.475 4.155 ;
        RECT 0.625 3.955 0.855 3.985 ;
        RECT 3.215 3.955 3.445 3.985 ;
        RECT 3.245 2.335 3.415 2.365 ;
        RECT 29.515 2.335 29.685 2.365 ;
        RECT 3.215 2.105 3.445 2.335 ;
        RECT 29.485 2.105 29.715 2.335 ;
        RECT 3.245 1.935 3.415 2.105 ;
        RECT 29.515 1.935 29.685 2.105 ;
        RECT 3.245 1.765 29.685 1.935 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 3.087750 ;
    PORT
      LAYER li1 ;
        RECT 6.575 4.275 6.745 4.865 ;
        RECT 4.355 1.920 4.525 3.125 ;
        RECT 10.275 1.920 10.445 4.975 ;
        RECT 28.775 4.715 28.945 4.895 ;
        RECT 28.695 4.545 29.025 4.715 ;
        RECT 28.775 1.915 28.945 4.545 ;
      LAYER mcon ;
        RECT 6.575 4.355 6.745 4.525 ;
        RECT 10.275 4.725 10.445 4.895 ;
        RECT 28.775 4.545 28.945 4.715 ;
        RECT 10.275 4.355 10.445 4.525 ;
        RECT 4.355 2.875 4.525 3.045 ;
        RECT 10.275 2.875 10.445 3.045 ;
      LAYER met1 ;
        RECT 10.245 4.895 10.475 4.925 ;
        RECT 10.215 4.745 28.945 4.895 ;
        RECT 10.215 4.725 28.975 4.745 ;
        RECT 10.245 4.695 10.475 4.725 ;
        RECT 6.545 4.525 6.775 4.555 ;
        RECT 10.245 4.525 10.475 4.555 ;
        RECT 6.515 4.355 10.505 4.525 ;
        RECT 28.745 4.515 28.975 4.725 ;
        RECT 28.775 4.485 28.945 4.515 ;
        RECT 6.545 4.325 6.775 4.355 ;
        RECT 10.245 4.325 10.475 4.355 ;
        RECT 4.325 3.045 4.555 3.075 ;
        RECT 10.245 3.045 10.475 3.075 ;
        RECT 4.295 2.875 10.505 3.045 ;
        RECT 4.325 2.845 4.555 2.875 ;
        RECT 10.245 2.845 10.475 2.875 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA 3.087750 ;
    PORT
      LAYER li1 ;
        RECT 17.675 4.275 17.845 4.865 ;
        RECT 15.455 1.920 15.625 3.125 ;
        RECT 21.375 1.920 21.545 4.865 ;
        RECT 23.225 1.915 23.395 4.865 ;
      LAYER mcon ;
        RECT 17.675 4.355 17.845 4.525 ;
        RECT 21.375 4.355 21.545 4.525 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 21.375 2.875 21.545 3.045 ;
        RECT 23.225 4.355 23.395 4.525 ;
      LAYER met1 ;
        RECT 17.645 4.525 17.875 4.555 ;
        RECT 21.345 4.525 21.575 4.555 ;
        RECT 23.195 4.525 23.425 4.555 ;
        RECT 17.615 4.355 23.455 4.525 ;
        RECT 17.645 4.325 17.875 4.355 ;
        RECT 21.345 4.325 21.575 4.355 ;
        RECT 23.195 4.325 23.425 4.355 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 21.345 3.045 21.575 3.075 ;
        RECT 15.395 2.875 21.605 3.045 ;
        RECT 15.425 2.845 15.655 2.875 ;
        RECT 21.345 2.845 21.575 2.875 ;
    END
  END CIN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 39.285 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 39.020 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
        RECT 3.365 5.550 3.535 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
        RECT 6.695 5.550 6.865 7.230 ;
        RECT 8.710 4.110 9.050 7.230 ;
        RECT 9.460 5.185 9.630 7.230 ;
        RECT 10.340 5.185 10.510 7.230 ;
        RECT 10.930 4.110 11.270 7.230 ;
        RECT 11.690 5.185 11.860 7.230 ;
        RECT 12.570 5.185 12.740 7.230 ;
        RECT 13.150 4.110 13.490 7.230 ;
        RECT 14.465 5.550 14.635 7.230 ;
        RECT 16.480 4.110 16.820 7.230 ;
        RECT 17.795 5.550 17.965 7.230 ;
        RECT 19.810 4.110 20.150 7.230 ;
        RECT 20.560 5.185 20.730 7.230 ;
        RECT 21.440 5.185 21.610 7.230 ;
        RECT 22.030 4.110 22.370 7.230 ;
        RECT 22.905 5.135 23.075 7.230 ;
        RECT 23.785 5.555 23.955 7.230 ;
        RECT 24.665 5.555 24.835 7.230 ;
        RECT 25.360 4.110 25.700 7.230 ;
        RECT 26.120 5.185 26.290 7.230 ;
        RECT 27.000 5.185 27.170 7.230 ;
        RECT 27.580 4.110 27.920 7.230 ;
        RECT 28.455 5.135 28.625 7.230 ;
        RECT 29.335 5.555 29.505 7.230 ;
        RECT 30.215 5.555 30.385 7.230 ;
        RECT 30.910 4.110 31.250 7.230 ;
        RECT 31.670 5.185 31.840 7.230 ;
        RECT 32.550 5.185 32.720 7.230 ;
        RECT 33.130 4.110 33.470 7.230 ;
        RECT 34.445 5.555 34.615 7.230 ;
        RECT 36.460 4.110 36.800 7.230 ;
        RECT 37.220 5.185 37.390 7.230 ;
        RECT 38.100 5.185 38.270 7.230 ;
        RECT 38.680 4.110 39.020 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.515 7.315 29.685 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.625 7.315 30.795 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 32.845 7.315 33.015 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.435 7.315 35.605 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.175 7.315 36.345 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 39.020 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 39.020 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT 3.315 0.170 3.485 1.125 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT 6.645 0.170 6.815 1.125 ;
        RECT 8.710 0.170 9.050 2.720 ;
        RECT 9.415 0.620 9.585 1.750 ;
        RECT 10.385 0.620 10.555 1.750 ;
        RECT 9.415 0.450 10.555 0.620 ;
        RECT 9.415 0.170 9.585 0.450 ;
        RECT 9.900 0.170 10.070 0.450 ;
        RECT 10.385 0.170 10.555 0.450 ;
        RECT 10.930 0.170 11.270 2.720 ;
        RECT 11.645 0.620 11.815 1.750 ;
        RECT 12.615 0.620 12.785 1.750 ;
        RECT 11.645 0.450 12.785 0.620 ;
        RECT 11.645 0.170 11.815 0.450 ;
        RECT 12.130 0.170 12.300 0.450 ;
        RECT 12.615 0.170 12.785 0.450 ;
        RECT 13.150 0.170 13.490 2.720 ;
        RECT 14.415 0.170 14.585 1.125 ;
        RECT 16.480 0.170 16.820 2.720 ;
        RECT 17.745 0.170 17.915 1.125 ;
        RECT 19.810 0.170 20.150 2.720 ;
        RECT 20.515 0.620 20.685 1.750 ;
        RECT 21.485 0.620 21.655 1.750 ;
        RECT 20.515 0.450 21.655 0.620 ;
        RECT 20.515 0.170 20.685 0.450 ;
        RECT 21.000 0.170 21.170 0.450 ;
        RECT 21.485 0.170 21.655 0.450 ;
        RECT 22.030 0.170 22.370 2.720 ;
        RECT 23.295 0.170 23.465 1.120 ;
        RECT 25.360 0.170 25.700 2.720 ;
        RECT 26.075 0.620 26.245 1.750 ;
        RECT 27.045 0.620 27.215 1.750 ;
        RECT 26.075 0.450 27.215 0.620 ;
        RECT 26.075 0.170 26.245 0.450 ;
        RECT 26.560 0.170 26.730 0.450 ;
        RECT 27.045 0.170 27.215 0.450 ;
        RECT 27.580 0.170 27.920 2.720 ;
        RECT 28.845 0.170 29.015 1.120 ;
        RECT 30.910 0.170 31.250 2.720 ;
        RECT 31.625 0.620 31.795 1.750 ;
        RECT 32.595 0.620 32.765 1.750 ;
        RECT 31.625 0.450 32.765 0.620 ;
        RECT 31.625 0.170 31.795 0.450 ;
        RECT 32.110 0.170 32.280 0.450 ;
        RECT 32.595 0.170 32.765 0.450 ;
        RECT 33.130 0.170 33.470 2.720 ;
        RECT 33.910 0.615 34.080 1.745 ;
        RECT 34.880 0.615 35.050 1.390 ;
        RECT 35.850 0.615 36.020 1.390 ;
        RECT 33.910 0.445 36.020 0.615 ;
        RECT 33.910 0.170 34.080 0.445 ;
        RECT 34.395 0.170 34.565 0.445 ;
        RECT 34.880 0.170 35.050 0.445 ;
        RECT 35.365 0.170 35.535 0.445 ;
        RECT 35.850 0.170 36.020 0.445 ;
        RECT 36.460 0.170 36.800 2.720 ;
        RECT 37.175 0.620 37.345 1.750 ;
        RECT 38.145 0.620 38.315 1.750 ;
        RECT 37.175 0.450 38.315 0.620 ;
        RECT 37.175 0.170 37.345 0.450 ;
        RECT 37.660 0.170 37.830 0.450 ;
        RECT 38.145 0.170 38.315 0.450 ;
        RECT 38.680 0.170 39.020 2.720 ;
        RECT -0.170 -0.170 39.020 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.515 -0.085 29.685 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.625 -0.085 30.795 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 32.845 -0.085 33.015 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.435 -0.085 35.605 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.175 -0.085 36.345 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 39.020 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 2.925 5.290 3.095 6.900 ;
        RECT 3.805 6.820 4.855 6.990 ;
        RECT 3.805 5.290 3.975 6.820 ;
        RECT 2.925 5.120 3.975 5.290 ;
        RECT 4.245 5.290 4.415 6.560 ;
        RECT 4.685 5.550 4.855 6.820 ;
        RECT 6.255 5.290 6.425 6.900 ;
        RECT 7.135 6.820 8.185 6.990 ;
        RECT 7.135 5.290 7.305 6.820 ;
        RECT 4.245 5.120 4.895 5.290 ;
        RECT 6.255 5.120 7.305 5.290 ;
        RECT 7.575 5.290 7.745 6.560 ;
        RECT 8.015 5.550 8.185 6.820 ;
        RECT 7.575 5.120 8.225 5.290 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 4.355 3.905 4.525 4.865 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
        RECT 2.830 1.670 3.000 1.750 ;
        RECT 3.800 1.670 3.970 1.750 ;
        RECT 4.725 1.740 4.895 5.120 ;
        RECT 6.575 1.920 6.745 3.495 ;
        RECT 7.685 1.920 7.855 4.865 ;
        RECT 2.830 1.500 3.970 1.670 ;
        RECT 2.830 0.370 3.000 1.500 ;
        RECT 3.800 0.620 3.970 1.500 ;
        RECT 4.285 1.570 4.895 1.740 ;
        RECT 6.160 1.670 6.330 1.750 ;
        RECT 7.130 1.670 7.300 1.750 ;
        RECT 8.055 1.740 8.225 5.120 ;
        RECT 9.900 4.665 10.070 7.020 ;
        RECT 9.535 4.495 10.070 4.665 ;
        RECT 9.535 2.165 9.705 4.495 ;
        RECT 9.535 1.995 10.075 2.165 ;
        RECT 4.285 0.840 4.455 1.570 ;
        RECT 6.160 1.500 7.300 1.670 ;
        RECT 4.770 0.620 4.940 1.390 ;
        RECT 3.800 0.450 4.940 0.620 ;
        RECT 3.800 0.370 3.970 0.450 ;
        RECT 4.770 0.370 4.940 0.450 ;
        RECT 6.160 0.370 6.330 1.500 ;
        RECT 7.130 0.620 7.300 1.500 ;
        RECT 7.615 1.570 8.225 1.740 ;
        RECT 7.615 0.840 7.785 1.570 ;
        RECT 8.100 0.620 8.270 1.390 ;
        RECT 9.905 0.840 10.075 1.995 ;
        RECT 11.755 1.920 11.925 4.865 ;
        RECT 12.130 4.665 12.300 7.020 ;
        RECT 14.025 5.290 14.195 6.900 ;
        RECT 14.905 6.820 15.955 6.990 ;
        RECT 14.905 5.290 15.075 6.820 ;
        RECT 15.785 5.550 15.955 6.820 ;
        RECT 14.025 5.120 15.075 5.290 ;
        RECT 17.355 5.290 17.525 6.900 ;
        RECT 18.235 6.820 19.285 6.990 ;
        RECT 18.235 5.290 18.405 6.820 ;
        RECT 19.115 5.550 19.285 6.820 ;
        RECT 17.355 5.120 18.405 5.290 ;
        RECT 12.130 4.495 12.665 4.665 ;
        RECT 12.495 2.165 12.665 4.495 ;
        RECT 12.125 1.995 12.665 2.165 ;
        RECT 12.125 0.840 12.295 1.995 ;
        RECT 14.345 1.920 14.515 4.865 ;
        RECT 15.455 3.905 15.625 4.865 ;
        RECT 17.675 1.920 17.845 3.495 ;
        RECT 18.785 1.920 18.955 4.865 ;
        RECT 21.000 4.665 21.170 7.020 ;
        RECT 23.345 5.285 23.515 7.020 ;
        RECT 24.225 5.285 24.395 7.020 ;
        RECT 23.345 5.115 24.875 5.285 ;
        RECT 23.995 4.710 24.165 4.865 ;
        RECT 20.635 4.495 21.170 4.665 ;
        RECT 23.965 4.535 24.165 4.710 ;
        RECT 20.635 2.165 20.805 4.495 ;
        RECT 20.635 1.995 21.175 2.165 ;
        RECT 13.930 1.670 14.100 1.750 ;
        RECT 14.900 1.670 15.070 1.750 ;
        RECT 13.930 1.500 15.070 1.670 ;
        RECT 7.130 0.450 8.270 0.620 ;
        RECT 7.130 0.370 7.300 0.450 ;
        RECT 8.100 0.370 8.270 0.450 ;
        RECT 13.930 0.370 14.100 1.500 ;
        RECT 14.900 0.620 15.070 1.500 ;
        RECT 17.260 1.670 17.430 1.750 ;
        RECT 18.230 1.670 18.400 1.750 ;
        RECT 17.260 1.500 18.400 1.670 ;
        RECT 15.870 0.620 16.040 1.390 ;
        RECT 14.900 0.450 16.040 0.620 ;
        RECT 14.900 0.370 15.070 0.450 ;
        RECT 15.870 0.370 16.040 0.450 ;
        RECT 17.260 0.370 17.430 1.500 ;
        RECT 18.230 0.620 18.400 1.500 ;
        RECT 19.200 0.620 19.370 1.390 ;
        RECT 21.005 0.840 21.175 1.995 ;
        RECT 23.965 1.915 24.135 4.535 ;
        RECT 22.810 1.665 22.980 1.745 ;
        RECT 23.780 1.665 23.950 1.745 ;
        RECT 24.705 1.740 24.875 5.115 ;
        RECT 26.185 1.920 26.355 4.865 ;
        RECT 26.560 4.665 26.730 7.020 ;
        RECT 28.895 5.285 29.065 7.020 ;
        RECT 29.775 5.285 29.945 7.020 ;
        RECT 28.895 5.115 30.425 5.285 ;
        RECT 26.560 4.495 27.095 4.665 ;
        RECT 26.925 2.165 27.095 4.495 ;
        RECT 26.555 1.995 27.095 2.165 ;
        RECT 22.810 1.495 23.950 1.665 ;
        RECT 18.230 0.450 19.370 0.620 ;
        RECT 18.230 0.370 18.400 0.450 ;
        RECT 19.200 0.370 19.370 0.450 ;
        RECT 22.810 0.365 22.980 1.495 ;
        RECT 23.780 0.615 23.950 1.495 ;
        RECT 24.265 1.570 24.875 1.740 ;
        RECT 24.265 0.835 24.435 1.570 ;
        RECT 24.750 0.615 24.920 1.385 ;
        RECT 26.555 0.840 26.725 1.995 ;
        RECT 28.360 1.665 28.530 1.745 ;
        RECT 29.330 1.665 29.500 1.745 ;
        RECT 30.255 1.740 30.425 5.115 ;
        RECT 31.735 1.920 31.905 4.865 ;
        RECT 32.110 4.665 32.280 7.020 ;
        RECT 34.005 5.295 34.175 7.025 ;
        RECT 34.885 6.825 35.935 6.995 ;
        RECT 34.885 5.295 35.055 6.825 ;
        RECT 34.005 5.125 35.055 5.295 ;
        RECT 35.325 5.295 35.495 6.565 ;
        RECT 35.765 5.555 35.935 6.825 ;
        RECT 35.325 5.125 35.975 5.295 ;
        RECT 34.170 4.710 34.340 4.870 ;
        RECT 35.100 4.710 35.270 4.870 ;
        RECT 32.110 4.495 32.645 4.665 ;
        RECT 34.170 4.540 34.495 4.710 ;
        RECT 32.475 2.165 32.645 4.495 ;
        RECT 32.105 1.995 32.645 2.165 ;
        RECT 28.360 1.495 29.500 1.665 ;
        RECT 23.780 0.445 24.920 0.615 ;
        RECT 23.780 0.365 23.950 0.445 ;
        RECT 24.750 0.365 24.920 0.445 ;
        RECT 28.360 0.365 28.530 1.495 ;
        RECT 29.330 0.615 29.500 1.495 ;
        RECT 29.815 1.570 30.425 1.740 ;
        RECT 29.815 0.835 29.985 1.570 ;
        RECT 30.300 0.615 30.470 1.385 ;
        RECT 32.105 0.840 32.275 1.995 ;
        RECT 34.325 1.915 34.495 4.540 ;
        RECT 35.065 4.540 35.270 4.710 ;
        RECT 35.065 1.915 35.235 4.540 ;
        RECT 35.805 1.740 35.975 5.125 ;
        RECT 37.285 1.920 37.455 4.865 ;
        RECT 37.660 4.665 37.830 7.020 ;
        RECT 37.660 4.495 38.195 4.665 ;
        RECT 38.025 2.165 38.195 4.495 ;
        RECT 37.655 1.995 38.195 2.165 ;
        RECT 34.395 1.570 35.975 1.740 ;
        RECT 34.395 0.835 34.565 1.570 ;
        RECT 35.365 0.835 35.535 1.570 ;
        RECT 37.655 0.840 37.825 1.995 ;
        RECT 29.330 0.445 30.470 0.615 ;
        RECT 29.330 0.365 29.500 0.445 ;
        RECT 30.300 0.365 30.470 0.445 ;
      LAYER mcon ;
        RECT 4.355 3.985 4.525 4.155 ;
        RECT 1.395 2.505 1.565 2.675 ;
        RECT 4.725 3.615 4.895 3.785 ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 7.685 2.505 7.855 2.675 ;
        RECT 8.055 3.615 8.225 3.785 ;
        RECT 9.535 3.985 9.705 4.155 ;
        RECT 9.535 3.245 9.705 3.415 ;
        RECT 11.755 3.985 11.925 4.155 ;
        RECT 11.755 3.615 11.925 3.785 ;
        RECT 11.755 2.135 11.925 2.305 ;
        RECT 12.495 2.505 12.665 2.675 ;
        RECT 14.345 3.985 14.515 4.155 ;
        RECT 15.455 3.985 15.625 4.155 ;
        RECT 17.675 3.245 17.845 3.415 ;
        RECT 18.785 2.505 18.955 2.675 ;
        RECT 20.635 3.985 20.805 4.155 ;
        RECT 20.635 3.245 20.805 3.415 ;
        RECT 23.965 2.135 24.135 2.305 ;
        RECT 24.705 3.245 24.875 3.415 ;
        RECT 26.185 3.245 26.355 3.415 ;
        RECT 26.925 2.875 27.095 3.045 ;
        RECT 30.255 3.245 30.425 3.415 ;
        RECT 31.735 3.245 31.905 3.415 ;
        RECT 32.475 3.245 32.645 3.415 ;
        RECT 34.325 2.875 34.495 3.045 ;
        RECT 35.065 3.245 35.235 3.415 ;
        RECT 35.805 3.245 35.975 3.415 ;
        RECT 37.285 3.245 37.455 3.415 ;
      LAYER met1 ;
        RECT 4.325 4.155 4.555 4.185 ;
        RECT 9.505 4.155 9.735 4.185 ;
        RECT 11.725 4.155 11.955 4.185 ;
        RECT 14.315 4.155 14.545 4.185 ;
        RECT 15.425 4.155 15.655 4.185 ;
        RECT 20.605 4.155 20.835 4.185 ;
        RECT 4.295 3.985 9.765 4.155 ;
        RECT 11.695 3.985 14.575 4.155 ;
        RECT 15.395 3.985 20.865 4.155 ;
        RECT 4.325 3.955 4.555 3.985 ;
        RECT 9.505 3.955 9.735 3.985 ;
        RECT 11.725 3.955 11.955 3.985 ;
        RECT 14.315 3.955 14.545 3.985 ;
        RECT 15.425 3.955 15.655 3.985 ;
        RECT 20.605 3.955 20.835 3.985 ;
        RECT 4.695 3.785 4.925 3.815 ;
        RECT 8.025 3.785 8.255 3.815 ;
        RECT 11.725 3.785 11.955 3.815 ;
        RECT 4.665 3.615 11.985 3.785 ;
        RECT 4.695 3.585 4.925 3.615 ;
        RECT 8.025 3.585 8.255 3.615 ;
        RECT 11.725 3.585 11.955 3.615 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 9.505 3.415 9.735 3.445 ;
        RECT 17.645 3.415 17.875 3.445 ;
        RECT 20.605 3.415 20.835 3.445 ;
        RECT 24.675 3.415 24.905 3.445 ;
        RECT 26.155 3.415 26.385 3.445 ;
        RECT 30.225 3.415 30.455 3.445 ;
        RECT 31.705 3.415 31.935 3.445 ;
        RECT 32.445 3.415 32.675 3.445 ;
        RECT 35.035 3.415 35.265 3.445 ;
        RECT 35.775 3.415 36.005 3.445 ;
        RECT 37.255 3.415 37.485 3.445 ;
        RECT 6.515 3.245 9.765 3.415 ;
        RECT 17.615 3.245 20.865 3.415 ;
        RECT 24.645 3.245 26.415 3.415 ;
        RECT 30.195 3.245 31.965 3.415 ;
        RECT 32.415 3.245 35.295 3.415 ;
        RECT 35.745 3.245 37.515 3.415 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 9.505 3.215 9.735 3.245 ;
        RECT 17.645 3.215 17.875 3.245 ;
        RECT 20.605 3.215 20.835 3.245 ;
        RECT 24.675 3.215 24.905 3.245 ;
        RECT 26.155 3.215 26.385 3.245 ;
        RECT 30.225 3.215 30.455 3.245 ;
        RECT 31.705 3.215 31.935 3.245 ;
        RECT 32.445 3.215 32.675 3.245 ;
        RECT 35.035 3.215 35.265 3.245 ;
        RECT 35.775 3.215 36.005 3.245 ;
        RECT 37.255 3.215 37.485 3.245 ;
        RECT 26.895 3.045 27.125 3.075 ;
        RECT 34.295 3.045 34.525 3.075 ;
        RECT 26.865 2.875 34.555 3.045 ;
        RECT 26.895 2.845 27.125 2.875 ;
        RECT 34.295 2.845 34.525 2.875 ;
        RECT 1.365 2.675 1.595 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 12.465 2.675 12.695 2.705 ;
        RECT 18.755 2.675 18.985 2.705 ;
        RECT 1.335 2.505 7.915 2.675 ;
        RECT 12.435 2.505 19.015 2.675 ;
        RECT 1.365 2.475 1.595 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
        RECT 12.465 2.475 12.695 2.505 ;
        RECT 18.755 2.475 18.985 2.505 ;
        RECT 11.725 2.305 11.955 2.335 ;
        RECT 23.935 2.305 24.165 2.335 ;
        RECT 11.695 2.135 24.195 2.305 ;
        RECT 11.725 2.105 11.955 2.135 ;
        RECT 23.935 2.105 24.165 2.135 ;
  END
END FA






MACRO FILL1
  CLASS CORE SPACER ;
  FOREIGN FILL1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.110 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT -0.170 7.230 1.280 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.170 -0.170 1.280 0.170 ;
    END
  END VGND
  PIN VPB
    ANTENNADIFFAREA 2.787850 ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 1.545 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 1.280 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.940 4.110 1.280 7.230 ;
    END
  END VPB
  PIN VNB
    ANTENNADIFFAREA 2.400250 ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 1.280 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.940 0.170 1.280 2.720 ;
        RECT -0.170 -0.170 1.280 0.170 ;
    END
  END VNB
END FILL1






MACRO HA
  CLASS CORE ;
  FOREIGN HA ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.650 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN SUM
    ANTENNADIFFAREA 1.543800 ;
    PORT
      LAYER li1 ;
        RECT 9.795 5.290 9.965 6.560 ;
        RECT 13.125 5.290 13.295 6.560 ;
        RECT 9.795 5.120 10.445 5.290 ;
        RECT 13.125 5.120 13.775 5.290 ;
        RECT 10.275 1.740 10.445 5.120 ;
        RECT 13.605 1.740 13.775 5.120 ;
        RECT 9.835 1.570 10.445 1.740 ;
        RECT 13.165 1.570 13.775 1.740 ;
        RECT 9.835 0.840 10.005 1.570 ;
        RECT 13.165 0.840 13.335 1.570 ;
      LAYER mcon ;
        RECT 10.275 3.615 10.445 3.785 ;
        RECT 13.605 3.615 13.775 3.785 ;
      LAYER met1 ;
        RECT 10.245 3.785 10.475 3.815 ;
        RECT 13.575 3.785 13.805 3.815 ;
        RECT 10.215 3.615 13.835 3.785 ;
        RECT 10.245 3.585 10.475 3.615 ;
        RECT 13.575 3.585 13.805 3.615 ;
    END
  END SUM
  PIN A
    ANTENNAGATEAREA 3.093750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 6.205 1.920 6.375 4.865 ;
        RECT 8.795 1.920 8.965 4.865 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 6.205 3.985 6.375 4.155 ;
        RECT 8.795 3.985 8.965 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 6.175 4.155 6.405 4.185 ;
        RECT 8.765 4.155 8.995 4.185 ;
        RECT 0.965 3.985 9.025 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 6.175 3.955 6.405 3.985 ;
        RECT 8.765 3.955 8.995 3.985 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 3.081750 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 9.535 3.535 9.705 4.605 ;
        RECT 12.125 4.275 12.295 4.865 ;
        RECT 9.905 1.920 10.075 3.125 ;
        RECT 15.825 1.920 15.995 4.865 ;
      LAYER mcon ;
        RECT 1.765 3.615 1.935 3.785 ;
        RECT 9.535 4.355 9.705 4.525 ;
        RECT 12.125 4.355 12.295 4.525 ;
        RECT 15.825 4.355 15.995 4.525 ;
        RECT 9.535 3.615 9.705 3.785 ;
        RECT 9.905 2.875 10.075 3.045 ;
        RECT 15.825 2.875 15.995 3.045 ;
      LAYER met1 ;
        RECT 9.505 4.525 9.735 4.555 ;
        RECT 12.095 4.525 12.325 4.555 ;
        RECT 15.795 4.525 16.025 4.555 ;
        RECT 9.475 4.355 16.055 4.525 ;
        RECT 9.505 4.325 9.735 4.355 ;
        RECT 12.095 4.325 12.325 4.355 ;
        RECT 15.795 4.325 16.025 4.355 ;
        RECT 1.735 3.785 1.965 3.815 ;
        RECT 9.505 3.785 9.735 3.815 ;
        RECT 1.705 3.615 9.765 3.785 ;
        RECT 1.735 3.585 1.965 3.615 ;
        RECT 9.505 3.585 9.735 3.615 ;
        RECT 9.875 3.045 10.105 3.075 ;
        RECT 15.795 3.045 16.025 3.075 ;
        RECT 9.845 2.875 16.055 3.045 ;
        RECT 9.875 2.845 10.105 2.875 ;
        RECT 15.795 2.845 16.025 2.875 ;
    END
  END B
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 17.085 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 16.820 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 3.920 5.185 4.090 7.230 ;
        RECT 4.800 5.185 4.970 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
        RECT 6.140 5.185 6.310 7.230 ;
        RECT 7.020 5.185 7.190 7.230 ;
        RECT 7.600 4.110 7.940 7.230 ;
        RECT 8.915 5.550 9.085 7.230 ;
        RECT 10.930 4.110 11.270 7.230 ;
        RECT 12.245 5.550 12.415 7.230 ;
        RECT 14.260 4.110 14.600 7.230 ;
        RECT 15.010 5.185 15.180 7.230 ;
        RECT 15.890 5.185 16.060 7.230 ;
        RECT 16.480 4.110 16.820 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 16.820 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 16.820 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 3.875 0.620 4.045 1.750 ;
        RECT 4.845 0.620 5.015 1.750 ;
        RECT 3.875 0.450 5.015 0.620 ;
        RECT 3.875 0.170 4.045 0.450 ;
        RECT 4.360 0.170 4.530 0.450 ;
        RECT 4.845 0.170 5.015 0.450 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT 6.095 0.620 6.265 1.750 ;
        RECT 7.065 0.620 7.235 1.750 ;
        RECT 6.095 0.450 7.235 0.620 ;
        RECT 6.095 0.170 6.265 0.450 ;
        RECT 6.580 0.170 6.750 0.450 ;
        RECT 7.065 0.170 7.235 0.450 ;
        RECT 7.600 0.170 7.940 2.720 ;
        RECT 8.865 0.170 9.035 1.125 ;
        RECT 10.930 0.170 11.270 2.720 ;
        RECT 12.195 0.170 12.365 1.125 ;
        RECT 14.260 0.170 14.600 2.720 ;
        RECT 14.965 0.620 15.135 1.750 ;
        RECT 15.935 0.620 16.105 1.750 ;
        RECT 14.965 0.450 16.105 0.620 ;
        RECT 14.965 0.170 15.135 0.450 ;
        RECT 15.450 0.170 15.620 0.450 ;
        RECT 15.935 0.170 16.105 0.450 ;
        RECT 16.480 0.170 16.820 2.720 ;
        RECT -0.170 -0.170 16.820 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 16.820 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 3.985 1.920 4.155 4.865 ;
        RECT 4.360 4.665 4.530 7.020 ;
        RECT 6.580 4.665 6.750 7.020 ;
        RECT 8.475 5.290 8.645 6.900 ;
        RECT 9.355 6.820 10.405 6.990 ;
        RECT 9.355 5.290 9.525 6.820 ;
        RECT 10.235 5.550 10.405 6.820 ;
        RECT 8.475 5.120 9.525 5.290 ;
        RECT 11.805 5.290 11.975 6.900 ;
        RECT 12.685 6.820 13.735 6.990 ;
        RECT 12.685 5.290 12.855 6.820 ;
        RECT 13.565 5.550 13.735 6.820 ;
        RECT 11.805 5.120 12.855 5.290 ;
        RECT 4.360 4.495 4.895 4.665 ;
        RECT 6.580 4.495 7.115 4.665 ;
        RECT 4.725 2.165 4.895 4.495 ;
        RECT 6.945 2.165 7.115 4.495 ;
        RECT 9.905 3.905 10.075 4.865 ;
        RECT 4.355 1.995 4.895 2.165 ;
        RECT 6.575 1.995 7.115 2.165 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 4.355 0.840 4.525 1.995 ;
        RECT 6.575 0.840 6.745 1.995 ;
        RECT 12.125 1.920 12.295 3.495 ;
        RECT 13.235 1.920 13.405 4.865 ;
        RECT 15.450 4.665 15.620 7.020 ;
        RECT 15.085 4.495 15.620 4.665 ;
        RECT 15.085 2.165 15.255 4.495 ;
        RECT 15.085 1.995 15.625 2.165 ;
        RECT 8.380 1.670 8.550 1.750 ;
        RECT 9.350 1.670 9.520 1.750 ;
        RECT 8.380 1.500 9.520 1.670 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 8.380 0.370 8.550 1.500 ;
        RECT 9.350 0.620 9.520 1.500 ;
        RECT 11.710 1.670 11.880 1.750 ;
        RECT 12.680 1.670 12.850 1.750 ;
        RECT 11.710 1.500 12.850 1.670 ;
        RECT 10.320 0.620 10.490 1.390 ;
        RECT 9.350 0.450 10.490 0.620 ;
        RECT 9.350 0.370 9.520 0.450 ;
        RECT 10.320 0.370 10.490 0.450 ;
        RECT 11.710 0.370 11.880 1.500 ;
        RECT 12.680 0.620 12.850 1.500 ;
        RECT 13.650 0.620 13.820 1.390 ;
        RECT 15.455 0.840 15.625 1.995 ;
        RECT 12.680 0.450 13.820 0.620 ;
        RECT 12.680 0.370 12.850 0.450 ;
        RECT 13.650 0.370 13.820 0.450 ;
      LAYER mcon ;
        RECT 2.505 3.245 2.675 3.415 ;
        RECT 3.985 3.245 4.155 3.415 ;
        RECT 9.905 3.985 10.075 4.155 ;
        RECT 6.945 2.505 7.115 2.675 ;
        RECT 12.125 3.245 12.295 3.415 ;
        RECT 13.235 2.505 13.405 2.675 ;
        RECT 15.085 3.985 15.255 4.155 ;
        RECT 15.085 3.245 15.255 3.415 ;
      LAYER met1 ;
        RECT 9.875 4.155 10.105 4.185 ;
        RECT 15.055 4.155 15.285 4.185 ;
        RECT 9.845 3.985 15.315 4.155 ;
        RECT 9.875 3.955 10.105 3.985 ;
        RECT 15.055 3.955 15.285 3.985 ;
        RECT 2.475 3.415 2.705 3.445 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 12.095 3.415 12.325 3.445 ;
        RECT 15.055 3.415 15.285 3.445 ;
        RECT 2.445 3.245 4.215 3.415 ;
        RECT 12.065 3.245 15.315 3.415 ;
        RECT 2.475 3.215 2.705 3.245 ;
        RECT 3.955 3.215 4.185 3.245 ;
        RECT 12.095 3.215 12.325 3.245 ;
        RECT 15.055 3.215 15.285 3.245 ;
        RECT 6.915 2.675 7.145 2.705 ;
        RECT 13.205 2.675 13.435 2.705 ;
        RECT 6.885 2.505 13.465 2.675 ;
        RECT 6.915 2.475 7.145 2.505 ;
        RECT 13.205 2.475 13.435 2.505 ;
  END
END HA






MACRO INVX1
  CLASS CORE ;
  FOREIGN INVX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.220 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 2.655 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 2.390 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 2.390 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 2.390 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT -0.170 -0.170 2.390 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 2.390 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
  END
END INVX1






MACRO INVX1_tmp
  CLASS BLOCK ;
  FOREIGN INVX1_tmp ;
  ORIGIN 0.435 0.170 ;
  SIZE 3.090 BY 7.920 ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 2.655 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 2.390 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 2.390 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 2.390 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT -0.170 -0.170 2.390 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 2.390 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
  END
END INVX1_tmp






MACRO MUX2X1
  CLASS CORE ;
  FOREIGN MUX2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.210 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN S
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
      LAYER mcon ;
        RECT 0.655 2.875 0.825 3.045 ;
        RECT 3.245 2.875 3.415 3.045 ;
      LAYER met1 ;
        RECT 0.625 3.045 0.855 3.075 ;
        RECT 3.215 3.045 3.445 3.075 ;
        RECT 0.595 2.875 3.475 3.045 ;
        RECT 0.625 2.845 0.855 2.875 ;
        RECT 3.215 2.845 3.445 2.875 ;
    END
  END S
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 12.645 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 12.380 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
        RECT 2.925 5.135 3.095 7.230 ;
        RECT 3.805 5.555 3.975 7.230 ;
        RECT 4.685 5.555 4.855 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
        RECT 6.255 5.135 6.425 7.230 ;
        RECT 7.135 5.555 7.305 7.230 ;
        RECT 8.015 5.555 8.185 7.230 ;
        RECT 8.710 4.110 9.050 7.230 ;
        RECT 9.585 5.135 9.755 7.230 ;
        RECT 10.465 5.555 10.635 7.230 ;
        RECT 11.345 5.555 11.515 7.230 ;
        RECT 12.040 4.110 12.380 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 12.380 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 12.380 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT 3.315 0.170 3.485 1.120 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT 6.645 0.170 6.815 1.120 ;
        RECT 8.710 0.170 9.050 2.720 ;
        RECT 9.975 0.170 10.145 1.120 ;
        RECT 12.040 0.170 12.380 2.720 ;
        RECT -0.170 -0.170 12.380 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 12.380 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 3.365 5.285 3.535 7.020 ;
        RECT 4.245 5.285 4.415 7.020 ;
        RECT 6.695 5.285 6.865 7.020 ;
        RECT 7.575 5.285 7.745 7.020 ;
        RECT 10.025 5.285 10.195 7.020 ;
        RECT 10.905 5.285 11.075 7.020 ;
        RECT 3.365 5.115 4.895 5.285 ;
        RECT 6.695 5.115 8.225 5.285 ;
        RECT 10.025 5.115 11.555 5.285 ;
        RECT 4.015 4.710 4.185 4.865 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 3.985 4.535 4.185 4.710 ;
        RECT 1.025 0.840 1.195 1.995 ;
        RECT 3.985 1.915 4.155 4.535 ;
        RECT 2.830 1.665 3.000 1.745 ;
        RECT 3.800 1.665 3.970 1.745 ;
        RECT 4.725 1.740 4.895 5.115 ;
        RECT 6.575 1.915 6.745 4.865 ;
        RECT 7.345 4.710 7.515 4.865 ;
        RECT 7.315 4.535 7.515 4.710 ;
        RECT 7.315 1.915 7.485 4.535 ;
        RECT 2.830 1.495 3.970 1.665 ;
        RECT 2.830 0.365 3.000 1.495 ;
        RECT 3.800 0.615 3.970 1.495 ;
        RECT 4.285 1.570 4.895 1.740 ;
        RECT 6.160 1.665 6.330 1.745 ;
        RECT 7.130 1.665 7.300 1.745 ;
        RECT 8.055 1.740 8.225 5.115 ;
        RECT 9.905 1.915 10.075 4.865 ;
        RECT 10.675 4.710 10.845 4.865 ;
        RECT 10.645 4.535 10.845 4.710 ;
        RECT 10.645 1.915 10.815 4.535 ;
        RECT 4.285 0.835 4.455 1.570 ;
        RECT 6.160 1.495 7.300 1.665 ;
        RECT 4.770 0.615 4.940 1.385 ;
        RECT 3.800 0.445 4.940 0.615 ;
        RECT 3.800 0.365 3.970 0.445 ;
        RECT 4.770 0.365 4.940 0.445 ;
        RECT 6.160 0.365 6.330 1.495 ;
        RECT 7.130 0.615 7.300 1.495 ;
        RECT 7.615 1.570 8.225 1.740 ;
        RECT 9.490 1.665 9.660 1.745 ;
        RECT 10.460 1.665 10.630 1.745 ;
        RECT 11.385 1.740 11.555 5.115 ;
        RECT 7.615 0.835 7.785 1.570 ;
        RECT 9.490 1.495 10.630 1.665 ;
        RECT 8.100 0.615 8.270 1.385 ;
        RECT 7.130 0.445 8.270 0.615 ;
        RECT 7.130 0.365 7.300 0.445 ;
        RECT 8.100 0.365 8.270 0.445 ;
        RECT 9.490 0.365 9.660 1.495 ;
        RECT 10.460 0.615 10.630 1.495 ;
        RECT 10.945 1.570 11.555 1.740 ;
        RECT 10.945 0.835 11.115 1.570 ;
        RECT 11.430 0.615 11.600 1.385 ;
        RECT 10.460 0.445 11.600 0.615 ;
        RECT 10.460 0.365 10.630 0.445 ;
        RECT 11.430 0.365 11.600 0.445 ;
      LAYER mcon ;
        RECT 1.395 3.245 1.565 3.415 ;
        RECT 4.725 2.875 4.895 3.045 ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 8.055 3.245 8.225 3.415 ;
        RECT 9.905 2.875 10.075 3.045 ;
        RECT 10.645 3.245 10.815 3.415 ;
      LAYER met1 ;
        RECT 1.365 3.415 1.595 3.445 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 8.025 3.415 8.255 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 1.335 3.245 6.805 3.415 ;
        RECT 7.995 3.245 10.875 3.415 ;
        RECT 1.365 3.215 1.595 3.245 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 8.025 3.215 8.255 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 4.695 3.045 4.925 3.075 ;
        RECT 9.875 3.045 10.105 3.075 ;
        RECT 4.665 2.875 10.135 3.045 ;
        RECT 4.695 2.845 4.925 2.875 ;
        RECT 9.875 2.845 10.105 2.875 ;
  END
END MUX2X1






MACRO NAND2X1
  CLASS CORE ;
  FOREIGN NAND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.330 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 3.765 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 3.500 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 3.500 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 3.500 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT -0.170 -0.170 3.500 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 3.500 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
  END
END NAND2X1






MACRO NAND3X1
  CLASS CORE ;
  FOREIGN NAND3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.810 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 5.245 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 4.980 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 4.980 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 4.980 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT -0.170 -0.170 4.980 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 4.980 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
  END
END NAND3X1






MACRO NOR2X1
  CLASS CORE ;
  FOREIGN NOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.330 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 3.765 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 3.500 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.145 5.555 1.315 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 3.500 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 3.500 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.610 0.615 0.780 1.745 ;
        RECT 1.580 0.615 1.750 1.390 ;
        RECT 2.550 0.615 2.720 1.390 ;
        RECT 0.610 0.445 2.720 0.615 ;
        RECT 0.610 0.170 0.780 0.445 ;
        RECT 1.095 0.170 1.265 0.445 ;
        RECT 1.580 0.170 1.750 0.445 ;
        RECT 2.065 0.170 2.235 0.445 ;
        RECT 2.550 0.170 2.720 0.445 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT -0.170 -0.170 3.500 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 3.500 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.705 5.295 0.875 7.025 ;
        RECT 1.585 6.825 2.635 6.995 ;
        RECT 1.585 5.295 1.755 6.825 ;
        RECT 0.705 5.125 1.755 5.295 ;
        RECT 2.025 5.295 2.195 6.565 ;
        RECT 2.465 5.555 2.635 6.825 ;
        RECT 2.025 5.125 2.675 5.295 ;
        RECT 0.870 4.710 1.040 4.870 ;
        RECT 1.800 4.710 1.970 4.870 ;
        RECT 0.870 4.540 1.195 4.710 ;
        RECT 1.025 1.915 1.195 4.540 ;
        RECT 1.765 4.540 1.970 4.710 ;
        RECT 1.765 1.915 1.935 4.540 ;
        RECT 2.505 1.740 2.675 5.125 ;
        RECT 1.095 1.570 2.675 1.740 ;
        RECT 1.095 0.835 1.265 1.570 ;
        RECT 2.065 0.835 2.235 1.570 ;
  END
END NOR2X1






MACRO OR2X1
  CLASS CORE ;
  FOREIGN OR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.550 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 5.985 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 5.720 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.145 5.555 1.315 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 3.920 5.185 4.090 7.230 ;
        RECT 4.800 5.185 4.970 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 5.720 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 5.720 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.610 0.615 0.780 1.745 ;
        RECT 1.580 0.615 1.750 1.390 ;
        RECT 2.550 0.615 2.720 1.390 ;
        RECT 0.610 0.445 2.720 0.615 ;
        RECT 0.610 0.170 0.780 0.445 ;
        RECT 1.095 0.170 1.265 0.445 ;
        RECT 1.580 0.170 1.750 0.445 ;
        RECT 2.065 0.170 2.235 0.445 ;
        RECT 2.550 0.170 2.720 0.445 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 3.875 0.620 4.045 1.750 ;
        RECT 4.845 0.620 5.015 1.750 ;
        RECT 3.875 0.450 5.015 0.620 ;
        RECT 3.875 0.170 4.045 0.450 ;
        RECT 4.360 0.170 4.530 0.450 ;
        RECT 4.845 0.170 5.015 0.450 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT -0.170 -0.170 5.720 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 5.720 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.705 5.295 0.875 7.025 ;
        RECT 1.585 6.825 2.635 6.995 ;
        RECT 1.585 5.295 1.755 6.825 ;
        RECT 0.705 5.125 1.755 5.295 ;
        RECT 2.025 5.295 2.195 6.565 ;
        RECT 2.465 5.555 2.635 6.825 ;
        RECT 2.025 5.125 2.675 5.295 ;
        RECT 0.870 4.710 1.040 4.870 ;
        RECT 1.800 4.710 1.970 4.870 ;
        RECT 0.870 4.540 1.195 4.710 ;
        RECT 1.025 1.915 1.195 4.540 ;
        RECT 1.765 4.540 1.970 4.710 ;
        RECT 1.765 1.915 1.935 4.540 ;
        RECT 2.505 1.740 2.675 5.125 ;
        RECT 3.985 1.920 4.155 4.865 ;
        RECT 4.360 4.665 4.530 7.020 ;
        RECT 4.360 4.495 4.895 4.665 ;
        RECT 4.725 2.165 4.895 4.495 ;
        RECT 4.355 1.995 4.895 2.165 ;
        RECT 1.095 1.570 2.675 1.740 ;
        RECT 1.095 0.835 1.265 1.570 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 4.355 0.840 4.525 1.995 ;
      LAYER mcon ;
        RECT 2.505 3.245 2.675 3.415 ;
        RECT 3.985 3.245 4.155 3.415 ;
      LAYER met1 ;
        RECT 2.475 3.415 2.705 3.445 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 2.445 3.245 4.215 3.415 ;
        RECT 2.475 3.215 2.705 3.245 ;
        RECT 3.955 3.215 4.185 3.245 ;
  END
END OR2X1






MACRO TIEHI
  CLASS CORE WELLTAP ;
  FOREIGN TIEHI ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.220 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 2.655 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 2.390 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.585 5.080 0.755 7.230 ;
        RECT 1.465 5.080 1.635 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 2.390 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 0.170 2.720 ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 2.050 -0.170 2.390 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.615 0.715 1.745 ;
        RECT 1.515 0.615 1.685 1.745 ;
        RECT 0.545 0.445 1.685 0.615 ;
        RECT 0.545 0.170 0.715 0.445 ;
        RECT 1.025 0.170 1.195 0.445 ;
        RECT 1.515 0.170 1.685 0.445 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT -0.170 -0.170 2.390 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 2.390 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.655 2.085 0.825 4.865 ;
        RECT 1.025 3.615 1.195 7.020 ;
        RECT 0.655 1.915 1.195 2.085 ;
        RECT 1.025 0.835 1.195 1.915 ;
  END
END TIEHI






MACRO TIELO
  CLASS CORE WELLTAP ;
  FOREIGN TIELO ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.220 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 2.655 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 2.390 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.585 5.080 0.755 7.230 ;
        RECT 1.465 5.080 1.635 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 2.390 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 0.170 2.720 ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 2.050 -0.170 2.390 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.615 0.715 1.745 ;
        RECT 1.515 0.615 1.685 1.745 ;
        RECT 0.545 0.445 1.685 0.615 ;
        RECT 0.545 0.170 0.715 0.445 ;
        RECT 1.025 0.170 1.195 0.445 ;
        RECT 1.515 0.170 1.685 0.445 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT -0.170 -0.170 2.390 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 2.390 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.655 4.785 0.825 4.865 ;
        RECT 1.025 4.785 1.195 7.020 ;
        RECT 0.655 4.615 1.195 4.785 ;
        RECT 0.655 1.915 0.825 4.615 ;
        RECT 1.025 0.835 1.195 3.045 ;
  END
END TIELO






MACRO TMRDFFQNX1
  CLASS CORE ;
  FOREIGN TMRDFFQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 74.370 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN D
    ANTENNAGATEAREA 3.081750 ;
    PORT
      LAYER li1 ;
        RECT 6.605 4.710 6.775 4.865 ;
        RECT 28.065 4.710 28.235 4.865 ;
        RECT 49.525 4.710 49.695 4.865 ;
        RECT 6.575 4.535 6.775 4.710 ;
        RECT 28.035 4.535 28.235 4.710 ;
        RECT 49.495 4.535 49.695 4.710 ;
        RECT 6.575 1.915 6.745 4.535 ;
        RECT 28.035 1.915 28.205 4.535 ;
        RECT 49.495 1.915 49.665 4.535 ;
      LAYER mcon ;
        RECT 6.575 2.505 6.745 2.675 ;
        RECT 28.035 2.505 28.205 2.675 ;
        RECT 49.495 2.505 49.665 2.675 ;
      LAYER met1 ;
        RECT 6.545 2.675 6.775 2.705 ;
        RECT 28.005 2.675 28.235 2.705 ;
        RECT 49.465 2.675 49.695 2.705 ;
        RECT 6.515 2.505 49.725 2.675 ;
        RECT 6.545 2.475 6.775 2.505 ;
        RECT 28.005 2.475 28.235 2.505 ;
        RECT 49.465 2.475 49.695 2.505 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.126300 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 13.265 4.710 13.435 4.865 ;
        RECT 13.235 4.535 13.435 4.710 ;
        RECT 13.235 1.915 13.405 4.535 ;
        RECT 23.595 1.915 23.765 4.865 ;
        RECT 34.725 4.710 34.895 4.865 ;
        RECT 34.695 4.535 34.895 4.710 ;
        RECT 34.695 1.915 34.865 4.535 ;
        RECT 45.055 1.915 45.225 4.865 ;
        RECT 56.185 4.710 56.355 4.865 ;
        RECT 56.155 4.535 56.355 4.710 ;
        RECT 56.155 1.915 56.325 4.535 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 13.235 4.355 13.405 4.525 ;
        RECT 23.595 4.355 23.765 4.525 ;
        RECT 34.695 4.355 34.865 4.525 ;
        RECT 45.055 4.355 45.225 4.525 ;
        RECT 56.155 4.355 56.325 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 13.205 4.525 13.435 4.555 ;
        RECT 23.565 4.525 23.795 4.555 ;
        RECT 34.665 4.525 34.895 4.555 ;
        RECT 45.025 4.525 45.255 4.555 ;
        RECT 56.125 4.525 56.355 4.555 ;
        RECT 2.075 4.520 13.465 4.525 ;
        RECT 16.745 4.520 56.385 4.525 ;
        RECT 2.075 4.365 56.385 4.520 ;
        RECT 2.075 4.355 13.465 4.365 ;
        RECT 16.745 4.355 56.385 4.365 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 13.205 4.325 13.435 4.355 ;
        RECT 23.565 4.325 23.795 4.355 ;
        RECT 34.665 4.325 34.895 4.355 ;
        RECT 45.025 4.325 45.255 4.355 ;
        RECT 56.125 4.325 56.355 4.355 ;
    END
  END CLK
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 74.805 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 74.540 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.515 5.135 5.685 7.230 ;
        RECT 6.395 5.555 6.565 7.230 ;
        RECT 7.275 5.555 7.445 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 8.845 5.135 9.015 7.230 ;
        RECT 9.725 5.555 9.895 7.230 ;
        RECT 10.605 5.555 10.775 7.230 ;
        RECT 11.300 4.110 11.640 7.230 ;
        RECT 12.175 5.135 12.345 7.230 ;
        RECT 13.055 5.555 13.225 7.230 ;
        RECT 13.935 5.555 14.105 7.230 ;
        RECT 14.630 4.110 14.970 7.230 ;
        RECT 15.505 5.135 15.675 7.230 ;
        RECT 16.385 5.555 16.555 7.230 ;
        RECT 17.265 5.555 17.435 7.230 ;
        RECT 17.960 4.110 18.300 7.230 ;
        RECT 18.835 5.135 19.005 7.230 ;
        RECT 19.715 5.555 19.885 7.230 ;
        RECT 20.595 5.555 20.765 7.230 ;
        RECT 21.290 4.110 21.630 7.230 ;
        RECT 22.465 5.215 22.635 7.230 ;
        RECT 23.345 5.555 23.515 7.230 ;
        RECT 24.225 5.555 24.395 7.230 ;
        RECT 25.105 5.555 25.275 7.230 ;
        RECT 26.100 4.110 26.440 7.230 ;
        RECT 26.975 5.135 27.145 7.230 ;
        RECT 27.855 5.555 28.025 7.230 ;
        RECT 28.735 5.555 28.905 7.230 ;
        RECT 29.430 4.110 29.770 7.230 ;
        RECT 30.305 5.135 30.475 7.230 ;
        RECT 31.185 5.555 31.355 7.230 ;
        RECT 32.065 5.555 32.235 7.230 ;
        RECT 32.760 4.110 33.100 7.230 ;
        RECT 33.635 5.135 33.805 7.230 ;
        RECT 34.515 5.555 34.685 7.230 ;
        RECT 35.395 5.555 35.565 7.230 ;
        RECT 36.090 4.110 36.430 7.230 ;
        RECT 36.965 5.135 37.135 7.230 ;
        RECT 37.845 5.555 38.015 7.230 ;
        RECT 38.725 5.555 38.895 7.230 ;
        RECT 39.420 4.110 39.760 7.230 ;
        RECT 40.295 5.135 40.465 7.230 ;
        RECT 41.175 5.555 41.345 7.230 ;
        RECT 42.055 5.555 42.225 7.230 ;
        RECT 42.750 4.110 43.090 7.230 ;
        RECT 43.925 5.215 44.095 7.230 ;
        RECT 44.805 5.555 44.975 7.230 ;
        RECT 45.685 5.555 45.855 7.230 ;
        RECT 46.565 5.555 46.735 7.230 ;
        RECT 47.560 4.110 47.900 7.230 ;
        RECT 48.435 5.135 48.605 7.230 ;
        RECT 49.315 5.555 49.485 7.230 ;
        RECT 50.195 5.555 50.365 7.230 ;
        RECT 50.890 4.110 51.230 7.230 ;
        RECT 51.765 5.135 51.935 7.230 ;
        RECT 52.645 5.555 52.815 7.230 ;
        RECT 53.525 5.555 53.695 7.230 ;
        RECT 54.220 4.110 54.560 7.230 ;
        RECT 55.095 5.135 55.265 7.230 ;
        RECT 55.975 5.555 56.145 7.230 ;
        RECT 56.855 5.555 57.025 7.230 ;
        RECT 57.550 4.110 57.890 7.230 ;
        RECT 58.425 5.135 58.595 7.230 ;
        RECT 59.305 5.555 59.475 7.230 ;
        RECT 60.185 5.555 60.355 7.230 ;
        RECT 60.880 4.110 61.220 7.230 ;
        RECT 61.755 5.135 61.925 7.230 ;
        RECT 62.635 5.555 62.805 7.230 ;
        RECT 63.515 5.555 63.685 7.230 ;
        RECT 64.210 4.110 64.550 7.230 ;
        RECT 65.085 5.125 65.255 7.230 ;
        RECT 65.965 5.555 66.135 7.230 ;
        RECT 66.845 5.125 67.015 7.230 ;
        RECT 67.540 4.110 67.880 7.230 ;
        RECT 70.870 4.110 71.210 7.230 ;
        RECT 74.200 4.110 74.540 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.625 7.315 30.795 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.435 7.315 35.605 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
        RECT 38.765 7.315 38.935 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.615 7.315 40.785 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 43.205 7.315 43.375 7.485 ;
        RECT 43.575 7.315 43.745 7.485 ;
        RECT 43.945 7.315 44.115 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 48.015 7.315 48.185 7.485 ;
        RECT 48.385 7.315 48.555 7.485 ;
        RECT 48.755 7.315 48.925 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 51.715 7.315 51.885 7.485 ;
        RECT 52.085 7.315 52.255 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 52.825 7.315 52.995 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.525 7.315 56.695 7.485 ;
        RECT 56.895 7.315 57.065 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 61.335 7.315 61.505 7.485 ;
        RECT 61.705 7.315 61.875 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.445 7.315 62.615 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.665 7.315 64.835 7.485 ;
        RECT 65.035 7.315 65.205 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.255 7.315 67.425 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.365 7.315 68.535 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.475 7.315 69.645 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.065 7.315 72.235 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.175 7.315 73.345 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 74.540 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 74.540 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.905 0.170 6.075 1.120 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.235 0.170 9.405 1.120 ;
        RECT 11.300 0.170 11.640 2.720 ;
        RECT 12.565 0.170 12.735 1.120 ;
        RECT 14.630 0.170 14.970 2.720 ;
        RECT 15.895 0.170 16.065 1.120 ;
        RECT 17.960 0.170 18.300 2.720 ;
        RECT 19.225 0.170 19.395 1.120 ;
        RECT 21.290 0.170 21.630 2.720 ;
        RECT 22.450 0.170 22.620 1.130 ;
        RECT 26.100 0.170 26.440 2.720 ;
        RECT 27.365 0.170 27.535 1.120 ;
        RECT 29.430 0.170 29.770 2.720 ;
        RECT 30.695 0.170 30.865 1.120 ;
        RECT 32.760 0.170 33.100 2.720 ;
        RECT 34.025 0.170 34.195 1.120 ;
        RECT 36.090 0.170 36.430 2.720 ;
        RECT 37.355 0.170 37.525 1.120 ;
        RECT 39.420 0.170 39.760 2.720 ;
        RECT 40.685 0.170 40.855 1.120 ;
        RECT 42.750 0.170 43.090 2.720 ;
        RECT 43.910 0.170 44.080 1.130 ;
        RECT 47.560 0.170 47.900 2.720 ;
        RECT 48.825 0.170 48.995 1.120 ;
        RECT 50.890 0.170 51.230 2.720 ;
        RECT 52.155 0.170 52.325 1.120 ;
        RECT 54.220 0.170 54.560 2.720 ;
        RECT 55.485 0.170 55.655 1.120 ;
        RECT 57.550 0.170 57.890 2.720 ;
        RECT 58.815 0.170 58.985 1.120 ;
        RECT 60.880 0.170 61.220 2.720 ;
        RECT 62.145 0.170 62.315 1.120 ;
        RECT 64.210 0.170 64.550 2.720 ;
        RECT 65.475 0.170 65.645 1.120 ;
        RECT 67.540 0.170 67.880 2.720 ;
        RECT 68.805 0.170 68.975 1.120 ;
        RECT 70.870 0.170 71.210 2.720 ;
        RECT 72.135 0.170 72.305 1.120 ;
        RECT 74.200 0.170 74.540 2.720 ;
        RECT -0.170 -0.170 74.540 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.625 -0.085 30.795 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.435 -0.085 35.605 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
        RECT 38.765 -0.085 38.935 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.615 -0.085 40.785 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 43.205 -0.085 43.375 0.085 ;
        RECT 43.575 -0.085 43.745 0.085 ;
        RECT 43.945 -0.085 44.115 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 48.015 -0.085 48.185 0.085 ;
        RECT 48.385 -0.085 48.555 0.085 ;
        RECT 48.755 -0.085 48.925 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 51.715 -0.085 51.885 0.085 ;
        RECT 52.085 -0.085 52.255 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 52.825 -0.085 52.995 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.525 -0.085 56.695 0.085 ;
        RECT 56.895 -0.085 57.065 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 61.335 -0.085 61.505 0.085 ;
        RECT 61.705 -0.085 61.875 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.445 -0.085 62.615 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.665 -0.085 64.835 0.085 ;
        RECT 65.035 -0.085 65.205 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.255 -0.085 67.425 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.365 -0.085 68.535 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.475 -0.085 69.645 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.065 -0.085 72.235 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.175 -0.085 73.345 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 74.540 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 5.955 5.285 6.125 7.020 ;
        RECT 6.835 5.285 7.005 7.020 ;
        RECT 9.285 5.285 9.455 7.020 ;
        RECT 10.165 5.285 10.335 7.020 ;
        RECT 12.615 5.285 12.785 7.020 ;
        RECT 13.495 5.285 13.665 7.020 ;
        RECT 15.945 5.285 16.115 7.020 ;
        RECT 16.825 5.285 16.995 7.020 ;
        RECT 19.275 5.285 19.445 7.020 ;
        RECT 20.155 5.285 20.325 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 5.955 5.115 7.485 5.285 ;
        RECT 9.285 5.115 10.815 5.285 ;
        RECT 12.615 5.115 14.145 5.285 ;
        RECT 15.945 5.115 17.475 5.285 ;
        RECT 19.275 5.115 20.805 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.420 1.665 5.590 1.745 ;
        RECT 6.390 1.665 6.560 1.745 ;
        RECT 7.315 1.740 7.485 5.115 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 9.935 4.710 10.105 4.865 ;
        RECT 9.905 4.535 10.105 4.710 ;
        RECT 9.905 1.915 10.075 4.535 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.420 1.495 6.560 1.665 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.420 0.365 5.590 1.495 ;
        RECT 6.390 0.615 6.560 1.495 ;
        RECT 6.875 1.570 7.485 1.740 ;
        RECT 8.750 1.665 8.920 1.745 ;
        RECT 9.720 1.665 9.890 1.745 ;
        RECT 10.645 1.740 10.815 5.115 ;
        RECT 12.495 1.915 12.665 4.865 ;
        RECT 6.875 0.835 7.045 1.570 ;
        RECT 8.750 1.495 9.890 1.665 ;
        RECT 7.360 0.615 7.530 1.385 ;
        RECT 6.390 0.445 7.530 0.615 ;
        RECT 6.390 0.365 6.560 0.445 ;
        RECT 7.360 0.365 7.530 0.445 ;
        RECT 8.750 0.365 8.920 1.495 ;
        RECT 9.720 0.615 9.890 1.495 ;
        RECT 10.205 1.570 10.815 1.740 ;
        RECT 12.080 1.665 12.250 1.745 ;
        RECT 13.050 1.665 13.220 1.745 ;
        RECT 13.975 1.740 14.145 5.115 ;
        RECT 15.825 1.915 15.995 4.865 ;
        RECT 16.595 4.710 16.765 4.865 ;
        RECT 16.565 4.535 16.765 4.710 ;
        RECT 16.565 1.915 16.735 4.535 ;
        RECT 10.205 0.835 10.375 1.570 ;
        RECT 12.080 1.495 13.220 1.665 ;
        RECT 10.690 0.615 10.860 1.385 ;
        RECT 9.720 0.445 10.860 0.615 ;
        RECT 9.720 0.365 9.890 0.445 ;
        RECT 10.690 0.365 10.860 0.445 ;
        RECT 12.080 0.365 12.250 1.495 ;
        RECT 13.050 0.615 13.220 1.495 ;
        RECT 13.535 1.570 14.145 1.740 ;
        RECT 15.410 1.665 15.580 1.745 ;
        RECT 16.380 1.665 16.550 1.745 ;
        RECT 17.305 1.740 17.475 5.115 ;
        RECT 19.155 1.915 19.325 4.865 ;
        RECT 19.925 4.710 20.095 4.865 ;
        RECT 19.895 4.535 20.095 4.710 ;
        RECT 19.895 1.915 20.065 4.535 ;
        RECT 13.535 0.835 13.705 1.570 ;
        RECT 15.410 1.495 16.550 1.665 ;
        RECT 14.020 0.615 14.190 1.385 ;
        RECT 13.050 0.445 14.190 0.615 ;
        RECT 13.050 0.365 13.220 0.445 ;
        RECT 14.020 0.365 14.190 0.445 ;
        RECT 15.410 0.365 15.580 1.495 ;
        RECT 16.380 0.615 16.550 1.495 ;
        RECT 16.865 1.570 17.475 1.740 ;
        RECT 18.740 1.665 18.910 1.745 ;
        RECT 19.710 1.665 19.880 1.745 ;
        RECT 20.635 1.740 20.805 5.115 ;
        RECT 22.905 5.240 23.075 7.020 ;
        RECT 23.785 5.240 23.955 7.020 ;
        RECT 24.665 5.240 24.835 7.020 ;
        RECT 27.415 5.285 27.585 7.020 ;
        RECT 28.295 5.285 28.465 7.020 ;
        RECT 30.745 5.285 30.915 7.020 ;
        RECT 31.625 5.285 31.795 7.020 ;
        RECT 34.075 5.285 34.245 7.020 ;
        RECT 34.955 5.285 35.125 7.020 ;
        RECT 37.405 5.285 37.575 7.020 ;
        RECT 38.285 5.285 38.455 7.020 ;
        RECT 40.735 5.285 40.905 7.020 ;
        RECT 41.615 5.285 41.785 7.020 ;
        RECT 22.905 5.070 25.615 5.240 ;
        RECT 27.415 5.115 28.945 5.285 ;
        RECT 30.745 5.115 32.275 5.285 ;
        RECT 34.075 5.115 35.605 5.285 ;
        RECT 37.405 5.115 38.935 5.285 ;
        RECT 40.735 5.115 42.265 5.285 ;
        RECT 22.485 1.915 22.655 4.865 ;
        RECT 24.705 1.915 24.875 4.865 ;
        RECT 16.865 0.835 17.035 1.570 ;
        RECT 18.740 1.495 19.880 1.665 ;
        RECT 17.350 0.615 17.520 1.385 ;
        RECT 16.380 0.445 17.520 0.615 ;
        RECT 16.380 0.365 16.550 0.445 ;
        RECT 17.350 0.365 17.520 0.445 ;
        RECT 18.740 0.365 18.910 1.495 ;
        RECT 19.710 0.615 19.880 1.495 ;
        RECT 20.195 1.570 20.805 1.740 ;
        RECT 21.965 1.675 22.135 1.755 ;
        RECT 22.935 1.675 23.105 1.755 ;
        RECT 23.905 1.675 24.075 1.755 ;
        RECT 20.195 0.835 20.365 1.570 ;
        RECT 21.965 1.505 24.075 1.675 ;
        RECT 20.680 0.615 20.850 1.385 ;
        RECT 19.710 0.445 20.850 0.615 ;
        RECT 19.710 0.365 19.880 0.445 ;
        RECT 20.680 0.365 20.850 0.445 ;
        RECT 21.965 0.375 22.135 1.505 ;
        RECT 22.935 0.625 23.105 1.505 ;
        RECT 23.905 1.425 24.075 1.505 ;
        RECT 23.425 1.080 23.595 1.160 ;
        RECT 24.475 1.080 24.645 1.755 ;
        RECT 25.445 1.750 25.615 5.070 ;
        RECT 27.295 1.915 27.465 4.865 ;
        RECT 23.425 0.910 24.645 1.080 ;
        RECT 23.425 0.830 23.595 0.910 ;
        RECT 23.905 0.625 24.075 0.705 ;
        RECT 22.935 0.455 24.075 0.625 ;
        RECT 22.935 0.375 23.105 0.455 ;
        RECT 23.905 0.375 24.075 0.455 ;
        RECT 24.475 0.625 24.645 0.910 ;
        RECT 24.960 1.580 25.615 1.750 ;
        RECT 26.880 1.665 27.050 1.745 ;
        RECT 27.850 1.665 28.020 1.745 ;
        RECT 28.775 1.740 28.945 5.115 ;
        RECT 30.625 1.915 30.795 4.865 ;
        RECT 31.395 4.710 31.565 4.865 ;
        RECT 31.365 4.535 31.565 4.710 ;
        RECT 31.365 1.915 31.535 4.535 ;
        RECT 24.960 0.845 25.130 1.580 ;
        RECT 26.880 1.495 28.020 1.665 ;
        RECT 25.445 0.625 25.615 1.395 ;
        RECT 24.475 0.455 25.615 0.625 ;
        RECT 24.475 0.375 24.645 0.455 ;
        RECT 25.445 0.375 25.615 0.455 ;
        RECT 26.880 0.365 27.050 1.495 ;
        RECT 27.850 0.615 28.020 1.495 ;
        RECT 28.335 1.570 28.945 1.740 ;
        RECT 30.210 1.665 30.380 1.745 ;
        RECT 31.180 1.665 31.350 1.745 ;
        RECT 32.105 1.740 32.275 5.115 ;
        RECT 33.955 1.915 34.125 4.865 ;
        RECT 28.335 0.835 28.505 1.570 ;
        RECT 30.210 1.495 31.350 1.665 ;
        RECT 28.820 0.615 28.990 1.385 ;
        RECT 27.850 0.445 28.990 0.615 ;
        RECT 27.850 0.365 28.020 0.445 ;
        RECT 28.820 0.365 28.990 0.445 ;
        RECT 30.210 0.365 30.380 1.495 ;
        RECT 31.180 0.615 31.350 1.495 ;
        RECT 31.665 1.570 32.275 1.740 ;
        RECT 33.540 1.665 33.710 1.745 ;
        RECT 34.510 1.665 34.680 1.745 ;
        RECT 35.435 1.740 35.605 5.115 ;
        RECT 37.285 1.915 37.455 4.865 ;
        RECT 38.055 4.710 38.225 4.865 ;
        RECT 38.025 4.535 38.225 4.710 ;
        RECT 38.025 1.915 38.195 4.535 ;
        RECT 31.665 0.835 31.835 1.570 ;
        RECT 33.540 1.495 34.680 1.665 ;
        RECT 32.150 0.615 32.320 1.385 ;
        RECT 31.180 0.445 32.320 0.615 ;
        RECT 31.180 0.365 31.350 0.445 ;
        RECT 32.150 0.365 32.320 0.445 ;
        RECT 33.540 0.365 33.710 1.495 ;
        RECT 34.510 0.615 34.680 1.495 ;
        RECT 34.995 1.570 35.605 1.740 ;
        RECT 36.870 1.665 37.040 1.745 ;
        RECT 37.840 1.665 38.010 1.745 ;
        RECT 38.765 1.740 38.935 5.115 ;
        RECT 40.615 1.915 40.785 4.865 ;
        RECT 41.385 4.710 41.555 4.865 ;
        RECT 41.355 4.535 41.555 4.710 ;
        RECT 41.355 1.915 41.525 4.535 ;
        RECT 34.995 0.835 35.165 1.570 ;
        RECT 36.870 1.495 38.010 1.665 ;
        RECT 35.480 0.615 35.650 1.385 ;
        RECT 34.510 0.445 35.650 0.615 ;
        RECT 34.510 0.365 34.680 0.445 ;
        RECT 35.480 0.365 35.650 0.445 ;
        RECT 36.870 0.365 37.040 1.495 ;
        RECT 37.840 0.615 38.010 1.495 ;
        RECT 38.325 1.570 38.935 1.740 ;
        RECT 40.200 1.665 40.370 1.745 ;
        RECT 41.170 1.665 41.340 1.745 ;
        RECT 42.095 1.740 42.265 5.115 ;
        RECT 44.365 5.240 44.535 7.020 ;
        RECT 45.245 5.240 45.415 7.020 ;
        RECT 46.125 5.240 46.295 7.020 ;
        RECT 48.875 5.285 49.045 7.020 ;
        RECT 49.755 5.285 49.925 7.020 ;
        RECT 52.205 5.285 52.375 7.020 ;
        RECT 53.085 5.285 53.255 7.020 ;
        RECT 55.535 5.285 55.705 7.020 ;
        RECT 56.415 5.285 56.585 7.020 ;
        RECT 58.865 5.285 59.035 7.020 ;
        RECT 59.745 5.285 59.915 7.020 ;
        RECT 62.195 5.285 62.365 7.020 ;
        RECT 63.075 5.285 63.245 7.020 ;
        RECT 65.525 6.825 65.705 6.995 ;
        RECT 65.525 5.295 65.695 6.825 ;
        RECT 66.405 5.295 66.575 6.995 ;
        RECT 44.365 5.070 47.075 5.240 ;
        RECT 48.875 5.115 50.405 5.285 ;
        RECT 52.205 5.115 53.735 5.285 ;
        RECT 55.535 5.115 57.065 5.285 ;
        RECT 58.865 5.115 60.395 5.285 ;
        RECT 62.195 5.115 63.725 5.285 ;
        RECT 65.525 5.125 66.575 5.295 ;
        RECT 43.945 1.915 44.115 4.865 ;
        RECT 46.165 1.915 46.335 4.865 ;
        RECT 38.325 0.835 38.495 1.570 ;
        RECT 40.200 1.495 41.340 1.665 ;
        RECT 38.810 0.615 38.980 1.385 ;
        RECT 37.840 0.445 38.980 0.615 ;
        RECT 37.840 0.365 38.010 0.445 ;
        RECT 38.810 0.365 38.980 0.445 ;
        RECT 40.200 0.365 40.370 1.495 ;
        RECT 41.170 0.615 41.340 1.495 ;
        RECT 41.655 1.570 42.265 1.740 ;
        RECT 43.425 1.675 43.595 1.755 ;
        RECT 44.395 1.675 44.565 1.755 ;
        RECT 45.365 1.675 45.535 1.755 ;
        RECT 41.655 0.835 41.825 1.570 ;
        RECT 43.425 1.505 45.535 1.675 ;
        RECT 42.140 0.615 42.310 1.385 ;
        RECT 41.170 0.445 42.310 0.615 ;
        RECT 41.170 0.365 41.340 0.445 ;
        RECT 42.140 0.365 42.310 0.445 ;
        RECT 43.425 0.375 43.595 1.505 ;
        RECT 44.395 0.625 44.565 1.505 ;
        RECT 45.365 1.425 45.535 1.505 ;
        RECT 44.885 1.080 45.055 1.160 ;
        RECT 45.935 1.080 46.105 1.755 ;
        RECT 46.905 1.750 47.075 5.070 ;
        RECT 48.755 1.915 48.925 4.865 ;
        RECT 44.885 0.910 46.105 1.080 ;
        RECT 44.885 0.830 45.055 0.910 ;
        RECT 45.365 0.625 45.535 0.705 ;
        RECT 44.395 0.455 45.535 0.625 ;
        RECT 44.395 0.375 44.565 0.455 ;
        RECT 45.365 0.375 45.535 0.455 ;
        RECT 45.935 0.625 46.105 0.910 ;
        RECT 46.420 1.580 47.075 1.750 ;
        RECT 48.340 1.665 48.510 1.745 ;
        RECT 49.310 1.665 49.480 1.745 ;
        RECT 50.235 1.740 50.405 5.115 ;
        RECT 52.085 1.915 52.255 4.865 ;
        RECT 52.855 4.710 53.025 4.865 ;
        RECT 52.825 4.535 53.025 4.710 ;
        RECT 52.825 1.915 52.995 4.535 ;
        RECT 46.420 0.845 46.590 1.580 ;
        RECT 48.340 1.495 49.480 1.665 ;
        RECT 46.905 0.625 47.075 1.395 ;
        RECT 45.935 0.455 47.075 0.625 ;
        RECT 45.935 0.375 46.105 0.455 ;
        RECT 46.905 0.375 47.075 0.455 ;
        RECT 48.340 0.365 48.510 1.495 ;
        RECT 49.310 0.615 49.480 1.495 ;
        RECT 49.795 1.570 50.405 1.740 ;
        RECT 51.670 1.665 51.840 1.745 ;
        RECT 52.640 1.665 52.810 1.745 ;
        RECT 53.565 1.740 53.735 5.115 ;
        RECT 55.415 1.915 55.585 4.865 ;
        RECT 49.795 0.835 49.965 1.570 ;
        RECT 51.670 1.495 52.810 1.665 ;
        RECT 50.280 0.615 50.450 1.385 ;
        RECT 49.310 0.445 50.450 0.615 ;
        RECT 49.310 0.365 49.480 0.445 ;
        RECT 50.280 0.365 50.450 0.445 ;
        RECT 51.670 0.365 51.840 1.495 ;
        RECT 52.640 0.615 52.810 1.495 ;
        RECT 53.125 1.570 53.735 1.740 ;
        RECT 55.000 1.665 55.170 1.745 ;
        RECT 55.970 1.665 56.140 1.745 ;
        RECT 56.895 1.740 57.065 5.115 ;
        RECT 58.745 1.915 58.915 4.865 ;
        RECT 59.515 4.710 59.685 4.865 ;
        RECT 59.485 4.535 59.685 4.710 ;
        RECT 59.485 1.915 59.655 4.535 ;
        RECT 53.125 0.835 53.295 1.570 ;
        RECT 55.000 1.495 56.140 1.665 ;
        RECT 53.610 0.615 53.780 1.385 ;
        RECT 52.640 0.445 53.780 0.615 ;
        RECT 52.640 0.365 52.810 0.445 ;
        RECT 53.610 0.365 53.780 0.445 ;
        RECT 55.000 0.365 55.170 1.495 ;
        RECT 55.970 0.615 56.140 1.495 ;
        RECT 56.455 1.570 57.065 1.740 ;
        RECT 58.330 1.665 58.500 1.745 ;
        RECT 59.300 1.665 59.470 1.745 ;
        RECT 60.225 1.740 60.395 5.115 ;
        RECT 62.075 1.915 62.245 4.865 ;
        RECT 62.845 4.710 63.015 4.865 ;
        RECT 62.815 4.535 63.015 4.710 ;
        RECT 62.815 1.915 62.985 4.535 ;
        RECT 56.455 0.835 56.625 1.570 ;
        RECT 58.330 1.495 59.470 1.665 ;
        RECT 56.940 0.615 57.110 1.385 ;
        RECT 55.970 0.445 57.110 0.615 ;
        RECT 55.970 0.365 56.140 0.445 ;
        RECT 56.940 0.365 57.110 0.445 ;
        RECT 58.330 0.365 58.500 1.495 ;
        RECT 59.300 0.615 59.470 1.495 ;
        RECT 59.785 1.570 60.395 1.740 ;
        RECT 61.660 1.665 61.830 1.745 ;
        RECT 62.630 1.665 62.800 1.745 ;
        RECT 63.555 1.740 63.725 5.115 ;
        RECT 66.405 5.045 66.575 5.125 ;
        RECT 68.405 6.825 70.335 6.995 ;
        RECT 68.405 5.045 68.575 6.825 ;
        RECT 68.845 5.295 69.015 6.565 ;
        RECT 69.285 5.555 69.455 6.825 ;
        RECT 69.725 5.295 69.895 6.565 ;
        RECT 70.165 5.375 70.335 6.825 ;
        RECT 71.745 6.825 73.675 6.995 ;
        RECT 68.845 5.125 69.895 5.295 ;
        RECT 69.725 5.045 69.895 5.125 ;
        RECT 71.745 5.045 71.915 6.825 ;
        RECT 72.185 5.295 72.355 6.565 ;
        RECT 72.625 5.555 72.795 6.825 ;
        RECT 73.065 5.295 73.235 6.565 ;
        RECT 73.505 5.555 73.675 6.825 ;
        RECT 72.185 5.125 73.715 5.295 ;
        RECT 65.035 1.915 65.205 4.870 ;
        RECT 66.185 4.710 66.355 4.870 ;
        RECT 66.145 4.540 66.355 4.710 ;
        RECT 66.145 1.915 66.315 4.540 ;
        RECT 68.735 1.915 68.905 4.870 ;
        RECT 70.215 1.915 70.385 4.870 ;
        RECT 71.695 1.915 71.865 4.870 ;
        RECT 72.805 4.540 72.995 4.870 ;
        RECT 72.805 1.915 72.975 4.540 ;
        RECT 59.785 0.835 59.955 1.570 ;
        RECT 61.660 1.495 62.800 1.665 ;
        RECT 60.270 0.615 60.440 1.385 ;
        RECT 59.300 0.445 60.440 0.615 ;
        RECT 59.300 0.365 59.470 0.445 ;
        RECT 60.270 0.365 60.440 0.445 ;
        RECT 61.660 0.365 61.830 1.495 ;
        RECT 62.630 0.615 62.800 1.495 ;
        RECT 63.115 1.570 63.725 1.740 ;
        RECT 64.990 1.665 65.160 1.745 ;
        RECT 65.960 1.665 66.130 1.745 ;
        RECT 63.115 0.835 63.285 1.570 ;
        RECT 64.990 1.495 66.130 1.665 ;
        RECT 63.600 0.615 63.770 1.385 ;
        RECT 62.630 0.445 63.770 0.615 ;
        RECT 62.630 0.365 62.800 0.445 ;
        RECT 63.600 0.365 63.770 0.445 ;
        RECT 64.990 0.365 65.160 1.495 ;
        RECT 65.960 0.615 66.130 1.495 ;
        RECT 66.445 1.170 66.615 1.345 ;
        RECT 66.440 1.015 66.615 1.170 ;
        RECT 66.440 0.835 66.610 1.015 ;
        RECT 66.930 0.615 67.100 1.745 ;
        RECT 65.960 0.445 67.100 0.615 ;
        RECT 65.960 0.365 66.130 0.445 ;
        RECT 66.930 0.365 67.100 0.445 ;
        RECT 68.320 1.665 68.490 1.745 ;
        RECT 69.290 1.665 69.460 1.745 ;
        RECT 68.320 1.495 69.460 1.665 ;
        RECT 68.320 0.365 68.490 1.495 ;
        RECT 69.290 0.615 69.460 1.495 ;
        RECT 69.775 0.835 69.945 1.345 ;
        RECT 70.260 0.615 70.430 1.745 ;
        RECT 69.290 0.445 70.430 0.615 ;
        RECT 69.290 0.365 69.460 0.445 ;
        RECT 70.260 0.365 70.430 0.445 ;
        RECT 71.650 1.665 71.820 1.745 ;
        RECT 72.620 1.665 72.790 1.745 ;
        RECT 73.545 1.730 73.715 5.125 ;
        RECT 71.650 1.495 72.790 1.665 ;
        RECT 71.650 0.365 71.820 1.495 ;
        RECT 72.620 0.615 72.790 1.495 ;
        RECT 73.105 1.560 73.715 1.730 ;
        RECT 73.105 0.835 73.275 1.560 ;
        RECT 73.590 0.615 73.760 1.390 ;
        RECT 72.620 0.445 73.760 0.615 ;
        RECT 72.620 0.365 72.790 0.445 ;
        RECT 73.590 0.365 73.760 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 7.315 3.245 7.485 3.415 ;
        RECT 9.165 3.245 9.335 3.415 ;
        RECT 9.905 3.985 10.075 4.155 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 12.495 3.245 12.665 3.415 ;
        RECT 13.975 3.985 14.145 4.155 ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 16.565 2.875 16.735 3.045 ;
        RECT 17.305 3.615 17.475 3.785 ;
        RECT 19.155 3.615 19.325 3.785 ;
        RECT 19.895 3.985 20.065 4.155 ;
        RECT 20.635 2.875 20.805 3.045 ;
        RECT 22.485 3.985 22.655 4.155 ;
        RECT 24.705 3.245 24.875 3.415 ;
        RECT 25.445 3.615 25.615 3.785 ;
        RECT 27.295 3.615 27.465 3.785 ;
        RECT 28.775 3.245 28.945 3.415 ;
        RECT 30.625 3.245 30.795 3.415 ;
        RECT 31.365 3.985 31.535 4.155 ;
        RECT 32.105 3.245 32.275 3.415 ;
        RECT 33.955 3.245 34.125 3.415 ;
        RECT 35.435 3.985 35.605 4.155 ;
        RECT 37.285 3.615 37.455 3.785 ;
        RECT 38.025 2.135 38.195 2.305 ;
        RECT 38.765 3.615 38.935 3.785 ;
        RECT 40.615 3.615 40.785 3.785 ;
        RECT 41.355 3.985 41.525 4.155 ;
        RECT 66.405 5.125 66.575 5.295 ;
        RECT 42.095 2.135 42.265 2.305 ;
        RECT 43.945 3.985 44.115 4.155 ;
        RECT 46.165 3.245 46.335 3.415 ;
        RECT 46.905 3.615 47.075 3.785 ;
        RECT 48.755 3.615 48.925 3.785 ;
        RECT 50.235 3.245 50.405 3.415 ;
        RECT 52.085 3.245 52.255 3.415 ;
        RECT 52.825 3.985 52.995 4.155 ;
        RECT 53.565 3.245 53.735 3.415 ;
        RECT 55.415 3.245 55.585 3.415 ;
        RECT 56.895 3.985 57.065 4.155 ;
        RECT 58.745 3.615 58.915 3.785 ;
        RECT 59.485 3.615 59.655 3.785 ;
        RECT 60.225 4.355 60.395 4.525 ;
        RECT 62.075 4.355 62.245 4.525 ;
        RECT 62.815 3.985 62.985 4.155 ;
        RECT 68.405 5.125 68.575 5.295 ;
        RECT 69.725 5.125 69.895 5.295 ;
        RECT 71.745 5.125 71.915 5.295 ;
        RECT 63.555 3.615 63.725 3.785 ;
        RECT 65.035 4.355 65.205 4.525 ;
        RECT 65.035 3.615 65.205 3.785 ;
        RECT 66.145 3.985 66.315 4.155 ;
        RECT 66.145 2.135 66.315 2.305 ;
        RECT 68.735 4.355 68.905 4.525 ;
        RECT 70.215 2.875 70.385 3.045 ;
        RECT 70.215 1.995 70.385 2.165 ;
        RECT 71.695 1.995 71.865 2.165 ;
        RECT 72.805 3.985 72.975 4.155 ;
        RECT 66.445 1.095 66.615 1.265 ;
        RECT 69.775 1.095 69.945 1.265 ;
        RECT 73.105 1.095 73.275 1.265 ;
      LAYER met1 ;
        RECT 66.375 5.295 66.605 5.325 ;
        RECT 68.375 5.295 68.605 5.325 ;
        RECT 69.695 5.295 69.925 5.325 ;
        RECT 71.715 5.295 71.945 5.325 ;
        RECT 66.345 5.125 68.635 5.295 ;
        RECT 69.665 5.125 71.975 5.295 ;
        RECT 66.375 5.095 66.605 5.125 ;
        RECT 68.375 5.095 68.605 5.125 ;
        RECT 69.695 5.095 69.925 5.125 ;
        RECT 71.715 5.095 71.945 5.125 ;
        RECT 60.195 4.525 60.425 4.555 ;
        RECT 62.045 4.525 62.275 4.555 ;
        RECT 65.005 4.525 65.235 4.555 ;
        RECT 68.705 4.525 68.935 4.555 ;
        RECT 60.165 4.355 62.305 4.525 ;
        RECT 64.975 4.355 68.965 4.525 ;
        RECT 60.195 4.325 60.425 4.355 ;
        RECT 62.045 4.325 62.275 4.355 ;
        RECT 65.005 4.325 65.235 4.355 ;
        RECT 68.705 4.325 68.935 4.355 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 9.875 4.155 10.105 4.185 ;
        RECT 13.945 4.155 14.175 4.185 ;
        RECT 19.865 4.155 20.095 4.185 ;
        RECT 22.455 4.155 22.685 4.185 ;
        RECT 31.335 4.155 31.565 4.185 ;
        RECT 35.405 4.155 35.635 4.185 ;
        RECT 41.325 4.155 41.555 4.185 ;
        RECT 43.915 4.155 44.145 4.185 ;
        RECT 52.795 4.155 53.025 4.185 ;
        RECT 56.865 4.155 57.095 4.185 ;
        RECT 62.785 4.155 63.015 4.185 ;
        RECT 66.115 4.155 66.345 4.185 ;
        RECT 72.775 4.155 73.005 4.185 ;
        RECT 0.965 3.985 20.125 4.155 ;
        RECT 22.425 3.985 41.585 4.155 ;
        RECT 43.885 3.985 63.045 4.155 ;
        RECT 66.085 3.985 73.035 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 9.875 3.955 10.105 3.985 ;
        RECT 13.945 3.955 14.175 3.985 ;
        RECT 19.865 3.955 20.095 3.985 ;
        RECT 22.455 3.955 22.685 3.985 ;
        RECT 31.335 3.955 31.565 3.985 ;
        RECT 35.405 3.955 35.635 3.985 ;
        RECT 41.325 3.955 41.555 3.985 ;
        RECT 43.915 3.955 44.145 3.985 ;
        RECT 52.795 3.955 53.025 3.985 ;
        RECT 56.865 3.955 57.095 3.985 ;
        RECT 62.785 3.955 63.015 3.985 ;
        RECT 66.115 3.955 66.345 3.985 ;
        RECT 72.775 3.955 73.005 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 17.275 3.785 17.505 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 25.415 3.785 25.645 3.815 ;
        RECT 27.265 3.785 27.495 3.815 ;
        RECT 37.255 3.785 37.485 3.815 ;
        RECT 38.735 3.785 38.965 3.815 ;
        RECT 40.585 3.785 40.815 3.815 ;
        RECT 46.875 3.785 47.105 3.815 ;
        RECT 48.725 3.785 48.955 3.815 ;
        RECT 58.715 3.785 58.945 3.815 ;
        RECT 59.455 3.785 59.685 3.815 ;
        RECT 63.525 3.785 63.755 3.815 ;
        RECT 65.005 3.785 65.235 3.815 ;
        RECT 3.925 3.615 16.055 3.785 ;
        RECT 17.245 3.615 19.385 3.785 ;
        RECT 25.385 3.615 37.515 3.785 ;
        RECT 38.705 3.615 40.845 3.785 ;
        RECT 46.845 3.615 58.975 3.785 ;
        RECT 59.425 3.615 65.265 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 17.275 3.585 17.505 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
        RECT 25.415 3.585 25.645 3.615 ;
        RECT 27.265 3.585 27.495 3.615 ;
        RECT 37.255 3.585 37.485 3.615 ;
        RECT 38.735 3.585 38.965 3.615 ;
        RECT 40.585 3.585 40.815 3.615 ;
        RECT 46.875 3.585 47.105 3.615 ;
        RECT 48.725 3.585 48.955 3.615 ;
        RECT 58.715 3.585 58.945 3.615 ;
        RECT 59.455 3.585 59.685 3.615 ;
        RECT 63.525 3.585 63.755 3.615 ;
        RECT 65.005 3.585 65.235 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 7.285 3.415 7.515 3.445 ;
        RECT 9.135 3.415 9.365 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.465 3.415 12.695 3.445 ;
        RECT 24.675 3.415 24.905 3.445 ;
        RECT 28.745 3.415 28.975 3.445 ;
        RECT 30.595 3.415 30.825 3.445 ;
        RECT 32.075 3.415 32.305 3.445 ;
        RECT 33.925 3.415 34.155 3.445 ;
        RECT 46.135 3.415 46.365 3.445 ;
        RECT 50.205 3.415 50.435 3.445 ;
        RECT 52.055 3.415 52.285 3.445 ;
        RECT 53.535 3.415 53.765 3.445 ;
        RECT 55.385 3.415 55.615 3.445 ;
        RECT 3.185 3.245 9.395 3.415 ;
        RECT 10.585 3.245 12.725 3.415 ;
        RECT 24.645 3.245 30.855 3.415 ;
        RECT 32.045 3.245 34.185 3.415 ;
        RECT 46.105 3.245 52.315 3.415 ;
        RECT 53.505 3.245 55.645 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 7.285 3.215 7.515 3.245 ;
        RECT 9.135 3.215 9.365 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.465 3.215 12.695 3.245 ;
        RECT 24.675 3.215 24.905 3.245 ;
        RECT 28.745 3.215 28.975 3.245 ;
        RECT 30.595 3.215 30.825 3.245 ;
        RECT 32.075 3.215 32.305 3.245 ;
        RECT 33.925 3.215 34.155 3.245 ;
        RECT 46.135 3.215 46.365 3.245 ;
        RECT 50.205 3.215 50.435 3.245 ;
        RECT 52.055 3.215 52.285 3.245 ;
        RECT 53.535 3.215 53.765 3.245 ;
        RECT 55.385 3.215 55.615 3.245 ;
        RECT 16.535 3.045 16.765 3.075 ;
        RECT 20.605 3.045 20.835 3.075 ;
        RECT 70.185 3.045 70.415 3.075 ;
        RECT 16.505 2.875 70.445 3.045 ;
        RECT 16.535 2.845 16.765 2.875 ;
        RECT 20.605 2.845 20.835 2.875 ;
        RECT 70.185 2.845 70.415 2.875 ;
        RECT 37.995 2.305 38.225 2.335 ;
        RECT 42.065 2.305 42.295 2.335 ;
        RECT 66.115 2.305 66.345 2.335 ;
        RECT 37.965 2.135 66.375 2.305 ;
        RECT 70.185 2.165 70.415 2.195 ;
        RECT 71.665 2.165 71.895 2.195 ;
        RECT 37.995 2.105 38.225 2.135 ;
        RECT 42.065 2.105 42.295 2.135 ;
        RECT 66.115 2.105 66.345 2.135 ;
        RECT 70.155 1.995 71.925 2.165 ;
        RECT 70.185 1.965 70.415 1.995 ;
        RECT 71.665 1.965 71.895 1.995 ;
        RECT 66.415 1.265 66.645 1.295 ;
        RECT 69.745 1.265 69.975 1.295 ;
        RECT 73.075 1.265 73.305 1.295 ;
        RECT 66.385 1.095 73.335 1.265 ;
        RECT 66.415 1.065 66.645 1.095 ;
        RECT 69.745 1.065 69.975 1.095 ;
        RECT 73.075 1.065 73.305 1.095 ;
  END
END TMRDFFQNX1






MACRO TMRDFFQX1
  CLASS CORE ;
  FOREIGN TMRDFFQX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 76.590 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN D
    ANTENNAGATEAREA 3.081750 ;
    PORT
      LAYER li1 ;
        RECT 6.605 4.710 6.775 4.865 ;
        RECT 28.065 4.710 28.235 4.865 ;
        RECT 49.525 4.710 49.695 4.865 ;
        RECT 6.575 4.535 6.775 4.710 ;
        RECT 28.035 4.535 28.235 4.710 ;
        RECT 49.495 4.535 49.695 4.710 ;
        RECT 6.575 1.915 6.745 4.535 ;
        RECT 28.035 1.915 28.205 4.535 ;
        RECT 49.495 1.915 49.665 4.535 ;
      LAYER mcon ;
        RECT 6.575 2.505 6.745 2.675 ;
        RECT 28.035 2.505 28.205 2.675 ;
        RECT 49.495 2.505 49.665 2.675 ;
      LAYER met1 ;
        RECT 6.545 2.675 6.775 2.705 ;
        RECT 28.005 2.675 28.235 2.705 ;
        RECT 49.465 2.675 49.695 2.705 ;
        RECT 6.515 2.505 49.725 2.675 ;
        RECT 6.545 2.475 6.775 2.505 ;
        RECT 28.005 2.475 28.235 2.505 ;
        RECT 49.465 2.475 49.695 2.505 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.126300 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 13.265 4.710 13.435 4.865 ;
        RECT 13.235 4.535 13.435 4.710 ;
        RECT 13.235 1.915 13.405 4.535 ;
        RECT 23.595 1.915 23.765 4.865 ;
        RECT 34.725 4.710 34.895 4.865 ;
        RECT 34.695 4.535 34.895 4.710 ;
        RECT 34.695 1.915 34.865 4.535 ;
        RECT 45.055 1.915 45.225 4.865 ;
        RECT 56.185 4.710 56.355 4.865 ;
        RECT 56.155 4.535 56.355 4.710 ;
        RECT 56.155 1.915 56.325 4.535 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 13.235 4.355 13.405 4.525 ;
        RECT 23.595 4.355 23.765 4.525 ;
        RECT 34.695 4.355 34.865 4.525 ;
        RECT 45.055 4.355 45.225 4.525 ;
        RECT 56.155 4.355 56.325 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 13.205 4.525 13.435 4.555 ;
        RECT 23.565 4.525 23.795 4.555 ;
        RECT 34.665 4.525 34.895 4.555 ;
        RECT 45.025 4.525 45.255 4.555 ;
        RECT 56.125 4.525 56.355 4.555 ;
        RECT 2.075 4.520 13.465 4.525 ;
        RECT 16.745 4.520 56.385 4.525 ;
        RECT 2.075 4.365 56.385 4.520 ;
        RECT 2.075 4.355 13.465 4.365 ;
        RECT 16.745 4.355 56.385 4.365 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 13.205 4.325 13.435 4.355 ;
        RECT 23.565 4.325 23.795 4.355 ;
        RECT 34.665 4.325 34.895 4.355 ;
        RECT 45.025 4.325 45.255 4.355 ;
        RECT 56.125 4.325 56.355 4.355 ;
    END
  END CLK
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 77.025 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 76.760 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.515 5.135 5.685 7.230 ;
        RECT 6.395 5.555 6.565 7.230 ;
        RECT 7.275 5.555 7.445 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 8.845 5.135 9.015 7.230 ;
        RECT 9.725 5.555 9.895 7.230 ;
        RECT 10.605 5.555 10.775 7.230 ;
        RECT 11.300 4.110 11.640 7.230 ;
        RECT 12.175 5.135 12.345 7.230 ;
        RECT 13.055 5.555 13.225 7.230 ;
        RECT 13.935 5.555 14.105 7.230 ;
        RECT 14.630 4.110 14.970 7.230 ;
        RECT 15.505 5.135 15.675 7.230 ;
        RECT 16.385 5.555 16.555 7.230 ;
        RECT 17.265 5.555 17.435 7.230 ;
        RECT 17.960 4.110 18.300 7.230 ;
        RECT 18.835 5.135 19.005 7.230 ;
        RECT 19.715 5.555 19.885 7.230 ;
        RECT 20.595 5.555 20.765 7.230 ;
        RECT 21.290 4.110 21.630 7.230 ;
        RECT 22.465 5.215 22.635 7.230 ;
        RECT 23.345 5.555 23.515 7.230 ;
        RECT 24.225 5.555 24.395 7.230 ;
        RECT 25.105 5.555 25.275 7.230 ;
        RECT 26.100 4.110 26.440 7.230 ;
        RECT 26.975 5.135 27.145 7.230 ;
        RECT 27.855 5.555 28.025 7.230 ;
        RECT 28.735 5.555 28.905 7.230 ;
        RECT 29.430 4.110 29.770 7.230 ;
        RECT 30.305 5.135 30.475 7.230 ;
        RECT 31.185 5.555 31.355 7.230 ;
        RECT 32.065 5.555 32.235 7.230 ;
        RECT 32.760 4.110 33.100 7.230 ;
        RECT 33.635 5.135 33.805 7.230 ;
        RECT 34.515 5.555 34.685 7.230 ;
        RECT 35.395 5.555 35.565 7.230 ;
        RECT 36.090 4.110 36.430 7.230 ;
        RECT 36.965 5.135 37.135 7.230 ;
        RECT 37.845 5.555 38.015 7.230 ;
        RECT 38.725 5.555 38.895 7.230 ;
        RECT 39.420 4.110 39.760 7.230 ;
        RECT 40.295 5.135 40.465 7.230 ;
        RECT 41.175 5.555 41.345 7.230 ;
        RECT 42.055 5.555 42.225 7.230 ;
        RECT 42.750 4.110 43.090 7.230 ;
        RECT 43.925 5.215 44.095 7.230 ;
        RECT 44.805 5.555 44.975 7.230 ;
        RECT 45.685 5.555 45.855 7.230 ;
        RECT 46.565 5.555 46.735 7.230 ;
        RECT 47.560 4.110 47.900 7.230 ;
        RECT 48.435 5.135 48.605 7.230 ;
        RECT 49.315 5.555 49.485 7.230 ;
        RECT 50.195 5.555 50.365 7.230 ;
        RECT 50.890 4.110 51.230 7.230 ;
        RECT 51.765 5.135 51.935 7.230 ;
        RECT 52.645 5.555 52.815 7.230 ;
        RECT 53.525 5.555 53.695 7.230 ;
        RECT 54.220 4.110 54.560 7.230 ;
        RECT 55.095 5.135 55.265 7.230 ;
        RECT 55.975 5.555 56.145 7.230 ;
        RECT 56.855 5.555 57.025 7.230 ;
        RECT 57.550 4.110 57.890 7.230 ;
        RECT 58.425 5.135 58.595 7.230 ;
        RECT 59.305 5.555 59.475 7.230 ;
        RECT 60.185 5.555 60.355 7.230 ;
        RECT 60.880 4.110 61.220 7.230 ;
        RECT 61.755 5.135 61.925 7.230 ;
        RECT 62.635 5.555 62.805 7.230 ;
        RECT 63.515 5.555 63.685 7.230 ;
        RECT 64.210 4.110 64.550 7.230 ;
        RECT 65.085 5.125 65.255 7.230 ;
        RECT 65.965 5.555 66.135 7.230 ;
        RECT 66.845 5.125 67.015 7.230 ;
        RECT 67.540 4.110 67.880 7.230 ;
        RECT 70.870 4.110 71.210 7.230 ;
        RECT 74.200 4.110 74.540 7.230 ;
        RECT 74.960 5.185 75.130 7.230 ;
        RECT 75.840 5.185 76.010 7.230 ;
        RECT 76.420 4.110 76.760 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.625 7.315 30.795 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.435 7.315 35.605 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
        RECT 38.765 7.315 38.935 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.615 7.315 40.785 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 43.205 7.315 43.375 7.485 ;
        RECT 43.575 7.315 43.745 7.485 ;
        RECT 43.945 7.315 44.115 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 48.015 7.315 48.185 7.485 ;
        RECT 48.385 7.315 48.555 7.485 ;
        RECT 48.755 7.315 48.925 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 51.715 7.315 51.885 7.485 ;
        RECT 52.085 7.315 52.255 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 52.825 7.315 52.995 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.525 7.315 56.695 7.485 ;
        RECT 56.895 7.315 57.065 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 61.335 7.315 61.505 7.485 ;
        RECT 61.705 7.315 61.875 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.445 7.315 62.615 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.665 7.315 64.835 7.485 ;
        RECT 65.035 7.315 65.205 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.255 7.315 67.425 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.365 7.315 68.535 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.475 7.315 69.645 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.065 7.315 72.235 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.175 7.315 73.345 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
        RECT 74.655 7.315 74.825 7.485 ;
        RECT 75.025 7.315 75.195 7.485 ;
        RECT 75.395 7.315 75.565 7.485 ;
        RECT 75.765 7.315 75.935 7.485 ;
        RECT 76.135 7.315 76.305 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 76.760 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 76.760 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.905 0.170 6.075 1.120 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.235 0.170 9.405 1.120 ;
        RECT 11.300 0.170 11.640 2.720 ;
        RECT 12.565 0.170 12.735 1.120 ;
        RECT 14.630 0.170 14.970 2.720 ;
        RECT 15.895 0.170 16.065 1.120 ;
        RECT 17.960 0.170 18.300 2.720 ;
        RECT 19.225 0.170 19.395 1.120 ;
        RECT 21.290 0.170 21.630 2.720 ;
        RECT 22.450 0.170 22.620 1.130 ;
        RECT 26.100 0.170 26.440 2.720 ;
        RECT 27.365 0.170 27.535 1.120 ;
        RECT 29.430 0.170 29.770 2.720 ;
        RECT 30.695 0.170 30.865 1.120 ;
        RECT 32.760 0.170 33.100 2.720 ;
        RECT 34.025 0.170 34.195 1.120 ;
        RECT 36.090 0.170 36.430 2.720 ;
        RECT 37.355 0.170 37.525 1.120 ;
        RECT 39.420 0.170 39.760 2.720 ;
        RECT 40.685 0.170 40.855 1.120 ;
        RECT 42.750 0.170 43.090 2.720 ;
        RECT 43.910 0.170 44.080 1.130 ;
        RECT 47.560 0.170 47.900 2.720 ;
        RECT 48.825 0.170 48.995 1.120 ;
        RECT 50.890 0.170 51.230 2.720 ;
        RECT 52.155 0.170 52.325 1.120 ;
        RECT 54.220 0.170 54.560 2.720 ;
        RECT 55.485 0.170 55.655 1.120 ;
        RECT 57.550 0.170 57.890 2.720 ;
        RECT 58.815 0.170 58.985 1.120 ;
        RECT 60.880 0.170 61.220 2.720 ;
        RECT 62.145 0.170 62.315 1.120 ;
        RECT 64.210 0.170 64.550 2.720 ;
        RECT 65.475 0.170 65.645 1.120 ;
        RECT 67.540 0.170 67.880 2.720 ;
        RECT 68.805 0.170 68.975 1.120 ;
        RECT 70.870 0.170 71.210 2.720 ;
        RECT 72.135 0.170 72.305 1.120 ;
        RECT 74.200 0.170 74.540 2.720 ;
        RECT 74.915 0.620 75.085 1.750 ;
        RECT 75.885 0.620 76.055 1.750 ;
        RECT 74.915 0.450 76.055 0.620 ;
        RECT 74.915 0.170 75.085 0.450 ;
        RECT 75.400 0.170 75.570 0.450 ;
        RECT 75.885 0.170 76.055 0.450 ;
        RECT 76.420 0.170 76.760 2.720 ;
        RECT -0.170 -0.170 76.760 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.625 -0.085 30.795 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.435 -0.085 35.605 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
        RECT 38.765 -0.085 38.935 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.615 -0.085 40.785 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 43.205 -0.085 43.375 0.085 ;
        RECT 43.575 -0.085 43.745 0.085 ;
        RECT 43.945 -0.085 44.115 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 48.015 -0.085 48.185 0.085 ;
        RECT 48.385 -0.085 48.555 0.085 ;
        RECT 48.755 -0.085 48.925 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 51.715 -0.085 51.885 0.085 ;
        RECT 52.085 -0.085 52.255 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 52.825 -0.085 52.995 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.525 -0.085 56.695 0.085 ;
        RECT 56.895 -0.085 57.065 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 61.335 -0.085 61.505 0.085 ;
        RECT 61.705 -0.085 61.875 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.445 -0.085 62.615 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.665 -0.085 64.835 0.085 ;
        RECT 65.035 -0.085 65.205 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.255 -0.085 67.425 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.365 -0.085 68.535 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.475 -0.085 69.645 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.065 -0.085 72.235 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.175 -0.085 73.345 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
        RECT 74.655 -0.085 74.825 0.085 ;
        RECT 75.025 -0.085 75.195 0.085 ;
        RECT 75.395 -0.085 75.565 0.085 ;
        RECT 75.765 -0.085 75.935 0.085 ;
        RECT 76.135 -0.085 76.305 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 76.760 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 5.955 5.285 6.125 7.020 ;
        RECT 6.835 5.285 7.005 7.020 ;
        RECT 9.285 5.285 9.455 7.020 ;
        RECT 10.165 5.285 10.335 7.020 ;
        RECT 12.615 5.285 12.785 7.020 ;
        RECT 13.495 5.285 13.665 7.020 ;
        RECT 15.945 5.285 16.115 7.020 ;
        RECT 16.825 5.285 16.995 7.020 ;
        RECT 19.275 5.285 19.445 7.020 ;
        RECT 20.155 5.285 20.325 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 5.955 5.115 7.485 5.285 ;
        RECT 9.285 5.115 10.815 5.285 ;
        RECT 12.615 5.115 14.145 5.285 ;
        RECT 15.945 5.115 17.475 5.285 ;
        RECT 19.275 5.115 20.805 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.420 1.665 5.590 1.745 ;
        RECT 6.390 1.665 6.560 1.745 ;
        RECT 7.315 1.740 7.485 5.115 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 9.935 4.710 10.105 4.865 ;
        RECT 9.905 4.535 10.105 4.710 ;
        RECT 9.905 1.915 10.075 4.535 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.420 1.495 6.560 1.665 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.420 0.365 5.590 1.495 ;
        RECT 6.390 0.615 6.560 1.495 ;
        RECT 6.875 1.570 7.485 1.740 ;
        RECT 8.750 1.665 8.920 1.745 ;
        RECT 9.720 1.665 9.890 1.745 ;
        RECT 10.645 1.740 10.815 5.115 ;
        RECT 12.495 1.915 12.665 4.865 ;
        RECT 6.875 0.835 7.045 1.570 ;
        RECT 8.750 1.495 9.890 1.665 ;
        RECT 7.360 0.615 7.530 1.385 ;
        RECT 6.390 0.445 7.530 0.615 ;
        RECT 6.390 0.365 6.560 0.445 ;
        RECT 7.360 0.365 7.530 0.445 ;
        RECT 8.750 0.365 8.920 1.495 ;
        RECT 9.720 0.615 9.890 1.495 ;
        RECT 10.205 1.570 10.815 1.740 ;
        RECT 12.080 1.665 12.250 1.745 ;
        RECT 13.050 1.665 13.220 1.745 ;
        RECT 13.975 1.740 14.145 5.115 ;
        RECT 15.825 1.915 15.995 4.865 ;
        RECT 16.595 4.710 16.765 4.865 ;
        RECT 16.565 4.535 16.765 4.710 ;
        RECT 16.565 1.915 16.735 4.535 ;
        RECT 10.205 0.835 10.375 1.570 ;
        RECT 12.080 1.495 13.220 1.665 ;
        RECT 10.690 0.615 10.860 1.385 ;
        RECT 9.720 0.445 10.860 0.615 ;
        RECT 9.720 0.365 9.890 0.445 ;
        RECT 10.690 0.365 10.860 0.445 ;
        RECT 12.080 0.365 12.250 1.495 ;
        RECT 13.050 0.615 13.220 1.495 ;
        RECT 13.535 1.570 14.145 1.740 ;
        RECT 15.410 1.665 15.580 1.745 ;
        RECT 16.380 1.665 16.550 1.745 ;
        RECT 17.305 1.740 17.475 5.115 ;
        RECT 19.155 1.915 19.325 4.865 ;
        RECT 19.925 4.710 20.095 4.865 ;
        RECT 19.895 4.535 20.095 4.710 ;
        RECT 19.895 1.915 20.065 4.535 ;
        RECT 13.535 0.835 13.705 1.570 ;
        RECT 15.410 1.495 16.550 1.665 ;
        RECT 14.020 0.615 14.190 1.385 ;
        RECT 13.050 0.445 14.190 0.615 ;
        RECT 13.050 0.365 13.220 0.445 ;
        RECT 14.020 0.365 14.190 0.445 ;
        RECT 15.410 0.365 15.580 1.495 ;
        RECT 16.380 0.615 16.550 1.495 ;
        RECT 16.865 1.570 17.475 1.740 ;
        RECT 18.740 1.665 18.910 1.745 ;
        RECT 19.710 1.665 19.880 1.745 ;
        RECT 20.635 1.740 20.805 5.115 ;
        RECT 22.905 5.240 23.075 7.020 ;
        RECT 23.785 5.240 23.955 7.020 ;
        RECT 24.665 5.240 24.835 7.020 ;
        RECT 27.415 5.285 27.585 7.020 ;
        RECT 28.295 5.285 28.465 7.020 ;
        RECT 30.745 5.285 30.915 7.020 ;
        RECT 31.625 5.285 31.795 7.020 ;
        RECT 34.075 5.285 34.245 7.020 ;
        RECT 34.955 5.285 35.125 7.020 ;
        RECT 37.405 5.285 37.575 7.020 ;
        RECT 38.285 5.285 38.455 7.020 ;
        RECT 40.735 5.285 40.905 7.020 ;
        RECT 41.615 5.285 41.785 7.020 ;
        RECT 22.905 5.070 25.615 5.240 ;
        RECT 27.415 5.115 28.945 5.285 ;
        RECT 30.745 5.115 32.275 5.285 ;
        RECT 34.075 5.115 35.605 5.285 ;
        RECT 37.405 5.115 38.935 5.285 ;
        RECT 40.735 5.115 42.265 5.285 ;
        RECT 22.485 1.915 22.655 4.865 ;
        RECT 24.705 1.915 24.875 4.865 ;
        RECT 16.865 0.835 17.035 1.570 ;
        RECT 18.740 1.495 19.880 1.665 ;
        RECT 17.350 0.615 17.520 1.385 ;
        RECT 16.380 0.445 17.520 0.615 ;
        RECT 16.380 0.365 16.550 0.445 ;
        RECT 17.350 0.365 17.520 0.445 ;
        RECT 18.740 0.365 18.910 1.495 ;
        RECT 19.710 0.615 19.880 1.495 ;
        RECT 20.195 1.570 20.805 1.740 ;
        RECT 21.965 1.675 22.135 1.755 ;
        RECT 22.935 1.675 23.105 1.755 ;
        RECT 23.905 1.675 24.075 1.755 ;
        RECT 20.195 0.835 20.365 1.570 ;
        RECT 21.965 1.505 24.075 1.675 ;
        RECT 20.680 0.615 20.850 1.385 ;
        RECT 19.710 0.445 20.850 0.615 ;
        RECT 19.710 0.365 19.880 0.445 ;
        RECT 20.680 0.365 20.850 0.445 ;
        RECT 21.965 0.375 22.135 1.505 ;
        RECT 22.935 0.625 23.105 1.505 ;
        RECT 23.905 1.425 24.075 1.505 ;
        RECT 23.425 1.080 23.595 1.160 ;
        RECT 24.475 1.080 24.645 1.755 ;
        RECT 25.445 1.750 25.615 5.070 ;
        RECT 27.295 1.915 27.465 4.865 ;
        RECT 23.425 0.910 24.645 1.080 ;
        RECT 23.425 0.830 23.595 0.910 ;
        RECT 23.905 0.625 24.075 0.705 ;
        RECT 22.935 0.455 24.075 0.625 ;
        RECT 22.935 0.375 23.105 0.455 ;
        RECT 23.905 0.375 24.075 0.455 ;
        RECT 24.475 0.625 24.645 0.910 ;
        RECT 24.960 1.580 25.615 1.750 ;
        RECT 26.880 1.665 27.050 1.745 ;
        RECT 27.850 1.665 28.020 1.745 ;
        RECT 28.775 1.740 28.945 5.115 ;
        RECT 30.625 1.915 30.795 4.865 ;
        RECT 31.395 4.710 31.565 4.865 ;
        RECT 31.365 4.535 31.565 4.710 ;
        RECT 31.365 1.915 31.535 4.535 ;
        RECT 24.960 0.845 25.130 1.580 ;
        RECT 26.880 1.495 28.020 1.665 ;
        RECT 25.445 0.625 25.615 1.395 ;
        RECT 24.475 0.455 25.615 0.625 ;
        RECT 24.475 0.375 24.645 0.455 ;
        RECT 25.445 0.375 25.615 0.455 ;
        RECT 26.880 0.365 27.050 1.495 ;
        RECT 27.850 0.615 28.020 1.495 ;
        RECT 28.335 1.570 28.945 1.740 ;
        RECT 30.210 1.665 30.380 1.745 ;
        RECT 31.180 1.665 31.350 1.745 ;
        RECT 32.105 1.740 32.275 5.115 ;
        RECT 33.955 1.915 34.125 4.865 ;
        RECT 28.335 0.835 28.505 1.570 ;
        RECT 30.210 1.495 31.350 1.665 ;
        RECT 28.820 0.615 28.990 1.385 ;
        RECT 27.850 0.445 28.990 0.615 ;
        RECT 27.850 0.365 28.020 0.445 ;
        RECT 28.820 0.365 28.990 0.445 ;
        RECT 30.210 0.365 30.380 1.495 ;
        RECT 31.180 0.615 31.350 1.495 ;
        RECT 31.665 1.570 32.275 1.740 ;
        RECT 33.540 1.665 33.710 1.745 ;
        RECT 34.510 1.665 34.680 1.745 ;
        RECT 35.435 1.740 35.605 5.115 ;
        RECT 37.285 1.915 37.455 4.865 ;
        RECT 38.055 4.710 38.225 4.865 ;
        RECT 38.025 4.535 38.225 4.710 ;
        RECT 38.025 1.915 38.195 4.535 ;
        RECT 31.665 0.835 31.835 1.570 ;
        RECT 33.540 1.495 34.680 1.665 ;
        RECT 32.150 0.615 32.320 1.385 ;
        RECT 31.180 0.445 32.320 0.615 ;
        RECT 31.180 0.365 31.350 0.445 ;
        RECT 32.150 0.365 32.320 0.445 ;
        RECT 33.540 0.365 33.710 1.495 ;
        RECT 34.510 0.615 34.680 1.495 ;
        RECT 34.995 1.570 35.605 1.740 ;
        RECT 36.870 1.665 37.040 1.745 ;
        RECT 37.840 1.665 38.010 1.745 ;
        RECT 38.765 1.740 38.935 5.115 ;
        RECT 40.615 1.915 40.785 4.865 ;
        RECT 41.385 4.710 41.555 4.865 ;
        RECT 41.355 4.535 41.555 4.710 ;
        RECT 41.355 1.915 41.525 4.535 ;
        RECT 34.995 0.835 35.165 1.570 ;
        RECT 36.870 1.495 38.010 1.665 ;
        RECT 35.480 0.615 35.650 1.385 ;
        RECT 34.510 0.445 35.650 0.615 ;
        RECT 34.510 0.365 34.680 0.445 ;
        RECT 35.480 0.365 35.650 0.445 ;
        RECT 36.870 0.365 37.040 1.495 ;
        RECT 37.840 0.615 38.010 1.495 ;
        RECT 38.325 1.570 38.935 1.740 ;
        RECT 40.200 1.665 40.370 1.745 ;
        RECT 41.170 1.665 41.340 1.745 ;
        RECT 42.095 1.740 42.265 5.115 ;
        RECT 44.365 5.240 44.535 7.020 ;
        RECT 45.245 5.240 45.415 7.020 ;
        RECT 46.125 5.240 46.295 7.020 ;
        RECT 48.875 5.285 49.045 7.020 ;
        RECT 49.755 5.285 49.925 7.020 ;
        RECT 52.205 5.285 52.375 7.020 ;
        RECT 53.085 5.285 53.255 7.020 ;
        RECT 55.535 5.285 55.705 7.020 ;
        RECT 56.415 5.285 56.585 7.020 ;
        RECT 58.865 5.285 59.035 7.020 ;
        RECT 59.745 5.285 59.915 7.020 ;
        RECT 62.195 5.285 62.365 7.020 ;
        RECT 63.075 5.285 63.245 7.020 ;
        RECT 65.525 6.825 65.705 6.995 ;
        RECT 65.525 5.295 65.695 6.825 ;
        RECT 66.405 5.295 66.575 6.995 ;
        RECT 44.365 5.070 47.075 5.240 ;
        RECT 48.875 5.115 50.405 5.285 ;
        RECT 52.205 5.115 53.735 5.285 ;
        RECT 55.535 5.115 57.065 5.285 ;
        RECT 58.865 5.115 60.395 5.285 ;
        RECT 62.195 5.115 63.725 5.285 ;
        RECT 65.525 5.125 66.575 5.295 ;
        RECT 43.945 1.915 44.115 4.865 ;
        RECT 46.165 1.915 46.335 4.865 ;
        RECT 38.325 0.835 38.495 1.570 ;
        RECT 40.200 1.495 41.340 1.665 ;
        RECT 38.810 0.615 38.980 1.385 ;
        RECT 37.840 0.445 38.980 0.615 ;
        RECT 37.840 0.365 38.010 0.445 ;
        RECT 38.810 0.365 38.980 0.445 ;
        RECT 40.200 0.365 40.370 1.495 ;
        RECT 41.170 0.615 41.340 1.495 ;
        RECT 41.655 1.570 42.265 1.740 ;
        RECT 43.425 1.675 43.595 1.755 ;
        RECT 44.395 1.675 44.565 1.755 ;
        RECT 45.365 1.675 45.535 1.755 ;
        RECT 41.655 0.835 41.825 1.570 ;
        RECT 43.425 1.505 45.535 1.675 ;
        RECT 42.140 0.615 42.310 1.385 ;
        RECT 41.170 0.445 42.310 0.615 ;
        RECT 41.170 0.365 41.340 0.445 ;
        RECT 42.140 0.365 42.310 0.445 ;
        RECT 43.425 0.375 43.595 1.505 ;
        RECT 44.395 0.625 44.565 1.505 ;
        RECT 45.365 1.425 45.535 1.505 ;
        RECT 44.885 1.080 45.055 1.160 ;
        RECT 45.935 1.080 46.105 1.755 ;
        RECT 46.905 1.750 47.075 5.070 ;
        RECT 48.755 1.915 48.925 4.865 ;
        RECT 44.885 0.910 46.105 1.080 ;
        RECT 44.885 0.830 45.055 0.910 ;
        RECT 45.365 0.625 45.535 0.705 ;
        RECT 44.395 0.455 45.535 0.625 ;
        RECT 44.395 0.375 44.565 0.455 ;
        RECT 45.365 0.375 45.535 0.455 ;
        RECT 45.935 0.625 46.105 0.910 ;
        RECT 46.420 1.580 47.075 1.750 ;
        RECT 48.340 1.665 48.510 1.745 ;
        RECT 49.310 1.665 49.480 1.745 ;
        RECT 50.235 1.740 50.405 5.115 ;
        RECT 52.085 1.915 52.255 4.865 ;
        RECT 52.855 4.710 53.025 4.865 ;
        RECT 52.825 4.535 53.025 4.710 ;
        RECT 52.825 1.915 52.995 4.535 ;
        RECT 46.420 0.845 46.590 1.580 ;
        RECT 48.340 1.495 49.480 1.665 ;
        RECT 46.905 0.625 47.075 1.395 ;
        RECT 45.935 0.455 47.075 0.625 ;
        RECT 45.935 0.375 46.105 0.455 ;
        RECT 46.905 0.375 47.075 0.455 ;
        RECT 48.340 0.365 48.510 1.495 ;
        RECT 49.310 0.615 49.480 1.495 ;
        RECT 49.795 1.570 50.405 1.740 ;
        RECT 51.670 1.665 51.840 1.745 ;
        RECT 52.640 1.665 52.810 1.745 ;
        RECT 53.565 1.740 53.735 5.115 ;
        RECT 55.415 1.915 55.585 4.865 ;
        RECT 49.795 0.835 49.965 1.570 ;
        RECT 51.670 1.495 52.810 1.665 ;
        RECT 50.280 0.615 50.450 1.385 ;
        RECT 49.310 0.445 50.450 0.615 ;
        RECT 49.310 0.365 49.480 0.445 ;
        RECT 50.280 0.365 50.450 0.445 ;
        RECT 51.670 0.365 51.840 1.495 ;
        RECT 52.640 0.615 52.810 1.495 ;
        RECT 53.125 1.570 53.735 1.740 ;
        RECT 55.000 1.665 55.170 1.745 ;
        RECT 55.970 1.665 56.140 1.745 ;
        RECT 56.895 1.740 57.065 5.115 ;
        RECT 58.745 1.915 58.915 4.865 ;
        RECT 59.515 4.710 59.685 4.865 ;
        RECT 59.485 4.535 59.685 4.710 ;
        RECT 59.485 1.915 59.655 4.535 ;
        RECT 53.125 0.835 53.295 1.570 ;
        RECT 55.000 1.495 56.140 1.665 ;
        RECT 53.610 0.615 53.780 1.385 ;
        RECT 52.640 0.445 53.780 0.615 ;
        RECT 52.640 0.365 52.810 0.445 ;
        RECT 53.610 0.365 53.780 0.445 ;
        RECT 55.000 0.365 55.170 1.495 ;
        RECT 55.970 0.615 56.140 1.495 ;
        RECT 56.455 1.570 57.065 1.740 ;
        RECT 58.330 1.665 58.500 1.745 ;
        RECT 59.300 1.665 59.470 1.745 ;
        RECT 60.225 1.740 60.395 5.115 ;
        RECT 62.075 1.915 62.245 4.865 ;
        RECT 62.845 4.710 63.015 4.865 ;
        RECT 62.815 4.535 63.015 4.710 ;
        RECT 62.815 1.915 62.985 4.535 ;
        RECT 56.455 0.835 56.625 1.570 ;
        RECT 58.330 1.495 59.470 1.665 ;
        RECT 56.940 0.615 57.110 1.385 ;
        RECT 55.970 0.445 57.110 0.615 ;
        RECT 55.970 0.365 56.140 0.445 ;
        RECT 56.940 0.365 57.110 0.445 ;
        RECT 58.330 0.365 58.500 1.495 ;
        RECT 59.300 0.615 59.470 1.495 ;
        RECT 59.785 1.570 60.395 1.740 ;
        RECT 61.660 1.665 61.830 1.745 ;
        RECT 62.630 1.665 62.800 1.745 ;
        RECT 63.555 1.740 63.725 5.115 ;
        RECT 66.405 5.045 66.575 5.125 ;
        RECT 68.405 6.825 70.335 6.995 ;
        RECT 68.405 5.045 68.575 6.825 ;
        RECT 68.845 5.295 69.015 6.565 ;
        RECT 69.285 5.555 69.455 6.825 ;
        RECT 69.725 5.295 69.895 6.565 ;
        RECT 70.165 5.375 70.335 6.825 ;
        RECT 71.745 6.825 73.675 6.995 ;
        RECT 68.845 5.125 69.895 5.295 ;
        RECT 69.725 5.045 69.895 5.125 ;
        RECT 71.745 5.045 71.915 6.825 ;
        RECT 72.185 5.295 72.355 6.565 ;
        RECT 72.625 5.555 72.795 6.825 ;
        RECT 73.065 5.295 73.235 6.565 ;
        RECT 73.505 5.555 73.675 6.825 ;
        RECT 72.185 5.125 73.715 5.295 ;
        RECT 65.035 1.915 65.205 4.870 ;
        RECT 66.185 4.710 66.355 4.870 ;
        RECT 66.145 4.540 66.355 4.710 ;
        RECT 66.145 1.915 66.315 4.540 ;
        RECT 68.735 1.915 68.905 4.870 ;
        RECT 70.215 1.915 70.385 4.870 ;
        RECT 71.695 1.915 71.865 4.870 ;
        RECT 72.805 4.540 72.995 4.870 ;
        RECT 72.805 1.915 72.975 4.540 ;
        RECT 59.785 0.835 59.955 1.570 ;
        RECT 61.660 1.495 62.800 1.665 ;
        RECT 60.270 0.615 60.440 1.385 ;
        RECT 59.300 0.445 60.440 0.615 ;
        RECT 59.300 0.365 59.470 0.445 ;
        RECT 60.270 0.365 60.440 0.445 ;
        RECT 61.660 0.365 61.830 1.495 ;
        RECT 62.630 0.615 62.800 1.495 ;
        RECT 63.115 1.570 63.725 1.740 ;
        RECT 64.990 1.665 65.160 1.745 ;
        RECT 65.960 1.665 66.130 1.745 ;
        RECT 63.115 0.835 63.285 1.570 ;
        RECT 64.990 1.495 66.130 1.665 ;
        RECT 63.600 0.615 63.770 1.385 ;
        RECT 62.630 0.445 63.770 0.615 ;
        RECT 62.630 0.365 62.800 0.445 ;
        RECT 63.600 0.365 63.770 0.445 ;
        RECT 64.990 0.365 65.160 1.495 ;
        RECT 65.960 0.615 66.130 1.495 ;
        RECT 66.445 1.170 66.615 1.345 ;
        RECT 66.440 1.015 66.615 1.170 ;
        RECT 66.440 0.835 66.610 1.015 ;
        RECT 66.930 0.615 67.100 1.745 ;
        RECT 65.960 0.445 67.100 0.615 ;
        RECT 65.960 0.365 66.130 0.445 ;
        RECT 66.930 0.365 67.100 0.445 ;
        RECT 68.320 1.665 68.490 1.745 ;
        RECT 69.290 1.665 69.460 1.745 ;
        RECT 68.320 1.495 69.460 1.665 ;
        RECT 68.320 0.365 68.490 1.495 ;
        RECT 69.290 0.615 69.460 1.495 ;
        RECT 69.775 0.835 69.945 1.345 ;
        RECT 70.260 0.615 70.430 1.745 ;
        RECT 69.290 0.445 70.430 0.615 ;
        RECT 69.290 0.365 69.460 0.445 ;
        RECT 70.260 0.365 70.430 0.445 ;
        RECT 71.650 1.665 71.820 1.745 ;
        RECT 72.620 1.665 72.790 1.745 ;
        RECT 73.545 1.730 73.715 5.125 ;
        RECT 75.025 1.920 75.195 4.865 ;
        RECT 75.400 4.665 75.570 7.020 ;
        RECT 75.400 4.495 75.935 4.665 ;
        RECT 75.765 2.165 75.935 4.495 ;
        RECT 75.395 1.995 75.935 2.165 ;
        RECT 71.650 1.495 72.790 1.665 ;
        RECT 71.650 0.365 71.820 1.495 ;
        RECT 72.620 0.615 72.790 1.495 ;
        RECT 73.105 1.560 73.715 1.730 ;
        RECT 73.105 0.835 73.275 1.560 ;
        RECT 73.590 0.615 73.760 1.390 ;
        RECT 75.395 0.840 75.565 1.995 ;
        RECT 72.620 0.445 73.760 0.615 ;
        RECT 72.620 0.365 72.790 0.445 ;
        RECT 73.590 0.365 73.760 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 7.315 3.245 7.485 3.415 ;
        RECT 9.165 3.245 9.335 3.415 ;
        RECT 9.905 3.985 10.075 4.155 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 12.495 3.245 12.665 3.415 ;
        RECT 13.975 3.985 14.145 4.155 ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 16.565 2.875 16.735 3.045 ;
        RECT 17.305 3.615 17.475 3.785 ;
        RECT 19.155 3.615 19.325 3.785 ;
        RECT 19.895 3.985 20.065 4.155 ;
        RECT 20.635 2.875 20.805 3.045 ;
        RECT 22.485 3.985 22.655 4.155 ;
        RECT 24.705 3.245 24.875 3.415 ;
        RECT 25.445 3.615 25.615 3.785 ;
        RECT 27.295 3.615 27.465 3.785 ;
        RECT 28.775 3.245 28.945 3.415 ;
        RECT 30.625 3.245 30.795 3.415 ;
        RECT 31.365 3.985 31.535 4.155 ;
        RECT 32.105 3.245 32.275 3.415 ;
        RECT 33.955 3.245 34.125 3.415 ;
        RECT 35.435 3.985 35.605 4.155 ;
        RECT 37.285 3.615 37.455 3.785 ;
        RECT 38.025 2.135 38.195 2.305 ;
        RECT 38.765 3.615 38.935 3.785 ;
        RECT 40.615 3.615 40.785 3.785 ;
        RECT 41.355 3.985 41.525 4.155 ;
        RECT 66.405 5.125 66.575 5.295 ;
        RECT 42.095 2.135 42.265 2.305 ;
        RECT 43.945 3.985 44.115 4.155 ;
        RECT 46.165 3.245 46.335 3.415 ;
        RECT 46.905 3.615 47.075 3.785 ;
        RECT 48.755 3.615 48.925 3.785 ;
        RECT 50.235 3.245 50.405 3.415 ;
        RECT 52.085 3.245 52.255 3.415 ;
        RECT 52.825 3.985 52.995 4.155 ;
        RECT 53.565 3.245 53.735 3.415 ;
        RECT 55.415 3.245 55.585 3.415 ;
        RECT 56.895 3.985 57.065 4.155 ;
        RECT 58.745 3.615 58.915 3.785 ;
        RECT 59.485 3.615 59.655 3.785 ;
        RECT 60.225 4.355 60.395 4.525 ;
        RECT 62.075 4.355 62.245 4.525 ;
        RECT 62.815 3.985 62.985 4.155 ;
        RECT 68.405 5.125 68.575 5.295 ;
        RECT 69.725 5.125 69.895 5.295 ;
        RECT 71.745 5.125 71.915 5.295 ;
        RECT 63.555 3.615 63.725 3.785 ;
        RECT 65.035 4.355 65.205 4.525 ;
        RECT 65.035 3.615 65.205 3.785 ;
        RECT 66.145 3.985 66.315 4.155 ;
        RECT 66.145 2.135 66.315 2.305 ;
        RECT 68.735 4.355 68.905 4.525 ;
        RECT 70.215 2.875 70.385 3.045 ;
        RECT 70.215 1.995 70.385 2.165 ;
        RECT 71.695 1.995 71.865 2.165 ;
        RECT 72.805 3.985 72.975 4.155 ;
        RECT 73.545 3.985 73.715 4.155 ;
        RECT 66.445 1.095 66.615 1.265 ;
        RECT 69.775 1.095 69.945 1.265 ;
        RECT 75.025 3.985 75.195 4.155 ;
        RECT 73.105 1.095 73.275 1.265 ;
      LAYER met1 ;
        RECT 66.375 5.295 66.605 5.325 ;
        RECT 68.375 5.295 68.605 5.325 ;
        RECT 69.695 5.295 69.925 5.325 ;
        RECT 71.715 5.295 71.945 5.325 ;
        RECT 66.345 5.125 68.635 5.295 ;
        RECT 69.665 5.125 71.975 5.295 ;
        RECT 66.375 5.095 66.605 5.125 ;
        RECT 68.375 5.095 68.605 5.125 ;
        RECT 69.695 5.095 69.925 5.125 ;
        RECT 71.715 5.095 71.945 5.125 ;
        RECT 60.195 4.525 60.425 4.555 ;
        RECT 62.045 4.525 62.275 4.555 ;
        RECT 65.005 4.525 65.235 4.555 ;
        RECT 68.705 4.525 68.935 4.555 ;
        RECT 60.165 4.355 62.305 4.525 ;
        RECT 64.975 4.355 68.965 4.525 ;
        RECT 60.195 4.325 60.425 4.355 ;
        RECT 62.045 4.325 62.275 4.355 ;
        RECT 65.005 4.325 65.235 4.355 ;
        RECT 68.705 4.325 68.935 4.355 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 9.875 4.155 10.105 4.185 ;
        RECT 13.945 4.155 14.175 4.185 ;
        RECT 19.865 4.155 20.095 4.185 ;
        RECT 22.455 4.155 22.685 4.185 ;
        RECT 31.335 4.155 31.565 4.185 ;
        RECT 35.405 4.155 35.635 4.185 ;
        RECT 41.325 4.155 41.555 4.185 ;
        RECT 43.915 4.155 44.145 4.185 ;
        RECT 52.795 4.155 53.025 4.185 ;
        RECT 56.865 4.155 57.095 4.185 ;
        RECT 62.785 4.155 63.015 4.185 ;
        RECT 66.115 4.155 66.345 4.185 ;
        RECT 72.775 4.155 73.005 4.185 ;
        RECT 73.515 4.155 73.745 4.185 ;
        RECT 74.995 4.155 75.225 4.185 ;
        RECT 0.965 3.985 20.125 4.155 ;
        RECT 22.425 3.985 41.585 4.155 ;
        RECT 43.885 3.985 63.045 4.155 ;
        RECT 66.085 3.985 73.035 4.155 ;
        RECT 73.485 3.985 75.255 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 9.875 3.955 10.105 3.985 ;
        RECT 13.945 3.955 14.175 3.985 ;
        RECT 19.865 3.955 20.095 3.985 ;
        RECT 22.455 3.955 22.685 3.985 ;
        RECT 31.335 3.955 31.565 3.985 ;
        RECT 35.405 3.955 35.635 3.985 ;
        RECT 41.325 3.955 41.555 3.985 ;
        RECT 43.915 3.955 44.145 3.985 ;
        RECT 52.795 3.955 53.025 3.985 ;
        RECT 56.865 3.955 57.095 3.985 ;
        RECT 62.785 3.955 63.015 3.985 ;
        RECT 66.115 3.955 66.345 3.985 ;
        RECT 72.775 3.955 73.005 3.985 ;
        RECT 73.515 3.955 73.745 3.985 ;
        RECT 74.995 3.955 75.225 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 17.275 3.785 17.505 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 25.415 3.785 25.645 3.815 ;
        RECT 27.265 3.785 27.495 3.815 ;
        RECT 37.255 3.785 37.485 3.815 ;
        RECT 38.735 3.785 38.965 3.815 ;
        RECT 40.585 3.785 40.815 3.815 ;
        RECT 46.875 3.785 47.105 3.815 ;
        RECT 48.725 3.785 48.955 3.815 ;
        RECT 58.715 3.785 58.945 3.815 ;
        RECT 59.455 3.785 59.685 3.815 ;
        RECT 63.525 3.785 63.755 3.815 ;
        RECT 65.005 3.785 65.235 3.815 ;
        RECT 3.925 3.615 16.055 3.785 ;
        RECT 17.245 3.615 19.385 3.785 ;
        RECT 25.385 3.615 37.515 3.785 ;
        RECT 38.705 3.615 40.845 3.785 ;
        RECT 46.845 3.615 58.975 3.785 ;
        RECT 59.425 3.615 65.265 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 17.275 3.585 17.505 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
        RECT 25.415 3.585 25.645 3.615 ;
        RECT 27.265 3.585 27.495 3.615 ;
        RECT 37.255 3.585 37.485 3.615 ;
        RECT 38.735 3.585 38.965 3.615 ;
        RECT 40.585 3.585 40.815 3.615 ;
        RECT 46.875 3.585 47.105 3.615 ;
        RECT 48.725 3.585 48.955 3.615 ;
        RECT 58.715 3.585 58.945 3.615 ;
        RECT 59.455 3.585 59.685 3.615 ;
        RECT 63.525 3.585 63.755 3.615 ;
        RECT 65.005 3.585 65.235 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 7.285 3.415 7.515 3.445 ;
        RECT 9.135 3.415 9.365 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.465 3.415 12.695 3.445 ;
        RECT 24.675 3.415 24.905 3.445 ;
        RECT 28.745 3.415 28.975 3.445 ;
        RECT 30.595 3.415 30.825 3.445 ;
        RECT 32.075 3.415 32.305 3.445 ;
        RECT 33.925 3.415 34.155 3.445 ;
        RECT 46.135 3.415 46.365 3.445 ;
        RECT 50.205 3.415 50.435 3.445 ;
        RECT 52.055 3.415 52.285 3.445 ;
        RECT 53.535 3.415 53.765 3.445 ;
        RECT 55.385 3.415 55.615 3.445 ;
        RECT 3.185 3.245 9.395 3.415 ;
        RECT 10.585 3.245 12.725 3.415 ;
        RECT 24.645 3.245 30.855 3.415 ;
        RECT 32.045 3.245 34.185 3.415 ;
        RECT 46.105 3.245 52.315 3.415 ;
        RECT 53.505 3.245 55.645 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 7.285 3.215 7.515 3.245 ;
        RECT 9.135 3.215 9.365 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.465 3.215 12.695 3.245 ;
        RECT 24.675 3.215 24.905 3.245 ;
        RECT 28.745 3.215 28.975 3.245 ;
        RECT 30.595 3.215 30.825 3.245 ;
        RECT 32.075 3.215 32.305 3.245 ;
        RECT 33.925 3.215 34.155 3.245 ;
        RECT 46.135 3.215 46.365 3.245 ;
        RECT 50.205 3.215 50.435 3.245 ;
        RECT 52.055 3.215 52.285 3.245 ;
        RECT 53.535 3.215 53.765 3.245 ;
        RECT 55.385 3.215 55.615 3.245 ;
        RECT 16.535 3.045 16.765 3.075 ;
        RECT 20.605 3.045 20.835 3.075 ;
        RECT 70.185 3.045 70.415 3.075 ;
        RECT 16.505 2.875 70.445 3.045 ;
        RECT 16.535 2.845 16.765 2.875 ;
        RECT 20.605 2.845 20.835 2.875 ;
        RECT 70.185 2.845 70.415 2.875 ;
        RECT 37.995 2.305 38.225 2.335 ;
        RECT 42.065 2.305 42.295 2.335 ;
        RECT 66.115 2.305 66.345 2.335 ;
        RECT 37.965 2.135 66.375 2.305 ;
        RECT 70.185 2.165 70.415 2.195 ;
        RECT 71.665 2.165 71.895 2.195 ;
        RECT 37.995 2.105 38.225 2.135 ;
        RECT 42.065 2.105 42.295 2.135 ;
        RECT 66.115 2.105 66.345 2.135 ;
        RECT 70.155 1.995 71.925 2.165 ;
        RECT 70.185 1.965 70.415 1.995 ;
        RECT 71.665 1.965 71.895 1.995 ;
        RECT 66.415 1.265 66.645 1.295 ;
        RECT 69.745 1.265 69.975 1.295 ;
        RECT 73.075 1.265 73.305 1.295 ;
        RECT 66.385 1.095 73.335 1.265 ;
        RECT 66.415 1.065 66.645 1.095 ;
        RECT 69.745 1.065 69.975 1.095 ;
        RECT 73.075 1.065 73.305 1.095 ;
  END
END TMRDFFQX1






MACRO TMRDFFRNQNX1
  CLASS CORE ;
  FOREIGN TMRDFFRNQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 87.690 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN D
    ANTENNAGATEAREA 3.044550 ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 32.845 1.915 33.015 4.865 ;
        RECT 58.745 1.915 58.915 4.865 ;
      LAYER mcon ;
        RECT 6.945 2.505 7.115 2.675 ;
        RECT 32.845 2.505 33.015 2.675 ;
        RECT 58.745 2.505 58.915 2.675 ;
      LAYER met1 ;
        RECT 6.915 2.675 7.145 2.705 ;
        RECT 32.815 2.675 33.045 2.705 ;
        RECT 58.715 2.675 58.945 2.705 ;
        RECT 6.885 2.505 59.095 2.675 ;
        RECT 6.915 2.475 7.145 2.505 ;
        RECT 32.815 2.475 33.045 2.505 ;
        RECT 58.715 2.475 58.945 2.505 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 15.085 1.915 15.255 4.865 ;
        RECT 28.035 1.915 28.205 4.865 ;
        RECT 40.985 1.915 41.155 4.865 ;
        RECT 53.935 1.915 54.105 4.865 ;
        RECT 66.885 1.915 67.055 4.865 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 15.085 4.355 15.255 4.525 ;
        RECT 28.035 4.355 28.205 4.525 ;
        RECT 40.985 4.355 41.155 4.525 ;
        RECT 53.935 4.355 54.105 4.525 ;
        RECT 66.885 4.355 67.055 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 15.055 4.525 15.285 4.555 ;
        RECT 28.005 4.525 28.235 4.555 ;
        RECT 40.955 4.525 41.185 4.555 ;
        RECT 53.905 4.525 54.135 4.555 ;
        RECT 66.855 4.525 67.085 4.555 ;
        RECT 2.075 4.355 67.115 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 15.055 4.325 15.285 4.355 ;
        RECT 28.005 4.325 28.235 4.355 ;
        RECT 40.955 4.325 41.185 4.355 ;
        RECT 53.905 4.325 54.135 4.355 ;
        RECT 66.855 4.325 67.085 4.355 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 9.208050 ;
    PORT
      LAYER li1 ;
        RECT 8.055 1.915 8.225 4.865 ;
        RECT 16.195 1.915 16.365 4.865 ;
        RECT 19.895 1.915 20.065 4.865 ;
        RECT 33.955 1.915 34.125 4.865 ;
        RECT 42.095 1.915 42.265 4.865 ;
        RECT 45.795 1.915 45.965 4.865 ;
        RECT 59.855 1.915 60.025 4.865 ;
        RECT 67.995 1.915 68.165 4.865 ;
        RECT 71.695 1.915 71.865 4.865 ;
      LAYER mcon ;
        RECT 8.055 2.135 8.225 2.305 ;
        RECT 16.195 2.135 16.365 2.305 ;
        RECT 19.895 2.135 20.065 2.305 ;
        RECT 33.955 2.135 34.125 2.305 ;
        RECT 42.095 2.135 42.265 2.305 ;
        RECT 45.795 2.135 45.965 2.305 ;
        RECT 59.855 2.135 60.025 2.305 ;
        RECT 67.995 2.135 68.165 2.305 ;
        RECT 71.695 2.135 71.865 2.305 ;
      LAYER met1 ;
        RECT 8.025 2.305 8.255 2.335 ;
        RECT 16.165 2.305 16.395 2.335 ;
        RECT 19.865 2.305 20.095 2.335 ;
        RECT 33.925 2.305 34.155 2.335 ;
        RECT 42.065 2.305 42.295 2.335 ;
        RECT 45.765 2.305 45.995 2.335 ;
        RECT 59.825 2.305 60.055 2.335 ;
        RECT 67.965 2.305 68.195 2.335 ;
        RECT 71.665 2.305 71.895 2.335 ;
        RECT 7.995 2.135 71.925 2.305 ;
        RECT 8.025 2.105 8.255 2.135 ;
        RECT 16.165 2.105 16.395 2.135 ;
        RECT 19.865 2.105 20.095 2.135 ;
        RECT 33.925 2.105 34.155 2.135 ;
        RECT 42.065 2.105 42.295 2.135 ;
        RECT 45.765 2.105 45.995 2.135 ;
        RECT 59.825 2.105 60.055 2.135 ;
        RECT 67.965 2.105 68.195 2.135 ;
        RECT 71.665 2.105 71.895 2.135 ;
    END
  END RN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 88.125 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 87.860 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.325 5.135 10.495 7.230 ;
        RECT 11.205 5.555 11.375 7.230 ;
        RECT 12.085 5.555 12.255 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.955 5.215 14.125 7.230 ;
        RECT 14.835 5.555 15.005 7.230 ;
        RECT 15.715 5.555 15.885 7.230 ;
        RECT 16.595 5.555 16.765 7.230 ;
        RECT 17.590 4.110 17.930 7.230 ;
        RECT 18.765 5.215 18.935 7.230 ;
        RECT 19.645 5.555 19.815 7.230 ;
        RECT 20.525 5.555 20.695 7.230 ;
        RECT 21.405 5.555 21.575 7.230 ;
        RECT 22.400 4.110 22.740 7.230 ;
        RECT 23.275 5.135 23.445 7.230 ;
        RECT 24.155 5.555 24.325 7.230 ;
        RECT 25.035 5.555 25.205 7.230 ;
        RECT 25.730 4.110 26.070 7.230 ;
        RECT 26.905 5.215 27.075 7.230 ;
        RECT 27.785 5.555 27.955 7.230 ;
        RECT 28.665 5.555 28.835 7.230 ;
        RECT 29.545 5.555 29.715 7.230 ;
        RECT 30.540 4.110 30.880 7.230 ;
        RECT 31.715 5.215 31.885 7.230 ;
        RECT 32.595 5.555 32.765 7.230 ;
        RECT 33.475 5.555 33.645 7.230 ;
        RECT 34.355 5.555 34.525 7.230 ;
        RECT 35.350 4.110 35.690 7.230 ;
        RECT 36.225 5.135 36.395 7.230 ;
        RECT 37.105 5.555 37.275 7.230 ;
        RECT 37.985 5.555 38.155 7.230 ;
        RECT 38.680 4.110 39.020 7.230 ;
        RECT 39.855 5.215 40.025 7.230 ;
        RECT 40.735 5.555 40.905 7.230 ;
        RECT 41.615 5.555 41.785 7.230 ;
        RECT 42.495 5.555 42.665 7.230 ;
        RECT 43.490 4.110 43.830 7.230 ;
        RECT 44.665 5.215 44.835 7.230 ;
        RECT 45.545 5.555 45.715 7.230 ;
        RECT 46.425 5.555 46.595 7.230 ;
        RECT 47.305 5.555 47.475 7.230 ;
        RECT 48.300 4.110 48.640 7.230 ;
        RECT 49.175 5.135 49.345 7.230 ;
        RECT 50.055 5.555 50.225 7.230 ;
        RECT 50.935 5.555 51.105 7.230 ;
        RECT 51.630 4.110 51.970 7.230 ;
        RECT 52.805 5.215 52.975 7.230 ;
        RECT 53.685 5.555 53.855 7.230 ;
        RECT 54.565 5.555 54.735 7.230 ;
        RECT 55.445 5.555 55.615 7.230 ;
        RECT 56.440 4.110 56.780 7.230 ;
        RECT 57.615 5.215 57.785 7.230 ;
        RECT 58.495 5.555 58.665 7.230 ;
        RECT 59.375 5.555 59.545 7.230 ;
        RECT 60.255 5.555 60.425 7.230 ;
        RECT 61.250 4.110 61.590 7.230 ;
        RECT 62.125 5.135 62.295 7.230 ;
        RECT 63.005 5.555 63.175 7.230 ;
        RECT 63.885 5.555 64.055 7.230 ;
        RECT 64.580 4.110 64.920 7.230 ;
        RECT 65.755 5.215 65.925 7.230 ;
        RECT 66.635 5.555 66.805 7.230 ;
        RECT 67.515 5.555 67.685 7.230 ;
        RECT 68.395 5.555 68.565 7.230 ;
        RECT 69.390 4.110 69.730 7.230 ;
        RECT 70.565 5.215 70.735 7.230 ;
        RECT 71.445 5.555 71.615 7.230 ;
        RECT 72.325 5.555 72.495 7.230 ;
        RECT 73.205 5.555 73.375 7.230 ;
        RECT 74.200 4.110 74.540 7.230 ;
        RECT 75.075 5.135 75.245 7.230 ;
        RECT 75.955 5.555 76.125 7.230 ;
        RECT 76.835 5.555 77.005 7.230 ;
        RECT 77.530 4.110 77.870 7.230 ;
        RECT 78.405 5.125 78.575 7.230 ;
        RECT 79.285 5.555 79.455 7.230 ;
        RECT 80.165 5.125 80.335 7.230 ;
        RECT 80.860 4.110 81.200 7.230 ;
        RECT 84.190 4.110 84.530 7.230 ;
        RECT 87.520 4.110 87.860 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.515 7.315 29.685 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 32.845 7.315 33.015 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.175 7.315 36.345 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.505 7.315 39.675 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.615 7.315 40.785 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 42.835 7.315 43.005 7.485 ;
        RECT 43.205 7.315 43.375 7.485 ;
        RECT 43.945 7.315 44.115 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 47.645 7.315 47.815 7.485 ;
        RECT 48.015 7.315 48.185 7.485 ;
        RECT 48.755 7.315 48.925 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 50.975 7.315 51.145 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 52.085 7.315 52.255 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 52.825 7.315 52.995 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.305 7.315 54.475 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.895 7.315 57.065 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 57.635 7.315 57.805 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 60.965 7.315 61.135 7.485 ;
        RECT 61.705 7.315 61.875 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.445 7.315 62.615 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.295 7.315 64.465 7.485 ;
        RECT 65.035 7.315 65.205 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.255 7.315 67.425 7.485 ;
        RECT 67.625 7.315 67.795 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.365 7.315 68.535 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 70.955 7.315 71.125 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.065 7.315 72.235 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.175 7.315 73.345 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
        RECT 74.655 7.315 74.825 7.485 ;
        RECT 75.025 7.315 75.195 7.485 ;
        RECT 75.395 7.315 75.565 7.485 ;
        RECT 75.765 7.315 75.935 7.485 ;
        RECT 76.135 7.315 76.305 7.485 ;
        RECT 76.505 7.315 76.675 7.485 ;
        RECT 76.875 7.315 77.045 7.485 ;
        RECT 77.245 7.315 77.415 7.485 ;
        RECT 77.985 7.315 78.155 7.485 ;
        RECT 78.355 7.315 78.525 7.485 ;
        RECT 78.725 7.315 78.895 7.485 ;
        RECT 79.095 7.315 79.265 7.485 ;
        RECT 79.465 7.315 79.635 7.485 ;
        RECT 79.835 7.315 80.005 7.485 ;
        RECT 80.205 7.315 80.375 7.485 ;
        RECT 80.575 7.315 80.745 7.485 ;
        RECT 81.315 7.315 81.485 7.485 ;
        RECT 81.685 7.315 81.855 7.485 ;
        RECT 82.055 7.315 82.225 7.485 ;
        RECT 82.425 7.315 82.595 7.485 ;
        RECT 82.795 7.315 82.965 7.485 ;
        RECT 83.165 7.315 83.335 7.485 ;
        RECT 83.535 7.315 83.705 7.485 ;
        RECT 83.905 7.315 84.075 7.485 ;
        RECT 84.645 7.315 84.815 7.485 ;
        RECT 85.015 7.315 85.185 7.485 ;
        RECT 85.385 7.315 85.555 7.485 ;
        RECT 85.755 7.315 85.925 7.485 ;
        RECT 86.125 7.315 86.295 7.485 ;
        RECT 86.495 7.315 86.665 7.485 ;
        RECT 86.865 7.315 87.035 7.485 ;
        RECT 87.235 7.315 87.405 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 87.860 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 87.860 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.715 0.170 10.885 1.120 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 13.940 0.170 14.110 1.130 ;
        RECT 17.590 0.170 17.930 2.720 ;
        RECT 18.750 0.170 18.920 1.130 ;
        RECT 22.400 0.170 22.740 2.720 ;
        RECT 23.665 0.170 23.835 1.120 ;
        RECT 25.730 0.170 26.070 2.720 ;
        RECT 26.890 0.170 27.060 1.130 ;
        RECT 30.540 0.170 30.880 2.720 ;
        RECT 31.700 0.170 31.870 1.130 ;
        RECT 35.350 0.170 35.690 2.720 ;
        RECT 36.615 0.170 36.785 1.120 ;
        RECT 38.680 0.170 39.020 2.720 ;
        RECT 39.840 0.170 40.010 1.130 ;
        RECT 43.490 0.170 43.830 2.720 ;
        RECT 44.650 0.170 44.820 1.130 ;
        RECT 48.300 0.170 48.640 2.720 ;
        RECT 49.565 0.170 49.735 1.120 ;
        RECT 51.630 0.170 51.970 2.720 ;
        RECT 52.790 0.170 52.960 1.130 ;
        RECT 56.440 0.170 56.780 2.720 ;
        RECT 57.600 0.170 57.770 1.130 ;
        RECT 61.250 0.170 61.590 2.720 ;
        RECT 62.515 0.170 62.685 1.120 ;
        RECT 64.580 0.170 64.920 2.720 ;
        RECT 65.740 0.170 65.910 1.130 ;
        RECT 69.390 0.170 69.730 2.720 ;
        RECT 70.550 0.170 70.720 1.130 ;
        RECT 74.200 0.170 74.540 2.720 ;
        RECT 75.465 0.170 75.635 1.120 ;
        RECT 77.530 0.170 77.870 2.720 ;
        RECT 78.795 0.170 78.965 1.120 ;
        RECT 80.860 0.170 81.200 2.720 ;
        RECT 82.125 0.170 82.295 1.120 ;
        RECT 84.190 0.170 84.530 2.720 ;
        RECT 85.455 0.170 85.625 1.120 ;
        RECT 87.520 0.170 87.860 2.720 ;
        RECT -0.170 -0.170 87.860 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.515 -0.085 29.685 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 32.845 -0.085 33.015 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.175 -0.085 36.345 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.505 -0.085 39.675 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.615 -0.085 40.785 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 42.835 -0.085 43.005 0.085 ;
        RECT 43.205 -0.085 43.375 0.085 ;
        RECT 43.945 -0.085 44.115 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 47.645 -0.085 47.815 0.085 ;
        RECT 48.015 -0.085 48.185 0.085 ;
        RECT 48.755 -0.085 48.925 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 50.975 -0.085 51.145 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 52.085 -0.085 52.255 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 52.825 -0.085 52.995 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.305 -0.085 54.475 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.895 -0.085 57.065 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 57.635 -0.085 57.805 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 60.965 -0.085 61.135 0.085 ;
        RECT 61.705 -0.085 61.875 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.445 -0.085 62.615 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.295 -0.085 64.465 0.085 ;
        RECT 65.035 -0.085 65.205 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.255 -0.085 67.425 0.085 ;
        RECT 67.625 -0.085 67.795 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.365 -0.085 68.535 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 70.955 -0.085 71.125 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.065 -0.085 72.235 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.175 -0.085 73.345 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
        RECT 74.655 -0.085 74.825 0.085 ;
        RECT 75.025 -0.085 75.195 0.085 ;
        RECT 75.395 -0.085 75.565 0.085 ;
        RECT 75.765 -0.085 75.935 0.085 ;
        RECT 76.135 -0.085 76.305 0.085 ;
        RECT 76.505 -0.085 76.675 0.085 ;
        RECT 76.875 -0.085 77.045 0.085 ;
        RECT 77.245 -0.085 77.415 0.085 ;
        RECT 77.985 -0.085 78.155 0.085 ;
        RECT 78.355 -0.085 78.525 0.085 ;
        RECT 78.725 -0.085 78.895 0.085 ;
        RECT 79.095 -0.085 79.265 0.085 ;
        RECT 79.465 -0.085 79.635 0.085 ;
        RECT 79.835 -0.085 80.005 0.085 ;
        RECT 80.205 -0.085 80.375 0.085 ;
        RECT 80.575 -0.085 80.745 0.085 ;
        RECT 81.315 -0.085 81.485 0.085 ;
        RECT 81.685 -0.085 81.855 0.085 ;
        RECT 82.055 -0.085 82.225 0.085 ;
        RECT 82.425 -0.085 82.595 0.085 ;
        RECT 82.795 -0.085 82.965 0.085 ;
        RECT 83.165 -0.085 83.335 0.085 ;
        RECT 83.535 -0.085 83.705 0.085 ;
        RECT 83.905 -0.085 84.075 0.085 ;
        RECT 84.645 -0.085 84.815 0.085 ;
        RECT 85.015 -0.085 85.185 0.085 ;
        RECT 85.385 -0.085 85.555 0.085 ;
        RECT 85.755 -0.085 85.925 0.085 ;
        RECT 86.125 -0.085 86.295 0.085 ;
        RECT 86.495 -0.085 86.665 0.085 ;
        RECT 86.865 -0.085 87.035 0.085 ;
        RECT 87.235 -0.085 87.405 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 87.860 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 10.765 5.285 10.935 7.020 ;
        RECT 11.645 5.285 11.815 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 10.765 5.115 12.295 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 11.415 4.710 11.585 4.865 ;
        RECT 11.385 4.535 11.585 4.710 ;
        RECT 11.385 1.915 11.555 4.535 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.230 1.665 10.400 1.745 ;
        RECT 11.200 1.665 11.370 1.745 ;
        RECT 12.125 1.740 12.295 5.115 ;
        RECT 14.395 5.240 14.565 7.020 ;
        RECT 15.275 5.240 15.445 7.020 ;
        RECT 16.155 5.240 16.325 7.020 ;
        RECT 19.205 5.240 19.375 7.020 ;
        RECT 20.085 5.240 20.255 7.020 ;
        RECT 20.965 5.240 21.135 7.020 ;
        RECT 23.715 5.285 23.885 7.020 ;
        RECT 24.595 5.285 24.765 7.020 ;
        RECT 14.395 5.070 17.105 5.240 ;
        RECT 19.205 5.070 21.915 5.240 ;
        RECT 23.715 5.115 25.245 5.285 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.230 1.495 11.370 1.665 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.230 0.365 10.400 1.495 ;
        RECT 11.200 0.615 11.370 1.495 ;
        RECT 11.685 1.570 12.295 1.740 ;
        RECT 13.455 1.675 13.625 1.755 ;
        RECT 14.425 1.675 14.595 1.755 ;
        RECT 15.395 1.675 15.565 1.755 ;
        RECT 11.685 0.835 11.855 1.570 ;
        RECT 13.455 1.505 15.565 1.675 ;
        RECT 12.170 0.615 12.340 1.385 ;
        RECT 11.200 0.445 12.340 0.615 ;
        RECT 11.200 0.365 11.370 0.445 ;
        RECT 12.170 0.365 12.340 0.445 ;
        RECT 13.455 0.375 13.625 1.505 ;
        RECT 14.425 0.625 14.595 1.505 ;
        RECT 15.395 1.425 15.565 1.505 ;
        RECT 14.915 1.080 15.085 1.160 ;
        RECT 15.965 1.080 16.135 1.755 ;
        RECT 16.935 1.750 17.105 5.070 ;
        RECT 18.785 1.915 18.955 4.865 ;
        RECT 21.005 1.915 21.175 4.865 ;
        RECT 14.915 0.910 16.135 1.080 ;
        RECT 14.915 0.830 15.085 0.910 ;
        RECT 15.395 0.625 15.565 0.705 ;
        RECT 14.425 0.455 15.565 0.625 ;
        RECT 14.425 0.375 14.595 0.455 ;
        RECT 15.395 0.375 15.565 0.455 ;
        RECT 15.965 0.625 16.135 0.910 ;
        RECT 16.450 1.580 17.105 1.750 ;
        RECT 18.265 1.675 18.435 1.755 ;
        RECT 19.235 1.675 19.405 1.755 ;
        RECT 20.205 1.675 20.375 1.755 ;
        RECT 16.450 0.845 16.620 1.580 ;
        RECT 18.265 1.505 20.375 1.675 ;
        RECT 16.935 0.625 17.105 1.395 ;
        RECT 15.965 0.455 17.105 0.625 ;
        RECT 15.965 0.375 16.135 0.455 ;
        RECT 16.935 0.375 17.105 0.455 ;
        RECT 18.265 0.375 18.435 1.505 ;
        RECT 19.235 0.625 19.405 1.505 ;
        RECT 20.205 1.425 20.375 1.505 ;
        RECT 19.725 1.080 19.895 1.160 ;
        RECT 20.775 1.080 20.945 1.755 ;
        RECT 21.745 1.750 21.915 5.070 ;
        RECT 23.595 1.915 23.765 4.865 ;
        RECT 24.365 4.710 24.535 4.865 ;
        RECT 24.335 4.535 24.535 4.710 ;
        RECT 24.335 1.915 24.505 4.535 ;
        RECT 19.725 0.910 20.945 1.080 ;
        RECT 19.725 0.830 19.895 0.910 ;
        RECT 20.205 0.625 20.375 0.705 ;
        RECT 19.235 0.455 20.375 0.625 ;
        RECT 19.235 0.375 19.405 0.455 ;
        RECT 20.205 0.375 20.375 0.455 ;
        RECT 20.775 0.625 20.945 0.910 ;
        RECT 21.260 1.580 21.915 1.750 ;
        RECT 23.180 1.665 23.350 1.745 ;
        RECT 24.150 1.665 24.320 1.745 ;
        RECT 25.075 1.740 25.245 5.115 ;
        RECT 27.345 5.240 27.515 7.020 ;
        RECT 28.225 5.240 28.395 7.020 ;
        RECT 29.105 5.240 29.275 7.020 ;
        RECT 32.155 5.240 32.325 7.020 ;
        RECT 33.035 5.240 33.205 7.020 ;
        RECT 33.915 5.240 34.085 7.020 ;
        RECT 36.665 5.285 36.835 7.020 ;
        RECT 37.545 5.285 37.715 7.020 ;
        RECT 27.345 5.070 30.055 5.240 ;
        RECT 32.155 5.070 34.865 5.240 ;
        RECT 36.665 5.115 38.195 5.285 ;
        RECT 26.925 1.915 27.095 4.865 ;
        RECT 29.145 1.915 29.315 4.865 ;
        RECT 21.260 0.845 21.430 1.580 ;
        RECT 23.180 1.495 24.320 1.665 ;
        RECT 21.745 0.625 21.915 1.395 ;
        RECT 20.775 0.455 21.915 0.625 ;
        RECT 20.775 0.375 20.945 0.455 ;
        RECT 21.745 0.375 21.915 0.455 ;
        RECT 23.180 0.365 23.350 1.495 ;
        RECT 24.150 0.615 24.320 1.495 ;
        RECT 24.635 1.570 25.245 1.740 ;
        RECT 26.405 1.675 26.575 1.755 ;
        RECT 27.375 1.675 27.545 1.755 ;
        RECT 28.345 1.675 28.515 1.755 ;
        RECT 24.635 0.835 24.805 1.570 ;
        RECT 26.405 1.505 28.515 1.675 ;
        RECT 25.120 0.615 25.290 1.385 ;
        RECT 24.150 0.445 25.290 0.615 ;
        RECT 24.150 0.365 24.320 0.445 ;
        RECT 25.120 0.365 25.290 0.445 ;
        RECT 26.405 0.375 26.575 1.505 ;
        RECT 27.375 0.625 27.545 1.505 ;
        RECT 28.345 1.425 28.515 1.505 ;
        RECT 27.865 1.080 28.035 1.160 ;
        RECT 28.915 1.080 29.085 1.755 ;
        RECT 29.885 1.750 30.055 5.070 ;
        RECT 31.735 1.915 31.905 4.865 ;
        RECT 27.865 0.910 29.085 1.080 ;
        RECT 27.865 0.830 28.035 0.910 ;
        RECT 28.345 0.625 28.515 0.705 ;
        RECT 27.375 0.455 28.515 0.625 ;
        RECT 27.375 0.375 27.545 0.455 ;
        RECT 28.345 0.375 28.515 0.455 ;
        RECT 28.915 0.625 29.085 0.910 ;
        RECT 29.400 1.580 30.055 1.750 ;
        RECT 31.215 1.675 31.385 1.755 ;
        RECT 32.185 1.675 32.355 1.755 ;
        RECT 33.155 1.675 33.325 1.755 ;
        RECT 29.400 0.845 29.570 1.580 ;
        RECT 31.215 1.505 33.325 1.675 ;
        RECT 29.885 0.625 30.055 1.395 ;
        RECT 28.915 0.455 30.055 0.625 ;
        RECT 28.915 0.375 29.085 0.455 ;
        RECT 29.885 0.375 30.055 0.455 ;
        RECT 31.215 0.375 31.385 1.505 ;
        RECT 32.185 0.625 32.355 1.505 ;
        RECT 33.155 1.425 33.325 1.505 ;
        RECT 32.675 1.080 32.845 1.160 ;
        RECT 33.725 1.080 33.895 1.755 ;
        RECT 34.695 1.750 34.865 5.070 ;
        RECT 36.545 1.915 36.715 4.865 ;
        RECT 37.315 4.710 37.485 4.865 ;
        RECT 37.285 4.535 37.485 4.710 ;
        RECT 37.285 1.915 37.455 4.535 ;
        RECT 32.675 0.910 33.895 1.080 ;
        RECT 32.675 0.830 32.845 0.910 ;
        RECT 33.155 0.625 33.325 0.705 ;
        RECT 32.185 0.455 33.325 0.625 ;
        RECT 32.185 0.375 32.355 0.455 ;
        RECT 33.155 0.375 33.325 0.455 ;
        RECT 33.725 0.625 33.895 0.910 ;
        RECT 34.210 1.580 34.865 1.750 ;
        RECT 36.130 1.665 36.300 1.745 ;
        RECT 37.100 1.665 37.270 1.745 ;
        RECT 38.025 1.740 38.195 5.115 ;
        RECT 40.295 5.240 40.465 7.020 ;
        RECT 41.175 5.240 41.345 7.020 ;
        RECT 42.055 5.240 42.225 7.020 ;
        RECT 45.105 5.240 45.275 7.020 ;
        RECT 45.985 5.240 46.155 7.020 ;
        RECT 46.865 5.240 47.035 7.020 ;
        RECT 49.615 5.285 49.785 7.020 ;
        RECT 50.495 5.285 50.665 7.020 ;
        RECT 40.295 5.070 43.005 5.240 ;
        RECT 45.105 5.070 47.815 5.240 ;
        RECT 49.615 5.115 51.145 5.285 ;
        RECT 39.875 1.915 40.045 4.865 ;
        RECT 34.210 0.845 34.380 1.580 ;
        RECT 36.130 1.495 37.270 1.665 ;
        RECT 34.695 0.625 34.865 1.395 ;
        RECT 33.725 0.455 34.865 0.625 ;
        RECT 33.725 0.375 33.895 0.455 ;
        RECT 34.695 0.375 34.865 0.455 ;
        RECT 36.130 0.365 36.300 1.495 ;
        RECT 37.100 0.615 37.270 1.495 ;
        RECT 37.585 1.570 38.195 1.740 ;
        RECT 39.355 1.675 39.525 1.755 ;
        RECT 40.325 1.675 40.495 1.755 ;
        RECT 41.295 1.675 41.465 1.755 ;
        RECT 37.585 0.835 37.755 1.570 ;
        RECT 39.355 1.505 41.465 1.675 ;
        RECT 38.070 0.615 38.240 1.385 ;
        RECT 37.100 0.445 38.240 0.615 ;
        RECT 37.100 0.365 37.270 0.445 ;
        RECT 38.070 0.365 38.240 0.445 ;
        RECT 39.355 0.375 39.525 1.505 ;
        RECT 40.325 0.625 40.495 1.505 ;
        RECT 41.295 1.425 41.465 1.505 ;
        RECT 40.815 1.080 40.985 1.160 ;
        RECT 41.865 1.080 42.035 1.755 ;
        RECT 42.835 1.750 43.005 5.070 ;
        RECT 44.685 1.915 44.855 4.865 ;
        RECT 46.905 1.915 47.075 4.865 ;
        RECT 40.815 0.910 42.035 1.080 ;
        RECT 40.815 0.830 40.985 0.910 ;
        RECT 41.295 0.625 41.465 0.705 ;
        RECT 40.325 0.455 41.465 0.625 ;
        RECT 40.325 0.375 40.495 0.455 ;
        RECT 41.295 0.375 41.465 0.455 ;
        RECT 41.865 0.625 42.035 0.910 ;
        RECT 42.350 1.580 43.005 1.750 ;
        RECT 44.165 1.675 44.335 1.755 ;
        RECT 45.135 1.675 45.305 1.755 ;
        RECT 46.105 1.675 46.275 1.755 ;
        RECT 42.350 0.845 42.520 1.580 ;
        RECT 44.165 1.505 46.275 1.675 ;
        RECT 42.835 0.625 43.005 1.395 ;
        RECT 41.865 0.455 43.005 0.625 ;
        RECT 41.865 0.375 42.035 0.455 ;
        RECT 42.835 0.375 43.005 0.455 ;
        RECT 44.165 0.375 44.335 1.505 ;
        RECT 45.135 0.625 45.305 1.505 ;
        RECT 46.105 1.425 46.275 1.505 ;
        RECT 45.625 1.080 45.795 1.160 ;
        RECT 46.675 1.080 46.845 1.755 ;
        RECT 47.645 1.750 47.815 5.070 ;
        RECT 49.495 1.915 49.665 4.865 ;
        RECT 50.265 4.710 50.435 4.865 ;
        RECT 50.235 4.535 50.435 4.710 ;
        RECT 50.235 1.915 50.405 4.535 ;
        RECT 45.625 0.910 46.845 1.080 ;
        RECT 45.625 0.830 45.795 0.910 ;
        RECT 46.105 0.625 46.275 0.705 ;
        RECT 45.135 0.455 46.275 0.625 ;
        RECT 45.135 0.375 45.305 0.455 ;
        RECT 46.105 0.375 46.275 0.455 ;
        RECT 46.675 0.625 46.845 0.910 ;
        RECT 47.160 1.580 47.815 1.750 ;
        RECT 49.080 1.665 49.250 1.745 ;
        RECT 50.050 1.665 50.220 1.745 ;
        RECT 50.975 1.740 51.145 5.115 ;
        RECT 53.245 5.240 53.415 7.020 ;
        RECT 54.125 5.240 54.295 7.020 ;
        RECT 55.005 5.240 55.175 7.020 ;
        RECT 58.055 5.240 58.225 7.020 ;
        RECT 58.935 5.240 59.105 7.020 ;
        RECT 59.815 5.240 59.985 7.020 ;
        RECT 62.565 5.285 62.735 7.020 ;
        RECT 63.445 5.285 63.615 7.020 ;
        RECT 53.245 5.070 55.955 5.240 ;
        RECT 58.055 5.070 60.765 5.240 ;
        RECT 62.565 5.115 64.095 5.285 ;
        RECT 52.825 1.915 52.995 4.865 ;
        RECT 55.045 1.915 55.215 4.865 ;
        RECT 47.160 0.845 47.330 1.580 ;
        RECT 49.080 1.495 50.220 1.665 ;
        RECT 47.645 0.625 47.815 1.395 ;
        RECT 46.675 0.455 47.815 0.625 ;
        RECT 46.675 0.375 46.845 0.455 ;
        RECT 47.645 0.375 47.815 0.455 ;
        RECT 49.080 0.365 49.250 1.495 ;
        RECT 50.050 0.615 50.220 1.495 ;
        RECT 50.535 1.570 51.145 1.740 ;
        RECT 52.305 1.675 52.475 1.755 ;
        RECT 53.275 1.675 53.445 1.755 ;
        RECT 54.245 1.675 54.415 1.755 ;
        RECT 50.535 0.835 50.705 1.570 ;
        RECT 52.305 1.505 54.415 1.675 ;
        RECT 51.020 0.615 51.190 1.385 ;
        RECT 50.050 0.445 51.190 0.615 ;
        RECT 50.050 0.365 50.220 0.445 ;
        RECT 51.020 0.365 51.190 0.445 ;
        RECT 52.305 0.375 52.475 1.505 ;
        RECT 53.275 0.625 53.445 1.505 ;
        RECT 54.245 1.425 54.415 1.505 ;
        RECT 53.765 1.080 53.935 1.160 ;
        RECT 54.815 1.080 54.985 1.755 ;
        RECT 55.785 1.750 55.955 5.070 ;
        RECT 57.635 1.915 57.805 4.865 ;
        RECT 53.765 0.910 54.985 1.080 ;
        RECT 53.765 0.830 53.935 0.910 ;
        RECT 54.245 0.625 54.415 0.705 ;
        RECT 53.275 0.455 54.415 0.625 ;
        RECT 53.275 0.375 53.445 0.455 ;
        RECT 54.245 0.375 54.415 0.455 ;
        RECT 54.815 0.625 54.985 0.910 ;
        RECT 55.300 1.580 55.955 1.750 ;
        RECT 57.115 1.675 57.285 1.755 ;
        RECT 58.085 1.675 58.255 1.755 ;
        RECT 59.055 1.675 59.225 1.755 ;
        RECT 55.300 0.845 55.470 1.580 ;
        RECT 57.115 1.505 59.225 1.675 ;
        RECT 55.785 0.625 55.955 1.395 ;
        RECT 54.815 0.455 55.955 0.625 ;
        RECT 54.815 0.375 54.985 0.455 ;
        RECT 55.785 0.375 55.955 0.455 ;
        RECT 57.115 0.375 57.285 1.505 ;
        RECT 58.085 0.625 58.255 1.505 ;
        RECT 59.055 1.425 59.225 1.505 ;
        RECT 58.575 1.080 58.745 1.160 ;
        RECT 59.625 1.080 59.795 1.755 ;
        RECT 60.595 1.750 60.765 5.070 ;
        RECT 62.445 1.915 62.615 4.865 ;
        RECT 63.215 4.710 63.385 4.865 ;
        RECT 63.185 4.535 63.385 4.710 ;
        RECT 63.185 1.915 63.355 4.535 ;
        RECT 58.575 0.910 59.795 1.080 ;
        RECT 58.575 0.830 58.745 0.910 ;
        RECT 59.055 0.625 59.225 0.705 ;
        RECT 58.085 0.455 59.225 0.625 ;
        RECT 58.085 0.375 58.255 0.455 ;
        RECT 59.055 0.375 59.225 0.455 ;
        RECT 59.625 0.625 59.795 0.910 ;
        RECT 60.110 1.580 60.765 1.750 ;
        RECT 62.030 1.665 62.200 1.745 ;
        RECT 63.000 1.665 63.170 1.745 ;
        RECT 63.925 1.740 64.095 5.115 ;
        RECT 66.195 5.240 66.365 7.020 ;
        RECT 67.075 5.240 67.245 7.020 ;
        RECT 67.955 5.240 68.125 7.020 ;
        RECT 71.005 5.240 71.175 7.020 ;
        RECT 71.885 5.240 72.055 7.020 ;
        RECT 72.765 5.240 72.935 7.020 ;
        RECT 75.515 5.285 75.685 7.020 ;
        RECT 76.395 5.285 76.565 7.020 ;
        RECT 78.845 6.825 79.025 6.995 ;
        RECT 78.845 5.295 79.015 6.825 ;
        RECT 79.725 5.295 79.895 6.995 ;
        RECT 66.195 5.070 68.905 5.240 ;
        RECT 71.005 5.070 73.715 5.240 ;
        RECT 75.515 5.115 77.045 5.285 ;
        RECT 78.845 5.125 79.895 5.295 ;
        RECT 65.775 1.915 65.945 4.865 ;
        RECT 60.110 0.845 60.280 1.580 ;
        RECT 62.030 1.495 63.170 1.665 ;
        RECT 60.595 0.625 60.765 1.395 ;
        RECT 59.625 0.455 60.765 0.625 ;
        RECT 59.625 0.375 59.795 0.455 ;
        RECT 60.595 0.375 60.765 0.455 ;
        RECT 62.030 0.365 62.200 1.495 ;
        RECT 63.000 0.615 63.170 1.495 ;
        RECT 63.485 1.570 64.095 1.740 ;
        RECT 65.255 1.675 65.425 1.755 ;
        RECT 66.225 1.675 66.395 1.755 ;
        RECT 67.195 1.675 67.365 1.755 ;
        RECT 63.485 0.835 63.655 1.570 ;
        RECT 65.255 1.505 67.365 1.675 ;
        RECT 63.970 0.615 64.140 1.385 ;
        RECT 63.000 0.445 64.140 0.615 ;
        RECT 63.000 0.365 63.170 0.445 ;
        RECT 63.970 0.365 64.140 0.445 ;
        RECT 65.255 0.375 65.425 1.505 ;
        RECT 66.225 0.625 66.395 1.505 ;
        RECT 67.195 1.425 67.365 1.505 ;
        RECT 66.715 1.080 66.885 1.160 ;
        RECT 67.765 1.080 67.935 1.755 ;
        RECT 68.735 1.750 68.905 5.070 ;
        RECT 70.585 1.915 70.755 4.865 ;
        RECT 72.805 1.915 72.975 4.865 ;
        RECT 66.715 0.910 67.935 1.080 ;
        RECT 66.715 0.830 66.885 0.910 ;
        RECT 67.195 0.625 67.365 0.705 ;
        RECT 66.225 0.455 67.365 0.625 ;
        RECT 66.225 0.375 66.395 0.455 ;
        RECT 67.195 0.375 67.365 0.455 ;
        RECT 67.765 0.625 67.935 0.910 ;
        RECT 68.250 1.580 68.905 1.750 ;
        RECT 70.065 1.675 70.235 1.755 ;
        RECT 71.035 1.675 71.205 1.755 ;
        RECT 72.005 1.675 72.175 1.755 ;
        RECT 68.250 0.845 68.420 1.580 ;
        RECT 70.065 1.505 72.175 1.675 ;
        RECT 68.735 0.625 68.905 1.395 ;
        RECT 67.765 0.455 68.905 0.625 ;
        RECT 67.765 0.375 67.935 0.455 ;
        RECT 68.735 0.375 68.905 0.455 ;
        RECT 70.065 0.375 70.235 1.505 ;
        RECT 71.035 0.625 71.205 1.505 ;
        RECT 72.005 1.425 72.175 1.505 ;
        RECT 71.525 1.080 71.695 1.160 ;
        RECT 72.575 1.080 72.745 1.755 ;
        RECT 73.545 1.750 73.715 5.070 ;
        RECT 75.395 1.915 75.565 4.865 ;
        RECT 76.165 4.710 76.335 4.865 ;
        RECT 76.135 4.535 76.335 4.710 ;
        RECT 76.135 1.915 76.305 4.535 ;
        RECT 71.525 0.910 72.745 1.080 ;
        RECT 71.525 0.830 71.695 0.910 ;
        RECT 72.005 0.625 72.175 0.705 ;
        RECT 71.035 0.455 72.175 0.625 ;
        RECT 71.035 0.375 71.205 0.455 ;
        RECT 72.005 0.375 72.175 0.455 ;
        RECT 72.575 0.625 72.745 0.910 ;
        RECT 73.060 1.580 73.715 1.750 ;
        RECT 74.980 1.665 75.150 1.745 ;
        RECT 75.950 1.665 76.120 1.745 ;
        RECT 76.875 1.740 77.045 5.115 ;
        RECT 79.725 5.045 79.895 5.125 ;
        RECT 81.725 6.825 83.655 6.995 ;
        RECT 81.725 5.045 81.895 6.825 ;
        RECT 82.165 5.295 82.335 6.565 ;
        RECT 82.605 5.555 82.775 6.825 ;
        RECT 83.045 5.295 83.215 6.565 ;
        RECT 83.485 5.375 83.655 6.825 ;
        RECT 85.065 6.825 86.995 6.995 ;
        RECT 82.165 5.125 83.215 5.295 ;
        RECT 83.045 5.045 83.215 5.125 ;
        RECT 85.065 5.045 85.235 6.825 ;
        RECT 85.505 5.295 85.675 6.565 ;
        RECT 85.945 5.555 86.115 6.825 ;
        RECT 86.385 5.295 86.555 6.565 ;
        RECT 86.825 5.555 86.995 6.825 ;
        RECT 85.505 5.125 87.035 5.295 ;
        RECT 78.355 1.915 78.525 4.870 ;
        RECT 79.505 4.710 79.675 4.870 ;
        RECT 79.465 4.540 79.675 4.710 ;
        RECT 79.465 1.915 79.635 4.540 ;
        RECT 82.055 1.915 82.225 4.870 ;
        RECT 83.535 1.915 83.705 4.870 ;
        RECT 85.015 1.915 85.185 4.870 ;
        RECT 86.125 4.540 86.315 4.870 ;
        RECT 86.125 1.915 86.295 4.540 ;
        RECT 73.060 0.845 73.230 1.580 ;
        RECT 74.980 1.495 76.120 1.665 ;
        RECT 73.545 0.625 73.715 1.395 ;
        RECT 72.575 0.455 73.715 0.625 ;
        RECT 72.575 0.375 72.745 0.455 ;
        RECT 73.545 0.375 73.715 0.455 ;
        RECT 74.980 0.365 75.150 1.495 ;
        RECT 75.950 0.615 76.120 1.495 ;
        RECT 76.435 1.570 77.045 1.740 ;
        RECT 78.310 1.665 78.480 1.745 ;
        RECT 79.280 1.665 79.450 1.745 ;
        RECT 76.435 0.835 76.605 1.570 ;
        RECT 78.310 1.495 79.450 1.665 ;
        RECT 76.920 0.615 77.090 1.385 ;
        RECT 75.950 0.445 77.090 0.615 ;
        RECT 75.950 0.365 76.120 0.445 ;
        RECT 76.920 0.365 77.090 0.445 ;
        RECT 78.310 0.365 78.480 1.495 ;
        RECT 79.280 0.615 79.450 1.495 ;
        RECT 79.765 1.170 79.935 1.345 ;
        RECT 79.760 1.015 79.935 1.170 ;
        RECT 79.760 0.835 79.930 1.015 ;
        RECT 80.250 0.615 80.420 1.745 ;
        RECT 79.280 0.445 80.420 0.615 ;
        RECT 79.280 0.365 79.450 0.445 ;
        RECT 80.250 0.365 80.420 0.445 ;
        RECT 81.640 1.665 81.810 1.745 ;
        RECT 82.610 1.665 82.780 1.745 ;
        RECT 81.640 1.495 82.780 1.665 ;
        RECT 81.640 0.365 81.810 1.495 ;
        RECT 82.610 0.615 82.780 1.495 ;
        RECT 83.095 0.835 83.265 1.345 ;
        RECT 83.580 0.615 83.750 1.745 ;
        RECT 82.610 0.445 83.750 0.615 ;
        RECT 82.610 0.365 82.780 0.445 ;
        RECT 83.580 0.365 83.750 0.445 ;
        RECT 84.970 1.665 85.140 1.745 ;
        RECT 85.940 1.665 86.110 1.745 ;
        RECT 86.865 1.730 87.035 5.125 ;
        RECT 84.970 1.495 86.110 1.665 ;
        RECT 84.970 0.365 85.140 1.495 ;
        RECT 85.940 0.615 86.110 1.495 ;
        RECT 86.425 1.560 87.035 1.730 ;
        RECT 86.425 0.835 86.595 1.560 ;
        RECT 86.910 0.615 87.080 1.390 ;
        RECT 85.940 0.445 87.080 0.615 ;
        RECT 85.940 0.365 86.110 0.445 ;
        RECT 86.910 0.365 87.080 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 3.245 12.295 3.415 ;
        RECT 13.975 3.245 14.145 3.415 ;
        RECT 16.935 3.985 17.105 4.155 ;
        RECT 18.785 3.615 18.955 3.785 ;
        RECT 21.005 2.875 21.175 3.045 ;
        RECT 21.745 3.985 21.915 4.155 ;
        RECT 23.595 3.985 23.765 4.155 ;
        RECT 24.335 3.985 24.505 4.155 ;
        RECT 25.075 2.875 25.245 3.045 ;
        RECT 26.925 3.985 27.095 4.155 ;
        RECT 29.145 3.245 29.315 3.415 ;
        RECT 29.885 3.615 30.055 3.785 ;
        RECT 31.735 3.615 31.905 3.785 ;
        RECT 34.695 3.245 34.865 3.415 ;
        RECT 36.545 3.245 36.715 3.415 ;
        RECT 37.285 3.985 37.455 4.155 ;
        RECT 38.025 3.245 38.195 3.415 ;
        RECT 39.875 3.245 40.045 3.415 ;
        RECT 42.835 3.985 43.005 4.155 ;
        RECT 44.685 3.615 44.855 3.785 ;
        RECT 46.905 3.245 47.075 3.415 ;
        RECT 47.645 3.615 47.815 3.785 ;
        RECT 49.495 3.615 49.665 3.785 ;
        RECT 50.235 3.985 50.405 4.155 ;
        RECT 50.975 3.245 51.145 3.415 ;
        RECT 52.825 3.985 52.995 4.155 ;
        RECT 55.045 3.245 55.215 3.415 ;
        RECT 55.785 3.615 55.955 3.785 ;
        RECT 57.635 3.615 57.805 3.785 ;
        RECT 60.595 3.245 60.765 3.415 ;
        RECT 62.445 3.245 62.615 3.415 ;
        RECT 63.185 3.985 63.355 4.155 ;
        RECT 79.725 5.125 79.895 5.295 ;
        RECT 63.925 3.245 64.095 3.415 ;
        RECT 65.775 3.245 65.945 3.415 ;
        RECT 68.735 3.985 68.905 4.155 ;
        RECT 70.585 3.615 70.755 3.785 ;
        RECT 72.805 3.615 72.975 3.785 ;
        RECT 73.545 3.985 73.715 4.155 ;
        RECT 75.395 3.985 75.565 4.155 ;
        RECT 76.135 3.985 76.305 4.155 ;
        RECT 81.725 5.125 81.895 5.295 ;
        RECT 83.045 5.125 83.215 5.295 ;
        RECT 85.065 5.125 85.235 5.295 ;
        RECT 76.875 3.615 77.045 3.785 ;
        RECT 78.355 4.355 78.525 4.525 ;
        RECT 78.355 3.245 78.525 3.415 ;
        RECT 79.465 3.985 79.635 4.155 ;
        RECT 79.465 3.615 79.635 3.785 ;
        RECT 82.055 4.355 82.225 4.525 ;
        RECT 83.535 2.875 83.705 3.045 ;
        RECT 83.535 1.995 83.705 2.165 ;
        RECT 85.015 1.995 85.185 2.165 ;
        RECT 86.125 3.985 86.295 4.155 ;
        RECT 79.765 1.095 79.935 1.265 ;
        RECT 83.095 1.095 83.265 1.265 ;
        RECT 86.425 1.095 86.595 1.265 ;
      LAYER met1 ;
        RECT 79.695 5.295 79.925 5.325 ;
        RECT 81.695 5.295 81.925 5.325 ;
        RECT 83.015 5.295 83.245 5.325 ;
        RECT 85.035 5.295 85.265 5.325 ;
        RECT 79.665 5.125 81.955 5.295 ;
        RECT 82.985 5.125 85.295 5.295 ;
        RECT 79.695 5.095 79.925 5.125 ;
        RECT 81.695 5.095 81.925 5.125 ;
        RECT 83.015 5.095 83.245 5.125 ;
        RECT 85.035 5.095 85.265 5.125 ;
        RECT 78.325 4.525 78.555 4.555 ;
        RECT 82.025 4.525 82.255 4.555 ;
        RECT 78.295 4.355 82.285 4.525 ;
        RECT 78.325 4.325 78.555 4.355 ;
        RECT 82.025 4.325 82.255 4.355 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 16.905 4.155 17.135 4.185 ;
        RECT 21.715 4.155 21.945 4.185 ;
        RECT 23.565 4.155 23.795 4.185 ;
        RECT 24.305 4.155 24.535 4.185 ;
        RECT 26.895 4.155 27.125 4.185 ;
        RECT 37.255 4.155 37.485 4.185 ;
        RECT 42.805 4.155 43.035 4.185 ;
        RECT 50.205 4.155 50.435 4.185 ;
        RECT 52.795 4.155 53.025 4.185 ;
        RECT 63.155 4.155 63.385 4.185 ;
        RECT 68.705 4.155 68.935 4.185 ;
        RECT 73.515 4.155 73.745 4.185 ;
        RECT 75.365 4.155 75.595 4.185 ;
        RECT 76.105 4.155 76.335 4.185 ;
        RECT 79.435 4.155 79.665 4.185 ;
        RECT 86.095 4.155 86.325 4.185 ;
        RECT 0.965 3.985 24.565 4.155 ;
        RECT 26.865 3.985 50.465 4.155 ;
        RECT 52.765 3.985 76.365 4.155 ;
        RECT 79.405 3.985 86.355 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 16.905 3.955 17.135 3.985 ;
        RECT 21.715 3.955 21.945 3.985 ;
        RECT 23.565 3.955 23.795 3.985 ;
        RECT 24.305 3.955 24.535 3.985 ;
        RECT 26.895 3.955 27.125 3.985 ;
        RECT 37.255 3.955 37.485 3.985 ;
        RECT 42.805 3.955 43.035 3.985 ;
        RECT 50.205 3.955 50.435 3.985 ;
        RECT 52.795 3.955 53.025 3.985 ;
        RECT 63.155 3.955 63.385 3.985 ;
        RECT 68.705 3.955 68.935 3.985 ;
        RECT 73.515 3.955 73.745 3.985 ;
        RECT 75.365 3.955 75.595 3.985 ;
        RECT 76.105 3.955 76.335 3.985 ;
        RECT 79.435 3.955 79.665 3.985 ;
        RECT 86.095 3.955 86.325 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 18.755 3.785 18.985 3.815 ;
        RECT 29.855 3.785 30.085 3.815 ;
        RECT 31.705 3.785 31.935 3.815 ;
        RECT 44.655 3.785 44.885 3.815 ;
        RECT 47.615 3.785 47.845 3.815 ;
        RECT 49.465 3.785 49.695 3.815 ;
        RECT 55.755 3.785 55.985 3.815 ;
        RECT 57.605 3.785 57.835 3.815 ;
        RECT 70.555 3.785 70.785 3.815 ;
        RECT 72.775 3.785 73.005 3.815 ;
        RECT 76.845 3.785 77.075 3.815 ;
        RECT 79.435 3.785 79.665 3.815 ;
        RECT 3.925 3.615 19.015 3.785 ;
        RECT 29.825 3.615 44.915 3.785 ;
        RECT 47.585 3.615 49.725 3.785 ;
        RECT 55.725 3.615 70.815 3.785 ;
        RECT 72.745 3.615 79.695 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 18.755 3.585 18.985 3.615 ;
        RECT 29.855 3.585 30.085 3.615 ;
        RECT 31.705 3.585 31.935 3.615 ;
        RECT 44.655 3.585 44.885 3.615 ;
        RECT 47.615 3.585 47.845 3.615 ;
        RECT 49.465 3.585 49.695 3.615 ;
        RECT 55.755 3.585 55.985 3.615 ;
        RECT 57.605 3.585 57.835 3.615 ;
        RECT 70.555 3.585 70.785 3.615 ;
        RECT 72.775 3.585 73.005 3.615 ;
        RECT 76.845 3.585 77.075 3.615 ;
        RECT 79.435 3.585 79.665 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 8.765 3.415 8.995 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.095 3.415 12.325 3.445 ;
        RECT 13.945 3.415 14.175 3.445 ;
        RECT 29.115 3.415 29.345 3.445 ;
        RECT 34.665 3.415 34.895 3.445 ;
        RECT 36.515 3.415 36.745 3.445 ;
        RECT 37.995 3.415 38.225 3.445 ;
        RECT 39.845 3.415 40.075 3.445 ;
        RECT 46.875 3.415 47.105 3.445 ;
        RECT 50.945 3.415 51.175 3.445 ;
        RECT 55.015 3.415 55.245 3.445 ;
        RECT 60.565 3.415 60.795 3.445 ;
        RECT 62.415 3.415 62.645 3.445 ;
        RECT 63.895 3.415 64.125 3.445 ;
        RECT 65.745 3.415 65.975 3.445 ;
        RECT 78.325 3.415 78.555 3.445 ;
        RECT 3.185 3.245 10.875 3.415 ;
        RECT 12.065 3.245 14.205 3.415 ;
        RECT 29.085 3.245 36.775 3.415 ;
        RECT 37.965 3.245 40.105 3.415 ;
        RECT 46.845 3.245 78.585 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 8.765 3.215 8.995 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.095 3.215 12.325 3.245 ;
        RECT 13.945 3.215 14.175 3.245 ;
        RECT 29.115 3.215 29.345 3.245 ;
        RECT 34.665 3.215 34.895 3.245 ;
        RECT 36.515 3.215 36.745 3.245 ;
        RECT 37.995 3.215 38.225 3.245 ;
        RECT 39.845 3.215 40.075 3.245 ;
        RECT 46.875 3.215 47.105 3.245 ;
        RECT 50.945 3.215 51.175 3.245 ;
        RECT 55.015 3.215 55.245 3.245 ;
        RECT 60.565 3.215 60.795 3.245 ;
        RECT 62.415 3.215 62.645 3.245 ;
        RECT 63.895 3.215 64.125 3.245 ;
        RECT 65.745 3.215 65.975 3.245 ;
        RECT 78.325 3.215 78.555 3.245 ;
        RECT 20.975 3.045 21.205 3.075 ;
        RECT 25.045 3.045 25.275 3.075 ;
        RECT 83.505 3.045 83.735 3.075 ;
        RECT 20.945 2.875 83.765 3.045 ;
        RECT 20.975 2.845 21.205 2.875 ;
        RECT 25.045 2.845 25.275 2.875 ;
        RECT 83.505 2.845 83.735 2.875 ;
        RECT 83.505 2.165 83.735 2.195 ;
        RECT 84.985 2.165 85.215 2.195 ;
        RECT 83.475 1.995 85.245 2.165 ;
        RECT 83.505 1.965 83.735 1.995 ;
        RECT 84.985 1.965 85.215 1.995 ;
        RECT 79.735 1.265 79.965 1.295 ;
        RECT 83.065 1.265 83.295 1.295 ;
        RECT 86.395 1.265 86.625 1.295 ;
        RECT 79.705 1.095 86.655 1.265 ;
        RECT 79.735 1.065 79.965 1.095 ;
        RECT 83.065 1.065 83.295 1.095 ;
        RECT 86.395 1.065 86.625 1.095 ;
  END
END TMRDFFRNQNX1






MACRO TMRDFFRNQX1
  CLASS CORE ;
  FOREIGN TMRDFFRNQX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 89.910 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN D
    ANTENNAGATEAREA 3.044550 ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 32.845 1.915 33.015 4.865 ;
        RECT 58.745 1.915 58.915 4.865 ;
      LAYER mcon ;
        RECT 6.945 2.505 7.115 2.675 ;
        RECT 32.845 2.505 33.015 2.675 ;
        RECT 58.745 2.505 58.915 2.675 ;
      LAYER met1 ;
        RECT 6.915 2.675 7.145 2.705 ;
        RECT 32.815 2.675 33.045 2.705 ;
        RECT 58.715 2.675 58.945 2.705 ;
        RECT 6.885 2.505 59.095 2.675 ;
        RECT 6.915 2.475 7.145 2.505 ;
        RECT 32.815 2.475 33.045 2.505 ;
        RECT 58.715 2.475 58.945 2.505 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 15.085 1.915 15.255 4.865 ;
        RECT 28.035 1.915 28.205 4.865 ;
        RECT 40.985 1.915 41.155 4.865 ;
        RECT 53.935 1.915 54.105 4.865 ;
        RECT 66.885 1.915 67.055 4.865 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 15.085 4.355 15.255 4.525 ;
        RECT 28.035 4.355 28.205 4.525 ;
        RECT 40.985 4.355 41.155 4.525 ;
        RECT 53.935 4.355 54.105 4.525 ;
        RECT 66.885 4.355 67.055 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 15.055 4.525 15.285 4.555 ;
        RECT 28.005 4.525 28.235 4.555 ;
        RECT 40.955 4.525 41.185 4.555 ;
        RECT 53.905 4.525 54.135 4.555 ;
        RECT 66.855 4.525 67.085 4.555 ;
        RECT 2.075 4.355 67.115 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 15.055 4.325 15.285 4.355 ;
        RECT 28.005 4.325 28.235 4.355 ;
        RECT 40.955 4.325 41.185 4.355 ;
        RECT 53.905 4.325 54.135 4.355 ;
        RECT 66.855 4.325 67.085 4.355 ;
    END
  END CLK
  PIN RN
    ANTENNAGATEAREA 9.208050 ;
    PORT
      LAYER li1 ;
        RECT 8.055 1.915 8.225 4.865 ;
        RECT 16.195 1.915 16.365 4.865 ;
        RECT 19.895 1.915 20.065 4.865 ;
        RECT 33.955 1.915 34.125 4.865 ;
        RECT 42.095 1.915 42.265 4.865 ;
        RECT 45.795 1.915 45.965 4.865 ;
        RECT 59.855 1.915 60.025 4.865 ;
        RECT 67.995 1.915 68.165 4.865 ;
        RECT 71.695 1.915 71.865 4.865 ;
      LAYER mcon ;
        RECT 8.055 2.135 8.225 2.305 ;
        RECT 16.195 2.135 16.365 2.305 ;
        RECT 19.895 2.135 20.065 2.305 ;
        RECT 33.955 2.135 34.125 2.305 ;
        RECT 42.095 2.135 42.265 2.305 ;
        RECT 45.795 2.135 45.965 2.305 ;
        RECT 59.855 2.135 60.025 2.305 ;
        RECT 67.995 2.135 68.165 2.305 ;
        RECT 71.695 2.135 71.865 2.305 ;
      LAYER met1 ;
        RECT 8.025 2.305 8.255 2.335 ;
        RECT 16.165 2.305 16.395 2.335 ;
        RECT 19.865 2.305 20.095 2.335 ;
        RECT 33.925 2.305 34.155 2.335 ;
        RECT 42.065 2.305 42.295 2.335 ;
        RECT 45.765 2.305 45.995 2.335 ;
        RECT 59.825 2.305 60.055 2.335 ;
        RECT 67.965 2.305 68.195 2.335 ;
        RECT 71.665 2.305 71.895 2.335 ;
        RECT 7.995 2.135 71.925 2.305 ;
        RECT 8.025 2.105 8.255 2.135 ;
        RECT 16.165 2.105 16.395 2.135 ;
        RECT 19.865 2.105 20.095 2.135 ;
        RECT 33.925 2.105 34.155 2.135 ;
        RECT 42.065 2.105 42.295 2.135 ;
        RECT 45.765 2.105 45.995 2.135 ;
        RECT 59.825 2.105 60.055 2.135 ;
        RECT 67.965 2.105 68.195 2.135 ;
        RECT 71.665 2.105 71.895 2.135 ;
    END
  END RN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 90.345 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 90.080 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.325 5.135 10.495 7.230 ;
        RECT 11.205 5.555 11.375 7.230 ;
        RECT 12.085 5.555 12.255 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.955 5.215 14.125 7.230 ;
        RECT 14.835 5.555 15.005 7.230 ;
        RECT 15.715 5.555 15.885 7.230 ;
        RECT 16.595 5.555 16.765 7.230 ;
        RECT 17.590 4.110 17.930 7.230 ;
        RECT 18.765 5.215 18.935 7.230 ;
        RECT 19.645 5.555 19.815 7.230 ;
        RECT 20.525 5.555 20.695 7.230 ;
        RECT 21.405 5.555 21.575 7.230 ;
        RECT 22.400 4.110 22.740 7.230 ;
        RECT 23.275 5.135 23.445 7.230 ;
        RECT 24.155 5.555 24.325 7.230 ;
        RECT 25.035 5.555 25.205 7.230 ;
        RECT 25.730 4.110 26.070 7.230 ;
        RECT 26.905 5.215 27.075 7.230 ;
        RECT 27.785 5.555 27.955 7.230 ;
        RECT 28.665 5.555 28.835 7.230 ;
        RECT 29.545 5.555 29.715 7.230 ;
        RECT 30.540 4.110 30.880 7.230 ;
        RECT 31.715 5.215 31.885 7.230 ;
        RECT 32.595 5.555 32.765 7.230 ;
        RECT 33.475 5.555 33.645 7.230 ;
        RECT 34.355 5.555 34.525 7.230 ;
        RECT 35.350 4.110 35.690 7.230 ;
        RECT 36.225 5.135 36.395 7.230 ;
        RECT 37.105 5.555 37.275 7.230 ;
        RECT 37.985 5.555 38.155 7.230 ;
        RECT 38.680 4.110 39.020 7.230 ;
        RECT 39.855 5.215 40.025 7.230 ;
        RECT 40.735 5.555 40.905 7.230 ;
        RECT 41.615 5.555 41.785 7.230 ;
        RECT 42.495 5.555 42.665 7.230 ;
        RECT 43.490 4.110 43.830 7.230 ;
        RECT 44.665 5.215 44.835 7.230 ;
        RECT 45.545 5.555 45.715 7.230 ;
        RECT 46.425 5.555 46.595 7.230 ;
        RECT 47.305 5.555 47.475 7.230 ;
        RECT 48.300 4.110 48.640 7.230 ;
        RECT 49.175 5.135 49.345 7.230 ;
        RECT 50.055 5.555 50.225 7.230 ;
        RECT 50.935 5.555 51.105 7.230 ;
        RECT 51.630 4.110 51.970 7.230 ;
        RECT 52.805 5.215 52.975 7.230 ;
        RECT 53.685 5.555 53.855 7.230 ;
        RECT 54.565 5.555 54.735 7.230 ;
        RECT 55.445 5.555 55.615 7.230 ;
        RECT 56.440 4.110 56.780 7.230 ;
        RECT 57.615 5.215 57.785 7.230 ;
        RECT 58.495 5.555 58.665 7.230 ;
        RECT 59.375 5.555 59.545 7.230 ;
        RECT 60.255 5.555 60.425 7.230 ;
        RECT 61.250 4.110 61.590 7.230 ;
        RECT 62.125 5.135 62.295 7.230 ;
        RECT 63.005 5.555 63.175 7.230 ;
        RECT 63.885 5.555 64.055 7.230 ;
        RECT 64.580 4.110 64.920 7.230 ;
        RECT 65.755 5.215 65.925 7.230 ;
        RECT 66.635 5.555 66.805 7.230 ;
        RECT 67.515 5.555 67.685 7.230 ;
        RECT 68.395 5.555 68.565 7.230 ;
        RECT 69.390 4.110 69.730 7.230 ;
        RECT 70.565 5.215 70.735 7.230 ;
        RECT 71.445 5.555 71.615 7.230 ;
        RECT 72.325 5.555 72.495 7.230 ;
        RECT 73.205 5.555 73.375 7.230 ;
        RECT 74.200 4.110 74.540 7.230 ;
        RECT 75.075 5.135 75.245 7.230 ;
        RECT 75.955 5.555 76.125 7.230 ;
        RECT 76.835 5.555 77.005 7.230 ;
        RECT 77.530 4.110 77.870 7.230 ;
        RECT 78.405 5.125 78.575 7.230 ;
        RECT 79.285 5.555 79.455 7.230 ;
        RECT 80.165 5.125 80.335 7.230 ;
        RECT 80.860 4.110 81.200 7.230 ;
        RECT 84.190 4.110 84.530 7.230 ;
        RECT 87.520 4.110 87.860 7.230 ;
        RECT 88.280 5.185 88.450 7.230 ;
        RECT 89.160 5.185 89.330 7.230 ;
        RECT 89.740 4.110 90.080 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.515 7.315 29.685 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 32.845 7.315 33.015 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.175 7.315 36.345 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.505 7.315 39.675 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.615 7.315 40.785 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 42.835 7.315 43.005 7.485 ;
        RECT 43.205 7.315 43.375 7.485 ;
        RECT 43.945 7.315 44.115 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 47.645 7.315 47.815 7.485 ;
        RECT 48.015 7.315 48.185 7.485 ;
        RECT 48.755 7.315 48.925 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 50.975 7.315 51.145 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 52.085 7.315 52.255 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 52.825 7.315 52.995 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.305 7.315 54.475 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.895 7.315 57.065 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 57.635 7.315 57.805 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 60.965 7.315 61.135 7.485 ;
        RECT 61.705 7.315 61.875 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.445 7.315 62.615 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.295 7.315 64.465 7.485 ;
        RECT 65.035 7.315 65.205 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.255 7.315 67.425 7.485 ;
        RECT 67.625 7.315 67.795 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.365 7.315 68.535 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 70.955 7.315 71.125 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.065 7.315 72.235 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.175 7.315 73.345 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
        RECT 74.655 7.315 74.825 7.485 ;
        RECT 75.025 7.315 75.195 7.485 ;
        RECT 75.395 7.315 75.565 7.485 ;
        RECT 75.765 7.315 75.935 7.485 ;
        RECT 76.135 7.315 76.305 7.485 ;
        RECT 76.505 7.315 76.675 7.485 ;
        RECT 76.875 7.315 77.045 7.485 ;
        RECT 77.245 7.315 77.415 7.485 ;
        RECT 77.985 7.315 78.155 7.485 ;
        RECT 78.355 7.315 78.525 7.485 ;
        RECT 78.725 7.315 78.895 7.485 ;
        RECT 79.095 7.315 79.265 7.485 ;
        RECT 79.465 7.315 79.635 7.485 ;
        RECT 79.835 7.315 80.005 7.485 ;
        RECT 80.205 7.315 80.375 7.485 ;
        RECT 80.575 7.315 80.745 7.485 ;
        RECT 81.315 7.315 81.485 7.485 ;
        RECT 81.685 7.315 81.855 7.485 ;
        RECT 82.055 7.315 82.225 7.485 ;
        RECT 82.425 7.315 82.595 7.485 ;
        RECT 82.795 7.315 82.965 7.485 ;
        RECT 83.165 7.315 83.335 7.485 ;
        RECT 83.535 7.315 83.705 7.485 ;
        RECT 83.905 7.315 84.075 7.485 ;
        RECT 84.645 7.315 84.815 7.485 ;
        RECT 85.015 7.315 85.185 7.485 ;
        RECT 85.385 7.315 85.555 7.485 ;
        RECT 85.755 7.315 85.925 7.485 ;
        RECT 86.125 7.315 86.295 7.485 ;
        RECT 86.495 7.315 86.665 7.485 ;
        RECT 86.865 7.315 87.035 7.485 ;
        RECT 87.235 7.315 87.405 7.485 ;
        RECT 87.975 7.315 88.145 7.485 ;
        RECT 88.345 7.315 88.515 7.485 ;
        RECT 88.715 7.315 88.885 7.485 ;
        RECT 89.085 7.315 89.255 7.485 ;
        RECT 89.455 7.315 89.625 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 90.080 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 90.080 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.715 0.170 10.885 1.120 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 13.940 0.170 14.110 1.130 ;
        RECT 17.590 0.170 17.930 2.720 ;
        RECT 18.750 0.170 18.920 1.130 ;
        RECT 22.400 0.170 22.740 2.720 ;
        RECT 23.665 0.170 23.835 1.120 ;
        RECT 25.730 0.170 26.070 2.720 ;
        RECT 26.890 0.170 27.060 1.130 ;
        RECT 30.540 0.170 30.880 2.720 ;
        RECT 31.700 0.170 31.870 1.130 ;
        RECT 35.350 0.170 35.690 2.720 ;
        RECT 36.615 0.170 36.785 1.120 ;
        RECT 38.680 0.170 39.020 2.720 ;
        RECT 39.840 0.170 40.010 1.130 ;
        RECT 43.490 0.170 43.830 2.720 ;
        RECT 44.650 0.170 44.820 1.130 ;
        RECT 48.300 0.170 48.640 2.720 ;
        RECT 49.565 0.170 49.735 1.120 ;
        RECT 51.630 0.170 51.970 2.720 ;
        RECT 52.790 0.170 52.960 1.130 ;
        RECT 56.440 0.170 56.780 2.720 ;
        RECT 57.600 0.170 57.770 1.130 ;
        RECT 61.250 0.170 61.590 2.720 ;
        RECT 62.515 0.170 62.685 1.120 ;
        RECT 64.580 0.170 64.920 2.720 ;
        RECT 65.740 0.170 65.910 1.130 ;
        RECT 69.390 0.170 69.730 2.720 ;
        RECT 70.550 0.170 70.720 1.130 ;
        RECT 74.200 0.170 74.540 2.720 ;
        RECT 75.465 0.170 75.635 1.120 ;
        RECT 77.530 0.170 77.870 2.720 ;
        RECT 78.795 0.170 78.965 1.120 ;
        RECT 80.860 0.170 81.200 2.720 ;
        RECT 82.125 0.170 82.295 1.120 ;
        RECT 84.190 0.170 84.530 2.720 ;
        RECT 85.455 0.170 85.625 1.120 ;
        RECT 87.520 0.170 87.860 2.720 ;
        RECT 88.235 0.620 88.405 1.750 ;
        RECT 89.205 0.620 89.375 1.750 ;
        RECT 88.235 0.450 89.375 0.620 ;
        RECT 88.235 0.170 88.405 0.450 ;
        RECT 88.720 0.170 88.890 0.450 ;
        RECT 89.205 0.170 89.375 0.450 ;
        RECT 89.740 0.170 90.080 2.720 ;
        RECT -0.170 -0.170 90.080 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.515 -0.085 29.685 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 32.845 -0.085 33.015 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.175 -0.085 36.345 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.505 -0.085 39.675 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.615 -0.085 40.785 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 42.835 -0.085 43.005 0.085 ;
        RECT 43.205 -0.085 43.375 0.085 ;
        RECT 43.945 -0.085 44.115 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 47.645 -0.085 47.815 0.085 ;
        RECT 48.015 -0.085 48.185 0.085 ;
        RECT 48.755 -0.085 48.925 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 50.975 -0.085 51.145 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 52.085 -0.085 52.255 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 52.825 -0.085 52.995 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.305 -0.085 54.475 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.895 -0.085 57.065 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 57.635 -0.085 57.805 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 60.965 -0.085 61.135 0.085 ;
        RECT 61.705 -0.085 61.875 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.445 -0.085 62.615 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.295 -0.085 64.465 0.085 ;
        RECT 65.035 -0.085 65.205 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.255 -0.085 67.425 0.085 ;
        RECT 67.625 -0.085 67.795 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.365 -0.085 68.535 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 70.955 -0.085 71.125 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.065 -0.085 72.235 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.175 -0.085 73.345 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
        RECT 74.655 -0.085 74.825 0.085 ;
        RECT 75.025 -0.085 75.195 0.085 ;
        RECT 75.395 -0.085 75.565 0.085 ;
        RECT 75.765 -0.085 75.935 0.085 ;
        RECT 76.135 -0.085 76.305 0.085 ;
        RECT 76.505 -0.085 76.675 0.085 ;
        RECT 76.875 -0.085 77.045 0.085 ;
        RECT 77.245 -0.085 77.415 0.085 ;
        RECT 77.985 -0.085 78.155 0.085 ;
        RECT 78.355 -0.085 78.525 0.085 ;
        RECT 78.725 -0.085 78.895 0.085 ;
        RECT 79.095 -0.085 79.265 0.085 ;
        RECT 79.465 -0.085 79.635 0.085 ;
        RECT 79.835 -0.085 80.005 0.085 ;
        RECT 80.205 -0.085 80.375 0.085 ;
        RECT 80.575 -0.085 80.745 0.085 ;
        RECT 81.315 -0.085 81.485 0.085 ;
        RECT 81.685 -0.085 81.855 0.085 ;
        RECT 82.055 -0.085 82.225 0.085 ;
        RECT 82.425 -0.085 82.595 0.085 ;
        RECT 82.795 -0.085 82.965 0.085 ;
        RECT 83.165 -0.085 83.335 0.085 ;
        RECT 83.535 -0.085 83.705 0.085 ;
        RECT 83.905 -0.085 84.075 0.085 ;
        RECT 84.645 -0.085 84.815 0.085 ;
        RECT 85.015 -0.085 85.185 0.085 ;
        RECT 85.385 -0.085 85.555 0.085 ;
        RECT 85.755 -0.085 85.925 0.085 ;
        RECT 86.125 -0.085 86.295 0.085 ;
        RECT 86.495 -0.085 86.665 0.085 ;
        RECT 86.865 -0.085 87.035 0.085 ;
        RECT 87.235 -0.085 87.405 0.085 ;
        RECT 87.975 -0.085 88.145 0.085 ;
        RECT 88.345 -0.085 88.515 0.085 ;
        RECT 88.715 -0.085 88.885 0.085 ;
        RECT 89.085 -0.085 89.255 0.085 ;
        RECT 89.455 -0.085 89.625 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 90.080 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 10.765 5.285 10.935 7.020 ;
        RECT 11.645 5.285 11.815 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 10.765 5.115 12.295 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 11.415 4.710 11.585 4.865 ;
        RECT 11.385 4.535 11.585 4.710 ;
        RECT 11.385 1.915 11.555 4.535 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.230 1.665 10.400 1.745 ;
        RECT 11.200 1.665 11.370 1.745 ;
        RECT 12.125 1.740 12.295 5.115 ;
        RECT 14.395 5.240 14.565 7.020 ;
        RECT 15.275 5.240 15.445 7.020 ;
        RECT 16.155 5.240 16.325 7.020 ;
        RECT 19.205 5.240 19.375 7.020 ;
        RECT 20.085 5.240 20.255 7.020 ;
        RECT 20.965 5.240 21.135 7.020 ;
        RECT 23.715 5.285 23.885 7.020 ;
        RECT 24.595 5.285 24.765 7.020 ;
        RECT 14.395 5.070 17.105 5.240 ;
        RECT 19.205 5.070 21.915 5.240 ;
        RECT 23.715 5.115 25.245 5.285 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.230 1.495 11.370 1.665 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.230 0.365 10.400 1.495 ;
        RECT 11.200 0.615 11.370 1.495 ;
        RECT 11.685 1.570 12.295 1.740 ;
        RECT 13.455 1.675 13.625 1.755 ;
        RECT 14.425 1.675 14.595 1.755 ;
        RECT 15.395 1.675 15.565 1.755 ;
        RECT 11.685 0.835 11.855 1.570 ;
        RECT 13.455 1.505 15.565 1.675 ;
        RECT 12.170 0.615 12.340 1.385 ;
        RECT 11.200 0.445 12.340 0.615 ;
        RECT 11.200 0.365 11.370 0.445 ;
        RECT 12.170 0.365 12.340 0.445 ;
        RECT 13.455 0.375 13.625 1.505 ;
        RECT 14.425 0.625 14.595 1.505 ;
        RECT 15.395 1.425 15.565 1.505 ;
        RECT 14.915 1.080 15.085 1.160 ;
        RECT 15.965 1.080 16.135 1.755 ;
        RECT 16.935 1.750 17.105 5.070 ;
        RECT 18.785 1.915 18.955 4.865 ;
        RECT 21.005 1.915 21.175 4.865 ;
        RECT 14.915 0.910 16.135 1.080 ;
        RECT 14.915 0.830 15.085 0.910 ;
        RECT 15.395 0.625 15.565 0.705 ;
        RECT 14.425 0.455 15.565 0.625 ;
        RECT 14.425 0.375 14.595 0.455 ;
        RECT 15.395 0.375 15.565 0.455 ;
        RECT 15.965 0.625 16.135 0.910 ;
        RECT 16.450 1.580 17.105 1.750 ;
        RECT 18.265 1.675 18.435 1.755 ;
        RECT 19.235 1.675 19.405 1.755 ;
        RECT 20.205 1.675 20.375 1.755 ;
        RECT 16.450 0.845 16.620 1.580 ;
        RECT 18.265 1.505 20.375 1.675 ;
        RECT 16.935 0.625 17.105 1.395 ;
        RECT 15.965 0.455 17.105 0.625 ;
        RECT 15.965 0.375 16.135 0.455 ;
        RECT 16.935 0.375 17.105 0.455 ;
        RECT 18.265 0.375 18.435 1.505 ;
        RECT 19.235 0.625 19.405 1.505 ;
        RECT 20.205 1.425 20.375 1.505 ;
        RECT 19.725 1.080 19.895 1.160 ;
        RECT 20.775 1.080 20.945 1.755 ;
        RECT 21.745 1.750 21.915 5.070 ;
        RECT 23.595 1.915 23.765 4.865 ;
        RECT 24.365 4.710 24.535 4.865 ;
        RECT 24.335 4.535 24.535 4.710 ;
        RECT 24.335 1.915 24.505 4.535 ;
        RECT 19.725 0.910 20.945 1.080 ;
        RECT 19.725 0.830 19.895 0.910 ;
        RECT 20.205 0.625 20.375 0.705 ;
        RECT 19.235 0.455 20.375 0.625 ;
        RECT 19.235 0.375 19.405 0.455 ;
        RECT 20.205 0.375 20.375 0.455 ;
        RECT 20.775 0.625 20.945 0.910 ;
        RECT 21.260 1.580 21.915 1.750 ;
        RECT 23.180 1.665 23.350 1.745 ;
        RECT 24.150 1.665 24.320 1.745 ;
        RECT 25.075 1.740 25.245 5.115 ;
        RECT 27.345 5.240 27.515 7.020 ;
        RECT 28.225 5.240 28.395 7.020 ;
        RECT 29.105 5.240 29.275 7.020 ;
        RECT 32.155 5.240 32.325 7.020 ;
        RECT 33.035 5.240 33.205 7.020 ;
        RECT 33.915 5.240 34.085 7.020 ;
        RECT 36.665 5.285 36.835 7.020 ;
        RECT 37.545 5.285 37.715 7.020 ;
        RECT 27.345 5.070 30.055 5.240 ;
        RECT 32.155 5.070 34.865 5.240 ;
        RECT 36.665 5.115 38.195 5.285 ;
        RECT 26.925 1.915 27.095 4.865 ;
        RECT 29.145 1.915 29.315 4.865 ;
        RECT 21.260 0.845 21.430 1.580 ;
        RECT 23.180 1.495 24.320 1.665 ;
        RECT 21.745 0.625 21.915 1.395 ;
        RECT 20.775 0.455 21.915 0.625 ;
        RECT 20.775 0.375 20.945 0.455 ;
        RECT 21.745 0.375 21.915 0.455 ;
        RECT 23.180 0.365 23.350 1.495 ;
        RECT 24.150 0.615 24.320 1.495 ;
        RECT 24.635 1.570 25.245 1.740 ;
        RECT 26.405 1.675 26.575 1.755 ;
        RECT 27.375 1.675 27.545 1.755 ;
        RECT 28.345 1.675 28.515 1.755 ;
        RECT 24.635 0.835 24.805 1.570 ;
        RECT 26.405 1.505 28.515 1.675 ;
        RECT 25.120 0.615 25.290 1.385 ;
        RECT 24.150 0.445 25.290 0.615 ;
        RECT 24.150 0.365 24.320 0.445 ;
        RECT 25.120 0.365 25.290 0.445 ;
        RECT 26.405 0.375 26.575 1.505 ;
        RECT 27.375 0.625 27.545 1.505 ;
        RECT 28.345 1.425 28.515 1.505 ;
        RECT 27.865 1.080 28.035 1.160 ;
        RECT 28.915 1.080 29.085 1.755 ;
        RECT 29.885 1.750 30.055 5.070 ;
        RECT 31.735 1.915 31.905 4.865 ;
        RECT 27.865 0.910 29.085 1.080 ;
        RECT 27.865 0.830 28.035 0.910 ;
        RECT 28.345 0.625 28.515 0.705 ;
        RECT 27.375 0.455 28.515 0.625 ;
        RECT 27.375 0.375 27.545 0.455 ;
        RECT 28.345 0.375 28.515 0.455 ;
        RECT 28.915 0.625 29.085 0.910 ;
        RECT 29.400 1.580 30.055 1.750 ;
        RECT 31.215 1.675 31.385 1.755 ;
        RECT 32.185 1.675 32.355 1.755 ;
        RECT 33.155 1.675 33.325 1.755 ;
        RECT 29.400 0.845 29.570 1.580 ;
        RECT 31.215 1.505 33.325 1.675 ;
        RECT 29.885 0.625 30.055 1.395 ;
        RECT 28.915 0.455 30.055 0.625 ;
        RECT 28.915 0.375 29.085 0.455 ;
        RECT 29.885 0.375 30.055 0.455 ;
        RECT 31.215 0.375 31.385 1.505 ;
        RECT 32.185 0.625 32.355 1.505 ;
        RECT 33.155 1.425 33.325 1.505 ;
        RECT 32.675 1.080 32.845 1.160 ;
        RECT 33.725 1.080 33.895 1.755 ;
        RECT 34.695 1.750 34.865 5.070 ;
        RECT 36.545 1.915 36.715 4.865 ;
        RECT 37.315 4.710 37.485 4.865 ;
        RECT 37.285 4.535 37.485 4.710 ;
        RECT 37.285 1.915 37.455 4.535 ;
        RECT 32.675 0.910 33.895 1.080 ;
        RECT 32.675 0.830 32.845 0.910 ;
        RECT 33.155 0.625 33.325 0.705 ;
        RECT 32.185 0.455 33.325 0.625 ;
        RECT 32.185 0.375 32.355 0.455 ;
        RECT 33.155 0.375 33.325 0.455 ;
        RECT 33.725 0.625 33.895 0.910 ;
        RECT 34.210 1.580 34.865 1.750 ;
        RECT 36.130 1.665 36.300 1.745 ;
        RECT 37.100 1.665 37.270 1.745 ;
        RECT 38.025 1.740 38.195 5.115 ;
        RECT 40.295 5.240 40.465 7.020 ;
        RECT 41.175 5.240 41.345 7.020 ;
        RECT 42.055 5.240 42.225 7.020 ;
        RECT 45.105 5.240 45.275 7.020 ;
        RECT 45.985 5.240 46.155 7.020 ;
        RECT 46.865 5.240 47.035 7.020 ;
        RECT 49.615 5.285 49.785 7.020 ;
        RECT 50.495 5.285 50.665 7.020 ;
        RECT 40.295 5.070 43.005 5.240 ;
        RECT 45.105 5.070 47.815 5.240 ;
        RECT 49.615 5.115 51.145 5.285 ;
        RECT 39.875 1.915 40.045 4.865 ;
        RECT 34.210 0.845 34.380 1.580 ;
        RECT 36.130 1.495 37.270 1.665 ;
        RECT 34.695 0.625 34.865 1.395 ;
        RECT 33.725 0.455 34.865 0.625 ;
        RECT 33.725 0.375 33.895 0.455 ;
        RECT 34.695 0.375 34.865 0.455 ;
        RECT 36.130 0.365 36.300 1.495 ;
        RECT 37.100 0.615 37.270 1.495 ;
        RECT 37.585 1.570 38.195 1.740 ;
        RECT 39.355 1.675 39.525 1.755 ;
        RECT 40.325 1.675 40.495 1.755 ;
        RECT 41.295 1.675 41.465 1.755 ;
        RECT 37.585 0.835 37.755 1.570 ;
        RECT 39.355 1.505 41.465 1.675 ;
        RECT 38.070 0.615 38.240 1.385 ;
        RECT 37.100 0.445 38.240 0.615 ;
        RECT 37.100 0.365 37.270 0.445 ;
        RECT 38.070 0.365 38.240 0.445 ;
        RECT 39.355 0.375 39.525 1.505 ;
        RECT 40.325 0.625 40.495 1.505 ;
        RECT 41.295 1.425 41.465 1.505 ;
        RECT 40.815 1.080 40.985 1.160 ;
        RECT 41.865 1.080 42.035 1.755 ;
        RECT 42.835 1.750 43.005 5.070 ;
        RECT 44.685 1.915 44.855 4.865 ;
        RECT 46.905 1.915 47.075 4.865 ;
        RECT 40.815 0.910 42.035 1.080 ;
        RECT 40.815 0.830 40.985 0.910 ;
        RECT 41.295 0.625 41.465 0.705 ;
        RECT 40.325 0.455 41.465 0.625 ;
        RECT 40.325 0.375 40.495 0.455 ;
        RECT 41.295 0.375 41.465 0.455 ;
        RECT 41.865 0.625 42.035 0.910 ;
        RECT 42.350 1.580 43.005 1.750 ;
        RECT 44.165 1.675 44.335 1.755 ;
        RECT 45.135 1.675 45.305 1.755 ;
        RECT 46.105 1.675 46.275 1.755 ;
        RECT 42.350 0.845 42.520 1.580 ;
        RECT 44.165 1.505 46.275 1.675 ;
        RECT 42.835 0.625 43.005 1.395 ;
        RECT 41.865 0.455 43.005 0.625 ;
        RECT 41.865 0.375 42.035 0.455 ;
        RECT 42.835 0.375 43.005 0.455 ;
        RECT 44.165 0.375 44.335 1.505 ;
        RECT 45.135 0.625 45.305 1.505 ;
        RECT 46.105 1.425 46.275 1.505 ;
        RECT 45.625 1.080 45.795 1.160 ;
        RECT 46.675 1.080 46.845 1.755 ;
        RECT 47.645 1.750 47.815 5.070 ;
        RECT 49.495 1.915 49.665 4.865 ;
        RECT 50.265 4.710 50.435 4.865 ;
        RECT 50.235 4.535 50.435 4.710 ;
        RECT 50.235 1.915 50.405 4.535 ;
        RECT 45.625 0.910 46.845 1.080 ;
        RECT 45.625 0.830 45.795 0.910 ;
        RECT 46.105 0.625 46.275 0.705 ;
        RECT 45.135 0.455 46.275 0.625 ;
        RECT 45.135 0.375 45.305 0.455 ;
        RECT 46.105 0.375 46.275 0.455 ;
        RECT 46.675 0.625 46.845 0.910 ;
        RECT 47.160 1.580 47.815 1.750 ;
        RECT 49.080 1.665 49.250 1.745 ;
        RECT 50.050 1.665 50.220 1.745 ;
        RECT 50.975 1.740 51.145 5.115 ;
        RECT 53.245 5.240 53.415 7.020 ;
        RECT 54.125 5.240 54.295 7.020 ;
        RECT 55.005 5.240 55.175 7.020 ;
        RECT 58.055 5.240 58.225 7.020 ;
        RECT 58.935 5.240 59.105 7.020 ;
        RECT 59.815 5.240 59.985 7.020 ;
        RECT 62.565 5.285 62.735 7.020 ;
        RECT 63.445 5.285 63.615 7.020 ;
        RECT 53.245 5.070 55.955 5.240 ;
        RECT 58.055 5.070 60.765 5.240 ;
        RECT 62.565 5.115 64.095 5.285 ;
        RECT 52.825 1.915 52.995 4.865 ;
        RECT 55.045 1.915 55.215 4.865 ;
        RECT 47.160 0.845 47.330 1.580 ;
        RECT 49.080 1.495 50.220 1.665 ;
        RECT 47.645 0.625 47.815 1.395 ;
        RECT 46.675 0.455 47.815 0.625 ;
        RECT 46.675 0.375 46.845 0.455 ;
        RECT 47.645 0.375 47.815 0.455 ;
        RECT 49.080 0.365 49.250 1.495 ;
        RECT 50.050 0.615 50.220 1.495 ;
        RECT 50.535 1.570 51.145 1.740 ;
        RECT 52.305 1.675 52.475 1.755 ;
        RECT 53.275 1.675 53.445 1.755 ;
        RECT 54.245 1.675 54.415 1.755 ;
        RECT 50.535 0.835 50.705 1.570 ;
        RECT 52.305 1.505 54.415 1.675 ;
        RECT 51.020 0.615 51.190 1.385 ;
        RECT 50.050 0.445 51.190 0.615 ;
        RECT 50.050 0.365 50.220 0.445 ;
        RECT 51.020 0.365 51.190 0.445 ;
        RECT 52.305 0.375 52.475 1.505 ;
        RECT 53.275 0.625 53.445 1.505 ;
        RECT 54.245 1.425 54.415 1.505 ;
        RECT 53.765 1.080 53.935 1.160 ;
        RECT 54.815 1.080 54.985 1.755 ;
        RECT 55.785 1.750 55.955 5.070 ;
        RECT 57.635 1.915 57.805 4.865 ;
        RECT 53.765 0.910 54.985 1.080 ;
        RECT 53.765 0.830 53.935 0.910 ;
        RECT 54.245 0.625 54.415 0.705 ;
        RECT 53.275 0.455 54.415 0.625 ;
        RECT 53.275 0.375 53.445 0.455 ;
        RECT 54.245 0.375 54.415 0.455 ;
        RECT 54.815 0.625 54.985 0.910 ;
        RECT 55.300 1.580 55.955 1.750 ;
        RECT 57.115 1.675 57.285 1.755 ;
        RECT 58.085 1.675 58.255 1.755 ;
        RECT 59.055 1.675 59.225 1.755 ;
        RECT 55.300 0.845 55.470 1.580 ;
        RECT 57.115 1.505 59.225 1.675 ;
        RECT 55.785 0.625 55.955 1.395 ;
        RECT 54.815 0.455 55.955 0.625 ;
        RECT 54.815 0.375 54.985 0.455 ;
        RECT 55.785 0.375 55.955 0.455 ;
        RECT 57.115 0.375 57.285 1.505 ;
        RECT 58.085 0.625 58.255 1.505 ;
        RECT 59.055 1.425 59.225 1.505 ;
        RECT 58.575 1.080 58.745 1.160 ;
        RECT 59.625 1.080 59.795 1.755 ;
        RECT 60.595 1.750 60.765 5.070 ;
        RECT 62.445 1.915 62.615 4.865 ;
        RECT 63.215 4.710 63.385 4.865 ;
        RECT 63.185 4.535 63.385 4.710 ;
        RECT 63.185 1.915 63.355 4.535 ;
        RECT 58.575 0.910 59.795 1.080 ;
        RECT 58.575 0.830 58.745 0.910 ;
        RECT 59.055 0.625 59.225 0.705 ;
        RECT 58.085 0.455 59.225 0.625 ;
        RECT 58.085 0.375 58.255 0.455 ;
        RECT 59.055 0.375 59.225 0.455 ;
        RECT 59.625 0.625 59.795 0.910 ;
        RECT 60.110 1.580 60.765 1.750 ;
        RECT 62.030 1.665 62.200 1.745 ;
        RECT 63.000 1.665 63.170 1.745 ;
        RECT 63.925 1.740 64.095 5.115 ;
        RECT 66.195 5.240 66.365 7.020 ;
        RECT 67.075 5.240 67.245 7.020 ;
        RECT 67.955 5.240 68.125 7.020 ;
        RECT 71.005 5.240 71.175 7.020 ;
        RECT 71.885 5.240 72.055 7.020 ;
        RECT 72.765 5.240 72.935 7.020 ;
        RECT 75.515 5.285 75.685 7.020 ;
        RECT 76.395 5.285 76.565 7.020 ;
        RECT 78.845 6.825 79.025 6.995 ;
        RECT 78.845 5.295 79.015 6.825 ;
        RECT 79.725 5.295 79.895 6.995 ;
        RECT 66.195 5.070 68.905 5.240 ;
        RECT 71.005 5.070 73.715 5.240 ;
        RECT 75.515 5.115 77.045 5.285 ;
        RECT 78.845 5.125 79.895 5.295 ;
        RECT 65.775 1.915 65.945 4.865 ;
        RECT 60.110 0.845 60.280 1.580 ;
        RECT 62.030 1.495 63.170 1.665 ;
        RECT 60.595 0.625 60.765 1.395 ;
        RECT 59.625 0.455 60.765 0.625 ;
        RECT 59.625 0.375 59.795 0.455 ;
        RECT 60.595 0.375 60.765 0.455 ;
        RECT 62.030 0.365 62.200 1.495 ;
        RECT 63.000 0.615 63.170 1.495 ;
        RECT 63.485 1.570 64.095 1.740 ;
        RECT 65.255 1.675 65.425 1.755 ;
        RECT 66.225 1.675 66.395 1.755 ;
        RECT 67.195 1.675 67.365 1.755 ;
        RECT 63.485 0.835 63.655 1.570 ;
        RECT 65.255 1.505 67.365 1.675 ;
        RECT 63.970 0.615 64.140 1.385 ;
        RECT 63.000 0.445 64.140 0.615 ;
        RECT 63.000 0.365 63.170 0.445 ;
        RECT 63.970 0.365 64.140 0.445 ;
        RECT 65.255 0.375 65.425 1.505 ;
        RECT 66.225 0.625 66.395 1.505 ;
        RECT 67.195 1.425 67.365 1.505 ;
        RECT 66.715 1.080 66.885 1.160 ;
        RECT 67.765 1.080 67.935 1.755 ;
        RECT 68.735 1.750 68.905 5.070 ;
        RECT 70.585 1.915 70.755 4.865 ;
        RECT 72.805 1.915 72.975 4.865 ;
        RECT 66.715 0.910 67.935 1.080 ;
        RECT 66.715 0.830 66.885 0.910 ;
        RECT 67.195 0.625 67.365 0.705 ;
        RECT 66.225 0.455 67.365 0.625 ;
        RECT 66.225 0.375 66.395 0.455 ;
        RECT 67.195 0.375 67.365 0.455 ;
        RECT 67.765 0.625 67.935 0.910 ;
        RECT 68.250 1.580 68.905 1.750 ;
        RECT 70.065 1.675 70.235 1.755 ;
        RECT 71.035 1.675 71.205 1.755 ;
        RECT 72.005 1.675 72.175 1.755 ;
        RECT 68.250 0.845 68.420 1.580 ;
        RECT 70.065 1.505 72.175 1.675 ;
        RECT 68.735 0.625 68.905 1.395 ;
        RECT 67.765 0.455 68.905 0.625 ;
        RECT 67.765 0.375 67.935 0.455 ;
        RECT 68.735 0.375 68.905 0.455 ;
        RECT 70.065 0.375 70.235 1.505 ;
        RECT 71.035 0.625 71.205 1.505 ;
        RECT 72.005 1.425 72.175 1.505 ;
        RECT 71.525 1.080 71.695 1.160 ;
        RECT 72.575 1.080 72.745 1.755 ;
        RECT 73.545 1.750 73.715 5.070 ;
        RECT 75.395 1.915 75.565 4.865 ;
        RECT 76.165 4.710 76.335 4.865 ;
        RECT 76.135 4.535 76.335 4.710 ;
        RECT 76.135 1.915 76.305 4.535 ;
        RECT 71.525 0.910 72.745 1.080 ;
        RECT 71.525 0.830 71.695 0.910 ;
        RECT 72.005 0.625 72.175 0.705 ;
        RECT 71.035 0.455 72.175 0.625 ;
        RECT 71.035 0.375 71.205 0.455 ;
        RECT 72.005 0.375 72.175 0.455 ;
        RECT 72.575 0.625 72.745 0.910 ;
        RECT 73.060 1.580 73.715 1.750 ;
        RECT 74.980 1.665 75.150 1.745 ;
        RECT 75.950 1.665 76.120 1.745 ;
        RECT 76.875 1.740 77.045 5.115 ;
        RECT 79.725 5.045 79.895 5.125 ;
        RECT 81.725 6.825 83.655 6.995 ;
        RECT 81.725 5.045 81.895 6.825 ;
        RECT 82.165 5.295 82.335 6.565 ;
        RECT 82.605 5.555 82.775 6.825 ;
        RECT 83.045 5.295 83.215 6.565 ;
        RECT 83.485 5.375 83.655 6.825 ;
        RECT 85.065 6.825 86.995 6.995 ;
        RECT 82.165 5.125 83.215 5.295 ;
        RECT 83.045 5.045 83.215 5.125 ;
        RECT 85.065 5.045 85.235 6.825 ;
        RECT 85.505 5.295 85.675 6.565 ;
        RECT 85.945 5.555 86.115 6.825 ;
        RECT 86.385 5.295 86.555 6.565 ;
        RECT 86.825 5.555 86.995 6.825 ;
        RECT 85.505 5.125 87.035 5.295 ;
        RECT 78.355 1.915 78.525 4.870 ;
        RECT 79.505 4.710 79.675 4.870 ;
        RECT 79.465 4.540 79.675 4.710 ;
        RECT 79.465 1.915 79.635 4.540 ;
        RECT 82.055 1.915 82.225 4.870 ;
        RECT 83.535 1.915 83.705 4.870 ;
        RECT 85.015 1.915 85.185 4.870 ;
        RECT 86.125 4.540 86.315 4.870 ;
        RECT 86.125 1.915 86.295 4.540 ;
        RECT 73.060 0.845 73.230 1.580 ;
        RECT 74.980 1.495 76.120 1.665 ;
        RECT 73.545 0.625 73.715 1.395 ;
        RECT 72.575 0.455 73.715 0.625 ;
        RECT 72.575 0.375 72.745 0.455 ;
        RECT 73.545 0.375 73.715 0.455 ;
        RECT 74.980 0.365 75.150 1.495 ;
        RECT 75.950 0.615 76.120 1.495 ;
        RECT 76.435 1.570 77.045 1.740 ;
        RECT 78.310 1.665 78.480 1.745 ;
        RECT 79.280 1.665 79.450 1.745 ;
        RECT 76.435 0.835 76.605 1.570 ;
        RECT 78.310 1.495 79.450 1.665 ;
        RECT 76.920 0.615 77.090 1.385 ;
        RECT 75.950 0.445 77.090 0.615 ;
        RECT 75.950 0.365 76.120 0.445 ;
        RECT 76.920 0.365 77.090 0.445 ;
        RECT 78.310 0.365 78.480 1.495 ;
        RECT 79.280 0.615 79.450 1.495 ;
        RECT 79.765 1.170 79.935 1.345 ;
        RECT 79.760 1.015 79.935 1.170 ;
        RECT 79.760 0.835 79.930 1.015 ;
        RECT 80.250 0.615 80.420 1.745 ;
        RECT 79.280 0.445 80.420 0.615 ;
        RECT 79.280 0.365 79.450 0.445 ;
        RECT 80.250 0.365 80.420 0.445 ;
        RECT 81.640 1.665 81.810 1.745 ;
        RECT 82.610 1.665 82.780 1.745 ;
        RECT 81.640 1.495 82.780 1.665 ;
        RECT 81.640 0.365 81.810 1.495 ;
        RECT 82.610 0.615 82.780 1.495 ;
        RECT 83.095 0.835 83.265 1.345 ;
        RECT 83.580 0.615 83.750 1.745 ;
        RECT 82.610 0.445 83.750 0.615 ;
        RECT 82.610 0.365 82.780 0.445 ;
        RECT 83.580 0.365 83.750 0.445 ;
        RECT 84.970 1.665 85.140 1.745 ;
        RECT 85.940 1.665 86.110 1.745 ;
        RECT 86.865 1.730 87.035 5.125 ;
        RECT 88.345 1.920 88.515 4.865 ;
        RECT 88.720 4.665 88.890 7.020 ;
        RECT 88.720 4.495 89.255 4.665 ;
        RECT 89.085 2.165 89.255 4.495 ;
        RECT 88.715 1.995 89.255 2.165 ;
        RECT 84.970 1.495 86.110 1.665 ;
        RECT 84.970 0.365 85.140 1.495 ;
        RECT 85.940 0.615 86.110 1.495 ;
        RECT 86.425 1.560 87.035 1.730 ;
        RECT 86.425 0.835 86.595 1.560 ;
        RECT 86.910 0.615 87.080 1.390 ;
        RECT 88.715 0.840 88.885 1.995 ;
        RECT 85.940 0.445 87.080 0.615 ;
        RECT 85.940 0.365 86.110 0.445 ;
        RECT 86.910 0.365 87.080 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 3.245 12.295 3.415 ;
        RECT 13.975 3.245 14.145 3.415 ;
        RECT 16.935 3.985 17.105 4.155 ;
        RECT 18.785 3.615 18.955 3.785 ;
        RECT 21.005 2.875 21.175 3.045 ;
        RECT 21.745 3.985 21.915 4.155 ;
        RECT 23.595 3.985 23.765 4.155 ;
        RECT 24.335 3.985 24.505 4.155 ;
        RECT 25.075 2.875 25.245 3.045 ;
        RECT 26.925 3.985 27.095 4.155 ;
        RECT 29.145 3.245 29.315 3.415 ;
        RECT 29.885 3.615 30.055 3.785 ;
        RECT 31.735 3.615 31.905 3.785 ;
        RECT 34.695 3.245 34.865 3.415 ;
        RECT 36.545 3.245 36.715 3.415 ;
        RECT 37.285 3.985 37.455 4.155 ;
        RECT 38.025 3.245 38.195 3.415 ;
        RECT 39.875 3.245 40.045 3.415 ;
        RECT 42.835 3.985 43.005 4.155 ;
        RECT 44.685 3.615 44.855 3.785 ;
        RECT 46.905 3.245 47.075 3.415 ;
        RECT 47.645 3.615 47.815 3.785 ;
        RECT 49.495 3.615 49.665 3.785 ;
        RECT 50.235 3.985 50.405 4.155 ;
        RECT 50.975 3.245 51.145 3.415 ;
        RECT 52.825 3.985 52.995 4.155 ;
        RECT 55.045 3.245 55.215 3.415 ;
        RECT 55.785 3.615 55.955 3.785 ;
        RECT 57.635 3.615 57.805 3.785 ;
        RECT 60.595 3.245 60.765 3.415 ;
        RECT 62.445 3.245 62.615 3.415 ;
        RECT 63.185 3.985 63.355 4.155 ;
        RECT 79.725 5.125 79.895 5.295 ;
        RECT 63.925 3.245 64.095 3.415 ;
        RECT 65.775 3.245 65.945 3.415 ;
        RECT 68.735 3.985 68.905 4.155 ;
        RECT 70.585 3.615 70.755 3.785 ;
        RECT 72.805 3.615 72.975 3.785 ;
        RECT 73.545 3.985 73.715 4.155 ;
        RECT 75.395 3.985 75.565 4.155 ;
        RECT 76.135 3.985 76.305 4.155 ;
        RECT 81.725 5.125 81.895 5.295 ;
        RECT 83.045 5.125 83.215 5.295 ;
        RECT 85.065 5.125 85.235 5.295 ;
        RECT 76.875 3.615 77.045 3.785 ;
        RECT 78.355 4.355 78.525 4.525 ;
        RECT 78.355 3.245 78.525 3.415 ;
        RECT 79.465 3.985 79.635 4.155 ;
        RECT 79.465 3.615 79.635 3.785 ;
        RECT 82.055 4.355 82.225 4.525 ;
        RECT 83.535 2.875 83.705 3.045 ;
        RECT 83.535 1.995 83.705 2.165 ;
        RECT 85.015 1.995 85.185 2.165 ;
        RECT 86.125 3.985 86.295 4.155 ;
        RECT 86.865 3.985 87.035 4.155 ;
        RECT 79.765 1.095 79.935 1.265 ;
        RECT 83.095 1.095 83.265 1.265 ;
        RECT 88.345 3.985 88.515 4.155 ;
        RECT 86.425 1.095 86.595 1.265 ;
      LAYER met1 ;
        RECT 79.695 5.295 79.925 5.325 ;
        RECT 81.695 5.295 81.925 5.325 ;
        RECT 83.015 5.295 83.245 5.325 ;
        RECT 85.035 5.295 85.265 5.325 ;
        RECT 79.665 5.125 81.955 5.295 ;
        RECT 82.985 5.125 85.295 5.295 ;
        RECT 79.695 5.095 79.925 5.125 ;
        RECT 81.695 5.095 81.925 5.125 ;
        RECT 83.015 5.095 83.245 5.125 ;
        RECT 85.035 5.095 85.265 5.125 ;
        RECT 78.325 4.525 78.555 4.555 ;
        RECT 82.025 4.525 82.255 4.555 ;
        RECT 78.295 4.355 82.285 4.525 ;
        RECT 78.325 4.325 78.555 4.355 ;
        RECT 82.025 4.325 82.255 4.355 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 16.905 4.155 17.135 4.185 ;
        RECT 21.715 4.155 21.945 4.185 ;
        RECT 23.565 4.155 23.795 4.185 ;
        RECT 24.305 4.155 24.535 4.185 ;
        RECT 26.895 4.155 27.125 4.185 ;
        RECT 37.255 4.155 37.485 4.185 ;
        RECT 42.805 4.155 43.035 4.185 ;
        RECT 50.205 4.155 50.435 4.185 ;
        RECT 52.795 4.155 53.025 4.185 ;
        RECT 63.155 4.155 63.385 4.185 ;
        RECT 68.705 4.155 68.935 4.185 ;
        RECT 73.515 4.155 73.745 4.185 ;
        RECT 75.365 4.155 75.595 4.185 ;
        RECT 76.105 4.155 76.335 4.185 ;
        RECT 79.435 4.155 79.665 4.185 ;
        RECT 86.095 4.155 86.325 4.185 ;
        RECT 86.835 4.155 87.065 4.185 ;
        RECT 88.315 4.155 88.545 4.185 ;
        RECT 0.965 3.985 24.565 4.155 ;
        RECT 26.865 3.985 50.465 4.155 ;
        RECT 52.765 3.985 76.365 4.155 ;
        RECT 79.405 3.985 86.355 4.155 ;
        RECT 86.805 3.985 88.575 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 16.905 3.955 17.135 3.985 ;
        RECT 21.715 3.955 21.945 3.985 ;
        RECT 23.565 3.955 23.795 3.985 ;
        RECT 24.305 3.955 24.535 3.985 ;
        RECT 26.895 3.955 27.125 3.985 ;
        RECT 37.255 3.955 37.485 3.985 ;
        RECT 42.805 3.955 43.035 3.985 ;
        RECT 50.205 3.955 50.435 3.985 ;
        RECT 52.795 3.955 53.025 3.985 ;
        RECT 63.155 3.955 63.385 3.985 ;
        RECT 68.705 3.955 68.935 3.985 ;
        RECT 73.515 3.955 73.745 3.985 ;
        RECT 75.365 3.955 75.595 3.985 ;
        RECT 76.105 3.955 76.335 3.985 ;
        RECT 79.435 3.955 79.665 3.985 ;
        RECT 86.095 3.955 86.325 3.985 ;
        RECT 86.835 3.955 87.065 3.985 ;
        RECT 88.315 3.955 88.545 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 18.755 3.785 18.985 3.815 ;
        RECT 29.855 3.785 30.085 3.815 ;
        RECT 31.705 3.785 31.935 3.815 ;
        RECT 44.655 3.785 44.885 3.815 ;
        RECT 47.615 3.785 47.845 3.815 ;
        RECT 49.465 3.785 49.695 3.815 ;
        RECT 55.755 3.785 55.985 3.815 ;
        RECT 57.605 3.785 57.835 3.815 ;
        RECT 70.555 3.785 70.785 3.815 ;
        RECT 72.775 3.785 73.005 3.815 ;
        RECT 76.845 3.785 77.075 3.815 ;
        RECT 79.435 3.785 79.665 3.815 ;
        RECT 3.925 3.615 19.015 3.785 ;
        RECT 29.825 3.615 44.915 3.785 ;
        RECT 47.585 3.615 49.725 3.785 ;
        RECT 55.725 3.615 70.815 3.785 ;
        RECT 72.745 3.615 79.695 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 18.755 3.585 18.985 3.615 ;
        RECT 29.855 3.585 30.085 3.615 ;
        RECT 31.705 3.585 31.935 3.615 ;
        RECT 44.655 3.585 44.885 3.615 ;
        RECT 47.615 3.585 47.845 3.615 ;
        RECT 49.465 3.585 49.695 3.615 ;
        RECT 55.755 3.585 55.985 3.615 ;
        RECT 57.605 3.585 57.835 3.615 ;
        RECT 70.555 3.585 70.785 3.615 ;
        RECT 72.775 3.585 73.005 3.615 ;
        RECT 76.845 3.585 77.075 3.615 ;
        RECT 79.435 3.585 79.665 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 8.765 3.415 8.995 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.095 3.415 12.325 3.445 ;
        RECT 13.945 3.415 14.175 3.445 ;
        RECT 29.115 3.415 29.345 3.445 ;
        RECT 34.665 3.415 34.895 3.445 ;
        RECT 36.515 3.415 36.745 3.445 ;
        RECT 37.995 3.415 38.225 3.445 ;
        RECT 39.845 3.415 40.075 3.445 ;
        RECT 46.875 3.415 47.105 3.445 ;
        RECT 50.945 3.415 51.175 3.445 ;
        RECT 55.015 3.415 55.245 3.445 ;
        RECT 60.565 3.415 60.795 3.445 ;
        RECT 62.415 3.415 62.645 3.445 ;
        RECT 63.895 3.415 64.125 3.445 ;
        RECT 65.745 3.415 65.975 3.445 ;
        RECT 78.325 3.415 78.555 3.445 ;
        RECT 3.185 3.245 10.875 3.415 ;
        RECT 12.065 3.245 14.205 3.415 ;
        RECT 29.085 3.245 36.775 3.415 ;
        RECT 37.965 3.245 40.105 3.415 ;
        RECT 46.845 3.245 78.585 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 8.765 3.215 8.995 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.095 3.215 12.325 3.245 ;
        RECT 13.945 3.215 14.175 3.245 ;
        RECT 29.115 3.215 29.345 3.245 ;
        RECT 34.665 3.215 34.895 3.245 ;
        RECT 36.515 3.215 36.745 3.245 ;
        RECT 37.995 3.215 38.225 3.245 ;
        RECT 39.845 3.215 40.075 3.245 ;
        RECT 46.875 3.215 47.105 3.245 ;
        RECT 50.945 3.215 51.175 3.245 ;
        RECT 55.015 3.215 55.245 3.245 ;
        RECT 60.565 3.215 60.795 3.245 ;
        RECT 62.415 3.215 62.645 3.245 ;
        RECT 63.895 3.215 64.125 3.245 ;
        RECT 65.745 3.215 65.975 3.245 ;
        RECT 78.325 3.215 78.555 3.245 ;
        RECT 20.975 3.045 21.205 3.075 ;
        RECT 25.045 3.045 25.275 3.075 ;
        RECT 83.505 3.045 83.735 3.075 ;
        RECT 20.945 2.875 83.765 3.045 ;
        RECT 20.975 2.845 21.205 2.875 ;
        RECT 25.045 2.845 25.275 2.875 ;
        RECT 83.505 2.845 83.735 2.875 ;
        RECT 83.505 2.165 83.735 2.195 ;
        RECT 84.985 2.165 85.215 2.195 ;
        RECT 83.475 1.995 85.245 2.165 ;
        RECT 83.505 1.965 83.735 1.995 ;
        RECT 84.985 1.965 85.215 1.995 ;
        RECT 79.735 1.265 79.965 1.295 ;
        RECT 83.065 1.265 83.295 1.295 ;
        RECT 86.395 1.265 86.625 1.295 ;
        RECT 79.705 1.095 86.655 1.265 ;
        RECT 79.735 1.065 79.965 1.095 ;
        RECT 83.065 1.065 83.295 1.095 ;
        RECT 86.395 1.065 86.625 1.095 ;
  END
END TMRDFFRNQX1






MACRO TMRDFFSNQNX1
  CLASS CORE ;
  FOREIGN TMRDFFSNQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 83.250 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN D
    ANTENNAGATEAREA 3.099750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 25.445 1.915 25.615 4.865 ;
        RECT 49.865 1.915 50.035 4.865 ;
      LAYER mcon ;
        RECT 1.025 2.875 1.195 3.045 ;
        RECT 25.445 2.875 25.615 3.045 ;
        RECT 49.865 2.875 50.035 3.045 ;
      LAYER met1 ;
        RECT 0.995 3.045 1.225 3.075 ;
        RECT 25.415 3.045 25.645 3.075 ;
        RECT 49.835 3.045 50.065 3.075 ;
        RECT 0.965 2.875 50.095 3.045 ;
        RECT 0.995 2.845 1.225 2.875 ;
        RECT 25.415 2.845 25.645 2.875 ;
        RECT 49.835 2.845 50.065 2.875 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.126300 ;
    PORT
      LAYER li1 ;
        RECT 5.465 1.915 5.635 4.865 ;
        RECT 14.745 4.710 14.915 4.865 ;
        RECT 14.715 4.535 14.915 4.710 ;
        RECT 14.715 1.915 14.885 4.535 ;
        RECT 29.885 1.915 30.055 4.865 ;
        RECT 39.165 4.710 39.335 4.865 ;
        RECT 39.135 4.535 39.335 4.710 ;
        RECT 39.135 1.915 39.305 4.535 ;
        RECT 54.305 1.915 54.475 4.865 ;
        RECT 63.585 4.710 63.755 4.865 ;
        RECT 63.555 4.535 63.755 4.710 ;
        RECT 63.555 1.915 63.725 4.535 ;
      LAYER mcon ;
        RECT 5.465 4.355 5.635 4.525 ;
        RECT 14.715 4.355 14.885 4.525 ;
        RECT 29.885 4.355 30.055 4.525 ;
        RECT 39.135 4.355 39.305 4.525 ;
        RECT 54.305 4.355 54.475 4.525 ;
        RECT 63.555 4.355 63.725 4.525 ;
      LAYER met1 ;
        RECT 5.435 4.525 5.665 4.555 ;
        RECT 14.685 4.525 14.915 4.555 ;
        RECT 29.855 4.525 30.085 4.555 ;
        RECT 39.105 4.525 39.335 4.555 ;
        RECT 54.275 4.525 54.505 4.555 ;
        RECT 63.525 4.525 63.755 4.555 ;
        RECT 5.405 4.355 63.785 4.525 ;
        RECT 5.435 4.325 5.665 4.355 ;
        RECT 14.685 4.325 14.915 4.355 ;
        RECT 29.855 4.325 30.085 4.355 ;
        RECT 39.105 4.325 39.335 4.355 ;
        RECT 54.275 4.325 54.505 4.355 ;
        RECT 63.525 4.325 63.755 4.355 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 10.275 1.915 10.445 4.865 ;
        RECT 21.745 1.915 21.915 4.865 ;
        RECT 34.695 1.915 34.865 4.865 ;
        RECT 46.165 1.915 46.335 4.865 ;
        RECT 59.115 1.915 59.285 4.865 ;
        RECT 70.585 1.915 70.755 4.865 ;
      LAYER mcon ;
        RECT 10.275 2.135 10.445 2.305 ;
        RECT 21.745 2.135 21.915 2.305 ;
        RECT 34.695 2.135 34.865 2.305 ;
        RECT 46.165 2.135 46.335 2.305 ;
        RECT 59.115 2.135 59.285 2.305 ;
        RECT 70.585 2.135 70.755 2.305 ;
      LAYER met1 ;
        RECT 10.245 2.305 10.475 2.335 ;
        RECT 21.715 2.305 21.945 2.335 ;
        RECT 34.665 2.305 34.895 2.335 ;
        RECT 46.135 2.305 46.365 2.335 ;
        RECT 59.085 2.305 59.315 2.335 ;
        RECT 70.555 2.305 70.785 2.335 ;
        RECT 10.215 2.135 70.815 2.305 ;
        RECT 10.245 2.105 10.475 2.135 ;
        RECT 21.715 2.105 21.945 2.135 ;
        RECT 34.665 2.105 34.895 2.135 ;
        RECT 46.135 2.105 46.365 2.135 ;
        RECT 59.085 2.105 59.315 2.135 ;
        RECT 70.555 2.105 70.785 2.135 ;
    END
  END SN
  PIN VPB
    ANTENNADIFFAREA 106.024750 ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 83.685 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 83.420 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.335 5.215 4.505 7.230 ;
        RECT 5.215 5.555 5.385 7.230 ;
        RECT 6.095 5.555 6.265 7.230 ;
        RECT 6.975 5.555 7.145 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 9.145 5.215 9.315 7.230 ;
        RECT 10.025 5.555 10.195 7.230 ;
        RECT 10.905 5.555 11.075 7.230 ;
        RECT 11.785 5.555 11.955 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.655 5.135 13.825 7.230 ;
        RECT 14.535 5.555 14.705 7.230 ;
        RECT 15.415 5.555 15.585 7.230 ;
        RECT 16.110 4.110 16.450 7.230 ;
        RECT 16.985 5.135 17.155 7.230 ;
        RECT 17.865 5.555 18.035 7.230 ;
        RECT 18.745 5.555 18.915 7.230 ;
        RECT 19.440 4.110 19.780 7.230 ;
        RECT 20.615 5.215 20.785 7.230 ;
        RECT 21.495 5.555 21.665 7.230 ;
        RECT 22.375 5.555 22.545 7.230 ;
        RECT 23.255 5.555 23.425 7.230 ;
        RECT 24.250 4.110 24.590 7.230 ;
        RECT 25.125 5.135 25.295 7.230 ;
        RECT 26.005 5.555 26.175 7.230 ;
        RECT 26.885 5.555 27.055 7.230 ;
        RECT 27.580 4.110 27.920 7.230 ;
        RECT 28.755 5.215 28.925 7.230 ;
        RECT 29.635 5.555 29.805 7.230 ;
        RECT 30.515 5.555 30.685 7.230 ;
        RECT 31.395 5.555 31.565 7.230 ;
        RECT 32.390 4.110 32.730 7.230 ;
        RECT 33.565 5.215 33.735 7.230 ;
        RECT 34.445 5.555 34.615 7.230 ;
        RECT 35.325 5.555 35.495 7.230 ;
        RECT 36.205 5.555 36.375 7.230 ;
        RECT 37.200 4.110 37.540 7.230 ;
        RECT 38.075 5.135 38.245 7.230 ;
        RECT 38.955 5.555 39.125 7.230 ;
        RECT 39.835 5.555 40.005 7.230 ;
        RECT 40.530 4.110 40.870 7.230 ;
        RECT 41.405 5.135 41.575 7.230 ;
        RECT 42.285 5.555 42.455 7.230 ;
        RECT 43.165 5.555 43.335 7.230 ;
        RECT 43.860 4.110 44.200 7.230 ;
        RECT 45.035 5.215 45.205 7.230 ;
        RECT 45.915 5.555 46.085 7.230 ;
        RECT 46.795 5.555 46.965 7.230 ;
        RECT 47.675 5.555 47.845 7.230 ;
        RECT 48.670 4.110 49.010 7.230 ;
        RECT 49.545 5.135 49.715 7.230 ;
        RECT 50.425 5.555 50.595 7.230 ;
        RECT 51.305 5.555 51.475 7.230 ;
        RECT 52.000 4.110 52.340 7.230 ;
        RECT 53.175 5.215 53.345 7.230 ;
        RECT 54.055 5.555 54.225 7.230 ;
        RECT 54.935 5.555 55.105 7.230 ;
        RECT 55.815 5.555 55.985 7.230 ;
        RECT 56.810 4.110 57.150 7.230 ;
        RECT 57.985 5.215 58.155 7.230 ;
        RECT 58.865 5.555 59.035 7.230 ;
        RECT 59.745 5.555 59.915 7.230 ;
        RECT 60.625 5.555 60.795 7.230 ;
        RECT 61.620 4.110 61.960 7.230 ;
        RECT 62.495 5.135 62.665 7.230 ;
        RECT 63.375 5.555 63.545 7.230 ;
        RECT 64.255 5.555 64.425 7.230 ;
        RECT 64.950 4.110 65.290 7.230 ;
        RECT 65.825 5.135 65.995 7.230 ;
        RECT 66.705 5.555 66.875 7.230 ;
        RECT 67.585 5.555 67.755 7.230 ;
        RECT 68.280 4.110 68.620 7.230 ;
        RECT 69.455 5.215 69.625 7.230 ;
        RECT 70.335 5.555 70.505 7.230 ;
        RECT 71.215 5.555 71.385 7.230 ;
        RECT 72.095 5.555 72.265 7.230 ;
        RECT 73.090 4.110 73.430 7.230 ;
        RECT 73.965 5.125 74.135 7.230 ;
        RECT 74.845 5.555 75.015 7.230 ;
        RECT 75.725 5.125 75.895 7.230 ;
        RECT 76.420 4.110 76.760 7.230 ;
        RECT 79.750 4.110 80.090 7.230 ;
        RECT 83.080 4.110 83.420 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.515 7.315 29.685 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.625 7.315 30.795 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.845 7.315 33.015 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.435 7.315 35.605 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.175 7.315 36.345 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
        RECT 38.765 7.315 38.935 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.505 7.315 39.675 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 42.835 7.315 43.005 7.485 ;
        RECT 43.205 7.315 43.375 7.485 ;
        RECT 43.575 7.315 43.745 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 47.645 7.315 47.815 7.485 ;
        RECT 48.015 7.315 48.185 7.485 ;
        RECT 48.385 7.315 48.555 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 50.975 7.315 51.145 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 51.715 7.315 51.885 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 52.825 7.315 52.995 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.305 7.315 54.475 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.525 7.315 56.695 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 57.635 7.315 57.805 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 60.965 7.315 61.135 7.485 ;
        RECT 61.335 7.315 61.505 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.445 7.315 62.615 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.295 7.315 64.465 7.485 ;
        RECT 64.665 7.315 64.835 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.255 7.315 67.425 7.485 ;
        RECT 67.625 7.315 67.795 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.475 7.315 69.645 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 70.955 7.315 71.125 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.065 7.315 72.235 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
        RECT 74.285 7.315 74.455 7.485 ;
        RECT 74.655 7.315 74.825 7.485 ;
        RECT 75.025 7.315 75.195 7.485 ;
        RECT 75.395 7.315 75.565 7.485 ;
        RECT 75.765 7.315 75.935 7.485 ;
        RECT 76.135 7.315 76.305 7.485 ;
        RECT 76.875 7.315 77.045 7.485 ;
        RECT 77.245 7.315 77.415 7.485 ;
        RECT 77.615 7.315 77.785 7.485 ;
        RECT 77.985 7.315 78.155 7.485 ;
        RECT 78.355 7.315 78.525 7.485 ;
        RECT 78.725 7.315 78.895 7.485 ;
        RECT 79.095 7.315 79.265 7.485 ;
        RECT 79.465 7.315 79.635 7.485 ;
        RECT 80.205 7.315 80.375 7.485 ;
        RECT 80.575 7.315 80.745 7.485 ;
        RECT 80.945 7.315 81.115 7.485 ;
        RECT 81.315 7.315 81.485 7.485 ;
        RECT 81.685 7.315 81.855 7.485 ;
        RECT 82.055 7.315 82.225 7.485 ;
        RECT 82.425 7.315 82.595 7.485 ;
        RECT 82.795 7.315 82.965 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 83.420 7.570 ;
    END
  END VPB
  PIN VNB
    ANTENNADIFFAREA 68.649246 ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 83.420 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 4.320 0.170 4.490 1.130 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.130 0.170 9.300 1.130 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 14.045 0.170 14.215 1.120 ;
        RECT 16.110 0.170 16.450 2.720 ;
        RECT 17.375 0.170 17.545 1.120 ;
        RECT 19.440 0.170 19.780 2.720 ;
        RECT 20.600 0.170 20.770 1.130 ;
        RECT 24.250 0.170 24.590 2.720 ;
        RECT 25.515 0.170 25.685 1.120 ;
        RECT 27.580 0.170 27.920 2.720 ;
        RECT 28.740 0.170 28.910 1.130 ;
        RECT 32.390 0.170 32.730 2.720 ;
        RECT 33.550 0.170 33.720 1.130 ;
        RECT 37.200 0.170 37.540 2.720 ;
        RECT 38.465 0.170 38.635 1.120 ;
        RECT 40.530 0.170 40.870 2.720 ;
        RECT 41.795 0.170 41.965 1.120 ;
        RECT 43.860 0.170 44.200 2.720 ;
        RECT 45.020 0.170 45.190 1.130 ;
        RECT 48.670 0.170 49.010 2.720 ;
        RECT 49.935 0.170 50.105 1.120 ;
        RECT 52.000 0.170 52.340 2.720 ;
        RECT 53.160 0.170 53.330 1.130 ;
        RECT 56.810 0.170 57.150 2.720 ;
        RECT 57.970 0.170 58.140 1.130 ;
        RECT 61.620 0.170 61.960 2.720 ;
        RECT 62.885 0.170 63.055 1.120 ;
        RECT 64.950 0.170 65.290 2.720 ;
        RECT 66.215 0.170 66.385 1.120 ;
        RECT 68.280 0.170 68.620 2.720 ;
        RECT 69.440 0.170 69.610 1.130 ;
        RECT 73.090 0.170 73.430 2.720 ;
        RECT 74.355 0.170 74.525 1.120 ;
        RECT 76.420 0.170 76.760 2.720 ;
        RECT 77.685 0.170 77.855 1.120 ;
        RECT 79.750 0.170 80.090 2.720 ;
        RECT 81.015 0.170 81.185 1.120 ;
        RECT 83.080 0.170 83.420 2.720 ;
        RECT -0.170 -0.170 83.420 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.515 -0.085 29.685 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.625 -0.085 30.795 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.845 -0.085 33.015 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.435 -0.085 35.605 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.175 -0.085 36.345 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
        RECT 38.765 -0.085 38.935 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.505 -0.085 39.675 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 42.835 -0.085 43.005 0.085 ;
        RECT 43.205 -0.085 43.375 0.085 ;
        RECT 43.575 -0.085 43.745 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 47.645 -0.085 47.815 0.085 ;
        RECT 48.015 -0.085 48.185 0.085 ;
        RECT 48.385 -0.085 48.555 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 50.975 -0.085 51.145 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 51.715 -0.085 51.885 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 52.825 -0.085 52.995 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.305 -0.085 54.475 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.525 -0.085 56.695 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 57.635 -0.085 57.805 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 60.965 -0.085 61.135 0.085 ;
        RECT 61.335 -0.085 61.505 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.445 -0.085 62.615 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.295 -0.085 64.465 0.085 ;
        RECT 64.665 -0.085 64.835 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.255 -0.085 67.425 0.085 ;
        RECT 67.625 -0.085 67.795 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.475 -0.085 69.645 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 70.955 -0.085 71.125 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.065 -0.085 72.235 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
        RECT 74.285 -0.085 74.455 0.085 ;
        RECT 74.655 -0.085 74.825 0.085 ;
        RECT 75.025 -0.085 75.195 0.085 ;
        RECT 75.395 -0.085 75.565 0.085 ;
        RECT 75.765 -0.085 75.935 0.085 ;
        RECT 76.135 -0.085 76.305 0.085 ;
        RECT 76.875 -0.085 77.045 0.085 ;
        RECT 77.245 -0.085 77.415 0.085 ;
        RECT 77.615 -0.085 77.785 0.085 ;
        RECT 77.985 -0.085 78.155 0.085 ;
        RECT 78.355 -0.085 78.525 0.085 ;
        RECT 78.725 -0.085 78.895 0.085 ;
        RECT 79.095 -0.085 79.265 0.085 ;
        RECT 79.465 -0.085 79.635 0.085 ;
        RECT 80.205 -0.085 80.375 0.085 ;
        RECT 80.575 -0.085 80.745 0.085 ;
        RECT 80.945 -0.085 81.115 0.085 ;
        RECT 81.315 -0.085 81.485 0.085 ;
        RECT 81.685 -0.085 81.855 0.085 ;
        RECT 82.055 -0.085 82.225 0.085 ;
        RECT 82.425 -0.085 82.595 0.085 ;
        RECT 82.795 -0.085 82.965 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 83.420 0.170 ;
    END
  END VNB
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.775 5.240 4.945 7.020 ;
        RECT 5.655 5.240 5.825 7.020 ;
        RECT 6.535 5.240 6.705 7.020 ;
        RECT 9.585 5.240 9.755 7.020 ;
        RECT 10.465 5.240 10.635 7.020 ;
        RECT 11.345 5.240 11.515 7.020 ;
        RECT 14.095 5.285 14.265 7.020 ;
        RECT 14.975 5.285 15.145 7.020 ;
        RECT 17.425 5.285 17.595 7.020 ;
        RECT 18.305 5.285 18.475 7.020 ;
        RECT 4.775 5.070 7.485 5.240 ;
        RECT 9.585 5.070 12.295 5.240 ;
        RECT 14.095 5.115 15.625 5.285 ;
        RECT 17.425 5.115 18.955 5.285 ;
        RECT 4.355 1.915 4.525 4.865 ;
        RECT 6.575 1.915 6.745 4.865 ;
        RECT 7.315 4.235 7.485 5.070 ;
        RECT 7.310 3.905 7.485 4.235 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 3.835 1.675 4.005 1.755 ;
        RECT 4.805 1.675 4.975 1.755 ;
        RECT 5.775 1.675 5.945 1.755 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 3.835 1.505 5.945 1.675 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 3.835 0.375 4.005 1.505 ;
        RECT 4.805 0.625 4.975 1.505 ;
        RECT 5.775 1.425 5.945 1.505 ;
        RECT 5.295 1.080 5.465 1.160 ;
        RECT 6.345 1.080 6.515 1.755 ;
        RECT 7.315 1.750 7.485 3.905 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 11.385 1.915 11.555 4.865 ;
        RECT 5.295 0.910 6.515 1.080 ;
        RECT 5.295 0.830 5.465 0.910 ;
        RECT 5.775 0.625 5.945 0.705 ;
        RECT 4.805 0.455 5.945 0.625 ;
        RECT 4.805 0.375 4.975 0.455 ;
        RECT 5.775 0.375 5.945 0.455 ;
        RECT 6.345 0.625 6.515 0.910 ;
        RECT 6.830 1.580 7.485 1.750 ;
        RECT 8.645 1.675 8.815 1.755 ;
        RECT 9.615 1.675 9.785 1.755 ;
        RECT 10.585 1.675 10.755 1.755 ;
        RECT 6.830 0.845 7.000 1.580 ;
        RECT 8.645 1.505 10.755 1.675 ;
        RECT 7.315 0.625 7.485 1.395 ;
        RECT 6.345 0.455 7.485 0.625 ;
        RECT 6.345 0.375 6.515 0.455 ;
        RECT 7.315 0.375 7.485 0.455 ;
        RECT 8.645 0.375 8.815 1.505 ;
        RECT 9.615 0.625 9.785 1.505 ;
        RECT 10.585 1.425 10.755 1.505 ;
        RECT 10.105 1.080 10.275 1.160 ;
        RECT 11.155 1.080 11.325 1.755 ;
        RECT 12.125 1.750 12.295 5.070 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 10.105 0.910 11.325 1.080 ;
        RECT 10.105 0.830 10.275 0.910 ;
        RECT 10.585 0.625 10.755 0.705 ;
        RECT 9.615 0.455 10.755 0.625 ;
        RECT 9.615 0.375 9.785 0.455 ;
        RECT 10.585 0.375 10.755 0.455 ;
        RECT 11.155 0.625 11.325 0.910 ;
        RECT 11.640 1.580 12.295 1.750 ;
        RECT 13.560 1.665 13.730 1.745 ;
        RECT 14.530 1.665 14.700 1.745 ;
        RECT 15.455 1.740 15.625 5.115 ;
        RECT 17.305 1.915 17.475 4.865 ;
        RECT 18.075 4.710 18.245 4.865 ;
        RECT 18.045 4.535 18.245 4.710 ;
        RECT 18.045 1.915 18.215 4.535 ;
        RECT 11.640 0.845 11.810 1.580 ;
        RECT 13.560 1.495 14.700 1.665 ;
        RECT 12.125 0.625 12.295 1.395 ;
        RECT 11.155 0.455 12.295 0.625 ;
        RECT 11.155 0.375 11.325 0.455 ;
        RECT 12.125 0.375 12.295 0.455 ;
        RECT 13.560 0.365 13.730 1.495 ;
        RECT 14.530 0.615 14.700 1.495 ;
        RECT 15.015 1.570 15.625 1.740 ;
        RECT 16.890 1.665 17.060 1.745 ;
        RECT 17.860 1.665 18.030 1.745 ;
        RECT 18.785 1.740 18.955 5.115 ;
        RECT 21.055 5.240 21.225 7.020 ;
        RECT 21.935 5.240 22.105 7.020 ;
        RECT 22.815 5.240 22.985 7.020 ;
        RECT 25.565 5.285 25.735 7.020 ;
        RECT 26.445 5.285 26.615 7.020 ;
        RECT 21.055 5.070 23.765 5.240 ;
        RECT 25.565 5.115 27.095 5.285 ;
        RECT 20.635 1.915 20.805 4.865 ;
        RECT 22.855 1.915 23.025 4.865 ;
        RECT 15.015 0.835 15.185 1.570 ;
        RECT 16.890 1.495 18.030 1.665 ;
        RECT 15.500 0.615 15.670 1.385 ;
        RECT 14.530 0.445 15.670 0.615 ;
        RECT 14.530 0.365 14.700 0.445 ;
        RECT 15.500 0.365 15.670 0.445 ;
        RECT 16.890 0.365 17.060 1.495 ;
        RECT 17.860 0.615 18.030 1.495 ;
        RECT 18.345 1.570 18.955 1.740 ;
        RECT 20.115 1.675 20.285 1.755 ;
        RECT 21.085 1.675 21.255 1.755 ;
        RECT 22.055 1.675 22.225 1.755 ;
        RECT 18.345 0.835 18.515 1.570 ;
        RECT 20.115 1.505 22.225 1.675 ;
        RECT 18.830 0.615 19.000 1.385 ;
        RECT 17.860 0.445 19.000 0.615 ;
        RECT 17.860 0.365 18.030 0.445 ;
        RECT 18.830 0.365 19.000 0.445 ;
        RECT 20.115 0.375 20.285 1.505 ;
        RECT 21.085 0.625 21.255 1.505 ;
        RECT 22.055 1.425 22.225 1.505 ;
        RECT 21.575 1.080 21.745 1.160 ;
        RECT 22.625 1.080 22.795 1.755 ;
        RECT 23.595 1.750 23.765 5.070 ;
        RECT 26.215 4.710 26.385 4.865 ;
        RECT 26.185 4.535 26.385 4.710 ;
        RECT 26.185 1.915 26.355 4.535 ;
        RECT 21.575 0.910 22.795 1.080 ;
        RECT 21.575 0.830 21.745 0.910 ;
        RECT 22.055 0.625 22.225 0.705 ;
        RECT 21.085 0.455 22.225 0.625 ;
        RECT 21.085 0.375 21.255 0.455 ;
        RECT 22.055 0.375 22.225 0.455 ;
        RECT 22.625 0.625 22.795 0.910 ;
        RECT 23.110 1.580 23.765 1.750 ;
        RECT 25.030 1.665 25.200 1.745 ;
        RECT 26.000 1.665 26.170 1.745 ;
        RECT 26.925 1.740 27.095 5.115 ;
        RECT 29.195 5.240 29.365 7.020 ;
        RECT 30.075 5.240 30.245 7.020 ;
        RECT 30.955 5.240 31.125 7.020 ;
        RECT 34.005 5.240 34.175 7.020 ;
        RECT 34.885 5.240 35.055 7.020 ;
        RECT 35.765 5.240 35.935 7.020 ;
        RECT 38.515 5.285 38.685 7.020 ;
        RECT 39.395 5.285 39.565 7.020 ;
        RECT 41.845 5.285 42.015 7.020 ;
        RECT 42.725 5.285 42.895 7.020 ;
        RECT 29.195 5.070 31.905 5.240 ;
        RECT 34.005 5.070 36.715 5.240 ;
        RECT 38.515 5.115 40.045 5.285 ;
        RECT 41.845 5.115 43.375 5.285 ;
        RECT 28.775 1.915 28.945 4.865 ;
        RECT 30.995 1.915 31.165 4.865 ;
        RECT 31.735 4.235 31.905 5.070 ;
        RECT 31.730 3.905 31.905 4.235 ;
        RECT 23.110 0.845 23.280 1.580 ;
        RECT 25.030 1.495 26.170 1.665 ;
        RECT 23.595 0.625 23.765 1.395 ;
        RECT 22.625 0.455 23.765 0.625 ;
        RECT 22.625 0.375 22.795 0.455 ;
        RECT 23.595 0.375 23.765 0.455 ;
        RECT 25.030 0.365 25.200 1.495 ;
        RECT 26.000 0.615 26.170 1.495 ;
        RECT 26.485 1.570 27.095 1.740 ;
        RECT 28.255 1.675 28.425 1.755 ;
        RECT 29.225 1.675 29.395 1.755 ;
        RECT 30.195 1.675 30.365 1.755 ;
        RECT 26.485 0.835 26.655 1.570 ;
        RECT 28.255 1.505 30.365 1.675 ;
        RECT 26.970 0.615 27.140 1.385 ;
        RECT 26.000 0.445 27.140 0.615 ;
        RECT 26.000 0.365 26.170 0.445 ;
        RECT 26.970 0.365 27.140 0.445 ;
        RECT 28.255 0.375 28.425 1.505 ;
        RECT 29.225 0.625 29.395 1.505 ;
        RECT 30.195 1.425 30.365 1.505 ;
        RECT 29.715 1.080 29.885 1.160 ;
        RECT 30.765 1.080 30.935 1.755 ;
        RECT 31.735 1.750 31.905 3.905 ;
        RECT 33.585 1.915 33.755 4.865 ;
        RECT 35.805 1.915 35.975 4.865 ;
        RECT 29.715 0.910 30.935 1.080 ;
        RECT 29.715 0.830 29.885 0.910 ;
        RECT 30.195 0.625 30.365 0.705 ;
        RECT 29.225 0.455 30.365 0.625 ;
        RECT 29.225 0.375 29.395 0.455 ;
        RECT 30.195 0.375 30.365 0.455 ;
        RECT 30.765 0.625 30.935 0.910 ;
        RECT 31.250 1.580 31.905 1.750 ;
        RECT 33.065 1.675 33.235 1.755 ;
        RECT 34.035 1.675 34.205 1.755 ;
        RECT 35.005 1.675 35.175 1.755 ;
        RECT 31.250 0.845 31.420 1.580 ;
        RECT 33.065 1.505 35.175 1.675 ;
        RECT 31.735 0.625 31.905 1.395 ;
        RECT 30.765 0.455 31.905 0.625 ;
        RECT 30.765 0.375 30.935 0.455 ;
        RECT 31.735 0.375 31.905 0.455 ;
        RECT 33.065 0.375 33.235 1.505 ;
        RECT 34.035 0.625 34.205 1.505 ;
        RECT 35.005 1.425 35.175 1.505 ;
        RECT 34.525 1.080 34.695 1.160 ;
        RECT 35.575 1.080 35.745 1.755 ;
        RECT 36.545 1.750 36.715 5.070 ;
        RECT 38.395 1.915 38.565 4.865 ;
        RECT 34.525 0.910 35.745 1.080 ;
        RECT 34.525 0.830 34.695 0.910 ;
        RECT 35.005 0.625 35.175 0.705 ;
        RECT 34.035 0.455 35.175 0.625 ;
        RECT 34.035 0.375 34.205 0.455 ;
        RECT 35.005 0.375 35.175 0.455 ;
        RECT 35.575 0.625 35.745 0.910 ;
        RECT 36.060 1.580 36.715 1.750 ;
        RECT 37.980 1.665 38.150 1.745 ;
        RECT 38.950 1.665 39.120 1.745 ;
        RECT 39.875 1.740 40.045 5.115 ;
        RECT 41.725 1.915 41.895 4.865 ;
        RECT 42.495 4.710 42.665 4.865 ;
        RECT 42.465 4.535 42.665 4.710 ;
        RECT 42.465 1.915 42.635 4.535 ;
        RECT 36.060 0.845 36.230 1.580 ;
        RECT 37.980 1.495 39.120 1.665 ;
        RECT 36.545 0.625 36.715 1.395 ;
        RECT 35.575 0.455 36.715 0.625 ;
        RECT 35.575 0.375 35.745 0.455 ;
        RECT 36.545 0.375 36.715 0.455 ;
        RECT 37.980 0.365 38.150 1.495 ;
        RECT 38.950 0.615 39.120 1.495 ;
        RECT 39.435 1.570 40.045 1.740 ;
        RECT 41.310 1.665 41.480 1.745 ;
        RECT 42.280 1.665 42.450 1.745 ;
        RECT 43.205 1.740 43.375 5.115 ;
        RECT 45.475 5.240 45.645 7.020 ;
        RECT 46.355 5.240 46.525 7.020 ;
        RECT 47.235 5.240 47.405 7.020 ;
        RECT 49.985 5.285 50.155 7.020 ;
        RECT 50.865 5.285 51.035 7.020 ;
        RECT 45.475 5.070 48.185 5.240 ;
        RECT 49.985 5.115 51.515 5.285 ;
        RECT 45.055 1.915 45.225 4.865 ;
        RECT 47.275 1.915 47.445 4.865 ;
        RECT 39.435 0.835 39.605 1.570 ;
        RECT 41.310 1.495 42.450 1.665 ;
        RECT 39.920 0.615 40.090 1.385 ;
        RECT 38.950 0.445 40.090 0.615 ;
        RECT 38.950 0.365 39.120 0.445 ;
        RECT 39.920 0.365 40.090 0.445 ;
        RECT 41.310 0.365 41.480 1.495 ;
        RECT 42.280 0.615 42.450 1.495 ;
        RECT 42.765 1.570 43.375 1.740 ;
        RECT 44.535 1.675 44.705 1.755 ;
        RECT 45.505 1.675 45.675 1.755 ;
        RECT 46.475 1.675 46.645 1.755 ;
        RECT 42.765 0.835 42.935 1.570 ;
        RECT 44.535 1.505 46.645 1.675 ;
        RECT 43.250 0.615 43.420 1.385 ;
        RECT 42.280 0.445 43.420 0.615 ;
        RECT 42.280 0.365 42.450 0.445 ;
        RECT 43.250 0.365 43.420 0.445 ;
        RECT 44.535 0.375 44.705 1.505 ;
        RECT 45.505 0.625 45.675 1.505 ;
        RECT 46.475 1.425 46.645 1.505 ;
        RECT 45.995 1.080 46.165 1.160 ;
        RECT 47.045 1.080 47.215 1.755 ;
        RECT 48.015 1.750 48.185 5.070 ;
        RECT 50.635 4.710 50.805 4.865 ;
        RECT 50.605 4.535 50.805 4.710 ;
        RECT 50.605 1.915 50.775 4.535 ;
        RECT 45.995 0.910 47.215 1.080 ;
        RECT 45.995 0.830 46.165 0.910 ;
        RECT 46.475 0.625 46.645 0.705 ;
        RECT 45.505 0.455 46.645 0.625 ;
        RECT 45.505 0.375 45.675 0.455 ;
        RECT 46.475 0.375 46.645 0.455 ;
        RECT 47.045 0.625 47.215 0.910 ;
        RECT 47.530 1.580 48.185 1.750 ;
        RECT 49.450 1.665 49.620 1.745 ;
        RECT 50.420 1.665 50.590 1.745 ;
        RECT 51.345 1.740 51.515 5.115 ;
        RECT 53.615 5.240 53.785 7.020 ;
        RECT 54.495 5.240 54.665 7.020 ;
        RECT 55.375 5.240 55.545 7.020 ;
        RECT 58.425 5.240 58.595 7.020 ;
        RECT 59.305 5.240 59.475 7.020 ;
        RECT 60.185 5.240 60.355 7.020 ;
        RECT 62.935 5.285 63.105 7.020 ;
        RECT 63.815 5.285 63.985 7.020 ;
        RECT 66.265 5.285 66.435 7.020 ;
        RECT 67.145 5.285 67.315 7.020 ;
        RECT 53.615 5.070 56.325 5.240 ;
        RECT 58.425 5.070 61.135 5.240 ;
        RECT 62.935 5.115 64.465 5.285 ;
        RECT 66.265 5.115 67.795 5.285 ;
        RECT 53.195 1.915 53.365 4.865 ;
        RECT 55.415 1.915 55.585 4.865 ;
        RECT 56.155 4.235 56.325 5.070 ;
        RECT 56.150 3.905 56.325 4.235 ;
        RECT 47.530 0.845 47.700 1.580 ;
        RECT 49.450 1.495 50.590 1.665 ;
        RECT 48.015 0.625 48.185 1.395 ;
        RECT 47.045 0.455 48.185 0.625 ;
        RECT 47.045 0.375 47.215 0.455 ;
        RECT 48.015 0.375 48.185 0.455 ;
        RECT 49.450 0.365 49.620 1.495 ;
        RECT 50.420 0.615 50.590 1.495 ;
        RECT 50.905 1.570 51.515 1.740 ;
        RECT 52.675 1.675 52.845 1.755 ;
        RECT 53.645 1.675 53.815 1.755 ;
        RECT 54.615 1.675 54.785 1.755 ;
        RECT 50.905 0.835 51.075 1.570 ;
        RECT 52.675 1.505 54.785 1.675 ;
        RECT 51.390 0.615 51.560 1.385 ;
        RECT 50.420 0.445 51.560 0.615 ;
        RECT 50.420 0.365 50.590 0.445 ;
        RECT 51.390 0.365 51.560 0.445 ;
        RECT 52.675 0.375 52.845 1.505 ;
        RECT 53.645 0.625 53.815 1.505 ;
        RECT 54.615 1.425 54.785 1.505 ;
        RECT 54.135 1.080 54.305 1.160 ;
        RECT 55.185 1.080 55.355 1.755 ;
        RECT 56.155 1.750 56.325 3.905 ;
        RECT 58.005 1.915 58.175 4.865 ;
        RECT 60.225 1.915 60.395 4.865 ;
        RECT 54.135 0.910 55.355 1.080 ;
        RECT 54.135 0.830 54.305 0.910 ;
        RECT 54.615 0.625 54.785 0.705 ;
        RECT 53.645 0.455 54.785 0.625 ;
        RECT 53.645 0.375 53.815 0.455 ;
        RECT 54.615 0.375 54.785 0.455 ;
        RECT 55.185 0.625 55.355 0.910 ;
        RECT 55.670 1.580 56.325 1.750 ;
        RECT 57.485 1.675 57.655 1.755 ;
        RECT 58.455 1.675 58.625 1.755 ;
        RECT 59.425 1.675 59.595 1.755 ;
        RECT 55.670 0.845 55.840 1.580 ;
        RECT 57.485 1.505 59.595 1.675 ;
        RECT 56.155 0.625 56.325 1.395 ;
        RECT 55.185 0.455 56.325 0.625 ;
        RECT 55.185 0.375 55.355 0.455 ;
        RECT 56.155 0.375 56.325 0.455 ;
        RECT 57.485 0.375 57.655 1.505 ;
        RECT 58.455 0.625 58.625 1.505 ;
        RECT 59.425 1.425 59.595 1.505 ;
        RECT 58.945 1.080 59.115 1.160 ;
        RECT 59.995 1.080 60.165 1.755 ;
        RECT 60.965 1.750 61.135 5.070 ;
        RECT 62.815 1.915 62.985 4.865 ;
        RECT 58.945 0.910 60.165 1.080 ;
        RECT 58.945 0.830 59.115 0.910 ;
        RECT 59.425 0.625 59.595 0.705 ;
        RECT 58.455 0.455 59.595 0.625 ;
        RECT 58.455 0.375 58.625 0.455 ;
        RECT 59.425 0.375 59.595 0.455 ;
        RECT 59.995 0.625 60.165 0.910 ;
        RECT 60.480 1.580 61.135 1.750 ;
        RECT 62.400 1.665 62.570 1.745 ;
        RECT 63.370 1.665 63.540 1.745 ;
        RECT 64.295 1.740 64.465 5.115 ;
        RECT 66.145 1.915 66.315 4.865 ;
        RECT 66.915 4.710 67.085 4.865 ;
        RECT 66.885 4.535 67.085 4.710 ;
        RECT 66.885 1.915 67.055 4.535 ;
        RECT 60.480 0.845 60.650 1.580 ;
        RECT 62.400 1.495 63.540 1.665 ;
        RECT 60.965 0.625 61.135 1.395 ;
        RECT 59.995 0.455 61.135 0.625 ;
        RECT 59.995 0.375 60.165 0.455 ;
        RECT 60.965 0.375 61.135 0.455 ;
        RECT 62.400 0.365 62.570 1.495 ;
        RECT 63.370 0.615 63.540 1.495 ;
        RECT 63.855 1.570 64.465 1.740 ;
        RECT 65.730 1.665 65.900 1.745 ;
        RECT 66.700 1.665 66.870 1.745 ;
        RECT 67.625 1.740 67.795 5.115 ;
        RECT 69.895 5.240 70.065 7.020 ;
        RECT 70.775 5.240 70.945 7.020 ;
        RECT 71.655 5.240 71.825 7.020 ;
        RECT 74.405 6.825 74.585 6.995 ;
        RECT 74.405 5.295 74.575 6.825 ;
        RECT 75.285 5.295 75.455 6.995 ;
        RECT 69.895 5.070 72.605 5.240 ;
        RECT 74.405 5.125 75.455 5.295 ;
        RECT 69.475 1.915 69.645 4.865 ;
        RECT 71.695 1.915 71.865 4.865 ;
        RECT 63.855 0.835 64.025 1.570 ;
        RECT 65.730 1.495 66.870 1.665 ;
        RECT 64.340 0.615 64.510 1.385 ;
        RECT 63.370 0.445 64.510 0.615 ;
        RECT 63.370 0.365 63.540 0.445 ;
        RECT 64.340 0.365 64.510 0.445 ;
        RECT 65.730 0.365 65.900 1.495 ;
        RECT 66.700 0.615 66.870 1.495 ;
        RECT 67.185 1.570 67.795 1.740 ;
        RECT 68.955 1.675 69.125 1.755 ;
        RECT 69.925 1.675 70.095 1.755 ;
        RECT 70.895 1.675 71.065 1.755 ;
        RECT 67.185 0.835 67.355 1.570 ;
        RECT 68.955 1.505 71.065 1.675 ;
        RECT 67.670 0.615 67.840 1.385 ;
        RECT 66.700 0.445 67.840 0.615 ;
        RECT 66.700 0.365 66.870 0.445 ;
        RECT 67.670 0.365 67.840 0.445 ;
        RECT 68.955 0.375 69.125 1.505 ;
        RECT 69.925 0.625 70.095 1.505 ;
        RECT 70.895 1.425 71.065 1.505 ;
        RECT 70.415 1.080 70.585 1.160 ;
        RECT 71.465 1.080 71.635 1.755 ;
        RECT 72.435 1.750 72.605 5.070 ;
        RECT 75.285 5.045 75.455 5.125 ;
        RECT 77.285 6.825 79.215 6.995 ;
        RECT 77.285 5.045 77.455 6.825 ;
        RECT 77.725 5.295 77.895 6.565 ;
        RECT 78.165 5.555 78.335 6.825 ;
        RECT 78.605 5.295 78.775 6.565 ;
        RECT 79.045 5.375 79.215 6.825 ;
        RECT 80.625 6.825 82.555 6.995 ;
        RECT 77.725 5.125 78.775 5.295 ;
        RECT 78.605 5.045 78.775 5.125 ;
        RECT 80.625 5.045 80.795 6.825 ;
        RECT 81.065 5.295 81.235 6.565 ;
        RECT 81.505 5.555 81.675 6.825 ;
        RECT 81.945 5.295 82.115 6.565 ;
        RECT 82.385 5.555 82.555 6.825 ;
        RECT 81.065 5.125 82.595 5.295 ;
        RECT 73.915 1.915 74.085 4.870 ;
        RECT 75.065 4.710 75.235 4.870 ;
        RECT 75.025 4.540 75.235 4.710 ;
        RECT 75.025 1.915 75.195 4.540 ;
        RECT 77.615 1.915 77.785 4.870 ;
        RECT 79.095 1.915 79.265 4.870 ;
        RECT 80.575 1.915 80.745 4.870 ;
        RECT 81.685 4.540 81.875 4.870 ;
        RECT 81.685 1.915 81.855 4.540 ;
        RECT 70.415 0.910 71.635 1.080 ;
        RECT 70.415 0.830 70.585 0.910 ;
        RECT 70.895 0.625 71.065 0.705 ;
        RECT 69.925 0.455 71.065 0.625 ;
        RECT 69.925 0.375 70.095 0.455 ;
        RECT 70.895 0.375 71.065 0.455 ;
        RECT 71.465 0.625 71.635 0.910 ;
        RECT 71.950 1.580 72.605 1.750 ;
        RECT 73.870 1.665 74.040 1.745 ;
        RECT 74.840 1.665 75.010 1.745 ;
        RECT 71.950 0.845 72.120 1.580 ;
        RECT 73.870 1.495 75.010 1.665 ;
        RECT 72.435 0.625 72.605 1.395 ;
        RECT 71.465 0.455 72.605 0.625 ;
        RECT 71.465 0.375 71.635 0.455 ;
        RECT 72.435 0.375 72.605 0.455 ;
        RECT 73.870 0.365 74.040 1.495 ;
        RECT 74.840 0.615 75.010 1.495 ;
        RECT 75.325 1.170 75.495 1.345 ;
        RECT 75.320 1.015 75.495 1.170 ;
        RECT 75.320 0.835 75.490 1.015 ;
        RECT 75.810 0.615 75.980 1.745 ;
        RECT 74.840 0.445 75.980 0.615 ;
        RECT 74.840 0.365 75.010 0.445 ;
        RECT 75.810 0.365 75.980 0.445 ;
        RECT 77.200 1.665 77.370 1.745 ;
        RECT 78.170 1.665 78.340 1.745 ;
        RECT 77.200 1.495 78.340 1.665 ;
        RECT 77.200 0.365 77.370 1.495 ;
        RECT 78.170 0.615 78.340 1.495 ;
        RECT 78.655 0.835 78.825 1.345 ;
        RECT 79.140 0.615 79.310 1.745 ;
        RECT 78.170 0.445 79.310 0.615 ;
        RECT 78.170 0.365 78.340 0.445 ;
        RECT 79.140 0.365 79.310 0.445 ;
        RECT 80.530 1.665 80.700 1.745 ;
        RECT 81.500 1.665 81.670 1.745 ;
        RECT 82.425 1.730 82.595 5.125 ;
        RECT 80.530 1.495 81.670 1.665 ;
        RECT 80.530 0.365 80.700 1.495 ;
        RECT 81.500 0.615 81.670 1.495 ;
        RECT 81.985 1.560 82.595 1.730 ;
        RECT 81.985 0.835 82.155 1.560 ;
        RECT 82.470 0.615 82.640 1.390 ;
        RECT 81.500 0.445 82.640 0.615 ;
        RECT 81.500 0.365 81.670 0.445 ;
        RECT 82.470 0.365 82.640 0.445 ;
      LAYER mcon ;
        RECT 1.765 3.985 1.935 4.155 ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.500 4.525 2.670 ;
        RECT 7.310 3.985 7.480 4.155 ;
        RECT 6.575 3.615 6.745 3.785 ;
        RECT 9.165 2.505 9.335 2.675 ;
        RECT 11.385 3.615 11.555 3.785 ;
        RECT 12.125 2.505 12.295 2.675 ;
        RECT 13.975 2.505 14.145 2.675 ;
        RECT 15.455 3.615 15.625 3.785 ;
        RECT 17.305 3.985 17.475 4.155 ;
        RECT 18.045 3.985 18.215 4.155 ;
        RECT 18.785 3.245 18.955 3.415 ;
        RECT 20.635 3.245 20.805 3.415 ;
        RECT 22.855 3.615 23.025 3.785 ;
        RECT 23.595 3.985 23.765 4.155 ;
        RECT 26.185 3.985 26.355 4.155 ;
        RECT 26.925 2.505 27.095 2.675 ;
        RECT 28.775 2.500 28.945 2.670 ;
        RECT 31.730 3.985 31.900 4.155 ;
        RECT 30.995 3.615 31.165 3.785 ;
        RECT 33.585 2.505 33.755 2.675 ;
        RECT 35.805 3.615 35.975 3.785 ;
        RECT 36.545 2.505 36.715 2.675 ;
        RECT 38.395 2.505 38.565 2.675 ;
        RECT 39.875 3.615 40.045 3.785 ;
        RECT 41.725 3.985 41.895 4.155 ;
        RECT 42.465 3.985 42.635 4.155 ;
        RECT 43.205 2.505 43.375 2.675 ;
        RECT 45.055 2.505 45.225 2.675 ;
        RECT 47.275 3.615 47.445 3.785 ;
        RECT 48.015 3.985 48.185 4.155 ;
        RECT 50.605 3.985 50.775 4.155 ;
        RECT 51.345 2.505 51.515 2.675 ;
        RECT 53.195 2.500 53.365 2.670 ;
        RECT 56.150 3.985 56.320 4.155 ;
        RECT 55.415 3.615 55.585 3.785 ;
        RECT 58.005 2.505 58.175 2.675 ;
        RECT 60.225 3.615 60.395 3.785 ;
        RECT 60.965 2.505 61.135 2.675 ;
        RECT 62.815 2.505 62.985 2.675 ;
        RECT 64.295 3.615 64.465 3.785 ;
        RECT 66.145 3.985 66.315 4.155 ;
        RECT 66.885 3.985 67.055 4.155 ;
        RECT 75.285 5.125 75.455 5.295 ;
        RECT 67.625 4.355 67.795 4.525 ;
        RECT 69.475 4.355 69.645 4.525 ;
        RECT 71.695 3.615 71.865 3.785 ;
        RECT 77.285 5.125 77.455 5.295 ;
        RECT 78.605 5.125 78.775 5.295 ;
        RECT 80.625 5.125 80.795 5.295 ;
        RECT 72.435 3.985 72.605 4.155 ;
        RECT 73.915 4.355 74.085 4.525 ;
        RECT 75.025 3.985 75.195 4.155 ;
        RECT 75.025 2.875 75.195 3.045 ;
        RECT 77.615 4.355 77.785 4.525 ;
        RECT 79.095 3.245 79.265 3.415 ;
        RECT 79.095 1.995 79.265 2.165 ;
        RECT 80.575 1.995 80.745 2.165 ;
        RECT 81.685 3.985 81.855 4.155 ;
        RECT 75.325 1.095 75.495 1.265 ;
        RECT 78.655 1.095 78.825 1.265 ;
        RECT 81.985 1.095 82.155 1.265 ;
      LAYER met1 ;
        RECT 75.255 5.295 75.485 5.325 ;
        RECT 77.255 5.295 77.485 5.325 ;
        RECT 78.575 5.295 78.805 5.325 ;
        RECT 80.595 5.295 80.825 5.325 ;
        RECT 75.225 5.125 77.515 5.295 ;
        RECT 78.545 5.125 80.855 5.295 ;
        RECT 75.255 5.095 75.485 5.125 ;
        RECT 77.255 5.095 77.485 5.125 ;
        RECT 78.575 5.095 78.805 5.125 ;
        RECT 80.595 5.095 80.825 5.125 ;
        RECT 67.595 4.525 67.825 4.555 ;
        RECT 69.445 4.525 69.675 4.555 ;
        RECT 73.885 4.525 74.115 4.555 ;
        RECT 77.585 4.525 77.815 4.555 ;
        RECT 67.565 4.355 77.845 4.525 ;
        RECT 67.595 4.325 67.825 4.355 ;
        RECT 69.445 4.325 69.675 4.355 ;
        RECT 73.885 4.325 74.115 4.355 ;
        RECT 77.585 4.325 77.815 4.355 ;
        RECT 1.735 4.155 1.965 4.185 ;
        RECT 7.280 4.155 7.510 4.185 ;
        RECT 17.275 4.155 17.505 4.185 ;
        RECT 18.015 4.155 18.245 4.185 ;
        RECT 23.565 4.155 23.795 4.185 ;
        RECT 26.155 4.155 26.385 4.185 ;
        RECT 31.700 4.155 31.930 4.185 ;
        RECT 41.695 4.155 41.925 4.185 ;
        RECT 42.435 4.155 42.665 4.185 ;
        RECT 47.985 4.155 48.215 4.185 ;
        RECT 50.575 4.155 50.805 4.185 ;
        RECT 56.120 4.155 56.350 4.185 ;
        RECT 66.115 4.155 66.345 4.185 ;
        RECT 66.855 4.155 67.085 4.185 ;
        RECT 72.405 4.155 72.635 4.185 ;
        RECT 74.995 4.155 75.225 4.185 ;
        RECT 81.655 4.155 81.885 4.185 ;
        RECT 1.705 3.985 17.535 4.155 ;
        RECT 17.985 3.985 23.945 4.155 ;
        RECT 26.125 3.985 41.955 4.155 ;
        RECT 42.405 3.985 48.245 4.155 ;
        RECT 50.545 3.985 66.375 4.155 ;
        RECT 66.825 3.985 72.665 4.155 ;
        RECT 74.965 3.985 81.915 4.155 ;
        RECT 1.735 3.955 1.965 3.985 ;
        RECT 7.280 3.955 7.510 3.985 ;
        RECT 17.275 3.955 17.505 3.985 ;
        RECT 18.015 3.955 18.245 3.985 ;
        RECT 23.565 3.955 23.795 3.985 ;
        RECT 26.155 3.955 26.385 3.985 ;
        RECT 31.700 3.955 31.930 3.985 ;
        RECT 41.695 3.955 41.925 3.985 ;
        RECT 42.435 3.955 42.665 3.985 ;
        RECT 47.985 3.955 48.215 3.985 ;
        RECT 50.575 3.955 50.805 3.985 ;
        RECT 56.120 3.955 56.350 3.985 ;
        RECT 66.115 3.955 66.345 3.985 ;
        RECT 66.855 3.955 67.085 3.985 ;
        RECT 72.405 3.955 72.635 3.985 ;
        RECT 74.995 3.955 75.225 3.985 ;
        RECT 81.655 3.955 81.885 3.985 ;
        RECT 6.545 3.785 6.775 3.815 ;
        RECT 11.355 3.785 11.585 3.815 ;
        RECT 15.425 3.785 15.655 3.815 ;
        RECT 22.825 3.785 23.055 3.815 ;
        RECT 30.965 3.785 31.195 3.815 ;
        RECT 35.775 3.785 36.005 3.815 ;
        RECT 39.845 3.785 40.075 3.815 ;
        RECT 47.245 3.785 47.475 3.815 ;
        RECT 55.385 3.785 55.615 3.815 ;
        RECT 60.195 3.785 60.425 3.815 ;
        RECT 64.265 3.785 64.495 3.815 ;
        RECT 71.665 3.785 71.895 3.815 ;
        RECT 6.515 3.615 23.085 3.785 ;
        RECT 30.935 3.615 47.505 3.785 ;
        RECT 55.355 3.615 71.925 3.785 ;
        RECT 6.545 3.585 6.775 3.615 ;
        RECT 11.355 3.585 11.585 3.615 ;
        RECT 15.425 3.585 15.655 3.615 ;
        RECT 22.825 3.585 23.055 3.615 ;
        RECT 30.965 3.585 31.195 3.615 ;
        RECT 35.775 3.585 36.005 3.615 ;
        RECT 39.845 3.585 40.075 3.615 ;
        RECT 47.245 3.585 47.475 3.615 ;
        RECT 55.385 3.585 55.615 3.615 ;
        RECT 60.195 3.585 60.425 3.615 ;
        RECT 64.265 3.585 64.495 3.615 ;
        RECT 71.665 3.585 71.895 3.615 ;
        RECT 18.755 3.415 18.985 3.445 ;
        RECT 20.605 3.415 20.835 3.445 ;
        RECT 79.065 3.415 79.295 3.445 ;
        RECT 18.725 3.245 79.325 3.415 ;
        RECT 18.755 3.215 18.985 3.245 ;
        RECT 20.605 3.215 20.835 3.245 ;
        RECT 79.065 3.215 79.295 3.245 ;
        RECT 74.995 3.045 75.225 3.075 ;
        RECT 50.605 2.875 75.255 3.045 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.700 ;
        RECT 9.135 2.675 9.365 2.705 ;
        RECT 12.095 2.675 12.325 2.705 ;
        RECT 13.945 2.675 14.175 2.705 ;
        RECT 26.895 2.675 27.125 2.705 ;
        RECT 28.745 2.675 28.975 2.700 ;
        RECT 33.555 2.675 33.785 2.705 ;
        RECT 36.515 2.675 36.745 2.705 ;
        RECT 38.365 2.675 38.595 2.705 ;
        RECT 43.175 2.675 43.405 2.705 ;
        RECT 45.025 2.675 45.255 2.705 ;
        RECT 50.605 2.675 50.775 2.875 ;
        RECT 74.995 2.845 75.225 2.875 ;
        RECT 51.315 2.675 51.545 2.705 ;
        RECT 53.165 2.675 53.395 2.700 ;
        RECT 57.975 2.675 58.205 2.705 ;
        RECT 60.935 2.675 61.165 2.705 ;
        RECT 62.785 2.675 63.015 2.705 ;
        RECT 2.445 2.505 9.395 2.675 ;
        RECT 12.065 2.505 14.205 2.675 ;
        RECT 26.865 2.505 33.815 2.675 ;
        RECT 36.485 2.505 38.625 2.675 ;
        RECT 43.145 2.505 50.775 2.675 ;
        RECT 51.285 2.505 58.235 2.675 ;
        RECT 60.905 2.505 63.045 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.295 2.500 4.705 2.505 ;
        RECT 4.325 2.470 4.555 2.500 ;
        RECT 9.135 2.475 9.365 2.505 ;
        RECT 12.095 2.475 12.325 2.505 ;
        RECT 13.945 2.475 14.175 2.505 ;
        RECT 26.895 2.475 27.125 2.505 ;
        RECT 28.715 2.500 29.125 2.505 ;
        RECT 28.745 2.470 28.975 2.500 ;
        RECT 33.555 2.475 33.785 2.505 ;
        RECT 36.515 2.475 36.745 2.505 ;
        RECT 38.365 2.475 38.595 2.505 ;
        RECT 43.175 2.475 43.405 2.505 ;
        RECT 45.025 2.475 45.255 2.505 ;
        RECT 51.315 2.475 51.545 2.505 ;
        RECT 53.135 2.500 53.545 2.505 ;
        RECT 53.165 2.470 53.395 2.500 ;
        RECT 57.975 2.475 58.205 2.505 ;
        RECT 60.935 2.475 61.165 2.505 ;
        RECT 62.785 2.475 63.015 2.505 ;
        RECT 79.065 2.165 79.295 2.195 ;
        RECT 80.545 2.165 80.775 2.195 ;
        RECT 79.035 1.995 80.805 2.165 ;
        RECT 79.065 1.965 79.295 1.995 ;
        RECT 80.545 1.965 80.775 1.995 ;
        RECT 75.295 1.265 75.525 1.295 ;
        RECT 78.625 1.265 78.855 1.295 ;
        RECT 81.955 1.265 82.185 1.295 ;
        RECT 75.265 1.095 82.215 1.265 ;
        RECT 75.295 1.065 75.525 1.095 ;
        RECT 78.625 1.065 78.855 1.095 ;
        RECT 81.955 1.065 82.185 1.095 ;
  END
END TMRDFFSNQNX1






MACRO TMRDFFSNQX1
  CLASS CORE ;
  FOREIGN TMRDFFSNQX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 85.470 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN D
    ANTENNAGATEAREA 3.099750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 25.445 1.915 25.615 4.865 ;
        RECT 49.865 1.915 50.035 4.865 ;
      LAYER mcon ;
        RECT 1.025 2.875 1.195 3.045 ;
        RECT 25.445 2.875 25.615 3.045 ;
        RECT 49.865 2.875 50.035 3.045 ;
      LAYER met1 ;
        RECT 0.995 3.045 1.225 3.075 ;
        RECT 25.415 3.045 25.645 3.075 ;
        RECT 49.835 3.045 50.065 3.075 ;
        RECT 0.965 2.875 50.095 3.045 ;
        RECT 0.995 2.845 1.225 2.875 ;
        RECT 25.415 2.845 25.645 2.875 ;
        RECT 49.835 2.845 50.065 2.875 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.126300 ;
    PORT
      LAYER li1 ;
        RECT 5.465 1.915 5.635 4.865 ;
        RECT 14.745 4.710 14.915 4.865 ;
        RECT 14.715 4.535 14.915 4.710 ;
        RECT 14.715 1.915 14.885 4.535 ;
        RECT 29.885 1.915 30.055 4.865 ;
        RECT 39.165 4.710 39.335 4.865 ;
        RECT 39.135 4.535 39.335 4.710 ;
        RECT 39.135 1.915 39.305 4.535 ;
        RECT 54.305 1.915 54.475 4.865 ;
        RECT 63.585 4.710 63.755 4.865 ;
        RECT 63.555 4.535 63.755 4.710 ;
        RECT 63.555 1.915 63.725 4.535 ;
      LAYER mcon ;
        RECT 5.465 4.355 5.635 4.525 ;
        RECT 14.715 4.355 14.885 4.525 ;
        RECT 29.885 4.355 30.055 4.525 ;
        RECT 39.135 4.355 39.305 4.525 ;
        RECT 54.305 4.355 54.475 4.525 ;
        RECT 63.555 4.355 63.725 4.525 ;
      LAYER met1 ;
        RECT 5.435 4.525 5.665 4.555 ;
        RECT 14.685 4.525 14.915 4.555 ;
        RECT 29.855 4.525 30.085 4.555 ;
        RECT 39.105 4.525 39.335 4.555 ;
        RECT 54.275 4.525 54.505 4.555 ;
        RECT 63.525 4.525 63.755 4.555 ;
        RECT 5.405 4.355 63.785 4.525 ;
        RECT 5.435 4.325 5.665 4.355 ;
        RECT 14.685 4.325 14.915 4.355 ;
        RECT 29.855 4.325 30.085 4.355 ;
        RECT 39.105 4.325 39.335 4.355 ;
        RECT 54.275 4.325 54.505 4.355 ;
        RECT 63.525 4.325 63.755 4.355 ;
    END
  END CLK
  PIN SN
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 10.275 1.915 10.445 4.865 ;
        RECT 21.745 1.915 21.915 4.865 ;
        RECT 34.695 1.915 34.865 4.865 ;
        RECT 46.165 1.915 46.335 4.865 ;
        RECT 59.115 1.915 59.285 4.865 ;
        RECT 70.585 1.915 70.755 4.865 ;
      LAYER mcon ;
        RECT 10.275 2.135 10.445 2.305 ;
        RECT 21.745 2.135 21.915 2.305 ;
        RECT 34.695 2.135 34.865 2.305 ;
        RECT 46.165 2.135 46.335 2.305 ;
        RECT 59.115 2.135 59.285 2.305 ;
        RECT 70.585 2.135 70.755 2.305 ;
      LAYER met1 ;
        RECT 10.245 2.305 10.475 2.335 ;
        RECT 21.715 2.305 21.945 2.335 ;
        RECT 34.665 2.305 34.895 2.335 ;
        RECT 46.135 2.305 46.365 2.335 ;
        RECT 59.085 2.305 59.315 2.335 ;
        RECT 70.555 2.305 70.785 2.335 ;
        RECT 10.215 2.135 70.815 2.305 ;
        RECT 10.245 2.105 10.475 2.135 ;
        RECT 21.715 2.105 21.945 2.135 ;
        RECT 34.665 2.105 34.895 2.135 ;
        RECT 46.135 2.105 46.365 2.135 ;
        RECT 59.085 2.105 59.315 2.135 ;
        RECT 70.555 2.105 70.785 2.135 ;
    END
  END SN
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 85.905 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 85.640 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.335 5.215 4.505 7.230 ;
        RECT 5.215 5.555 5.385 7.230 ;
        RECT 6.095 5.555 6.265 7.230 ;
        RECT 6.975 5.555 7.145 7.230 ;
        RECT 7.970 4.110 8.310 7.230 ;
        RECT 9.145 5.215 9.315 7.230 ;
        RECT 10.025 5.555 10.195 7.230 ;
        RECT 10.905 5.555 11.075 7.230 ;
        RECT 11.785 5.555 11.955 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.655 5.135 13.825 7.230 ;
        RECT 14.535 5.555 14.705 7.230 ;
        RECT 15.415 5.555 15.585 7.230 ;
        RECT 16.110 4.110 16.450 7.230 ;
        RECT 16.985 5.135 17.155 7.230 ;
        RECT 17.865 5.555 18.035 7.230 ;
        RECT 18.745 5.555 18.915 7.230 ;
        RECT 19.440 4.110 19.780 7.230 ;
        RECT 20.615 5.215 20.785 7.230 ;
        RECT 21.495 5.555 21.665 7.230 ;
        RECT 22.375 5.555 22.545 7.230 ;
        RECT 23.255 5.555 23.425 7.230 ;
        RECT 24.250 4.110 24.590 7.230 ;
        RECT 25.125 5.135 25.295 7.230 ;
        RECT 26.005 5.555 26.175 7.230 ;
        RECT 26.885 5.555 27.055 7.230 ;
        RECT 27.580 4.110 27.920 7.230 ;
        RECT 28.755 5.215 28.925 7.230 ;
        RECT 29.635 5.555 29.805 7.230 ;
        RECT 30.515 5.555 30.685 7.230 ;
        RECT 31.395 5.555 31.565 7.230 ;
        RECT 32.390 4.110 32.730 7.230 ;
        RECT 33.565 5.215 33.735 7.230 ;
        RECT 34.445 5.555 34.615 7.230 ;
        RECT 35.325 5.555 35.495 7.230 ;
        RECT 36.205 5.555 36.375 7.230 ;
        RECT 37.200 4.110 37.540 7.230 ;
        RECT 38.075 5.135 38.245 7.230 ;
        RECT 38.955 5.555 39.125 7.230 ;
        RECT 39.835 5.555 40.005 7.230 ;
        RECT 40.530 4.110 40.870 7.230 ;
        RECT 41.405 5.135 41.575 7.230 ;
        RECT 42.285 5.555 42.455 7.230 ;
        RECT 43.165 5.555 43.335 7.230 ;
        RECT 43.860 4.110 44.200 7.230 ;
        RECT 45.035 5.215 45.205 7.230 ;
        RECT 45.915 5.555 46.085 7.230 ;
        RECT 46.795 5.555 46.965 7.230 ;
        RECT 47.675 5.555 47.845 7.230 ;
        RECT 48.670 4.110 49.010 7.230 ;
        RECT 49.545 5.135 49.715 7.230 ;
        RECT 50.425 5.555 50.595 7.230 ;
        RECT 51.305 5.555 51.475 7.230 ;
        RECT 52.000 4.110 52.340 7.230 ;
        RECT 53.175 5.215 53.345 7.230 ;
        RECT 54.055 5.555 54.225 7.230 ;
        RECT 54.935 5.555 55.105 7.230 ;
        RECT 55.815 5.555 55.985 7.230 ;
        RECT 56.810 4.110 57.150 7.230 ;
        RECT 57.985 5.215 58.155 7.230 ;
        RECT 58.865 5.555 59.035 7.230 ;
        RECT 59.745 5.555 59.915 7.230 ;
        RECT 60.625 5.555 60.795 7.230 ;
        RECT 61.620 4.110 61.960 7.230 ;
        RECT 62.495 5.135 62.665 7.230 ;
        RECT 63.375 5.555 63.545 7.230 ;
        RECT 64.255 5.555 64.425 7.230 ;
        RECT 64.950 4.110 65.290 7.230 ;
        RECT 65.825 5.135 65.995 7.230 ;
        RECT 66.705 5.555 66.875 7.230 ;
        RECT 67.585 5.555 67.755 7.230 ;
        RECT 68.280 4.110 68.620 7.230 ;
        RECT 69.455 5.215 69.625 7.230 ;
        RECT 70.335 5.555 70.505 7.230 ;
        RECT 71.215 5.555 71.385 7.230 ;
        RECT 72.095 5.555 72.265 7.230 ;
        RECT 73.090 4.110 73.430 7.230 ;
        RECT 73.965 5.125 74.135 7.230 ;
        RECT 74.845 5.555 75.015 7.230 ;
        RECT 75.725 5.125 75.895 7.230 ;
        RECT 76.420 4.110 76.760 7.230 ;
        RECT 79.750 4.110 80.090 7.230 ;
        RECT 83.080 4.110 83.420 7.230 ;
        RECT 83.840 5.185 84.010 7.230 ;
        RECT 84.720 5.185 84.890 7.230 ;
        RECT 85.300 4.110 85.640 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.515 7.315 29.685 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.625 7.315 30.795 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.845 7.315 33.015 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.435 7.315 35.605 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.175 7.315 36.345 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
        RECT 38.765 7.315 38.935 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.505 7.315 39.675 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 42.835 7.315 43.005 7.485 ;
        RECT 43.205 7.315 43.375 7.485 ;
        RECT 43.575 7.315 43.745 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 47.645 7.315 47.815 7.485 ;
        RECT 48.015 7.315 48.185 7.485 ;
        RECT 48.385 7.315 48.555 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 50.975 7.315 51.145 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 51.715 7.315 51.885 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 52.825 7.315 52.995 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.305 7.315 54.475 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.525 7.315 56.695 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 57.635 7.315 57.805 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 60.965 7.315 61.135 7.485 ;
        RECT 61.335 7.315 61.505 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.445 7.315 62.615 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.295 7.315 64.465 7.485 ;
        RECT 64.665 7.315 64.835 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.255 7.315 67.425 7.485 ;
        RECT 67.625 7.315 67.795 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.475 7.315 69.645 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 70.955 7.315 71.125 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.065 7.315 72.235 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
        RECT 74.285 7.315 74.455 7.485 ;
        RECT 74.655 7.315 74.825 7.485 ;
        RECT 75.025 7.315 75.195 7.485 ;
        RECT 75.395 7.315 75.565 7.485 ;
        RECT 75.765 7.315 75.935 7.485 ;
        RECT 76.135 7.315 76.305 7.485 ;
        RECT 76.875 7.315 77.045 7.485 ;
        RECT 77.245 7.315 77.415 7.485 ;
        RECT 77.615 7.315 77.785 7.485 ;
        RECT 77.985 7.315 78.155 7.485 ;
        RECT 78.355 7.315 78.525 7.485 ;
        RECT 78.725 7.315 78.895 7.485 ;
        RECT 79.095 7.315 79.265 7.485 ;
        RECT 79.465 7.315 79.635 7.485 ;
        RECT 80.205 7.315 80.375 7.485 ;
        RECT 80.575 7.315 80.745 7.485 ;
        RECT 80.945 7.315 81.115 7.485 ;
        RECT 81.315 7.315 81.485 7.485 ;
        RECT 81.685 7.315 81.855 7.485 ;
        RECT 82.055 7.315 82.225 7.485 ;
        RECT 82.425 7.315 82.595 7.485 ;
        RECT 82.795 7.315 82.965 7.485 ;
        RECT 83.535 7.315 83.705 7.485 ;
        RECT 83.905 7.315 84.075 7.485 ;
        RECT 84.275 7.315 84.445 7.485 ;
        RECT 84.645 7.315 84.815 7.485 ;
        RECT 85.015 7.315 85.185 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 85.640 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 85.640 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 4.320 0.170 4.490 1.130 ;
        RECT 7.970 0.170 8.310 2.720 ;
        RECT 9.130 0.170 9.300 1.130 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 14.045 0.170 14.215 1.120 ;
        RECT 16.110 0.170 16.450 2.720 ;
        RECT 17.375 0.170 17.545 1.120 ;
        RECT 19.440 0.170 19.780 2.720 ;
        RECT 20.600 0.170 20.770 1.130 ;
        RECT 24.250 0.170 24.590 2.720 ;
        RECT 25.515 0.170 25.685 1.120 ;
        RECT 27.580 0.170 27.920 2.720 ;
        RECT 28.740 0.170 28.910 1.130 ;
        RECT 32.390 0.170 32.730 2.720 ;
        RECT 33.550 0.170 33.720 1.130 ;
        RECT 37.200 0.170 37.540 2.720 ;
        RECT 38.465 0.170 38.635 1.120 ;
        RECT 40.530 0.170 40.870 2.720 ;
        RECT 41.795 0.170 41.965 1.120 ;
        RECT 43.860 0.170 44.200 2.720 ;
        RECT 45.020 0.170 45.190 1.130 ;
        RECT 48.670 0.170 49.010 2.720 ;
        RECT 49.935 0.170 50.105 1.120 ;
        RECT 52.000 0.170 52.340 2.720 ;
        RECT 53.160 0.170 53.330 1.130 ;
        RECT 56.810 0.170 57.150 2.720 ;
        RECT 57.970 0.170 58.140 1.130 ;
        RECT 61.620 0.170 61.960 2.720 ;
        RECT 62.885 0.170 63.055 1.120 ;
        RECT 64.950 0.170 65.290 2.720 ;
        RECT 66.215 0.170 66.385 1.120 ;
        RECT 68.280 0.170 68.620 2.720 ;
        RECT 69.440 0.170 69.610 1.130 ;
        RECT 73.090 0.170 73.430 2.720 ;
        RECT 74.355 0.170 74.525 1.120 ;
        RECT 76.420 0.170 76.760 2.720 ;
        RECT 77.685 0.170 77.855 1.120 ;
        RECT 79.750 0.170 80.090 2.720 ;
        RECT 81.015 0.170 81.185 1.120 ;
        RECT 83.080 0.170 83.420 2.720 ;
        RECT 83.795 0.620 83.965 1.750 ;
        RECT 84.765 0.620 84.935 1.750 ;
        RECT 83.795 0.450 84.935 0.620 ;
        RECT 83.795 0.170 83.965 0.450 ;
        RECT 84.280 0.170 84.450 0.450 ;
        RECT 84.765 0.170 84.935 0.450 ;
        RECT 85.300 0.170 85.640 2.720 ;
        RECT -0.170 -0.170 85.640 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.515 -0.085 29.685 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.625 -0.085 30.795 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.845 -0.085 33.015 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.435 -0.085 35.605 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.175 -0.085 36.345 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
        RECT 38.765 -0.085 38.935 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.505 -0.085 39.675 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 42.835 -0.085 43.005 0.085 ;
        RECT 43.205 -0.085 43.375 0.085 ;
        RECT 43.575 -0.085 43.745 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 47.645 -0.085 47.815 0.085 ;
        RECT 48.015 -0.085 48.185 0.085 ;
        RECT 48.385 -0.085 48.555 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 50.975 -0.085 51.145 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 51.715 -0.085 51.885 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 52.825 -0.085 52.995 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.305 -0.085 54.475 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.525 -0.085 56.695 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 57.635 -0.085 57.805 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 60.965 -0.085 61.135 0.085 ;
        RECT 61.335 -0.085 61.505 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.445 -0.085 62.615 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.295 -0.085 64.465 0.085 ;
        RECT 64.665 -0.085 64.835 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.255 -0.085 67.425 0.085 ;
        RECT 67.625 -0.085 67.795 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.475 -0.085 69.645 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 70.955 -0.085 71.125 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.065 -0.085 72.235 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
        RECT 74.285 -0.085 74.455 0.085 ;
        RECT 74.655 -0.085 74.825 0.085 ;
        RECT 75.025 -0.085 75.195 0.085 ;
        RECT 75.395 -0.085 75.565 0.085 ;
        RECT 75.765 -0.085 75.935 0.085 ;
        RECT 76.135 -0.085 76.305 0.085 ;
        RECT 76.875 -0.085 77.045 0.085 ;
        RECT 77.245 -0.085 77.415 0.085 ;
        RECT 77.615 -0.085 77.785 0.085 ;
        RECT 77.985 -0.085 78.155 0.085 ;
        RECT 78.355 -0.085 78.525 0.085 ;
        RECT 78.725 -0.085 78.895 0.085 ;
        RECT 79.095 -0.085 79.265 0.085 ;
        RECT 79.465 -0.085 79.635 0.085 ;
        RECT 80.205 -0.085 80.375 0.085 ;
        RECT 80.575 -0.085 80.745 0.085 ;
        RECT 80.945 -0.085 81.115 0.085 ;
        RECT 81.315 -0.085 81.485 0.085 ;
        RECT 81.685 -0.085 81.855 0.085 ;
        RECT 82.055 -0.085 82.225 0.085 ;
        RECT 82.425 -0.085 82.595 0.085 ;
        RECT 82.795 -0.085 82.965 0.085 ;
        RECT 83.535 -0.085 83.705 0.085 ;
        RECT 83.905 -0.085 84.075 0.085 ;
        RECT 84.275 -0.085 84.445 0.085 ;
        RECT 84.645 -0.085 84.815 0.085 ;
        RECT 85.015 -0.085 85.185 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 85.640 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.775 5.240 4.945 7.020 ;
        RECT 5.655 5.240 5.825 7.020 ;
        RECT 6.535 5.240 6.705 7.020 ;
        RECT 9.585 5.240 9.755 7.020 ;
        RECT 10.465 5.240 10.635 7.020 ;
        RECT 11.345 5.240 11.515 7.020 ;
        RECT 14.095 5.285 14.265 7.020 ;
        RECT 14.975 5.285 15.145 7.020 ;
        RECT 17.425 5.285 17.595 7.020 ;
        RECT 18.305 5.285 18.475 7.020 ;
        RECT 4.775 5.070 7.485 5.240 ;
        RECT 9.585 5.070 12.295 5.240 ;
        RECT 14.095 5.115 15.625 5.285 ;
        RECT 17.425 5.115 18.955 5.285 ;
        RECT 4.355 1.915 4.525 4.865 ;
        RECT 6.575 1.915 6.745 4.865 ;
        RECT 7.315 4.235 7.485 5.070 ;
        RECT 7.310 3.905 7.485 4.235 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 3.835 1.675 4.005 1.755 ;
        RECT 4.805 1.675 4.975 1.755 ;
        RECT 5.775 1.675 5.945 1.755 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 3.835 1.505 5.945 1.675 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 3.835 0.375 4.005 1.505 ;
        RECT 4.805 0.625 4.975 1.505 ;
        RECT 5.775 1.425 5.945 1.505 ;
        RECT 5.295 1.080 5.465 1.160 ;
        RECT 6.345 1.080 6.515 1.755 ;
        RECT 7.315 1.750 7.485 3.905 ;
        RECT 9.165 1.915 9.335 4.865 ;
        RECT 11.385 1.915 11.555 4.865 ;
        RECT 5.295 0.910 6.515 1.080 ;
        RECT 5.295 0.830 5.465 0.910 ;
        RECT 5.775 0.625 5.945 0.705 ;
        RECT 4.805 0.455 5.945 0.625 ;
        RECT 4.805 0.375 4.975 0.455 ;
        RECT 5.775 0.375 5.945 0.455 ;
        RECT 6.345 0.625 6.515 0.910 ;
        RECT 6.830 1.580 7.485 1.750 ;
        RECT 8.645 1.675 8.815 1.755 ;
        RECT 9.615 1.675 9.785 1.755 ;
        RECT 10.585 1.675 10.755 1.755 ;
        RECT 6.830 0.845 7.000 1.580 ;
        RECT 8.645 1.505 10.755 1.675 ;
        RECT 7.315 0.625 7.485 1.395 ;
        RECT 6.345 0.455 7.485 0.625 ;
        RECT 6.345 0.375 6.515 0.455 ;
        RECT 7.315 0.375 7.485 0.455 ;
        RECT 8.645 0.375 8.815 1.505 ;
        RECT 9.615 0.625 9.785 1.505 ;
        RECT 10.585 1.425 10.755 1.505 ;
        RECT 10.105 1.080 10.275 1.160 ;
        RECT 11.155 1.080 11.325 1.755 ;
        RECT 12.125 1.750 12.295 5.070 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 10.105 0.910 11.325 1.080 ;
        RECT 10.105 0.830 10.275 0.910 ;
        RECT 10.585 0.625 10.755 0.705 ;
        RECT 9.615 0.455 10.755 0.625 ;
        RECT 9.615 0.375 9.785 0.455 ;
        RECT 10.585 0.375 10.755 0.455 ;
        RECT 11.155 0.625 11.325 0.910 ;
        RECT 11.640 1.580 12.295 1.750 ;
        RECT 13.560 1.665 13.730 1.745 ;
        RECT 14.530 1.665 14.700 1.745 ;
        RECT 15.455 1.740 15.625 5.115 ;
        RECT 17.305 1.915 17.475 4.865 ;
        RECT 18.075 4.710 18.245 4.865 ;
        RECT 18.045 4.535 18.245 4.710 ;
        RECT 18.045 1.915 18.215 4.535 ;
        RECT 11.640 0.845 11.810 1.580 ;
        RECT 13.560 1.495 14.700 1.665 ;
        RECT 12.125 0.625 12.295 1.395 ;
        RECT 11.155 0.455 12.295 0.625 ;
        RECT 11.155 0.375 11.325 0.455 ;
        RECT 12.125 0.375 12.295 0.455 ;
        RECT 13.560 0.365 13.730 1.495 ;
        RECT 14.530 0.615 14.700 1.495 ;
        RECT 15.015 1.570 15.625 1.740 ;
        RECT 16.890 1.665 17.060 1.745 ;
        RECT 17.860 1.665 18.030 1.745 ;
        RECT 18.785 1.740 18.955 5.115 ;
        RECT 21.055 5.240 21.225 7.020 ;
        RECT 21.935 5.240 22.105 7.020 ;
        RECT 22.815 5.240 22.985 7.020 ;
        RECT 25.565 5.285 25.735 7.020 ;
        RECT 26.445 5.285 26.615 7.020 ;
        RECT 21.055 5.070 23.765 5.240 ;
        RECT 25.565 5.115 27.095 5.285 ;
        RECT 20.635 1.915 20.805 4.865 ;
        RECT 22.855 1.915 23.025 4.865 ;
        RECT 15.015 0.835 15.185 1.570 ;
        RECT 16.890 1.495 18.030 1.665 ;
        RECT 15.500 0.615 15.670 1.385 ;
        RECT 14.530 0.445 15.670 0.615 ;
        RECT 14.530 0.365 14.700 0.445 ;
        RECT 15.500 0.365 15.670 0.445 ;
        RECT 16.890 0.365 17.060 1.495 ;
        RECT 17.860 0.615 18.030 1.495 ;
        RECT 18.345 1.570 18.955 1.740 ;
        RECT 20.115 1.675 20.285 1.755 ;
        RECT 21.085 1.675 21.255 1.755 ;
        RECT 22.055 1.675 22.225 1.755 ;
        RECT 18.345 0.835 18.515 1.570 ;
        RECT 20.115 1.505 22.225 1.675 ;
        RECT 18.830 0.615 19.000 1.385 ;
        RECT 17.860 0.445 19.000 0.615 ;
        RECT 17.860 0.365 18.030 0.445 ;
        RECT 18.830 0.365 19.000 0.445 ;
        RECT 20.115 0.375 20.285 1.505 ;
        RECT 21.085 0.625 21.255 1.505 ;
        RECT 22.055 1.425 22.225 1.505 ;
        RECT 21.575 1.080 21.745 1.160 ;
        RECT 22.625 1.080 22.795 1.755 ;
        RECT 23.595 1.750 23.765 5.070 ;
        RECT 26.215 4.710 26.385 4.865 ;
        RECT 26.185 4.535 26.385 4.710 ;
        RECT 26.185 1.915 26.355 4.535 ;
        RECT 21.575 0.910 22.795 1.080 ;
        RECT 21.575 0.830 21.745 0.910 ;
        RECT 22.055 0.625 22.225 0.705 ;
        RECT 21.085 0.455 22.225 0.625 ;
        RECT 21.085 0.375 21.255 0.455 ;
        RECT 22.055 0.375 22.225 0.455 ;
        RECT 22.625 0.625 22.795 0.910 ;
        RECT 23.110 1.580 23.765 1.750 ;
        RECT 25.030 1.665 25.200 1.745 ;
        RECT 26.000 1.665 26.170 1.745 ;
        RECT 26.925 1.740 27.095 5.115 ;
        RECT 29.195 5.240 29.365 7.020 ;
        RECT 30.075 5.240 30.245 7.020 ;
        RECT 30.955 5.240 31.125 7.020 ;
        RECT 34.005 5.240 34.175 7.020 ;
        RECT 34.885 5.240 35.055 7.020 ;
        RECT 35.765 5.240 35.935 7.020 ;
        RECT 38.515 5.285 38.685 7.020 ;
        RECT 39.395 5.285 39.565 7.020 ;
        RECT 41.845 5.285 42.015 7.020 ;
        RECT 42.725 5.285 42.895 7.020 ;
        RECT 29.195 5.070 31.905 5.240 ;
        RECT 34.005 5.070 36.715 5.240 ;
        RECT 38.515 5.115 40.045 5.285 ;
        RECT 41.845 5.115 43.375 5.285 ;
        RECT 28.775 1.915 28.945 4.865 ;
        RECT 30.995 1.915 31.165 4.865 ;
        RECT 31.735 4.235 31.905 5.070 ;
        RECT 31.730 3.905 31.905 4.235 ;
        RECT 23.110 0.845 23.280 1.580 ;
        RECT 25.030 1.495 26.170 1.665 ;
        RECT 23.595 0.625 23.765 1.395 ;
        RECT 22.625 0.455 23.765 0.625 ;
        RECT 22.625 0.375 22.795 0.455 ;
        RECT 23.595 0.375 23.765 0.455 ;
        RECT 25.030 0.365 25.200 1.495 ;
        RECT 26.000 0.615 26.170 1.495 ;
        RECT 26.485 1.570 27.095 1.740 ;
        RECT 28.255 1.675 28.425 1.755 ;
        RECT 29.225 1.675 29.395 1.755 ;
        RECT 30.195 1.675 30.365 1.755 ;
        RECT 26.485 0.835 26.655 1.570 ;
        RECT 28.255 1.505 30.365 1.675 ;
        RECT 26.970 0.615 27.140 1.385 ;
        RECT 26.000 0.445 27.140 0.615 ;
        RECT 26.000 0.365 26.170 0.445 ;
        RECT 26.970 0.365 27.140 0.445 ;
        RECT 28.255 0.375 28.425 1.505 ;
        RECT 29.225 0.625 29.395 1.505 ;
        RECT 30.195 1.425 30.365 1.505 ;
        RECT 29.715 1.080 29.885 1.160 ;
        RECT 30.765 1.080 30.935 1.755 ;
        RECT 31.735 1.750 31.905 3.905 ;
        RECT 33.585 1.915 33.755 4.865 ;
        RECT 35.805 1.915 35.975 4.865 ;
        RECT 29.715 0.910 30.935 1.080 ;
        RECT 29.715 0.830 29.885 0.910 ;
        RECT 30.195 0.625 30.365 0.705 ;
        RECT 29.225 0.455 30.365 0.625 ;
        RECT 29.225 0.375 29.395 0.455 ;
        RECT 30.195 0.375 30.365 0.455 ;
        RECT 30.765 0.625 30.935 0.910 ;
        RECT 31.250 1.580 31.905 1.750 ;
        RECT 33.065 1.675 33.235 1.755 ;
        RECT 34.035 1.675 34.205 1.755 ;
        RECT 35.005 1.675 35.175 1.755 ;
        RECT 31.250 0.845 31.420 1.580 ;
        RECT 33.065 1.505 35.175 1.675 ;
        RECT 31.735 0.625 31.905 1.395 ;
        RECT 30.765 0.455 31.905 0.625 ;
        RECT 30.765 0.375 30.935 0.455 ;
        RECT 31.735 0.375 31.905 0.455 ;
        RECT 33.065 0.375 33.235 1.505 ;
        RECT 34.035 0.625 34.205 1.505 ;
        RECT 35.005 1.425 35.175 1.505 ;
        RECT 34.525 1.080 34.695 1.160 ;
        RECT 35.575 1.080 35.745 1.755 ;
        RECT 36.545 1.750 36.715 5.070 ;
        RECT 38.395 1.915 38.565 4.865 ;
        RECT 34.525 0.910 35.745 1.080 ;
        RECT 34.525 0.830 34.695 0.910 ;
        RECT 35.005 0.625 35.175 0.705 ;
        RECT 34.035 0.455 35.175 0.625 ;
        RECT 34.035 0.375 34.205 0.455 ;
        RECT 35.005 0.375 35.175 0.455 ;
        RECT 35.575 0.625 35.745 0.910 ;
        RECT 36.060 1.580 36.715 1.750 ;
        RECT 37.980 1.665 38.150 1.745 ;
        RECT 38.950 1.665 39.120 1.745 ;
        RECT 39.875 1.740 40.045 5.115 ;
        RECT 41.725 1.915 41.895 4.865 ;
        RECT 42.495 4.710 42.665 4.865 ;
        RECT 42.465 4.535 42.665 4.710 ;
        RECT 42.465 1.915 42.635 4.535 ;
        RECT 36.060 0.845 36.230 1.580 ;
        RECT 37.980 1.495 39.120 1.665 ;
        RECT 36.545 0.625 36.715 1.395 ;
        RECT 35.575 0.455 36.715 0.625 ;
        RECT 35.575 0.375 35.745 0.455 ;
        RECT 36.545 0.375 36.715 0.455 ;
        RECT 37.980 0.365 38.150 1.495 ;
        RECT 38.950 0.615 39.120 1.495 ;
        RECT 39.435 1.570 40.045 1.740 ;
        RECT 41.310 1.665 41.480 1.745 ;
        RECT 42.280 1.665 42.450 1.745 ;
        RECT 43.205 1.740 43.375 5.115 ;
        RECT 45.475 5.240 45.645 7.020 ;
        RECT 46.355 5.240 46.525 7.020 ;
        RECT 47.235 5.240 47.405 7.020 ;
        RECT 49.985 5.285 50.155 7.020 ;
        RECT 50.865 5.285 51.035 7.020 ;
        RECT 45.475 5.070 48.185 5.240 ;
        RECT 49.985 5.115 51.515 5.285 ;
        RECT 45.055 1.915 45.225 4.865 ;
        RECT 47.275 1.915 47.445 4.865 ;
        RECT 39.435 0.835 39.605 1.570 ;
        RECT 41.310 1.495 42.450 1.665 ;
        RECT 39.920 0.615 40.090 1.385 ;
        RECT 38.950 0.445 40.090 0.615 ;
        RECT 38.950 0.365 39.120 0.445 ;
        RECT 39.920 0.365 40.090 0.445 ;
        RECT 41.310 0.365 41.480 1.495 ;
        RECT 42.280 0.615 42.450 1.495 ;
        RECT 42.765 1.570 43.375 1.740 ;
        RECT 44.535 1.675 44.705 1.755 ;
        RECT 45.505 1.675 45.675 1.755 ;
        RECT 46.475 1.675 46.645 1.755 ;
        RECT 42.765 0.835 42.935 1.570 ;
        RECT 44.535 1.505 46.645 1.675 ;
        RECT 43.250 0.615 43.420 1.385 ;
        RECT 42.280 0.445 43.420 0.615 ;
        RECT 42.280 0.365 42.450 0.445 ;
        RECT 43.250 0.365 43.420 0.445 ;
        RECT 44.535 0.375 44.705 1.505 ;
        RECT 45.505 0.625 45.675 1.505 ;
        RECT 46.475 1.425 46.645 1.505 ;
        RECT 45.995 1.080 46.165 1.160 ;
        RECT 47.045 1.080 47.215 1.755 ;
        RECT 48.015 1.750 48.185 5.070 ;
        RECT 50.635 4.710 50.805 4.865 ;
        RECT 50.605 4.535 50.805 4.710 ;
        RECT 50.605 1.915 50.775 4.535 ;
        RECT 45.995 0.910 47.215 1.080 ;
        RECT 45.995 0.830 46.165 0.910 ;
        RECT 46.475 0.625 46.645 0.705 ;
        RECT 45.505 0.455 46.645 0.625 ;
        RECT 45.505 0.375 45.675 0.455 ;
        RECT 46.475 0.375 46.645 0.455 ;
        RECT 47.045 0.625 47.215 0.910 ;
        RECT 47.530 1.580 48.185 1.750 ;
        RECT 49.450 1.665 49.620 1.745 ;
        RECT 50.420 1.665 50.590 1.745 ;
        RECT 51.345 1.740 51.515 5.115 ;
        RECT 53.615 5.240 53.785 7.020 ;
        RECT 54.495 5.240 54.665 7.020 ;
        RECT 55.375 5.240 55.545 7.020 ;
        RECT 58.425 5.240 58.595 7.020 ;
        RECT 59.305 5.240 59.475 7.020 ;
        RECT 60.185 5.240 60.355 7.020 ;
        RECT 62.935 5.285 63.105 7.020 ;
        RECT 63.815 5.285 63.985 7.020 ;
        RECT 66.265 5.285 66.435 7.020 ;
        RECT 67.145 5.285 67.315 7.020 ;
        RECT 53.615 5.070 56.325 5.240 ;
        RECT 58.425 5.070 61.135 5.240 ;
        RECT 62.935 5.115 64.465 5.285 ;
        RECT 66.265 5.115 67.795 5.285 ;
        RECT 53.195 1.915 53.365 4.865 ;
        RECT 55.415 1.915 55.585 4.865 ;
        RECT 56.155 4.235 56.325 5.070 ;
        RECT 56.150 3.905 56.325 4.235 ;
        RECT 47.530 0.845 47.700 1.580 ;
        RECT 49.450 1.495 50.590 1.665 ;
        RECT 48.015 0.625 48.185 1.395 ;
        RECT 47.045 0.455 48.185 0.625 ;
        RECT 47.045 0.375 47.215 0.455 ;
        RECT 48.015 0.375 48.185 0.455 ;
        RECT 49.450 0.365 49.620 1.495 ;
        RECT 50.420 0.615 50.590 1.495 ;
        RECT 50.905 1.570 51.515 1.740 ;
        RECT 52.675 1.675 52.845 1.755 ;
        RECT 53.645 1.675 53.815 1.755 ;
        RECT 54.615 1.675 54.785 1.755 ;
        RECT 50.905 0.835 51.075 1.570 ;
        RECT 52.675 1.505 54.785 1.675 ;
        RECT 51.390 0.615 51.560 1.385 ;
        RECT 50.420 0.445 51.560 0.615 ;
        RECT 50.420 0.365 50.590 0.445 ;
        RECT 51.390 0.365 51.560 0.445 ;
        RECT 52.675 0.375 52.845 1.505 ;
        RECT 53.645 0.625 53.815 1.505 ;
        RECT 54.615 1.425 54.785 1.505 ;
        RECT 54.135 1.080 54.305 1.160 ;
        RECT 55.185 1.080 55.355 1.755 ;
        RECT 56.155 1.750 56.325 3.905 ;
        RECT 58.005 1.915 58.175 4.865 ;
        RECT 60.225 1.915 60.395 4.865 ;
        RECT 54.135 0.910 55.355 1.080 ;
        RECT 54.135 0.830 54.305 0.910 ;
        RECT 54.615 0.625 54.785 0.705 ;
        RECT 53.645 0.455 54.785 0.625 ;
        RECT 53.645 0.375 53.815 0.455 ;
        RECT 54.615 0.375 54.785 0.455 ;
        RECT 55.185 0.625 55.355 0.910 ;
        RECT 55.670 1.580 56.325 1.750 ;
        RECT 57.485 1.675 57.655 1.755 ;
        RECT 58.455 1.675 58.625 1.755 ;
        RECT 59.425 1.675 59.595 1.755 ;
        RECT 55.670 0.845 55.840 1.580 ;
        RECT 57.485 1.505 59.595 1.675 ;
        RECT 56.155 0.625 56.325 1.395 ;
        RECT 55.185 0.455 56.325 0.625 ;
        RECT 55.185 0.375 55.355 0.455 ;
        RECT 56.155 0.375 56.325 0.455 ;
        RECT 57.485 0.375 57.655 1.505 ;
        RECT 58.455 0.625 58.625 1.505 ;
        RECT 59.425 1.425 59.595 1.505 ;
        RECT 58.945 1.080 59.115 1.160 ;
        RECT 59.995 1.080 60.165 1.755 ;
        RECT 60.965 1.750 61.135 5.070 ;
        RECT 62.815 1.915 62.985 4.865 ;
        RECT 58.945 0.910 60.165 1.080 ;
        RECT 58.945 0.830 59.115 0.910 ;
        RECT 59.425 0.625 59.595 0.705 ;
        RECT 58.455 0.455 59.595 0.625 ;
        RECT 58.455 0.375 58.625 0.455 ;
        RECT 59.425 0.375 59.595 0.455 ;
        RECT 59.995 0.625 60.165 0.910 ;
        RECT 60.480 1.580 61.135 1.750 ;
        RECT 62.400 1.665 62.570 1.745 ;
        RECT 63.370 1.665 63.540 1.745 ;
        RECT 64.295 1.740 64.465 5.115 ;
        RECT 66.145 1.915 66.315 4.865 ;
        RECT 66.915 4.710 67.085 4.865 ;
        RECT 66.885 4.535 67.085 4.710 ;
        RECT 66.885 1.915 67.055 4.535 ;
        RECT 60.480 0.845 60.650 1.580 ;
        RECT 62.400 1.495 63.540 1.665 ;
        RECT 60.965 0.625 61.135 1.395 ;
        RECT 59.995 0.455 61.135 0.625 ;
        RECT 59.995 0.375 60.165 0.455 ;
        RECT 60.965 0.375 61.135 0.455 ;
        RECT 62.400 0.365 62.570 1.495 ;
        RECT 63.370 0.615 63.540 1.495 ;
        RECT 63.855 1.570 64.465 1.740 ;
        RECT 65.730 1.665 65.900 1.745 ;
        RECT 66.700 1.665 66.870 1.745 ;
        RECT 67.625 1.740 67.795 5.115 ;
        RECT 69.895 5.240 70.065 7.020 ;
        RECT 70.775 5.240 70.945 7.020 ;
        RECT 71.655 5.240 71.825 7.020 ;
        RECT 74.405 6.825 74.585 6.995 ;
        RECT 74.405 5.295 74.575 6.825 ;
        RECT 75.285 5.295 75.455 6.995 ;
        RECT 69.895 5.070 72.605 5.240 ;
        RECT 74.405 5.125 75.455 5.295 ;
        RECT 69.475 1.915 69.645 4.975 ;
        RECT 71.695 1.915 71.865 4.865 ;
        RECT 63.855 0.835 64.025 1.570 ;
        RECT 65.730 1.495 66.870 1.665 ;
        RECT 64.340 0.615 64.510 1.385 ;
        RECT 63.370 0.445 64.510 0.615 ;
        RECT 63.370 0.365 63.540 0.445 ;
        RECT 64.340 0.365 64.510 0.445 ;
        RECT 65.730 0.365 65.900 1.495 ;
        RECT 66.700 0.615 66.870 1.495 ;
        RECT 67.185 1.570 67.795 1.740 ;
        RECT 68.955 1.675 69.125 1.755 ;
        RECT 69.925 1.675 70.095 1.755 ;
        RECT 70.895 1.675 71.065 1.755 ;
        RECT 67.185 0.835 67.355 1.570 ;
        RECT 68.955 1.505 71.065 1.675 ;
        RECT 67.670 0.615 67.840 1.385 ;
        RECT 66.700 0.445 67.840 0.615 ;
        RECT 66.700 0.365 66.870 0.445 ;
        RECT 67.670 0.365 67.840 0.445 ;
        RECT 68.955 0.375 69.125 1.505 ;
        RECT 69.925 0.625 70.095 1.505 ;
        RECT 70.895 1.425 71.065 1.505 ;
        RECT 70.415 1.080 70.585 1.160 ;
        RECT 71.465 1.080 71.635 1.755 ;
        RECT 72.435 1.750 72.605 5.070 ;
        RECT 75.285 5.045 75.455 5.125 ;
        RECT 77.285 6.825 79.215 6.995 ;
        RECT 77.285 5.045 77.455 6.825 ;
        RECT 77.725 5.295 77.895 6.565 ;
        RECT 78.165 5.555 78.335 6.825 ;
        RECT 78.605 5.295 78.775 6.565 ;
        RECT 79.045 5.375 79.215 6.825 ;
        RECT 80.625 6.825 82.555 6.995 ;
        RECT 77.725 5.125 78.775 5.295 ;
        RECT 78.605 5.045 78.775 5.125 ;
        RECT 80.625 5.045 80.795 6.825 ;
        RECT 81.065 5.295 81.235 6.565 ;
        RECT 81.505 5.555 81.675 6.825 ;
        RECT 81.945 5.295 82.115 6.565 ;
        RECT 82.385 5.555 82.555 6.825 ;
        RECT 81.065 5.125 82.595 5.295 ;
        RECT 73.915 1.915 74.085 4.870 ;
        RECT 75.065 4.710 75.235 4.870 ;
        RECT 75.025 4.540 75.235 4.710 ;
        RECT 75.025 1.915 75.195 4.540 ;
        RECT 77.615 1.915 77.785 4.870 ;
        RECT 79.095 1.915 79.265 4.870 ;
        RECT 80.575 1.915 80.745 4.870 ;
        RECT 81.685 4.540 81.875 4.870 ;
        RECT 81.685 1.915 81.855 4.540 ;
        RECT 70.415 0.910 71.635 1.080 ;
        RECT 70.415 0.830 70.585 0.910 ;
        RECT 70.895 0.625 71.065 0.705 ;
        RECT 69.925 0.455 71.065 0.625 ;
        RECT 69.925 0.375 70.095 0.455 ;
        RECT 70.895 0.375 71.065 0.455 ;
        RECT 71.465 0.625 71.635 0.910 ;
        RECT 71.950 1.580 72.605 1.750 ;
        RECT 73.870 1.665 74.040 1.745 ;
        RECT 74.840 1.665 75.010 1.745 ;
        RECT 71.950 0.845 72.120 1.580 ;
        RECT 73.870 1.495 75.010 1.665 ;
        RECT 72.435 0.625 72.605 1.395 ;
        RECT 71.465 0.455 72.605 0.625 ;
        RECT 71.465 0.375 71.635 0.455 ;
        RECT 72.435 0.375 72.605 0.455 ;
        RECT 73.870 0.365 74.040 1.495 ;
        RECT 74.840 0.615 75.010 1.495 ;
        RECT 75.325 1.170 75.495 1.345 ;
        RECT 75.320 1.015 75.495 1.170 ;
        RECT 75.320 0.835 75.490 1.015 ;
        RECT 75.810 0.615 75.980 1.745 ;
        RECT 74.840 0.445 75.980 0.615 ;
        RECT 74.840 0.365 75.010 0.445 ;
        RECT 75.810 0.365 75.980 0.445 ;
        RECT 77.200 1.665 77.370 1.745 ;
        RECT 78.170 1.665 78.340 1.745 ;
        RECT 77.200 1.495 78.340 1.665 ;
        RECT 77.200 0.365 77.370 1.495 ;
        RECT 78.170 0.615 78.340 1.495 ;
        RECT 78.655 0.835 78.825 1.345 ;
        RECT 79.140 0.615 79.310 1.745 ;
        RECT 78.170 0.445 79.310 0.615 ;
        RECT 78.170 0.365 78.340 0.445 ;
        RECT 79.140 0.365 79.310 0.445 ;
        RECT 80.530 1.665 80.700 1.745 ;
        RECT 81.500 1.665 81.670 1.745 ;
        RECT 82.425 1.730 82.595 5.125 ;
        RECT 83.905 1.920 84.075 4.865 ;
        RECT 84.280 4.665 84.450 7.020 ;
        RECT 84.280 4.495 84.815 4.665 ;
        RECT 84.645 2.165 84.815 4.495 ;
        RECT 84.275 1.995 84.815 2.165 ;
        RECT 80.530 1.495 81.670 1.665 ;
        RECT 80.530 0.365 80.700 1.495 ;
        RECT 81.500 0.615 81.670 1.495 ;
        RECT 81.985 1.560 82.595 1.730 ;
        RECT 81.985 0.835 82.155 1.560 ;
        RECT 82.470 0.615 82.640 1.390 ;
        RECT 84.275 0.840 84.445 1.995 ;
        RECT 81.500 0.445 82.640 0.615 ;
        RECT 81.500 0.365 81.670 0.445 ;
        RECT 82.470 0.365 82.640 0.445 ;
      LAYER mcon ;
        RECT 1.765 3.985 1.935 4.155 ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.500 4.525 2.670 ;
        RECT 7.310 3.985 7.480 4.155 ;
        RECT 6.575 3.615 6.745 3.785 ;
        RECT 9.165 2.505 9.335 2.675 ;
        RECT 11.385 3.615 11.555 3.785 ;
        RECT 12.125 2.505 12.295 2.675 ;
        RECT 13.975 2.505 14.145 2.675 ;
        RECT 15.455 3.615 15.625 3.785 ;
        RECT 17.305 3.985 17.475 4.155 ;
        RECT 18.045 3.245 18.215 3.415 ;
        RECT 18.785 3.985 18.955 4.155 ;
        RECT 20.635 3.985 20.805 4.155 ;
        RECT 22.855 3.615 23.025 3.785 ;
        RECT 23.595 3.245 23.765 3.415 ;
        RECT 26.185 3.985 26.355 4.155 ;
        RECT 26.925 2.505 27.095 2.675 ;
        RECT 28.775 2.500 28.945 2.670 ;
        RECT 31.730 3.985 31.900 4.155 ;
        RECT 30.995 3.615 31.165 3.785 ;
        RECT 33.585 2.505 33.755 2.675 ;
        RECT 35.805 3.615 35.975 3.785 ;
        RECT 36.545 2.505 36.715 2.675 ;
        RECT 38.395 2.505 38.565 2.675 ;
        RECT 39.875 3.615 40.045 3.785 ;
        RECT 41.725 3.985 41.895 4.155 ;
        RECT 42.465 3.985 42.635 4.155 ;
        RECT 43.205 2.505 43.375 2.675 ;
        RECT 45.055 2.505 45.225 2.675 ;
        RECT 47.275 3.615 47.445 3.785 ;
        RECT 48.015 3.985 48.185 4.155 ;
        RECT 48.015 2.505 48.185 2.675 ;
        RECT 50.605 3.985 50.775 4.155 ;
        RECT 51.345 2.505 51.515 2.675 ;
        RECT 53.195 2.500 53.365 2.670 ;
        RECT 56.150 3.985 56.320 4.155 ;
        RECT 55.415 3.615 55.585 3.785 ;
        RECT 58.005 2.505 58.175 2.675 ;
        RECT 60.225 3.615 60.395 3.785 ;
        RECT 60.965 2.505 61.135 2.675 ;
        RECT 62.815 2.505 62.985 2.675 ;
        RECT 75.285 5.125 75.455 5.295 ;
        RECT 64.295 3.615 64.465 3.785 ;
        RECT 66.145 3.985 66.315 4.155 ;
        RECT 67.625 4.725 67.795 4.895 ;
        RECT 66.885 4.355 67.055 4.525 ;
        RECT 69.475 4.725 69.645 4.895 ;
        RECT 71.695 3.615 71.865 3.785 ;
        RECT 77.285 5.125 77.455 5.295 ;
        RECT 78.605 5.125 78.775 5.295 ;
        RECT 80.625 5.125 80.795 5.295 ;
        RECT 72.435 4.355 72.605 4.525 ;
        RECT 73.915 4.355 74.085 4.525 ;
        RECT 75.025 3.985 75.195 4.155 ;
        RECT 75.025 2.875 75.195 3.045 ;
        RECT 77.615 4.355 77.785 4.525 ;
        RECT 79.095 3.245 79.265 3.415 ;
        RECT 79.095 1.995 79.265 2.165 ;
        RECT 80.575 1.995 80.745 2.165 ;
        RECT 81.685 3.985 81.855 4.155 ;
        RECT 82.425 3.985 82.595 4.155 ;
        RECT 75.325 1.095 75.495 1.265 ;
        RECT 78.655 1.095 78.825 1.265 ;
        RECT 83.905 3.985 84.075 4.155 ;
        RECT 81.985 1.095 82.155 1.265 ;
      LAYER met1 ;
        RECT 75.255 5.295 75.485 5.325 ;
        RECT 77.255 5.295 77.485 5.325 ;
        RECT 78.575 5.295 78.805 5.325 ;
        RECT 80.595 5.295 80.825 5.325 ;
        RECT 75.225 5.125 77.515 5.295 ;
        RECT 78.545 5.125 80.855 5.295 ;
        RECT 75.255 5.095 75.485 5.125 ;
        RECT 77.255 5.095 77.485 5.125 ;
        RECT 78.575 5.095 78.805 5.125 ;
        RECT 80.595 5.095 80.825 5.125 ;
        RECT 67.595 4.895 67.825 4.925 ;
        RECT 69.445 4.895 69.675 4.925 ;
        RECT 67.565 4.725 69.705 4.895 ;
        RECT 67.595 4.695 67.825 4.725 ;
        RECT 69.445 4.695 69.675 4.725 ;
        RECT 66.855 4.525 67.085 4.555 ;
        RECT 72.405 4.525 72.635 4.555 ;
        RECT 73.885 4.525 74.115 4.555 ;
        RECT 77.585 4.525 77.815 4.555 ;
        RECT 66.825 4.355 77.845 4.525 ;
        RECT 66.855 4.325 67.085 4.355 ;
        RECT 72.405 4.325 72.635 4.355 ;
        RECT 73.885 4.325 74.115 4.355 ;
        RECT 77.585 4.325 77.815 4.355 ;
        RECT 1.735 4.155 1.965 4.185 ;
        RECT 7.280 4.155 7.510 4.185 ;
        RECT 17.275 4.155 17.505 4.185 ;
        RECT 18.755 4.155 18.985 4.185 ;
        RECT 20.605 4.155 20.835 4.185 ;
        RECT 26.155 4.155 26.385 4.185 ;
        RECT 31.700 4.155 31.930 4.185 ;
        RECT 41.695 4.155 41.925 4.185 ;
        RECT 42.435 4.155 42.665 4.185 ;
        RECT 47.985 4.155 48.215 4.185 ;
        RECT 50.575 4.155 50.805 4.185 ;
        RECT 56.120 4.155 56.350 4.185 ;
        RECT 66.115 4.155 66.345 4.185 ;
        RECT 74.995 4.155 75.225 4.185 ;
        RECT 81.655 4.155 81.885 4.185 ;
        RECT 82.395 4.155 82.625 4.185 ;
        RECT 83.875 4.155 84.105 4.185 ;
        RECT 1.705 3.985 17.535 4.155 ;
        RECT 18.725 3.985 20.865 4.155 ;
        RECT 26.125 3.985 41.955 4.155 ;
        RECT 42.405 3.985 48.245 4.155 ;
        RECT 50.545 3.985 66.375 4.155 ;
        RECT 74.965 3.985 81.915 4.155 ;
        RECT 82.365 3.985 84.135 4.155 ;
        RECT 1.735 3.955 1.965 3.985 ;
        RECT 7.280 3.955 7.510 3.985 ;
        RECT 17.275 3.955 17.505 3.985 ;
        RECT 18.755 3.955 18.985 3.985 ;
        RECT 20.605 3.955 20.835 3.985 ;
        RECT 26.155 3.955 26.385 3.985 ;
        RECT 31.700 3.955 31.930 3.985 ;
        RECT 41.695 3.955 41.925 3.985 ;
        RECT 42.435 3.955 42.665 3.985 ;
        RECT 47.985 3.955 48.215 3.985 ;
        RECT 50.575 3.955 50.805 3.985 ;
        RECT 56.120 3.955 56.350 3.985 ;
        RECT 66.115 3.955 66.345 3.985 ;
        RECT 74.995 3.955 75.225 3.985 ;
        RECT 81.655 3.955 81.885 3.985 ;
        RECT 82.395 3.955 82.625 3.985 ;
        RECT 83.875 3.955 84.105 3.985 ;
        RECT 6.545 3.785 6.775 3.815 ;
        RECT 11.355 3.785 11.585 3.815 ;
        RECT 15.425 3.785 15.655 3.815 ;
        RECT 22.825 3.785 23.055 3.815 ;
        RECT 30.965 3.785 31.195 3.815 ;
        RECT 35.775 3.785 36.005 3.815 ;
        RECT 39.845 3.785 40.075 3.815 ;
        RECT 47.245 3.785 47.475 3.815 ;
        RECT 55.385 3.785 55.615 3.815 ;
        RECT 60.195 3.785 60.425 3.815 ;
        RECT 64.265 3.785 64.495 3.815 ;
        RECT 71.665 3.785 71.895 3.815 ;
        RECT 6.515 3.615 23.085 3.785 ;
        RECT 30.935 3.615 47.505 3.785 ;
        RECT 55.355 3.615 71.925 3.785 ;
        RECT 6.545 3.585 6.775 3.615 ;
        RECT 11.355 3.585 11.585 3.615 ;
        RECT 15.425 3.585 15.655 3.615 ;
        RECT 22.825 3.585 23.055 3.615 ;
        RECT 30.965 3.585 31.195 3.615 ;
        RECT 35.775 3.585 36.005 3.615 ;
        RECT 39.845 3.585 40.075 3.615 ;
        RECT 47.245 3.585 47.475 3.615 ;
        RECT 55.385 3.585 55.615 3.615 ;
        RECT 60.195 3.585 60.425 3.615 ;
        RECT 64.265 3.585 64.495 3.615 ;
        RECT 71.665 3.585 71.895 3.615 ;
        RECT 18.015 3.415 18.245 3.445 ;
        RECT 23.565 3.415 23.795 3.445 ;
        RECT 79.065 3.415 79.295 3.445 ;
        RECT 17.985 3.245 79.325 3.415 ;
        RECT 18.015 3.215 18.245 3.245 ;
        RECT 23.565 3.215 23.795 3.245 ;
        RECT 79.065 3.215 79.295 3.245 ;
        RECT 74.995 3.045 75.225 3.075 ;
        RECT 50.605 2.875 75.255 3.045 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.700 ;
        RECT 9.135 2.675 9.365 2.705 ;
        RECT 12.095 2.675 12.325 2.705 ;
        RECT 13.945 2.675 14.175 2.705 ;
        RECT 26.895 2.675 27.125 2.705 ;
        RECT 28.745 2.675 28.975 2.700 ;
        RECT 33.555 2.675 33.785 2.705 ;
        RECT 36.515 2.675 36.745 2.705 ;
        RECT 38.365 2.675 38.595 2.705 ;
        RECT 43.175 2.675 43.405 2.705 ;
        RECT 45.025 2.675 45.255 2.705 ;
        RECT 47.985 2.675 48.215 2.705 ;
        RECT 50.605 2.675 50.775 2.875 ;
        RECT 74.995 2.845 75.225 2.875 ;
        RECT 51.315 2.675 51.545 2.705 ;
        RECT 53.165 2.675 53.395 2.700 ;
        RECT 57.975 2.675 58.205 2.705 ;
        RECT 60.935 2.675 61.165 2.705 ;
        RECT 62.785 2.675 63.015 2.705 ;
        RECT 2.445 2.505 9.395 2.675 ;
        RECT 12.065 2.505 14.205 2.675 ;
        RECT 26.865 2.505 33.815 2.675 ;
        RECT 36.485 2.505 38.625 2.675 ;
        RECT 43.145 2.505 45.285 2.675 ;
        RECT 47.955 2.505 50.775 2.675 ;
        RECT 51.285 2.505 58.235 2.675 ;
        RECT 60.905 2.505 63.045 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.295 2.500 4.705 2.505 ;
        RECT 4.325 2.470 4.555 2.500 ;
        RECT 9.135 2.475 9.365 2.505 ;
        RECT 12.095 2.475 12.325 2.505 ;
        RECT 13.945 2.475 14.175 2.505 ;
        RECT 26.895 2.475 27.125 2.505 ;
        RECT 28.715 2.500 29.125 2.505 ;
        RECT 28.745 2.470 28.975 2.500 ;
        RECT 33.555 2.475 33.785 2.505 ;
        RECT 36.515 2.475 36.745 2.505 ;
        RECT 38.365 2.475 38.595 2.505 ;
        RECT 43.175 2.475 43.405 2.505 ;
        RECT 45.025 2.475 45.255 2.505 ;
        RECT 47.985 2.475 48.215 2.505 ;
        RECT 51.315 2.475 51.545 2.505 ;
        RECT 53.135 2.500 53.545 2.505 ;
        RECT 53.165 2.470 53.395 2.500 ;
        RECT 57.975 2.475 58.205 2.505 ;
        RECT 60.935 2.475 61.165 2.505 ;
        RECT 62.785 2.475 63.015 2.505 ;
        RECT 79.065 2.165 79.295 2.195 ;
        RECT 80.545 2.165 80.775 2.195 ;
        RECT 79.035 1.995 80.805 2.165 ;
        RECT 79.065 1.965 79.295 1.995 ;
        RECT 80.545 1.965 80.775 1.995 ;
        RECT 75.295 1.265 75.525 1.295 ;
        RECT 78.625 1.265 78.855 1.295 ;
        RECT 81.955 1.265 82.185 1.295 ;
        RECT 75.265 1.095 82.215 1.265 ;
        RECT 75.295 1.065 75.525 1.095 ;
        RECT 78.625 1.065 78.855 1.095 ;
        RECT 81.955 1.065 82.185 1.095 ;
  END
END TMRDFFSNQX1






MACRO TMRDFFSNRNQNX1
  CLASS CORE ;
  FOREIGN TMRDFFSNRNQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 96.570 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN SN
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 11.755 1.915 11.925 4.865 ;
        RECT 26.185 1.915 26.355 4.865 ;
        RECT 40.615 1.915 40.785 4.865 ;
        RECT 55.045 1.915 55.215 4.865 ;
        RECT 69.475 1.915 69.645 4.865 ;
        RECT 83.905 1.915 84.075 4.865 ;
      LAYER mcon ;
        RECT 11.755 2.875 11.925 3.045 ;
        RECT 26.185 2.875 26.355 3.045 ;
        RECT 40.615 2.875 40.785 3.045 ;
        RECT 55.045 2.875 55.215 3.045 ;
        RECT 69.475 2.875 69.645 3.045 ;
        RECT 83.905 2.875 84.075 3.045 ;
      LAYER met1 ;
        RECT 11.725 3.045 11.955 3.075 ;
        RECT 26.155 3.045 26.385 3.075 ;
        RECT 40.585 3.045 40.815 3.075 ;
        RECT 55.015 3.045 55.245 3.075 ;
        RECT 69.445 3.045 69.675 3.075 ;
        RECT 83.875 3.045 84.105 3.075 ;
        RECT 11.695 2.875 84.135 3.045 ;
        RECT 11.725 2.845 11.955 2.875 ;
        RECT 26.155 2.845 26.385 2.875 ;
        RECT 40.585 2.845 40.815 2.875 ;
        RECT 55.015 2.845 55.245 2.875 ;
        RECT 69.445 2.845 69.675 2.875 ;
        RECT 83.875 2.845 84.105 2.875 ;
    END
  END SN
  PIN RN
    ANTENNAGATEAREA 9.170850 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 17.675 1.915 17.845 4.865 ;
        RECT 21.375 1.915 21.545 4.865 ;
        RECT 30.995 1.915 31.165 4.865 ;
        RECT 46.535 1.915 46.705 4.865 ;
        RECT 50.235 1.915 50.405 4.865 ;
        RECT 59.855 1.915 60.025 4.865 ;
        RECT 75.395 1.915 75.565 4.865 ;
        RECT 79.095 1.915 79.265 4.865 ;
      LAYER mcon ;
        RECT 2.135 2.135 2.305 2.305 ;
        RECT 17.675 2.135 17.845 2.305 ;
        RECT 21.375 2.135 21.545 2.305 ;
        RECT 30.995 2.135 31.165 2.305 ;
        RECT 46.535 2.135 46.705 2.305 ;
        RECT 50.235 2.135 50.405 2.305 ;
        RECT 59.855 2.135 60.025 2.305 ;
        RECT 75.395 2.135 75.565 2.305 ;
        RECT 79.095 2.135 79.265 2.305 ;
      LAYER met1 ;
        RECT 2.105 2.305 2.335 2.335 ;
        RECT 17.645 2.305 17.875 2.335 ;
        RECT 21.345 2.305 21.575 2.335 ;
        RECT 30.965 2.305 31.195 2.335 ;
        RECT 46.505 2.305 46.735 2.335 ;
        RECT 50.205 2.305 50.435 2.335 ;
        RECT 59.825 2.305 60.055 2.335 ;
        RECT 75.365 2.305 75.595 2.335 ;
        RECT 79.065 2.305 79.295 2.335 ;
        RECT 2.075 2.135 79.325 2.305 ;
        RECT 2.105 2.105 2.335 2.135 ;
        RECT 17.645 2.105 17.875 2.135 ;
        RECT 21.345 2.105 21.575 2.135 ;
        RECT 30.965 2.105 31.195 2.135 ;
        RECT 46.505 2.105 46.735 2.135 ;
        RECT 50.205 2.105 50.435 2.135 ;
        RECT 59.825 2.105 60.055 2.135 ;
        RECT 75.365 2.105 75.595 2.135 ;
        RECT 79.065 2.105 79.295 2.135 ;
    END
  END RN
  PIN D
    ANTENNAGATEAREA 3.099750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 29.885 1.915 30.055 4.865 ;
        RECT 58.745 1.915 58.915 4.865 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 29.885 3.985 30.055 4.155 ;
        RECT 58.745 3.985 58.915 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 29.855 4.155 30.085 4.185 ;
        RECT 58.715 4.155 58.945 4.185 ;
        RECT 0.845 3.985 58.975 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 29.855 3.955 30.085 3.985 ;
        RECT 58.715 3.955 58.945 3.985 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 16.565 1.915 16.735 4.865 ;
        RECT 35.805 1.915 35.975 4.865 ;
        RECT 45.425 1.915 45.595 4.865 ;
        RECT 64.665 1.915 64.835 4.865 ;
        RECT 74.285 1.915 74.455 4.865 ;
      LAYER mcon ;
        RECT 6.945 4.355 7.115 4.525 ;
        RECT 16.565 4.355 16.735 4.525 ;
        RECT 35.805 4.355 35.975 4.525 ;
        RECT 45.425 4.355 45.595 4.525 ;
        RECT 64.665 4.355 64.835 4.525 ;
        RECT 74.285 4.355 74.455 4.525 ;
      LAYER met1 ;
        RECT 6.915 4.525 7.145 4.555 ;
        RECT 16.535 4.525 16.765 4.555 ;
        RECT 35.775 4.525 36.005 4.555 ;
        RECT 45.395 4.525 45.625 4.555 ;
        RECT 64.635 4.525 64.865 4.555 ;
        RECT 74.255 4.525 74.485 4.555 ;
        RECT 6.885 4.355 74.515 4.525 ;
        RECT 6.915 4.325 7.145 4.355 ;
        RECT 16.535 4.325 16.765 4.355 ;
        RECT 35.775 4.325 36.005 4.355 ;
        RECT 45.395 4.325 45.625 4.355 ;
        RECT 64.635 4.325 64.865 4.355 ;
        RECT 74.255 4.325 74.485 4.355 ;
    END
  END CLK
  PIN Q
    ANTENNADIFFAREA 1.734950 ;
    PORT
      LAYER li1 ;
        RECT 94.385 5.295 94.555 6.565 ;
        RECT 95.265 5.295 95.435 6.565 ;
        RECT 94.385 5.125 95.915 5.295 ;
        RECT 95.745 1.730 95.915 5.125 ;
        RECT 95.305 1.560 95.915 1.730 ;
        RECT 88.645 1.170 88.815 1.345 ;
        RECT 88.640 1.015 88.815 1.170 ;
        RECT 88.640 0.835 88.810 1.015 ;
        RECT 91.975 0.835 92.145 1.345 ;
        RECT 95.305 0.835 95.475 1.560 ;
      LAYER mcon ;
        RECT 95.745 3.985 95.915 4.155 ;
        RECT 88.645 1.095 88.815 1.265 ;
        RECT 91.975 1.095 92.145 1.265 ;
        RECT 95.305 1.095 95.475 1.265 ;
      LAYER met1 ;
        RECT 95.715 4.155 95.945 4.185 ;
        RECT 95.685 3.985 96.095 4.155 ;
        RECT 95.715 3.955 95.945 3.985 ;
        RECT 88.615 1.265 88.845 1.295 ;
        RECT 91.945 1.265 92.175 1.295 ;
        RECT 95.275 1.265 95.505 1.295 ;
        RECT 88.585 1.095 95.535 1.265 ;
        RECT 88.615 1.065 88.845 1.095 ;
        RECT 91.945 1.065 92.175 1.095 ;
        RECT 95.275 1.065 95.505 1.095 ;
    END
  END Q
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 97.005 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 96.740 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.625 5.215 10.795 7.230 ;
        RECT 11.505 5.555 11.675 7.230 ;
        RECT 12.385 5.555 12.555 7.230 ;
        RECT 13.265 5.555 13.435 7.230 ;
        RECT 14.260 4.110 14.600 7.230 ;
        RECT 15.435 5.215 15.605 7.230 ;
        RECT 16.315 5.555 16.485 7.230 ;
        RECT 17.195 5.555 17.365 7.230 ;
        RECT 18.075 5.555 18.245 7.230 ;
        RECT 19.070 4.110 19.410 7.230 ;
        RECT 20.245 5.215 20.415 7.230 ;
        RECT 21.125 5.555 21.295 7.230 ;
        RECT 22.005 5.555 22.175 7.230 ;
        RECT 22.885 5.555 23.055 7.230 ;
        RECT 23.880 4.110 24.220 7.230 ;
        RECT 25.055 5.215 25.225 7.230 ;
        RECT 25.935 5.555 26.105 7.230 ;
        RECT 26.815 5.555 26.985 7.230 ;
        RECT 27.695 5.555 27.865 7.230 ;
        RECT 28.690 4.110 29.030 7.230 ;
        RECT 29.865 5.215 30.035 7.230 ;
        RECT 30.745 5.555 30.915 7.230 ;
        RECT 31.625 5.555 31.795 7.230 ;
        RECT 32.505 5.555 32.675 7.230 ;
        RECT 33.500 4.110 33.840 7.230 ;
        RECT 34.675 5.215 34.845 7.230 ;
        RECT 35.555 5.555 35.725 7.230 ;
        RECT 36.435 5.555 36.605 7.230 ;
        RECT 37.315 5.555 37.485 7.230 ;
        RECT 38.310 4.110 38.650 7.230 ;
        RECT 39.485 5.215 39.655 7.230 ;
        RECT 40.365 5.555 40.535 7.230 ;
        RECT 41.245 5.555 41.415 7.230 ;
        RECT 42.125 5.555 42.295 7.230 ;
        RECT 43.120 4.110 43.460 7.230 ;
        RECT 44.295 5.215 44.465 7.230 ;
        RECT 45.175 5.555 45.345 7.230 ;
        RECT 46.055 5.555 46.225 7.230 ;
        RECT 46.935 5.555 47.105 7.230 ;
        RECT 47.930 4.110 48.270 7.230 ;
        RECT 49.105 5.215 49.275 7.230 ;
        RECT 49.985 5.555 50.155 7.230 ;
        RECT 50.865 5.555 51.035 7.230 ;
        RECT 51.745 5.555 51.915 7.230 ;
        RECT 52.740 4.110 53.080 7.230 ;
        RECT 53.915 5.215 54.085 7.230 ;
        RECT 54.795 5.555 54.965 7.230 ;
        RECT 55.675 5.555 55.845 7.230 ;
        RECT 56.555 5.555 56.725 7.230 ;
        RECT 57.550 4.110 57.890 7.230 ;
        RECT 58.725 5.215 58.895 7.230 ;
        RECT 59.605 5.555 59.775 7.230 ;
        RECT 60.485 5.555 60.655 7.230 ;
        RECT 61.365 5.555 61.535 7.230 ;
        RECT 62.360 4.110 62.700 7.230 ;
        RECT 63.535 5.215 63.705 7.230 ;
        RECT 64.415 5.555 64.585 7.230 ;
        RECT 65.295 5.555 65.465 7.230 ;
        RECT 66.175 5.555 66.345 7.230 ;
        RECT 67.170 4.110 67.510 7.230 ;
        RECT 68.345 5.215 68.515 7.230 ;
        RECT 69.225 5.555 69.395 7.230 ;
        RECT 70.105 5.555 70.275 7.230 ;
        RECT 70.985 5.555 71.155 7.230 ;
        RECT 71.980 4.110 72.320 7.230 ;
        RECT 73.155 5.215 73.325 7.230 ;
        RECT 74.035 5.555 74.205 7.230 ;
        RECT 74.915 5.555 75.085 7.230 ;
        RECT 75.795 5.555 75.965 7.230 ;
        RECT 76.790 4.110 77.130 7.230 ;
        RECT 77.965 5.215 78.135 7.230 ;
        RECT 78.845 5.555 79.015 7.230 ;
        RECT 79.725 5.555 79.895 7.230 ;
        RECT 80.605 5.555 80.775 7.230 ;
        RECT 81.600 4.110 81.940 7.230 ;
        RECT 82.775 5.215 82.945 7.230 ;
        RECT 83.655 5.555 83.825 7.230 ;
        RECT 84.535 5.555 84.705 7.230 ;
        RECT 85.415 5.555 85.585 7.230 ;
        RECT 86.410 4.110 86.750 7.230 ;
        RECT 87.285 5.125 87.455 7.230 ;
        RECT 88.165 5.555 88.335 7.230 ;
        RECT 89.045 5.125 89.215 7.230 ;
        RECT 89.740 4.110 90.080 7.230 ;
        RECT 93.070 4.110 93.410 7.230 ;
        RECT 96.400 4.110 96.740 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.515 7.315 29.685 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.625 7.315 30.795 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 32.845 7.315 33.015 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.435 7.315 35.605 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.175 7.315 36.345 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.765 7.315 38.935 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.505 7.315 39.675 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.615 7.315 40.785 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 42.835 7.315 43.005 7.485 ;
        RECT 43.575 7.315 43.745 7.485 ;
        RECT 43.945 7.315 44.115 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 47.645 7.315 47.815 7.485 ;
        RECT 48.385 7.315 48.555 7.485 ;
        RECT 48.755 7.315 48.925 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 50.975 7.315 51.145 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 51.715 7.315 51.885 7.485 ;
        RECT 52.085 7.315 52.255 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.305 7.315 54.475 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.525 7.315 56.695 7.485 ;
        RECT 56.895 7.315 57.065 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 60.965 7.315 61.135 7.485 ;
        RECT 61.335 7.315 61.505 7.485 ;
        RECT 61.705 7.315 61.875 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.295 7.315 64.465 7.485 ;
        RECT 64.665 7.315 64.835 7.485 ;
        RECT 65.035 7.315 65.205 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.625 7.315 67.795 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.365 7.315 68.535 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.475 7.315 69.645 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 70.955 7.315 71.125 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.175 7.315 73.345 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
        RECT 74.285 7.315 74.455 7.485 ;
        RECT 74.655 7.315 74.825 7.485 ;
        RECT 75.025 7.315 75.195 7.485 ;
        RECT 75.395 7.315 75.565 7.485 ;
        RECT 75.765 7.315 75.935 7.485 ;
        RECT 76.135 7.315 76.305 7.485 ;
        RECT 76.505 7.315 76.675 7.485 ;
        RECT 77.245 7.315 77.415 7.485 ;
        RECT 77.615 7.315 77.785 7.485 ;
        RECT 77.985 7.315 78.155 7.485 ;
        RECT 78.355 7.315 78.525 7.485 ;
        RECT 78.725 7.315 78.895 7.485 ;
        RECT 79.095 7.315 79.265 7.485 ;
        RECT 79.465 7.315 79.635 7.485 ;
        RECT 79.835 7.315 80.005 7.485 ;
        RECT 80.205 7.315 80.375 7.485 ;
        RECT 80.575 7.315 80.745 7.485 ;
        RECT 80.945 7.315 81.115 7.485 ;
        RECT 81.315 7.315 81.485 7.485 ;
        RECT 82.055 7.315 82.225 7.485 ;
        RECT 82.425 7.315 82.595 7.485 ;
        RECT 82.795 7.315 82.965 7.485 ;
        RECT 83.165 7.315 83.335 7.485 ;
        RECT 83.535 7.315 83.705 7.485 ;
        RECT 83.905 7.315 84.075 7.485 ;
        RECT 84.275 7.315 84.445 7.485 ;
        RECT 84.645 7.315 84.815 7.485 ;
        RECT 85.015 7.315 85.185 7.485 ;
        RECT 85.385 7.315 85.555 7.485 ;
        RECT 85.755 7.315 85.925 7.485 ;
        RECT 86.125 7.315 86.295 7.485 ;
        RECT 86.865 7.315 87.035 7.485 ;
        RECT 87.235 7.315 87.405 7.485 ;
        RECT 87.605 7.315 87.775 7.485 ;
        RECT 87.975 7.315 88.145 7.485 ;
        RECT 88.345 7.315 88.515 7.485 ;
        RECT 88.715 7.315 88.885 7.485 ;
        RECT 89.085 7.315 89.255 7.485 ;
        RECT 89.455 7.315 89.625 7.485 ;
        RECT 90.195 7.315 90.365 7.485 ;
        RECT 90.565 7.315 90.735 7.485 ;
        RECT 90.935 7.315 91.105 7.485 ;
        RECT 91.305 7.315 91.475 7.485 ;
        RECT 91.675 7.315 91.845 7.485 ;
        RECT 92.045 7.315 92.215 7.485 ;
        RECT 92.415 7.315 92.585 7.485 ;
        RECT 92.785 7.315 92.955 7.485 ;
        RECT 93.525 7.315 93.695 7.485 ;
        RECT 93.895 7.315 94.065 7.485 ;
        RECT 94.265 7.315 94.435 7.485 ;
        RECT 94.635 7.315 94.805 7.485 ;
        RECT 95.005 7.315 95.175 7.485 ;
        RECT 95.375 7.315 95.545 7.485 ;
        RECT 95.745 7.315 95.915 7.485 ;
        RECT 96.115 7.315 96.285 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 96.740 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 96.740 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.610 0.170 10.780 1.130 ;
        RECT 14.260 0.170 14.600 2.720 ;
        RECT 15.420 0.170 15.590 1.130 ;
        RECT 19.070 0.170 19.410 2.720 ;
        RECT 20.230 0.170 20.400 1.130 ;
        RECT 23.880 0.170 24.220 2.720 ;
        RECT 25.040 0.170 25.210 1.130 ;
        RECT 28.690 0.170 29.030 2.720 ;
        RECT 29.850 0.170 30.020 1.130 ;
        RECT 33.500 0.170 33.840 2.720 ;
        RECT 34.660 0.170 34.830 1.130 ;
        RECT 38.310 0.170 38.650 2.720 ;
        RECT 39.470 0.170 39.640 1.130 ;
        RECT 43.120 0.170 43.460 2.720 ;
        RECT 44.280 0.170 44.450 1.130 ;
        RECT 47.930 0.170 48.270 2.720 ;
        RECT 49.090 0.170 49.260 1.130 ;
        RECT 52.740 0.170 53.080 2.720 ;
        RECT 53.900 0.170 54.070 1.130 ;
        RECT 57.550 0.170 57.890 2.720 ;
        RECT 58.710 0.170 58.880 1.130 ;
        RECT 62.360 0.170 62.700 2.720 ;
        RECT 63.520 0.170 63.690 1.130 ;
        RECT 67.170 0.170 67.510 2.720 ;
        RECT 68.330 0.170 68.500 1.130 ;
        RECT 71.980 0.170 72.320 2.720 ;
        RECT 73.140 0.170 73.310 1.130 ;
        RECT 76.790 0.170 77.130 2.720 ;
        RECT 77.950 0.170 78.120 1.130 ;
        RECT 81.600 0.170 81.940 2.720 ;
        RECT 82.760 0.170 82.930 1.130 ;
        RECT 86.410 0.170 86.750 2.720 ;
        RECT 87.675 0.170 87.845 1.120 ;
        RECT 89.740 0.170 90.080 2.720 ;
        RECT 91.005 0.170 91.175 1.120 ;
        RECT 93.070 0.170 93.410 2.720 ;
        RECT 94.335 0.170 94.505 1.120 ;
        RECT 96.400 0.170 96.740 2.720 ;
        RECT -0.170 -0.170 96.740 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.515 -0.085 29.685 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.625 -0.085 30.795 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 32.845 -0.085 33.015 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.435 -0.085 35.605 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.175 -0.085 36.345 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.765 -0.085 38.935 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.505 -0.085 39.675 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.615 -0.085 40.785 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 42.835 -0.085 43.005 0.085 ;
        RECT 43.575 -0.085 43.745 0.085 ;
        RECT 43.945 -0.085 44.115 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 47.645 -0.085 47.815 0.085 ;
        RECT 48.385 -0.085 48.555 0.085 ;
        RECT 48.755 -0.085 48.925 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 50.975 -0.085 51.145 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 51.715 -0.085 51.885 0.085 ;
        RECT 52.085 -0.085 52.255 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.305 -0.085 54.475 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.525 -0.085 56.695 0.085 ;
        RECT 56.895 -0.085 57.065 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 60.965 -0.085 61.135 0.085 ;
        RECT 61.335 -0.085 61.505 0.085 ;
        RECT 61.705 -0.085 61.875 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.295 -0.085 64.465 0.085 ;
        RECT 64.665 -0.085 64.835 0.085 ;
        RECT 65.035 -0.085 65.205 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.625 -0.085 67.795 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.365 -0.085 68.535 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.475 -0.085 69.645 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 70.955 -0.085 71.125 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.175 -0.085 73.345 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
        RECT 74.285 -0.085 74.455 0.085 ;
        RECT 74.655 -0.085 74.825 0.085 ;
        RECT 75.025 -0.085 75.195 0.085 ;
        RECT 75.395 -0.085 75.565 0.085 ;
        RECT 75.765 -0.085 75.935 0.085 ;
        RECT 76.135 -0.085 76.305 0.085 ;
        RECT 76.505 -0.085 76.675 0.085 ;
        RECT 77.245 -0.085 77.415 0.085 ;
        RECT 77.615 -0.085 77.785 0.085 ;
        RECT 77.985 -0.085 78.155 0.085 ;
        RECT 78.355 -0.085 78.525 0.085 ;
        RECT 78.725 -0.085 78.895 0.085 ;
        RECT 79.095 -0.085 79.265 0.085 ;
        RECT 79.465 -0.085 79.635 0.085 ;
        RECT 79.835 -0.085 80.005 0.085 ;
        RECT 80.205 -0.085 80.375 0.085 ;
        RECT 80.575 -0.085 80.745 0.085 ;
        RECT 80.945 -0.085 81.115 0.085 ;
        RECT 81.315 -0.085 81.485 0.085 ;
        RECT 82.055 -0.085 82.225 0.085 ;
        RECT 82.425 -0.085 82.595 0.085 ;
        RECT 82.795 -0.085 82.965 0.085 ;
        RECT 83.165 -0.085 83.335 0.085 ;
        RECT 83.535 -0.085 83.705 0.085 ;
        RECT 83.905 -0.085 84.075 0.085 ;
        RECT 84.275 -0.085 84.445 0.085 ;
        RECT 84.645 -0.085 84.815 0.085 ;
        RECT 85.015 -0.085 85.185 0.085 ;
        RECT 85.385 -0.085 85.555 0.085 ;
        RECT 85.755 -0.085 85.925 0.085 ;
        RECT 86.125 -0.085 86.295 0.085 ;
        RECT 86.865 -0.085 87.035 0.085 ;
        RECT 87.235 -0.085 87.405 0.085 ;
        RECT 87.605 -0.085 87.775 0.085 ;
        RECT 87.975 -0.085 88.145 0.085 ;
        RECT 88.345 -0.085 88.515 0.085 ;
        RECT 88.715 -0.085 88.885 0.085 ;
        RECT 89.085 -0.085 89.255 0.085 ;
        RECT 89.455 -0.085 89.625 0.085 ;
        RECT 90.195 -0.085 90.365 0.085 ;
        RECT 90.565 -0.085 90.735 0.085 ;
        RECT 90.935 -0.085 91.105 0.085 ;
        RECT 91.305 -0.085 91.475 0.085 ;
        RECT 91.675 -0.085 91.845 0.085 ;
        RECT 92.045 -0.085 92.215 0.085 ;
        RECT 92.415 -0.085 92.585 0.085 ;
        RECT 92.785 -0.085 92.955 0.085 ;
        RECT 93.525 -0.085 93.695 0.085 ;
        RECT 93.895 -0.085 94.065 0.085 ;
        RECT 94.265 -0.085 94.435 0.085 ;
        RECT 94.635 -0.085 94.805 0.085 ;
        RECT 95.005 -0.085 95.175 0.085 ;
        RECT 95.375 -0.085 95.545 0.085 ;
        RECT 95.745 -0.085 95.915 0.085 ;
        RECT 96.115 -0.085 96.285 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 96.740 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 11.065 5.240 11.235 7.020 ;
        RECT 11.945 5.240 12.115 7.020 ;
        RECT 12.825 5.240 12.995 7.020 ;
        RECT 15.875 5.240 16.045 7.020 ;
        RECT 16.755 5.240 16.925 7.020 ;
        RECT 17.635 5.240 17.805 7.020 ;
        RECT 20.685 5.240 20.855 7.020 ;
        RECT 21.565 5.240 21.735 7.020 ;
        RECT 22.445 5.240 22.615 7.020 ;
        RECT 25.495 5.240 25.665 7.020 ;
        RECT 26.375 5.240 26.545 7.020 ;
        RECT 27.255 5.240 27.425 7.020 ;
        RECT 30.305 5.240 30.475 7.020 ;
        RECT 31.185 5.240 31.355 7.020 ;
        RECT 32.065 5.240 32.235 7.020 ;
        RECT 35.115 5.240 35.285 7.020 ;
        RECT 35.995 5.240 36.165 7.020 ;
        RECT 36.875 5.240 37.045 7.020 ;
        RECT 39.925 5.240 40.095 7.020 ;
        RECT 40.805 5.240 40.975 7.020 ;
        RECT 41.685 5.240 41.855 7.020 ;
        RECT 44.735 5.240 44.905 7.020 ;
        RECT 45.615 5.240 45.785 7.020 ;
        RECT 46.495 5.240 46.665 7.020 ;
        RECT 49.545 5.240 49.715 7.020 ;
        RECT 50.425 5.240 50.595 7.020 ;
        RECT 51.305 5.240 51.475 7.020 ;
        RECT 54.355 5.240 54.525 7.020 ;
        RECT 55.235 5.240 55.405 7.020 ;
        RECT 56.115 5.240 56.285 7.020 ;
        RECT 59.165 5.240 59.335 7.020 ;
        RECT 60.045 5.240 60.215 7.020 ;
        RECT 60.925 5.240 61.095 7.020 ;
        RECT 63.975 5.240 64.145 7.020 ;
        RECT 64.855 5.240 65.025 7.020 ;
        RECT 65.735 5.240 65.905 7.020 ;
        RECT 68.785 5.240 68.955 7.020 ;
        RECT 69.665 5.240 69.835 7.020 ;
        RECT 70.545 5.240 70.715 7.020 ;
        RECT 73.595 5.240 73.765 7.020 ;
        RECT 74.475 5.240 74.645 7.020 ;
        RECT 75.355 5.240 75.525 7.020 ;
        RECT 78.405 5.240 78.575 7.020 ;
        RECT 79.285 5.240 79.455 7.020 ;
        RECT 80.165 5.240 80.335 7.020 ;
        RECT 83.215 5.240 83.385 7.020 ;
        RECT 84.095 5.240 84.265 7.020 ;
        RECT 84.975 5.240 85.145 7.020 ;
        RECT 87.725 6.825 87.905 6.995 ;
        RECT 87.725 5.295 87.895 6.825 ;
        RECT 88.605 5.295 88.775 6.995 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 11.065 5.070 13.775 5.240 ;
        RECT 15.875 5.070 18.585 5.240 ;
        RECT 20.685 5.070 23.395 5.240 ;
        RECT 25.495 5.070 28.205 5.240 ;
        RECT 30.305 5.070 33.015 5.240 ;
        RECT 35.115 5.070 37.825 5.240 ;
        RECT 39.925 5.070 42.635 5.240 ;
        RECT 44.735 5.070 47.445 5.240 ;
        RECT 49.545 5.070 52.255 5.240 ;
        RECT 54.355 5.070 57.065 5.240 ;
        RECT 59.165 5.070 61.875 5.240 ;
        RECT 63.975 5.070 66.685 5.240 ;
        RECT 68.785 5.070 71.495 5.240 ;
        RECT 73.595 5.070 76.305 5.240 ;
        RECT 78.405 5.070 81.115 5.240 ;
        RECT 83.215 5.070 85.925 5.240 ;
        RECT 87.725 5.125 88.775 5.295 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 8.055 1.915 8.225 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 12.865 1.915 13.035 4.865 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.125 1.675 10.295 1.755 ;
        RECT 11.095 1.675 11.265 1.755 ;
        RECT 12.065 1.675 12.235 1.755 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.125 1.505 12.235 1.675 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.125 0.375 10.295 1.505 ;
        RECT 11.095 0.625 11.265 1.505 ;
        RECT 12.065 1.425 12.235 1.505 ;
        RECT 11.585 1.080 11.755 1.160 ;
        RECT 12.635 1.080 12.805 1.755 ;
        RECT 13.605 1.750 13.775 5.070 ;
        RECT 15.455 1.915 15.625 4.865 ;
        RECT 11.585 0.910 12.805 1.080 ;
        RECT 11.585 0.830 11.755 0.910 ;
        RECT 12.065 0.625 12.235 0.705 ;
        RECT 11.095 0.455 12.235 0.625 ;
        RECT 11.095 0.375 11.265 0.455 ;
        RECT 12.065 0.375 12.235 0.455 ;
        RECT 12.635 0.625 12.805 0.910 ;
        RECT 13.120 1.580 13.775 1.750 ;
        RECT 14.935 1.675 15.105 1.755 ;
        RECT 15.905 1.675 16.075 1.755 ;
        RECT 16.875 1.675 17.045 1.755 ;
        RECT 13.120 0.845 13.290 1.580 ;
        RECT 14.935 1.505 17.045 1.675 ;
        RECT 13.605 0.625 13.775 1.395 ;
        RECT 12.635 0.455 13.775 0.625 ;
        RECT 12.635 0.375 12.805 0.455 ;
        RECT 13.605 0.375 13.775 0.455 ;
        RECT 14.935 0.375 15.105 1.505 ;
        RECT 15.905 0.625 16.075 1.505 ;
        RECT 16.875 1.425 17.045 1.505 ;
        RECT 16.395 1.080 16.565 1.160 ;
        RECT 17.445 1.080 17.615 1.755 ;
        RECT 18.415 1.750 18.585 5.070 ;
        RECT 20.265 1.915 20.435 4.865 ;
        RECT 22.485 1.915 22.655 4.865 ;
        RECT 16.395 0.910 17.615 1.080 ;
        RECT 16.395 0.830 16.565 0.910 ;
        RECT 16.875 0.625 17.045 0.705 ;
        RECT 15.905 0.455 17.045 0.625 ;
        RECT 15.905 0.375 16.075 0.455 ;
        RECT 16.875 0.375 17.045 0.455 ;
        RECT 17.445 0.625 17.615 0.910 ;
        RECT 17.930 1.580 18.585 1.750 ;
        RECT 19.745 1.675 19.915 1.755 ;
        RECT 20.715 1.675 20.885 1.755 ;
        RECT 21.685 1.675 21.855 1.755 ;
        RECT 17.930 0.845 18.100 1.580 ;
        RECT 19.745 1.505 21.855 1.675 ;
        RECT 18.415 0.625 18.585 1.395 ;
        RECT 17.445 0.455 18.585 0.625 ;
        RECT 17.445 0.375 17.615 0.455 ;
        RECT 18.415 0.375 18.585 0.455 ;
        RECT 19.745 0.375 19.915 1.505 ;
        RECT 20.715 0.625 20.885 1.505 ;
        RECT 21.685 1.425 21.855 1.505 ;
        RECT 21.205 1.080 21.375 1.160 ;
        RECT 22.255 1.080 22.425 1.755 ;
        RECT 23.225 1.750 23.395 5.070 ;
        RECT 25.075 1.915 25.245 4.865 ;
        RECT 27.295 1.915 27.465 4.865 ;
        RECT 21.205 0.910 22.425 1.080 ;
        RECT 21.205 0.830 21.375 0.910 ;
        RECT 21.685 0.625 21.855 0.705 ;
        RECT 20.715 0.455 21.855 0.625 ;
        RECT 20.715 0.375 20.885 0.455 ;
        RECT 21.685 0.375 21.855 0.455 ;
        RECT 22.255 0.625 22.425 0.910 ;
        RECT 22.740 1.580 23.395 1.750 ;
        RECT 24.555 1.675 24.725 1.755 ;
        RECT 25.525 1.675 25.695 1.755 ;
        RECT 26.495 1.675 26.665 1.755 ;
        RECT 22.740 0.845 22.910 1.580 ;
        RECT 24.555 1.505 26.665 1.675 ;
        RECT 23.225 0.625 23.395 1.395 ;
        RECT 22.255 0.455 23.395 0.625 ;
        RECT 22.255 0.375 22.425 0.455 ;
        RECT 23.225 0.375 23.395 0.455 ;
        RECT 24.555 0.375 24.725 1.505 ;
        RECT 25.525 0.625 25.695 1.505 ;
        RECT 26.495 1.425 26.665 1.505 ;
        RECT 26.015 1.080 26.185 1.160 ;
        RECT 27.065 1.080 27.235 1.755 ;
        RECT 28.035 1.750 28.205 5.070 ;
        RECT 32.105 1.915 32.275 4.865 ;
        RECT 26.015 0.910 27.235 1.080 ;
        RECT 26.015 0.830 26.185 0.910 ;
        RECT 26.495 0.625 26.665 0.705 ;
        RECT 25.525 0.455 26.665 0.625 ;
        RECT 25.525 0.375 25.695 0.455 ;
        RECT 26.495 0.375 26.665 0.455 ;
        RECT 27.065 0.625 27.235 0.910 ;
        RECT 27.550 1.580 28.205 1.750 ;
        RECT 29.365 1.675 29.535 1.755 ;
        RECT 30.335 1.675 30.505 1.755 ;
        RECT 31.305 1.675 31.475 1.755 ;
        RECT 27.550 0.845 27.720 1.580 ;
        RECT 29.365 1.505 31.475 1.675 ;
        RECT 28.035 0.625 28.205 1.395 ;
        RECT 27.065 0.455 28.205 0.625 ;
        RECT 27.065 0.375 27.235 0.455 ;
        RECT 28.035 0.375 28.205 0.455 ;
        RECT 29.365 0.375 29.535 1.505 ;
        RECT 30.335 0.625 30.505 1.505 ;
        RECT 31.305 1.425 31.475 1.505 ;
        RECT 30.825 1.080 30.995 1.160 ;
        RECT 31.875 1.080 32.045 1.755 ;
        RECT 32.845 1.750 33.015 5.070 ;
        RECT 34.695 1.915 34.865 4.865 ;
        RECT 36.915 1.915 37.085 4.865 ;
        RECT 30.825 0.910 32.045 1.080 ;
        RECT 30.825 0.830 30.995 0.910 ;
        RECT 31.305 0.625 31.475 0.705 ;
        RECT 30.335 0.455 31.475 0.625 ;
        RECT 30.335 0.375 30.505 0.455 ;
        RECT 31.305 0.375 31.475 0.455 ;
        RECT 31.875 0.625 32.045 0.910 ;
        RECT 32.360 1.580 33.015 1.750 ;
        RECT 34.175 1.675 34.345 1.755 ;
        RECT 35.145 1.675 35.315 1.755 ;
        RECT 36.115 1.675 36.285 1.755 ;
        RECT 32.360 0.845 32.530 1.580 ;
        RECT 34.175 1.505 36.285 1.675 ;
        RECT 32.845 0.625 33.015 1.395 ;
        RECT 31.875 0.455 33.015 0.625 ;
        RECT 31.875 0.375 32.045 0.455 ;
        RECT 32.845 0.375 33.015 0.455 ;
        RECT 34.175 0.375 34.345 1.505 ;
        RECT 35.145 0.625 35.315 1.505 ;
        RECT 36.115 1.425 36.285 1.505 ;
        RECT 35.635 1.080 35.805 1.160 ;
        RECT 36.685 1.080 36.855 1.755 ;
        RECT 37.655 1.750 37.825 5.070 ;
        RECT 39.505 1.915 39.675 4.865 ;
        RECT 41.725 1.915 41.895 4.865 ;
        RECT 35.635 0.910 36.855 1.080 ;
        RECT 35.635 0.830 35.805 0.910 ;
        RECT 36.115 0.625 36.285 0.705 ;
        RECT 35.145 0.455 36.285 0.625 ;
        RECT 35.145 0.375 35.315 0.455 ;
        RECT 36.115 0.375 36.285 0.455 ;
        RECT 36.685 0.625 36.855 0.910 ;
        RECT 37.170 1.580 37.825 1.750 ;
        RECT 38.985 1.675 39.155 1.755 ;
        RECT 39.955 1.675 40.125 1.755 ;
        RECT 40.925 1.675 41.095 1.755 ;
        RECT 37.170 0.845 37.340 1.580 ;
        RECT 38.985 1.505 41.095 1.675 ;
        RECT 37.655 0.625 37.825 1.395 ;
        RECT 36.685 0.455 37.825 0.625 ;
        RECT 36.685 0.375 36.855 0.455 ;
        RECT 37.655 0.375 37.825 0.455 ;
        RECT 38.985 0.375 39.155 1.505 ;
        RECT 39.955 0.625 40.125 1.505 ;
        RECT 40.925 1.425 41.095 1.505 ;
        RECT 40.445 1.080 40.615 1.160 ;
        RECT 41.495 1.080 41.665 1.755 ;
        RECT 42.465 1.750 42.635 5.070 ;
        RECT 44.315 1.915 44.485 4.865 ;
        RECT 40.445 0.910 41.665 1.080 ;
        RECT 40.445 0.830 40.615 0.910 ;
        RECT 40.925 0.625 41.095 0.705 ;
        RECT 39.955 0.455 41.095 0.625 ;
        RECT 39.955 0.375 40.125 0.455 ;
        RECT 40.925 0.375 41.095 0.455 ;
        RECT 41.495 0.625 41.665 0.910 ;
        RECT 41.980 1.580 42.635 1.750 ;
        RECT 43.795 1.675 43.965 1.755 ;
        RECT 44.765 1.675 44.935 1.755 ;
        RECT 45.735 1.675 45.905 1.755 ;
        RECT 41.980 0.845 42.150 1.580 ;
        RECT 43.795 1.505 45.905 1.675 ;
        RECT 42.465 0.625 42.635 1.395 ;
        RECT 41.495 0.455 42.635 0.625 ;
        RECT 41.495 0.375 41.665 0.455 ;
        RECT 42.465 0.375 42.635 0.455 ;
        RECT 43.795 0.375 43.965 1.505 ;
        RECT 44.765 0.625 44.935 1.505 ;
        RECT 45.735 1.425 45.905 1.505 ;
        RECT 45.255 1.080 45.425 1.160 ;
        RECT 46.305 1.080 46.475 1.755 ;
        RECT 47.275 1.750 47.445 5.070 ;
        RECT 49.125 1.915 49.295 4.865 ;
        RECT 51.345 1.915 51.515 4.865 ;
        RECT 45.255 0.910 46.475 1.080 ;
        RECT 45.255 0.830 45.425 0.910 ;
        RECT 45.735 0.625 45.905 0.705 ;
        RECT 44.765 0.455 45.905 0.625 ;
        RECT 44.765 0.375 44.935 0.455 ;
        RECT 45.735 0.375 45.905 0.455 ;
        RECT 46.305 0.625 46.475 0.910 ;
        RECT 46.790 1.580 47.445 1.750 ;
        RECT 48.605 1.675 48.775 1.755 ;
        RECT 49.575 1.675 49.745 1.755 ;
        RECT 50.545 1.675 50.715 1.755 ;
        RECT 46.790 0.845 46.960 1.580 ;
        RECT 48.605 1.505 50.715 1.675 ;
        RECT 47.275 0.625 47.445 1.395 ;
        RECT 46.305 0.455 47.445 0.625 ;
        RECT 46.305 0.375 46.475 0.455 ;
        RECT 47.275 0.375 47.445 0.455 ;
        RECT 48.605 0.375 48.775 1.505 ;
        RECT 49.575 0.625 49.745 1.505 ;
        RECT 50.545 1.425 50.715 1.505 ;
        RECT 50.065 1.080 50.235 1.160 ;
        RECT 51.115 1.080 51.285 1.755 ;
        RECT 52.085 1.750 52.255 5.070 ;
        RECT 53.935 1.915 54.105 4.865 ;
        RECT 56.155 1.915 56.325 4.865 ;
        RECT 50.065 0.910 51.285 1.080 ;
        RECT 50.065 0.830 50.235 0.910 ;
        RECT 50.545 0.625 50.715 0.705 ;
        RECT 49.575 0.455 50.715 0.625 ;
        RECT 49.575 0.375 49.745 0.455 ;
        RECT 50.545 0.375 50.715 0.455 ;
        RECT 51.115 0.625 51.285 0.910 ;
        RECT 51.600 1.580 52.255 1.750 ;
        RECT 53.415 1.675 53.585 1.755 ;
        RECT 54.385 1.675 54.555 1.755 ;
        RECT 55.355 1.675 55.525 1.755 ;
        RECT 51.600 0.845 51.770 1.580 ;
        RECT 53.415 1.505 55.525 1.675 ;
        RECT 52.085 0.625 52.255 1.395 ;
        RECT 51.115 0.455 52.255 0.625 ;
        RECT 51.115 0.375 51.285 0.455 ;
        RECT 52.085 0.375 52.255 0.455 ;
        RECT 53.415 0.375 53.585 1.505 ;
        RECT 54.385 0.625 54.555 1.505 ;
        RECT 55.355 1.425 55.525 1.505 ;
        RECT 54.875 1.080 55.045 1.160 ;
        RECT 55.925 1.080 56.095 1.755 ;
        RECT 56.895 1.750 57.065 5.070 ;
        RECT 60.965 1.915 61.135 4.865 ;
        RECT 54.875 0.910 56.095 1.080 ;
        RECT 54.875 0.830 55.045 0.910 ;
        RECT 55.355 0.625 55.525 0.705 ;
        RECT 54.385 0.455 55.525 0.625 ;
        RECT 54.385 0.375 54.555 0.455 ;
        RECT 55.355 0.375 55.525 0.455 ;
        RECT 55.925 0.625 56.095 0.910 ;
        RECT 56.410 1.580 57.065 1.750 ;
        RECT 58.225 1.675 58.395 1.755 ;
        RECT 59.195 1.675 59.365 1.755 ;
        RECT 60.165 1.675 60.335 1.755 ;
        RECT 56.410 0.845 56.580 1.580 ;
        RECT 58.225 1.505 60.335 1.675 ;
        RECT 56.895 0.625 57.065 1.395 ;
        RECT 55.925 0.455 57.065 0.625 ;
        RECT 55.925 0.375 56.095 0.455 ;
        RECT 56.895 0.375 57.065 0.455 ;
        RECT 58.225 0.375 58.395 1.505 ;
        RECT 59.195 0.625 59.365 1.505 ;
        RECT 60.165 1.425 60.335 1.505 ;
        RECT 59.685 1.080 59.855 1.160 ;
        RECT 60.735 1.080 60.905 1.755 ;
        RECT 61.705 1.750 61.875 5.070 ;
        RECT 63.555 1.915 63.725 4.865 ;
        RECT 65.775 1.915 65.945 4.865 ;
        RECT 59.685 0.910 60.905 1.080 ;
        RECT 59.685 0.830 59.855 0.910 ;
        RECT 60.165 0.625 60.335 0.705 ;
        RECT 59.195 0.455 60.335 0.625 ;
        RECT 59.195 0.375 59.365 0.455 ;
        RECT 60.165 0.375 60.335 0.455 ;
        RECT 60.735 0.625 60.905 0.910 ;
        RECT 61.220 1.580 61.875 1.750 ;
        RECT 63.035 1.675 63.205 1.755 ;
        RECT 64.005 1.675 64.175 1.755 ;
        RECT 64.975 1.675 65.145 1.755 ;
        RECT 61.220 0.845 61.390 1.580 ;
        RECT 63.035 1.505 65.145 1.675 ;
        RECT 61.705 0.625 61.875 1.395 ;
        RECT 60.735 0.455 61.875 0.625 ;
        RECT 60.735 0.375 60.905 0.455 ;
        RECT 61.705 0.375 61.875 0.455 ;
        RECT 63.035 0.375 63.205 1.505 ;
        RECT 64.005 0.625 64.175 1.505 ;
        RECT 64.975 1.425 65.145 1.505 ;
        RECT 64.495 1.080 64.665 1.160 ;
        RECT 65.545 1.080 65.715 1.755 ;
        RECT 66.515 1.750 66.685 5.070 ;
        RECT 68.365 1.915 68.535 4.865 ;
        RECT 70.585 1.915 70.755 4.865 ;
        RECT 64.495 0.910 65.715 1.080 ;
        RECT 64.495 0.830 64.665 0.910 ;
        RECT 64.975 0.625 65.145 0.705 ;
        RECT 64.005 0.455 65.145 0.625 ;
        RECT 64.005 0.375 64.175 0.455 ;
        RECT 64.975 0.375 65.145 0.455 ;
        RECT 65.545 0.625 65.715 0.910 ;
        RECT 66.030 1.580 66.685 1.750 ;
        RECT 67.845 1.675 68.015 1.755 ;
        RECT 68.815 1.675 68.985 1.755 ;
        RECT 69.785 1.675 69.955 1.755 ;
        RECT 66.030 0.845 66.200 1.580 ;
        RECT 67.845 1.505 69.955 1.675 ;
        RECT 66.515 0.625 66.685 1.395 ;
        RECT 65.545 0.455 66.685 0.625 ;
        RECT 65.545 0.375 65.715 0.455 ;
        RECT 66.515 0.375 66.685 0.455 ;
        RECT 67.845 0.375 68.015 1.505 ;
        RECT 68.815 0.625 68.985 1.505 ;
        RECT 69.785 1.425 69.955 1.505 ;
        RECT 69.305 1.080 69.475 1.160 ;
        RECT 70.355 1.080 70.525 1.755 ;
        RECT 71.325 1.750 71.495 5.070 ;
        RECT 73.175 1.915 73.345 4.865 ;
        RECT 69.305 0.910 70.525 1.080 ;
        RECT 69.305 0.830 69.475 0.910 ;
        RECT 69.785 0.625 69.955 0.705 ;
        RECT 68.815 0.455 69.955 0.625 ;
        RECT 68.815 0.375 68.985 0.455 ;
        RECT 69.785 0.375 69.955 0.455 ;
        RECT 70.355 0.625 70.525 0.910 ;
        RECT 70.840 1.580 71.495 1.750 ;
        RECT 72.655 1.675 72.825 1.755 ;
        RECT 73.625 1.675 73.795 1.755 ;
        RECT 74.595 1.675 74.765 1.755 ;
        RECT 70.840 0.845 71.010 1.580 ;
        RECT 72.655 1.505 74.765 1.675 ;
        RECT 71.325 0.625 71.495 1.395 ;
        RECT 70.355 0.455 71.495 0.625 ;
        RECT 70.355 0.375 70.525 0.455 ;
        RECT 71.325 0.375 71.495 0.455 ;
        RECT 72.655 0.375 72.825 1.505 ;
        RECT 73.625 0.625 73.795 1.505 ;
        RECT 74.595 1.425 74.765 1.505 ;
        RECT 74.115 1.080 74.285 1.160 ;
        RECT 75.165 1.080 75.335 1.755 ;
        RECT 76.135 1.750 76.305 5.070 ;
        RECT 77.985 1.915 78.155 4.865 ;
        RECT 80.205 1.915 80.375 4.865 ;
        RECT 74.115 0.910 75.335 1.080 ;
        RECT 74.115 0.830 74.285 0.910 ;
        RECT 74.595 0.625 74.765 0.705 ;
        RECT 73.625 0.455 74.765 0.625 ;
        RECT 73.625 0.375 73.795 0.455 ;
        RECT 74.595 0.375 74.765 0.455 ;
        RECT 75.165 0.625 75.335 0.910 ;
        RECT 75.650 1.580 76.305 1.750 ;
        RECT 77.465 1.675 77.635 1.755 ;
        RECT 78.435 1.675 78.605 1.755 ;
        RECT 79.405 1.675 79.575 1.755 ;
        RECT 75.650 0.845 75.820 1.580 ;
        RECT 77.465 1.505 79.575 1.675 ;
        RECT 76.135 0.625 76.305 1.395 ;
        RECT 75.165 0.455 76.305 0.625 ;
        RECT 75.165 0.375 75.335 0.455 ;
        RECT 76.135 0.375 76.305 0.455 ;
        RECT 77.465 0.375 77.635 1.505 ;
        RECT 78.435 0.625 78.605 1.505 ;
        RECT 79.405 1.425 79.575 1.505 ;
        RECT 78.925 1.080 79.095 1.160 ;
        RECT 79.975 1.080 80.145 1.755 ;
        RECT 80.945 1.750 81.115 5.070 ;
        RECT 82.795 1.915 82.965 4.865 ;
        RECT 85.015 1.915 85.185 4.865 ;
        RECT 78.925 0.910 80.145 1.080 ;
        RECT 78.925 0.830 79.095 0.910 ;
        RECT 79.405 0.625 79.575 0.705 ;
        RECT 78.435 0.455 79.575 0.625 ;
        RECT 78.435 0.375 78.605 0.455 ;
        RECT 79.405 0.375 79.575 0.455 ;
        RECT 79.975 0.625 80.145 0.910 ;
        RECT 80.460 1.580 81.115 1.750 ;
        RECT 82.275 1.675 82.445 1.755 ;
        RECT 83.245 1.675 83.415 1.755 ;
        RECT 84.215 1.675 84.385 1.755 ;
        RECT 80.460 0.845 80.630 1.580 ;
        RECT 82.275 1.505 84.385 1.675 ;
        RECT 80.945 0.625 81.115 1.395 ;
        RECT 79.975 0.455 81.115 0.625 ;
        RECT 79.975 0.375 80.145 0.455 ;
        RECT 80.945 0.375 81.115 0.455 ;
        RECT 82.275 0.375 82.445 1.505 ;
        RECT 83.245 0.625 83.415 1.505 ;
        RECT 84.215 1.425 84.385 1.505 ;
        RECT 83.735 1.080 83.905 1.160 ;
        RECT 84.785 1.080 84.955 1.755 ;
        RECT 85.755 1.750 85.925 5.070 ;
        RECT 88.605 5.045 88.775 5.125 ;
        RECT 90.605 6.825 92.535 6.995 ;
        RECT 90.605 5.045 90.775 6.825 ;
        RECT 91.045 5.295 91.215 6.565 ;
        RECT 91.485 5.555 91.655 6.825 ;
        RECT 91.925 5.295 92.095 6.565 ;
        RECT 92.365 5.375 92.535 6.825 ;
        RECT 93.945 6.825 95.875 6.995 ;
        RECT 91.045 5.125 92.095 5.295 ;
        RECT 91.925 5.045 92.095 5.125 ;
        RECT 93.945 5.045 94.115 6.825 ;
        RECT 94.825 5.555 94.995 6.825 ;
        RECT 95.705 5.555 95.875 6.825 ;
        RECT 87.235 1.915 87.405 4.870 ;
        RECT 88.385 4.710 88.555 4.870 ;
        RECT 88.345 4.540 88.555 4.710 ;
        RECT 88.345 1.915 88.515 4.540 ;
        RECT 90.935 1.915 91.105 4.870 ;
        RECT 92.415 1.915 92.585 4.870 ;
        RECT 93.895 1.915 94.065 4.870 ;
        RECT 95.005 4.540 95.195 4.870 ;
        RECT 95.005 1.915 95.175 4.540 ;
        RECT 83.735 0.910 84.955 1.080 ;
        RECT 83.735 0.830 83.905 0.910 ;
        RECT 84.215 0.625 84.385 0.705 ;
        RECT 83.245 0.455 84.385 0.625 ;
        RECT 83.245 0.375 83.415 0.455 ;
        RECT 84.215 0.375 84.385 0.455 ;
        RECT 84.785 0.625 84.955 0.910 ;
        RECT 85.270 1.580 85.925 1.750 ;
        RECT 87.190 1.665 87.360 1.745 ;
        RECT 88.160 1.665 88.330 1.745 ;
        RECT 85.270 0.845 85.440 1.580 ;
        RECT 87.190 1.495 88.330 1.665 ;
        RECT 85.755 0.625 85.925 1.395 ;
        RECT 84.785 0.455 85.925 0.625 ;
        RECT 84.785 0.375 84.955 0.455 ;
        RECT 85.755 0.375 85.925 0.455 ;
        RECT 87.190 0.365 87.360 1.495 ;
        RECT 88.160 0.615 88.330 1.495 ;
        RECT 89.130 0.615 89.300 1.745 ;
        RECT 88.160 0.445 89.300 0.615 ;
        RECT 88.160 0.365 88.330 0.445 ;
        RECT 89.130 0.365 89.300 0.445 ;
        RECT 90.520 1.665 90.690 1.745 ;
        RECT 91.490 1.665 91.660 1.745 ;
        RECT 90.520 1.495 91.660 1.665 ;
        RECT 90.520 0.365 90.690 1.495 ;
        RECT 91.490 0.615 91.660 1.495 ;
        RECT 92.460 0.615 92.630 1.745 ;
        RECT 91.490 0.445 92.630 0.615 ;
        RECT 91.490 0.365 91.660 0.445 ;
        RECT 92.460 0.365 92.630 0.445 ;
        RECT 93.850 1.665 94.020 1.745 ;
        RECT 94.820 1.665 94.990 1.745 ;
        RECT 93.850 1.495 94.990 1.665 ;
        RECT 93.850 0.365 94.020 1.495 ;
        RECT 94.820 0.615 94.990 1.495 ;
        RECT 95.790 0.615 95.960 1.390 ;
        RECT 94.820 0.445 95.960 0.615 ;
        RECT 94.820 0.365 94.990 0.445 ;
        RECT 95.790 0.365 95.960 0.445 ;
      LAYER mcon ;
        RECT 88.605 5.125 88.775 5.295 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 2.505 4.155 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 8.055 3.615 8.225 3.785 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 10.645 2.505 10.815 2.675 ;
        RECT 12.865 3.615 13.035 3.785 ;
        RECT 13.605 2.505 13.775 2.675 ;
        RECT 15.455 2.505 15.625 2.675 ;
        RECT 18.415 3.615 18.585 3.785 ;
        RECT 20.265 3.245 20.435 3.415 ;
        RECT 22.485 3.245 22.655 3.415 ;
        RECT 23.225 4.725 23.395 4.895 ;
        RECT 23.225 2.505 23.395 2.675 ;
        RECT 25.075 2.505 25.245 2.675 ;
        RECT 27.295 3.615 27.465 3.785 ;
        RECT 28.035 3.245 28.205 3.415 ;
        RECT 32.105 3.245 32.275 3.415 ;
        RECT 32.845 2.505 33.015 2.675 ;
        RECT 34.695 2.505 34.865 2.675 ;
        RECT 36.915 3.615 37.085 3.785 ;
        RECT 37.655 3.245 37.825 3.415 ;
        RECT 39.505 2.505 39.675 2.675 ;
        RECT 41.725 3.615 41.895 3.785 ;
        RECT 42.465 2.505 42.635 2.675 ;
        RECT 44.315 2.505 44.485 2.675 ;
        RECT 47.275 3.615 47.445 3.785 ;
        RECT 49.125 3.245 49.295 3.415 ;
        RECT 51.345 2.505 51.515 2.675 ;
        RECT 52.085 3.245 52.255 3.415 ;
        RECT 53.935 3.245 54.105 3.415 ;
        RECT 56.155 3.615 56.325 3.785 ;
        RECT 56.895 2.505 57.065 2.675 ;
        RECT 60.965 3.245 61.135 3.415 ;
        RECT 61.705 2.505 61.875 2.675 ;
        RECT 63.555 2.505 63.725 2.675 ;
        RECT 65.775 3.615 65.945 3.785 ;
        RECT 66.515 3.245 66.685 3.415 ;
        RECT 68.365 2.505 68.535 2.675 ;
        RECT 70.585 3.615 70.755 3.785 ;
        RECT 71.325 2.505 71.495 2.675 ;
        RECT 73.175 2.505 73.345 2.675 ;
        RECT 76.135 3.615 76.305 3.785 ;
        RECT 77.985 3.245 78.155 3.415 ;
        RECT 80.205 2.505 80.375 2.675 ;
        RECT 80.945 2.135 81.115 2.305 ;
        RECT 82.795 2.135 82.965 2.305 ;
        RECT 85.015 3.615 85.185 3.785 ;
        RECT 90.605 5.125 90.775 5.295 ;
        RECT 91.925 5.125 92.095 5.295 ;
        RECT 93.945 5.125 94.115 5.295 ;
        RECT 85.755 2.505 85.925 2.675 ;
        RECT 87.235 4.355 87.405 4.525 ;
        RECT 88.345 3.985 88.515 4.155 ;
        RECT 90.935 4.355 91.105 4.525 ;
        RECT 92.415 1.995 92.585 2.165 ;
        RECT 93.895 1.995 94.065 2.165 ;
        RECT 95.005 3.985 95.175 4.155 ;
      LAYER met1 ;
        RECT 88.575 5.295 88.805 5.325 ;
        RECT 90.575 5.295 90.805 5.325 ;
        RECT 91.895 5.295 92.125 5.325 ;
        RECT 93.915 5.295 94.145 5.325 ;
        RECT 88.545 5.125 90.835 5.295 ;
        RECT 91.865 5.125 94.175 5.295 ;
        RECT 88.575 5.095 88.805 5.125 ;
        RECT 90.575 5.095 90.805 5.125 ;
        RECT 91.895 5.095 92.125 5.125 ;
        RECT 93.915 5.095 94.145 5.125 ;
        RECT 23.195 4.895 23.425 4.925 ;
        RECT 23.165 4.725 75.195 4.895 ;
        RECT 23.195 4.695 23.425 4.725 ;
        RECT 75.025 4.525 75.195 4.725 ;
        RECT 87.205 4.525 87.435 4.555 ;
        RECT 90.905 4.525 91.135 4.555 ;
        RECT 75.025 4.365 91.165 4.525 ;
        RECT 75.105 4.355 91.165 4.365 ;
        RECT 87.205 4.325 87.435 4.355 ;
        RECT 90.905 4.325 91.135 4.355 ;
        RECT 88.315 4.155 88.545 4.185 ;
        RECT 94.975 4.155 95.205 4.185 ;
        RECT 65.035 3.985 95.235 4.155 ;
        RECT 8.025 3.785 8.255 3.815 ;
        RECT 12.835 3.785 13.065 3.815 ;
        RECT 18.385 3.785 18.615 3.815 ;
        RECT 27.265 3.785 27.495 3.815 ;
        RECT 36.885 3.785 37.115 3.815 ;
        RECT 41.695 3.785 41.925 3.815 ;
        RECT 47.245 3.785 47.475 3.815 ;
        RECT 56.125 3.785 56.355 3.815 ;
        RECT 65.035 3.785 65.205 3.985 ;
        RECT 88.315 3.955 88.545 3.985 ;
        RECT 94.975 3.955 95.205 3.985 ;
        RECT 65.745 3.785 65.975 3.815 ;
        RECT 70.555 3.785 70.785 3.815 ;
        RECT 76.105 3.785 76.335 3.815 ;
        RECT 84.985 3.785 85.215 3.815 ;
        RECT 7.995 3.615 27.525 3.785 ;
        RECT 36.855 3.615 56.385 3.785 ;
        RECT 56.895 3.615 65.205 3.785 ;
        RECT 65.715 3.615 85.245 3.785 ;
        RECT 8.025 3.585 8.255 3.615 ;
        RECT 12.835 3.585 13.065 3.615 ;
        RECT 18.385 3.585 18.615 3.615 ;
        RECT 27.265 3.585 27.495 3.615 ;
        RECT 36.885 3.585 37.115 3.615 ;
        RECT 41.695 3.585 41.925 3.615 ;
        RECT 47.245 3.585 47.475 3.615 ;
        RECT 56.125 3.585 56.355 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 8.765 3.415 8.995 3.445 ;
        RECT 20.235 3.415 20.465 3.445 ;
        RECT 22.455 3.415 22.685 3.445 ;
        RECT 28.005 3.415 28.235 3.445 ;
        RECT 32.075 3.415 32.305 3.445 ;
        RECT 37.625 3.415 37.855 3.445 ;
        RECT 49.095 3.415 49.325 3.445 ;
        RECT 52.055 3.415 52.285 3.445 ;
        RECT 53.905 3.415 54.135 3.445 ;
        RECT 56.895 3.415 57.065 3.615 ;
        RECT 65.745 3.585 65.975 3.615 ;
        RECT 70.555 3.585 70.785 3.615 ;
        RECT 76.105 3.585 76.335 3.615 ;
        RECT 84.985 3.585 85.215 3.615 ;
        RECT 60.935 3.415 61.165 3.445 ;
        RECT 66.485 3.415 66.715 3.445 ;
        RECT 77.955 3.415 78.185 3.445 ;
        RECT 3.185 3.245 20.495 3.415 ;
        RECT 22.425 3.245 28.265 3.415 ;
        RECT 32.045 3.245 49.355 3.415 ;
        RECT 52.025 3.245 57.065 3.415 ;
        RECT 60.905 3.245 78.215 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 8.765 3.215 8.995 3.245 ;
        RECT 20.235 3.215 20.465 3.245 ;
        RECT 22.455 3.215 22.685 3.245 ;
        RECT 28.005 3.215 28.235 3.245 ;
        RECT 32.075 3.215 32.305 3.245 ;
        RECT 37.625 3.215 37.855 3.245 ;
        RECT 49.095 3.215 49.325 3.245 ;
        RECT 52.055 3.215 52.285 3.245 ;
        RECT 53.905 3.215 54.135 3.245 ;
        RECT 60.935 3.215 61.165 3.245 ;
        RECT 66.485 3.215 66.715 3.245 ;
        RECT 77.955 3.215 78.185 3.245 ;
        RECT 3.955 2.675 4.185 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 10.615 2.675 10.845 2.705 ;
        RECT 13.575 2.675 13.805 2.705 ;
        RECT 15.425 2.675 15.655 2.705 ;
        RECT 23.195 2.675 23.425 2.705 ;
        RECT 25.045 2.675 25.275 2.705 ;
        RECT 32.815 2.675 33.045 2.705 ;
        RECT 34.665 2.675 34.895 2.705 ;
        RECT 39.475 2.675 39.705 2.705 ;
        RECT 42.435 2.675 42.665 2.705 ;
        RECT 44.285 2.675 44.515 2.705 ;
        RECT 51.315 2.675 51.545 2.705 ;
        RECT 56.865 2.675 57.095 2.705 ;
        RECT 61.675 2.675 61.905 2.705 ;
        RECT 63.525 2.675 63.755 2.705 ;
        RECT 68.335 2.675 68.565 2.705 ;
        RECT 71.295 2.675 71.525 2.705 ;
        RECT 73.145 2.675 73.375 2.705 ;
        RECT 80.175 2.675 80.405 2.705 ;
        RECT 85.725 2.675 85.955 2.705 ;
        RECT 3.925 2.505 10.875 2.675 ;
        RECT 13.545 2.505 15.685 2.675 ;
        RECT 23.165 2.505 25.305 2.675 ;
        RECT 32.785 2.505 39.735 2.675 ;
        RECT 42.405 2.505 44.545 2.675 ;
        RECT 51.285 2.505 57.125 2.675 ;
        RECT 61.645 2.505 68.595 2.675 ;
        RECT 71.265 2.505 73.405 2.675 ;
        RECT 80.145 2.505 85.985 2.675 ;
        RECT 3.955 2.475 4.185 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 10.615 2.475 10.845 2.505 ;
        RECT 13.575 2.475 13.805 2.505 ;
        RECT 15.425 2.475 15.655 2.505 ;
        RECT 23.195 2.475 23.425 2.505 ;
        RECT 25.045 2.475 25.275 2.505 ;
        RECT 32.815 2.475 33.045 2.505 ;
        RECT 34.665 2.475 34.895 2.505 ;
        RECT 39.475 2.475 39.705 2.505 ;
        RECT 42.435 2.475 42.665 2.505 ;
        RECT 44.285 2.475 44.515 2.505 ;
        RECT 51.315 2.475 51.545 2.505 ;
        RECT 56.865 2.475 57.095 2.505 ;
        RECT 61.675 2.475 61.905 2.505 ;
        RECT 63.525 2.475 63.755 2.505 ;
        RECT 68.335 2.475 68.565 2.505 ;
        RECT 71.295 2.475 71.525 2.505 ;
        RECT 73.145 2.475 73.375 2.505 ;
        RECT 80.175 2.475 80.405 2.505 ;
        RECT 85.725 2.475 85.955 2.505 ;
        RECT 80.915 2.305 81.145 2.335 ;
        RECT 82.765 2.305 82.995 2.335 ;
        RECT 80.885 2.165 92.615 2.305 ;
        RECT 93.865 2.165 94.095 2.195 ;
        RECT 80.885 2.135 94.125 2.165 ;
        RECT 80.915 2.105 81.145 2.135 ;
        RECT 82.765 2.105 82.995 2.135 ;
        RECT 92.355 1.995 94.125 2.135 ;
        RECT 92.385 1.965 92.615 1.995 ;
        RECT 93.865 1.965 94.095 1.995 ;
  END
END TMRDFFSNRNQNX1






MACRO TMRDFFSNRNQX1
  CLASS CORE ;
  FOREIGN TMRDFFSNRNQX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 98.790 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 97.600 4.665 97.770 7.020 ;
        RECT 97.600 4.495 98.135 4.665 ;
        RECT 97.965 2.165 98.135 4.495 ;
        RECT 97.595 1.995 98.135 2.165 ;
        RECT 97.595 0.840 97.765 1.995 ;
      LAYER mcon ;
        RECT 97.965 3.985 98.135 4.155 ;
      LAYER met1 ;
        RECT 97.935 4.155 98.165 4.185 ;
        RECT 97.905 3.985 98.315 4.155 ;
        RECT 97.935 3.955 98.165 3.985 ;
    END
  END Q
  PIN SN
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 11.755 1.915 11.925 4.865 ;
        RECT 26.185 1.915 26.355 4.865 ;
        RECT 40.615 1.915 40.785 4.865 ;
        RECT 55.045 1.915 55.215 4.865 ;
        RECT 69.475 1.915 69.645 4.865 ;
        RECT 83.905 1.915 84.075 4.865 ;
      LAYER mcon ;
        RECT 11.755 2.875 11.925 3.045 ;
        RECT 26.185 2.875 26.355 3.045 ;
        RECT 40.615 2.875 40.785 3.045 ;
        RECT 55.045 2.875 55.215 3.045 ;
        RECT 69.475 2.875 69.645 3.045 ;
        RECT 83.905 2.875 84.075 3.045 ;
      LAYER met1 ;
        RECT 11.725 3.045 11.955 3.075 ;
        RECT 26.155 3.045 26.385 3.075 ;
        RECT 40.585 3.045 40.815 3.075 ;
        RECT 55.015 3.045 55.245 3.075 ;
        RECT 69.445 3.045 69.675 3.075 ;
        RECT 83.875 3.045 84.105 3.075 ;
        RECT 11.695 2.875 84.135 3.045 ;
        RECT 11.725 2.845 11.955 2.875 ;
        RECT 26.155 2.845 26.385 2.875 ;
        RECT 40.585 2.845 40.815 2.875 ;
        RECT 55.015 2.845 55.245 2.875 ;
        RECT 69.445 2.845 69.675 2.875 ;
        RECT 83.875 2.845 84.105 2.875 ;
    END
  END SN
  PIN RN
    ANTENNAGATEAREA 9.170850 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 17.675 1.915 17.845 4.865 ;
        RECT 21.375 1.915 21.545 4.865 ;
        RECT 30.995 1.915 31.165 4.865 ;
        RECT 46.535 1.915 46.705 4.865 ;
        RECT 50.235 1.915 50.405 4.865 ;
        RECT 59.855 1.915 60.025 4.865 ;
        RECT 75.395 1.915 75.565 4.865 ;
        RECT 79.095 1.915 79.265 4.865 ;
      LAYER mcon ;
        RECT 2.135 2.135 2.305 2.305 ;
        RECT 17.675 2.135 17.845 2.305 ;
        RECT 21.375 2.135 21.545 2.305 ;
        RECT 30.995 2.135 31.165 2.305 ;
        RECT 46.535 2.135 46.705 2.305 ;
        RECT 50.235 2.135 50.405 2.305 ;
        RECT 59.855 2.135 60.025 2.305 ;
        RECT 75.395 2.135 75.565 2.305 ;
        RECT 79.095 2.135 79.265 2.305 ;
      LAYER met1 ;
        RECT 2.105 2.305 2.335 2.335 ;
        RECT 17.645 2.305 17.875 2.335 ;
        RECT 21.345 2.305 21.575 2.335 ;
        RECT 30.965 2.305 31.195 2.335 ;
        RECT 46.505 2.305 46.735 2.335 ;
        RECT 50.205 2.305 50.435 2.335 ;
        RECT 59.825 2.305 60.055 2.335 ;
        RECT 75.365 2.305 75.595 2.335 ;
        RECT 79.065 2.305 79.295 2.335 ;
        RECT 2.075 2.135 79.325 2.305 ;
        RECT 2.105 2.105 2.335 2.135 ;
        RECT 17.645 2.105 17.875 2.135 ;
        RECT 21.345 2.105 21.575 2.135 ;
        RECT 30.965 2.105 31.195 2.135 ;
        RECT 46.505 2.105 46.735 2.135 ;
        RECT 50.205 2.105 50.435 2.135 ;
        RECT 59.825 2.105 60.055 2.135 ;
        RECT 75.365 2.105 75.595 2.135 ;
        RECT 79.065 2.105 79.295 2.135 ;
    END
  END RN
  PIN D
    ANTENNAGATEAREA 3.099750 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 29.885 1.915 30.055 4.865 ;
        RECT 58.745 1.915 58.915 4.865 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 29.885 3.985 30.055 4.155 ;
        RECT 58.745 3.985 58.915 4.155 ;
      LAYER met1 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 29.855 4.155 30.085 4.185 ;
        RECT 58.715 4.155 58.945 4.185 ;
        RECT 0.845 3.985 58.975 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 29.855 3.955 30.085 3.985 ;
        RECT 58.715 3.955 58.945 3.985 ;
    END
  END D
  PIN CLK
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 16.565 1.915 16.735 4.865 ;
        RECT 35.805 1.915 35.975 4.865 ;
        RECT 45.425 1.915 45.595 4.865 ;
        RECT 64.665 1.915 64.835 4.865 ;
        RECT 74.285 1.915 74.455 4.865 ;
      LAYER mcon ;
        RECT 6.945 4.355 7.115 4.525 ;
        RECT 16.565 4.355 16.735 4.525 ;
        RECT 35.805 4.355 35.975 4.525 ;
        RECT 45.425 4.355 45.595 4.525 ;
        RECT 64.665 4.355 64.835 4.525 ;
        RECT 74.285 4.355 74.455 4.525 ;
      LAYER met1 ;
        RECT 6.915 4.525 7.145 4.555 ;
        RECT 16.535 4.525 16.765 4.555 ;
        RECT 35.775 4.525 36.005 4.555 ;
        RECT 45.395 4.525 45.625 4.555 ;
        RECT 64.635 4.525 64.865 4.555 ;
        RECT 74.255 4.525 74.485 4.555 ;
        RECT 6.885 4.355 74.515 4.525 ;
        RECT 6.915 4.325 7.145 4.355 ;
        RECT 16.535 4.325 16.765 4.355 ;
        RECT 35.775 4.325 36.005 4.355 ;
        RECT 45.395 4.325 45.625 4.355 ;
        RECT 64.635 4.325 64.865 4.355 ;
        RECT 74.255 4.325 74.485 4.355 ;
    END
  END CLK
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 99.225 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 98.960 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.625 5.215 10.795 7.230 ;
        RECT 11.505 5.555 11.675 7.230 ;
        RECT 12.385 5.555 12.555 7.230 ;
        RECT 13.265 5.555 13.435 7.230 ;
        RECT 14.260 4.110 14.600 7.230 ;
        RECT 15.435 5.215 15.605 7.230 ;
        RECT 16.315 5.555 16.485 7.230 ;
        RECT 17.195 5.555 17.365 7.230 ;
        RECT 18.075 5.555 18.245 7.230 ;
        RECT 19.070 4.110 19.410 7.230 ;
        RECT 20.245 5.215 20.415 7.230 ;
        RECT 21.125 5.555 21.295 7.230 ;
        RECT 22.005 5.555 22.175 7.230 ;
        RECT 22.885 5.555 23.055 7.230 ;
        RECT 23.880 4.110 24.220 7.230 ;
        RECT 25.055 5.215 25.225 7.230 ;
        RECT 25.935 5.555 26.105 7.230 ;
        RECT 26.815 5.555 26.985 7.230 ;
        RECT 27.695 5.555 27.865 7.230 ;
        RECT 28.690 4.110 29.030 7.230 ;
        RECT 29.865 5.215 30.035 7.230 ;
        RECT 30.745 5.555 30.915 7.230 ;
        RECT 31.625 5.555 31.795 7.230 ;
        RECT 32.505 5.555 32.675 7.230 ;
        RECT 33.500 4.110 33.840 7.230 ;
        RECT 34.675 5.215 34.845 7.230 ;
        RECT 35.555 5.555 35.725 7.230 ;
        RECT 36.435 5.555 36.605 7.230 ;
        RECT 37.315 5.555 37.485 7.230 ;
        RECT 38.310 4.110 38.650 7.230 ;
        RECT 39.485 5.215 39.655 7.230 ;
        RECT 40.365 5.555 40.535 7.230 ;
        RECT 41.245 5.555 41.415 7.230 ;
        RECT 42.125 5.555 42.295 7.230 ;
        RECT 43.120 4.110 43.460 7.230 ;
        RECT 44.295 5.215 44.465 7.230 ;
        RECT 45.175 5.555 45.345 7.230 ;
        RECT 46.055 5.555 46.225 7.230 ;
        RECT 46.935 5.555 47.105 7.230 ;
        RECT 47.930 4.110 48.270 7.230 ;
        RECT 49.105 5.215 49.275 7.230 ;
        RECT 49.985 5.555 50.155 7.230 ;
        RECT 50.865 5.555 51.035 7.230 ;
        RECT 51.745 5.555 51.915 7.230 ;
        RECT 52.740 4.110 53.080 7.230 ;
        RECT 53.915 5.215 54.085 7.230 ;
        RECT 54.795 5.555 54.965 7.230 ;
        RECT 55.675 5.555 55.845 7.230 ;
        RECT 56.555 5.555 56.725 7.230 ;
        RECT 57.550 4.110 57.890 7.230 ;
        RECT 58.725 5.215 58.895 7.230 ;
        RECT 59.605 5.555 59.775 7.230 ;
        RECT 60.485 5.555 60.655 7.230 ;
        RECT 61.365 5.555 61.535 7.230 ;
        RECT 62.360 4.110 62.700 7.230 ;
        RECT 63.535 5.215 63.705 7.230 ;
        RECT 64.415 5.555 64.585 7.230 ;
        RECT 65.295 5.555 65.465 7.230 ;
        RECT 66.175 5.555 66.345 7.230 ;
        RECT 67.170 4.110 67.510 7.230 ;
        RECT 68.345 5.215 68.515 7.230 ;
        RECT 69.225 5.555 69.395 7.230 ;
        RECT 70.105 5.555 70.275 7.230 ;
        RECT 70.985 5.555 71.155 7.230 ;
        RECT 71.980 4.110 72.320 7.230 ;
        RECT 73.155 5.215 73.325 7.230 ;
        RECT 74.035 5.555 74.205 7.230 ;
        RECT 74.915 5.555 75.085 7.230 ;
        RECT 75.795 5.555 75.965 7.230 ;
        RECT 76.790 4.110 77.130 7.230 ;
        RECT 77.965 5.215 78.135 7.230 ;
        RECT 78.845 5.555 79.015 7.230 ;
        RECT 79.725 5.555 79.895 7.230 ;
        RECT 80.605 5.555 80.775 7.230 ;
        RECT 81.600 4.110 81.940 7.230 ;
        RECT 82.775 5.215 82.945 7.230 ;
        RECT 83.655 5.555 83.825 7.230 ;
        RECT 84.535 5.555 84.705 7.230 ;
        RECT 85.415 5.555 85.585 7.230 ;
        RECT 86.410 4.110 86.750 7.230 ;
        RECT 87.285 5.125 87.455 7.230 ;
        RECT 88.165 5.555 88.335 7.230 ;
        RECT 89.045 5.125 89.215 7.230 ;
        RECT 89.740 4.110 90.080 7.230 ;
        RECT 93.070 4.110 93.410 7.230 ;
        RECT 96.400 4.110 96.740 7.230 ;
        RECT 97.160 5.185 97.330 7.230 ;
        RECT 98.040 5.185 98.210 7.230 ;
        RECT 98.620 4.110 98.960 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.515 7.315 29.685 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.625 7.315 30.795 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 32.845 7.315 33.015 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.435 7.315 35.605 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.175 7.315 36.345 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.765 7.315 38.935 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.505 7.315 39.675 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.615 7.315 40.785 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 42.835 7.315 43.005 7.485 ;
        RECT 43.575 7.315 43.745 7.485 ;
        RECT 43.945 7.315 44.115 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 47.645 7.315 47.815 7.485 ;
        RECT 48.385 7.315 48.555 7.485 ;
        RECT 48.755 7.315 48.925 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 50.975 7.315 51.145 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 51.715 7.315 51.885 7.485 ;
        RECT 52.085 7.315 52.255 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.305 7.315 54.475 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.525 7.315 56.695 7.485 ;
        RECT 56.895 7.315 57.065 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 60.965 7.315 61.135 7.485 ;
        RECT 61.335 7.315 61.505 7.485 ;
        RECT 61.705 7.315 61.875 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.295 7.315 64.465 7.485 ;
        RECT 64.665 7.315 64.835 7.485 ;
        RECT 65.035 7.315 65.205 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.625 7.315 67.795 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.365 7.315 68.535 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.475 7.315 69.645 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 70.955 7.315 71.125 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.175 7.315 73.345 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
        RECT 74.285 7.315 74.455 7.485 ;
        RECT 74.655 7.315 74.825 7.485 ;
        RECT 75.025 7.315 75.195 7.485 ;
        RECT 75.395 7.315 75.565 7.485 ;
        RECT 75.765 7.315 75.935 7.485 ;
        RECT 76.135 7.315 76.305 7.485 ;
        RECT 76.505 7.315 76.675 7.485 ;
        RECT 77.245 7.315 77.415 7.485 ;
        RECT 77.615 7.315 77.785 7.485 ;
        RECT 77.985 7.315 78.155 7.485 ;
        RECT 78.355 7.315 78.525 7.485 ;
        RECT 78.725 7.315 78.895 7.485 ;
        RECT 79.095 7.315 79.265 7.485 ;
        RECT 79.465 7.315 79.635 7.485 ;
        RECT 79.835 7.315 80.005 7.485 ;
        RECT 80.205 7.315 80.375 7.485 ;
        RECT 80.575 7.315 80.745 7.485 ;
        RECT 80.945 7.315 81.115 7.485 ;
        RECT 81.315 7.315 81.485 7.485 ;
        RECT 82.055 7.315 82.225 7.485 ;
        RECT 82.425 7.315 82.595 7.485 ;
        RECT 82.795 7.315 82.965 7.485 ;
        RECT 83.165 7.315 83.335 7.485 ;
        RECT 83.535 7.315 83.705 7.485 ;
        RECT 83.905 7.315 84.075 7.485 ;
        RECT 84.275 7.315 84.445 7.485 ;
        RECT 84.645 7.315 84.815 7.485 ;
        RECT 85.015 7.315 85.185 7.485 ;
        RECT 85.385 7.315 85.555 7.485 ;
        RECT 85.755 7.315 85.925 7.485 ;
        RECT 86.125 7.315 86.295 7.485 ;
        RECT 86.865 7.315 87.035 7.485 ;
        RECT 87.235 7.315 87.405 7.485 ;
        RECT 87.605 7.315 87.775 7.485 ;
        RECT 87.975 7.315 88.145 7.485 ;
        RECT 88.345 7.315 88.515 7.485 ;
        RECT 88.715 7.315 88.885 7.485 ;
        RECT 89.085 7.315 89.255 7.485 ;
        RECT 89.455 7.315 89.625 7.485 ;
        RECT 90.195 7.315 90.365 7.485 ;
        RECT 90.565 7.315 90.735 7.485 ;
        RECT 90.935 7.315 91.105 7.485 ;
        RECT 91.305 7.315 91.475 7.485 ;
        RECT 91.675 7.315 91.845 7.485 ;
        RECT 92.045 7.315 92.215 7.485 ;
        RECT 92.415 7.315 92.585 7.485 ;
        RECT 92.785 7.315 92.955 7.485 ;
        RECT 93.525 7.315 93.695 7.485 ;
        RECT 93.895 7.315 94.065 7.485 ;
        RECT 94.265 7.315 94.435 7.485 ;
        RECT 94.635 7.315 94.805 7.485 ;
        RECT 95.005 7.315 95.175 7.485 ;
        RECT 95.375 7.315 95.545 7.485 ;
        RECT 95.745 7.315 95.915 7.485 ;
        RECT 96.115 7.315 96.285 7.485 ;
        RECT 96.855 7.315 97.025 7.485 ;
        RECT 97.225 7.315 97.395 7.485 ;
        RECT 97.595 7.315 97.765 7.485 ;
        RECT 97.965 7.315 98.135 7.485 ;
        RECT 98.335 7.315 98.505 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 98.960 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 98.960 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.610 0.170 10.780 1.130 ;
        RECT 14.260 0.170 14.600 2.720 ;
        RECT 15.420 0.170 15.590 1.130 ;
        RECT 19.070 0.170 19.410 2.720 ;
        RECT 20.230 0.170 20.400 1.130 ;
        RECT 23.880 0.170 24.220 2.720 ;
        RECT 25.040 0.170 25.210 1.130 ;
        RECT 28.690 0.170 29.030 2.720 ;
        RECT 29.850 0.170 30.020 1.130 ;
        RECT 33.500 0.170 33.840 2.720 ;
        RECT 34.660 0.170 34.830 1.130 ;
        RECT 38.310 0.170 38.650 2.720 ;
        RECT 39.470 0.170 39.640 1.130 ;
        RECT 43.120 0.170 43.460 2.720 ;
        RECT 44.280 0.170 44.450 1.130 ;
        RECT 47.930 0.170 48.270 2.720 ;
        RECT 49.090 0.170 49.260 1.130 ;
        RECT 52.740 0.170 53.080 2.720 ;
        RECT 53.900 0.170 54.070 1.130 ;
        RECT 57.550 0.170 57.890 2.720 ;
        RECT 58.710 0.170 58.880 1.130 ;
        RECT 62.360 0.170 62.700 2.720 ;
        RECT 63.520 0.170 63.690 1.130 ;
        RECT 67.170 0.170 67.510 2.720 ;
        RECT 68.330 0.170 68.500 1.130 ;
        RECT 71.980 0.170 72.320 2.720 ;
        RECT 73.140 0.170 73.310 1.130 ;
        RECT 76.790 0.170 77.130 2.720 ;
        RECT 77.950 0.170 78.120 1.130 ;
        RECT 81.600 0.170 81.940 2.720 ;
        RECT 82.760 0.170 82.930 1.130 ;
        RECT 86.410 0.170 86.750 2.720 ;
        RECT 87.675 0.170 87.845 1.120 ;
        RECT 89.740 0.170 90.080 2.720 ;
        RECT 91.005 0.170 91.175 1.120 ;
        RECT 93.070 0.170 93.410 2.720 ;
        RECT 94.335 0.170 94.505 1.120 ;
        RECT 96.400 0.170 96.740 2.720 ;
        RECT 97.115 0.620 97.285 1.750 ;
        RECT 98.085 0.620 98.255 1.750 ;
        RECT 97.115 0.450 98.255 0.620 ;
        RECT 97.115 0.170 97.285 0.450 ;
        RECT 97.600 0.170 97.770 0.450 ;
        RECT 98.085 0.170 98.255 0.450 ;
        RECT 98.620 0.170 98.960 2.720 ;
        RECT -0.170 -0.170 98.960 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.515 -0.085 29.685 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.625 -0.085 30.795 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 32.845 -0.085 33.015 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.435 -0.085 35.605 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.175 -0.085 36.345 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.765 -0.085 38.935 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.505 -0.085 39.675 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.615 -0.085 40.785 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 42.835 -0.085 43.005 0.085 ;
        RECT 43.575 -0.085 43.745 0.085 ;
        RECT 43.945 -0.085 44.115 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 47.645 -0.085 47.815 0.085 ;
        RECT 48.385 -0.085 48.555 0.085 ;
        RECT 48.755 -0.085 48.925 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 50.975 -0.085 51.145 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 51.715 -0.085 51.885 0.085 ;
        RECT 52.085 -0.085 52.255 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.305 -0.085 54.475 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.525 -0.085 56.695 0.085 ;
        RECT 56.895 -0.085 57.065 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 60.965 -0.085 61.135 0.085 ;
        RECT 61.335 -0.085 61.505 0.085 ;
        RECT 61.705 -0.085 61.875 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.295 -0.085 64.465 0.085 ;
        RECT 64.665 -0.085 64.835 0.085 ;
        RECT 65.035 -0.085 65.205 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.625 -0.085 67.795 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.365 -0.085 68.535 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.475 -0.085 69.645 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 70.955 -0.085 71.125 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.175 -0.085 73.345 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
        RECT 74.285 -0.085 74.455 0.085 ;
        RECT 74.655 -0.085 74.825 0.085 ;
        RECT 75.025 -0.085 75.195 0.085 ;
        RECT 75.395 -0.085 75.565 0.085 ;
        RECT 75.765 -0.085 75.935 0.085 ;
        RECT 76.135 -0.085 76.305 0.085 ;
        RECT 76.505 -0.085 76.675 0.085 ;
        RECT 77.245 -0.085 77.415 0.085 ;
        RECT 77.615 -0.085 77.785 0.085 ;
        RECT 77.985 -0.085 78.155 0.085 ;
        RECT 78.355 -0.085 78.525 0.085 ;
        RECT 78.725 -0.085 78.895 0.085 ;
        RECT 79.095 -0.085 79.265 0.085 ;
        RECT 79.465 -0.085 79.635 0.085 ;
        RECT 79.835 -0.085 80.005 0.085 ;
        RECT 80.205 -0.085 80.375 0.085 ;
        RECT 80.575 -0.085 80.745 0.085 ;
        RECT 80.945 -0.085 81.115 0.085 ;
        RECT 81.315 -0.085 81.485 0.085 ;
        RECT 82.055 -0.085 82.225 0.085 ;
        RECT 82.425 -0.085 82.595 0.085 ;
        RECT 82.795 -0.085 82.965 0.085 ;
        RECT 83.165 -0.085 83.335 0.085 ;
        RECT 83.535 -0.085 83.705 0.085 ;
        RECT 83.905 -0.085 84.075 0.085 ;
        RECT 84.275 -0.085 84.445 0.085 ;
        RECT 84.645 -0.085 84.815 0.085 ;
        RECT 85.015 -0.085 85.185 0.085 ;
        RECT 85.385 -0.085 85.555 0.085 ;
        RECT 85.755 -0.085 85.925 0.085 ;
        RECT 86.125 -0.085 86.295 0.085 ;
        RECT 86.865 -0.085 87.035 0.085 ;
        RECT 87.235 -0.085 87.405 0.085 ;
        RECT 87.605 -0.085 87.775 0.085 ;
        RECT 87.975 -0.085 88.145 0.085 ;
        RECT 88.345 -0.085 88.515 0.085 ;
        RECT 88.715 -0.085 88.885 0.085 ;
        RECT 89.085 -0.085 89.255 0.085 ;
        RECT 89.455 -0.085 89.625 0.085 ;
        RECT 90.195 -0.085 90.365 0.085 ;
        RECT 90.565 -0.085 90.735 0.085 ;
        RECT 90.935 -0.085 91.105 0.085 ;
        RECT 91.305 -0.085 91.475 0.085 ;
        RECT 91.675 -0.085 91.845 0.085 ;
        RECT 92.045 -0.085 92.215 0.085 ;
        RECT 92.415 -0.085 92.585 0.085 ;
        RECT 92.785 -0.085 92.955 0.085 ;
        RECT 93.525 -0.085 93.695 0.085 ;
        RECT 93.895 -0.085 94.065 0.085 ;
        RECT 94.265 -0.085 94.435 0.085 ;
        RECT 94.635 -0.085 94.805 0.085 ;
        RECT 95.005 -0.085 95.175 0.085 ;
        RECT 95.375 -0.085 95.545 0.085 ;
        RECT 95.745 -0.085 95.915 0.085 ;
        RECT 96.115 -0.085 96.285 0.085 ;
        RECT 96.855 -0.085 97.025 0.085 ;
        RECT 97.225 -0.085 97.395 0.085 ;
        RECT 97.595 -0.085 97.765 0.085 ;
        RECT 97.965 -0.085 98.135 0.085 ;
        RECT 98.335 -0.085 98.505 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 98.960 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 11.065 5.240 11.235 7.020 ;
        RECT 11.945 5.240 12.115 7.020 ;
        RECT 12.825 5.240 12.995 7.020 ;
        RECT 15.875 5.240 16.045 7.020 ;
        RECT 16.755 5.240 16.925 7.020 ;
        RECT 17.635 5.240 17.805 7.020 ;
        RECT 20.685 5.240 20.855 7.020 ;
        RECT 21.565 5.240 21.735 7.020 ;
        RECT 22.445 5.240 22.615 7.020 ;
        RECT 25.495 5.240 25.665 7.020 ;
        RECT 26.375 5.240 26.545 7.020 ;
        RECT 27.255 5.240 27.425 7.020 ;
        RECT 30.305 5.240 30.475 7.020 ;
        RECT 31.185 5.240 31.355 7.020 ;
        RECT 32.065 5.240 32.235 7.020 ;
        RECT 35.115 5.240 35.285 7.020 ;
        RECT 35.995 5.240 36.165 7.020 ;
        RECT 36.875 5.240 37.045 7.020 ;
        RECT 39.925 5.240 40.095 7.020 ;
        RECT 40.805 5.240 40.975 7.020 ;
        RECT 41.685 5.240 41.855 7.020 ;
        RECT 44.735 5.240 44.905 7.020 ;
        RECT 45.615 5.240 45.785 7.020 ;
        RECT 46.495 5.240 46.665 7.020 ;
        RECT 49.545 5.240 49.715 7.020 ;
        RECT 50.425 5.240 50.595 7.020 ;
        RECT 51.305 5.240 51.475 7.020 ;
        RECT 54.355 5.240 54.525 7.020 ;
        RECT 55.235 5.240 55.405 7.020 ;
        RECT 56.115 5.240 56.285 7.020 ;
        RECT 59.165 5.240 59.335 7.020 ;
        RECT 60.045 5.240 60.215 7.020 ;
        RECT 60.925 5.240 61.095 7.020 ;
        RECT 63.975 5.240 64.145 7.020 ;
        RECT 64.855 5.240 65.025 7.020 ;
        RECT 65.735 5.240 65.905 7.020 ;
        RECT 68.785 5.240 68.955 7.020 ;
        RECT 69.665 5.240 69.835 7.020 ;
        RECT 70.545 5.240 70.715 7.020 ;
        RECT 73.595 5.240 73.765 7.020 ;
        RECT 74.475 5.240 74.645 7.020 ;
        RECT 75.355 5.240 75.525 7.020 ;
        RECT 78.405 5.240 78.575 7.020 ;
        RECT 79.285 5.240 79.455 7.020 ;
        RECT 80.165 5.240 80.335 7.020 ;
        RECT 83.215 5.240 83.385 7.020 ;
        RECT 84.095 5.240 84.265 7.020 ;
        RECT 84.975 5.240 85.145 7.020 ;
        RECT 87.725 6.825 87.905 6.995 ;
        RECT 87.725 5.295 87.895 6.825 ;
        RECT 88.605 5.295 88.775 6.995 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 11.065 5.070 13.775 5.240 ;
        RECT 15.875 5.070 18.585 5.240 ;
        RECT 20.685 5.070 23.395 5.240 ;
        RECT 25.495 5.070 28.205 5.240 ;
        RECT 30.305 5.070 33.015 5.240 ;
        RECT 35.115 5.070 37.825 5.240 ;
        RECT 39.925 5.070 42.635 5.240 ;
        RECT 44.735 5.070 47.445 5.240 ;
        RECT 49.545 5.070 52.255 5.240 ;
        RECT 54.355 5.070 57.065 5.240 ;
        RECT 59.165 5.070 61.875 5.240 ;
        RECT 63.975 5.070 66.685 5.240 ;
        RECT 68.785 5.070 71.495 5.240 ;
        RECT 73.595 5.070 76.305 5.240 ;
        RECT 78.405 5.070 81.115 5.240 ;
        RECT 83.215 5.070 85.925 5.240 ;
        RECT 87.725 5.125 88.775 5.295 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 8.055 1.915 8.225 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 12.865 1.915 13.035 4.865 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.125 1.675 10.295 1.755 ;
        RECT 11.095 1.675 11.265 1.755 ;
        RECT 12.065 1.675 12.235 1.755 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.125 1.505 12.235 1.675 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.125 0.375 10.295 1.505 ;
        RECT 11.095 0.625 11.265 1.505 ;
        RECT 12.065 1.425 12.235 1.505 ;
        RECT 11.585 1.080 11.755 1.160 ;
        RECT 12.635 1.080 12.805 1.755 ;
        RECT 13.605 1.750 13.775 5.070 ;
        RECT 15.455 1.915 15.625 4.865 ;
        RECT 11.585 0.910 12.805 1.080 ;
        RECT 11.585 0.830 11.755 0.910 ;
        RECT 12.065 0.625 12.235 0.705 ;
        RECT 11.095 0.455 12.235 0.625 ;
        RECT 11.095 0.375 11.265 0.455 ;
        RECT 12.065 0.375 12.235 0.455 ;
        RECT 12.635 0.625 12.805 0.910 ;
        RECT 13.120 1.580 13.775 1.750 ;
        RECT 14.935 1.675 15.105 1.755 ;
        RECT 15.905 1.675 16.075 1.755 ;
        RECT 16.875 1.675 17.045 1.755 ;
        RECT 13.120 0.845 13.290 1.580 ;
        RECT 14.935 1.505 17.045 1.675 ;
        RECT 13.605 0.625 13.775 1.395 ;
        RECT 12.635 0.455 13.775 0.625 ;
        RECT 12.635 0.375 12.805 0.455 ;
        RECT 13.605 0.375 13.775 0.455 ;
        RECT 14.935 0.375 15.105 1.505 ;
        RECT 15.905 0.625 16.075 1.505 ;
        RECT 16.875 1.425 17.045 1.505 ;
        RECT 16.395 1.080 16.565 1.160 ;
        RECT 17.445 1.080 17.615 1.755 ;
        RECT 18.415 1.750 18.585 5.070 ;
        RECT 20.265 1.915 20.435 4.865 ;
        RECT 22.485 1.915 22.655 4.865 ;
        RECT 16.395 0.910 17.615 1.080 ;
        RECT 16.395 0.830 16.565 0.910 ;
        RECT 16.875 0.625 17.045 0.705 ;
        RECT 15.905 0.455 17.045 0.625 ;
        RECT 15.905 0.375 16.075 0.455 ;
        RECT 16.875 0.375 17.045 0.455 ;
        RECT 17.445 0.625 17.615 0.910 ;
        RECT 17.930 1.580 18.585 1.750 ;
        RECT 19.745 1.675 19.915 1.755 ;
        RECT 20.715 1.675 20.885 1.755 ;
        RECT 21.685 1.675 21.855 1.755 ;
        RECT 17.930 0.845 18.100 1.580 ;
        RECT 19.745 1.505 21.855 1.675 ;
        RECT 18.415 0.625 18.585 1.395 ;
        RECT 17.445 0.455 18.585 0.625 ;
        RECT 17.445 0.375 17.615 0.455 ;
        RECT 18.415 0.375 18.585 0.455 ;
        RECT 19.745 0.375 19.915 1.505 ;
        RECT 20.715 0.625 20.885 1.505 ;
        RECT 21.685 1.425 21.855 1.505 ;
        RECT 21.205 1.080 21.375 1.160 ;
        RECT 22.255 1.080 22.425 1.755 ;
        RECT 23.225 1.750 23.395 5.070 ;
        RECT 25.075 1.915 25.245 4.865 ;
        RECT 27.295 1.915 27.465 4.865 ;
        RECT 21.205 0.910 22.425 1.080 ;
        RECT 21.205 0.830 21.375 0.910 ;
        RECT 21.685 0.625 21.855 0.705 ;
        RECT 20.715 0.455 21.855 0.625 ;
        RECT 20.715 0.375 20.885 0.455 ;
        RECT 21.685 0.375 21.855 0.455 ;
        RECT 22.255 0.625 22.425 0.910 ;
        RECT 22.740 1.580 23.395 1.750 ;
        RECT 24.555 1.675 24.725 1.755 ;
        RECT 25.525 1.675 25.695 1.755 ;
        RECT 26.495 1.675 26.665 1.755 ;
        RECT 22.740 0.845 22.910 1.580 ;
        RECT 24.555 1.505 26.665 1.675 ;
        RECT 23.225 0.625 23.395 1.395 ;
        RECT 22.255 0.455 23.395 0.625 ;
        RECT 22.255 0.375 22.425 0.455 ;
        RECT 23.225 0.375 23.395 0.455 ;
        RECT 24.555 0.375 24.725 1.505 ;
        RECT 25.525 0.625 25.695 1.505 ;
        RECT 26.495 1.425 26.665 1.505 ;
        RECT 26.015 1.080 26.185 1.160 ;
        RECT 27.065 1.080 27.235 1.755 ;
        RECT 28.035 1.750 28.205 5.070 ;
        RECT 32.105 1.915 32.275 4.865 ;
        RECT 26.015 0.910 27.235 1.080 ;
        RECT 26.015 0.830 26.185 0.910 ;
        RECT 26.495 0.625 26.665 0.705 ;
        RECT 25.525 0.455 26.665 0.625 ;
        RECT 25.525 0.375 25.695 0.455 ;
        RECT 26.495 0.375 26.665 0.455 ;
        RECT 27.065 0.625 27.235 0.910 ;
        RECT 27.550 1.580 28.205 1.750 ;
        RECT 29.365 1.675 29.535 1.755 ;
        RECT 30.335 1.675 30.505 1.755 ;
        RECT 31.305 1.675 31.475 1.755 ;
        RECT 27.550 0.845 27.720 1.580 ;
        RECT 29.365 1.505 31.475 1.675 ;
        RECT 28.035 0.625 28.205 1.395 ;
        RECT 27.065 0.455 28.205 0.625 ;
        RECT 27.065 0.375 27.235 0.455 ;
        RECT 28.035 0.375 28.205 0.455 ;
        RECT 29.365 0.375 29.535 1.505 ;
        RECT 30.335 0.625 30.505 1.505 ;
        RECT 31.305 1.425 31.475 1.505 ;
        RECT 30.825 1.080 30.995 1.160 ;
        RECT 31.875 1.080 32.045 1.755 ;
        RECT 32.845 1.750 33.015 5.070 ;
        RECT 34.695 1.915 34.865 4.865 ;
        RECT 36.915 1.915 37.085 4.865 ;
        RECT 30.825 0.910 32.045 1.080 ;
        RECT 30.825 0.830 30.995 0.910 ;
        RECT 31.305 0.625 31.475 0.705 ;
        RECT 30.335 0.455 31.475 0.625 ;
        RECT 30.335 0.375 30.505 0.455 ;
        RECT 31.305 0.375 31.475 0.455 ;
        RECT 31.875 0.625 32.045 0.910 ;
        RECT 32.360 1.580 33.015 1.750 ;
        RECT 34.175 1.675 34.345 1.755 ;
        RECT 35.145 1.675 35.315 1.755 ;
        RECT 36.115 1.675 36.285 1.755 ;
        RECT 32.360 0.845 32.530 1.580 ;
        RECT 34.175 1.505 36.285 1.675 ;
        RECT 32.845 0.625 33.015 1.395 ;
        RECT 31.875 0.455 33.015 0.625 ;
        RECT 31.875 0.375 32.045 0.455 ;
        RECT 32.845 0.375 33.015 0.455 ;
        RECT 34.175 0.375 34.345 1.505 ;
        RECT 35.145 0.625 35.315 1.505 ;
        RECT 36.115 1.425 36.285 1.505 ;
        RECT 35.635 1.080 35.805 1.160 ;
        RECT 36.685 1.080 36.855 1.755 ;
        RECT 37.655 1.750 37.825 5.070 ;
        RECT 39.505 1.915 39.675 4.865 ;
        RECT 41.725 1.915 41.895 4.865 ;
        RECT 35.635 0.910 36.855 1.080 ;
        RECT 35.635 0.830 35.805 0.910 ;
        RECT 36.115 0.625 36.285 0.705 ;
        RECT 35.145 0.455 36.285 0.625 ;
        RECT 35.145 0.375 35.315 0.455 ;
        RECT 36.115 0.375 36.285 0.455 ;
        RECT 36.685 0.625 36.855 0.910 ;
        RECT 37.170 1.580 37.825 1.750 ;
        RECT 38.985 1.675 39.155 1.755 ;
        RECT 39.955 1.675 40.125 1.755 ;
        RECT 40.925 1.675 41.095 1.755 ;
        RECT 37.170 0.845 37.340 1.580 ;
        RECT 38.985 1.505 41.095 1.675 ;
        RECT 37.655 0.625 37.825 1.395 ;
        RECT 36.685 0.455 37.825 0.625 ;
        RECT 36.685 0.375 36.855 0.455 ;
        RECT 37.655 0.375 37.825 0.455 ;
        RECT 38.985 0.375 39.155 1.505 ;
        RECT 39.955 0.625 40.125 1.505 ;
        RECT 40.925 1.425 41.095 1.505 ;
        RECT 40.445 1.080 40.615 1.160 ;
        RECT 41.495 1.080 41.665 1.755 ;
        RECT 42.465 1.750 42.635 5.070 ;
        RECT 44.315 1.915 44.485 4.865 ;
        RECT 40.445 0.910 41.665 1.080 ;
        RECT 40.445 0.830 40.615 0.910 ;
        RECT 40.925 0.625 41.095 0.705 ;
        RECT 39.955 0.455 41.095 0.625 ;
        RECT 39.955 0.375 40.125 0.455 ;
        RECT 40.925 0.375 41.095 0.455 ;
        RECT 41.495 0.625 41.665 0.910 ;
        RECT 41.980 1.580 42.635 1.750 ;
        RECT 43.795 1.675 43.965 1.755 ;
        RECT 44.765 1.675 44.935 1.755 ;
        RECT 45.735 1.675 45.905 1.755 ;
        RECT 41.980 0.845 42.150 1.580 ;
        RECT 43.795 1.505 45.905 1.675 ;
        RECT 42.465 0.625 42.635 1.395 ;
        RECT 41.495 0.455 42.635 0.625 ;
        RECT 41.495 0.375 41.665 0.455 ;
        RECT 42.465 0.375 42.635 0.455 ;
        RECT 43.795 0.375 43.965 1.505 ;
        RECT 44.765 0.625 44.935 1.505 ;
        RECT 45.735 1.425 45.905 1.505 ;
        RECT 45.255 1.080 45.425 1.160 ;
        RECT 46.305 1.080 46.475 1.755 ;
        RECT 47.275 1.750 47.445 5.070 ;
        RECT 49.125 1.915 49.295 4.865 ;
        RECT 51.345 1.915 51.515 4.865 ;
        RECT 45.255 0.910 46.475 1.080 ;
        RECT 45.255 0.830 45.425 0.910 ;
        RECT 45.735 0.625 45.905 0.705 ;
        RECT 44.765 0.455 45.905 0.625 ;
        RECT 44.765 0.375 44.935 0.455 ;
        RECT 45.735 0.375 45.905 0.455 ;
        RECT 46.305 0.625 46.475 0.910 ;
        RECT 46.790 1.580 47.445 1.750 ;
        RECT 48.605 1.675 48.775 1.755 ;
        RECT 49.575 1.675 49.745 1.755 ;
        RECT 50.545 1.675 50.715 1.755 ;
        RECT 46.790 0.845 46.960 1.580 ;
        RECT 48.605 1.505 50.715 1.675 ;
        RECT 47.275 0.625 47.445 1.395 ;
        RECT 46.305 0.455 47.445 0.625 ;
        RECT 46.305 0.375 46.475 0.455 ;
        RECT 47.275 0.375 47.445 0.455 ;
        RECT 48.605 0.375 48.775 1.505 ;
        RECT 49.575 0.625 49.745 1.505 ;
        RECT 50.545 1.425 50.715 1.505 ;
        RECT 50.065 1.080 50.235 1.160 ;
        RECT 51.115 1.080 51.285 1.755 ;
        RECT 52.085 1.750 52.255 5.070 ;
        RECT 53.935 1.915 54.105 4.865 ;
        RECT 56.155 1.915 56.325 4.865 ;
        RECT 50.065 0.910 51.285 1.080 ;
        RECT 50.065 0.830 50.235 0.910 ;
        RECT 50.545 0.625 50.715 0.705 ;
        RECT 49.575 0.455 50.715 0.625 ;
        RECT 49.575 0.375 49.745 0.455 ;
        RECT 50.545 0.375 50.715 0.455 ;
        RECT 51.115 0.625 51.285 0.910 ;
        RECT 51.600 1.580 52.255 1.750 ;
        RECT 53.415 1.675 53.585 1.755 ;
        RECT 54.385 1.675 54.555 1.755 ;
        RECT 55.355 1.675 55.525 1.755 ;
        RECT 51.600 0.845 51.770 1.580 ;
        RECT 53.415 1.505 55.525 1.675 ;
        RECT 52.085 0.625 52.255 1.395 ;
        RECT 51.115 0.455 52.255 0.625 ;
        RECT 51.115 0.375 51.285 0.455 ;
        RECT 52.085 0.375 52.255 0.455 ;
        RECT 53.415 0.375 53.585 1.505 ;
        RECT 54.385 0.625 54.555 1.505 ;
        RECT 55.355 1.425 55.525 1.505 ;
        RECT 54.875 1.080 55.045 1.160 ;
        RECT 55.925 1.080 56.095 1.755 ;
        RECT 56.895 1.750 57.065 5.070 ;
        RECT 60.965 1.915 61.135 4.865 ;
        RECT 54.875 0.910 56.095 1.080 ;
        RECT 54.875 0.830 55.045 0.910 ;
        RECT 55.355 0.625 55.525 0.705 ;
        RECT 54.385 0.455 55.525 0.625 ;
        RECT 54.385 0.375 54.555 0.455 ;
        RECT 55.355 0.375 55.525 0.455 ;
        RECT 55.925 0.625 56.095 0.910 ;
        RECT 56.410 1.580 57.065 1.750 ;
        RECT 58.225 1.675 58.395 1.755 ;
        RECT 59.195 1.675 59.365 1.755 ;
        RECT 60.165 1.675 60.335 1.755 ;
        RECT 56.410 0.845 56.580 1.580 ;
        RECT 58.225 1.505 60.335 1.675 ;
        RECT 56.895 0.625 57.065 1.395 ;
        RECT 55.925 0.455 57.065 0.625 ;
        RECT 55.925 0.375 56.095 0.455 ;
        RECT 56.895 0.375 57.065 0.455 ;
        RECT 58.225 0.375 58.395 1.505 ;
        RECT 59.195 0.625 59.365 1.505 ;
        RECT 60.165 1.425 60.335 1.505 ;
        RECT 59.685 1.080 59.855 1.160 ;
        RECT 60.735 1.080 60.905 1.755 ;
        RECT 61.705 1.750 61.875 5.070 ;
        RECT 63.555 1.915 63.725 4.865 ;
        RECT 65.775 1.915 65.945 4.865 ;
        RECT 59.685 0.910 60.905 1.080 ;
        RECT 59.685 0.830 59.855 0.910 ;
        RECT 60.165 0.625 60.335 0.705 ;
        RECT 59.195 0.455 60.335 0.625 ;
        RECT 59.195 0.375 59.365 0.455 ;
        RECT 60.165 0.375 60.335 0.455 ;
        RECT 60.735 0.625 60.905 0.910 ;
        RECT 61.220 1.580 61.875 1.750 ;
        RECT 63.035 1.675 63.205 1.755 ;
        RECT 64.005 1.675 64.175 1.755 ;
        RECT 64.975 1.675 65.145 1.755 ;
        RECT 61.220 0.845 61.390 1.580 ;
        RECT 63.035 1.505 65.145 1.675 ;
        RECT 61.705 0.625 61.875 1.395 ;
        RECT 60.735 0.455 61.875 0.625 ;
        RECT 60.735 0.375 60.905 0.455 ;
        RECT 61.705 0.375 61.875 0.455 ;
        RECT 63.035 0.375 63.205 1.505 ;
        RECT 64.005 0.625 64.175 1.505 ;
        RECT 64.975 1.425 65.145 1.505 ;
        RECT 64.495 1.080 64.665 1.160 ;
        RECT 65.545 1.080 65.715 1.755 ;
        RECT 66.515 1.750 66.685 5.070 ;
        RECT 68.365 1.915 68.535 4.865 ;
        RECT 70.585 1.915 70.755 4.865 ;
        RECT 64.495 0.910 65.715 1.080 ;
        RECT 64.495 0.830 64.665 0.910 ;
        RECT 64.975 0.625 65.145 0.705 ;
        RECT 64.005 0.455 65.145 0.625 ;
        RECT 64.005 0.375 64.175 0.455 ;
        RECT 64.975 0.375 65.145 0.455 ;
        RECT 65.545 0.625 65.715 0.910 ;
        RECT 66.030 1.580 66.685 1.750 ;
        RECT 67.845 1.675 68.015 1.755 ;
        RECT 68.815 1.675 68.985 1.755 ;
        RECT 69.785 1.675 69.955 1.755 ;
        RECT 66.030 0.845 66.200 1.580 ;
        RECT 67.845 1.505 69.955 1.675 ;
        RECT 66.515 0.625 66.685 1.395 ;
        RECT 65.545 0.455 66.685 0.625 ;
        RECT 65.545 0.375 65.715 0.455 ;
        RECT 66.515 0.375 66.685 0.455 ;
        RECT 67.845 0.375 68.015 1.505 ;
        RECT 68.815 0.625 68.985 1.505 ;
        RECT 69.785 1.425 69.955 1.505 ;
        RECT 69.305 1.080 69.475 1.160 ;
        RECT 70.355 1.080 70.525 1.755 ;
        RECT 71.325 1.750 71.495 5.070 ;
        RECT 73.175 1.915 73.345 4.865 ;
        RECT 69.305 0.910 70.525 1.080 ;
        RECT 69.305 0.830 69.475 0.910 ;
        RECT 69.785 0.625 69.955 0.705 ;
        RECT 68.815 0.455 69.955 0.625 ;
        RECT 68.815 0.375 68.985 0.455 ;
        RECT 69.785 0.375 69.955 0.455 ;
        RECT 70.355 0.625 70.525 0.910 ;
        RECT 70.840 1.580 71.495 1.750 ;
        RECT 72.655 1.675 72.825 1.755 ;
        RECT 73.625 1.675 73.795 1.755 ;
        RECT 74.595 1.675 74.765 1.755 ;
        RECT 70.840 0.845 71.010 1.580 ;
        RECT 72.655 1.505 74.765 1.675 ;
        RECT 71.325 0.625 71.495 1.395 ;
        RECT 70.355 0.455 71.495 0.625 ;
        RECT 70.355 0.375 70.525 0.455 ;
        RECT 71.325 0.375 71.495 0.455 ;
        RECT 72.655 0.375 72.825 1.505 ;
        RECT 73.625 0.625 73.795 1.505 ;
        RECT 74.595 1.425 74.765 1.505 ;
        RECT 74.115 1.080 74.285 1.160 ;
        RECT 75.165 1.080 75.335 1.755 ;
        RECT 76.135 1.750 76.305 5.070 ;
        RECT 77.985 1.915 78.155 4.865 ;
        RECT 80.205 1.915 80.375 4.865 ;
        RECT 74.115 0.910 75.335 1.080 ;
        RECT 74.115 0.830 74.285 0.910 ;
        RECT 74.595 0.625 74.765 0.705 ;
        RECT 73.625 0.455 74.765 0.625 ;
        RECT 73.625 0.375 73.795 0.455 ;
        RECT 74.595 0.375 74.765 0.455 ;
        RECT 75.165 0.625 75.335 0.910 ;
        RECT 75.650 1.580 76.305 1.750 ;
        RECT 77.465 1.675 77.635 1.755 ;
        RECT 78.435 1.675 78.605 1.755 ;
        RECT 79.405 1.675 79.575 1.755 ;
        RECT 75.650 0.845 75.820 1.580 ;
        RECT 77.465 1.505 79.575 1.675 ;
        RECT 76.135 0.625 76.305 1.395 ;
        RECT 75.165 0.455 76.305 0.625 ;
        RECT 75.165 0.375 75.335 0.455 ;
        RECT 76.135 0.375 76.305 0.455 ;
        RECT 77.465 0.375 77.635 1.505 ;
        RECT 78.435 0.625 78.605 1.505 ;
        RECT 79.405 1.425 79.575 1.505 ;
        RECT 78.925 1.080 79.095 1.160 ;
        RECT 79.975 1.080 80.145 1.755 ;
        RECT 80.945 1.750 81.115 5.070 ;
        RECT 82.795 1.915 82.965 4.865 ;
        RECT 85.015 1.915 85.185 4.865 ;
        RECT 78.925 0.910 80.145 1.080 ;
        RECT 78.925 0.830 79.095 0.910 ;
        RECT 79.405 0.625 79.575 0.705 ;
        RECT 78.435 0.455 79.575 0.625 ;
        RECT 78.435 0.375 78.605 0.455 ;
        RECT 79.405 0.375 79.575 0.455 ;
        RECT 79.975 0.625 80.145 0.910 ;
        RECT 80.460 1.580 81.115 1.750 ;
        RECT 82.275 1.675 82.445 1.755 ;
        RECT 83.245 1.675 83.415 1.755 ;
        RECT 84.215 1.675 84.385 1.755 ;
        RECT 80.460 0.845 80.630 1.580 ;
        RECT 82.275 1.505 84.385 1.675 ;
        RECT 80.945 0.625 81.115 1.395 ;
        RECT 79.975 0.455 81.115 0.625 ;
        RECT 79.975 0.375 80.145 0.455 ;
        RECT 80.945 0.375 81.115 0.455 ;
        RECT 82.275 0.375 82.445 1.505 ;
        RECT 83.245 0.625 83.415 1.505 ;
        RECT 84.215 1.425 84.385 1.505 ;
        RECT 83.735 1.080 83.905 1.160 ;
        RECT 84.785 1.080 84.955 1.755 ;
        RECT 85.755 1.750 85.925 5.070 ;
        RECT 88.605 5.045 88.775 5.125 ;
        RECT 90.605 6.825 92.535 6.995 ;
        RECT 90.605 5.045 90.775 6.825 ;
        RECT 91.045 5.295 91.215 6.565 ;
        RECT 91.485 5.555 91.655 6.825 ;
        RECT 91.925 5.295 92.095 6.565 ;
        RECT 92.365 5.375 92.535 6.825 ;
        RECT 93.945 6.825 95.875 6.995 ;
        RECT 91.045 5.125 92.095 5.295 ;
        RECT 91.925 5.045 92.095 5.125 ;
        RECT 93.945 5.045 94.115 6.825 ;
        RECT 94.385 5.295 94.555 6.565 ;
        RECT 94.825 5.555 94.995 6.825 ;
        RECT 95.265 5.295 95.435 6.565 ;
        RECT 95.705 5.555 95.875 6.825 ;
        RECT 94.385 5.125 95.915 5.295 ;
        RECT 87.235 1.915 87.405 4.870 ;
        RECT 88.385 4.710 88.555 4.870 ;
        RECT 88.345 4.540 88.555 4.710 ;
        RECT 88.345 1.915 88.515 4.540 ;
        RECT 90.935 1.915 91.105 4.870 ;
        RECT 92.415 1.915 92.585 4.870 ;
        RECT 93.895 1.915 94.065 4.870 ;
        RECT 95.005 4.540 95.195 4.870 ;
        RECT 95.005 1.915 95.175 4.540 ;
        RECT 83.735 0.910 84.955 1.080 ;
        RECT 83.735 0.830 83.905 0.910 ;
        RECT 84.215 0.625 84.385 0.705 ;
        RECT 83.245 0.455 84.385 0.625 ;
        RECT 83.245 0.375 83.415 0.455 ;
        RECT 84.215 0.375 84.385 0.455 ;
        RECT 84.785 0.625 84.955 0.910 ;
        RECT 85.270 1.580 85.925 1.750 ;
        RECT 87.190 1.665 87.360 1.745 ;
        RECT 88.160 1.665 88.330 1.745 ;
        RECT 85.270 0.845 85.440 1.580 ;
        RECT 87.190 1.495 88.330 1.665 ;
        RECT 85.755 0.625 85.925 1.395 ;
        RECT 84.785 0.455 85.925 0.625 ;
        RECT 84.785 0.375 84.955 0.455 ;
        RECT 85.755 0.375 85.925 0.455 ;
        RECT 87.190 0.365 87.360 1.495 ;
        RECT 88.160 0.615 88.330 1.495 ;
        RECT 88.645 1.170 88.815 1.345 ;
        RECT 88.640 1.015 88.815 1.170 ;
        RECT 88.640 0.835 88.810 1.015 ;
        RECT 89.130 0.615 89.300 1.745 ;
        RECT 88.160 0.445 89.300 0.615 ;
        RECT 88.160 0.365 88.330 0.445 ;
        RECT 89.130 0.365 89.300 0.445 ;
        RECT 90.520 1.665 90.690 1.745 ;
        RECT 91.490 1.665 91.660 1.745 ;
        RECT 90.520 1.495 91.660 1.665 ;
        RECT 90.520 0.365 90.690 1.495 ;
        RECT 91.490 0.615 91.660 1.495 ;
        RECT 91.975 0.835 92.145 1.345 ;
        RECT 92.460 0.615 92.630 1.745 ;
        RECT 91.490 0.445 92.630 0.615 ;
        RECT 91.490 0.365 91.660 0.445 ;
        RECT 92.460 0.365 92.630 0.445 ;
        RECT 93.850 1.665 94.020 1.745 ;
        RECT 94.820 1.665 94.990 1.745 ;
        RECT 95.745 1.730 95.915 5.125 ;
        RECT 97.225 1.920 97.395 4.865 ;
        RECT 93.850 1.495 94.990 1.665 ;
        RECT 93.850 0.365 94.020 1.495 ;
        RECT 94.820 0.615 94.990 1.495 ;
        RECT 95.305 1.560 95.915 1.730 ;
        RECT 95.305 0.835 95.475 1.560 ;
        RECT 95.790 0.615 95.960 1.390 ;
        RECT 94.820 0.445 95.960 0.615 ;
        RECT 94.820 0.365 94.990 0.445 ;
        RECT 95.790 0.365 95.960 0.445 ;
      LAYER mcon ;
        RECT 88.605 5.125 88.775 5.295 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 2.505 4.155 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 8.055 3.615 8.225 3.785 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 10.645 2.505 10.815 2.675 ;
        RECT 12.865 3.615 13.035 3.785 ;
        RECT 13.605 2.505 13.775 2.675 ;
        RECT 15.455 2.505 15.625 2.675 ;
        RECT 18.415 3.615 18.585 3.785 ;
        RECT 20.265 3.245 20.435 3.415 ;
        RECT 22.485 3.245 22.655 3.415 ;
        RECT 23.225 2.505 23.395 2.675 ;
        RECT 25.075 2.505 25.245 2.675 ;
        RECT 27.295 3.615 27.465 3.785 ;
        RECT 28.035 4.725 28.205 4.895 ;
        RECT 28.035 3.245 28.205 3.415 ;
        RECT 32.105 3.245 32.275 3.415 ;
        RECT 32.845 2.505 33.015 2.675 ;
        RECT 34.695 2.505 34.865 2.675 ;
        RECT 36.915 3.615 37.085 3.785 ;
        RECT 37.655 3.245 37.825 3.415 ;
        RECT 39.505 2.505 39.675 2.675 ;
        RECT 41.725 3.615 41.895 3.785 ;
        RECT 42.465 2.505 42.635 2.675 ;
        RECT 44.315 2.505 44.485 2.675 ;
        RECT 47.275 3.615 47.445 3.785 ;
        RECT 49.125 3.245 49.295 3.415 ;
        RECT 51.345 3.245 51.515 3.415 ;
        RECT 52.085 2.505 52.255 2.675 ;
        RECT 53.935 2.505 54.105 2.675 ;
        RECT 56.155 3.615 56.325 3.785 ;
        RECT 56.895 3.615 57.065 3.785 ;
        RECT 56.895 3.245 57.065 3.415 ;
        RECT 60.965 3.245 61.135 3.415 ;
        RECT 61.705 2.505 61.875 2.675 ;
        RECT 63.555 2.505 63.725 2.675 ;
        RECT 65.775 3.615 65.945 3.785 ;
        RECT 66.515 3.245 66.685 3.415 ;
        RECT 68.365 2.505 68.535 2.675 ;
        RECT 70.585 3.615 70.755 3.785 ;
        RECT 71.325 2.505 71.495 2.675 ;
        RECT 73.175 2.505 73.345 2.675 ;
        RECT 76.135 3.615 76.305 3.785 ;
        RECT 77.985 3.245 78.155 3.415 ;
        RECT 80.205 2.135 80.375 2.305 ;
        RECT 80.945 2.505 81.115 2.675 ;
        RECT 82.795 2.505 82.965 2.675 ;
        RECT 85.015 3.615 85.185 3.785 ;
        RECT 90.605 5.125 90.775 5.295 ;
        RECT 91.925 5.125 92.095 5.295 ;
        RECT 93.945 5.125 94.115 5.295 ;
        RECT 85.755 2.135 85.925 2.305 ;
        RECT 87.235 4.355 87.405 4.525 ;
        RECT 88.345 3.985 88.515 4.155 ;
        RECT 90.935 4.355 91.105 4.525 ;
        RECT 92.415 1.995 92.585 2.165 ;
        RECT 93.895 1.995 94.065 2.165 ;
        RECT 95.005 3.985 95.175 4.155 ;
        RECT 95.745 3.985 95.915 4.155 ;
        RECT 88.645 1.095 88.815 1.265 ;
        RECT 91.975 1.095 92.145 1.265 ;
        RECT 97.225 3.985 97.395 4.155 ;
        RECT 95.305 1.095 95.475 1.265 ;
      LAYER met1 ;
        RECT 88.575 5.295 88.805 5.325 ;
        RECT 90.575 5.295 90.805 5.325 ;
        RECT 91.895 5.295 92.125 5.325 ;
        RECT 93.915 5.295 94.145 5.325 ;
        RECT 88.545 5.125 90.835 5.295 ;
        RECT 91.865 5.125 94.175 5.295 ;
        RECT 88.575 5.095 88.805 5.125 ;
        RECT 90.575 5.095 90.805 5.125 ;
        RECT 91.895 5.095 92.125 5.125 ;
        RECT 93.915 5.095 94.145 5.125 ;
        RECT 28.005 4.895 28.235 4.925 ;
        RECT 27.975 4.725 75.195 4.895 ;
        RECT 28.005 4.695 28.235 4.725 ;
        RECT 75.025 4.525 75.195 4.725 ;
        RECT 87.205 4.525 87.435 4.555 ;
        RECT 90.905 4.525 91.135 4.555 ;
        RECT 75.025 4.365 91.165 4.525 ;
        RECT 75.105 4.355 91.165 4.365 ;
        RECT 87.205 4.325 87.435 4.355 ;
        RECT 90.905 4.325 91.135 4.355 ;
        RECT 88.315 4.155 88.545 4.185 ;
        RECT 94.975 4.155 95.205 4.185 ;
        RECT 95.715 4.155 95.945 4.185 ;
        RECT 97.195 4.155 97.425 4.185 ;
        RECT 65.035 3.985 95.235 4.155 ;
        RECT 95.685 3.985 97.455 4.155 ;
        RECT 8.025 3.785 8.255 3.815 ;
        RECT 12.835 3.785 13.065 3.815 ;
        RECT 18.385 3.785 18.615 3.815 ;
        RECT 27.265 3.785 27.495 3.815 ;
        RECT 36.885 3.785 37.115 3.815 ;
        RECT 41.695 3.785 41.925 3.815 ;
        RECT 47.245 3.785 47.475 3.815 ;
        RECT 56.125 3.785 56.355 3.815 ;
        RECT 56.865 3.785 57.095 3.815 ;
        RECT 65.035 3.785 65.205 3.985 ;
        RECT 88.315 3.955 88.545 3.985 ;
        RECT 94.975 3.955 95.205 3.985 ;
        RECT 95.715 3.955 95.945 3.985 ;
        RECT 97.195 3.955 97.425 3.985 ;
        RECT 65.745 3.785 65.975 3.815 ;
        RECT 70.555 3.785 70.785 3.815 ;
        RECT 76.105 3.785 76.335 3.815 ;
        RECT 84.985 3.785 85.215 3.815 ;
        RECT 7.995 3.615 27.525 3.785 ;
        RECT 36.855 3.615 56.385 3.785 ;
        RECT 56.835 3.615 65.205 3.785 ;
        RECT 65.715 3.615 85.245 3.785 ;
        RECT 8.025 3.585 8.255 3.615 ;
        RECT 12.835 3.585 13.065 3.615 ;
        RECT 18.385 3.585 18.615 3.615 ;
        RECT 27.265 3.585 27.495 3.615 ;
        RECT 36.885 3.585 37.115 3.615 ;
        RECT 41.695 3.585 41.925 3.615 ;
        RECT 47.245 3.585 47.475 3.615 ;
        RECT 56.125 3.585 56.355 3.615 ;
        RECT 56.865 3.585 57.095 3.615 ;
        RECT 65.745 3.585 65.975 3.615 ;
        RECT 70.555 3.585 70.785 3.615 ;
        RECT 76.105 3.585 76.335 3.615 ;
        RECT 84.985 3.585 85.215 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 8.765 3.415 8.995 3.445 ;
        RECT 20.235 3.415 20.465 3.445 ;
        RECT 22.455 3.415 22.685 3.445 ;
        RECT 28.005 3.415 28.235 3.445 ;
        RECT 32.075 3.415 32.305 3.445 ;
        RECT 37.625 3.415 37.855 3.445 ;
        RECT 49.095 3.415 49.325 3.445 ;
        RECT 51.315 3.415 51.545 3.445 ;
        RECT 56.865 3.415 57.095 3.445 ;
        RECT 60.935 3.415 61.165 3.445 ;
        RECT 66.485 3.415 66.715 3.445 ;
        RECT 77.955 3.415 78.185 3.445 ;
        RECT 3.185 3.245 20.495 3.415 ;
        RECT 22.425 3.245 28.265 3.415 ;
        RECT 32.045 3.245 49.355 3.415 ;
        RECT 51.285 3.245 57.125 3.415 ;
        RECT 60.905 3.245 78.215 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 8.765 3.215 8.995 3.245 ;
        RECT 20.235 3.215 20.465 3.245 ;
        RECT 22.455 3.215 22.685 3.245 ;
        RECT 28.005 3.215 28.235 3.245 ;
        RECT 32.075 3.215 32.305 3.245 ;
        RECT 37.625 3.215 37.855 3.245 ;
        RECT 49.095 3.215 49.325 3.245 ;
        RECT 51.315 3.215 51.545 3.245 ;
        RECT 56.865 3.215 57.095 3.245 ;
        RECT 60.935 3.215 61.165 3.245 ;
        RECT 66.485 3.215 66.715 3.245 ;
        RECT 77.955 3.215 78.185 3.245 ;
        RECT 3.955 2.675 4.185 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 10.615 2.675 10.845 2.705 ;
        RECT 13.575 2.675 13.805 2.705 ;
        RECT 15.425 2.675 15.655 2.705 ;
        RECT 23.195 2.675 23.425 2.705 ;
        RECT 25.045 2.675 25.275 2.705 ;
        RECT 32.815 2.675 33.045 2.705 ;
        RECT 34.665 2.675 34.895 2.705 ;
        RECT 39.475 2.675 39.705 2.705 ;
        RECT 42.435 2.675 42.665 2.705 ;
        RECT 44.285 2.675 44.515 2.705 ;
        RECT 52.055 2.675 52.285 2.705 ;
        RECT 53.905 2.675 54.135 2.705 ;
        RECT 61.675 2.675 61.905 2.705 ;
        RECT 63.525 2.675 63.755 2.705 ;
        RECT 68.335 2.675 68.565 2.705 ;
        RECT 71.295 2.675 71.525 2.705 ;
        RECT 73.145 2.675 73.375 2.705 ;
        RECT 80.915 2.675 81.145 2.705 ;
        RECT 82.765 2.675 82.995 2.705 ;
        RECT 3.925 2.505 10.875 2.675 ;
        RECT 13.545 2.505 15.685 2.675 ;
        RECT 23.165 2.505 25.305 2.675 ;
        RECT 32.785 2.505 39.735 2.675 ;
        RECT 42.405 2.505 44.545 2.675 ;
        RECT 52.025 2.505 54.165 2.675 ;
        RECT 61.645 2.505 68.595 2.675 ;
        RECT 71.265 2.505 73.405 2.675 ;
        RECT 80.885 2.505 83.025 2.675 ;
        RECT 3.955 2.475 4.185 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 10.615 2.475 10.845 2.505 ;
        RECT 13.575 2.475 13.805 2.505 ;
        RECT 15.425 2.475 15.655 2.505 ;
        RECT 23.195 2.475 23.425 2.505 ;
        RECT 25.045 2.475 25.275 2.505 ;
        RECT 32.815 2.475 33.045 2.505 ;
        RECT 34.665 2.475 34.895 2.505 ;
        RECT 39.475 2.475 39.705 2.505 ;
        RECT 42.435 2.475 42.665 2.505 ;
        RECT 44.285 2.475 44.515 2.505 ;
        RECT 52.055 2.475 52.285 2.505 ;
        RECT 53.905 2.475 54.135 2.505 ;
        RECT 61.675 2.475 61.905 2.505 ;
        RECT 63.525 2.475 63.755 2.505 ;
        RECT 68.335 2.475 68.565 2.505 ;
        RECT 71.295 2.475 71.525 2.505 ;
        RECT 73.145 2.475 73.375 2.505 ;
        RECT 80.915 2.475 81.145 2.505 ;
        RECT 82.765 2.475 82.995 2.505 ;
        RECT 80.175 2.305 80.405 2.335 ;
        RECT 85.725 2.305 85.955 2.335 ;
        RECT 80.145 2.165 92.615 2.305 ;
        RECT 93.865 2.165 94.095 2.195 ;
        RECT 80.145 2.135 94.125 2.165 ;
        RECT 80.175 2.105 80.405 2.135 ;
        RECT 85.725 2.105 85.955 2.135 ;
        RECT 92.355 1.995 94.125 2.135 ;
        RECT 92.385 1.965 92.615 1.995 ;
        RECT 93.865 1.965 94.095 1.995 ;
        RECT 88.615 1.265 88.845 1.295 ;
        RECT 91.945 1.265 92.175 1.295 ;
        RECT 95.275 1.265 95.505 1.295 ;
        RECT 88.585 1.095 95.535 1.265 ;
        RECT 88.615 1.065 88.845 1.095 ;
        RECT 91.945 1.065 92.175 1.095 ;
        RECT 95.275 1.065 95.505 1.095 ;
  END
END TMRDFFSNRNQX1






MACRO VOTER3X1
  CLASS CORE ;
  FOREIGN VOTER3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.210 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN A
    ANTENNAGATEAREA 2.053700 ;
    PORT
      LAYER li1 ;
        RECT 1.805 4.710 1.975 4.870 ;
        RECT 1.765 4.540 1.975 4.710 ;
        RECT 8.425 4.540 8.615 4.870 ;
        RECT 1.765 1.915 1.935 4.540 ;
        RECT 8.425 1.915 8.595 4.540 ;
      LAYER mcon ;
        RECT 1.765 3.985 1.935 4.155 ;
        RECT 8.425 3.985 8.595 4.155 ;
      LAYER met1 ;
        RECT 1.735 4.155 1.965 4.185 ;
        RECT 8.395 4.155 8.625 4.185 ;
        RECT 1.705 3.985 8.655 4.155 ;
        RECT 1.735 3.955 1.965 3.985 ;
        RECT 8.395 3.955 8.625 3.985 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 2.066500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.915 0.825 4.870 ;
        RECT 4.355 1.915 4.525 4.870 ;
      LAYER mcon ;
        RECT 0.655 4.355 0.825 4.525 ;
        RECT 4.355 4.355 4.525 4.525 ;
      LAYER met1 ;
        RECT 0.625 4.525 0.855 4.555 ;
        RECT 4.325 4.525 4.555 4.555 ;
        RECT 0.595 4.355 4.585 4.525 ;
        RECT 0.625 4.325 0.855 4.355 ;
        RECT 4.325 4.325 4.555 4.355 ;
    END
  END B
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 12.645 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 12.380 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.125 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.125 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 6.490 4.110 6.830 7.230 ;
        RECT 9.820 4.110 10.160 7.230 ;
        RECT 10.580 5.185 10.750 7.230 ;
        RECT 11.460 5.185 11.630 7.230 ;
        RECT 12.040 4.110 12.380 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 12.380 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 12.380 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 4.425 0.170 4.595 1.120 ;
        RECT 6.490 0.170 6.830 2.720 ;
        RECT 7.755 0.170 7.925 1.120 ;
        RECT 9.820 0.170 10.160 2.720 ;
        RECT 10.535 0.620 10.705 1.750 ;
        RECT 11.505 0.620 11.675 1.750 ;
        RECT 10.535 0.450 11.675 0.620 ;
        RECT 10.535 0.170 10.705 0.450 ;
        RECT 11.020 0.170 11.190 0.450 ;
        RECT 11.505 0.170 11.675 0.450 ;
        RECT 12.040 0.170 12.380 2.720 ;
        RECT -0.170 -0.170 12.380 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 12.380 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 6.825 1.325 6.995 ;
        RECT 1.145 5.295 1.315 6.825 ;
        RECT 2.025 5.295 2.195 6.995 ;
        RECT 1.145 5.125 2.195 5.295 ;
        RECT 2.025 5.045 2.195 5.125 ;
        RECT 4.025 6.825 5.955 6.995 ;
        RECT 4.025 5.045 4.195 6.825 ;
        RECT 4.465 5.295 4.635 6.565 ;
        RECT 4.905 5.555 5.075 6.825 ;
        RECT 5.345 5.295 5.515 6.565 ;
        RECT 5.785 5.375 5.955 6.825 ;
        RECT 7.365 6.825 9.295 6.995 ;
        RECT 4.465 5.125 5.515 5.295 ;
        RECT 5.345 5.045 5.515 5.125 ;
        RECT 7.365 5.045 7.535 6.825 ;
        RECT 7.805 5.295 7.975 6.565 ;
        RECT 8.245 5.555 8.415 6.825 ;
        RECT 8.685 5.295 8.855 6.565 ;
        RECT 9.125 5.555 9.295 6.825 ;
        RECT 7.805 5.125 9.335 5.295 ;
        RECT 5.835 1.915 6.005 4.870 ;
        RECT 7.315 1.915 7.485 4.870 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.170 2.235 1.345 ;
        RECT 2.060 1.015 2.235 1.170 ;
        RECT 2.060 0.835 2.230 1.015 ;
        RECT 2.550 0.615 2.720 1.745 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 3.940 1.665 4.110 1.745 ;
        RECT 4.910 1.665 5.080 1.745 ;
        RECT 3.940 1.495 5.080 1.665 ;
        RECT 3.940 0.365 4.110 1.495 ;
        RECT 4.910 0.615 5.080 1.495 ;
        RECT 5.395 0.835 5.565 1.345 ;
        RECT 5.880 0.615 6.050 1.745 ;
        RECT 4.910 0.445 6.050 0.615 ;
        RECT 4.910 0.365 5.080 0.445 ;
        RECT 5.880 0.365 6.050 0.445 ;
        RECT 7.270 1.665 7.440 1.745 ;
        RECT 8.240 1.665 8.410 1.745 ;
        RECT 9.165 1.730 9.335 5.125 ;
        RECT 10.645 1.920 10.815 4.865 ;
        RECT 11.020 4.665 11.190 7.020 ;
        RECT 11.020 4.495 11.555 4.665 ;
        RECT 11.385 2.165 11.555 4.495 ;
        RECT 11.015 1.995 11.555 2.165 ;
        RECT 7.270 1.495 8.410 1.665 ;
        RECT 7.270 0.365 7.440 1.495 ;
        RECT 8.240 0.615 8.410 1.495 ;
        RECT 8.725 1.560 9.335 1.730 ;
        RECT 8.725 0.835 8.895 1.560 ;
        RECT 9.210 0.615 9.380 1.390 ;
        RECT 11.015 0.840 11.185 1.995 ;
        RECT 8.240 0.445 9.380 0.615 ;
        RECT 8.240 0.365 8.410 0.445 ;
        RECT 9.210 0.365 9.380 0.445 ;
      LAYER mcon ;
        RECT 2.025 5.125 2.195 5.295 ;
        RECT 4.025 5.125 4.195 5.295 ;
        RECT 5.345 5.125 5.515 5.295 ;
        RECT 7.365 5.125 7.535 5.295 ;
        RECT 5.835 1.995 6.005 2.165 ;
        RECT 7.315 1.995 7.485 2.165 ;
        RECT 9.165 3.985 9.335 4.155 ;
        RECT 2.065 1.095 2.235 1.265 ;
        RECT 5.395 1.095 5.565 1.265 ;
        RECT 10.645 3.985 10.815 4.155 ;
        RECT 8.725 1.095 8.895 1.265 ;
      LAYER met1 ;
        RECT 1.995 5.295 2.225 5.325 ;
        RECT 3.995 5.295 4.225 5.325 ;
        RECT 5.315 5.295 5.545 5.325 ;
        RECT 7.335 5.295 7.565 5.325 ;
        RECT 1.965 5.125 4.255 5.295 ;
        RECT 5.285 5.125 7.595 5.295 ;
        RECT 1.995 5.095 2.225 5.125 ;
        RECT 3.995 5.095 4.225 5.125 ;
        RECT 5.315 5.095 5.545 5.125 ;
        RECT 7.335 5.095 7.565 5.125 ;
        RECT 9.135 4.155 9.365 4.185 ;
        RECT 10.615 4.155 10.845 4.185 ;
        RECT 9.105 3.985 10.875 4.155 ;
        RECT 9.135 3.955 9.365 3.985 ;
        RECT 10.615 3.955 10.845 3.985 ;
        RECT 5.805 2.165 6.035 2.195 ;
        RECT 7.285 2.165 7.515 2.195 ;
        RECT 5.775 1.995 7.545 2.165 ;
        RECT 5.805 1.965 6.035 1.995 ;
        RECT 7.285 1.965 7.515 1.995 ;
        RECT 2.035 1.265 2.265 1.295 ;
        RECT 5.365 1.265 5.595 1.295 ;
        RECT 8.695 1.265 8.925 1.295 ;
        RECT 2.005 1.095 8.955 1.265 ;
        RECT 2.035 1.065 2.265 1.095 ;
        RECT 5.365 1.065 5.595 1.095 ;
        RECT 8.695 1.065 8.925 1.095 ;
  END
END VOTER3X1






MACRO VOTERN3X1
  CLASS CORE ;
  FOREIGN VOTERN3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.990 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN A
    ANTENNAGATEAREA 2.053700 ;
    PORT
      LAYER li1 ;
        RECT 1.805 4.710 1.975 4.870 ;
        RECT 1.765 4.540 1.975 4.710 ;
        RECT 8.425 4.540 8.615 4.870 ;
        RECT 1.765 1.915 1.935 4.540 ;
        RECT 8.425 1.915 8.595 4.540 ;
      LAYER mcon ;
        RECT 1.765 3.985 1.935 4.155 ;
        RECT 8.425 3.985 8.595 4.155 ;
      LAYER met1 ;
        RECT 1.735 4.155 1.965 4.185 ;
        RECT 8.395 4.155 8.625 4.185 ;
        RECT 1.705 3.985 8.655 4.155 ;
        RECT 1.735 3.955 1.965 3.985 ;
        RECT 8.395 3.955 8.625 3.985 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 2.066500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.915 0.825 4.870 ;
        RECT 4.355 1.915 4.525 4.870 ;
      LAYER mcon ;
        RECT 0.655 4.355 0.825 4.525 ;
        RECT 4.355 4.355 4.525 4.525 ;
      LAYER met1 ;
        RECT 0.625 4.525 0.855 4.555 ;
        RECT 4.325 4.525 4.555 4.555 ;
        RECT 0.595 4.355 4.585 4.525 ;
        RECT 0.625 4.325 0.855 4.355 ;
        RECT 4.325 4.325 4.555 4.355 ;
    END
  END B
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 10.425 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 10.160 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.125 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.125 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 6.490 4.110 6.830 7.230 ;
        RECT 9.820 4.110 10.160 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 10.160 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 10.160 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 4.425 0.170 4.595 1.120 ;
        RECT 6.490 0.170 6.830 2.720 ;
        RECT 7.755 0.170 7.925 1.120 ;
        RECT 9.820 0.170 10.160 2.720 ;
        RECT -0.170 -0.170 10.160 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 10.160 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.145 6.825 1.325 6.995 ;
        RECT 1.145 5.295 1.315 6.825 ;
        RECT 2.025 5.295 2.195 6.995 ;
        RECT 1.145 5.125 2.195 5.295 ;
        RECT 2.025 5.045 2.195 5.125 ;
        RECT 4.025 6.825 5.955 6.995 ;
        RECT 4.025 5.045 4.195 6.825 ;
        RECT 4.465 5.295 4.635 6.565 ;
        RECT 4.905 5.555 5.075 6.825 ;
        RECT 5.345 5.295 5.515 6.565 ;
        RECT 5.785 5.375 5.955 6.825 ;
        RECT 7.365 6.825 9.295 6.995 ;
        RECT 4.465 5.125 5.515 5.295 ;
        RECT 5.345 5.045 5.515 5.125 ;
        RECT 7.365 5.045 7.535 6.825 ;
        RECT 7.805 5.295 7.975 6.565 ;
        RECT 8.245 5.555 8.415 6.825 ;
        RECT 8.685 5.295 8.855 6.565 ;
        RECT 9.125 5.555 9.295 6.825 ;
        RECT 7.805 5.125 9.335 5.295 ;
        RECT 5.835 1.915 6.005 4.870 ;
        RECT 7.315 1.915 7.485 4.870 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.170 2.235 1.345 ;
        RECT 2.060 1.015 2.235 1.170 ;
        RECT 2.060 0.835 2.230 1.015 ;
        RECT 2.550 0.615 2.720 1.745 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 3.940 1.665 4.110 1.745 ;
        RECT 4.910 1.665 5.080 1.745 ;
        RECT 3.940 1.495 5.080 1.665 ;
        RECT 3.940 0.365 4.110 1.495 ;
        RECT 4.910 0.615 5.080 1.495 ;
        RECT 5.395 0.835 5.565 1.345 ;
        RECT 5.880 0.615 6.050 1.745 ;
        RECT 4.910 0.445 6.050 0.615 ;
        RECT 4.910 0.365 5.080 0.445 ;
        RECT 5.880 0.365 6.050 0.445 ;
        RECT 7.270 1.665 7.440 1.745 ;
        RECT 8.240 1.665 8.410 1.745 ;
        RECT 9.165 1.730 9.335 5.125 ;
        RECT 7.270 1.495 8.410 1.665 ;
        RECT 7.270 0.365 7.440 1.495 ;
        RECT 8.240 0.615 8.410 1.495 ;
        RECT 8.725 1.560 9.335 1.730 ;
        RECT 8.725 0.835 8.895 1.560 ;
        RECT 9.210 0.615 9.380 1.390 ;
        RECT 8.240 0.445 9.380 0.615 ;
        RECT 8.240 0.365 8.410 0.445 ;
        RECT 9.210 0.365 9.380 0.445 ;
      LAYER mcon ;
        RECT 2.025 5.125 2.195 5.295 ;
        RECT 4.025 5.125 4.195 5.295 ;
        RECT 5.345 5.125 5.515 5.295 ;
        RECT 7.365 5.125 7.535 5.295 ;
        RECT 5.835 1.995 6.005 2.165 ;
        RECT 7.315 1.995 7.485 2.165 ;
        RECT 2.065 1.095 2.235 1.265 ;
        RECT 5.395 1.095 5.565 1.265 ;
        RECT 8.725 1.095 8.895 1.265 ;
      LAYER met1 ;
        RECT 1.995 5.295 2.225 5.325 ;
        RECT 3.995 5.295 4.225 5.325 ;
        RECT 5.315 5.295 5.545 5.325 ;
        RECT 7.335 5.295 7.565 5.325 ;
        RECT 1.965 5.125 4.255 5.295 ;
        RECT 5.285 5.125 7.595 5.295 ;
        RECT 1.995 5.095 2.225 5.125 ;
        RECT 3.995 5.095 4.225 5.125 ;
        RECT 5.315 5.095 5.545 5.125 ;
        RECT 7.335 5.095 7.565 5.125 ;
        RECT 5.805 2.165 6.035 2.195 ;
        RECT 7.285 2.165 7.515 2.195 ;
        RECT 5.775 1.995 7.545 2.165 ;
        RECT 5.805 1.965 6.035 1.995 ;
        RECT 7.285 1.965 7.515 1.995 ;
        RECT 2.035 1.265 2.265 1.295 ;
        RECT 5.365 1.265 5.595 1.295 ;
        RECT 8.695 1.265 8.925 1.295 ;
        RECT 2.005 1.095 8.955 1.265 ;
        RECT 2.035 1.065 2.265 1.095 ;
        RECT 5.365 1.065 5.595 1.095 ;
        RECT 8.695 1.065 8.925 1.095 ;
  END
END VOTERN3X1






MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.100 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Y
    ANTENNADIFFAREA 1.543800 ;
    PORT
      LAYER li1 ;
        RECT 4.245 5.290 4.415 6.560 ;
        RECT 7.575 5.290 7.745 6.560 ;
        RECT 4.245 5.120 4.895 5.290 ;
        RECT 7.575 5.120 8.225 5.290 ;
        RECT 4.725 1.735 4.895 5.120 ;
        RECT 8.055 1.735 8.225 5.120 ;
        RECT 4.285 1.565 4.895 1.735 ;
        RECT 7.615 1.565 8.225 1.735 ;
        RECT 4.285 0.835 4.455 1.565 ;
        RECT 7.615 0.835 7.785 1.565 ;
      LAYER mcon ;
        RECT 4.725 3.615 4.895 3.785 ;
        RECT 8.055 3.615 8.225 3.785 ;
      LAYER met1 ;
        RECT 4.695 3.785 4.925 3.815 ;
        RECT 8.025 3.785 8.255 3.815 ;
        RECT 4.665 3.615 8.285 3.785 ;
        RECT 4.695 3.585 4.925 3.615 ;
        RECT 8.025 3.585 8.255 3.615 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
      LAYER mcon ;
        RECT 0.655 3.985 0.825 4.155 ;
        RECT 3.245 3.985 3.415 4.155 ;
      LAYER met1 ;
        RECT 0.625 4.155 0.855 4.185 ;
        RECT 3.215 4.155 3.445 4.185 ;
        RECT 0.595 3.985 3.475 4.155 ;
        RECT 0.625 3.955 0.855 3.985 ;
        RECT 3.215 3.955 3.445 3.985 ;
    END
  END A
  PIN A
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
        RECT 7.685 1.915 7.855 4.865 ;
      LAYER mcon ;
        RECT 1.395 2.505 1.565 2.675 ;
        RECT 7.685 2.505 7.855 2.675 ;
      LAYER met1 ;
        RECT 1.365 2.675 1.595 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 1.335 2.505 7.915 2.675 ;
        RECT 1.365 2.475 1.595 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 4.355 3.905 4.525 4.865 ;
        RECT 6.575 1.915 6.745 3.495 ;
        RECT 10.275 1.920 10.445 4.865 ;
      LAYER mcon ;
        RECT 4.355 3.985 4.525 4.155 ;
        RECT 10.275 3.985 10.445 4.155 ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 10.275 3.245 10.445 3.415 ;
      LAYER met1 ;
        RECT 4.325 4.155 4.555 4.185 ;
        RECT 10.245 4.155 10.475 4.185 ;
        RECT 4.295 3.985 10.505 4.155 ;
        RECT 4.325 3.955 4.555 3.985 ;
        RECT 10.245 3.955 10.475 3.985 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 10.245 3.415 10.475 3.445 ;
        RECT 6.515 3.245 10.505 3.415 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 10.245 3.215 10.475 3.245 ;
    END
  END B
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 11.535 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 11.270 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
        RECT 3.365 5.550 3.535 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
        RECT 6.695 5.550 6.865 7.230 ;
        RECT 8.710 4.110 9.050 7.230 ;
        RECT 9.460 5.185 9.630 7.230 ;
        RECT 10.340 5.185 10.510 7.230 ;
        RECT 10.930 4.110 11.270 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 11.270 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 11.270 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT 3.315 0.170 3.485 1.120 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT 6.645 0.170 6.815 1.120 ;
        RECT 8.710 0.170 9.050 2.720 ;
        RECT 9.415 0.620 9.585 1.750 ;
        RECT 10.385 0.620 10.555 1.750 ;
        RECT 9.415 0.450 10.555 0.620 ;
        RECT 9.415 0.170 9.585 0.450 ;
        RECT 9.900 0.170 10.070 0.450 ;
        RECT 10.385 0.170 10.555 0.450 ;
        RECT 10.930 0.170 11.270 2.720 ;
        RECT -0.170 -0.170 11.270 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 11.270 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 2.925 5.290 3.095 6.900 ;
        RECT 3.805 6.820 4.855 6.990 ;
        RECT 3.805 5.290 3.975 6.820 ;
        RECT 4.685 5.550 4.855 6.820 ;
        RECT 2.925 5.120 3.975 5.290 ;
        RECT 6.255 5.290 6.425 6.900 ;
        RECT 7.135 6.820 8.185 6.990 ;
        RECT 7.135 5.290 7.305 6.820 ;
        RECT 8.015 5.550 8.185 6.820 ;
        RECT 6.255 5.120 7.305 5.290 ;
        RECT 6.575 4.275 6.745 4.865 ;
        RECT 9.900 4.665 10.070 7.020 ;
        RECT 9.535 4.495 10.070 4.665 ;
        RECT 4.355 1.915 4.525 3.125 ;
        RECT 9.535 2.165 9.705 4.495 ;
        RECT 9.535 1.995 10.075 2.165 ;
        RECT 2.830 1.665 3.000 1.745 ;
        RECT 3.800 1.665 3.970 1.745 ;
        RECT 2.830 1.495 3.970 1.665 ;
        RECT 2.830 0.365 3.000 1.495 ;
        RECT 3.800 0.615 3.970 1.495 ;
        RECT 6.160 1.665 6.330 1.745 ;
        RECT 7.130 1.665 7.300 1.745 ;
        RECT 6.160 1.495 7.300 1.665 ;
        RECT 4.770 0.615 4.940 1.385 ;
        RECT 3.800 0.445 4.940 0.615 ;
        RECT 3.800 0.365 3.970 0.445 ;
        RECT 4.770 0.365 4.940 0.445 ;
        RECT 6.160 0.365 6.330 1.495 ;
        RECT 7.130 0.615 7.300 1.495 ;
        RECT 8.100 0.615 8.270 1.385 ;
        RECT 9.905 0.840 10.075 1.995 ;
        RECT 7.130 0.445 8.270 0.615 ;
        RECT 7.130 0.365 7.300 0.445 ;
        RECT 8.100 0.365 8.270 0.445 ;
      LAYER mcon ;
        RECT 6.575 4.355 6.745 4.525 ;
        RECT 9.535 4.355 9.705 4.525 ;
        RECT 4.355 2.875 4.525 3.045 ;
        RECT 9.535 2.875 9.705 3.045 ;
      LAYER met1 ;
        RECT 6.545 4.525 6.775 4.555 ;
        RECT 9.505 4.525 9.735 4.555 ;
        RECT 6.515 4.355 9.765 4.525 ;
        RECT 6.545 4.325 6.775 4.355 ;
        RECT 9.505 4.325 9.735 4.355 ;
        RECT 4.325 3.045 4.555 3.075 ;
        RECT 9.505 3.045 9.735 3.075 ;
        RECT 4.295 2.875 9.765 3.045 ;
        RECT 4.325 2.845 4.555 2.875 ;
        RECT 9.505 2.845 9.735 2.875 ;
  END
END XNOR2X1






MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.100 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Y
    ANTENNADIFFAREA 1.543800 ;
    PORT
      LAYER li1 ;
        RECT 4.245 5.290 4.415 6.560 ;
        RECT 7.575 5.290 7.745 6.560 ;
        RECT 4.245 5.120 4.895 5.290 ;
        RECT 7.575 5.120 8.225 5.290 ;
        RECT 4.725 1.740 4.895 5.120 ;
        RECT 8.055 1.740 8.225 5.120 ;
        RECT 4.285 1.570 4.895 1.740 ;
        RECT 7.615 1.570 8.225 1.740 ;
        RECT 4.285 0.840 4.455 1.570 ;
        RECT 7.615 0.840 7.785 1.570 ;
      LAYER mcon ;
        RECT 4.725 3.615 4.895 3.785 ;
        RECT 8.055 3.615 8.225 3.785 ;
      LAYER met1 ;
        RECT 4.695 3.785 4.925 3.815 ;
        RECT 8.025 3.785 8.255 3.815 ;
        RECT 4.665 3.615 8.285 3.785 ;
        RECT 4.695 3.585 4.925 3.615 ;
        RECT 8.025 3.585 8.255 3.615 ;
    END
  END Y
  PIN A
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 3.245 1.920 3.415 4.865 ;
      LAYER mcon ;
        RECT 0.655 3.985 0.825 4.155 ;
        RECT 3.245 3.985 3.415 4.155 ;
      LAYER met1 ;
        RECT 0.625 4.155 0.855 4.185 ;
        RECT 3.215 4.155 3.445 4.185 ;
        RECT 0.595 3.985 3.475 4.155 ;
        RECT 0.625 3.955 0.855 3.985 ;
        RECT 3.215 3.955 3.445 3.985 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA 2.054500 ;
    PORT
      LAYER li1 ;
        RECT 6.575 4.275 6.745 4.865 ;
        RECT 4.355 1.920 4.525 3.125 ;
        RECT 10.275 1.920 10.445 4.865 ;
      LAYER mcon ;
        RECT 6.575 4.355 6.745 4.525 ;
        RECT 10.275 4.355 10.445 4.525 ;
        RECT 4.355 2.875 4.525 3.045 ;
        RECT 10.275 2.875 10.445 3.045 ;
      LAYER met1 ;
        RECT 6.545 4.525 6.775 4.555 ;
        RECT 10.245 4.525 10.475 4.555 ;
        RECT 6.515 4.355 10.505 4.525 ;
        RECT 6.545 4.325 6.775 4.355 ;
        RECT 10.245 4.325 10.475 4.355 ;
        RECT 4.325 3.045 4.555 3.075 ;
        RECT 10.245 3.045 10.475 3.075 ;
        RECT 4.295 2.875 10.505 3.045 ;
        RECT 4.325 2.845 4.555 2.875 ;
        RECT 10.245 2.845 10.475 2.875 ;
    END
  END B
  PIN VPWR
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 11.535 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 11.270 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
        RECT 3.365 5.550 3.535 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
        RECT 6.695 5.550 6.865 7.230 ;
        RECT 8.710 4.110 9.050 7.230 ;
        RECT 9.460 5.185 9.630 7.230 ;
        RECT 10.340 5.185 10.510 7.230 ;
        RECT 10.930 4.110 11.270 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 11.270 7.570 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 11.270 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT 3.315 0.170 3.485 1.125 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT 6.645 0.170 6.815 1.125 ;
        RECT 8.710 0.170 9.050 2.720 ;
        RECT 9.415 0.620 9.585 1.750 ;
        RECT 10.385 0.620 10.555 1.750 ;
        RECT 9.415 0.450 10.555 0.620 ;
        RECT 9.415 0.170 9.585 0.450 ;
        RECT 9.900 0.170 10.070 0.450 ;
        RECT 10.385 0.170 10.555 0.450 ;
        RECT 10.930 0.170 11.270 2.720 ;
        RECT -0.170 -0.170 11.270 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 11.270 0.170 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 2.925 5.290 3.095 6.900 ;
        RECT 3.805 6.820 4.855 6.990 ;
        RECT 3.805 5.290 3.975 6.820 ;
        RECT 4.685 5.550 4.855 6.820 ;
        RECT 2.925 5.120 3.975 5.290 ;
        RECT 6.255 5.290 6.425 6.900 ;
        RECT 7.135 6.820 8.185 6.990 ;
        RECT 7.135 5.290 7.305 6.820 ;
        RECT 8.015 5.550 8.185 6.820 ;
        RECT 6.255 5.120 7.305 5.290 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 4.355 3.905 4.525 4.865 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
        RECT 6.575 1.920 6.745 3.495 ;
        RECT 7.685 1.920 7.855 4.865 ;
        RECT 9.900 4.665 10.070 7.020 ;
        RECT 9.535 4.495 10.070 4.665 ;
        RECT 9.535 2.165 9.705 4.495 ;
        RECT 9.535 1.995 10.075 2.165 ;
        RECT 2.830 1.670 3.000 1.750 ;
        RECT 3.800 1.670 3.970 1.750 ;
        RECT 2.830 1.500 3.970 1.670 ;
        RECT 2.830 0.370 3.000 1.500 ;
        RECT 3.800 0.620 3.970 1.500 ;
        RECT 6.160 1.670 6.330 1.750 ;
        RECT 7.130 1.670 7.300 1.750 ;
        RECT 6.160 1.500 7.300 1.670 ;
        RECT 4.770 0.620 4.940 1.390 ;
        RECT 3.800 0.450 4.940 0.620 ;
        RECT 3.800 0.370 3.970 0.450 ;
        RECT 4.770 0.370 4.940 0.450 ;
        RECT 6.160 0.370 6.330 1.500 ;
        RECT 7.130 0.620 7.300 1.500 ;
        RECT 8.100 0.620 8.270 1.390 ;
        RECT 9.905 0.840 10.075 1.995 ;
        RECT 7.130 0.450 8.270 0.620 ;
        RECT 7.130 0.370 7.300 0.450 ;
        RECT 8.100 0.370 8.270 0.450 ;
      LAYER mcon ;
        RECT 4.355 3.985 4.525 4.155 ;
        RECT 1.395 2.505 1.565 2.675 ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 7.685 2.505 7.855 2.675 ;
        RECT 9.535 3.985 9.705 4.155 ;
        RECT 9.535 3.245 9.705 3.415 ;
      LAYER met1 ;
        RECT 4.325 4.155 4.555 4.185 ;
        RECT 9.505 4.155 9.735 4.185 ;
        RECT 4.295 3.985 9.765 4.155 ;
        RECT 4.325 3.955 4.555 3.985 ;
        RECT 9.505 3.955 9.735 3.985 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 9.505 3.415 9.735 3.445 ;
        RECT 6.515 3.245 9.765 3.415 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 9.505 3.215 9.735 3.245 ;
        RECT 1.365 2.675 1.595 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 1.335 2.505 7.915 2.675 ;
        RECT 1.365 2.475 1.595 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
  END
END XOR2X1


END LIBRARY
