VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO FA
  CLASS CORE ;
  FOREIGN FA ;
  ORIGIN 0.000 0.000 ;
  SIZE 38.850 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.543800 ;
    PORT
      LAYER li1 ;
        RECT 15.345 5.290 15.515 6.560 ;
        RECT 18.675 5.290 18.845 6.560 ;
        RECT 15.345 5.120 15.995 5.290 ;
        RECT 18.675 5.120 19.325 5.290 ;
        RECT 15.825 1.740 15.995 5.120 ;
        RECT 19.155 1.740 19.325 5.120 ;
        RECT 15.385 1.570 15.995 1.740 ;
        RECT 18.715 1.570 19.325 1.740 ;
        RECT 15.385 0.840 15.555 1.570 ;
        RECT 18.715 0.840 18.885 1.570 ;
      LAYER mcon ;
        RECT 15.825 3.615 15.995 3.785 ;
        RECT 19.155 3.615 19.325 3.785 ;
      LAYER met1 ;
        RECT 15.795 3.785 16.025 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 15.765 3.615 19.385 3.785 ;
        RECT 15.795 3.585 16.025 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
    END
  END SUM
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 37.660 4.665 37.830 7.020 ;
        RECT 37.660 4.495 38.195 4.665 ;
        RECT 38.025 2.165 38.195 4.495 ;
        RECT 37.655 1.995 38.195 2.165 ;
        RECT 37.655 0.840 37.825 1.995 ;
    END
  END COUT
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.087750 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 3.245 2.305 3.415 4.865 ;
        RECT 29.545 4.710 29.715 4.865 ;
        RECT 29.515 4.535 29.715 4.710 ;
        RECT 29.515 2.305 29.685 4.535 ;
        RECT 3.165 2.135 3.495 2.305 ;
        RECT 29.435 2.135 29.765 2.305 ;
        RECT 3.245 1.920 3.415 2.135 ;
        RECT 29.515 1.915 29.685 2.135 ;
      LAYER mcon ;
        RECT 0.655 3.985 0.825 4.155 ;
        RECT 3.245 3.985 3.415 4.155 ;
        RECT 3.245 2.135 3.415 2.305 ;
        RECT 29.515 2.135 29.685 2.305 ;
      LAYER met1 ;
        RECT 0.625 4.155 0.855 4.185 ;
        RECT 3.215 4.155 3.445 4.185 ;
        RECT 0.595 3.985 3.475 4.155 ;
        RECT 0.625 3.955 0.855 3.985 ;
        RECT 3.215 3.955 3.445 3.985 ;
        RECT 3.245 2.335 3.415 2.365 ;
        RECT 29.515 2.335 29.685 2.365 ;
        RECT 3.215 2.105 3.445 2.335 ;
        RECT 29.485 2.105 29.715 2.335 ;
        RECT 3.245 1.935 3.415 2.105 ;
        RECT 29.515 1.935 29.685 2.105 ;
        RECT 3.245 1.765 29.685 1.935 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.087750 ;
    PORT
      LAYER li1 ;
        RECT 6.575 4.275 6.745 4.865 ;
        RECT 4.355 1.920 4.525 3.125 ;
        RECT 10.275 1.920 10.445 4.975 ;
        RECT 28.775 4.715 28.945 4.895 ;
        RECT 28.695 4.545 29.025 4.715 ;
        RECT 28.775 1.915 28.945 4.545 ;
      LAYER mcon ;
        RECT 6.575 4.355 6.745 4.525 ;
        RECT 10.275 4.725 10.445 4.895 ;
        RECT 28.775 4.545 28.945 4.715 ;
        RECT 10.275 4.355 10.445 4.525 ;
        RECT 4.355 2.875 4.525 3.045 ;
        RECT 10.275 2.875 10.445 3.045 ;
      LAYER met1 ;
        RECT 10.245 4.895 10.475 4.925 ;
        RECT 10.215 4.745 28.945 4.895 ;
        RECT 10.215 4.725 28.975 4.745 ;
        RECT 10.245 4.695 10.475 4.725 ;
        RECT 6.545 4.525 6.775 4.555 ;
        RECT 10.245 4.525 10.475 4.555 ;
        RECT 6.515 4.355 10.505 4.525 ;
        RECT 28.745 4.515 28.975 4.725 ;
        RECT 28.775 4.485 28.945 4.515 ;
        RECT 6.545 4.325 6.775 4.355 ;
        RECT 10.245 4.325 10.475 4.355 ;
        RECT 4.325 3.045 4.555 3.075 ;
        RECT 10.245 3.045 10.475 3.075 ;
        RECT 4.295 2.875 10.505 3.045 ;
        RECT 4.325 2.845 4.555 2.875 ;
        RECT 10.245 2.845 10.475 2.875 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.087750 ;
    PORT
      LAYER li1 ;
        RECT 17.675 4.275 17.845 4.865 ;
        RECT 15.455 1.920 15.625 3.125 ;
        RECT 21.375 1.920 21.545 4.865 ;
        RECT 23.225 1.915 23.395 4.865 ;
      LAYER mcon ;
        RECT 17.675 4.355 17.845 4.525 ;
        RECT 21.375 4.355 21.545 4.525 ;
        RECT 15.455 2.875 15.625 3.045 ;
        RECT 21.375 2.875 21.545 3.045 ;
        RECT 23.225 4.355 23.395 4.525 ;
      LAYER met1 ;
        RECT 17.645 4.525 17.875 4.555 ;
        RECT 21.345 4.525 21.575 4.555 ;
        RECT 23.195 4.525 23.425 4.555 ;
        RECT 17.615 4.355 23.455 4.525 ;
        RECT 17.645 4.325 17.875 4.355 ;
        RECT 21.345 4.325 21.575 4.355 ;
        RECT 23.195 4.325 23.425 4.355 ;
        RECT 15.425 3.045 15.655 3.075 ;
        RECT 21.345 3.045 21.575 3.075 ;
        RECT 15.395 2.875 21.605 3.045 ;
        RECT 15.425 2.845 15.655 2.875 ;
        RECT 21.345 2.845 21.575 2.875 ;
    END
  END CIN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 39.285 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 39.020 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
        RECT 3.365 5.550 3.535 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
        RECT 6.695 5.550 6.865 7.230 ;
        RECT 8.710 4.110 9.050 7.230 ;
        RECT 9.460 5.185 9.630 7.230 ;
        RECT 10.340 5.185 10.510 7.230 ;
        RECT 10.930 4.110 11.270 7.230 ;
        RECT 11.690 5.185 11.860 7.230 ;
        RECT 12.570 5.185 12.740 7.230 ;
        RECT 13.150 4.110 13.490 7.230 ;
        RECT 14.465 5.550 14.635 7.230 ;
        RECT 16.480 4.110 16.820 7.230 ;
        RECT 17.795 5.550 17.965 7.230 ;
        RECT 19.810 4.110 20.150 7.230 ;
        RECT 20.560 5.185 20.730 7.230 ;
        RECT 21.440 5.185 21.610 7.230 ;
        RECT 22.030 4.110 22.370 7.230 ;
        RECT 22.905 5.135 23.075 7.230 ;
        RECT 23.785 5.555 23.955 7.230 ;
        RECT 24.665 5.555 24.835 7.230 ;
        RECT 25.360 4.110 25.700 7.230 ;
        RECT 26.120 5.185 26.290 7.230 ;
        RECT 27.000 5.185 27.170 7.230 ;
        RECT 27.580 4.110 27.920 7.230 ;
        RECT 28.455 5.135 28.625 7.230 ;
        RECT 29.335 5.555 29.505 7.230 ;
        RECT 30.215 5.555 30.385 7.230 ;
        RECT 30.910 4.110 31.250 7.230 ;
        RECT 31.670 5.185 31.840 7.230 ;
        RECT 32.550 5.185 32.720 7.230 ;
        RECT 33.130 4.110 33.470 7.230 ;
        RECT 34.445 5.555 34.615 7.230 ;
        RECT 36.460 4.110 36.800 7.230 ;
        RECT 37.220 5.185 37.390 7.230 ;
        RECT 38.100 5.185 38.270 7.230 ;
        RECT 38.680 4.110 39.020 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.485 7.315 22.655 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.815 7.315 25.985 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.515 7.315 29.685 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.625 7.315 30.795 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 32.845 7.315 33.015 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.435 7.315 35.605 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.175 7.315 36.345 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 39.020 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 39.020 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT 3.315 0.170 3.485 1.125 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT 6.645 0.170 6.815 1.125 ;
        RECT 8.710 0.170 9.050 2.720 ;
        RECT 9.415 0.620 9.585 1.750 ;
        RECT 10.385 0.620 10.555 1.750 ;
        RECT 9.415 0.450 10.555 0.620 ;
        RECT 9.415 0.170 9.585 0.450 ;
        RECT 9.900 0.170 10.070 0.450 ;
        RECT 10.385 0.170 10.555 0.450 ;
        RECT 10.930 0.170 11.270 2.720 ;
        RECT 11.645 0.620 11.815 1.750 ;
        RECT 12.615 0.620 12.785 1.750 ;
        RECT 11.645 0.450 12.785 0.620 ;
        RECT 11.645 0.170 11.815 0.450 ;
        RECT 12.130 0.170 12.300 0.450 ;
        RECT 12.615 0.170 12.785 0.450 ;
        RECT 13.150 0.170 13.490 2.720 ;
        RECT 14.415 0.170 14.585 1.125 ;
        RECT 16.480 0.170 16.820 2.720 ;
        RECT 17.745 0.170 17.915 1.125 ;
        RECT 19.810 0.170 20.150 2.720 ;
        RECT 20.515 0.620 20.685 1.750 ;
        RECT 21.485 0.620 21.655 1.750 ;
        RECT 20.515 0.450 21.655 0.620 ;
        RECT 20.515 0.170 20.685 0.450 ;
        RECT 21.000 0.170 21.170 0.450 ;
        RECT 21.485 0.170 21.655 0.450 ;
        RECT 22.030 0.170 22.370 2.720 ;
        RECT 23.295 0.170 23.465 1.120 ;
        RECT 25.360 0.170 25.700 2.720 ;
        RECT 26.075 0.620 26.245 1.750 ;
        RECT 27.045 0.620 27.215 1.750 ;
        RECT 26.075 0.450 27.215 0.620 ;
        RECT 26.075 0.170 26.245 0.450 ;
        RECT 26.560 0.170 26.730 0.450 ;
        RECT 27.045 0.170 27.215 0.450 ;
        RECT 27.580 0.170 27.920 2.720 ;
        RECT 28.845 0.170 29.015 1.120 ;
        RECT 30.910 0.170 31.250 2.720 ;
        RECT 31.625 0.620 31.795 1.750 ;
        RECT 32.595 0.620 32.765 1.750 ;
        RECT 31.625 0.450 32.765 0.620 ;
        RECT 31.625 0.170 31.795 0.450 ;
        RECT 32.110 0.170 32.280 0.450 ;
        RECT 32.595 0.170 32.765 0.450 ;
        RECT 33.130 0.170 33.470 2.720 ;
        RECT 33.910 0.615 34.080 1.745 ;
        RECT 34.880 0.615 35.050 1.390 ;
        RECT 35.850 0.615 36.020 1.390 ;
        RECT 33.910 0.445 36.020 0.615 ;
        RECT 33.910 0.170 34.080 0.445 ;
        RECT 34.395 0.170 34.565 0.445 ;
        RECT 34.880 0.170 35.050 0.445 ;
        RECT 35.365 0.170 35.535 0.445 ;
        RECT 35.850 0.170 36.020 0.445 ;
        RECT 36.460 0.170 36.800 2.720 ;
        RECT 37.175 0.620 37.345 1.750 ;
        RECT 38.145 0.620 38.315 1.750 ;
        RECT 37.175 0.450 38.315 0.620 ;
        RECT 37.175 0.170 37.345 0.450 ;
        RECT 37.660 0.170 37.830 0.450 ;
        RECT 38.145 0.170 38.315 0.450 ;
        RECT 38.680 0.170 39.020 2.720 ;
        RECT -0.170 -0.170 39.020 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.485 -0.085 22.655 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.815 -0.085 25.985 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.515 -0.085 29.685 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.625 -0.085 30.795 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 32.845 -0.085 33.015 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.435 -0.085 35.605 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.175 -0.085 36.345 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 39.020 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 2.925 5.290 3.095 6.900 ;
        RECT 3.805 6.820 4.855 6.990 ;
        RECT 3.805 5.290 3.975 6.820 ;
        RECT 2.925 5.120 3.975 5.290 ;
        RECT 4.245 5.290 4.415 6.560 ;
        RECT 4.685 5.550 4.855 6.820 ;
        RECT 6.255 5.290 6.425 6.900 ;
        RECT 7.135 6.820 8.185 6.990 ;
        RECT 7.135 5.290 7.305 6.820 ;
        RECT 4.245 5.120 4.895 5.290 ;
        RECT 6.255 5.120 7.305 5.290 ;
        RECT 7.575 5.290 7.745 6.560 ;
        RECT 8.015 5.550 8.185 6.820 ;
        RECT 7.575 5.120 8.225 5.290 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 4.355 3.905 4.525 4.865 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
        RECT 2.830 1.670 3.000 1.750 ;
        RECT 3.800 1.670 3.970 1.750 ;
        RECT 4.725 1.740 4.895 5.120 ;
        RECT 6.575 1.920 6.745 3.495 ;
        RECT 7.685 1.920 7.855 4.865 ;
        RECT 2.830 1.500 3.970 1.670 ;
        RECT 2.830 0.370 3.000 1.500 ;
        RECT 3.800 0.620 3.970 1.500 ;
        RECT 4.285 1.570 4.895 1.740 ;
        RECT 6.160 1.670 6.330 1.750 ;
        RECT 7.130 1.670 7.300 1.750 ;
        RECT 8.055 1.740 8.225 5.120 ;
        RECT 9.900 4.665 10.070 7.020 ;
        RECT 9.535 4.495 10.070 4.665 ;
        RECT 9.535 2.165 9.705 4.495 ;
        RECT 9.535 1.995 10.075 2.165 ;
        RECT 4.285 0.840 4.455 1.570 ;
        RECT 6.160 1.500 7.300 1.670 ;
        RECT 4.770 0.620 4.940 1.390 ;
        RECT 3.800 0.450 4.940 0.620 ;
        RECT 3.800 0.370 3.970 0.450 ;
        RECT 4.770 0.370 4.940 0.450 ;
        RECT 6.160 0.370 6.330 1.500 ;
        RECT 7.130 0.620 7.300 1.500 ;
        RECT 7.615 1.570 8.225 1.740 ;
        RECT 7.615 0.840 7.785 1.570 ;
        RECT 8.100 0.620 8.270 1.390 ;
        RECT 9.905 0.840 10.075 1.995 ;
        RECT 11.755 1.920 11.925 4.865 ;
        RECT 12.130 4.665 12.300 7.020 ;
        RECT 14.025 5.290 14.195 6.900 ;
        RECT 14.905 6.820 15.955 6.990 ;
        RECT 14.905 5.290 15.075 6.820 ;
        RECT 15.785 5.550 15.955 6.820 ;
        RECT 14.025 5.120 15.075 5.290 ;
        RECT 17.355 5.290 17.525 6.900 ;
        RECT 18.235 6.820 19.285 6.990 ;
        RECT 18.235 5.290 18.405 6.820 ;
        RECT 19.115 5.550 19.285 6.820 ;
        RECT 17.355 5.120 18.405 5.290 ;
        RECT 12.130 4.495 12.665 4.665 ;
        RECT 12.495 2.165 12.665 4.495 ;
        RECT 12.125 1.995 12.665 2.165 ;
        RECT 12.125 0.840 12.295 1.995 ;
        RECT 14.345 1.920 14.515 4.865 ;
        RECT 15.455 3.905 15.625 4.865 ;
        RECT 17.675 1.920 17.845 3.495 ;
        RECT 18.785 1.920 18.955 4.865 ;
        RECT 21.000 4.665 21.170 7.020 ;
        RECT 23.345 5.285 23.515 7.020 ;
        RECT 24.225 5.285 24.395 7.020 ;
        RECT 23.345 5.115 24.875 5.285 ;
        RECT 23.995 4.710 24.165 4.865 ;
        RECT 20.635 4.495 21.170 4.665 ;
        RECT 23.965 4.535 24.165 4.710 ;
        RECT 20.635 2.165 20.805 4.495 ;
        RECT 20.635 1.995 21.175 2.165 ;
        RECT 13.930 1.670 14.100 1.750 ;
        RECT 14.900 1.670 15.070 1.750 ;
        RECT 13.930 1.500 15.070 1.670 ;
        RECT 7.130 0.450 8.270 0.620 ;
        RECT 7.130 0.370 7.300 0.450 ;
        RECT 8.100 0.370 8.270 0.450 ;
        RECT 13.930 0.370 14.100 1.500 ;
        RECT 14.900 0.620 15.070 1.500 ;
        RECT 17.260 1.670 17.430 1.750 ;
        RECT 18.230 1.670 18.400 1.750 ;
        RECT 17.260 1.500 18.400 1.670 ;
        RECT 15.870 0.620 16.040 1.390 ;
        RECT 14.900 0.450 16.040 0.620 ;
        RECT 14.900 0.370 15.070 0.450 ;
        RECT 15.870 0.370 16.040 0.450 ;
        RECT 17.260 0.370 17.430 1.500 ;
        RECT 18.230 0.620 18.400 1.500 ;
        RECT 19.200 0.620 19.370 1.390 ;
        RECT 21.005 0.840 21.175 1.995 ;
        RECT 23.965 1.915 24.135 4.535 ;
        RECT 22.810 1.665 22.980 1.745 ;
        RECT 23.780 1.665 23.950 1.745 ;
        RECT 24.705 1.740 24.875 5.115 ;
        RECT 26.185 1.920 26.355 4.865 ;
        RECT 26.560 4.665 26.730 7.020 ;
        RECT 28.895 5.285 29.065 7.020 ;
        RECT 29.775 5.285 29.945 7.020 ;
        RECT 28.895 5.115 30.425 5.285 ;
        RECT 26.560 4.495 27.095 4.665 ;
        RECT 26.925 2.165 27.095 4.495 ;
        RECT 26.555 1.995 27.095 2.165 ;
        RECT 22.810 1.495 23.950 1.665 ;
        RECT 18.230 0.450 19.370 0.620 ;
        RECT 18.230 0.370 18.400 0.450 ;
        RECT 19.200 0.370 19.370 0.450 ;
        RECT 22.810 0.365 22.980 1.495 ;
        RECT 23.780 0.615 23.950 1.495 ;
        RECT 24.265 1.570 24.875 1.740 ;
        RECT 24.265 0.835 24.435 1.570 ;
        RECT 24.750 0.615 24.920 1.385 ;
        RECT 26.555 0.840 26.725 1.995 ;
        RECT 28.360 1.665 28.530 1.745 ;
        RECT 29.330 1.665 29.500 1.745 ;
        RECT 30.255 1.740 30.425 5.115 ;
        RECT 31.735 1.920 31.905 4.865 ;
        RECT 32.110 4.665 32.280 7.020 ;
        RECT 34.005 5.295 34.175 7.025 ;
        RECT 34.885 6.825 35.935 6.995 ;
        RECT 34.885 5.295 35.055 6.825 ;
        RECT 34.005 5.125 35.055 5.295 ;
        RECT 35.325 5.295 35.495 6.565 ;
        RECT 35.765 5.555 35.935 6.825 ;
        RECT 35.325 5.125 35.975 5.295 ;
        RECT 34.170 4.710 34.340 4.870 ;
        RECT 35.100 4.710 35.270 4.870 ;
        RECT 32.110 4.495 32.645 4.665 ;
        RECT 34.170 4.540 34.495 4.710 ;
        RECT 32.475 2.165 32.645 4.495 ;
        RECT 32.105 1.995 32.645 2.165 ;
        RECT 28.360 1.495 29.500 1.665 ;
        RECT 23.780 0.445 24.920 0.615 ;
        RECT 23.780 0.365 23.950 0.445 ;
        RECT 24.750 0.365 24.920 0.445 ;
        RECT 28.360 0.365 28.530 1.495 ;
        RECT 29.330 0.615 29.500 1.495 ;
        RECT 29.815 1.570 30.425 1.740 ;
        RECT 29.815 0.835 29.985 1.570 ;
        RECT 30.300 0.615 30.470 1.385 ;
        RECT 32.105 0.840 32.275 1.995 ;
        RECT 34.325 1.915 34.495 4.540 ;
        RECT 35.065 4.540 35.270 4.710 ;
        RECT 35.065 1.915 35.235 4.540 ;
        RECT 35.805 1.740 35.975 5.125 ;
        RECT 37.285 1.920 37.455 4.865 ;
        RECT 34.395 1.570 35.975 1.740 ;
        RECT 34.395 0.835 34.565 1.570 ;
        RECT 35.365 0.835 35.535 1.570 ;
        RECT 29.330 0.445 30.470 0.615 ;
        RECT 29.330 0.365 29.500 0.445 ;
        RECT 30.300 0.365 30.470 0.445 ;
      LAYER mcon ;
        RECT 4.355 3.985 4.525 4.155 ;
        RECT 1.395 2.505 1.565 2.675 ;
        RECT 4.725 3.615 4.895 3.785 ;
        RECT 6.575 3.245 6.745 3.415 ;
        RECT 7.685 2.505 7.855 2.675 ;
        RECT 8.055 3.615 8.225 3.785 ;
        RECT 9.535 3.985 9.705 4.155 ;
        RECT 9.535 3.245 9.705 3.415 ;
        RECT 11.755 3.985 11.925 4.155 ;
        RECT 11.755 3.615 11.925 3.785 ;
        RECT 11.755 2.135 11.925 2.305 ;
        RECT 12.495 2.505 12.665 2.675 ;
        RECT 14.345 3.985 14.515 4.155 ;
        RECT 15.455 3.985 15.625 4.155 ;
        RECT 17.675 3.245 17.845 3.415 ;
        RECT 18.785 2.505 18.955 2.675 ;
        RECT 20.635 3.985 20.805 4.155 ;
        RECT 20.635 3.245 20.805 3.415 ;
        RECT 23.965 2.135 24.135 2.305 ;
        RECT 24.705 3.245 24.875 3.415 ;
        RECT 26.185 3.245 26.355 3.415 ;
        RECT 26.925 2.875 27.095 3.045 ;
        RECT 30.255 3.245 30.425 3.415 ;
        RECT 31.735 3.245 31.905 3.415 ;
        RECT 32.475 3.245 32.645 3.415 ;
        RECT 34.325 2.875 34.495 3.045 ;
        RECT 35.065 3.245 35.235 3.415 ;
        RECT 35.805 3.245 35.975 3.415 ;
        RECT 37.285 3.245 37.455 3.415 ;
      LAYER met1 ;
        RECT 4.325 4.155 4.555 4.185 ;
        RECT 9.505 4.155 9.735 4.185 ;
        RECT 11.725 4.155 11.955 4.185 ;
        RECT 14.315 4.155 14.545 4.185 ;
        RECT 15.425 4.155 15.655 4.185 ;
        RECT 20.605 4.155 20.835 4.185 ;
        RECT 4.295 3.985 9.765 4.155 ;
        RECT 11.695 3.985 14.575 4.155 ;
        RECT 15.395 3.985 20.865 4.155 ;
        RECT 4.325 3.955 4.555 3.985 ;
        RECT 9.505 3.955 9.735 3.985 ;
        RECT 11.725 3.955 11.955 3.985 ;
        RECT 14.315 3.955 14.545 3.985 ;
        RECT 15.425 3.955 15.655 3.985 ;
        RECT 20.605 3.955 20.835 3.985 ;
        RECT 4.695 3.785 4.925 3.815 ;
        RECT 8.025 3.785 8.255 3.815 ;
        RECT 11.725 3.785 11.955 3.815 ;
        RECT 4.665 3.615 11.985 3.785 ;
        RECT 4.695 3.585 4.925 3.615 ;
        RECT 8.025 3.585 8.255 3.615 ;
        RECT 11.725 3.585 11.955 3.615 ;
        RECT 6.545 3.415 6.775 3.445 ;
        RECT 9.505 3.415 9.735 3.445 ;
        RECT 17.645 3.415 17.875 3.445 ;
        RECT 20.605 3.415 20.835 3.445 ;
        RECT 24.675 3.415 24.905 3.445 ;
        RECT 26.155 3.415 26.385 3.445 ;
        RECT 30.225 3.415 30.455 3.445 ;
        RECT 31.705 3.415 31.935 3.445 ;
        RECT 32.445 3.415 32.675 3.445 ;
        RECT 35.035 3.415 35.265 3.445 ;
        RECT 35.775 3.415 36.005 3.445 ;
        RECT 37.255 3.415 37.485 3.445 ;
        RECT 6.515 3.245 9.765 3.415 ;
        RECT 17.615 3.245 20.865 3.415 ;
        RECT 24.645 3.245 26.415 3.415 ;
        RECT 30.195 3.245 31.965 3.415 ;
        RECT 32.415 3.245 35.295 3.415 ;
        RECT 35.745 3.245 37.515 3.415 ;
        RECT 6.545 3.215 6.775 3.245 ;
        RECT 9.505 3.215 9.735 3.245 ;
        RECT 17.645 3.215 17.875 3.245 ;
        RECT 20.605 3.215 20.835 3.245 ;
        RECT 24.675 3.215 24.905 3.245 ;
        RECT 26.155 3.215 26.385 3.245 ;
        RECT 30.225 3.215 30.455 3.245 ;
        RECT 31.705 3.215 31.935 3.245 ;
        RECT 32.445 3.215 32.675 3.245 ;
        RECT 35.035 3.215 35.265 3.245 ;
        RECT 35.775 3.215 36.005 3.245 ;
        RECT 37.255 3.215 37.485 3.245 ;
        RECT 26.895 3.045 27.125 3.075 ;
        RECT 34.295 3.045 34.525 3.075 ;
        RECT 26.865 2.875 34.555 3.045 ;
        RECT 26.895 2.845 27.125 2.875 ;
        RECT 34.295 2.845 34.525 2.875 ;
        RECT 1.365 2.675 1.595 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 12.465 2.675 12.695 2.705 ;
        RECT 18.755 2.675 18.985 2.705 ;
        RECT 1.335 2.505 7.915 2.675 ;
        RECT 12.435 2.505 19.015 2.675 ;
        RECT 1.365 2.475 1.595 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
        RECT 12.465 2.475 12.695 2.505 ;
        RECT 18.755 2.475 18.985 2.505 ;
        RECT 11.725 2.305 11.955 2.335 ;
        RECT 23.935 2.305 24.165 2.335 ;
        RECT 11.695 2.135 24.195 2.305 ;
        RECT 11.725 2.105 11.955 2.135 ;
        RECT 23.935 2.105 24.165 2.135 ;
  END
END FA
END LIBRARY

