* SPICE3 file created from AO3X1.ext - technology: sky130A

.subckt AO3X1 Y A B C VDD GND
M1000 a_864_209.t3 C.t0 a_797_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 GND A.t1 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=3.2565p pd=22.61u as=0p ps=0u
M1002 VDD.t5 a_217_1050.t5 a_797_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t2 A.t0 a_217_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD.t7 a_864_209.t4 Y.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD.t0 B.t0 a_217_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_217_1050.t4 A.t2 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_797_1051.t2 C.t1 a_864_209.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y.t1 a_864_209.t5 VDD.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_864_209.t6 GND.t3 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1010 a_797_1051.t1 a_217_1050.t7 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_217_1050.t1 B.t2 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD B 0.07fF
C1 A B 0.27fF
C2 VDD C 0.07fF
C3 VDD Y 0.76fF
C4 VDD A 0.08fF
R0 C.n0 C.t1 470.752
R1 C.n0 C.t0 384.527
R2 C.n1 C.t2 241.172
R3 C.n1 C.n0 110.173
R4 C.n2 C.n1 76
R5 C.n2 C 0.046
R6 a_797_1051.t0 a_797_1051.n0 101.66
R7 a_797_1051.n0 a_797_1051.t2 101.659
R8 a_797_1051.n0 a_797_1051.t3 14.294
R9 a_797_1051.n0 a_797_1051.t1 14.282
R10 a_864_209.n0 a_864_209.t4 512.525
R11 a_864_209.n0 a_864_209.t5 371.139
R12 a_864_209.n10 a_864_209.n9 244.994
R13 a_864_209.n1 a_864_209.n0 226.306
R14 a_864_209.n1 a_864_209.t6 157.328
R15 a_864_209.n9 a_864_209.n1 153.043
R16 a_864_209.n8 a_864_209.n7 133.539
R17 a_864_209.n9 a_864_209.n8 82.528
R18 a_864_209.n4 a_864_209.n2 80.526
R19 a_864_209.n8 a_864_209.n4 48.405
R20 a_864_209.n4 a_864_209.n3 30
R21 a_864_209.n7 a_864_209.n6 22.578
R22 a_864_209.n10 a_864_209.t2 14.282
R23 a_864_209.t3 a_864_209.n10 14.282
R24 a_864_209.n7 a_864_209.n5 8.58
R25 a_217_1050.n4 a_217_1050.t7 486.819
R26 a_217_1050.n4 a_217_1050.t5 384.527
R27 a_217_1050.n6 a_217_1050.n3 232.158
R28 a_217_1050.n5 a_217_1050.t6 197.395
R29 a_217_1050.n5 a_217_1050.n4 186.206
R30 a_217_1050.n6 a_217_1050.n5 153.315
R31 a_217_1050.n8 a_217_1050.n6 130.933
R32 a_217_1050.n3 a_217_1050.n2 76.002
R33 a_217_1050.n8 a_217_1050.n7 30
R34 a_217_1050.n9 a_217_1050.n0 24.383
R35 a_217_1050.n9 a_217_1050.n8 23.684
R36 a_217_1050.n1 a_217_1050.t0 14.282
R37 a_217_1050.n1 a_217_1050.t1 14.282
R38 a_217_1050.n2 a_217_1050.t3 14.282
R39 a_217_1050.n2 a_217_1050.t4 14.282
R40 a_217_1050.n3 a_217_1050.n1 12.85
R41 VDD.n68 VDD.n66 144.705
R42 VDD.n170 VDD.n168 144.705
R43 VDD.n26 VDD.n25 77.792
R44 VDD.n35 VDD.n34 77.792
R45 VDD.n29 VDD.n23 76.145
R46 VDD.n29 VDD.n28 76
R47 VDD.n33 VDD.n32 76
R48 VDD.n39 VDD.n38 76
R49 VDD.n43 VDD.n42 76
R50 VDD.n70 VDD.n69 76
R51 VDD.n74 VDD.n73 76
R52 VDD.n78 VDD.n77 76
R53 VDD.n82 VDD.n81 76
R54 VDD.n87 VDD.n86 76
R55 VDD.n183 VDD.n182 76
R56 VDD.n176 VDD.n175 76
R57 VDD.n172 VDD.n171 76
R58 VDD.n145 VDD.n144 76
R59 VDD.n141 VDD.n140 76
R60 VDD.n136 VDD.n135 76
R61 VDD.n131 VDD.n130 76
R62 VDD.n125 VDD.n124 76
R63 VDD.n120 VDD.n119 76
R64 VDD.n115 VDD.n114 76
R65 VDD.n110 VDD.n109 76
R66 VDD.n111 VDD.t3 55.106
R67 VDD.n37 VDD.t6 55.106
R68 VDD.n24 VDD.t7 55.106
R69 VDD.n137 VDD.t0 55.106
R70 VDD.n178 VDD.n177 41.183
R71 VDD.n127 VDD.n126 40.824
R72 VDD.n48 VDD.n47 36.774
R73 VDD.n161 VDD.n160 36.774
R74 VDD.n133 VDD.n132 36.608
R75 VDD.n180 VDD.n179 32.032
R76 VDD.n117 VDD.n116 32.032
R77 VDD.n109 VDD.n106 21.841
R78 VDD.n23 VDD.n20 21.841
R79 VDD.n126 VDD.t1 14.282
R80 VDD.n126 VDD.t2 14.282
R81 VDD.n177 VDD.t4 14.282
R82 VDD.n177 VDD.t5 14.282
R83 VDD.n106 VDD.n89 14.167
R84 VDD.n89 VDD.n88 14.167
R85 VDD.n64 VDD.n45 14.167
R86 VDD.n45 VDD.n44 14.167
R87 VDD.n166 VDD.n147 14.167
R88 VDD.n147 VDD.n146 14.167
R89 VDD.n20 VDD.n19 14.167
R90 VDD.n19 VDD.n17 14.167
R91 VDD.n69 VDD.n65 14.167
R92 VDD.n171 VDD.n167 14.167
R93 VDD.n23 VDD.n22 13.653
R94 VDD.n22 VDD.n21 13.653
R95 VDD.n28 VDD.n27 13.653
R96 VDD.n27 VDD.n26 13.653
R97 VDD.n32 VDD.n31 13.653
R98 VDD.n31 VDD.n30 13.653
R99 VDD.n38 VDD.n36 13.653
R100 VDD.n36 VDD.n35 13.653
R101 VDD.n42 VDD.n41 13.653
R102 VDD.n41 VDD.n40 13.653
R103 VDD.n69 VDD.n68 13.653
R104 VDD.n68 VDD.n67 13.653
R105 VDD.n73 VDD.n72 13.653
R106 VDD.n72 VDD.n71 13.653
R107 VDD.n77 VDD.n76 13.653
R108 VDD.n76 VDD.n75 13.653
R109 VDD.n81 VDD.n80 13.653
R110 VDD.n80 VDD.n79 13.653
R111 VDD.n86 VDD.n85 13.653
R112 VDD.n85 VDD.n84 13.653
R113 VDD.n182 VDD.n181 13.653
R114 VDD.n181 VDD.n180 13.653
R115 VDD.n175 VDD.n174 13.653
R116 VDD.n174 VDD.n173 13.653
R117 VDD.n171 VDD.n170 13.653
R118 VDD.n170 VDD.n169 13.653
R119 VDD.n144 VDD.n143 13.653
R120 VDD.n143 VDD.n142 13.653
R121 VDD.n140 VDD.n139 13.653
R122 VDD.n139 VDD.n138 13.653
R123 VDD.n135 VDD.n134 13.653
R124 VDD.n134 VDD.n133 13.653
R125 VDD.n130 VDD.n129 13.653
R126 VDD.n129 VDD.n128 13.653
R127 VDD.n124 VDD.n123 13.653
R128 VDD.n123 VDD.n122 13.653
R129 VDD.n119 VDD.n118 13.653
R130 VDD.n118 VDD.n117 13.653
R131 VDD.n114 VDD.n113 13.653
R132 VDD.n113 VDD.n112 13.653
R133 VDD.n109 VDD.n108 13.653
R134 VDD.n108 VDD.n107 13.653
R135 VDD.n4 VDD.n2 12.915
R136 VDD.n4 VDD.n3 12.66
R137 VDD.n12 VDD.n11 12.343
R138 VDD.n8 VDD.n7 12.343
R139 VDD.n12 VDD.n9 12.343
R140 VDD.n130 VDD.n127 8.658
R141 VDD.n65 VDD.n64 7.674
R142 VDD.n167 VDD.n166 7.674
R143 VDD.n59 VDD.n58 7.5
R144 VDD.n53 VDD.n52 7.5
R145 VDD.n55 VDD.n54 7.5
R146 VDD.n50 VDD.n49 7.5
R147 VDD.n64 VDD.n63 7.5
R148 VDD.n151 VDD.n150 7.5
R149 VDD.n154 VDD.n153 7.5
R150 VDD.n156 VDD.n155 7.5
R151 VDD.n159 VDD.n158 7.5
R152 VDD.n166 VDD.n165 7.5
R153 VDD.n101 VDD.n100 7.5
R154 VDD.n95 VDD.n94 7.5
R155 VDD.n97 VDD.n96 7.5
R156 VDD.n103 VDD.n93 7.5
R157 VDD.n103 VDD.n91 7.5
R158 VDD.n106 VDD.n105 7.5
R159 VDD.n20 VDD.n16 7.5
R160 VDD.n2 VDD.n1 7.5
R161 VDD.n7 VDD.n6 7.5
R162 VDD.n11 VDD.n10 7.5
R163 VDD.n19 VDD.n18 7.5
R164 VDD.n14 VDD.n0 7.5
R165 VDD.n51 VDD.n48 6.772
R166 VDD.n62 VDD.n46 6.772
R167 VDD.n60 VDD.n57 6.772
R168 VDD.n56 VDD.n53 6.772
R169 VDD.n104 VDD.n90 6.772
R170 VDD.n102 VDD.n99 6.772
R171 VDD.n98 VDD.n95 6.772
R172 VDD.n51 VDD.n50 6.772
R173 VDD.n56 VDD.n55 6.772
R174 VDD.n60 VDD.n59 6.772
R175 VDD.n63 VDD.n62 6.772
R176 VDD.n98 VDD.n97 6.772
R177 VDD.n102 VDD.n101 6.772
R178 VDD.n105 VDD.n104 6.772
R179 VDD.n165 VDD.n164 6.772
R180 VDD.n152 VDD.n149 6.772
R181 VDD.n157 VDD.n154 6.772
R182 VDD.n162 VDD.n159 6.772
R183 VDD.n162 VDD.n161 6.772
R184 VDD.n157 VDD.n156 6.772
R185 VDD.n152 VDD.n151 6.772
R186 VDD.n164 VDD.n148 6.772
R187 VDD.n16 VDD.n15 6.458
R188 VDD.n93 VDD.n92 6.202
R189 VDD.n182 VDD.n178 5.903
R190 VDD.n84 VDD.n83 4.576
R191 VDD.n122 VDD.n121 4.576
R192 VDD.n114 VDD.n111 2.754
R193 VDD.n140 VDD.n137 2.361
R194 VDD.n28 VDD.n24 1.967
R195 VDD.n38 VDD.n37 1.967
R196 VDD.n14 VDD.n5 1.329
R197 VDD.n14 VDD.n8 1.329
R198 VDD.n14 VDD.n12 1.329
R199 VDD.n14 VDD.n13 1.329
R200 VDD.n15 VDD.n14 0.696
R201 VDD.n14 VDD.n4 0.696
R202 VDD.n61 VDD.n60 0.365
R203 VDD.n61 VDD.n56 0.365
R204 VDD.n61 VDD.n51 0.365
R205 VDD.n62 VDD.n61 0.365
R206 VDD.n103 VDD.n102 0.365
R207 VDD.n103 VDD.n98 0.365
R208 VDD.n104 VDD.n103 0.365
R209 VDD.n163 VDD.n162 0.365
R210 VDD.n163 VDD.n157 0.365
R211 VDD.n163 VDD.n152 0.365
R212 VDD.n164 VDD.n163 0.365
R213 VDD.n70 VDD.n43 0.29
R214 VDD.n172 VDD.n145 0.29
R215 VDD.n110 VDD 0.207
R216 VDD.n87 VDD.n82 0.181
R217 VDD.n131 VDD.n125 0.181
R218 VDD.n33 VDD.n29 0.157
R219 VDD.n39 VDD.n33 0.157
R220 VDD.n43 VDD.n39 0.145
R221 VDD.n74 VDD.n70 0.145
R222 VDD.n78 VDD.n74 0.145
R223 VDD.n82 VDD.n78 0.145
R224 VDD.n183 VDD.n176 0.145
R225 VDD.n176 VDD.n172 0.145
R226 VDD.n145 VDD.n141 0.145
R227 VDD.n141 VDD.n136 0.145
R228 VDD.n136 VDD.n131 0.145
R229 VDD.n125 VDD.n120 0.145
R230 VDD.n120 VDD.n115 0.145
R231 VDD.n115 VDD.n110 0.145
R232 VDD VDD.n87 0.133
R233 VDD VDD.n183 0.012
R234 A.n0 A.t0 480.392
R235 A.n0 A.t2 403.272
R236 A.n1 A.t1 230.374
R237 A.n1 A.n0 151.553
R238 A.n2 A.n1 76
R239 A.n2 A 0.046
R240 Y.n5 Y.n4 232.121
R241 Y.n5 Y.n0 130.901
R242 Y.n6 Y.n5 76
R243 Y.n4 Y.n3 30
R244 Y.n2 Y.n1 24.383
R245 Y.n4 Y.n2 23.684
R246 Y.n0 Y.t2 14.282
R247 Y.n0 Y.t1 14.282
R248 Y.n6 Y 0.046
R249 GND.n30 GND.n28 219.745
R250 GND.n89 GND.n88 219.745
R251 GND.n30 GND.n29 85.529
R252 GND.n89 GND.n87 85.529
R253 GND.n9 GND.n1 76.145
R254 GND.n59 GND.n58 76
R255 GND.n9 GND.n8 76
R256 GND.n17 GND.n16 76
R257 GND.n24 GND.n23 76
R258 GND.n27 GND.n26 76
R259 GND.n34 GND.n33 76
R260 GND.n41 GND.n40 76
R261 GND.n47 GND.n46 76
R262 GND.n50 GND.n49 76
R263 GND.n56 GND.n55 76
R264 GND.n104 GND.n103 76
R265 GND.n99 GND.n98 76
R266 GND.n92 GND.n91 76
R267 GND.n85 GND.n84 76
R268 GND.n82 GND.n81 76
R269 GND.n79 GND.n78 76
R270 GND.n76 GND.n75 76
R271 GND.n73 GND.n72 76
R272 GND.n70 GND.n69 76
R273 GND.n62 GND.n61 76
R274 GND.n67 GND.n66 63.835
R275 GND.n5 GND.n4 35.01
R276 GND.n3 GND.n2 29.127
R277 GND.n66 GND.n65 28.421
R278 GND.n66 GND.n64 25.263
R279 GND.n64 GND.n63 24.383
R280 GND.n12 GND.t3 20.794
R281 GND.n6 GND.n5 19.735
R282 GND.n14 GND.n13 19.735
R283 GND.n22 GND.n21 19.735
R284 GND.n101 GND.n100 19.735
R285 GND.n53 GND.n52 19.735
R286 GND.n45 GND.n44 19.735
R287 GND.n38 GND.n37 19.735
R288 GND.n97 GND.n96 19.735
R289 GND.n44 GND.t2 19.724
R290 GND.n100 GND.t1 19.724
R291 GND.n5 GND.n3 19.017
R292 GND.n33 GND.n31 14.167
R293 GND.n91 GND.n90 14.167
R294 GND.n61 GND.n60 13.653
R295 GND.n69 GND.n68 13.653
R296 GND.n72 GND.n71 13.653
R297 GND.n75 GND.n74 13.653
R298 GND.n78 GND.n77 13.653
R299 GND.n81 GND.n80 13.653
R300 GND.n84 GND.n83 13.653
R301 GND.n91 GND.n86 13.653
R302 GND.n98 GND.n93 13.653
R303 GND.n103 GND.n102 13.653
R304 GND.n55 GND.n54 13.653
R305 GND.n49 GND.n48 13.653
R306 GND.n46 GND.n42 13.653
R307 GND.n40 GND.n39 13.653
R308 GND.n33 GND.n32 13.653
R309 GND.n26 GND.n25 13.653
R310 GND.n23 GND.n18 13.653
R311 GND.n16 GND.n15 13.653
R312 GND.n8 GND.n7 13.653
R313 GND.n21 GND.n20 12.837
R314 GND.n96 GND.n95 12.837
R315 GND.n37 GND.n36 11.605
R316 GND.n36 GND.n35 9.809
R317 GND.n55 GND.n53 8.854
R318 GND.n20 GND.n19 7.566
R319 GND.n95 GND.n94 7.566
R320 GND.n31 GND.n30 7.312
R321 GND.n90 GND.n89 7.312
R322 GND.t2 GND.n43 7.04
R323 GND.n52 GND.n51 5.774
R324 GND.n11 GND.n10 4.551
R325 GND.n8 GND.n6 3.935
R326 GND.n46 GND.n45 3.935
R327 GND.n103 GND.n101 3.935
R328 GND.n69 GND.n67 3.935
R329 GND.n23 GND.n22 3.541
R330 GND.t3 GND.n11 2.238
R331 GND.n40 GND.n38 0.983
R332 GND.n98 GND.n97 0.983
R333 GND.n1 GND.n0 0.596
R334 GND.n58 GND.n57 0.596
R335 GND.n13 GND.n12 0.358
R336 GND.n34 GND.n27 0.29
R337 GND.n92 GND.n85 0.29
R338 GND.n59 GND 0.207
R339 GND.n16 GND.n14 0.196
R340 GND.n56 GND.n50 0.181
R341 GND.n76 GND.n73 0.181
R342 GND.n17 GND.n9 0.157
R343 GND.n24 GND.n17 0.157
R344 GND.n27 GND.n24 0.145
R345 GND.n41 GND.n34 0.145
R346 GND.n47 GND.n41 0.145
R347 GND.n50 GND.n47 0.145
R348 GND.n104 GND.n99 0.145
R349 GND.n99 GND.n92 0.145
R350 GND.n85 GND.n82 0.145
R351 GND.n82 GND.n79 0.145
R352 GND.n79 GND.n76 0.145
R353 GND.n73 GND.n70 0.145
R354 GND.n70 GND.n62 0.145
R355 GND.n62 GND.n59 0.145
R356 GND GND.n56 0.133
R357 GND GND.n104 0.012
R358 a_112_101.n12 a_112_101.n11 26.811
R359 a_112_101.n6 a_112_101.n5 24.977
R360 a_112_101.n2 a_112_101.n1 24.877
R361 a_112_101.t0 a_112_101.n2 12.677
R362 a_112_101.t0 a_112_101.n3 11.595
R363 a_112_101.t1 a_112_101.n8 8.137
R364 a_112_101.t0 a_112_101.n4 7.273
R365 a_112_101.t0 a_112_101.n0 6.109
R366 a_112_101.t1 a_112_101.n7 4.864
R367 a_112_101.t0 a_112_101.n12 2.074
R368 a_112_101.n7 a_112_101.n6 1.13
R369 a_112_101.n12 a_112_101.t1 0.937
R370 a_112_101.t1 a_112_101.n10 0.804
R371 a_112_101.n10 a_112_101.n9 0.136
R372 B.n0 B.t0 472.359
R373 B.n0 B.t2 384.527
R374 B.n1 B.t1 214.619
R375 B.n1 B.n0 136.613
R376 B.n2 B.n1 76
R377 B.n2 B 0.046
C5 VDD GND 7.42fF
C6 a_112_101.n0 GND 0.02fF
C7 a_112_101.n1 GND 0.10fF
C8 a_112_101.n2 GND 0.06fF
C9 a_112_101.n3 GND 0.06fF
C10 a_112_101.n4 GND 0.00fF
C11 a_112_101.n5 GND 0.04fF
C12 a_112_101.n6 GND 0.05fF
C13 a_112_101.n7 GND 0.02fF
C14 a_112_101.n8 GND 0.05fF
C15 a_112_101.n9 GND 0.07fF
C16 a_112_101.n10 GND 0.17fF
C17 a_112_101.t1 GND 0.22fF
C18 a_112_101.n11 GND 0.09fF
C19 a_112_101.n12 GND 0.00fF
C20 Y.n0 GND 0.74fF
C21 Y.n1 GND 0.04fF
C22 Y.n2 GND 0.06fF
C23 Y.n3 GND 0.04fF
C24 Y.n4 GND 0.34fF
C25 Y.n5 GND 0.47fF
C26 Y.n6 GND 0.01fF
C27 VDD.n0 GND 0.11fF
C28 VDD.n1 GND 0.02fF
C29 VDD.n2 GND 0.02fF
C30 VDD.n3 GND 0.04fF
C31 VDD.n4 GND 0.01fF
C32 VDD.n6 GND 0.02fF
C33 VDD.n7 GND 0.02fF
C34 VDD.n9 GND 0.02fF
C35 VDD.n10 GND 0.02fF
C36 VDD.n11 GND 0.02fF
C37 VDD.n14 GND 0.42fF
C38 VDD.n16 GND 0.03fF
C39 VDD.n17 GND 0.02fF
C40 VDD.n18 GND 0.02fF
C41 VDD.n19 GND 0.02fF
C42 VDD.n20 GND 0.03fF
C43 VDD.n21 GND 0.25fF
C44 VDD.n22 GND 0.02fF
C45 VDD.n23 GND 0.03fF
C46 VDD.n24 GND 0.05fF
C47 VDD.n25 GND 0.14fF
C48 VDD.n26 GND 0.19fF
C49 VDD.n27 GND 0.01fF
C50 VDD.n28 GND 0.01fF
C51 VDD.n29 GND 0.06fF
C52 VDD.n30 GND 0.15fF
C53 VDD.n31 GND 0.01fF
C54 VDD.n32 GND 0.02fF
C55 VDD.n33 GND 0.02fF
C56 VDD.n34 GND 0.14fF
C57 VDD.n35 GND 0.19fF
C58 VDD.n36 GND 0.01fF
C59 VDD.n37 GND 0.06fF
C60 VDD.n38 GND 0.01fF
C61 VDD.n39 GND 0.02fF
C62 VDD.n40 GND 0.25fF
C63 VDD.n41 GND 0.01fF
C64 VDD.n42 GND 0.02fF
C65 VDD.n43 GND 0.03fF
C66 VDD.n44 GND 0.02fF
C67 VDD.n45 GND 0.02fF
C68 VDD.n46 GND 0.02fF
C69 VDD.n47 GND 0.17fF
C70 VDD.n48 GND 0.04fF
C71 VDD.n49 GND 0.03fF
C72 VDD.n50 GND 0.02fF
C73 VDD.n52 GND 0.02fF
C74 VDD.n53 GND 0.02fF
C75 VDD.n54 GND 0.02fF
C76 VDD.n55 GND 0.02fF
C77 VDD.n57 GND 0.02fF
C78 VDD.n58 GND 0.02fF
C79 VDD.n59 GND 0.02fF
C80 VDD.n61 GND 0.25fF
C81 VDD.n63 GND 0.02fF
C82 VDD.n64 GND 0.02fF
C83 VDD.n65 GND 0.03fF
C84 VDD.n66 GND 0.02fF
C85 VDD.n67 GND 0.25fF
C86 VDD.n68 GND 0.01fF
C87 VDD.n69 GND 0.02fF
C88 VDD.n70 GND 0.03fF
C89 VDD.n71 GND 0.25fF
C90 VDD.n72 GND 0.01fF
C91 VDD.n73 GND 0.02fF
C92 VDD.n74 GND 0.02fF
C93 VDD.n75 GND 0.25fF
C94 VDD.n76 GND 0.01fF
C95 VDD.n77 GND 0.02fF
C96 VDD.n78 GND 0.02fF
C97 VDD.n79 GND 0.28fF
C98 VDD.n80 GND 0.01fF
C99 VDD.n81 GND 0.02fF
C100 VDD.n82 GND 0.02fF
C101 VDD.n83 GND 0.16fF
C102 VDD.n84 GND 0.13fF
C103 VDD.n85 GND 0.01fF
C104 VDD.n86 GND 0.02fF
C105 VDD.n87 GND 0.02fF
C106 VDD.n88 GND 0.02fF
C107 VDD.n89 GND 0.02fF
C108 VDD.n90 GND 0.02fF
C109 VDD.n91 GND 0.14fF
C110 VDD.n92 GND 0.03fF
C111 VDD.n93 GND 0.02fF
C112 VDD.n94 GND 0.02fF
C113 VDD.n95 GND 0.02fF
C114 VDD.n96 GND 0.02fF
C115 VDD.n97 GND 0.02fF
C116 VDD.n99 GND 0.02fF
C117 VDD.n100 GND 0.02fF
C118 VDD.n101 GND 0.02fF
C119 VDD.n103 GND 0.42fF
C120 VDD.n105 GND 0.03fF
C121 VDD.n106 GND 0.03fF
C122 VDD.n107 GND 0.25fF
C123 VDD.n108 GND 0.02fF
C124 VDD.n109 GND 0.03fF
C125 VDD.n110 GND 0.03fF
C126 VDD.n111 GND 0.06fF
C127 VDD.n112 GND 0.23fF
C128 VDD.n113 GND 0.01fF
C129 VDD.n114 GND 0.01fF
C130 VDD.n115 GND 0.02fF
C131 VDD.n116 GND 0.13fF
C132 VDD.n117 GND 0.15fF
C133 VDD.n118 GND 0.01fF
C134 VDD.n119 GND 0.02fF
C135 VDD.n120 GND 0.02fF
C136 VDD.n121 GND 0.16fF
C137 VDD.n122 GND 0.13fF
C138 VDD.n123 GND 0.01fF
C139 VDD.n124 GND 0.02fF
C140 VDD.n125 GND 0.02fF
C141 VDD.n126 GND 0.10fF
C142 VDD.n127 GND 0.02fF
C143 VDD.n128 GND 0.28fF
C144 VDD.n129 GND 0.01fF
C145 VDD.n130 GND 0.02fF
C146 VDD.n131 GND 0.02fF
C147 VDD.n132 GND 0.13fF
C148 VDD.n133 GND 0.15fF
C149 VDD.n134 GND 0.01fF
C150 VDD.n135 GND 0.02fF
C151 VDD.n136 GND 0.02fF
C152 VDD.n137 GND 0.05fF
C153 VDD.n138 GND 0.23fF
C154 VDD.n139 GND 0.01fF
C155 VDD.n140 GND 0.01fF
C156 VDD.n141 GND 0.02fF
C157 VDD.n142 GND 0.25fF
C158 VDD.n143 GND 0.01fF
C159 VDD.n144 GND 0.02fF
C160 VDD.n145 GND 0.03fF
C161 VDD.n146 GND 0.02fF
C162 VDD.n147 GND 0.02fF
C163 VDD.n148 GND 0.02fF
C164 VDD.n149 GND 0.02fF
C165 VDD.n150 GND 0.02fF
C166 VDD.n151 GND 0.02fF
C167 VDD.n153 GND 0.02fF
C168 VDD.n154 GND 0.02fF
C169 VDD.n155 GND 0.02fF
C170 VDD.n156 GND 0.02fF
C171 VDD.n158 GND 0.03fF
C172 VDD.n159 GND 0.02fF
C173 VDD.n160 GND 0.20fF
C174 VDD.n161 GND 0.04fF
C175 VDD.n163 GND 0.25fF
C176 VDD.n165 GND 0.02fF
C177 VDD.n166 GND 0.02fF
C178 VDD.n167 GND 0.03fF
C179 VDD.n168 GND 0.02fF
C180 VDD.n169 GND 0.25fF
C181 VDD.n170 GND 0.01fF
C182 VDD.n171 GND 0.02fF
C183 VDD.n172 GND 0.03fF
C184 VDD.n173 GND 0.23fF
C185 VDD.n174 GND 0.01fF
C186 VDD.n175 GND 0.02fF
C187 VDD.n176 GND 0.02fF
C188 VDD.n177 GND 0.10fF
C189 VDD.n178 GND 0.02fF
C190 VDD.n179 GND 0.13fF
C191 VDD.n180 GND 0.15fF
C192 VDD.n181 GND 0.01fF
C193 VDD.n182 GND 0.01fF
C194 VDD.n183 GND 0.01fF
C195 a_217_1050.n0 GND 0.03fF
C196 a_217_1050.n1 GND 0.42fF
C197 a_217_1050.n2 GND 0.50fF
C198 a_217_1050.n3 GND 0.32fF
C199 a_217_1050.n4 GND 0.36fF
C200 a_217_1050.t6 GND 0.37fF
C201 a_217_1050.n5 GND 0.45fF
C202 a_217_1050.n6 GND 0.48fF
C203 a_217_1050.n7 GND 0.03fF
C204 a_217_1050.n8 GND 0.16fF
C205 a_217_1050.n9 GND 0.04fF
C206 a_864_209.n0 GND 0.36fF
C207 a_864_209.n1 GND 0.47fF
C208 a_864_209.n2 GND 0.05fF
C209 a_864_209.n3 GND 0.03fF
C210 a_864_209.n4 GND 0.10fF
C211 a_864_209.n5 GND 0.04fF
C212 a_864_209.n6 GND 0.04fF
C213 a_864_209.n7 GND 0.16fF
C214 a_864_209.n8 GND 0.27fF
C215 a_864_209.n9 GND 0.44fF
C216 a_864_209.n10 GND 0.63fF
C217 a_797_1051.n0 GND 0.54fF
.ends
