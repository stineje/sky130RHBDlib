* SPICE3 file created from AOA4X1.ext - technology: sky130A

.subckt AOA4X1 Y A B C D VPB VNB
X0 a_864_181# a_217_1004# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.4356e+12p ps=2.418e+07u w=3e+06u l=150000u
X1 VPB a_343_383# a_217_1004# VPB sky130_fd_pr__pfet_01v8 ad=5.04e+12p pd=4.104e+07u as=0p ps=0u w=2e+06u l=150000u M=2
X2 VNB a_168_157# a_112_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 VNB a_864_181# a_1444_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4 VPB a_864_181# a_1549_1004# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X5 a_1549_1004# a_1675_383# a_1444_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X6 VPB a_1549_1004# a_2183_182# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X7 a_797_1005# a_1009_383# a_864_181# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X8 a_217_1004# a_168_157# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X9 a_217_1004# a_343_383# a_112_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X10 VPB a_1675_383# a_1549_1004# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X11 a_864_181# a_1009_383# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X12 a_797_1005# a_217_1004# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X13 a_2183_182# a_1549_1004# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends
