* SPICE3 file created from TIELO.ext - technology: sky130A

.subckt TIELO YN VDD GND
M1000 a_121_411.t1 a_121_411.t0 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VDD.t0 a_121_411.t2 a_121_411.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 YN a_121_411.t4 GND.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
R0 a_121_411.n0 a_121_411.t2 512.525
R1 a_121_411.n0 a_121_411.t0 371.139
R2 a_121_411.n1 a_121_411.t4 319.158
R3 a_121_411.n2 a_121_411.n1 75.63
R4 a_121_411.n1 a_121_411.n0 58.377
R5 a_121_411.n2 a_121_411.t3 14.282
R6 a_121_411.t1 a_121_411.n2 14.282
R7 GND.n9 GND.n1 76.145
R8 GND.n12 GND.n11 76
R9 GND.n9 GND.n8 76
R10 GND.n27 GND.n26 76
R11 GND.n21 GND.n20 76
R12 GND.n17 GND.t0 39.412
R13 GND.n5 GND.n4 35.01
R14 GND.n26 GND.n24 19.735
R15 GND.n6 GND.n5 19.735
R16 GND.n19 GND.n18 19.735
R17 GND.n5 GND.n3 19.017
R18 GND.n17 GND.n16 17.185
R19 GND.n20 GND.n13 13.653
R20 GND.n26 GND.n25 13.653
R21 GND.n8 GND.n7 13.653
R22 GND.n3 GND.n2 7.5
R23 GND.n24 GND.n23 7.5
R24 GND.n18 GND.n17 6.139
R25 GND.n15 GND.n14 4.551
R26 GND.n8 GND.n6 3.935
R27 GND.n20 GND.n19 3.541
R28 GND.t0 GND.n15 2.238
R29 GND.n23 GND.n22 1.935
R30 GND.n1 GND.n0 0.596
R31 GND.n11 GND.n10 0.596
R32 GND.n12 GND 0.207
R33 GND.n27 GND.n9 0.157
R34 GND.n27 GND.n21 0.157
R35 GND.n21 GND.n12 0.145
R36 YN.n1 YN.n0 235.85
R37 YN.n1 YN 0.046
R38 VDD.n26 VDD.n25 77.792
R39 VDD.n55 VDD.n54 77.792
R40 VDD.n29 VDD.n23 76.145
R41 VDD.n29 VDD.n28 76
R42 VDD.n63 VDD.n62 76
R43 VDD.n59 VDD.n58 76
R44 VDD.n53 VDD.n52 76
R45 VDD.n57 VDD.t1 55.106
R46 VDD.n24 VDD.t0 55.106
R47 VDD.n52 VDD.n49 21.841
R48 VDD.n23 VDD.n20 21.841
R49 VDD.n49 VDD.n31 14.167
R50 VDD.n31 VDD.n30 14.167
R51 VDD.n20 VDD.n19 14.167
R52 VDD.n19 VDD.n17 14.167
R53 VDD.n23 VDD.n22 13.653
R54 VDD.n22 VDD.n21 13.653
R55 VDD.n28 VDD.n27 13.653
R56 VDD.n27 VDD.n26 13.653
R57 VDD.n62 VDD.n61 13.653
R58 VDD.n61 VDD.n60 13.653
R59 VDD.n58 VDD.n56 13.653
R60 VDD.n56 VDD.n55 13.653
R61 VDD.n52 VDD.n51 13.653
R62 VDD.n51 VDD.n50 13.653
R63 VDD.n4 VDD.n2 12.915
R64 VDD.n4 VDD.n3 12.66
R65 VDD.n12 VDD.n11 12.343
R66 VDD.n10 VDD.n9 12.343
R67 VDD.n7 VDD.n6 12.343
R68 VDD.n35 VDD.n34 7.5
R69 VDD.n38 VDD.n37 7.5
R70 VDD.n40 VDD.n39 7.5
R71 VDD.n43 VDD.n42 7.5
R72 VDD.n49 VDD.n48 7.5
R73 VDD.n20 VDD.n16 7.5
R74 VDD.n2 VDD.n1 7.5
R75 VDD.n6 VDD.n5 7.5
R76 VDD.n9 VDD.n8 7.5
R77 VDD.n19 VDD.n18 7.5
R78 VDD.n14 VDD.n0 7.5
R79 VDD.n48 VDD.n47 6.772
R80 VDD.n36 VDD.n33 6.772
R81 VDD.n41 VDD.n38 6.772
R82 VDD.n45 VDD.n43 6.772
R83 VDD.n45 VDD.n44 6.772
R84 VDD.n41 VDD.n40 6.772
R85 VDD.n36 VDD.n35 6.772
R86 VDD.n47 VDD.n32 6.772
R87 VDD.n16 VDD.n15 6.458
R88 VDD.n28 VDD.n24 1.967
R89 VDD.n58 VDD.n57 1.967
R90 VDD.n14 VDD.n7 1.329
R91 VDD.n14 VDD.n10 1.329
R92 VDD.n14 VDD.n12 1.329
R93 VDD.n14 VDD.n13 1.329
R94 VDD.n15 VDD.n14 0.696
R95 VDD.n14 VDD.n4 0.696
R96 VDD.n46 VDD.n45 0.365
R97 VDD.n46 VDD.n41 0.365
R98 VDD.n46 VDD.n36 0.365
R99 VDD.n47 VDD.n46 0.365
R100 VDD.n53 VDD 0.207
R101 VDD.n63 VDD.n29 0.157
R102 VDD.n63 VDD.n59 0.157
R103 VDD.n59 VDD.n53 0.145
C0 VDD GND 2.55fF
C1 VDD.n0 GND 0.10fF
C2 VDD.n1 GND 0.02fF
C3 VDD.n2 GND 0.02fF
C4 VDD.n3 GND 0.04fF
C5 VDD.n4 GND 0.01fF
C6 VDD.n5 GND 0.02fF
C7 VDD.n6 GND 0.02fF
C8 VDD.n8 GND 0.02fF
C9 VDD.n9 GND 0.02fF
C10 VDD.n11 GND 0.02fF
C11 VDD.n14 GND 0.38fF
C12 VDD.n16 GND 0.03fF
C13 VDD.n17 GND 0.02fF
C14 VDD.n18 GND 0.02fF
C15 VDD.n19 GND 0.02fF
C16 VDD.n20 GND 0.03fF
C17 VDD.n21 GND 0.23fF
C18 VDD.n22 GND 0.02fF
C19 VDD.n23 GND 0.03fF
C20 VDD.n24 GND 0.05fF
C21 VDD.n25 GND 0.12fF
C22 VDD.n26 GND 0.17fF
C23 VDD.n27 GND 0.01fF
C24 VDD.n28 GND 0.01fF
C25 VDD.n29 GND 0.06fF
C26 VDD.n30 GND 0.02fF
C27 VDD.n31 GND 0.02fF
C28 VDD.n32 GND 0.02fF
C29 VDD.n33 GND 0.02fF
C30 VDD.n34 GND 0.02fF
C31 VDD.n35 GND 0.02fF
C32 VDD.n37 GND 0.02fF
C33 VDD.n38 GND 0.02fF
C34 VDD.n39 GND 0.02fF
C35 VDD.n40 GND 0.02fF
C36 VDD.n42 GND 0.03fF
C37 VDD.n43 GND 0.02fF
C38 VDD.n44 GND 0.10fF
C39 VDD.n46 GND 0.38fF
C40 VDD.n48 GND 0.03fF
C41 VDD.n49 GND 0.03fF
C42 VDD.n50 GND 0.23fF
C43 VDD.n51 GND 0.02fF
C44 VDD.n52 GND 0.03fF
C45 VDD.n53 GND 0.02fF
C46 VDD.n54 GND 0.12fF
C47 VDD.n55 GND 0.17fF
C48 VDD.n56 GND 0.01fF
C49 VDD.n57 GND 0.05fF
C50 VDD.n58 GND 0.01fF
C51 VDD.n59 GND 0.02fF
C52 VDD.n60 GND 0.14fF
C53 VDD.n61 GND 0.01fF
C54 VDD.n62 GND 0.02fF
C55 VDD.n63 GND 0.02fF
C56 YN.n0 GND 0.53fF
C57 YN.n1 GND 0.23fF
C58 a_121_411.n0 GND 0.14fF
C59 a_121_411.n1 GND 0.32fF
C60 a_121_411.n2 GND 0.39fF
.ends
