* SPICE3 file created from TMRDFFRNQNX1.ext - technology: sky130A

.subckt TMRDFFRNQNX1 QN D CLK RN VDD VSS
X0 VDD RN a_10507_187 VDD sky130_fd_pr__pfet_01v8 ad=0.003888 pd=3.1488 as=0 ps=0 w=2 l=0.15 M=2
X1 a_14189_1050 a_10637_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X2 a_10959_989 a_10637_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X3 a_599_989 D VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X4 VSS a_10637_1050 a_11413_103 VSS sky130_fd_pr__nfet_01v8 ad=0.0037611 pd=3.297 as=0 ps=0 w=3 l=0.15
X5 a_16421_1051 a_14511_989 QN VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.00116 ps=9.16 w=2 l=0.15 M=2
X6 a_5327_187 RN a_8142_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X7 a_5327_187 CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X8 VDD a_599_989 a_2141_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X9 a_9331_989 a_9009_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X10 a_4151_989 a_147_187 a_4626_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X11 a_1334_210 D a_1053_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X12 VDD CLK a_277_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X13 VDD a_5457_1050 a_5779_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X14 VDD a_5457_1050 a_9009_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X15 VSS a_10959_989 a_12396_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X16 VDD a_277_1050 a_3829_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X17 VDD RN a_5779_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X18 VDD a_9331_989 a_9009_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X19 a_2141_1050 a_147_187 a_2036_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X20 VDD CLK a_10507_187 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X21 VDD CLK a_10637_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X22 a_9331_989 a_5327_187 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X23 VSS a_10507_187 a_10451_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X24 a_14189_1050 RN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X25 a_10959_989 D VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X26 a_599_989 RN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X27 a_3829_1050 a_4151_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X28 VDD a_14511_989 a_15757_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X29 a_10637_1050 a_10507_187 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X30 a_147_187 CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X31 QN a_14511_989 a_15652_101 VSS sky130_fd_pr__nfet_01v8 ad=0.005373 pd=4.72 as=0 ps=0 w=3 l=0.15
X32 a_5779_989 RN a_6514_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X33 a_4151_989 a_3829_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X34 a_11694_210 D a_11413_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X35 a_15757_1051 a_9331_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X36 a_14511_989 a_10507_187 a_14986_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X37 VDD a_14189_1050 a_14511_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X38 VDD a_10959_989 a_12501_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X39 VDD a_147_187 a_2141_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X40 VDD a_599_989 a_277_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X41 VDD D a_5779_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X42 VDD RN a_9009_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X43 VDD a_2141_1050 a_147_187 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X44 VDD a_5327_187 a_5457_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X45 VDD a_7321_1050 a_5327_187 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X46 a_9104_210 RN a_8823_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X47 VSS a_9331_989 a_16318_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X48 a_14189_1050 a_14511_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X49 a_10959_989 RN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X50 a_147_187 RN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X51 a_4151_989 a_147_187 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X52 a_7321_1050 a_5327_187 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X53 a_277_1050 a_599_989 a_372_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X54 QN a_4151_989 a_16421_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X55 a_10732_210 CLK a_10451_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X56 VSS a_5457_1050 a_8823_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X57 VDD a_10959_989 a_10637_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X58 VSS a_5457_1050 a_6233_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X59 a_5457_1050 a_5779_989 a_5552_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X60 VDD a_10507_187 a_14511_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X61 VDD a_10507_187 a_12501_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X62 QN a_14511_989 a_16984_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X63 a_147_187 RN a_2962_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X64 a_8142_210 CLK a_7861_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X65 a_277_1050 a_147_187 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X66 a_16421_1051 a_4151_989 a_15757_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X67 VSS a_9009_1050 a_9806_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X68 a_10507_187 a_12501_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X69 VSS a_5779_989 a_7216_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X70 a_7321_1050 a_5779_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X71 VSS a_147_187 a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X72 VDD a_277_1050 a_599_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X73 VSS a_7321_1050 a_7861_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X74 VSS a_5327_187 a_5271_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X75 a_3829_1050 a_4151_989 a_3924_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X76 a_10507_187 RN a_13322_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X77 a_12501_1050 a_10507_187 a_12396_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X78 a_9331_989 a_5327_187 a_9806_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X79 VDD a_5779_989 a_5457_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X80 VDD RN a_5327_187 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X81 a_16421_1051 a_9331_989 a_15757_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X82 a_6514_210 D a_6233_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X83 VDD RN a_3829_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X84 a_14189_1050 a_14511_989 a_14284_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X85 VSS a_12501_1050 a_13041_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X86 a_372_210 CLK a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X87 VSS a_277_1050 a_3643_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X88 VDD CLK a_5457_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X89 a_5552_210 CLK a_5271_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X90 QN a_4151_989 a_16318_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X91 VSS a_3829_1050 a_4626_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X92 VSS a_599_989 a_2036_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X93 VSS a_10637_1050 a_14003_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X94 VSS a_2141_1050 a_2681_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X95 a_599_989 RN a_1334_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X96 a_10637_1050 a_10959_989 a_10732_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X97 a_13322_210 CLK a_13041_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X98 a_3924_210 RN a_3643_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X99 a_7321_1050 a_5327_187 a_7216_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X100 VSS a_9331_989 a_15652_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X101 VSS a_14189_1050 a_14986_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X102 a_10959_989 RN a_11694_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X103 a_9009_1050 a_9331_989 a_9104_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X104 VSS a_277_1050 a_1053_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X105 a_14284_210 RN a_14003_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X106 a_2962_210 CLK a_2681_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X107 VSS a_4151_989 a_16984_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 VDD a_5327_187 7.74f
C1 a_4151_989 a_9331_989 7.56f
C2 a_10507_187 VDD 7.74f
C3 VDD a_5779_989 3.11f
C4 a_10959_989 VDD 3.11f
C5 a_15757_1051 VDD 3.14f
C6 a_9331_989 a_14511_989 2.55f
C7 VDD a_3829_1050 2.84f
C8 a_4151_989 VDD 2.85f
C9 VDD a_14511_989 4.10f
C10 a_599_989 a_277_1050 2.02f
C11 VDD a_2141_1050 2.17f
C12 VDD a_14189_1050 2.84f
C13 a_277_1050 a_147_187 3.69f
C14 a_10507_187 a_10637_1050 3.69f
C15 CLK a_147_187 5.64f
C16 a_4151_989 D 3.19f
C17 a_10959_989 a_10637_1050 2.02f
C18 RN a_9331_989 2.34f
C19 VDD a_10637_1050 3.23f
C20 a_5327_187 CLK 5.96f
C21 RN VDD 2.66f
C22 VDD a_277_1050 3.23f
C23 a_10507_187 CLK 3.76f
C24 a_5327_187 a_5457_1050 3.69f
C25 VDD CLK 8.54f
C26 VDD a_7321_1050 2.17f
C27 a_5457_1050 a_5779_989 2.02f
C28 a_9009_1050 VDD 2.84f
C29 VDD a_599_989 3.11f
C30 a_4151_989 RN 12.01f
C31 VDD a_147_187 7.74f
C32 VDD a_5457_1050 3.23f
C33 a_12501_1050 VDD 2.17f
C34 VDD a_9331_989 3.26f
C35 D RN 12.60f
C36 RN VSS 7.34f
C37 VDD VSS 28.66f
C38 a_9331_989 VSS 3.02f **FLOATING
C39 a_4151_989 VSS 5.62f **FLOATING
.ends
