* SPICE3 file created from DFFRNQX1.ext - technology: sky130A

.subckt DFFRNQX1 Q D CLK RN VDD VSS
M1000 VDD.t14 RN.t0 a_147_187.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VDD.t7 a_147_187.t8 Q.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t4 a_147_187.t9 a_277_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VSS a_147_187.t10 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1004 a_599_989.t6 D.t0 VDD.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD.t24 CLK.t0 a_277_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VDD.t2 a_599_989.t8 a_2141_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t3 a_277_1050.t7 a_3829_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_599_989.t5 RN.t2 VDD.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_147_187.t6 CLK.t1 VDD.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_3829_1050.t4 Q.t5 VDD.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VSS a_277_1050.t8 a_3643_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1012 Q.t4 a_3829_1050.t7 VDD.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VDD.t6 a_147_187.t11 a_2141_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t1 a_599_989.t9 a_277_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD.t21 a_2141_1050.t5 a_147_187.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VSS a_3829_1050.t8 a_4626_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1017 VSS a_599_989.t10 a_2036_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1018 VSS a_2141_1050.t6 a_2681_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_147_187.t4 RN.t3 VDD.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q.t1 a_147_187.t12 VDD.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_277_1050.t1 a_147_187.t13 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t26 a_277_1050.t9 a_599_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VSS a_277_1050.t11 a_1053_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 VDD.t15 RN.t5 a_599_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 VDD.t28 Q.t7 a_3829_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_277_1050.t5 CLK.t3 VDD.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_2141_1050.t4 a_599_989.t11 VDD.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_3829_1050.t0 a_277_1050.t10 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VDD.t0 D.t1 a_599_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VDD.t12 RN.t7 a_3829_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_599_989.t1 a_277_1050.t12 VDD.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 Q a_147_187.t15 a_4626_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1033 a_277_1050.t6 a_599_989.t12 VDD.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2141_1050.t2 a_147_187.t14 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_147_187.t3 a_2141_1050.t7 VDD.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_3829_1050.t5 RN.t8 VDD.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VDD.t10 CLK.t5 a_147_187.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VDD.t17 a_3829_1050.t9 Q.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 CLK VDD 0.38fF
C1 D VDD 0.05fF
C2 RN VDD 0.17fF
C3 Q VDD 1.39fF
C4 CLK D 0.07fF
C5 RN CLK 0.28fF
C6 RN D 0.18fF
C7 RN Q 0.18fF
R0 a_147_187.n10 a_147_187.t9 512.525
R1 a_147_187.n8 a_147_187.t11 472.359
R2 a_147_187.n6 a_147_187.t8 472.359
R3 a_147_187.n8 a_147_187.t14 384.527
R4 a_147_187.n6 a_147_187.t12 384.527
R5 a_147_187.n10 a_147_187.t13 371.139
R6 a_147_187.n11 a_147_187.t10 340.774
R7 a_147_187.n9 a_147_187.t7 294.278
R8 a_147_187.n7 a_147_187.t15 294.278
R9 a_147_187.n16 a_147_187.n14 266.21
R10 a_147_187.n14 a_147_187.n5 117.693
R11 a_147_187.n11 a_147_187.n10 109.607
R12 a_147_187.n12 a_147_187.n11 83.572
R13 a_147_187.n13 a_147_187.n7 81.396
R14 a_147_187.n4 a_147_187.n3 79.232
R15 a_147_187.n12 a_147_187.n9 76
R16 a_147_187.n14 a_147_187.n13 76
R17 a_147_187.n5 a_147_187.n4 63.152
R18 a_147_187.n9 a_147_187.n8 56.954
R19 a_147_187.n7 a_147_187.n6 56.954
R20 a_147_187.n17 a_147_187.n0 55.263
R21 a_147_187.n16 a_147_187.n15 30
R22 a_147_187.n17 a_147_187.n16 23.684
R23 a_147_187.n5 a_147_187.n1 16.08
R24 a_147_187.n4 a_147_187.n2 16.08
R25 a_147_187.n1 a_147_187.t5 14.282
R26 a_147_187.n1 a_147_187.t4 14.282
R27 a_147_187.n2 a_147_187.t0 14.282
R28 a_147_187.n2 a_147_187.t6 14.282
R29 a_147_187.n3 a_147_187.t1 14.282
R30 a_147_187.n3 a_147_187.t3 14.282
R31 a_147_187.n13 a_147_187.n12 4.035
R32 a_2036_101.n5 a_2036_101.n4 24.877
R33 a_2036_101.t0 a_2036_101.n5 12.677
R34 a_2036_101.t0 a_2036_101.n3 11.595
R35 a_2036_101.t0 a_2036_101.n6 8.137
R36 a_2036_101.n2 a_2036_101.n0 4.031
R37 a_2036_101.n2 a_2036_101.n1 3.644
R38 a_2036_101.t0 a_2036_101.n2 1.093
R39 a_2141_1050.n3 a_2141_1050.t5 512.525
R40 a_2141_1050.n3 a_2141_1050.t7 371.139
R41 a_2141_1050.n4 a_2141_1050.t6 287.668
R42 a_2141_1050.n7 a_2141_1050.n5 217.114
R43 a_2141_1050.n4 a_2141_1050.n3 162.713
R44 a_2141_1050.n5 a_2141_1050.n4 153.315
R45 a_2141_1050.n5 a_2141_1050.n2 152.499
R46 a_2141_1050.n2 a_2141_1050.n1 76.002
R47 a_2141_1050.n7 a_2141_1050.n6 15.218
R48 a_2141_1050.n0 a_2141_1050.t3 14.282
R49 a_2141_1050.n0 a_2141_1050.t2 14.282
R50 a_2141_1050.n1 a_2141_1050.t0 14.282
R51 a_2141_1050.n1 a_2141_1050.t4 14.282
R52 a_2141_1050.n2 a_2141_1050.n0 12.85
R53 a_2141_1050.n8 a_2141_1050.n7 12.014
R54 RN.n0 RN.t7 479.223
R55 RN.n5 RN.t2 454.685
R56 RN.n2 RN.t3 454.685
R57 RN.n5 RN.t5 428.979
R58 RN.n2 RN.t0 428.979
R59 RN.n0 RN.t8 375.52
R60 RN.n6 RN.n5 178.106
R61 RN.n3 RN.n2 178.106
R62 RN.n1 RN.n0 175.429
R63 RN.n1 RN.t6 162.048
R64 RN.n6 RN.t4 158.3
R65 RN.n3 RN.t1 158.3
R66 RN.n4 RN.n1 78.675
R67 RN.n4 RN.n3 76
R68 RN.n7 RN.n6 76
R69 RN.n7 RN.n4 5.94
R70 RN.n7 RN 0.046
R71 VDD.n306 VDD.n304 144.705
R72 VDD.n245 VDD.n243 144.705
R73 VDD.n164 VDD.n162 144.705
R74 VDD.n83 VDD.n81 144.705
R75 VDD.n388 VDD.n386 144.705
R76 VDD.n44 VDD.n43 76
R77 VDD.n49 VDD.n48 76
R78 VDD.n54 VDD.n53 76
R79 VDD.n58 VDD.n57 76
R80 VDD.n85 VDD.n84 76
R81 VDD.n89 VDD.n88 76
R82 VDD.n93 VDD.n92 76
R83 VDD.n98 VDD.n97 76
R84 VDD.n105 VDD.n104 76
R85 VDD.n110 VDD.n109 76
R86 VDD.n115 VDD.n114 76
R87 VDD.n122 VDD.n121 76
R88 VDD.n127 VDD.n126 76
R89 VDD.n132 VDD.n131 76
R90 VDD.n136 VDD.n135 76
R91 VDD.n140 VDD.n139 76
R92 VDD.n166 VDD.n165 76
R93 VDD.n170 VDD.n169 76
R94 VDD.n174 VDD.n173 76
R95 VDD.n179 VDD.n178 76
R96 VDD.n186 VDD.n185 76
R97 VDD.n191 VDD.n190 76
R98 VDD.n196 VDD.n195 76
R99 VDD.n203 VDD.n202 76
R100 VDD.n208 VDD.n207 76
R101 VDD.n213 VDD.n212 76
R102 VDD.n217 VDD.n216 76
R103 VDD.n221 VDD.n220 76
R104 VDD.n247 VDD.n246 76
R105 VDD.n252 VDD.n251 76
R106 VDD.n257 VDD.n256 76
R107 VDD.n263 VDD.n262 76
R108 VDD.n268 VDD.n267 76
R109 VDD.n273 VDD.n272 76
R110 VDD.n278 VDD.n277 76
R111 VDD.n282 VDD.n281 76
R112 VDD.n308 VDD.n307 76
R113 VDD.n312 VDD.n311 76
R114 VDD.n316 VDD.n315 76
R115 VDD.n321 VDD.n320 76
R116 VDD.n328 VDD.n327 76
R117 VDD.n333 VDD.n332 76
R118 VDD.n338 VDD.n337 76
R119 VDD.n345 VDD.n344 76
R120 VDD.n350 VDD.n349 76
R121 VDD.n355 VDD.n354 76
R122 VDD.n359 VDD.n358 76
R123 VDD.n363 VDD.n362 76
R124 VDD.n390 VDD.n389 76
R125 VDD.n394 VDD.n393 76
R126 VDD.n398 VDD.n397 76
R127 VDD.n403 VDD.n402 76
R128 VDD.n410 VDD.n409 76
R129 VDD.n415 VDD.n414 76
R130 VDD.n420 VDD.n419 76
R131 VDD.n427 VDD.n426 76
R132 VDD.n432 VDD.n431 76
R133 VDD.n437 VDD.n436 76
R134 VDD.n441 VDD.n440 76
R135 VDD.n464 VDD.n463 76
R136 VDD.n95 VDD.n94 64.064
R137 VDD.n176 VDD.n175 64.064
R138 VDD.n318 VDD.n317 64.064
R139 VDD.n400 VDD.n399 64.064
R140 VDD.n124 VDD.n123 59.488
R141 VDD.n205 VDD.n204 59.488
R142 VDD.n347 VDD.n346 59.488
R143 VDD.n429 VDD.n428 59.488
R144 VDD.n433 VDD.t8 55.106
R145 VDD.n351 VDD.t22 55.106
R146 VDD.n274 VDD.t27 55.106
R147 VDD.n209 VDD.t20 55.106
R148 VDD.n128 VDD.t18 55.106
R149 VDD.n50 VDD.t23 55.106
R150 VDD.n397 VDD.t1 55.106
R151 VDD.n315 VDD.t15 55.106
R152 VDD.n173 VDD.t14 55.106
R153 VDD.n92 VDD.t28 55.106
R154 VDD.n248 VDD.t6 55.106
R155 VDD.n33 VDD.t7 55.106
R156 VDD.n422 VDD.n421 40.824
R157 VDD.n408 VDD.n407 40.824
R158 VDD.n340 VDD.n339 40.824
R159 VDD.n326 VDD.n325 40.824
R160 VDD.n259 VDD.n258 40.824
R161 VDD.n198 VDD.n197 40.824
R162 VDD.n184 VDD.n183 40.824
R163 VDD.n117 VDD.n116 40.824
R164 VDD.n103 VDD.n102 40.824
R165 VDD.n28 VDD.n27 40.824
R166 VDD.n287 VDD.n286 36.774
R167 VDD.n226 VDD.n225 36.774
R168 VDD.n145 VDD.n144 36.774
R169 VDD.n63 VDD.n62 36.774
R170 VDD.n379 VDD.n378 36.774
R171 VDD.n25 VDD.n24 36.608
R172 VDD.n254 VDD.n253 36.608
R173 VDD.n38 VDD.n37 34.942
R174 VDD.n46 VDD.n45 32.032
R175 VDD.n270 VDD.n269 32.032
R176 VDD.n100 VDD.n99 27.456
R177 VDD.n181 VDD.n180 27.456
R178 VDD.n323 VDD.n322 27.456
R179 VDD.n405 VDD.n404 27.456
R180 VDD.n119 VDD.n118 22.88
R181 VDD.n200 VDD.n199 22.88
R182 VDD.n342 VDD.n341 22.88
R183 VDD.n424 VDD.n423 22.88
R184 VDD.n463 VDD.n460 21.841
R185 VDD.n23 VDD.n20 21.841
R186 VDD.n421 VDD.t29 14.282
R187 VDD.n421 VDD.t4 14.282
R188 VDD.n407 VDD.t30 14.282
R189 VDD.n407 VDD.t24 14.282
R190 VDD.n339 VDD.t19 14.282
R191 VDD.n339 VDD.t26 14.282
R192 VDD.n325 VDD.t16 14.282
R193 VDD.n325 VDD.t0 14.282
R194 VDD.n258 VDD.t5 14.282
R195 VDD.n258 VDD.t2 14.282
R196 VDD.n197 VDD.t31 14.282
R197 VDD.n197 VDD.t21 14.282
R198 VDD.n183 VDD.t13 14.282
R199 VDD.n183 VDD.t10 14.282
R200 VDD.n116 VDD.t11 14.282
R201 VDD.n116 VDD.t3 14.282
R202 VDD.n102 VDD.t25 14.282
R203 VDD.n102 VDD.t12 14.282
R204 VDD.n27 VDD.t9 14.282
R205 VDD.n27 VDD.t17 14.282
R206 VDD.n460 VDD.n443 14.167
R207 VDD.n443 VDD.n442 14.167
R208 VDD.n302 VDD.n284 14.167
R209 VDD.n284 VDD.n283 14.167
R210 VDD.n241 VDD.n223 14.167
R211 VDD.n223 VDD.n222 14.167
R212 VDD.n160 VDD.n142 14.167
R213 VDD.n142 VDD.n141 14.167
R214 VDD.n79 VDD.n60 14.167
R215 VDD.n60 VDD.n59 14.167
R216 VDD.n384 VDD.n365 14.167
R217 VDD.n365 VDD.n364 14.167
R218 VDD.n20 VDD.n19 14.167
R219 VDD.n19 VDD.n17 14.167
R220 VDD.n32 VDD.n31 14.167
R221 VDD.n84 VDD.n80 14.167
R222 VDD.n165 VDD.n161 14.167
R223 VDD.n246 VDD.n242 14.167
R224 VDD.n307 VDD.n303 14.167
R225 VDD.n389 VDD.n385 14.167
R226 VDD.n112 VDD.n111 13.728
R227 VDD.n193 VDD.n192 13.728
R228 VDD.n335 VDD.n334 13.728
R229 VDD.n417 VDD.n416 13.728
R230 VDD.n23 VDD.n22 13.653
R231 VDD.n22 VDD.n21 13.653
R232 VDD.n36 VDD.n35 13.653
R233 VDD.n35 VDD.n34 13.653
R234 VDD.n32 VDD.n26 13.653
R235 VDD.n26 VDD.n25 13.653
R236 VDD.n31 VDD.n30 13.653
R237 VDD.n30 VDD.n29 13.653
R238 VDD.n43 VDD.n42 13.653
R239 VDD.n42 VDD.n41 13.653
R240 VDD.n48 VDD.n47 13.653
R241 VDD.n47 VDD.n46 13.653
R242 VDD.n53 VDD.n52 13.653
R243 VDD.n52 VDD.n51 13.653
R244 VDD.n57 VDD.n56 13.653
R245 VDD.n56 VDD.n55 13.653
R246 VDD.n84 VDD.n83 13.653
R247 VDD.n83 VDD.n82 13.653
R248 VDD.n88 VDD.n87 13.653
R249 VDD.n87 VDD.n86 13.653
R250 VDD.n92 VDD.n91 13.653
R251 VDD.n91 VDD.n90 13.653
R252 VDD.n97 VDD.n96 13.653
R253 VDD.n96 VDD.n95 13.653
R254 VDD.n104 VDD.n101 13.653
R255 VDD.n101 VDD.n100 13.653
R256 VDD.n109 VDD.n108 13.653
R257 VDD.n108 VDD.n107 13.653
R258 VDD.n114 VDD.n113 13.653
R259 VDD.n113 VDD.n112 13.653
R260 VDD.n121 VDD.n120 13.653
R261 VDD.n120 VDD.n119 13.653
R262 VDD.n126 VDD.n125 13.653
R263 VDD.n125 VDD.n124 13.653
R264 VDD.n131 VDD.n130 13.653
R265 VDD.n130 VDD.n129 13.653
R266 VDD.n135 VDD.n134 13.653
R267 VDD.n134 VDD.n133 13.653
R268 VDD.n139 VDD.n138 13.653
R269 VDD.n138 VDD.n137 13.653
R270 VDD.n165 VDD.n164 13.653
R271 VDD.n164 VDD.n163 13.653
R272 VDD.n169 VDD.n168 13.653
R273 VDD.n168 VDD.n167 13.653
R274 VDD.n173 VDD.n172 13.653
R275 VDD.n172 VDD.n171 13.653
R276 VDD.n178 VDD.n177 13.653
R277 VDD.n177 VDD.n176 13.653
R278 VDD.n185 VDD.n182 13.653
R279 VDD.n182 VDD.n181 13.653
R280 VDD.n190 VDD.n189 13.653
R281 VDD.n189 VDD.n188 13.653
R282 VDD.n195 VDD.n194 13.653
R283 VDD.n194 VDD.n193 13.653
R284 VDD.n202 VDD.n201 13.653
R285 VDD.n201 VDD.n200 13.653
R286 VDD.n207 VDD.n206 13.653
R287 VDD.n206 VDD.n205 13.653
R288 VDD.n212 VDD.n211 13.653
R289 VDD.n211 VDD.n210 13.653
R290 VDD.n216 VDD.n215 13.653
R291 VDD.n215 VDD.n214 13.653
R292 VDD.n220 VDD.n219 13.653
R293 VDD.n219 VDD.n218 13.653
R294 VDD.n246 VDD.n245 13.653
R295 VDD.n245 VDD.n244 13.653
R296 VDD.n251 VDD.n250 13.653
R297 VDD.n250 VDD.n249 13.653
R298 VDD.n256 VDD.n255 13.653
R299 VDD.n255 VDD.n254 13.653
R300 VDD.n262 VDD.n261 13.653
R301 VDD.n261 VDD.n260 13.653
R302 VDD.n267 VDD.n266 13.653
R303 VDD.n266 VDD.n265 13.653
R304 VDD.n272 VDD.n271 13.653
R305 VDD.n271 VDD.n270 13.653
R306 VDD.n277 VDD.n276 13.653
R307 VDD.n276 VDD.n275 13.653
R308 VDD.n281 VDD.n280 13.653
R309 VDD.n280 VDD.n279 13.653
R310 VDD.n307 VDD.n306 13.653
R311 VDD.n306 VDD.n305 13.653
R312 VDD.n311 VDD.n310 13.653
R313 VDD.n310 VDD.n309 13.653
R314 VDD.n315 VDD.n314 13.653
R315 VDD.n314 VDD.n313 13.653
R316 VDD.n320 VDD.n319 13.653
R317 VDD.n319 VDD.n318 13.653
R318 VDD.n327 VDD.n324 13.653
R319 VDD.n324 VDD.n323 13.653
R320 VDD.n332 VDD.n331 13.653
R321 VDD.n331 VDD.n330 13.653
R322 VDD.n337 VDD.n336 13.653
R323 VDD.n336 VDD.n335 13.653
R324 VDD.n344 VDD.n343 13.653
R325 VDD.n343 VDD.n342 13.653
R326 VDD.n349 VDD.n348 13.653
R327 VDD.n348 VDD.n347 13.653
R328 VDD.n354 VDD.n353 13.653
R329 VDD.n353 VDD.n352 13.653
R330 VDD.n358 VDD.n357 13.653
R331 VDD.n357 VDD.n356 13.653
R332 VDD.n362 VDD.n361 13.653
R333 VDD.n361 VDD.n360 13.653
R334 VDD.n389 VDD.n388 13.653
R335 VDD.n388 VDD.n387 13.653
R336 VDD.n393 VDD.n392 13.653
R337 VDD.n392 VDD.n391 13.653
R338 VDD.n397 VDD.n396 13.653
R339 VDD.n396 VDD.n395 13.653
R340 VDD.n402 VDD.n401 13.653
R341 VDD.n401 VDD.n400 13.653
R342 VDD.n409 VDD.n406 13.653
R343 VDD.n406 VDD.n405 13.653
R344 VDD.n414 VDD.n413 13.653
R345 VDD.n413 VDD.n412 13.653
R346 VDD.n419 VDD.n418 13.653
R347 VDD.n418 VDD.n417 13.653
R348 VDD.n426 VDD.n425 13.653
R349 VDD.n425 VDD.n424 13.653
R350 VDD.n431 VDD.n430 13.653
R351 VDD.n430 VDD.n429 13.653
R352 VDD.n436 VDD.n435 13.653
R353 VDD.n435 VDD.n434 13.653
R354 VDD.n440 VDD.n439 13.653
R355 VDD.n439 VDD.n438 13.653
R356 VDD.n463 VDD.n462 13.653
R357 VDD.n462 VDD.n461 13.653
R358 VDD.n4 VDD.n2 12.915
R359 VDD.n4 VDD.n3 12.66
R360 VDD.n10 VDD.n9 12.343
R361 VDD.n12 VDD.n11 12.343
R362 VDD.n10 VDD.n7 12.343
R363 VDD.n33 VDD.n32 11.806
R364 VDD.n107 VDD.n106 9.152
R365 VDD.n188 VDD.n187 9.152
R366 VDD.n330 VDD.n329 9.152
R367 VDD.n412 VDD.n411 9.152
R368 VDD.n31 VDD.n28 8.658
R369 VDD.n262 VDD.n259 8.658
R370 VDD.n303 VDD.n302 7.674
R371 VDD.n242 VDD.n241 7.674
R372 VDD.n161 VDD.n160 7.674
R373 VDD.n80 VDD.n79 7.674
R374 VDD.n385 VDD.n384 7.674
R375 VDD.n74 VDD.n73 7.5
R376 VDD.n68 VDD.n67 7.5
R377 VDD.n70 VDD.n69 7.5
R378 VDD.n65 VDD.n64 7.5
R379 VDD.n79 VDD.n78 7.5
R380 VDD.n155 VDD.n154 7.5
R381 VDD.n149 VDD.n148 7.5
R382 VDD.n151 VDD.n150 7.5
R383 VDD.n157 VDD.n147 7.5
R384 VDD.n157 VDD.n145 7.5
R385 VDD.n160 VDD.n159 7.5
R386 VDD.n236 VDD.n235 7.5
R387 VDD.n230 VDD.n229 7.5
R388 VDD.n232 VDD.n231 7.5
R389 VDD.n238 VDD.n228 7.5
R390 VDD.n238 VDD.n226 7.5
R391 VDD.n241 VDD.n240 7.5
R392 VDD.n297 VDD.n296 7.5
R393 VDD.n291 VDD.n290 7.5
R394 VDD.n293 VDD.n292 7.5
R395 VDD.n299 VDD.n289 7.5
R396 VDD.n299 VDD.n287 7.5
R397 VDD.n302 VDD.n301 7.5
R398 VDD.n369 VDD.n368 7.5
R399 VDD.n372 VDD.n371 7.5
R400 VDD.n374 VDD.n373 7.5
R401 VDD.n377 VDD.n376 7.5
R402 VDD.n384 VDD.n383 7.5
R403 VDD.n455 VDD.n454 7.5
R404 VDD.n449 VDD.n448 7.5
R405 VDD.n451 VDD.n450 7.5
R406 VDD.n457 VDD.n447 7.5
R407 VDD.n457 VDD.n445 7.5
R408 VDD.n460 VDD.n459 7.5
R409 VDD.n20 VDD.n16 7.5
R410 VDD.n2 VDD.n1 7.5
R411 VDD.n9 VDD.n8 7.5
R412 VDD.n7 VDD.n6 7.5
R413 VDD.n19 VDD.n18 7.5
R414 VDD.n14 VDD.n0 7.5
R415 VDD.n66 VDD.n63 6.772
R416 VDD.n77 VDD.n61 6.772
R417 VDD.n75 VDD.n72 6.772
R418 VDD.n71 VDD.n68 6.772
R419 VDD.n158 VDD.n143 6.772
R420 VDD.n156 VDD.n153 6.772
R421 VDD.n152 VDD.n149 6.772
R422 VDD.n239 VDD.n224 6.772
R423 VDD.n237 VDD.n234 6.772
R424 VDD.n233 VDD.n230 6.772
R425 VDD.n300 VDD.n285 6.772
R426 VDD.n298 VDD.n295 6.772
R427 VDD.n294 VDD.n291 6.772
R428 VDD.n458 VDD.n444 6.772
R429 VDD.n456 VDD.n453 6.772
R430 VDD.n452 VDD.n449 6.772
R431 VDD.n66 VDD.n65 6.772
R432 VDD.n71 VDD.n70 6.772
R433 VDD.n75 VDD.n74 6.772
R434 VDD.n78 VDD.n77 6.772
R435 VDD.n152 VDD.n151 6.772
R436 VDD.n156 VDD.n155 6.772
R437 VDD.n159 VDD.n158 6.772
R438 VDD.n233 VDD.n232 6.772
R439 VDD.n237 VDD.n236 6.772
R440 VDD.n240 VDD.n239 6.772
R441 VDD.n294 VDD.n293 6.772
R442 VDD.n298 VDD.n297 6.772
R443 VDD.n301 VDD.n300 6.772
R444 VDD.n452 VDD.n451 6.772
R445 VDD.n456 VDD.n455 6.772
R446 VDD.n459 VDD.n458 6.772
R447 VDD.n383 VDD.n382 6.772
R448 VDD.n370 VDD.n367 6.772
R449 VDD.n375 VDD.n372 6.772
R450 VDD.n380 VDD.n377 6.772
R451 VDD.n380 VDD.n379 6.772
R452 VDD.n375 VDD.n374 6.772
R453 VDD.n370 VDD.n369 6.772
R454 VDD.n382 VDD.n366 6.772
R455 VDD.n121 VDD.n117 6.69
R456 VDD.n202 VDD.n198 6.69
R457 VDD.n344 VDD.n340 6.69
R458 VDD.n426 VDD.n422 6.69
R459 VDD.n37 VDD.n23 6.487
R460 VDD.n37 VDD.n36 6.475
R461 VDD.n16 VDD.n15 6.458
R462 VDD.n104 VDD.n103 6.296
R463 VDD.n185 VDD.n184 6.296
R464 VDD.n327 VDD.n326 6.296
R465 VDD.n409 VDD.n408 6.296
R466 VDD.n147 VDD.n146 6.202
R467 VDD.n228 VDD.n227 6.202
R468 VDD.n289 VDD.n288 6.202
R469 VDD.n447 VDD.n446 6.202
R470 VDD.n41 VDD.n40 4.576
R471 VDD.n265 VDD.n264 4.576
R472 VDD.n53 VDD.n50 2.754
R473 VDD.n277 VDD.n274 2.754
R474 VDD.n36 VDD.n33 2.361
R475 VDD.n251 VDD.n248 2.361
R476 VDD.n14 VDD.n5 1.329
R477 VDD.n14 VDD.n10 1.329
R478 VDD.n14 VDD.n12 1.329
R479 VDD.n14 VDD.n13 1.329
R480 VDD.n15 VDD.n14 0.696
R481 VDD.n14 VDD.n4 0.696
R482 VDD.n131 VDD.n128 0.393
R483 VDD.n212 VDD.n209 0.393
R484 VDD.n354 VDD.n351 0.393
R485 VDD.n436 VDD.n433 0.393
R486 VDD.n76 VDD.n75 0.365
R487 VDD.n76 VDD.n71 0.365
R488 VDD.n76 VDD.n66 0.365
R489 VDD.n77 VDD.n76 0.365
R490 VDD.n157 VDD.n156 0.365
R491 VDD.n157 VDD.n152 0.365
R492 VDD.n158 VDD.n157 0.365
R493 VDD.n238 VDD.n237 0.365
R494 VDD.n238 VDD.n233 0.365
R495 VDD.n239 VDD.n238 0.365
R496 VDD.n299 VDD.n298 0.365
R497 VDD.n299 VDD.n294 0.365
R498 VDD.n300 VDD.n299 0.365
R499 VDD.n457 VDD.n456 0.365
R500 VDD.n457 VDD.n452 0.365
R501 VDD.n458 VDD.n457 0.365
R502 VDD.n381 VDD.n380 0.365
R503 VDD.n381 VDD.n375 0.365
R504 VDD.n381 VDD.n370 0.365
R505 VDD.n382 VDD.n381 0.365
R506 VDD.n85 VDD.n58 0.29
R507 VDD.n166 VDD.n140 0.29
R508 VDD.n247 VDD.n221 0.29
R509 VDD.n308 VDD.n282 0.29
R510 VDD.n390 VDD.n363 0.29
R511 VDD.n115 VDD.n110 0.197
R512 VDD.n196 VDD.n191 0.197
R513 VDD.n338 VDD.n333 0.197
R514 VDD.n420 VDD.n415 0.197
R515 VDD.n44 VDD.n39 0.181
R516 VDD.n268 VDD.n263 0.181
R517 VDD.n39 VDD.n38 0.145
R518 VDD.n49 VDD.n44 0.145
R519 VDD.n54 VDD.n49 0.145
R520 VDD.n58 VDD.n54 0.145
R521 VDD.n89 VDD.n85 0.145
R522 VDD.n93 VDD.n89 0.145
R523 VDD.n98 VDD.n93 0.145
R524 VDD.n105 VDD.n98 0.145
R525 VDD.n110 VDD.n105 0.145
R526 VDD.n122 VDD.n115 0.145
R527 VDD.n127 VDD.n122 0.145
R528 VDD.n132 VDD.n127 0.145
R529 VDD.n136 VDD.n132 0.145
R530 VDD.n140 VDD.n136 0.145
R531 VDD.n170 VDD.n166 0.145
R532 VDD.n174 VDD.n170 0.145
R533 VDD.n179 VDD.n174 0.145
R534 VDD.n186 VDD.n179 0.145
R535 VDD.n191 VDD.n186 0.145
R536 VDD.n203 VDD.n196 0.145
R537 VDD.n208 VDD.n203 0.145
R538 VDD.n213 VDD.n208 0.145
R539 VDD.n217 VDD.n213 0.145
R540 VDD.n221 VDD.n217 0.145
R541 VDD.n252 VDD.n247 0.145
R542 VDD.n257 VDD.n252 0.145
R543 VDD.n263 VDD.n257 0.145
R544 VDD.n273 VDD.n268 0.145
R545 VDD.n278 VDD.n273 0.145
R546 VDD.n282 VDD.n278 0.145
R547 VDD.n312 VDD.n308 0.145
R548 VDD.n316 VDD.n312 0.145
R549 VDD.n321 VDD.n316 0.145
R550 VDD.n328 VDD.n321 0.145
R551 VDD.n333 VDD.n328 0.145
R552 VDD.n345 VDD.n338 0.145
R553 VDD.n350 VDD.n345 0.145
R554 VDD.n355 VDD.n350 0.145
R555 VDD.n359 VDD.n355 0.145
R556 VDD.n363 VDD.n359 0.145
R557 VDD.n394 VDD.n390 0.145
R558 VDD.n398 VDD.n394 0.145
R559 VDD.n403 VDD.n398 0.145
R560 VDD.n410 VDD.n403 0.145
R561 VDD.n415 VDD.n410 0.145
R562 VDD.n427 VDD.n420 0.145
R563 VDD.n432 VDD.n427 0.145
R564 VDD.n437 VDD.n432 0.145
R565 VDD.n441 VDD.n437 0.145
R566 VDD.n464 VDD.n441 0.145
R567 VDD.n464 VDD 0.034
R568 Q.n8 Q.t5 454.685
R569 Q.n8 Q.t7 428.979
R570 Q.n9 Q.t6 264.512
R571 Q.n7 Q.n6 237.145
R572 Q.n7 Q.n2 125.947
R573 Q Q.n9 78.901
R574 Q.n2 Q.n1 76.002
R575 Q.n10 Q.n7 76
R576 Q.n9 Q.n8 71.894
R577 Q.n6 Q.n5 30
R578 Q.n4 Q.n3 24.383
R579 Q.n6 Q.n4 23.684
R580 Q.n0 Q.t2 14.282
R581 Q.n0 Q.t1 14.282
R582 Q.n1 Q.t3 14.282
R583 Q.n1 Q.t4 14.282
R584 Q.n2 Q.n0 12.85
R585 Q.n10 Q 0.046
R586 a_277_1050.n4 a_277_1050.t9 512.525
R587 a_277_1050.n2 a_277_1050.t7 512.525
R588 a_277_1050.n4 a_277_1050.t12 371.139
R589 a_277_1050.n2 a_277_1050.t10 371.139
R590 a_277_1050.n5 a_277_1050.t11 314.221
R591 a_277_1050.n3 a_277_1050.t8 314.221
R592 a_277_1050.n8 a_277_1050.n7 261.396
R593 a_277_1050.n9 a_277_1050.n8 144.246
R594 a_277_1050.n5 a_277_1050.n4 136.16
R595 a_277_1050.n3 a_277_1050.n2 136.16
R596 a_277_1050.n6 a_277_1050.n3 85.476
R597 a_277_1050.n11 a_277_1050.n10 79.231
R598 a_277_1050.n8 a_277_1050.n6 77.315
R599 a_277_1050.n6 a_277_1050.n5 76
R600 a_277_1050.n10 a_277_1050.n9 63.152
R601 a_277_1050.n9 a_277_1050.n1 16.08
R602 a_277_1050.n10 a_277_1050.n0 16.08
R603 a_277_1050.n1 a_277_1050.t0 14.282
R604 a_277_1050.n1 a_277_1050.t6 14.282
R605 a_277_1050.n0 a_277_1050.t4 14.282
R606 a_277_1050.n0 a_277_1050.t5 14.282
R607 a_277_1050.t2 a_277_1050.n11 14.282
R608 a_277_1050.n11 a_277_1050.t1 14.282
R609 a_599_989.n2 a_599_989.t8 480.392
R610 a_599_989.n4 a_599_989.t12 454.685
R611 a_599_989.n4 a_599_989.t9 428.979
R612 a_599_989.n2 a_599_989.t11 403.272
R613 a_599_989.n3 a_599_989.t10 283.48
R614 a_599_989.n5 a_599_989.t7 237.959
R615 a_599_989.n11 a_599_989.n10 213.104
R616 a_599_989.n12 a_599_989.n11 170.799
R617 a_599_989.n5 a_599_989.n4 98.447
R618 a_599_989.n3 a_599_989.n2 98.447
R619 a_599_989.n6 a_599_989.n5 80.035
R620 a_599_989.n14 a_599_989.n13 79.231
R621 a_599_989.n6 a_599_989.n3 77.315
R622 a_599_989.n11 a_599_989.n6 76
R623 a_599_989.n13 a_599_989.n12 63.152
R624 a_599_989.n10 a_599_989.n9 30
R625 a_599_989.n8 a_599_989.n7 24.383
R626 a_599_989.n10 a_599_989.n8 23.684
R627 a_599_989.n12 a_599_989.n1 16.08
R628 a_599_989.n13 a_599_989.n0 16.08
R629 a_599_989.n1 a_599_989.t4 14.282
R630 a_599_989.n1 a_599_989.t5 14.282
R631 a_599_989.n0 a_599_989.t0 14.282
R632 a_599_989.n0 a_599_989.t6 14.282
R633 a_599_989.t2 a_599_989.n14 14.282
R634 a_599_989.n14 a_599_989.t1 14.282
R635 a_372_210.n10 a_372_210.n8 82.852
R636 a_372_210.n11 a_372_210.n0 49.6
R637 a_372_210.n7 a_372_210.n6 32.833
R638 a_372_210.n8 a_372_210.t1 32.416
R639 a_372_210.n10 a_372_210.n9 27.2
R640 a_372_210.n3 a_372_210.n2 23.284
R641 a_372_210.n11 a_372_210.n10 22.4
R642 a_372_210.n7 a_372_210.n4 19.017
R643 a_372_210.n6 a_372_210.n5 13.494
R644 a_372_210.t1 a_372_210.n1 7.04
R645 a_372_210.t1 a_372_210.n3 5.727
R646 a_372_210.n8 a_372_210.n7 1.435
R647 D.n0 D.t1 479.223
R648 D.n0 D.t0 375.52
R649 D.n1 D.t2 215.154
R650 D.n1 D.n0 122.323
R651 D.n2 D.n1 76
R652 D.n2 D 0.046
R653 a_2962_210.n10 a_2962_210.n8 82.852
R654 a_2962_210.n11 a_2962_210.n0 49.6
R655 a_2962_210.n7 a_2962_210.n6 32.833
R656 a_2962_210.n8 a_2962_210.t1 32.416
R657 a_2962_210.n10 a_2962_210.n9 27.2
R658 a_2962_210.n3 a_2962_210.n2 23.284
R659 a_2962_210.n11 a_2962_210.n10 22.4
R660 a_2962_210.n7 a_2962_210.n4 19.017
R661 a_2962_210.n6 a_2962_210.n5 13.494
R662 a_2962_210.t1 a_2962_210.n1 7.04
R663 a_2962_210.t1 a_2962_210.n3 5.727
R664 a_2962_210.n8 a_2962_210.n7 1.435
R665 CLK.n2 CLK.t0 459.505
R666 CLK.n0 CLK.t5 459.505
R667 CLK.n2 CLK.t3 384.527
R668 CLK.n0 CLK.t1 384.527
R669 CLK.n3 CLK.t2 322.152
R670 CLK.n1 CLK.t4 322.151
R671 CLK.n4 CLK.n1 58.818
R672 CLK.n4 CLK.n3 49.342
R673 CLK.n3 CLK.n2 27.599
R674 CLK.n1 CLK.n0 27.599
R675 CLK.n4 CLK 0.046
R676 a_3829_1050.n2 a_3829_1050.t9 480.392
R677 a_3829_1050.n2 a_3829_1050.t7 403.272
R678 a_3829_1050.n3 a_3829_1050.t8 283.48
R679 a_3829_1050.n8 a_3829_1050.n7 213.104
R680 a_3829_1050.n9 a_3829_1050.n8 170.799
R681 a_3829_1050.n8 a_3829_1050.n3 153.315
R682 a_3829_1050.n3 a_3829_1050.n2 98.447
R683 a_3829_1050.n11 a_3829_1050.n10 79.231
R684 a_3829_1050.n10 a_3829_1050.n9 63.152
R685 a_3829_1050.n7 a_3829_1050.n6 30
R686 a_3829_1050.n5 a_3829_1050.n4 24.383
R687 a_3829_1050.n7 a_3829_1050.n5 23.684
R688 a_3829_1050.n9 a_3829_1050.n1 16.08
R689 a_3829_1050.n10 a_3829_1050.n0 16.08
R690 a_3829_1050.n1 a_3829_1050.t3 14.282
R691 a_3829_1050.n1 a_3829_1050.t4 14.282
R692 a_3829_1050.n0 a_3829_1050.t6 14.282
R693 a_3829_1050.n0 a_3829_1050.t5 14.282
R694 a_3829_1050.t1 a_3829_1050.n11 14.282
R695 a_3829_1050.n11 a_3829_1050.t0 14.282
R696 a_91_103.t0 a_91_103.n3 117.777
R697 a_91_103.n6 a_91_103.n5 45.444
R698 a_91_103.t0 a_91_103.n6 21.213
R699 a_91_103.t0 a_91_103.n4 11.595
R700 a_91_103.n2 a_91_103.n1 2.455
R701 a_91_103.n2 a_91_103.n0 1.32
R702 a_91_103.t0 a_91_103.n2 0.246
R703 VSS.n29 VSS.n27 219.745
R704 VSS.n194 VSS.n193 219.745
R705 VSS.n149 VSS.n147 219.745
R706 VSS.n119 VSS.n117 219.745
R707 VSS.n74 VSS.n73 219.745
R708 VSS.n225 VSS.n224 85.559
R709 VSS.n29 VSS.n28 85.529
R710 VSS.n194 VSS.n192 85.529
R711 VSS.n149 VSS.n148 85.529
R712 VSS.n119 VSS.n118 85.529
R713 VSS.n74 VSS.n72 85.529
R714 VSS.n137 VSS.n136 84.842
R715 VSS.n233 VSS.n232 76
R716 VSS.n12 VSS.n11 76
R717 VSS.n20 VSS.n19 76
R718 VSS.n23 VSS.n22 76
R719 VSS.n26 VSS.n25 76
R720 VSS.n33 VSS.n32 76
R721 VSS.n36 VSS.n35 76
R722 VSS.n39 VSS.n38 76
R723 VSS.n42 VSS.n41 76
R724 VSS.n45 VSS.n44 76
R725 VSS.n48 VSS.n47 76
R726 VSS.n51 VSS.n50 76
R727 VSS.n54 VSS.n53 76
R728 VSS.n57 VSS.n56 76
R729 VSS.n65 VSS.n64 76
R730 VSS.n68 VSS.n67 76
R731 VSS.n71 VSS.n70 76
R732 VSS.n78 VSS.n77 76
R733 VSS.n81 VSS.n80 76
R734 VSS.n84 VSS.n83 76
R735 VSS.n87 VSS.n86 76
R736 VSS.n90 VSS.n89 76
R737 VSS.n93 VSS.n92 76
R738 VSS.n96 VSS.n95 76
R739 VSS.n99 VSS.n98 76
R740 VSS.n102 VSS.n101 76
R741 VSS.n110 VSS.n109 76
R742 VSS.n113 VSS.n112 76
R743 VSS.n116 VSS.n115 76
R744 VSS.n123 VSS.n122 76
R745 VSS.n126 VSS.n125 76
R746 VSS.n129 VSS.n128 76
R747 VSS.n132 VSS.n131 76
R748 VSS.n135 VSS.n134 76
R749 VSS.n140 VSS.n139 76
R750 VSS.n143 VSS.n142 76
R751 VSS.n146 VSS.n145 76
R752 VSS.n153 VSS.n152 76
R753 VSS.n156 VSS.n155 76
R754 VSS.n159 VSS.n158 76
R755 VSS.n162 VSS.n161 76
R756 VSS.n165 VSS.n164 76
R757 VSS.n168 VSS.n167 76
R758 VSS.n171 VSS.n170 76
R759 VSS.n174 VSS.n173 76
R760 VSS.n177 VSS.n176 76
R761 VSS.n185 VSS.n184 76
R762 VSS.n188 VSS.n187 76
R763 VSS.n191 VSS.n190 76
R764 VSS.n198 VSS.n197 76
R765 VSS.n201 VSS.n200 76
R766 VSS.n204 VSS.n203 76
R767 VSS.n207 VSS.n206 76
R768 VSS.n210 VSS.n209 76
R769 VSS.n213 VSS.n212 76
R770 VSS.n216 VSS.n215 76
R771 VSS.n219 VSS.n218 76
R772 VSS.n222 VSS.n221 76
R773 VSS.n227 VSS.n226 76
R774 VSS.n230 VSS.n229 76
R775 VSS.n63 VSS.n62 64.552
R776 VSS.n108 VSS.n107 64.552
R777 VSS.n183 VSS.n182 64.552
R778 VSS.n17 VSS.n16 63.835
R779 VSS.n8 VSS.n7 34.942
R780 VSS.n16 VSS.n15 28.421
R781 VSS.n62 VSS.n61 28.421
R782 VSS.n107 VSS.n106 28.421
R783 VSS.n182 VSS.n181 28.421
R784 VSS.n16 VSS.n14 25.263
R785 VSS.n62 VSS.n60 25.263
R786 VSS.n107 VSS.n105 25.263
R787 VSS.n182 VSS.n180 25.263
R788 VSS.n14 VSS.n13 24.383
R789 VSS.n60 VSS.n59 24.383
R790 VSS.n105 VSS.n104 24.383
R791 VSS.n180 VSS.n179 24.383
R792 VSS.n6 VSS.n5 14.167
R793 VSS.n5 VSS.n4 14.167
R794 VSS.n32 VSS.n30 14.167
R795 VSS.n77 VSS.n75 14.167
R796 VSS.n122 VSS.n120 14.167
R797 VSS.n152 VSS.n150 14.167
R798 VSS.n197 VSS.n195 14.167
R799 VSS.n229 VSS.n228 13.653
R800 VSS.n226 VSS.n223 13.653
R801 VSS.n221 VSS.n220 13.653
R802 VSS.n218 VSS.n217 13.653
R803 VSS.n215 VSS.n214 13.653
R804 VSS.n212 VSS.n211 13.653
R805 VSS.n209 VSS.n208 13.653
R806 VSS.n206 VSS.n205 13.653
R807 VSS.n203 VSS.n202 13.653
R808 VSS.n200 VSS.n199 13.653
R809 VSS.n197 VSS.n196 13.653
R810 VSS.n190 VSS.n189 13.653
R811 VSS.n187 VSS.n186 13.653
R812 VSS.n184 VSS.n178 13.653
R813 VSS.n176 VSS.n175 13.653
R814 VSS.n173 VSS.n172 13.653
R815 VSS.n170 VSS.n169 13.653
R816 VSS.n167 VSS.n166 13.653
R817 VSS.n164 VSS.n163 13.653
R818 VSS.n161 VSS.n160 13.653
R819 VSS.n158 VSS.n157 13.653
R820 VSS.n155 VSS.n154 13.653
R821 VSS.n152 VSS.n151 13.653
R822 VSS.n145 VSS.n144 13.653
R823 VSS.n142 VSS.n141 13.653
R824 VSS.n139 VSS.n138 13.653
R825 VSS.n134 VSS.n133 13.653
R826 VSS.n131 VSS.n130 13.653
R827 VSS.n128 VSS.n127 13.653
R828 VSS.n125 VSS.n124 13.653
R829 VSS.n122 VSS.n121 13.653
R830 VSS.n115 VSS.n114 13.653
R831 VSS.n112 VSS.n111 13.653
R832 VSS.n109 VSS.n103 13.653
R833 VSS.n101 VSS.n100 13.653
R834 VSS.n98 VSS.n97 13.653
R835 VSS.n95 VSS.n94 13.653
R836 VSS.n92 VSS.n91 13.653
R837 VSS.n89 VSS.n88 13.653
R838 VSS.n86 VSS.n85 13.653
R839 VSS.n83 VSS.n82 13.653
R840 VSS.n80 VSS.n79 13.653
R841 VSS.n77 VSS.n76 13.653
R842 VSS.n70 VSS.n69 13.653
R843 VSS.n67 VSS.n66 13.653
R844 VSS.n64 VSS.n58 13.653
R845 VSS.n56 VSS.n55 13.653
R846 VSS.n53 VSS.n52 13.653
R847 VSS.n50 VSS.n49 13.653
R848 VSS.n47 VSS.n46 13.653
R849 VSS.n44 VSS.n43 13.653
R850 VSS.n41 VSS.n40 13.653
R851 VSS.n38 VSS.n37 13.653
R852 VSS.n35 VSS.n34 13.653
R853 VSS.n32 VSS.n31 13.653
R854 VSS.n25 VSS.n24 13.653
R855 VSS.n22 VSS.n21 13.653
R856 VSS.n19 VSS.n18 13.653
R857 VSS.n11 VSS.n10 13.653
R858 VSS.n4 VSS.n3 13.653
R859 VSS.n5 VSS.n2 13.653
R860 VSS.n6 VSS.n1 13.653
R861 VSS.n30 VSS.n29 7.312
R862 VSS.n195 VSS.n194 7.312
R863 VSS.n150 VSS.n149 7.312
R864 VSS.n120 VSS.n119 7.312
R865 VSS.n75 VSS.n74 7.312
R866 VSS.n7 VSS.n0 7.083
R867 VSS.n7 VSS.n6 6.474
R868 VSS.n19 VSS.n17 3.935
R869 VSS.n139 VSS.n137 3.935
R870 VSS.n232 VSS.n231 0.596
R871 VSS.n33 VSS.n26 0.29
R872 VSS.n78 VSS.n71 0.29
R873 VSS.n123 VSS.n116 0.29
R874 VSS.n153 VSS.n146 0.29
R875 VSS.n198 VSS.n191 0.29
R876 VSS.n51 VSS.n48 0.197
R877 VSS.n96 VSS.n93 0.197
R878 VSS.n171 VSS.n168 0.197
R879 VSS.n216 VSS.n213 0.197
R880 VSS.n64 VSS.n63 0.196
R881 VSS.n109 VSS.n108 0.196
R882 VSS.n184 VSS.n183 0.196
R883 VSS.n226 VSS.n225 0.196
R884 VSS.n12 VSS.n9 0.181
R885 VSS.n135 VSS.n132 0.181
R886 VSS.n9 VSS.n8 0.145
R887 VSS.n20 VSS.n12 0.145
R888 VSS.n23 VSS.n20 0.145
R889 VSS.n26 VSS.n23 0.145
R890 VSS.n36 VSS.n33 0.145
R891 VSS.n39 VSS.n36 0.145
R892 VSS.n42 VSS.n39 0.145
R893 VSS.n45 VSS.n42 0.145
R894 VSS.n48 VSS.n45 0.145
R895 VSS.n54 VSS.n51 0.145
R896 VSS.n57 VSS.n54 0.145
R897 VSS.n65 VSS.n57 0.145
R898 VSS.n68 VSS.n65 0.145
R899 VSS.n71 VSS.n68 0.145
R900 VSS.n81 VSS.n78 0.145
R901 VSS.n84 VSS.n81 0.145
R902 VSS.n87 VSS.n84 0.145
R903 VSS.n90 VSS.n87 0.145
R904 VSS.n93 VSS.n90 0.145
R905 VSS.n99 VSS.n96 0.145
R906 VSS.n102 VSS.n99 0.145
R907 VSS.n110 VSS.n102 0.145
R908 VSS.n113 VSS.n110 0.145
R909 VSS.n116 VSS.n113 0.145
R910 VSS.n126 VSS.n123 0.145
R911 VSS.n129 VSS.n126 0.145
R912 VSS.n132 VSS.n129 0.145
R913 VSS.n140 VSS.n135 0.145
R914 VSS.n143 VSS.n140 0.145
R915 VSS.n146 VSS.n143 0.145
R916 VSS.n156 VSS.n153 0.145
R917 VSS.n159 VSS.n156 0.145
R918 VSS.n162 VSS.n159 0.145
R919 VSS.n165 VSS.n162 0.145
R920 VSS.n168 VSS.n165 0.145
R921 VSS.n174 VSS.n171 0.145
R922 VSS.n177 VSS.n174 0.145
R923 VSS.n185 VSS.n177 0.145
R924 VSS.n188 VSS.n185 0.145
R925 VSS.n191 VSS.n188 0.145
R926 VSS.n201 VSS.n198 0.145
R927 VSS.n204 VSS.n201 0.145
R928 VSS.n207 VSS.n204 0.145
R929 VSS.n210 VSS.n207 0.145
R930 VSS.n213 VSS.n210 0.145
R931 VSS.n219 VSS.n216 0.145
R932 VSS.n222 VSS.n219 0.145
R933 VSS.n227 VSS.n222 0.145
R934 VSS.n230 VSS.n227 0.145
R935 VSS.n233 VSS.n230 0.145
R936 VSS.n233 VSS 0.034
R937 a_3924_210.n9 a_3924_210.n7 82.852
R938 a_3924_210.n3 a_3924_210.n1 44.628
R939 a_3924_210.t0 a_3924_210.n9 32.417
R940 a_3924_210.n7 a_3924_210.n6 27.2
R941 a_3924_210.n5 a_3924_210.n4 23.498
R942 a_3924_210.n3 a_3924_210.n2 23.284
R943 a_3924_210.n7 a_3924_210.n5 22.4
R944 a_3924_210.t0 a_3924_210.n11 20.241
R945 a_3924_210.n11 a_3924_210.n10 13.494
R946 a_3924_210.t0 a_3924_210.n0 8.137
R947 a_3924_210.t0 a_3924_210.n3 5.727
R948 a_3924_210.n9 a_3924_210.n8 1.435
R949 a_3643_103.n5 a_3643_103.n4 19.724
R950 a_3643_103.t0 a_3643_103.n3 11.595
R951 a_3643_103.t0 a_3643_103.n5 9.207
R952 a_3643_103.n2 a_3643_103.n1 2.455
R953 a_3643_103.n2 a_3643_103.n0 1.32
R954 a_3643_103.t0 a_3643_103.n2 0.246
R955 a_4626_101.t0 a_4626_101.n1 34.62
R956 a_4626_101.t0 a_4626_101.n0 8.137
R957 a_4626_101.t0 a_4626_101.n2 4.69
R958 a_1334_210.n9 a_1334_210.n7 82.852
R959 a_1334_210.n3 a_1334_210.n1 44.628
R960 a_1334_210.t0 a_1334_210.n9 32.417
R961 a_1334_210.n7 a_1334_210.n6 27.2
R962 a_1334_210.n5 a_1334_210.n4 23.498
R963 a_1334_210.n3 a_1334_210.n2 23.284
R964 a_1334_210.n7 a_1334_210.n5 22.4
R965 a_1334_210.t0 a_1334_210.n11 20.241
R966 a_1334_210.n11 a_1334_210.n10 13.494
R967 a_1334_210.t0 a_1334_210.n0 8.137
R968 a_1334_210.t0 a_1334_210.n3 5.727
R969 a_1334_210.n9 a_1334_210.n8 1.435
R970 a_2681_103.n5 a_2681_103.n4 19.724
R971 a_2681_103.t0 a_2681_103.n3 11.595
R972 a_2681_103.t0 a_2681_103.n5 9.207
R973 a_2681_103.n2 a_2681_103.n1 2.455
R974 a_2681_103.n2 a_2681_103.n0 1.32
R975 a_2681_103.t0 a_2681_103.n2 0.246
R976 a_1053_103.n5 a_1053_103.n4 19.724
R977 a_1053_103.t0 a_1053_103.n3 11.595
R978 a_1053_103.t0 a_1053_103.n5 9.207
R979 a_1053_103.n2 a_1053_103.n1 2.455
R980 a_1053_103.n2 a_1053_103.n0 1.32
R981 a_1053_103.t0 a_1053_103.n2 0.246
C8 RN VSS 2.65fF
C9 VDD VSS 19.26fF
C10 a_1053_103.n0 VSS 0.10fF
C11 a_1053_103.n1 VSS 0.04fF
C12 a_1053_103.n2 VSS 0.03fF
C13 a_1053_103.n3 VSS 0.07fF
C14 a_1053_103.n4 VSS 0.08fF
C15 a_1053_103.n5 VSS 0.06fF
C16 a_2681_103.n0 VSS 0.10fF
C17 a_2681_103.n1 VSS 0.04fF
C18 a_2681_103.n2 VSS 0.03fF
C19 a_2681_103.n3 VSS 0.07fF
C20 a_2681_103.n4 VSS 0.08fF
C21 a_2681_103.n5 VSS 0.06fF
C22 a_1334_210.n0 VSS 0.07fF
C23 a_1334_210.n1 VSS 0.09fF
C24 a_1334_210.n2 VSS 0.13fF
C25 a_1334_210.n3 VSS 0.11fF
C26 a_1334_210.n4 VSS 0.02fF
C27 a_1334_210.n5 VSS 0.03fF
C28 a_1334_210.n6 VSS 0.02fF
C29 a_1334_210.n7 VSS 0.05fF
C30 a_1334_210.n8 VSS 0.03fF
C31 a_1334_210.n9 VSS 0.11fF
C32 a_1334_210.n10 VSS 0.06fF
C33 a_1334_210.n11 VSS 0.01fF
C34 a_1334_210.t0 VSS 0.33fF
C35 a_4626_101.n0 VSS 0.05fF
C36 a_4626_101.n1 VSS 0.12fF
C37 a_4626_101.n2 VSS 0.04fF
C38 a_3643_103.n0 VSS 0.10fF
C39 a_3643_103.n1 VSS 0.04fF
C40 a_3643_103.n2 VSS 0.03fF
C41 a_3643_103.n3 VSS 0.07fF
C42 a_3643_103.n4 VSS 0.08fF
C43 a_3643_103.n5 VSS 0.06fF
C44 a_3924_210.n0 VSS 0.07fF
C45 a_3924_210.n1 VSS 0.09fF
C46 a_3924_210.n2 VSS 0.13fF
C47 a_3924_210.n3 VSS 0.11fF
C48 a_3924_210.n4 VSS 0.02fF
C49 a_3924_210.n5 VSS 0.03fF
C50 a_3924_210.n6 VSS 0.02fF
C51 a_3924_210.n7 VSS 0.05fF
C52 a_3924_210.n8 VSS 0.03fF
C53 a_3924_210.n9 VSS 0.11fF
C54 a_3924_210.n10 VSS 0.06fF
C55 a_3924_210.n11 VSS 0.01fF
C56 a_3924_210.t0 VSS 0.33fF
C57 a_91_103.n0 VSS 0.10fF
C58 a_91_103.n1 VSS 0.04fF
C59 a_91_103.n2 VSS 0.03fF
C60 a_91_103.n3 VSS 0.03fF
C61 a_91_103.n4 VSS 0.05fF
C62 a_91_103.n5 VSS 0.08fF
C63 a_91_103.n6 VSS 0.07fF
C64 a_3829_1050.n0 VSS 0.46fF
C65 a_3829_1050.n1 VSS 0.46fF
C66 a_3829_1050.n2 VSS 0.32fF
C67 a_3829_1050.n3 VSS 0.49fF
C68 a_3829_1050.n4 VSS 0.03fF
C69 a_3829_1050.n5 VSS 0.05fF
C70 a_3829_1050.n6 VSS 0.03fF
C71 a_3829_1050.n7 VSS 0.26fF
C72 a_3829_1050.n8 VSS 0.54fF
C73 a_3829_1050.n9 VSS 0.26fF
C74 a_3829_1050.n10 VSS 0.17fF
C75 a_3829_1050.n11 VSS 0.54fF
C76 a_2962_210.n0 VSS 0.02fF
C77 a_2962_210.n1 VSS 0.09fF
C78 a_2962_210.n2 VSS 0.13fF
C79 a_2962_210.n3 VSS 0.11fF
C80 a_2962_210.t1 VSS 0.30fF
C81 a_2962_210.n4 VSS 0.09fF
C82 a_2962_210.n5 VSS 0.06fF
C83 a_2962_210.n6 VSS 0.01fF
C84 a_2962_210.n7 VSS 0.03fF
C85 a_2962_210.n8 VSS 0.11fF
C86 a_2962_210.n9 VSS 0.02fF
C87 a_2962_210.n10 VSS 0.05fF
C88 a_2962_210.n11 VSS 0.02fF
C89 a_372_210.n0 VSS 0.02fF
C90 a_372_210.n1 VSS 0.09fF
C91 a_372_210.n2 VSS 0.13fF
C92 a_372_210.n3 VSS 0.11fF
C93 a_372_210.t1 VSS 0.30fF
C94 a_372_210.n4 VSS 0.09fF
C95 a_372_210.n5 VSS 0.06fF
C96 a_372_210.n6 VSS 0.01fF
C97 a_372_210.n7 VSS 0.03fF
C98 a_372_210.n8 VSS 0.11fF
C99 a_372_210.n9 VSS 0.02fF
C100 a_372_210.n10 VSS 0.05fF
C101 a_372_210.n11 VSS 0.02fF
C102 a_599_989.n0 VSS 0.57fF
C103 a_599_989.n1 VSS 0.57fF
C104 a_599_989.n2 VSS 0.40fF
C105 a_599_989.n3 VSS 0.42fF
C106 a_599_989.n4 VSS 0.40fF
C107 a_599_989.t7 VSS 0.57fF
C108 a_599_989.n5 VSS 0.42fF
C109 a_599_989.n6 VSS 1.32fF
C110 a_599_989.n7 VSS 0.04fF
C111 a_599_989.n8 VSS 0.06fF
C112 a_599_989.n9 VSS 0.04fF
C113 a_599_989.n10 VSS 0.32fF
C114 a_599_989.n11 VSS 0.48fF
C115 a_599_989.n12 VSS 0.32fF
C116 a_599_989.n13 VSS 0.21fF
C117 a_599_989.n14 VSS 0.67fF
C118 a_277_1050.n0 VSS 0.74fF
C119 a_277_1050.n1 VSS 0.74fF
C120 a_277_1050.n2 VSS 0.42fF
C121 a_277_1050.n3 VSS 0.83fF
C122 a_277_1050.n4 VSS 0.42fF
C123 a_277_1050.n5 VSS 0.66fF
C124 a_277_1050.n6 VSS 3.24fF
C125 a_277_1050.n7 VSS 0.59fF
C126 a_277_1050.n8 VSS 0.66fF
C127 a_277_1050.n9 VSS 0.38fF
C128 a_277_1050.n10 VSS 0.27fF
C129 a_277_1050.n11 VSS 0.87fF
C130 Q.n0 VSS 0.54fF
C131 Q.n1 VSS 0.64fF
C132 Q.n2 VSS 0.28fF
C133 Q.n3 VSS 0.04fF
C134 Q.n4 VSS 0.05fF
C135 Q.n5 VSS 0.03fF
C136 Q.n6 VSS 0.34fF
C137 Q.n7 VSS 0.43fF
C138 Q.n8 VSS 0.35fF
C139 Q.t6 VSS 0.57fF
C140 Q.n9 VSS 0.39fF
C141 Q.n10 VSS 0.03fF
C142 VDD.n0 VSS 0.15fF
C143 VDD.n1 VSS 0.02fF
C144 VDD.n2 VSS 0.02fF
C145 VDD.n3 VSS 0.04fF
C146 VDD.n4 VSS 0.01fF
C147 VDD.n6 VSS 0.02fF
C148 VDD.n7 VSS 0.02fF
C149 VDD.n8 VSS 0.02fF
C150 VDD.n9 VSS 0.02fF
C151 VDD.n11 VSS 0.02fF
C152 VDD.n14 VSS 0.45fF
C153 VDD.n16 VSS 0.03fF
C154 VDD.n17 VSS 0.02fF
C155 VDD.n18 VSS 0.02fF
C156 VDD.n19 VSS 0.02fF
C157 VDD.n20 VSS 0.04fF
C158 VDD.n21 VSS 0.27fF
C159 VDD.n22 VSS 0.02fF
C160 VDD.n23 VSS 0.03fF
C161 VDD.n24 VSS 0.14fF
C162 VDD.n25 VSS 0.17fF
C163 VDD.n26 VSS 0.01fF
C164 VDD.n27 VSS 0.11fF
C165 VDD.n28 VSS 0.03fF
C166 VDD.n29 VSS 0.30fF
C167 VDD.n30 VSS 0.01fF
C168 VDD.n31 VSS 0.02fF
C169 VDD.n32 VSS 0.02fF
C170 VDD.n33 VSS 0.06fF
C171 VDD.n34 VSS 0.24fF
C172 VDD.n35 VSS 0.01fF
C173 VDD.n36 VSS 0.01fF
C174 VDD.n37 VSS 0.00fF
C175 VDD.n38 VSS 0.09fF
C176 VDD.n39 VSS 0.03fF
C177 VDD.n40 VSS 0.17fF
C178 VDD.n41 VSS 0.14fF
C179 VDD.n42 VSS 0.01fF
C180 VDD.n43 VSS 0.02fF
C181 VDD.n44 VSS 0.03fF
C182 VDD.n45 VSS 0.14fF
C183 VDD.n46 VSS 0.16fF
C184 VDD.n47 VSS 0.01fF
C185 VDD.n48 VSS 0.02fF
C186 VDD.n49 VSS 0.02fF
C187 VDD.n50 VSS 0.06fF
C188 VDD.n51 VSS 0.25fF
C189 VDD.n52 VSS 0.01fF
C190 VDD.n53 VSS 0.01fF
C191 VDD.n54 VSS 0.02fF
C192 VDD.n55 VSS 0.27fF
C193 VDD.n56 VSS 0.01fF
C194 VDD.n57 VSS 0.02fF
C195 VDD.n58 VSS 0.03fF
C196 VDD.n59 VSS 0.02fF
C197 VDD.n60 VSS 0.02fF
C198 VDD.n61 VSS 0.02fF
C199 VDD.n62 VSS 0.26fF
C200 VDD.n63 VSS 0.04fF
C201 VDD.n64 VSS 0.04fF
C202 VDD.n65 VSS 0.02fF
C203 VDD.n67 VSS 0.02fF
C204 VDD.n68 VSS 0.02fF
C205 VDD.n69 VSS 0.02fF
C206 VDD.n70 VSS 0.02fF
C207 VDD.n72 VSS 0.02fF
C208 VDD.n73 VSS 0.02fF
C209 VDD.n74 VSS 0.02fF
C210 VDD.n76 VSS 0.27fF
C211 VDD.n78 VSS 0.02fF
C212 VDD.n79 VSS 0.02fF
C213 VDD.n80 VSS 0.03fF
C214 VDD.n81 VSS 0.02fF
C215 VDD.n82 VSS 0.27fF
C216 VDD.n83 VSS 0.01fF
C217 VDD.n84 VSS 0.02fF
C218 VDD.n85 VSS 0.03fF
C219 VDD.n86 VSS 0.27fF
C220 VDD.n87 VSS 0.01fF
C221 VDD.n88 VSS 0.02fF
C222 VDD.n89 VSS 0.02fF
C223 VDD.n90 VSS 0.22fF
C224 VDD.n91 VSS 0.01fF
C225 VDD.n92 VSS 0.07fF
C226 VDD.n93 VSS 0.02fF
C227 VDD.n94 VSS 0.14fF
C228 VDD.n95 VSS 0.17fF
C229 VDD.n96 VSS 0.01fF
C230 VDD.n97 VSS 0.02fF
C231 VDD.n98 VSS 0.02fF
C232 VDD.n99 VSS 0.14fF
C233 VDD.n100 VSS 0.16fF
C234 VDD.n101 VSS 0.01fF
C235 VDD.n102 VSS 0.11fF
C236 VDD.n103 VSS 0.02fF
C237 VDD.n104 VSS 0.02fF
C238 VDD.n105 VSS 0.02fF
C239 VDD.n106 VSS 0.17fF
C240 VDD.n107 VSS 0.14fF
C241 VDD.n108 VSS 0.01fF
C242 VDD.n109 VSS 0.02fF
C243 VDD.n110 VSS 0.03fF
C244 VDD.n111 VSS 0.18fF
C245 VDD.n112 VSS 0.15fF
C246 VDD.n113 VSS 0.01fF
C247 VDD.n114 VSS 0.02fF
C248 VDD.n115 VSS 0.03fF
C249 VDD.n116 VSS 0.11fF
C250 VDD.n117 VSS 0.02fF
C251 VDD.n118 VSS 0.14fF
C252 VDD.n119 VSS 0.15fF
C253 VDD.n120 VSS 0.01fF
C254 VDD.n121 VSS 0.02fF
C255 VDD.n122 VSS 0.02fF
C256 VDD.n123 VSS 0.14fF
C257 VDD.n124 VSS 0.17fF
C258 VDD.n125 VSS 0.01fF
C259 VDD.n126 VSS 0.02fF
C260 VDD.n127 VSS 0.02fF
C261 VDD.n128 VSS 0.06fF
C262 VDD.n129 VSS 0.22fF
C263 VDD.n130 VSS 0.01fF
C264 VDD.n131 VSS 0.01fF
C265 VDD.n132 VSS 0.02fF
C266 VDD.n133 VSS 0.27fF
C267 VDD.n134 VSS 0.01fF
C268 VDD.n135 VSS 0.02fF
C269 VDD.n136 VSS 0.02fF
C270 VDD.n137 VSS 0.27fF
C271 VDD.n138 VSS 0.01fF
C272 VDD.n139 VSS 0.02fF
C273 VDD.n140 VSS 0.03fF
C274 VDD.n141 VSS 0.02fF
C275 VDD.n142 VSS 0.02fF
C276 VDD.n143 VSS 0.02fF
C277 VDD.n144 VSS 0.31fF
C278 VDD.n145 VSS 0.04fF
C279 VDD.n146 VSS 0.03fF
C280 VDD.n147 VSS 0.02fF
C281 VDD.n148 VSS 0.02fF
C282 VDD.n149 VSS 0.02fF
C283 VDD.n150 VSS 0.02fF
C284 VDD.n151 VSS 0.02fF
C285 VDD.n153 VSS 0.02fF
C286 VDD.n154 VSS 0.02fF
C287 VDD.n155 VSS 0.02fF
C288 VDD.n157 VSS 0.27fF
C289 VDD.n159 VSS 0.02fF
C290 VDD.n160 VSS 0.02fF
C291 VDD.n161 VSS 0.03fF
C292 VDD.n162 VSS 0.02fF
C293 VDD.n163 VSS 0.27fF
C294 VDD.n164 VSS 0.01fF
C295 VDD.n165 VSS 0.02fF
C296 VDD.n166 VSS 0.03fF
C297 VDD.n167 VSS 0.27fF
C298 VDD.n168 VSS 0.01fF
C299 VDD.n169 VSS 0.02fF
C300 VDD.n170 VSS 0.02fF
C301 VDD.n171 VSS 0.22fF
C302 VDD.n172 VSS 0.01fF
C303 VDD.n173 VSS 0.07fF
C304 VDD.n174 VSS 0.02fF
C305 VDD.n175 VSS 0.14fF
C306 VDD.n176 VSS 0.17fF
C307 VDD.n177 VSS 0.01fF
C308 VDD.n178 VSS 0.02fF
C309 VDD.n179 VSS 0.02fF
C310 VDD.n180 VSS 0.14fF
C311 VDD.n181 VSS 0.16fF
C312 VDD.n182 VSS 0.01fF
C313 VDD.n183 VSS 0.11fF
C314 VDD.n184 VSS 0.02fF
C315 VDD.n185 VSS 0.02fF
C316 VDD.n186 VSS 0.02fF
C317 VDD.n187 VSS 0.17fF
C318 VDD.n188 VSS 0.14fF
C319 VDD.n189 VSS 0.01fF
C320 VDD.n190 VSS 0.02fF
C321 VDD.n191 VSS 0.03fF
C322 VDD.n192 VSS 0.18fF
C323 VDD.n193 VSS 0.15fF
C324 VDD.n194 VSS 0.01fF
C325 VDD.n195 VSS 0.02fF
C326 VDD.n196 VSS 0.03fF
C327 VDD.n197 VSS 0.11fF
C328 VDD.n198 VSS 0.02fF
C329 VDD.n199 VSS 0.14fF
C330 VDD.n200 VSS 0.15fF
C331 VDD.n201 VSS 0.01fF
C332 VDD.n202 VSS 0.02fF
C333 VDD.n203 VSS 0.02fF
C334 VDD.n204 VSS 0.14fF
C335 VDD.n205 VSS 0.17fF
C336 VDD.n206 VSS 0.01fF
C337 VDD.n207 VSS 0.02fF
C338 VDD.n208 VSS 0.02fF
C339 VDD.n209 VSS 0.06fF
C340 VDD.n210 VSS 0.22fF
C341 VDD.n211 VSS 0.01fF
C342 VDD.n212 VSS 0.01fF
C343 VDD.n213 VSS 0.02fF
C344 VDD.n214 VSS 0.27fF
C345 VDD.n215 VSS 0.01fF
C346 VDD.n216 VSS 0.02fF
C347 VDD.n217 VSS 0.02fF
C348 VDD.n218 VSS 0.27fF
C349 VDD.n219 VSS 0.01fF
C350 VDD.n220 VSS 0.02fF
C351 VDD.n221 VSS 0.03fF
C352 VDD.n222 VSS 0.02fF
C353 VDD.n223 VSS 0.02fF
C354 VDD.n224 VSS 0.02fF
C355 VDD.n225 VSS 0.26fF
C356 VDD.n226 VSS 0.04fF
C357 VDD.n227 VSS 0.03fF
C358 VDD.n228 VSS 0.02fF
C359 VDD.n229 VSS 0.02fF
C360 VDD.n230 VSS 0.02fF
C361 VDD.n231 VSS 0.02fF
C362 VDD.n232 VSS 0.02fF
C363 VDD.n234 VSS 0.02fF
C364 VDD.n235 VSS 0.02fF
C365 VDD.n236 VSS 0.02fF
C366 VDD.n238 VSS 0.27fF
C367 VDD.n240 VSS 0.02fF
C368 VDD.n241 VSS 0.02fF
C369 VDD.n242 VSS 0.03fF
C370 VDD.n243 VSS 0.02fF
C371 VDD.n244 VSS 0.27fF
C372 VDD.n245 VSS 0.01fF
C373 VDD.n246 VSS 0.02fF
C374 VDD.n247 VSS 0.03fF
C375 VDD.n248 VSS 0.06fF
C376 VDD.n249 VSS 0.24fF
C377 VDD.n250 VSS 0.01fF
C378 VDD.n251 VSS 0.01fF
C379 VDD.n252 VSS 0.02fF
C380 VDD.n253 VSS 0.14fF
C381 VDD.n254 VSS 0.17fF
C382 VDD.n255 VSS 0.01fF
C383 VDD.n256 VSS 0.02fF
C384 VDD.n257 VSS 0.02fF
C385 VDD.n258 VSS 0.11fF
C386 VDD.n259 VSS 0.03fF
C387 VDD.n260 VSS 0.30fF
C388 VDD.n261 VSS 0.01fF
C389 VDD.n262 VSS 0.02fF
C390 VDD.n263 VSS 0.03fF
C391 VDD.n264 VSS 0.17fF
C392 VDD.n265 VSS 0.14fF
C393 VDD.n266 VSS 0.01fF
C394 VDD.n267 VSS 0.02fF
C395 VDD.n268 VSS 0.03fF
C396 VDD.n269 VSS 0.14fF
C397 VDD.n270 VSS 0.16fF
C398 VDD.n271 VSS 0.01fF
C399 VDD.n272 VSS 0.02fF
C400 VDD.n273 VSS 0.02fF
C401 VDD.n274 VSS 0.06fF
C402 VDD.n275 VSS 0.25fF
C403 VDD.n276 VSS 0.01fF
C404 VDD.n277 VSS 0.01fF
C405 VDD.n278 VSS 0.02fF
C406 VDD.n279 VSS 0.27fF
C407 VDD.n280 VSS 0.01fF
C408 VDD.n281 VSS 0.02fF
C409 VDD.n282 VSS 0.03fF
C410 VDD.n283 VSS 0.02fF
C411 VDD.n284 VSS 0.02fF
C412 VDD.n285 VSS 0.02fF
C413 VDD.n286 VSS 0.26fF
C414 VDD.n287 VSS 0.04fF
C415 VDD.n288 VSS 0.03fF
C416 VDD.n289 VSS 0.02fF
C417 VDD.n290 VSS 0.02fF
C418 VDD.n291 VSS 0.02fF
C419 VDD.n292 VSS 0.02fF
C420 VDD.n293 VSS 0.02fF
C421 VDD.n295 VSS 0.02fF
C422 VDD.n296 VSS 0.02fF
C423 VDD.n297 VSS 0.02fF
C424 VDD.n299 VSS 0.27fF
C425 VDD.n301 VSS 0.02fF
C426 VDD.n302 VSS 0.02fF
C427 VDD.n303 VSS 0.03fF
C428 VDD.n304 VSS 0.02fF
C429 VDD.n305 VSS 0.27fF
C430 VDD.n306 VSS 0.01fF
C431 VDD.n307 VSS 0.02fF
C432 VDD.n308 VSS 0.03fF
C433 VDD.n309 VSS 0.27fF
C434 VDD.n310 VSS 0.01fF
C435 VDD.n311 VSS 0.02fF
C436 VDD.n312 VSS 0.02fF
C437 VDD.n313 VSS 0.22fF
C438 VDD.n314 VSS 0.01fF
C439 VDD.n315 VSS 0.07fF
C440 VDD.n316 VSS 0.02fF
C441 VDD.n317 VSS 0.14fF
C442 VDD.n318 VSS 0.17fF
C443 VDD.n319 VSS 0.01fF
C444 VDD.n320 VSS 0.02fF
C445 VDD.n321 VSS 0.02fF
C446 VDD.n322 VSS 0.14fF
C447 VDD.n323 VSS 0.16fF
C448 VDD.n324 VSS 0.01fF
C449 VDD.n325 VSS 0.11fF
C450 VDD.n326 VSS 0.02fF
C451 VDD.n327 VSS 0.02fF
C452 VDD.n328 VSS 0.02fF
C453 VDD.n329 VSS 0.17fF
C454 VDD.n330 VSS 0.14fF
C455 VDD.n331 VSS 0.01fF
C456 VDD.n332 VSS 0.02fF
C457 VDD.n333 VSS 0.03fF
C458 VDD.n334 VSS 0.18fF
C459 VDD.n335 VSS 0.15fF
C460 VDD.n336 VSS 0.01fF
C461 VDD.n337 VSS 0.02fF
C462 VDD.n338 VSS 0.03fF
C463 VDD.n339 VSS 0.11fF
C464 VDD.n340 VSS 0.02fF
C465 VDD.n341 VSS 0.14fF
C466 VDD.n342 VSS 0.15fF
C467 VDD.n343 VSS 0.01fF
C468 VDD.n344 VSS 0.02fF
C469 VDD.n345 VSS 0.02fF
C470 VDD.n346 VSS 0.14fF
C471 VDD.n347 VSS 0.17fF
C472 VDD.n348 VSS 0.01fF
C473 VDD.n349 VSS 0.02fF
C474 VDD.n350 VSS 0.02fF
C475 VDD.n351 VSS 0.06fF
C476 VDD.n352 VSS 0.22fF
C477 VDD.n353 VSS 0.01fF
C478 VDD.n354 VSS 0.01fF
C479 VDD.n355 VSS 0.02fF
C480 VDD.n356 VSS 0.27fF
C481 VDD.n357 VSS 0.01fF
C482 VDD.n358 VSS 0.02fF
C483 VDD.n359 VSS 0.02fF
C484 VDD.n360 VSS 0.27fF
C485 VDD.n361 VSS 0.01fF
C486 VDD.n362 VSS 0.02fF
C487 VDD.n363 VSS 0.03fF
C488 VDD.n364 VSS 0.02fF
C489 VDD.n365 VSS 0.02fF
C490 VDD.n366 VSS 0.02fF
C491 VDD.n367 VSS 0.02fF
C492 VDD.n368 VSS 0.02fF
C493 VDD.n369 VSS 0.02fF
C494 VDD.n371 VSS 0.02fF
C495 VDD.n372 VSS 0.02fF
C496 VDD.n373 VSS 0.02fF
C497 VDD.n374 VSS 0.02fF
C498 VDD.n376 VSS 0.04fF
C499 VDD.n377 VSS 0.02fF
C500 VDD.n378 VSS 0.31fF
C501 VDD.n379 VSS 0.04fF
C502 VDD.n381 VSS 0.27fF
C503 VDD.n383 VSS 0.02fF
C504 VDD.n384 VSS 0.02fF
C505 VDD.n385 VSS 0.03fF
C506 VDD.n386 VSS 0.02fF
C507 VDD.n387 VSS 0.27fF
C508 VDD.n388 VSS 0.01fF
C509 VDD.n389 VSS 0.02fF
C510 VDD.n390 VSS 0.03fF
C511 VDD.n391 VSS 0.27fF
C512 VDD.n392 VSS 0.01fF
C513 VDD.n393 VSS 0.02fF
C514 VDD.n394 VSS 0.02fF
C515 VDD.n395 VSS 0.22fF
C516 VDD.n396 VSS 0.01fF
C517 VDD.n397 VSS 0.07fF
C518 VDD.n398 VSS 0.02fF
C519 VDD.n399 VSS 0.14fF
C520 VDD.n400 VSS 0.17fF
C521 VDD.n401 VSS 0.01fF
C522 VDD.n402 VSS 0.02fF
C523 VDD.n403 VSS 0.02fF
C524 VDD.n404 VSS 0.14fF
C525 VDD.n405 VSS 0.16fF
C526 VDD.n406 VSS 0.01fF
C527 VDD.n407 VSS 0.11fF
C528 VDD.n408 VSS 0.02fF
C529 VDD.n409 VSS 0.02fF
C530 VDD.n410 VSS 0.02fF
C531 VDD.n411 VSS 0.17fF
C532 VDD.n412 VSS 0.14fF
C533 VDD.n413 VSS 0.01fF
C534 VDD.n414 VSS 0.02fF
C535 VDD.n415 VSS 0.03fF
C536 VDD.n416 VSS 0.18fF
C537 VDD.n417 VSS 0.15fF
C538 VDD.n418 VSS 0.01fF
C539 VDD.n419 VSS 0.02fF
C540 VDD.n420 VSS 0.03fF
C541 VDD.n421 VSS 0.11fF
C542 VDD.n422 VSS 0.02fF
C543 VDD.n423 VSS 0.14fF
C544 VDD.n424 VSS 0.15fF
C545 VDD.n425 VSS 0.01fF
C546 VDD.n426 VSS 0.02fF
C547 VDD.n427 VSS 0.02fF
C548 VDD.n428 VSS 0.14fF
C549 VDD.n429 VSS 0.17fF
C550 VDD.n430 VSS 0.01fF
C551 VDD.n431 VSS 0.02fF
C552 VDD.n432 VSS 0.02fF
C553 VDD.n433 VSS 0.06fF
C554 VDD.n434 VSS 0.22fF
C555 VDD.n435 VSS 0.01fF
C556 VDD.n436 VSS 0.01fF
C557 VDD.n437 VSS 0.02fF
C558 VDD.n438 VSS 0.27fF
C559 VDD.n439 VSS 0.01fF
C560 VDD.n440 VSS 0.02fF
C561 VDD.n441 VSS 0.02fF
C562 VDD.n442 VSS 0.02fF
C563 VDD.n443 VSS 0.02fF
C564 VDD.n444 VSS 0.02fF
C565 VDD.n445 VSS 0.20fF
C566 VDD.n446 VSS 0.03fF
C567 VDD.n447 VSS 0.02fF
C568 VDD.n448 VSS 0.02fF
C569 VDD.n449 VSS 0.02fF
C570 VDD.n450 VSS 0.02fF
C571 VDD.n451 VSS 0.02fF
C572 VDD.n453 VSS 0.02fF
C573 VDD.n454 VSS 0.02fF
C574 VDD.n455 VSS 0.02fF
C575 VDD.n457 VSS 0.45fF
C576 VDD.n459 VSS 0.03fF
C577 VDD.n460 VSS 0.04fF
C578 VDD.n461 VSS 0.27fF
C579 VDD.n462 VSS 0.02fF
C580 VDD.n463 VSS 0.03fF
C581 VDD.n464 VSS 0.01fF
C582 RN.n0 VSS 0.39fF
C583 RN.t6 VSS 0.35fF
C584 RN.n1 VSS 0.30fF
C585 RN.n2 VSS 0.38fF
C586 RN.t1 VSS 0.36fF
C587 RN.n3 VSS 0.29fF
C588 RN.n4 VSS 1.05fF
C589 RN.n5 VSS 0.38fF
C590 RN.t4 VSS 0.37fF
C591 RN.n6 VSS 0.29fF
C592 RN.n7 VSS 0.55fF
C593 a_2141_1050.n0 VSS 0.52fF
C594 a_2141_1050.n1 VSS 0.61fF
C595 a_2141_1050.n2 VSS 0.30fF
C596 a_2141_1050.n3 VSS 0.33fF
C597 a_2141_1050.n4 VSS 0.64fF
C598 a_2141_1050.n5 VSS 0.60fF
C599 a_2141_1050.n6 VSS 0.08fF
C600 a_2141_1050.n7 VSS 0.28fF
C601 a_2141_1050.n8 VSS 0.04fF
C602 a_2036_101.n0 VSS 0.08fF
C603 a_2036_101.n1 VSS 0.02fF
C604 a_2036_101.n2 VSS 0.01fF
C605 a_2036_101.n3 VSS 0.06fF
C606 a_2036_101.n4 VSS 0.10fF
C607 a_2036_101.n5 VSS 0.06fF
C608 a_2036_101.n6 VSS 0.05fF
C609 a_147_187.n0 VSS 0.06fF
C610 a_147_187.n1 VSS 0.73fF
C611 a_147_187.n2 VSS 0.73fF
C612 a_147_187.n3 VSS 0.86fF
C613 a_147_187.n4 VSS 0.27fF
C614 a_147_187.n5 VSS 0.33fF
C615 a_147_187.n6 VSS 0.38fF
C616 a_147_187.n7 VSS 0.58fF
C617 a_147_187.n8 VSS 0.38fF
C618 a_147_187.t7 VSS 0.81fF
C619 a_147_187.n9 VSS 0.52fF
C620 a_147_187.n10 VSS 0.37fF
C621 a_147_187.n11 VSS 0.77fF
C622 a_147_187.n12 VSS 2.88fF
C623 a_147_187.n13 VSS 2.27fF
C624 a_147_187.n14 VSS 0.62fF
C625 a_147_187.n15 VSS 0.06fF
C626 a_147_187.n16 VSS 0.50fF
C627 a_147_187.n17 VSS 0.06fF
.ends
