* SPICE3 file created from TMRDFFRNQX1.ext - technology: sky130A

.subckt TMRDFFRNQX1 Q D CLK RN VDD GND
X0 VDD a_5457_1004 a_9009_1004 VDD pshort w=2 l=0.15 M=2
X1 a_9331_943 a_9009_1004 VDD VDD pshort w=2 l=0.15 M=2
X2 VDD CLK a_277_1004 VDD pshort w=2 l=0.15 M=2
X3 VDD a_277_1004 a_147_159 VDD pshort w=2 l=0.15 M=2
X4 VDD a_5457_1004 a_5779_943 VDD pshort w=2 l=0.15 M=2
X5 VDD RN a_5779_943 VDD pshort w=2 l=0.15 M=2
X6 VDD a_9331_943 a_9009_1004 VDD pshort w=2 l=0.15 M=2
X7 VDD CLK a_10637_1004 VDD pshort w=2 l=0.15 M=2
X8 GND a_9009_1004 a_9806_73 GND nshort w=3 l=0.15
X9 VDD CLK a_10507_159 VDD pshort w=2 l=0.15 M=2
X10 a_9331_943 a_5327_159 VDD VDD pshort w=2 l=0.15 M=2
X11 GND a_5779_943 a_7216_73 GND nshort w=3 l=0.15
X12 GND a_147_159 a_91_75 GND nshort w=3 l=0.15
X13 a_10507_159 RN VDD VDD pshort w=2 l=0.15 M=2
X14 a_9331_943 D VDD VDD pshort w=2 l=0.15 M=2
X15 a_147_159 a_4151_943 VDD VDD pshort w=2 l=0.15 M=2
X16 a_599_943 RN VDD VDD pshort w=2 l=0.15 M=2
X17 GND a_7321_1004 a_7861_75 GND nshort w=3 l=0.15
X18 a_10637_1004 a_10507_159 VDD VDD pshort w=2 l=0.15 M=2
X19 VDD a_14511_943 a_15757_1005 VDD pshort w=2 l=0.15 M=2
X20 a_147_159 CLK VDD VDD pshort w=2 l=0.15 M=2
X21 a_147_159 a_4151_943 a_3924_182 GND nshort w=3 l=0.15
X22 GND a_5327_159 a_5271_75 GND nshort w=3 l=0.15
X23 a_4151_943 a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X24 a_10507_159 RN a_13322_182 GND nshort w=3 l=0.15
X25 a_9331_943 a_10507_159 a_12396_73 GND nshort w=3 l=0.15
X26 a_15757_1005 a_9331_943 VDD VDD pshort w=2 l=0.15 M=2
X27 VDD a_10507_159 a_14511_943 VDD pshort w=2 l=0.15 M=2
X28 a_9331_943 a_5327_159 a_9806_73 GND nshort w=3 l=0.15
X29 VDD a_9331_943 a_9331_943 VDD pshort w=2 l=0.15 M=2
X30 VDD a_147_159 a_2141_1004 VDD pshort w=2 l=0.15 M=2
X31 VDD a_599_943 a_277_1004 VDD pshort w=2 l=0.15 M=2
X32 VDD D a_5779_943 VDD pshort w=2 l=0.15 M=2
X33 VDD RN a_9009_1004 VDD pshort w=2 l=0.15 M=2
X34 a_6514_182 D a_6233_75 GND nshort w=3 l=0.15
X35 VDD a_5327_159 a_5457_1004 VDD pshort w=2 l=0.15 M=2
X36 VDD a_7321_1004 a_5327_159 VDD pshort w=2 l=0.15 M=2
X37 VDD a_2141_1004 a_147_159 VDD pshort w=2 l=0.15 M=2
X38 a_10507_159 a_14511_943 VDD VDD pshort w=2 l=0.15 M=2
X39 a_9331_943 RN VDD VDD pshort w=2 l=0.15 M=2
X40 a_10507_159 a_14511_943 a_14284_182 GND nshort w=3 l=0.15
X41 a_147_159 RN VDD VDD pshort w=2 l=0.15 M=2
X42 a_7321_1004 a_5327_159 VDD VDD pshort w=2 l=0.15 M=2
X43 GND a_9331_943 a_13041_75 GND nshort w=3 l=0.15
X44 a_15932_181 a_4151_943 a_16421_1005 VDD pshort w=2 l=0.15 M=2
X45 a_372_182 CLK a_91_75 GND nshort w=3 l=0.15
X46 GND a_277_1004 a_3643_75 GND nshort w=3 l=0.15
X47 VDD a_9331_943 a_10637_1004 VDD pshort w=2 l=0.15 M=2
X48 VDD a_10507_159 a_9331_943 VDD pshort w=2 l=0.15 M=2
X49 a_5552_182 CLK a_5271_75 GND nshort w=3 l=0.15
X50 a_15932_181 a_4151_943 a_16318_73 GND nshort w=3 l=0.15
X51 VDD a_15932_181 Q VDD pshort w=2 l=0.15 M=2
X52 a_277_1004 a_147_159 VDD VDD pshort w=2 l=0.15 M=2
X53 a_16421_1005 a_4151_943 a_15757_1005 VDD pshort w=2 l=0.15 M=2
X54 GND a_147_159 a_4626_73 GND nshort w=3 l=0.15
X55 a_10507_159 a_9331_943 VDD VDD pshort w=2 l=0.15 M=2
X56 a_7321_1004 a_5779_943 VDD VDD pshort w=2 l=0.15 M=2
X57 VDD a_277_1004 a_599_943 VDD pshort w=2 l=0.15 M=2
X58 GND a_599_943 a_2036_73 GND nshort w=3 l=0.15
X59 GND a_10637_1004 a_14003_75 GND nshort w=3 l=0.15
X60 GND a_2141_1004 a_2681_75 GND nshort w=3 l=0.15
X61 a_599_943 RN a_1334_182 GND nshort w=3 l=0.15
X62 a_15932_181 a_14511_943 a_16421_1005 VDD pshort w=2 l=0.15 M=2
X63 a_10637_1004 a_9331_943 a_10732_182 GND nshort w=3 l=0.15
X64 a_13322_182 CLK a_13041_75 GND nshort w=3 l=0.15
X65 Q a_15932_181 GND GND nshort w=3 l=0.15
X66 a_3924_182 RN a_3643_75 GND nshort w=3 l=0.15
X67 VDD a_5779_943 a_5457_1004 VDD pshort w=2 l=0.15 M=2
X68 VDD RN a_5327_159 VDD pshort w=2 l=0.15 M=2
X69 a_7321_1004 a_5327_159 a_7216_73 GND nshort w=3 l=0.15
X70 a_2141_1004 a_599_943 VDD VDD pshort w=2 l=0.15 M=2
X71 GND a_9331_943 a_15652_73 GND nshort w=3 l=0.15
X72 a_16421_1005 a_9331_943 a_15757_1005 VDD pshort w=2 l=0.15 M=2
X73 GND a_10507_159 a_14986_73 GND nshort w=3 l=0.15
X74 a_9331_943 RN a_11694_182 GND nshort w=3 l=0.15
X75 VDD a_10637_1004 a_10507_159 VDD pshort w=2 l=0.15 M=2
X76 VDD a_10637_1004 a_9331_943 VDD pshort w=2 l=0.15 M=2
X77 VDD D a_599_943 VDD pshort w=2 l=0.15 M=2
X78 a_9009_1004 a_9331_943 a_9104_182 GND nshort w=3 l=0.15
X79 GND a_277_1004 a_1053_75 GND nshort w=3 l=0.15
X80 a_14284_182 RN a_14003_75 GND nshort w=3 l=0.15
X81 a_2962_182 CLK a_2681_75 GND nshort w=3 l=0.15
X82 VDD CLK a_5457_1004 VDD pshort w=2 l=0.15 M=2
X83 VDD CLK a_5327_159 VDD pshort w=2 l=0.15 M=2
X84 GND a_4151_943 a_16984_73 GND nshort w=3 l=0.15
X85 GND a_10637_1004 a_11413_75 GND nshort w=3 l=0.15
X86 a_5327_159 RN a_8142_182 GND nshort w=3 l=0.15
X87 a_4151_943 a_147_159 a_4626_73 GND nshort w=3 l=0.15
X88 a_1334_182 D a_1053_75 GND nshort w=3 l=0.15
X89 GND a_9331_943 a_12396_73 GND nshort w=3 l=0.15
X90 a_2141_1004 a_147_159 a_2036_73 GND nshort w=3 l=0.15
X91 GND a_10507_159 a_10451_75 GND nshort w=3 l=0.15
X92 a_15932_181 a_14511_943 a_15652_73 GND nshort w=3 l=0.15
X93 a_5779_943 RN a_6514_182 GND nshort w=3 l=0.15
X94 a_11694_182 D a_11413_75 GND nshort w=3 l=0.15
X95 a_14511_943 a_10507_159 a_14986_73 GND nshort w=3 l=0.15
X96 a_9104_182 RN a_8823_75 GND nshort w=3 l=0.15
X97 GND a_9331_943 a_16318_73 GND nshort w=3 l=0.15
X98 a_277_1004 a_599_943 a_372_182 GND nshort w=3 l=0.15
X99 a_10732_182 CLK a_10451_75 GND nshort w=3 l=0.15
X100 GND a_5457_1004 a_8823_75 GND nshort w=3 l=0.15
X101 GND a_5457_1004 a_6233_75 GND nshort w=3 l=0.15
X102 a_5457_1004 a_5779_943 a_5552_182 GND nshort w=3 l=0.15
X103 a_15932_181 a_14511_943 a_16984_73 GND nshort w=3 l=0.15
X104 a_147_159 RN a_2962_182 GND nshort w=3 l=0.15
X105 a_8142_182 CLK a_7861_75 GND nshort w=3 l=0.15
C0 VDD a_5779_943 2.36fF
C1 a_5457_1004 VDD 2.55fF
C2 VDD a_5327_159 3.67fF
C3 a_10637_1004 a_10507_159 3.69fF
C4 a_10507_159 a_9331_943 2.98fF
C5 a_147_159 CLK 5.49fF
C6 a_14511_943 a_9331_943 2.50fF
C7 a_4151_943 VDD 2.71fF
C8 CLK a_5327_159 5.65fF
C9 a_147_159 a_277_1004 3.68fF
C10 RN VDD 2.46fF
C11 CLK VDD 5.84fF
C12 D a_4151_943 8.50fF
C13 a_599_943 a_277_1004 2.06fF
C14 VDD a_10637_1004 2.55fF
C15 VDD a_9331_943 6.51fF
C16 RN a_4151_943 4.25fF
C17 VDD a_10507_159 5.91fF
C18 RN D 11.85fF
C19 a_277_1004 VDD 2.39fF
C20 a_4151_943 a_9331_943 7.52fF
C21 a_14511_943 VDD 2.40fF
C22 RN CLK 2.13fF
C23 a_147_159 VDD 5.76fF
C24 VDD a_15757_1005 2.00fF
C25 VDD a_9009_1004 2.08fF
C26 a_5457_1004 a_5779_943 2.06fF
C27 a_599_943 VDD 2.34fF
C28 a_5457_1004 a_5327_159 3.62fF
C29 CLK a_10507_159 3.54fF
C30 a_10637_1004 a_9331_943 4.14fF
C31 RN GND 4.65fF
C32 VDD GND 42.64fF
C33 a_9331_943 GND 3.59fF **FLOATING
C34 a_4151_943 GND 3.64fF **FLOATING
.ends
