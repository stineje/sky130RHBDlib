magic
tech sky130A
magscale 1 2
timestamp 1669564307
<< nwell >>
rect -87 786 753 1550
<< pwell >>
rect -34 -34 700 544
<< nmos >>
rect 168 296 198 349
tri 198 296 214 312 sw
rect 362 296 392 349
tri 392 296 408 312 sw
rect 168 266 274 296
tri 274 266 304 296 sw
rect 168 165 198 266
tri 198 250 214 266 nw
tri 258 250 274 266 ne
tri 198 165 214 181 sw
tri 258 165 274 181 se
rect 274 165 304 266
rect 362 266 468 296
tri 468 266 498 296 sw
rect 362 251 393 266
tri 393 251 408 266 nw
tri 452 251 467 266 ne
rect 467 251 498 266
tri 168 135 198 165 ne
rect 198 135 274 165
tri 274 135 304 165 nw
rect 362 165 392 251
tri 392 165 408 181 sw
tri 452 165 468 181 se
rect 468 165 498 251
tri 362 135 392 165 ne
rect 392 135 468 165
tri 468 135 498 165 nw
<< pmos >>
rect 187 1005 217 1405
rect 275 1005 305 1405
rect 363 1005 393 1405
rect 451 1005 481 1405
<< ndiff >>
rect 112 333 168 349
rect 112 299 122 333
rect 156 299 168 333
rect 112 261 168 299
rect 198 312 362 349
tri 198 296 214 312 ne
rect 214 296 362 312
rect 392 312 554 349
tri 392 296 408 312 ne
rect 408 296 554 312
tri 274 266 304 296 ne
rect 112 227 122 261
rect 156 227 168 261
rect 112 193 168 227
rect 112 159 122 193
rect 156 159 168 193
tri 198 250 214 266 se
rect 214 250 258 266
tri 258 250 274 266 sw
rect 198 217 274 250
rect 198 183 219 217
rect 253 183 274 217
rect 198 181 274 183
tri 198 165 214 181 ne
rect 214 165 258 181
tri 258 165 274 181 nw
rect 304 261 362 296
tri 468 266 498 296 ne
rect 304 227 316 261
rect 350 227 362 261
tri 393 251 408 266 se
rect 408 251 452 266
tri 452 251 467 266 sw
rect 498 261 554 296
rect 304 193 362 227
rect 112 135 168 159
tri 168 135 198 165 sw
tri 274 135 304 165 se
rect 304 159 316 193
rect 350 159 362 193
rect 392 217 468 251
rect 392 183 413 217
rect 447 183 468 217
rect 392 181 468 183
tri 392 165 408 181 ne
rect 408 165 452 181
tri 452 165 468 181 nw
rect 498 227 510 261
rect 544 227 554 261
rect 498 193 554 227
rect 304 135 362 159
tri 362 135 392 165 sw
tri 468 135 498 165 se
rect 498 159 510 193
rect 544 159 554 193
rect 498 135 554 159
rect 112 123 554 135
rect 112 89 122 123
rect 156 89 219 123
rect 253 89 316 123
rect 350 89 413 123
rect 447 89 510 123
rect 544 89 554 123
rect 112 73 554 89
<< pdiff >>
rect 131 1365 187 1405
rect 131 1331 141 1365
rect 175 1331 187 1365
rect 131 1297 187 1331
rect 131 1263 141 1297
rect 175 1263 187 1297
rect 131 1229 187 1263
rect 131 1195 141 1229
rect 175 1195 187 1229
rect 131 1161 187 1195
rect 131 1127 141 1161
rect 175 1127 187 1161
rect 131 1093 187 1127
rect 131 1059 141 1093
rect 175 1059 187 1093
rect 131 1005 187 1059
rect 217 1365 275 1405
rect 217 1331 229 1365
rect 263 1331 275 1365
rect 217 1297 275 1331
rect 217 1263 229 1297
rect 263 1263 275 1297
rect 217 1229 275 1263
rect 217 1195 229 1229
rect 263 1195 275 1229
rect 217 1161 275 1195
rect 217 1127 229 1161
rect 263 1127 275 1161
rect 217 1005 275 1127
rect 305 1365 363 1405
rect 305 1331 317 1365
rect 351 1331 363 1365
rect 305 1297 363 1331
rect 305 1263 317 1297
rect 351 1263 363 1297
rect 305 1229 363 1263
rect 305 1195 317 1229
rect 351 1195 363 1229
rect 305 1161 363 1195
rect 305 1127 317 1161
rect 351 1127 363 1161
rect 305 1093 363 1127
rect 305 1059 317 1093
rect 351 1059 363 1093
rect 305 1005 363 1059
rect 393 1297 451 1405
rect 393 1263 405 1297
rect 439 1263 451 1297
rect 393 1229 451 1263
rect 393 1195 405 1229
rect 439 1195 451 1229
rect 393 1161 451 1195
rect 393 1127 405 1161
rect 439 1127 451 1161
rect 393 1093 451 1127
rect 393 1059 405 1093
rect 439 1059 451 1093
rect 393 1005 451 1059
rect 481 1365 535 1405
rect 481 1331 493 1365
rect 527 1331 535 1365
rect 481 1297 535 1331
rect 481 1263 493 1297
rect 527 1263 535 1297
rect 481 1229 535 1263
rect 481 1195 493 1229
rect 527 1195 535 1229
rect 481 1161 535 1195
rect 481 1127 493 1161
rect 527 1127 535 1161
rect 481 1005 535 1127
<< ndiffc >>
rect 122 299 156 333
rect 122 227 156 261
rect 122 159 156 193
rect 219 183 253 217
rect 316 227 350 261
rect 316 159 350 193
rect 413 183 447 217
rect 510 227 544 261
rect 510 159 544 193
rect 122 89 156 123
rect 219 89 253 123
rect 316 89 350 123
rect 413 89 447 123
rect 510 89 544 123
<< pdiffc >>
rect 141 1331 175 1365
rect 141 1263 175 1297
rect 141 1195 175 1229
rect 141 1127 175 1161
rect 141 1059 175 1093
rect 229 1331 263 1365
rect 229 1263 263 1297
rect 229 1195 263 1229
rect 229 1127 263 1161
rect 317 1331 351 1365
rect 317 1263 351 1297
rect 317 1195 351 1229
rect 317 1127 351 1161
rect 317 1059 351 1093
rect 405 1263 439 1297
rect 405 1195 439 1229
rect 405 1127 439 1161
rect 405 1059 439 1093
rect 493 1331 527 1365
rect 493 1263 527 1297
rect 493 1195 527 1229
rect 493 1127 527 1161
<< psubdiff >>
rect -34 482 700 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 632 461 700 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 632 427 649 461
rect 683 427 700 461
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 632 313 700 353
rect 632 279 649 313
rect 683 279 700 313
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect -34 17 34 57
rect 632 57 649 91
rect 683 57 700 91
rect 632 17 700 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 700 17
rect -34 -34 700 -17
<< nsubdiff >>
rect -34 1497 700 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 700 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 632 1423 700 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 632 979 700 1019
rect 632 945 649 979
rect 683 945 700 979
rect -34 871 -17 905
rect 17 884 34 905
rect 632 905 700 945
rect 632 884 649 905
rect 17 871 649 884
rect 683 871 700 905
rect -34 822 700 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 649 427 683 461
rect 649 353 683 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 649 279 683 313
rect 649 205 683 239
rect 649 131 683 165
rect 649 57 683 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 649 1389 683 1423
rect 649 1315 683 1349
rect 649 1241 683 1275
rect 649 1167 683 1201
rect 649 1093 683 1127
rect 649 1019 683 1053
rect -17 945 17 979
rect 649 945 683 979
rect -17 871 17 905
rect 649 871 683 905
<< poly >>
rect 187 1405 217 1431
rect 275 1405 305 1431
rect 363 1405 393 1431
rect 451 1405 481 1431
rect 187 974 217 1005
rect 275 974 305 1005
rect 363 974 393 1005
rect 451 974 481 1005
rect 164 958 305 974
rect 164 924 174 958
rect 208 944 305 958
rect 350 958 481 974
rect 208 924 218 944
rect 164 908 218 924
rect 350 924 360 958
rect 394 944 481 958
rect 394 924 404 944
rect 350 908 404 924
rect 195 433 249 449
rect 195 413 205 433
rect 168 399 205 413
rect 239 399 249 433
rect 168 383 249 399
rect 343 433 397 449
rect 343 399 353 433
rect 387 399 397 433
rect 343 383 397 399
rect 168 349 198 383
rect 362 349 392 383
<< polycont >>
rect 174 924 208 958
rect 360 924 394 958
rect 205 399 239 433
rect 353 399 387 433
<< locali >>
rect -34 1497 700 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 700 1497
rect -34 1446 700 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 141 1365 175 1405
rect 141 1297 175 1331
rect 141 1229 175 1263
rect 141 1161 175 1195
rect 141 1093 175 1127
rect 229 1365 263 1446
rect 632 1423 700 1446
rect 229 1297 263 1331
rect 229 1229 263 1263
rect 229 1161 263 1195
rect 229 1111 263 1127
rect 317 1365 527 1399
rect 317 1297 351 1331
rect 317 1229 351 1263
rect 317 1161 351 1195
rect 317 1093 351 1127
rect 141 1025 351 1059
rect 405 1297 439 1313
rect 405 1229 439 1263
rect 405 1161 439 1195
rect 405 1093 439 1127
rect 493 1297 527 1331
rect 493 1229 527 1263
rect 493 1161 527 1195
rect 493 1111 527 1127
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 405 1025 535 1059
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 174 958 208 974
rect 360 958 394 974
rect 208 924 239 942
rect 174 908 239 924
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 908
rect 205 383 239 399
rect 353 924 360 942
rect 353 908 394 924
rect 353 433 387 908
rect 353 383 387 399
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 122 333 156 349
rect 501 348 535 1025
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect 632 979 700 1019
rect 632 945 649 979
rect 683 945 700 979
rect 632 905 700 945
rect 632 871 649 905
rect 683 871 700 905
rect 632 822 700 871
rect 122 261 156 299
rect 122 193 156 227
rect 219 314 535 348
rect 632 461 700 544
rect 632 427 649 461
rect 683 427 700 461
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect 219 217 253 314
rect 219 167 253 183
rect 316 261 350 278
rect 316 193 350 227
rect 122 123 156 159
rect 413 217 447 314
rect 632 313 700 353
rect 632 279 649 313
rect 683 279 700 313
rect 413 167 447 183
rect 510 261 544 278
rect 510 193 544 227
rect 316 123 350 159
rect 510 123 544 159
rect 156 89 219 123
rect 253 89 316 123
rect 350 89 413 123
rect 447 89 510 123
rect 122 34 156 89
rect 219 34 253 89
rect 316 34 350 89
rect 413 34 447 89
rect 510 34 544 89
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect 632 57 649 91
rect 683 57 700 91
rect 632 34 700 57
rect -34 17 700 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 700 17
rect -34 -34 700 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
<< metal1 >>
rect -34 1497 700 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 700 1497
rect -34 1446 700 1463
rect -34 17 700 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 700 17
rect -34 -34 700 -17
<< labels >>
rlabel metal1 501 427 535 461 1 Y
port 1 n
rlabel metal1 501 501 535 535 1 Y
port 2 n
rlabel metal1 501 575 535 609 1 Y
port 3 n
rlabel metal1 501 649 535 683 1 Y
port 4 n
rlabel metal1 501 723 535 757 1 Y
port 5 n
rlabel metal1 501 797 535 831 1 Y
port 6 n
rlabel metal1 501 871 535 905 1 Y
port 7 n
rlabel metal1 205 427 239 461 1 A
port 8 n
rlabel metal1 205 501 239 535 1 A
port 9 n
rlabel metal1 205 575 239 609 1 A
port 10 n
rlabel metal1 205 649 239 683 1 A
port 11 n
rlabel metal1 205 723 239 757 1 A
port 12 n
rlabel metal1 205 797 239 831 1 A
port 13 n
rlabel metal1 205 871 239 905 1 A
port 14 n
rlabel metal1 353 427 387 461 1 B
port 15 n
rlabel metal1 353 501 387 535 1 B
port 16 n
rlabel metal1 353 575 387 609 1 B
port 17 n
rlabel metal1 353 649 387 683 1 B
port 18 n
rlabel metal1 353 723 387 757 1 B
port 19 n
rlabel metal1 353 797 387 831 1 B
port 20 n
rlabel metal1 353 871 387 905 1 B
port 21 n
rlabel metal1 -34 1446 700 1514 1 VPWR
port 22 n
rlabel metal1 -34 -34 700 34 1 VGND
port 23 n
rlabel nwell 57 1463 91 1497 1 VPB
port 24 n
rlabel pwell 57 -17 91 17 1 VNB
port 25 n
<< end >>
