* SPICE3 file created from TMRDFFRNQX1.ext - technology: sky130A

.subckt TMRDFFRNQX1 Q D CLK RN VPB VNB
M1000 a_14511_943.t4 a_10507_159.t14 VPB.t47 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_9331_943.t7 a_9331_943.t6 VPB.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VNB a_9009_1004.t9 a_9806_73.t0 nshort w=-1.605u l=1.765u
+  ad=4.9019p pd=41.07u as=0p ps=0u
M1003 VPB.t85 RN a_9331_943.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VNB a_5779_943.t12 a_7216_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1005 VNB a_10507_159.t21 a_10451_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_5457_1004.t5 a_5779_943.t7 VPB.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_5327_159.t4 RN VPB.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t101 a_147_159.t14 a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_15757_1005.t7 a_4151_943.t5 a_16421_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t49 a_10507_159.t15 a_10637_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPB.t0 a_9331_943.t19 a_10507_159.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t90 RN a_10507_159.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_10507_159.t1 a_10637_1004.t7 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_9331_943.t14 a_10637_1004.t8 VPB.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_599_943.t1 D VPB.t41 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_16421_1005.t0 a_14511_943.t6 a_15932_181.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_5327_159.t2 CLK VPB.t63 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPB.t33 a_599_943.t7 a_2141_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_9331_943.t1 a_9009_1004.t7 VPB.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPB.t57 CLK a_277_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPB.t28 a_5457_1004.t7 a_9009_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t30 a_277_1004.t8 a_147_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPB.t4 a_5457_1004.t8 a_5779_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPB.t93 RN a_5779_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPB.t79 a_9331_943.t21 a_9009_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPB.t56 CLK a_10637_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPB.t61 CLK a_10507_159.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_9331_943.t15 a_5327_159.t8 VPB.t78 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VNB a_5457_1004.t11 a_8823_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_10507_159.t12 RN VPB.t89 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_9331_943.t3 D VPB.t36 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_599_943.t5 RN VPB.t96 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_147_159.t8 a_4151_943.t7 VPB.t68 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VNB a_5457_1004.t12 a_6233_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPB.t2 a_14511_943.t7 a_15757_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_10637_1004.t3 a_10507_159.t16 VPB.t50 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_147_159.t7 CLK VPB.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_4151_943.t3 a_147_159.t16 VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_9009_1004.t3 a_5457_1004.t9 VPB.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_15757_1005.t3 a_9331_943.t23 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPB.t52 a_10507_159.t17 a_14511_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPB.t5 a_9331_943.t4 a_9331_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 VNB a_147_159.t15 a_4626_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPB.t7 a_147_159.t17 a_2141_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPB.t74 a_599_943.t9 a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 VNB a_147_159.t24 a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPB.t38 D a_5779_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 VPB.t97 RN a_9009_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 VNB a_599_943.t8 a_2036_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1050 VNB a_7321_1004.t7 a_7861_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1051 VPB.t77 a_5327_159.t10 a_5457_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 VPB.t43 a_7321_1004.t5 a_5327_159.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 VPB.t42 a_2141_1004.t6 a_147_159.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_10507_159.t4 a_14511_943.t8 VPB.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 VNB a_5327_159.t14 a_5271_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_9331_943.t16 RN VPB.t83 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_147_159.t12 RN VPB.t82 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_4151_943.t2 a_147_159.t18 VPB.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 a_7321_1004.t1 a_5327_159.t11 VPB.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 a_15932_181.t6 a_4151_943.t8 a_16421_1005.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 VPB.t10 a_9331_943.t26 a_10637_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 VNB a_9331_943.t24 a_15652_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1063 VNB a_10507_159.t18 a_14986_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_15757_1005.t0 a_14511_943.t9 VPB.t54 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 VPB.t51 a_10507_159.t19 a_14511_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 VPB.t53 a_10507_159.t20 a_9331_943.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1067 VPB.t100 a_15932_181.t8 a_17723_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_277_1004.t5 a_147_159.t19 VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 VPB.t67 a_9009_1004.t8 a_9331_943.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_16421_1005.t4 a_4151_943.t10 a_15757_1005.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 VNB a_9331_943.t20 a_13041_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_10507_159.t2 a_9331_943.t27 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 a_10637_1004.t1 a_9331_943.t28 VPB.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 a_10507_159.t11 RN VPB.t88 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 VNB a_277_1004.t7 a_3643_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1076 a_7321_1004.t4 a_5779_943.t8 VPB.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 VPB.t32 a_277_1004.t10 a_599_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 a_15932_181.t2 a_14511_943.t10 a_16421_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VPB.t94 RN a_599_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 VPB.t26 a_4151_943.t11 a_147_159.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 VNB a_4151_943.t9 a_16984_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1082 VPB.t70 a_5779_943.t9 a_5457_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 VPB.t95 RN a_5327_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_16421_1005.t3 a_9331_943.t30 a_15757_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_2141_1004.t0 a_599_943.t10 VPB.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_277_1004.t2 CLK VPB.t59 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 a_147_159.t2 a_277_1004.t11 VPB.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_5779_943.t1 a_5457_1004.t10 VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_10637_1004.t5 CLK VPB.t55 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 a_10507_159.t6 CLK VPB.t60 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 VNB a_10637_1004.t9 a_14003_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1092 VNB a_2141_1004.t5 a_2681_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_17723_182.t0 a_15932_181.t9 VPB.t99 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 VPB.t76 a_10637_1004.t11 a_10507_159.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 VPB.t71 a_10637_1004.t12 a_9331_943.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 VPB.t39 D a_599_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 VPB.t92 RN a_147_159.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 VNB a_9331_943.t29 a_12396_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1099 a_599_943.t2 a_277_1004.t12 VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 VPB.t66 CLK a_5457_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 VPB.t64 CLK a_5327_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_2141_1004.t2 a_147_159.t22 VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_277_1004.t0 a_599_943.t11 VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_147_159.t10 RN VPB.t81 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 a_5779_943.t2 D VPB.t37 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 a_9009_1004.t5 RN VPB.t86 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 a_5327_159.t6 a_7321_1004.t6 VPB.t98 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 VPB.t21 a_5327_159.t12 a_9331_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 a_147_159.t5 a_2141_1004.t7 VPB.t44 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_5457_1004.t0 a_5327_159.t13 VPB.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 VPB.t87 RN a_10507_159.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1112 VPB.t40 D a_9331_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 VNB a_277_1004.t9 a_1053_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1114 VPB.t58 CLK a_147_159.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 VPB.t69 a_5779_943.t10 a_7321_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 VPB.t13 a_147_159.t23 a_4151_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1117 VPB.t24 a_9331_943.t32 a_15757_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_14511_943.t1 a_10507_159.t23 VPB.t46 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_9331_943.t8 a_10507_159.t24 VPB.t48 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 VNB a_9331_943.t31 a_16318_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1121 a_9009_1004.t0 a_9331_943.t33 VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 a_5779_943.t4 RN VPB.t91 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 VNB a_10637_1004.t10 a_11413_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1124 a_5457_1004.t2 CLK VPB.t65 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1125 a_15757_1005.t4 a_9331_943.t34 a_16421_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1126 VPB.t27 a_14511_943.t13 a_10507_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1127 VPB.t80 RN a_147_159.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1128 VPB.t15 a_147_159.t25 a_4151_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1129 VPB.t72 a_5327_159.t15 a_7321_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1130 a_16421_1005.t5 a_4151_943.t13 a_15932_181.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB RN 0.50fF
C1 D CLK 1.65fF
C2 D RN 12.41fF
C3 CLK RN 1.02fF
C4 VPB D 0.15fF
C5 VPB CLK 3.49fF
R0 a_10507_159.n23 a_10507_159.t15 512.525
R1 a_10507_159.n8 a_10507_159.t17 480.392
R2 a_10507_159.n21 a_10507_159.t20 472.359
R3 a_10507_159.n6 a_10507_159.t19 472.359
R4 a_10507_159.n8 a_10507_159.t14 403.272
R5 a_10507_159.n21 a_10507_159.t24 384.527
R6 a_10507_159.n6 a_10507_159.t23 384.527
R7 a_10507_159.n23 a_10507_159.t16 371.139
R8 a_10507_159.n24 a_10507_159.t21 324.268
R9 a_10507_159.n9 a_10507_159.t18 320.08
R10 a_10507_159.n22 a_10507_159.t25 277.772
R11 a_10507_159.n7 a_10507_159.t22 277.772
R12 a_10507_159.n20 a_10507_159.n19 249.704
R13 a_10507_159.n30 a_10507_159.n28 249.704
R14 a_10507_159.n20 a_10507_159.n15 127.74
R15 a_10507_159.n28 a_10507_159.n5 127.74
R16 a_10507_159.n24 a_10507_159.n23 119.654
R17 a_10507_159.n25 a_10507_159.n24 83.572
R18 a_10507_159.n4 a_10507_159.n3 79.232
R19 a_10507_159.n14 a_10507_159.n13 79.232
R20 a_10507_159.n10 a_10507_159.n7 76.499
R21 a_10507_159.n25 a_10507_159.n22 76
R22 a_10507_159.n26 a_10507_159.n20 76
R23 a_10507_159.n10 a_10507_159.n9 76
R24 a_10507_159.n28 a_10507_159.n27 76
R25 a_10507_159.n22 a_10507_159.n21 67.001
R26 a_10507_159.n7 a_10507_159.n6 67.001
R27 a_10507_159.n15 a_10507_159.n14 63.152
R28 a_10507_159.n5 a_10507_159.n4 63.152
R29 a_10507_159.n9 a_10507_159.n8 55.388
R30 a_10507_159.n31 a_10507_159.n0 55.263
R31 a_10507_159.n19 a_10507_159.n18 30
R32 a_10507_159.n30 a_10507_159.n29 30
R33 a_10507_159.n17 a_10507_159.n16 24.383
R34 a_10507_159.n19 a_10507_159.n17 23.684
R35 a_10507_159.n31 a_10507_159.n30 23.684
R36 a_10507_159.n15 a_10507_159.n11 16.08
R37 a_10507_159.n14 a_10507_159.n12 16.08
R38 a_10507_159.n5 a_10507_159.n1 16.08
R39 a_10507_159.n4 a_10507_159.n2 16.08
R40 a_10507_159.n11 a_10507_159.t13 14.282
R41 a_10507_159.n11 a_10507_159.t11 14.282
R42 a_10507_159.n12 a_10507_159.t7 14.282
R43 a_10507_159.n12 a_10507_159.t6 14.282
R44 a_10507_159.n13 a_10507_159.t0 14.282
R45 a_10507_159.n13 a_10507_159.t2 14.282
R46 a_10507_159.n1 a_10507_159.t3 14.282
R47 a_10507_159.n1 a_10507_159.t4 14.282
R48 a_10507_159.n2 a_10507_159.t10 14.282
R49 a_10507_159.n2 a_10507_159.t12 14.282
R50 a_10507_159.n3 a_10507_159.t8 14.282
R51 a_10507_159.n3 a_10507_159.t1 14.282
R52 a_10507_159.n26 a_10507_159.n25 4.035
R53 a_10507_159.n27 a_10507_159.n26 3.491
R54 a_10507_159.n27 a_10507_159.n10 1.315
R55 VPB VPB.n1609 126.832
R56 VPB.n40 VPB.n38 94.117
R57 VPB.n1531 VPB.n1529 94.117
R58 VPB.n1468 VPB.n1466 94.117
R59 VPB.n1385 VPB.n1383 94.117
R60 VPB.n1302 VPB.n1300 94.117
R61 VPB.n1239 VPB.n1237 94.117
R62 VPB.n1156 VPB.n1154 94.117
R63 VPB.n1073 VPB.n1071 94.117
R64 VPB.n1010 VPB.n1008 94.117
R65 VPB.n927 VPB.n925 94.117
R66 VPB.n115 VPB.n113 94.117
R67 VPB.n845 VPB.n843 94.117
R68 VPB.n762 VPB.n760 94.117
R69 VPB.n679 VPB.n677 94.117
R70 VPB.n616 VPB.n614 94.117
R71 VPB.n533 VPB.n531 94.117
R72 VPB.n450 VPB.n448 94.117
R73 VPB.n387 VPB.n385 94.117
R74 VPB.n324 VPB.n322 94.117
R75 VPB.n269 VPB.n267 94.117
R76 VPB.n214 VPB.n212 91.036
R77 VPB.n463 VPB.n462 80.104
R78 VPB.n546 VPB.n545 80.104
R79 VPB.n692 VPB.n691 80.104
R80 VPB.n775 VPB.n774 80.104
R81 VPB.n125 VPB.n124 80.104
R82 VPB.n940 VPB.n939 80.104
R83 VPB.n1086 VPB.n1085 80.104
R84 VPB.n1169 VPB.n1168 80.104
R85 VPB.n1315 VPB.n1314 80.104
R86 VPB.n1398 VPB.n1397 80.104
R87 VPB.n1544 VPB.n1543 80.104
R88 VPB.n50 VPB.n49 80.104
R89 VPB.n175 VPB.n169 76.136
R90 VPB.n175 VPB.n174 76
R91 VPB.n179 VPB.n178 76
R92 VPB.n185 VPB.n184 76
R93 VPB.n189 VPB.n188 76
R94 VPB.n216 VPB.n215 76
R95 VPB.n220 VPB.n219 76
R96 VPB.n224 VPB.n223 76
R97 VPB.n228 VPB.n227 76
R98 VPB.n232 VPB.n231 76
R99 VPB.n236 VPB.n235 76
R100 VPB.n240 VPB.n239 76
R101 VPB.n244 VPB.n243 76
R102 VPB.n271 VPB.n270 76
R103 VPB.n275 VPB.n274 76
R104 VPB.n279 VPB.n278 76
R105 VPB.n283 VPB.n282 76
R106 VPB.n287 VPB.n286 76
R107 VPB.n291 VPB.n290 76
R108 VPB.n295 VPB.n294 76
R109 VPB.n299 VPB.n298 76
R110 VPB.n326 VPB.n325 76
R111 VPB.n331 VPB.n330 76
R112 VPB.n336 VPB.n335 76
R113 VPB.n343 VPB.n342 76
R114 VPB.n348 VPB.n347 76
R115 VPB.n353 VPB.n352 76
R116 VPB.n358 VPB.n357 76
R117 VPB.n362 VPB.n361 76
R118 VPB.n389 VPB.n388 76
R119 VPB.n394 VPB.n393 76
R120 VPB.n399 VPB.n398 76
R121 VPB.n406 VPB.n405 76
R122 VPB.n411 VPB.n410 76
R123 VPB.n416 VPB.n415 76
R124 VPB.n421 VPB.n420 76
R125 VPB.n425 VPB.n424 76
R126 VPB.n452 VPB.n451 76
R127 VPB.n456 VPB.n455 76
R128 VPB.n461 VPB.n460 76
R129 VPB.n466 VPB.n465 76
R130 VPB.n473 VPB.n472 76
R131 VPB.n478 VPB.n477 76
R132 VPB.n483 VPB.n482 76
R133 VPB.n490 VPB.n489 76
R134 VPB.n495 VPB.n494 76
R135 VPB.n500 VPB.n499 76
R136 VPB.n504 VPB.n503 76
R137 VPB.n508 VPB.n507 76
R138 VPB.n535 VPB.n534 76
R139 VPB.n539 VPB.n538 76
R140 VPB.n544 VPB.n543 76
R141 VPB.n549 VPB.n548 76
R142 VPB.n556 VPB.n555 76
R143 VPB.n561 VPB.n560 76
R144 VPB.n566 VPB.n565 76
R145 VPB.n573 VPB.n572 76
R146 VPB.n578 VPB.n577 76
R147 VPB.n583 VPB.n582 76
R148 VPB.n587 VPB.n586 76
R149 VPB.n591 VPB.n590 76
R150 VPB.n618 VPB.n617 76
R151 VPB.n623 VPB.n622 76
R152 VPB.n628 VPB.n627 76
R153 VPB.n635 VPB.n634 76
R154 VPB.n640 VPB.n639 76
R155 VPB.n645 VPB.n644 76
R156 VPB.n650 VPB.n649 76
R157 VPB.n654 VPB.n653 76
R158 VPB.n681 VPB.n680 76
R159 VPB.n685 VPB.n684 76
R160 VPB.n690 VPB.n689 76
R161 VPB.n695 VPB.n694 76
R162 VPB.n702 VPB.n701 76
R163 VPB.n707 VPB.n706 76
R164 VPB.n712 VPB.n711 76
R165 VPB.n719 VPB.n718 76
R166 VPB.n724 VPB.n723 76
R167 VPB.n729 VPB.n728 76
R168 VPB.n733 VPB.n732 76
R169 VPB.n737 VPB.n736 76
R170 VPB.n764 VPB.n763 76
R171 VPB.n768 VPB.n767 76
R172 VPB.n773 VPB.n772 76
R173 VPB.n778 VPB.n777 76
R174 VPB.n785 VPB.n784 76
R175 VPB.n790 VPB.n789 76
R176 VPB.n795 VPB.n794 76
R177 VPB.n802 VPB.n801 76
R178 VPB.n807 VPB.n806 76
R179 VPB.n812 VPB.n811 76
R180 VPB.n816 VPB.n815 76
R181 VPB.n820 VPB.n819 76
R182 VPB.n847 VPB.n846 76
R183 VPB.n852 VPB.n851 76
R184 VPB.n857 VPB.n856 76
R185 VPB.n864 VPB.n863 76
R186 VPB.n869 VPB.n868 76
R187 VPB.n874 VPB.n873 76
R188 VPB.n889 VPB.n885 76
R189 VPB.n894 VPB.n893 76
R190 VPB.n898 VPB.n897 76
R191 VPB.n902 VPB.n901 76
R192 VPB.n929 VPB.n928 76
R193 VPB.n933 VPB.n932 76
R194 VPB.n938 VPB.n937 76
R195 VPB.n943 VPB.n942 76
R196 VPB.n950 VPB.n949 76
R197 VPB.n955 VPB.n954 76
R198 VPB.n960 VPB.n959 76
R199 VPB.n967 VPB.n966 76
R200 VPB.n972 VPB.n971 76
R201 VPB.n977 VPB.n976 76
R202 VPB.n981 VPB.n980 76
R203 VPB.n985 VPB.n984 76
R204 VPB.n1012 VPB.n1011 76
R205 VPB.n1017 VPB.n1016 76
R206 VPB.n1022 VPB.n1021 76
R207 VPB.n1029 VPB.n1028 76
R208 VPB.n1034 VPB.n1033 76
R209 VPB.n1039 VPB.n1038 76
R210 VPB.n1044 VPB.n1043 76
R211 VPB.n1048 VPB.n1047 76
R212 VPB.n1075 VPB.n1074 76
R213 VPB.n1079 VPB.n1078 76
R214 VPB.n1084 VPB.n1083 76
R215 VPB.n1089 VPB.n1088 76
R216 VPB.n1096 VPB.n1095 76
R217 VPB.n1101 VPB.n1100 76
R218 VPB.n1106 VPB.n1105 76
R219 VPB.n1113 VPB.n1112 76
R220 VPB.n1118 VPB.n1117 76
R221 VPB.n1123 VPB.n1122 76
R222 VPB.n1127 VPB.n1126 76
R223 VPB.n1131 VPB.n1130 76
R224 VPB.n1158 VPB.n1157 76
R225 VPB.n1162 VPB.n1161 76
R226 VPB.n1167 VPB.n1166 76
R227 VPB.n1172 VPB.n1171 76
R228 VPB.n1179 VPB.n1178 76
R229 VPB.n1184 VPB.n1183 76
R230 VPB.n1189 VPB.n1188 76
R231 VPB.n1196 VPB.n1195 76
R232 VPB.n1201 VPB.n1200 76
R233 VPB.n1206 VPB.n1205 76
R234 VPB.n1210 VPB.n1209 76
R235 VPB.n1214 VPB.n1213 76
R236 VPB.n1241 VPB.n1240 76
R237 VPB.n1246 VPB.n1245 76
R238 VPB.n1251 VPB.n1250 76
R239 VPB.n1258 VPB.n1257 76
R240 VPB.n1263 VPB.n1262 76
R241 VPB.n1268 VPB.n1267 76
R242 VPB.n1273 VPB.n1272 76
R243 VPB.n1277 VPB.n1276 76
R244 VPB.n1304 VPB.n1303 76
R245 VPB.n1308 VPB.n1307 76
R246 VPB.n1313 VPB.n1312 76
R247 VPB.n1318 VPB.n1317 76
R248 VPB.n1325 VPB.n1324 76
R249 VPB.n1330 VPB.n1329 76
R250 VPB.n1335 VPB.n1334 76
R251 VPB.n1342 VPB.n1341 76
R252 VPB.n1347 VPB.n1346 76
R253 VPB.n1352 VPB.n1351 76
R254 VPB.n1356 VPB.n1355 76
R255 VPB.n1360 VPB.n1359 76
R256 VPB.n1387 VPB.n1386 76
R257 VPB.n1391 VPB.n1390 76
R258 VPB.n1396 VPB.n1395 76
R259 VPB.n1401 VPB.n1400 76
R260 VPB.n1408 VPB.n1407 76
R261 VPB.n1413 VPB.n1412 76
R262 VPB.n1418 VPB.n1417 76
R263 VPB.n1425 VPB.n1424 76
R264 VPB.n1430 VPB.n1429 76
R265 VPB.n1435 VPB.n1434 76
R266 VPB.n1439 VPB.n1438 76
R267 VPB.n1443 VPB.n1442 76
R268 VPB.n1470 VPB.n1469 76
R269 VPB.n1475 VPB.n1474 76
R270 VPB.n1480 VPB.n1479 76
R271 VPB.n1487 VPB.n1486 76
R272 VPB.n1492 VPB.n1491 76
R273 VPB.n1497 VPB.n1496 76
R274 VPB.n1502 VPB.n1501 76
R275 VPB.n1506 VPB.n1505 76
R276 VPB.n1533 VPB.n1532 76
R277 VPB.n1537 VPB.n1536 76
R278 VPB.n1542 VPB.n1541 76
R279 VPB.n1547 VPB.n1546 76
R280 VPB.n1554 VPB.n1553 76
R281 VPB.n1559 VPB.n1558 76
R282 VPB.n1564 VPB.n1563 76
R283 VPB.n1571 VPB.n1570 76
R284 VPB.n1576 VPB.n1575 76
R285 VPB.n1581 VPB.n1580 76
R286 VPB.n1585 VPB.n1584 76
R287 VPB.n1589 VPB.n1588 76
R288 VPB.n1602 VPB.n1601 76
R289 VPB.n492 VPB.n491 75.654
R290 VPB.n575 VPB.n574 75.654
R291 VPB.n721 VPB.n720 75.654
R292 VPB.n804 VPB.n803 75.654
R293 VPB.n887 VPB.n886 75.654
R294 VPB.n969 VPB.n968 75.654
R295 VPB.n1115 VPB.n1114 75.654
R296 VPB.n1198 VPB.n1197 75.654
R297 VPB.n1344 VPB.n1343 75.654
R298 VPB.n1427 VPB.n1426 75.654
R299 VPB.n1573 VPB.n1572 75.654
R300 VPB.n72 VPB.n71 75.654
R301 VPB.n182 VPB.n181 68.979
R302 VPB.n172 VPB.n171 64.528
R303 VPB.n22 VPB.n21 61.764
R304 VPB.n1513 VPB.n1512 61.764
R305 VPB.n1450 VPB.n1449 61.764
R306 VPB.n1367 VPB.n1366 61.764
R307 VPB.n1284 VPB.n1283 61.764
R308 VPB.n1221 VPB.n1220 61.764
R309 VPB.n1138 VPB.n1137 61.764
R310 VPB.n1055 VPB.n1054 61.764
R311 VPB.n992 VPB.n991 61.764
R312 VPB.n909 VPB.n908 61.764
R313 VPB.n90 VPB.n89 61.764
R314 VPB.n827 VPB.n826 61.764
R315 VPB.n744 VPB.n743 61.764
R316 VPB.n661 VPB.n660 61.764
R317 VPB.n598 VPB.n597 61.764
R318 VPB.n515 VPB.n514 61.764
R319 VPB.n432 VPB.n431 61.764
R320 VPB.n369 VPB.n368 61.764
R321 VPB.n306 VPB.n305 61.764
R322 VPB.n251 VPB.n250 61.764
R323 VPB.n196 VPB.n195 61.764
R324 VPB.n354 VPB.t1 55.465
R325 VPB.n327 VPB.t2 55.465
R326 VPB.n78 VPB.t9 55.106
R327 VPB.n1577 VPB.t3 55.106
R328 VPB.n1498 VPB.t29 55.106
R329 VPB.n1431 VPB.t44 55.106
R330 VPB.n1348 VPB.t31 55.106
R331 VPB.n1269 VPB.t14 55.106
R332 VPB.n1202 VPB.t73 55.106
R333 VPB.n1119 VPB.t20 55.106
R334 VPB.n1040 VPB.t19 55.106
R335 VPB.n973 VPB.t98 55.106
R336 VPB.n890 VPB.t16 55.106
R337 VPB.n105 VPB.t34 55.106
R338 VPB.n808 VPB.t50 55.106
R339 VPB.n725 VPB.t75 55.106
R340 VPB.n646 VPB.t22 55.106
R341 VPB.n579 VPB.t12 55.106
R342 VPB.n496 VPB.t6 55.106
R343 VPB.n417 VPB.t47 55.106
R344 VPB.n180 VPB.t99 55.106
R345 VPB.n170 VPB.t100 55.106
R346 VPB.n45 VPB.t74 55.106
R347 VPB.n1538 VPB.t94 55.106
R348 VPB.n1471 VPB.t7 55.106
R349 VPB.n1392 VPB.t80 55.106
R350 VPB.n1309 VPB.t26 55.106
R351 VPB.n1242 VPB.t15 55.106
R352 VPB.n1163 VPB.t70 55.106
R353 VPB.n1080 VPB.t93 55.106
R354 VPB.n1013 VPB.t72 55.106
R355 VPB.n934 VPB.t95 55.106
R356 VPB.n120 VPB.t79 55.106
R357 VPB.n848 VPB.t21 55.106
R358 VPB.n769 VPB.t10 55.106
R359 VPB.n686 VPB.t85 55.106
R360 VPB.n619 VPB.t53 55.106
R361 VPB.n540 VPB.t90 55.106
R362 VPB.n457 VPB.t27 55.106
R363 VPB.n390 VPB.t51 55.106
R364 VPB.n333 VPB.n332 48.952
R365 VPB.n396 VPB.n395 48.952
R366 VPB.n470 VPB.n469 48.952
R367 VPB.n553 VPB.n552 48.952
R368 VPB.n625 VPB.n624 48.952
R369 VPB.n699 VPB.n698 48.952
R370 VPB.n782 VPB.n781 48.952
R371 VPB.n854 VPB.n853 48.952
R372 VPB.n129 VPB.n128 48.952
R373 VPB.n947 VPB.n946 48.952
R374 VPB.n1019 VPB.n1018 48.952
R375 VPB.n1093 VPB.n1092 48.952
R376 VPB.n1176 VPB.n1175 48.952
R377 VPB.n1248 VPB.n1247 48.952
R378 VPB.n1322 VPB.n1321 48.952
R379 VPB.n1405 VPB.n1404 48.952
R380 VPB.n1477 VPB.n1476 48.952
R381 VPB.n1551 VPB.n1550 48.952
R382 VPB.n54 VPB.n53 48.952
R383 VPB.n350 VPB.n349 44.502
R384 VPB.n413 VPB.n412 44.502
R385 VPB.n487 VPB.n486 44.502
R386 VPB.n570 VPB.n569 44.502
R387 VPB.n642 VPB.n641 44.502
R388 VPB.n716 VPB.n715 44.502
R389 VPB.n799 VPB.n798 44.502
R390 VPB.n871 VPB.n870 44.502
R391 VPB.n143 VPB.n142 44.502
R392 VPB.n964 VPB.n963 44.502
R393 VPB.n1036 VPB.n1035 44.502
R394 VPB.n1110 VPB.n1109 44.502
R395 VPB.n1193 VPB.n1192 44.502
R396 VPB.n1265 VPB.n1264 44.502
R397 VPB.n1339 VPB.n1338 44.502
R398 VPB.n1422 VPB.n1421 44.502
R399 VPB.n1494 VPB.n1493 44.502
R400 VPB.n1568 VPB.n1567 44.502
R401 VPB.n68 VPB.n67 44.502
R402 VPB.n338 VPB.n337 41.183
R403 VPB.n66 VPB.n14 40.824
R404 VPB.n57 VPB.n15 40.824
R405 VPB.n1566 VPB.n1565 40.824
R406 VPB.n1549 VPB.n1548 40.824
R407 VPB.n1482 VPB.n1481 40.824
R408 VPB.n1420 VPB.n1419 40.824
R409 VPB.n1403 VPB.n1402 40.824
R410 VPB.n1337 VPB.n1336 40.824
R411 VPB.n1320 VPB.n1319 40.824
R412 VPB.n1253 VPB.n1252 40.824
R413 VPB.n1191 VPB.n1190 40.824
R414 VPB.n1174 VPB.n1173 40.824
R415 VPB.n1108 VPB.n1107 40.824
R416 VPB.n1091 VPB.n1090 40.824
R417 VPB.n1024 VPB.n1023 40.824
R418 VPB.n962 VPB.n961 40.824
R419 VPB.n945 VPB.n944 40.824
R420 VPB.n141 VPB.n82 40.824
R421 VPB.n132 VPB.n83 40.824
R422 VPB.n859 VPB.n858 40.824
R423 VPB.n797 VPB.n796 40.824
R424 VPB.n780 VPB.n779 40.824
R425 VPB.n714 VPB.n713 40.824
R426 VPB.n697 VPB.n696 40.824
R427 VPB.n630 VPB.n629 40.824
R428 VPB.n568 VPB.n567 40.824
R429 VPB.n551 VPB.n550 40.824
R430 VPB.n485 VPB.n484 40.824
R431 VPB.n468 VPB.n467 40.824
R432 VPB.n401 VPB.n400 40.824
R433 VPB.n1606 VPB.n1602 20.452
R434 VPB.n169 VPB.n166 20.452
R435 VPB.n340 VPB.n339 17.801
R436 VPB.n403 VPB.n402 17.801
R437 VPB.n475 VPB.n474 17.801
R438 VPB.n558 VPB.n557 17.801
R439 VPB.n632 VPB.n631 17.801
R440 VPB.n704 VPB.n703 17.801
R441 VPB.n787 VPB.n786 17.801
R442 VPB.n861 VPB.n860 17.801
R443 VPB.n134 VPB.n133 17.801
R444 VPB.n952 VPB.n951 17.801
R445 VPB.n1026 VPB.n1025 17.801
R446 VPB.n1098 VPB.n1097 17.801
R447 VPB.n1181 VPB.n1180 17.801
R448 VPB.n1255 VPB.n1254 17.801
R449 VPB.n1327 VPB.n1326 17.801
R450 VPB.n1410 VPB.n1409 17.801
R451 VPB.n1484 VPB.n1483 17.801
R452 VPB.n1556 VPB.n1555 17.801
R453 VPB.n59 VPB.n58 17.801
R454 VPB.n14 VPB.t59 14.282
R455 VPB.n14 VPB.t101 14.282
R456 VPB.n15 VPB.t17 14.282
R457 VPB.n15 VPB.t57 14.282
R458 VPB.n1565 VPB.t41 14.282
R459 VPB.n1565 VPB.t32 14.282
R460 VPB.n1548 VPB.t96 14.282
R461 VPB.n1548 VPB.t39 14.282
R462 VPB.n1481 VPB.t11 14.282
R463 VPB.n1481 VPB.t33 14.282
R464 VPB.n1419 VPB.t62 14.282
R465 VPB.n1419 VPB.t42 14.282
R466 VPB.n1402 VPB.t82 14.282
R467 VPB.n1402 VPB.t58 14.282
R468 VPB.n1336 VPB.t81 14.282
R469 VPB.n1336 VPB.t30 14.282
R470 VPB.n1319 VPB.t68 14.282
R471 VPB.n1319 VPB.t92 14.282
R472 VPB.n1252 VPB.t8 14.282
R473 VPB.n1252 VPB.t13 14.282
R474 VPB.n1190 VPB.t65 14.282
R475 VPB.n1190 VPB.t77 14.282
R476 VPB.n1173 VPB.t25 14.282
R477 VPB.n1173 VPB.t66 14.282
R478 VPB.n1107 VPB.t37 14.282
R479 VPB.n1107 VPB.t4 14.282
R480 VPB.n1090 VPB.t91 14.282
R481 VPB.n1090 VPB.t38 14.282
R482 VPB.n1023 VPB.t23 14.282
R483 VPB.n1023 VPB.t69 14.282
R484 VPB.n961 VPB.t63 14.282
R485 VPB.n961 VPB.t43 14.282
R486 VPB.n944 VPB.t84 14.282
R487 VPB.n944 VPB.t64 14.282
R488 VPB.n82 VPB.t86 14.282
R489 VPB.n82 VPB.t28 14.282
R490 VPB.n83 VPB.t18 14.282
R491 VPB.n83 VPB.t97 14.282
R492 VPB.n858 VPB.t78 14.282
R493 VPB.n858 VPB.t67 14.282
R494 VPB.n796 VPB.t55 14.282
R495 VPB.n796 VPB.t49 14.282
R496 VPB.n779 VPB.t45 14.282
R497 VPB.n779 VPB.t56 14.282
R498 VPB.n713 VPB.t36 14.282
R499 VPB.n713 VPB.t71 14.282
R500 VPB.n696 VPB.t83 14.282
R501 VPB.n696 VPB.t40 14.282
R502 VPB.n629 VPB.t48 14.282
R503 VPB.n629 VPB.t5 14.282
R504 VPB.n567 VPB.t60 14.282
R505 VPB.n567 VPB.t0 14.282
R506 VPB.n550 VPB.t88 14.282
R507 VPB.n550 VPB.t61 14.282
R508 VPB.n484 VPB.t89 14.282
R509 VPB.n484 VPB.t76 14.282
R510 VPB.n467 VPB.t35 14.282
R511 VPB.n467 VPB.t87 14.282
R512 VPB.n400 VPB.t46 14.282
R513 VPB.n400 VPB.t52 14.282
R514 VPB.n337 VPB.t54 14.282
R515 VPB.n337 VPB.t24 14.282
R516 VPB.n169 VPB.n168 13.653
R517 VPB.n168 VPB.n167 13.653
R518 VPB.n174 VPB.n173 13.653
R519 VPB.n173 VPB.n172 13.653
R520 VPB.n178 VPB.n177 13.653
R521 VPB.n177 VPB.n176 13.653
R522 VPB.n184 VPB.n183 13.653
R523 VPB.n183 VPB.n182 13.653
R524 VPB.n188 VPB.n187 13.653
R525 VPB.n187 VPB.n186 13.653
R526 VPB.n215 VPB.n214 13.653
R527 VPB.n214 VPB.n213 13.653
R528 VPB.n219 VPB.n218 13.653
R529 VPB.n218 VPB.n217 13.653
R530 VPB.n223 VPB.n222 13.653
R531 VPB.n222 VPB.n221 13.653
R532 VPB.n227 VPB.n226 13.653
R533 VPB.n226 VPB.n225 13.653
R534 VPB.n231 VPB.n230 13.653
R535 VPB.n230 VPB.n229 13.653
R536 VPB.n235 VPB.n234 13.653
R537 VPB.n234 VPB.n233 13.653
R538 VPB.n239 VPB.n238 13.653
R539 VPB.n238 VPB.n237 13.653
R540 VPB.n243 VPB.n242 13.653
R541 VPB.n242 VPB.n241 13.653
R542 VPB.n270 VPB.n269 13.653
R543 VPB.n269 VPB.n268 13.653
R544 VPB.n274 VPB.n273 13.653
R545 VPB.n273 VPB.n272 13.653
R546 VPB.n278 VPB.n277 13.653
R547 VPB.n277 VPB.n276 13.653
R548 VPB.n282 VPB.n281 13.653
R549 VPB.n281 VPB.n280 13.653
R550 VPB.n286 VPB.n285 13.653
R551 VPB.n285 VPB.n284 13.653
R552 VPB.n290 VPB.n289 13.653
R553 VPB.n289 VPB.n288 13.653
R554 VPB.n294 VPB.n293 13.653
R555 VPB.n293 VPB.n292 13.653
R556 VPB.n298 VPB.n297 13.653
R557 VPB.n297 VPB.n296 13.653
R558 VPB.n325 VPB.n324 13.653
R559 VPB.n324 VPB.n323 13.653
R560 VPB.n330 VPB.n329 13.653
R561 VPB.n329 VPB.n328 13.653
R562 VPB.n335 VPB.n334 13.653
R563 VPB.n334 VPB.n333 13.653
R564 VPB.n342 VPB.n341 13.653
R565 VPB.n341 VPB.n340 13.653
R566 VPB.n347 VPB.n346 13.653
R567 VPB.n346 VPB.n345 13.653
R568 VPB.n352 VPB.n351 13.653
R569 VPB.n351 VPB.n350 13.653
R570 VPB.n357 VPB.n356 13.653
R571 VPB.n356 VPB.n355 13.653
R572 VPB.n361 VPB.n360 13.653
R573 VPB.n360 VPB.n359 13.653
R574 VPB.n388 VPB.n387 13.653
R575 VPB.n387 VPB.n386 13.653
R576 VPB.n393 VPB.n392 13.653
R577 VPB.n392 VPB.n391 13.653
R578 VPB.n398 VPB.n397 13.653
R579 VPB.n397 VPB.n396 13.653
R580 VPB.n405 VPB.n404 13.653
R581 VPB.n404 VPB.n403 13.653
R582 VPB.n410 VPB.n409 13.653
R583 VPB.n409 VPB.n408 13.653
R584 VPB.n415 VPB.n414 13.653
R585 VPB.n414 VPB.n413 13.653
R586 VPB.n420 VPB.n419 13.653
R587 VPB.n419 VPB.n418 13.653
R588 VPB.n424 VPB.n423 13.653
R589 VPB.n423 VPB.n422 13.653
R590 VPB.n451 VPB.n450 13.653
R591 VPB.n450 VPB.n449 13.653
R592 VPB.n455 VPB.n454 13.653
R593 VPB.n454 VPB.n453 13.653
R594 VPB.n460 VPB.n459 13.653
R595 VPB.n459 VPB.n458 13.653
R596 VPB.n465 VPB.n464 13.653
R597 VPB.n464 VPB.n463 13.653
R598 VPB.n472 VPB.n471 13.653
R599 VPB.n471 VPB.n470 13.653
R600 VPB.n477 VPB.n476 13.653
R601 VPB.n476 VPB.n475 13.653
R602 VPB.n482 VPB.n481 13.653
R603 VPB.n481 VPB.n480 13.653
R604 VPB.n489 VPB.n488 13.653
R605 VPB.n488 VPB.n487 13.653
R606 VPB.n494 VPB.n493 13.653
R607 VPB.n493 VPB.n492 13.653
R608 VPB.n499 VPB.n498 13.653
R609 VPB.n498 VPB.n497 13.653
R610 VPB.n503 VPB.n502 13.653
R611 VPB.n502 VPB.n501 13.653
R612 VPB.n507 VPB.n506 13.653
R613 VPB.n506 VPB.n505 13.653
R614 VPB.n534 VPB.n533 13.653
R615 VPB.n533 VPB.n532 13.653
R616 VPB.n538 VPB.n537 13.653
R617 VPB.n537 VPB.n536 13.653
R618 VPB.n543 VPB.n542 13.653
R619 VPB.n542 VPB.n541 13.653
R620 VPB.n548 VPB.n547 13.653
R621 VPB.n547 VPB.n546 13.653
R622 VPB.n555 VPB.n554 13.653
R623 VPB.n554 VPB.n553 13.653
R624 VPB.n560 VPB.n559 13.653
R625 VPB.n559 VPB.n558 13.653
R626 VPB.n565 VPB.n564 13.653
R627 VPB.n564 VPB.n563 13.653
R628 VPB.n572 VPB.n571 13.653
R629 VPB.n571 VPB.n570 13.653
R630 VPB.n577 VPB.n576 13.653
R631 VPB.n576 VPB.n575 13.653
R632 VPB.n582 VPB.n581 13.653
R633 VPB.n581 VPB.n580 13.653
R634 VPB.n586 VPB.n585 13.653
R635 VPB.n585 VPB.n584 13.653
R636 VPB.n590 VPB.n589 13.653
R637 VPB.n589 VPB.n588 13.653
R638 VPB.n617 VPB.n616 13.653
R639 VPB.n616 VPB.n615 13.653
R640 VPB.n622 VPB.n621 13.653
R641 VPB.n621 VPB.n620 13.653
R642 VPB.n627 VPB.n626 13.653
R643 VPB.n626 VPB.n625 13.653
R644 VPB.n634 VPB.n633 13.653
R645 VPB.n633 VPB.n632 13.653
R646 VPB.n639 VPB.n638 13.653
R647 VPB.n638 VPB.n637 13.653
R648 VPB.n644 VPB.n643 13.653
R649 VPB.n643 VPB.n642 13.653
R650 VPB.n649 VPB.n648 13.653
R651 VPB.n648 VPB.n647 13.653
R652 VPB.n653 VPB.n652 13.653
R653 VPB.n652 VPB.n651 13.653
R654 VPB.n680 VPB.n679 13.653
R655 VPB.n679 VPB.n678 13.653
R656 VPB.n684 VPB.n683 13.653
R657 VPB.n683 VPB.n682 13.653
R658 VPB.n689 VPB.n688 13.653
R659 VPB.n688 VPB.n687 13.653
R660 VPB.n694 VPB.n693 13.653
R661 VPB.n693 VPB.n692 13.653
R662 VPB.n701 VPB.n700 13.653
R663 VPB.n700 VPB.n699 13.653
R664 VPB.n706 VPB.n705 13.653
R665 VPB.n705 VPB.n704 13.653
R666 VPB.n711 VPB.n710 13.653
R667 VPB.n710 VPB.n709 13.653
R668 VPB.n718 VPB.n717 13.653
R669 VPB.n717 VPB.n716 13.653
R670 VPB.n723 VPB.n722 13.653
R671 VPB.n722 VPB.n721 13.653
R672 VPB.n728 VPB.n727 13.653
R673 VPB.n727 VPB.n726 13.653
R674 VPB.n732 VPB.n731 13.653
R675 VPB.n731 VPB.n730 13.653
R676 VPB.n736 VPB.n735 13.653
R677 VPB.n735 VPB.n734 13.653
R678 VPB.n763 VPB.n762 13.653
R679 VPB.n762 VPB.n761 13.653
R680 VPB.n767 VPB.n766 13.653
R681 VPB.n766 VPB.n765 13.653
R682 VPB.n772 VPB.n771 13.653
R683 VPB.n771 VPB.n770 13.653
R684 VPB.n777 VPB.n776 13.653
R685 VPB.n776 VPB.n775 13.653
R686 VPB.n784 VPB.n783 13.653
R687 VPB.n783 VPB.n782 13.653
R688 VPB.n789 VPB.n788 13.653
R689 VPB.n788 VPB.n787 13.653
R690 VPB.n794 VPB.n793 13.653
R691 VPB.n793 VPB.n792 13.653
R692 VPB.n801 VPB.n800 13.653
R693 VPB.n800 VPB.n799 13.653
R694 VPB.n806 VPB.n805 13.653
R695 VPB.n805 VPB.n804 13.653
R696 VPB.n811 VPB.n810 13.653
R697 VPB.n810 VPB.n809 13.653
R698 VPB.n815 VPB.n814 13.653
R699 VPB.n814 VPB.n813 13.653
R700 VPB.n819 VPB.n818 13.653
R701 VPB.n818 VPB.n817 13.653
R702 VPB.n846 VPB.n845 13.653
R703 VPB.n845 VPB.n844 13.653
R704 VPB.n851 VPB.n850 13.653
R705 VPB.n850 VPB.n849 13.653
R706 VPB.n856 VPB.n855 13.653
R707 VPB.n855 VPB.n854 13.653
R708 VPB.n863 VPB.n862 13.653
R709 VPB.n862 VPB.n861 13.653
R710 VPB.n868 VPB.n867 13.653
R711 VPB.n867 VPB.n866 13.653
R712 VPB.n873 VPB.n872 13.653
R713 VPB.n872 VPB.n871 13.653
R714 VPB.n108 VPB.n107 13.653
R715 VPB.n107 VPB.n106 13.653
R716 VPB.n111 VPB.n110 13.653
R717 VPB.n110 VPB.n109 13.653
R718 VPB.n116 VPB.n115 13.653
R719 VPB.n115 VPB.n114 13.653
R720 VPB.n119 VPB.n118 13.653
R721 VPB.n118 VPB.n117 13.653
R722 VPB.n123 VPB.n122 13.653
R723 VPB.n122 VPB.n121 13.653
R724 VPB.n127 VPB.n126 13.653
R725 VPB.n126 VPB.n125 13.653
R726 VPB.n131 VPB.n130 13.653
R727 VPB.n130 VPB.n129 13.653
R728 VPB.n136 VPB.n135 13.653
R729 VPB.n135 VPB.n134 13.653
R730 VPB.n140 VPB.n139 13.653
R731 VPB.n139 VPB.n138 13.653
R732 VPB.n145 VPB.n144 13.653
R733 VPB.n144 VPB.n143 13.653
R734 VPB.n889 VPB.n888 13.653
R735 VPB.n888 VPB.n887 13.653
R736 VPB.n893 VPB.n892 13.653
R737 VPB.n892 VPB.n891 13.653
R738 VPB.n897 VPB.n896 13.653
R739 VPB.n896 VPB.n895 13.653
R740 VPB.n901 VPB.n900 13.653
R741 VPB.n900 VPB.n899 13.653
R742 VPB.n928 VPB.n927 13.653
R743 VPB.n927 VPB.n926 13.653
R744 VPB.n932 VPB.n931 13.653
R745 VPB.n931 VPB.n930 13.653
R746 VPB.n937 VPB.n936 13.653
R747 VPB.n936 VPB.n935 13.653
R748 VPB.n942 VPB.n941 13.653
R749 VPB.n941 VPB.n940 13.653
R750 VPB.n949 VPB.n948 13.653
R751 VPB.n948 VPB.n947 13.653
R752 VPB.n954 VPB.n953 13.653
R753 VPB.n953 VPB.n952 13.653
R754 VPB.n959 VPB.n958 13.653
R755 VPB.n958 VPB.n957 13.653
R756 VPB.n966 VPB.n965 13.653
R757 VPB.n965 VPB.n964 13.653
R758 VPB.n971 VPB.n970 13.653
R759 VPB.n970 VPB.n969 13.653
R760 VPB.n976 VPB.n975 13.653
R761 VPB.n975 VPB.n974 13.653
R762 VPB.n980 VPB.n979 13.653
R763 VPB.n979 VPB.n978 13.653
R764 VPB.n984 VPB.n983 13.653
R765 VPB.n983 VPB.n982 13.653
R766 VPB.n1011 VPB.n1010 13.653
R767 VPB.n1010 VPB.n1009 13.653
R768 VPB.n1016 VPB.n1015 13.653
R769 VPB.n1015 VPB.n1014 13.653
R770 VPB.n1021 VPB.n1020 13.653
R771 VPB.n1020 VPB.n1019 13.653
R772 VPB.n1028 VPB.n1027 13.653
R773 VPB.n1027 VPB.n1026 13.653
R774 VPB.n1033 VPB.n1032 13.653
R775 VPB.n1032 VPB.n1031 13.653
R776 VPB.n1038 VPB.n1037 13.653
R777 VPB.n1037 VPB.n1036 13.653
R778 VPB.n1043 VPB.n1042 13.653
R779 VPB.n1042 VPB.n1041 13.653
R780 VPB.n1047 VPB.n1046 13.653
R781 VPB.n1046 VPB.n1045 13.653
R782 VPB.n1074 VPB.n1073 13.653
R783 VPB.n1073 VPB.n1072 13.653
R784 VPB.n1078 VPB.n1077 13.653
R785 VPB.n1077 VPB.n1076 13.653
R786 VPB.n1083 VPB.n1082 13.653
R787 VPB.n1082 VPB.n1081 13.653
R788 VPB.n1088 VPB.n1087 13.653
R789 VPB.n1087 VPB.n1086 13.653
R790 VPB.n1095 VPB.n1094 13.653
R791 VPB.n1094 VPB.n1093 13.653
R792 VPB.n1100 VPB.n1099 13.653
R793 VPB.n1099 VPB.n1098 13.653
R794 VPB.n1105 VPB.n1104 13.653
R795 VPB.n1104 VPB.n1103 13.653
R796 VPB.n1112 VPB.n1111 13.653
R797 VPB.n1111 VPB.n1110 13.653
R798 VPB.n1117 VPB.n1116 13.653
R799 VPB.n1116 VPB.n1115 13.653
R800 VPB.n1122 VPB.n1121 13.653
R801 VPB.n1121 VPB.n1120 13.653
R802 VPB.n1126 VPB.n1125 13.653
R803 VPB.n1125 VPB.n1124 13.653
R804 VPB.n1130 VPB.n1129 13.653
R805 VPB.n1129 VPB.n1128 13.653
R806 VPB.n1157 VPB.n1156 13.653
R807 VPB.n1156 VPB.n1155 13.653
R808 VPB.n1161 VPB.n1160 13.653
R809 VPB.n1160 VPB.n1159 13.653
R810 VPB.n1166 VPB.n1165 13.653
R811 VPB.n1165 VPB.n1164 13.653
R812 VPB.n1171 VPB.n1170 13.653
R813 VPB.n1170 VPB.n1169 13.653
R814 VPB.n1178 VPB.n1177 13.653
R815 VPB.n1177 VPB.n1176 13.653
R816 VPB.n1183 VPB.n1182 13.653
R817 VPB.n1182 VPB.n1181 13.653
R818 VPB.n1188 VPB.n1187 13.653
R819 VPB.n1187 VPB.n1186 13.653
R820 VPB.n1195 VPB.n1194 13.653
R821 VPB.n1194 VPB.n1193 13.653
R822 VPB.n1200 VPB.n1199 13.653
R823 VPB.n1199 VPB.n1198 13.653
R824 VPB.n1205 VPB.n1204 13.653
R825 VPB.n1204 VPB.n1203 13.653
R826 VPB.n1209 VPB.n1208 13.653
R827 VPB.n1208 VPB.n1207 13.653
R828 VPB.n1213 VPB.n1212 13.653
R829 VPB.n1212 VPB.n1211 13.653
R830 VPB.n1240 VPB.n1239 13.653
R831 VPB.n1239 VPB.n1238 13.653
R832 VPB.n1245 VPB.n1244 13.653
R833 VPB.n1244 VPB.n1243 13.653
R834 VPB.n1250 VPB.n1249 13.653
R835 VPB.n1249 VPB.n1248 13.653
R836 VPB.n1257 VPB.n1256 13.653
R837 VPB.n1256 VPB.n1255 13.653
R838 VPB.n1262 VPB.n1261 13.653
R839 VPB.n1261 VPB.n1260 13.653
R840 VPB.n1267 VPB.n1266 13.653
R841 VPB.n1266 VPB.n1265 13.653
R842 VPB.n1272 VPB.n1271 13.653
R843 VPB.n1271 VPB.n1270 13.653
R844 VPB.n1276 VPB.n1275 13.653
R845 VPB.n1275 VPB.n1274 13.653
R846 VPB.n1303 VPB.n1302 13.653
R847 VPB.n1302 VPB.n1301 13.653
R848 VPB.n1307 VPB.n1306 13.653
R849 VPB.n1306 VPB.n1305 13.653
R850 VPB.n1312 VPB.n1311 13.653
R851 VPB.n1311 VPB.n1310 13.653
R852 VPB.n1317 VPB.n1316 13.653
R853 VPB.n1316 VPB.n1315 13.653
R854 VPB.n1324 VPB.n1323 13.653
R855 VPB.n1323 VPB.n1322 13.653
R856 VPB.n1329 VPB.n1328 13.653
R857 VPB.n1328 VPB.n1327 13.653
R858 VPB.n1334 VPB.n1333 13.653
R859 VPB.n1333 VPB.n1332 13.653
R860 VPB.n1341 VPB.n1340 13.653
R861 VPB.n1340 VPB.n1339 13.653
R862 VPB.n1346 VPB.n1345 13.653
R863 VPB.n1345 VPB.n1344 13.653
R864 VPB.n1351 VPB.n1350 13.653
R865 VPB.n1350 VPB.n1349 13.653
R866 VPB.n1355 VPB.n1354 13.653
R867 VPB.n1354 VPB.n1353 13.653
R868 VPB.n1359 VPB.n1358 13.653
R869 VPB.n1358 VPB.n1357 13.653
R870 VPB.n1386 VPB.n1385 13.653
R871 VPB.n1385 VPB.n1384 13.653
R872 VPB.n1390 VPB.n1389 13.653
R873 VPB.n1389 VPB.n1388 13.653
R874 VPB.n1395 VPB.n1394 13.653
R875 VPB.n1394 VPB.n1393 13.653
R876 VPB.n1400 VPB.n1399 13.653
R877 VPB.n1399 VPB.n1398 13.653
R878 VPB.n1407 VPB.n1406 13.653
R879 VPB.n1406 VPB.n1405 13.653
R880 VPB.n1412 VPB.n1411 13.653
R881 VPB.n1411 VPB.n1410 13.653
R882 VPB.n1417 VPB.n1416 13.653
R883 VPB.n1416 VPB.n1415 13.653
R884 VPB.n1424 VPB.n1423 13.653
R885 VPB.n1423 VPB.n1422 13.653
R886 VPB.n1429 VPB.n1428 13.653
R887 VPB.n1428 VPB.n1427 13.653
R888 VPB.n1434 VPB.n1433 13.653
R889 VPB.n1433 VPB.n1432 13.653
R890 VPB.n1438 VPB.n1437 13.653
R891 VPB.n1437 VPB.n1436 13.653
R892 VPB.n1442 VPB.n1441 13.653
R893 VPB.n1441 VPB.n1440 13.653
R894 VPB.n1469 VPB.n1468 13.653
R895 VPB.n1468 VPB.n1467 13.653
R896 VPB.n1474 VPB.n1473 13.653
R897 VPB.n1473 VPB.n1472 13.653
R898 VPB.n1479 VPB.n1478 13.653
R899 VPB.n1478 VPB.n1477 13.653
R900 VPB.n1486 VPB.n1485 13.653
R901 VPB.n1485 VPB.n1484 13.653
R902 VPB.n1491 VPB.n1490 13.653
R903 VPB.n1490 VPB.n1489 13.653
R904 VPB.n1496 VPB.n1495 13.653
R905 VPB.n1495 VPB.n1494 13.653
R906 VPB.n1501 VPB.n1500 13.653
R907 VPB.n1500 VPB.n1499 13.653
R908 VPB.n1505 VPB.n1504 13.653
R909 VPB.n1504 VPB.n1503 13.653
R910 VPB.n1532 VPB.n1531 13.653
R911 VPB.n1531 VPB.n1530 13.653
R912 VPB.n1536 VPB.n1535 13.653
R913 VPB.n1535 VPB.n1534 13.653
R914 VPB.n1541 VPB.n1540 13.653
R915 VPB.n1540 VPB.n1539 13.653
R916 VPB.n1546 VPB.n1545 13.653
R917 VPB.n1545 VPB.n1544 13.653
R918 VPB.n1553 VPB.n1552 13.653
R919 VPB.n1552 VPB.n1551 13.653
R920 VPB.n1558 VPB.n1557 13.653
R921 VPB.n1557 VPB.n1556 13.653
R922 VPB.n1563 VPB.n1562 13.653
R923 VPB.n1562 VPB.n1561 13.653
R924 VPB.n1570 VPB.n1569 13.653
R925 VPB.n1569 VPB.n1568 13.653
R926 VPB.n1575 VPB.n1574 13.653
R927 VPB.n1574 VPB.n1573 13.653
R928 VPB.n1580 VPB.n1579 13.653
R929 VPB.n1579 VPB.n1578 13.653
R930 VPB.n1584 VPB.n1583 13.653
R931 VPB.n1583 VPB.n1582 13.653
R932 VPB.n1588 VPB.n1587 13.653
R933 VPB.n1587 VPB.n1586 13.653
R934 VPB.n41 VPB.n40 13.653
R935 VPB.n40 VPB.n39 13.653
R936 VPB.n44 VPB.n43 13.653
R937 VPB.n43 VPB.n42 13.653
R938 VPB.n48 VPB.n47 13.653
R939 VPB.n47 VPB.n46 13.653
R940 VPB.n52 VPB.n51 13.653
R941 VPB.n51 VPB.n50 13.653
R942 VPB.n56 VPB.n55 13.653
R943 VPB.n55 VPB.n54 13.653
R944 VPB.n61 VPB.n60 13.653
R945 VPB.n60 VPB.n59 13.653
R946 VPB.n65 VPB.n64 13.653
R947 VPB.n64 VPB.n63 13.653
R948 VPB.n70 VPB.n69 13.653
R949 VPB.n69 VPB.n68 13.653
R950 VPB.n74 VPB.n73 13.653
R951 VPB.n73 VPB.n72 13.653
R952 VPB.n77 VPB.n76 13.653
R953 VPB.n76 VPB.n75 13.653
R954 VPB.n81 VPB.n80 13.653
R955 VPB.n80 VPB.n79 13.653
R956 VPB.n1602 VPB.n0 13.653
R957 VPB VPB.n0 13.653
R958 VPB.n345 VPB.n344 13.35
R959 VPB.n408 VPB.n407 13.35
R960 VPB.n480 VPB.n479 13.35
R961 VPB.n563 VPB.n562 13.35
R962 VPB.n637 VPB.n636 13.35
R963 VPB.n709 VPB.n708 13.35
R964 VPB.n792 VPB.n791 13.35
R965 VPB.n866 VPB.n865 13.35
R966 VPB.n138 VPB.n137 13.35
R967 VPB.n957 VPB.n956 13.35
R968 VPB.n1031 VPB.n1030 13.35
R969 VPB.n1103 VPB.n1102 13.35
R970 VPB.n1186 VPB.n1185 13.35
R971 VPB.n1260 VPB.n1259 13.35
R972 VPB.n1332 VPB.n1331 13.35
R973 VPB.n1415 VPB.n1414 13.35
R974 VPB.n1489 VPB.n1488 13.35
R975 VPB.n1561 VPB.n1560 13.35
R976 VPB.n63 VPB.n62 13.35
R977 VPB.n1606 VPB.n1605 13.276
R978 VPB.n1605 VPB.n1603 13.276
R979 VPB.n36 VPB.n18 13.276
R980 VPB.n18 VPB.n16 13.276
R981 VPB.n1527 VPB.n1509 13.276
R982 VPB.n1509 VPB.n1507 13.276
R983 VPB.n1464 VPB.n1446 13.276
R984 VPB.n1446 VPB.n1444 13.276
R985 VPB.n1381 VPB.n1363 13.276
R986 VPB.n1363 VPB.n1361 13.276
R987 VPB.n1298 VPB.n1280 13.276
R988 VPB.n1280 VPB.n1278 13.276
R989 VPB.n1235 VPB.n1217 13.276
R990 VPB.n1217 VPB.n1215 13.276
R991 VPB.n1152 VPB.n1134 13.276
R992 VPB.n1134 VPB.n1132 13.276
R993 VPB.n1069 VPB.n1051 13.276
R994 VPB.n1051 VPB.n1049 13.276
R995 VPB.n1006 VPB.n988 13.276
R996 VPB.n988 VPB.n986 13.276
R997 VPB.n923 VPB.n905 13.276
R998 VPB.n905 VPB.n903 13.276
R999 VPB.n104 VPB.n86 13.276
R1000 VPB.n86 VPB.n84 13.276
R1001 VPB.n841 VPB.n823 13.276
R1002 VPB.n823 VPB.n821 13.276
R1003 VPB.n758 VPB.n740 13.276
R1004 VPB.n740 VPB.n738 13.276
R1005 VPB.n675 VPB.n657 13.276
R1006 VPB.n657 VPB.n655 13.276
R1007 VPB.n612 VPB.n594 13.276
R1008 VPB.n594 VPB.n592 13.276
R1009 VPB.n529 VPB.n511 13.276
R1010 VPB.n511 VPB.n509 13.276
R1011 VPB.n446 VPB.n428 13.276
R1012 VPB.n428 VPB.n426 13.276
R1013 VPB.n383 VPB.n365 13.276
R1014 VPB.n365 VPB.n363 13.276
R1015 VPB.n320 VPB.n302 13.276
R1016 VPB.n302 VPB.n300 13.276
R1017 VPB.n265 VPB.n247 13.276
R1018 VPB.n247 VPB.n245 13.276
R1019 VPB.n210 VPB.n192 13.276
R1020 VPB.n192 VPB.n190 13.276
R1021 VPB.n215 VPB.n211 13.276
R1022 VPB.n270 VPB.n266 13.276
R1023 VPB.n325 VPB.n321 13.276
R1024 VPB.n388 VPB.n384 13.276
R1025 VPB.n451 VPB.n447 13.276
R1026 VPB.n534 VPB.n530 13.276
R1027 VPB.n617 VPB.n613 13.276
R1028 VPB.n680 VPB.n676 13.276
R1029 VPB.n763 VPB.n759 13.276
R1030 VPB.n846 VPB.n842 13.276
R1031 VPB.n111 VPB.n108 13.276
R1032 VPB.n112 VPB.n111 13.276
R1033 VPB.n116 VPB.n112 13.276
R1034 VPB.n119 VPB.n116 13.276
R1035 VPB.n127 VPB.n123 13.276
R1036 VPB.n131 VPB.n127 13.276
R1037 VPB.n140 VPB.n136 13.276
R1038 VPB.n889 VPB.n145 13.276
R1039 VPB.n893 VPB.n889 13.276
R1040 VPB.n928 VPB.n924 13.276
R1041 VPB.n1011 VPB.n1007 13.276
R1042 VPB.n1074 VPB.n1070 13.276
R1043 VPB.n1157 VPB.n1153 13.276
R1044 VPB.n1240 VPB.n1236 13.276
R1045 VPB.n1303 VPB.n1299 13.276
R1046 VPB.n1386 VPB.n1382 13.276
R1047 VPB.n1469 VPB.n1465 13.276
R1048 VPB.n1532 VPB.n1528 13.276
R1049 VPB.n41 VPB.n37 13.276
R1050 VPB.n44 VPB.n41 13.276
R1051 VPB.n52 VPB.n48 13.276
R1052 VPB.n56 VPB.n52 13.276
R1053 VPB.n65 VPB.n61 13.276
R1054 VPB.n74 VPB.n70 13.276
R1055 VPB.n77 VPB.n74 13.276
R1056 VPB.n1602 VPB.n81 13.276
R1057 VPB.n166 VPB.n148 13.276
R1058 VPB.n148 VPB.n146 13.276
R1059 VPB.n153 VPB.n151 12.796
R1060 VPB.n153 VPB.n152 12.564
R1061 VPB.n81 VPB.n78 12.558
R1062 VPB.n120 VPB.n119 12.2
R1063 VPB.n45 VPB.n44 12.2
R1064 VPB.n161 VPB.n160 12.198
R1065 VPB.n161 VPB.n158 12.198
R1066 VPB.n156 VPB.n155 12.198
R1067 VPB.n136 VPB.n132 9.329
R1068 VPB.n61 VPB.n57 9.329
R1069 VPB.n141 VPB.n140 8.97
R1070 VPB.n66 VPB.n65 8.97
R1071 VPB.n166 VPB.n165 7.5
R1072 VPB.n151 VPB.n150 7.5
R1073 VPB.n155 VPB.n154 7.5
R1074 VPB.n160 VPB.n159 7.5
R1075 VPB.n148 VPB.n147 7.5
R1076 VPB.n163 VPB.n149 7.5
R1077 VPB.n192 VPB.n191 7.5
R1078 VPB.n205 VPB.n204 7.5
R1079 VPB.n199 VPB.n198 7.5
R1080 VPB.n201 VPB.n200 7.5
R1081 VPB.n194 VPB.n193 7.5
R1082 VPB.n210 VPB.n209 7.5
R1083 VPB.n247 VPB.n246 7.5
R1084 VPB.n260 VPB.n259 7.5
R1085 VPB.n254 VPB.n253 7.5
R1086 VPB.n256 VPB.n255 7.5
R1087 VPB.n249 VPB.n248 7.5
R1088 VPB.n265 VPB.n264 7.5
R1089 VPB.n302 VPB.n301 7.5
R1090 VPB.n315 VPB.n314 7.5
R1091 VPB.n309 VPB.n308 7.5
R1092 VPB.n311 VPB.n310 7.5
R1093 VPB.n304 VPB.n303 7.5
R1094 VPB.n320 VPB.n319 7.5
R1095 VPB.n365 VPB.n364 7.5
R1096 VPB.n378 VPB.n377 7.5
R1097 VPB.n372 VPB.n371 7.5
R1098 VPB.n374 VPB.n373 7.5
R1099 VPB.n367 VPB.n366 7.5
R1100 VPB.n383 VPB.n382 7.5
R1101 VPB.n428 VPB.n427 7.5
R1102 VPB.n441 VPB.n440 7.5
R1103 VPB.n435 VPB.n434 7.5
R1104 VPB.n437 VPB.n436 7.5
R1105 VPB.n430 VPB.n429 7.5
R1106 VPB.n446 VPB.n445 7.5
R1107 VPB.n511 VPB.n510 7.5
R1108 VPB.n524 VPB.n523 7.5
R1109 VPB.n518 VPB.n517 7.5
R1110 VPB.n520 VPB.n519 7.5
R1111 VPB.n513 VPB.n512 7.5
R1112 VPB.n529 VPB.n528 7.5
R1113 VPB.n594 VPB.n593 7.5
R1114 VPB.n607 VPB.n606 7.5
R1115 VPB.n601 VPB.n600 7.5
R1116 VPB.n603 VPB.n602 7.5
R1117 VPB.n596 VPB.n595 7.5
R1118 VPB.n612 VPB.n611 7.5
R1119 VPB.n657 VPB.n656 7.5
R1120 VPB.n670 VPB.n669 7.5
R1121 VPB.n664 VPB.n663 7.5
R1122 VPB.n666 VPB.n665 7.5
R1123 VPB.n659 VPB.n658 7.5
R1124 VPB.n675 VPB.n674 7.5
R1125 VPB.n740 VPB.n739 7.5
R1126 VPB.n753 VPB.n752 7.5
R1127 VPB.n747 VPB.n746 7.5
R1128 VPB.n749 VPB.n748 7.5
R1129 VPB.n742 VPB.n741 7.5
R1130 VPB.n758 VPB.n757 7.5
R1131 VPB.n823 VPB.n822 7.5
R1132 VPB.n836 VPB.n835 7.5
R1133 VPB.n830 VPB.n829 7.5
R1134 VPB.n832 VPB.n831 7.5
R1135 VPB.n825 VPB.n824 7.5
R1136 VPB.n841 VPB.n840 7.5
R1137 VPB.n86 VPB.n85 7.5
R1138 VPB.n99 VPB.n98 7.5
R1139 VPB.n93 VPB.n92 7.5
R1140 VPB.n95 VPB.n94 7.5
R1141 VPB.n88 VPB.n87 7.5
R1142 VPB.n104 VPB.n103 7.5
R1143 VPB.n905 VPB.n904 7.5
R1144 VPB.n918 VPB.n917 7.5
R1145 VPB.n912 VPB.n911 7.5
R1146 VPB.n914 VPB.n913 7.5
R1147 VPB.n907 VPB.n906 7.5
R1148 VPB.n923 VPB.n922 7.5
R1149 VPB.n988 VPB.n987 7.5
R1150 VPB.n1001 VPB.n1000 7.5
R1151 VPB.n995 VPB.n994 7.5
R1152 VPB.n997 VPB.n996 7.5
R1153 VPB.n990 VPB.n989 7.5
R1154 VPB.n1006 VPB.n1005 7.5
R1155 VPB.n1051 VPB.n1050 7.5
R1156 VPB.n1064 VPB.n1063 7.5
R1157 VPB.n1058 VPB.n1057 7.5
R1158 VPB.n1060 VPB.n1059 7.5
R1159 VPB.n1053 VPB.n1052 7.5
R1160 VPB.n1069 VPB.n1068 7.5
R1161 VPB.n1134 VPB.n1133 7.5
R1162 VPB.n1147 VPB.n1146 7.5
R1163 VPB.n1141 VPB.n1140 7.5
R1164 VPB.n1143 VPB.n1142 7.5
R1165 VPB.n1136 VPB.n1135 7.5
R1166 VPB.n1152 VPB.n1151 7.5
R1167 VPB.n1217 VPB.n1216 7.5
R1168 VPB.n1230 VPB.n1229 7.5
R1169 VPB.n1224 VPB.n1223 7.5
R1170 VPB.n1226 VPB.n1225 7.5
R1171 VPB.n1219 VPB.n1218 7.5
R1172 VPB.n1235 VPB.n1234 7.5
R1173 VPB.n1280 VPB.n1279 7.5
R1174 VPB.n1293 VPB.n1292 7.5
R1175 VPB.n1287 VPB.n1286 7.5
R1176 VPB.n1289 VPB.n1288 7.5
R1177 VPB.n1282 VPB.n1281 7.5
R1178 VPB.n1298 VPB.n1297 7.5
R1179 VPB.n1363 VPB.n1362 7.5
R1180 VPB.n1376 VPB.n1375 7.5
R1181 VPB.n1370 VPB.n1369 7.5
R1182 VPB.n1372 VPB.n1371 7.5
R1183 VPB.n1365 VPB.n1364 7.5
R1184 VPB.n1381 VPB.n1380 7.5
R1185 VPB.n1446 VPB.n1445 7.5
R1186 VPB.n1459 VPB.n1458 7.5
R1187 VPB.n1453 VPB.n1452 7.5
R1188 VPB.n1455 VPB.n1454 7.5
R1189 VPB.n1448 VPB.n1447 7.5
R1190 VPB.n1464 VPB.n1463 7.5
R1191 VPB.n1509 VPB.n1508 7.5
R1192 VPB.n1522 VPB.n1521 7.5
R1193 VPB.n1516 VPB.n1515 7.5
R1194 VPB.n1518 VPB.n1517 7.5
R1195 VPB.n1511 VPB.n1510 7.5
R1196 VPB.n1527 VPB.n1526 7.5
R1197 VPB.n18 VPB.n17 7.5
R1198 VPB.n31 VPB.n30 7.5
R1199 VPB.n25 VPB.n24 7.5
R1200 VPB.n27 VPB.n26 7.5
R1201 VPB.n20 VPB.n19 7.5
R1202 VPB.n36 VPB.n35 7.5
R1203 VPB.n1605 VPB.n1604 7.5
R1204 VPB.n12 VPB.n11 7.5
R1205 VPB.n6 VPB.n5 7.5
R1206 VPB.n8 VPB.n7 7.5
R1207 VPB.n2 VPB.n1 7.5
R1208 VPB.n1607 VPB.n1606 7.5
R1209 VPB.n37 VPB.n36 7.176
R1210 VPB.n1528 VPB.n1527 7.176
R1211 VPB.n1465 VPB.n1464 7.176
R1212 VPB.n1382 VPB.n1381 7.176
R1213 VPB.n1299 VPB.n1298 7.176
R1214 VPB.n1236 VPB.n1235 7.176
R1215 VPB.n1153 VPB.n1152 7.176
R1216 VPB.n1070 VPB.n1069 7.176
R1217 VPB.n1007 VPB.n1006 7.176
R1218 VPB.n924 VPB.n923 7.176
R1219 VPB.n112 VPB.n104 7.176
R1220 VPB.n842 VPB.n841 7.176
R1221 VPB.n759 VPB.n758 7.176
R1222 VPB.n676 VPB.n675 7.176
R1223 VPB.n613 VPB.n612 7.176
R1224 VPB.n530 VPB.n529 7.176
R1225 VPB.n447 VPB.n446 7.176
R1226 VPB.n384 VPB.n383 7.176
R1227 VPB.n321 VPB.n320 7.176
R1228 VPB.n266 VPB.n265 7.176
R1229 VPB.n211 VPB.n210 7.176
R1230 VPB.n206 VPB.n203 6.729
R1231 VPB.n202 VPB.n199 6.729
R1232 VPB.n197 VPB.n194 6.729
R1233 VPB.n261 VPB.n258 6.729
R1234 VPB.n257 VPB.n254 6.729
R1235 VPB.n252 VPB.n249 6.729
R1236 VPB.n316 VPB.n313 6.729
R1237 VPB.n312 VPB.n309 6.729
R1238 VPB.n307 VPB.n304 6.729
R1239 VPB.n379 VPB.n376 6.729
R1240 VPB.n375 VPB.n372 6.729
R1241 VPB.n370 VPB.n367 6.729
R1242 VPB.n442 VPB.n439 6.729
R1243 VPB.n438 VPB.n435 6.729
R1244 VPB.n433 VPB.n430 6.729
R1245 VPB.n525 VPB.n522 6.729
R1246 VPB.n521 VPB.n518 6.729
R1247 VPB.n516 VPB.n513 6.729
R1248 VPB.n608 VPB.n605 6.729
R1249 VPB.n604 VPB.n601 6.729
R1250 VPB.n599 VPB.n596 6.729
R1251 VPB.n671 VPB.n668 6.729
R1252 VPB.n667 VPB.n664 6.729
R1253 VPB.n662 VPB.n659 6.729
R1254 VPB.n754 VPB.n751 6.729
R1255 VPB.n750 VPB.n747 6.729
R1256 VPB.n745 VPB.n742 6.729
R1257 VPB.n837 VPB.n834 6.729
R1258 VPB.n833 VPB.n830 6.729
R1259 VPB.n828 VPB.n825 6.729
R1260 VPB.n100 VPB.n97 6.729
R1261 VPB.n96 VPB.n93 6.729
R1262 VPB.n91 VPB.n88 6.729
R1263 VPB.n919 VPB.n916 6.729
R1264 VPB.n915 VPB.n912 6.729
R1265 VPB.n910 VPB.n907 6.729
R1266 VPB.n1002 VPB.n999 6.729
R1267 VPB.n998 VPB.n995 6.729
R1268 VPB.n993 VPB.n990 6.729
R1269 VPB.n1065 VPB.n1062 6.729
R1270 VPB.n1061 VPB.n1058 6.729
R1271 VPB.n1056 VPB.n1053 6.729
R1272 VPB.n1148 VPB.n1145 6.729
R1273 VPB.n1144 VPB.n1141 6.729
R1274 VPB.n1139 VPB.n1136 6.729
R1275 VPB.n1231 VPB.n1228 6.729
R1276 VPB.n1227 VPB.n1224 6.729
R1277 VPB.n1222 VPB.n1219 6.729
R1278 VPB.n1294 VPB.n1291 6.729
R1279 VPB.n1290 VPB.n1287 6.729
R1280 VPB.n1285 VPB.n1282 6.729
R1281 VPB.n1377 VPB.n1374 6.729
R1282 VPB.n1373 VPB.n1370 6.729
R1283 VPB.n1368 VPB.n1365 6.729
R1284 VPB.n1460 VPB.n1457 6.729
R1285 VPB.n1456 VPB.n1453 6.729
R1286 VPB.n1451 VPB.n1448 6.729
R1287 VPB.n1523 VPB.n1520 6.729
R1288 VPB.n1519 VPB.n1516 6.729
R1289 VPB.n1514 VPB.n1511 6.729
R1290 VPB.n32 VPB.n29 6.729
R1291 VPB.n28 VPB.n25 6.729
R1292 VPB.n23 VPB.n20 6.729
R1293 VPB.n13 VPB.n10 6.729
R1294 VPB.n9 VPB.n6 6.729
R1295 VPB.n4 VPB.n2 6.729
R1296 VPB.n197 VPB.n196 6.728
R1297 VPB.n202 VPB.n201 6.728
R1298 VPB.n206 VPB.n205 6.728
R1299 VPB.n209 VPB.n208 6.728
R1300 VPB.n252 VPB.n251 6.728
R1301 VPB.n257 VPB.n256 6.728
R1302 VPB.n261 VPB.n260 6.728
R1303 VPB.n264 VPB.n263 6.728
R1304 VPB.n307 VPB.n306 6.728
R1305 VPB.n312 VPB.n311 6.728
R1306 VPB.n316 VPB.n315 6.728
R1307 VPB.n319 VPB.n318 6.728
R1308 VPB.n370 VPB.n369 6.728
R1309 VPB.n375 VPB.n374 6.728
R1310 VPB.n379 VPB.n378 6.728
R1311 VPB.n382 VPB.n381 6.728
R1312 VPB.n433 VPB.n432 6.728
R1313 VPB.n438 VPB.n437 6.728
R1314 VPB.n442 VPB.n441 6.728
R1315 VPB.n445 VPB.n444 6.728
R1316 VPB.n516 VPB.n515 6.728
R1317 VPB.n521 VPB.n520 6.728
R1318 VPB.n525 VPB.n524 6.728
R1319 VPB.n528 VPB.n527 6.728
R1320 VPB.n599 VPB.n598 6.728
R1321 VPB.n604 VPB.n603 6.728
R1322 VPB.n608 VPB.n607 6.728
R1323 VPB.n611 VPB.n610 6.728
R1324 VPB.n662 VPB.n661 6.728
R1325 VPB.n667 VPB.n666 6.728
R1326 VPB.n671 VPB.n670 6.728
R1327 VPB.n674 VPB.n673 6.728
R1328 VPB.n745 VPB.n744 6.728
R1329 VPB.n750 VPB.n749 6.728
R1330 VPB.n754 VPB.n753 6.728
R1331 VPB.n757 VPB.n756 6.728
R1332 VPB.n828 VPB.n827 6.728
R1333 VPB.n833 VPB.n832 6.728
R1334 VPB.n837 VPB.n836 6.728
R1335 VPB.n840 VPB.n839 6.728
R1336 VPB.n91 VPB.n90 6.728
R1337 VPB.n96 VPB.n95 6.728
R1338 VPB.n100 VPB.n99 6.728
R1339 VPB.n103 VPB.n102 6.728
R1340 VPB.n910 VPB.n909 6.728
R1341 VPB.n915 VPB.n914 6.728
R1342 VPB.n919 VPB.n918 6.728
R1343 VPB.n922 VPB.n921 6.728
R1344 VPB.n993 VPB.n992 6.728
R1345 VPB.n998 VPB.n997 6.728
R1346 VPB.n1002 VPB.n1001 6.728
R1347 VPB.n1005 VPB.n1004 6.728
R1348 VPB.n1056 VPB.n1055 6.728
R1349 VPB.n1061 VPB.n1060 6.728
R1350 VPB.n1065 VPB.n1064 6.728
R1351 VPB.n1068 VPB.n1067 6.728
R1352 VPB.n1139 VPB.n1138 6.728
R1353 VPB.n1144 VPB.n1143 6.728
R1354 VPB.n1148 VPB.n1147 6.728
R1355 VPB.n1151 VPB.n1150 6.728
R1356 VPB.n1222 VPB.n1221 6.728
R1357 VPB.n1227 VPB.n1226 6.728
R1358 VPB.n1231 VPB.n1230 6.728
R1359 VPB.n1234 VPB.n1233 6.728
R1360 VPB.n1285 VPB.n1284 6.728
R1361 VPB.n1290 VPB.n1289 6.728
R1362 VPB.n1294 VPB.n1293 6.728
R1363 VPB.n1297 VPB.n1296 6.728
R1364 VPB.n1368 VPB.n1367 6.728
R1365 VPB.n1373 VPB.n1372 6.728
R1366 VPB.n1377 VPB.n1376 6.728
R1367 VPB.n1380 VPB.n1379 6.728
R1368 VPB.n1451 VPB.n1450 6.728
R1369 VPB.n1456 VPB.n1455 6.728
R1370 VPB.n1460 VPB.n1459 6.728
R1371 VPB.n1463 VPB.n1462 6.728
R1372 VPB.n1514 VPB.n1513 6.728
R1373 VPB.n1519 VPB.n1518 6.728
R1374 VPB.n1523 VPB.n1522 6.728
R1375 VPB.n1526 VPB.n1525 6.728
R1376 VPB.n23 VPB.n22 6.728
R1377 VPB.n28 VPB.n27 6.728
R1378 VPB.n32 VPB.n31 6.728
R1379 VPB.n35 VPB.n34 6.728
R1380 VPB.n4 VPB.n3 6.728
R1381 VPB.n9 VPB.n8 6.728
R1382 VPB.n13 VPB.n12 6.728
R1383 VPB.n1608 VPB.n1607 6.728
R1384 VPB.n342 VPB.n338 6.458
R1385 VPB.n405 VPB.n401 6.458
R1386 VPB.n634 VPB.n630 6.458
R1387 VPB.n863 VPB.n859 6.458
R1388 VPB.n1028 VPB.n1024 6.458
R1389 VPB.n1257 VPB.n1253 6.458
R1390 VPB.n1486 VPB.n1482 6.458
R1391 VPB.n165 VPB.n164 6.398
R1392 VPB.n489 VPB.n485 4.305
R1393 VPB.n572 VPB.n568 4.305
R1394 VPB.n718 VPB.n714 4.305
R1395 VPB.n801 VPB.n797 4.305
R1396 VPB.n145 VPB.n141 4.305
R1397 VPB.n966 VPB.n962 4.305
R1398 VPB.n1112 VPB.n1108 4.305
R1399 VPB.n1195 VPB.n1191 4.305
R1400 VPB.n1341 VPB.n1337 4.305
R1401 VPB.n1424 VPB.n1420 4.305
R1402 VPB.n1570 VPB.n1566 4.305
R1403 VPB.n70 VPB.n66 4.305
R1404 VPB.n472 VPB.n468 3.947
R1405 VPB.n555 VPB.n551 3.947
R1406 VPB.n701 VPB.n697 3.947
R1407 VPB.n784 VPB.n780 3.947
R1408 VPB.n132 VPB.n131 3.947
R1409 VPB.n949 VPB.n945 3.947
R1410 VPB.n1095 VPB.n1091 3.947
R1411 VPB.n1178 VPB.n1174 3.947
R1412 VPB.n1324 VPB.n1320 3.947
R1413 VPB.n1407 VPB.n1403 3.947
R1414 VPB.n1553 VPB.n1549 3.947
R1415 VPB.n57 VPB.n56 3.947
R1416 VPB.n174 VPB.n170 2.691
R1417 VPB.n184 VPB.n180 2.332
R1418 VPB.n357 VPB.n354 1.794
R1419 VPB.n420 VPB.n417 1.794
R1420 VPB.n649 VPB.n646 1.794
R1421 VPB.n108 VPB.n105 1.794
R1422 VPB.n1043 VPB.n1040 1.794
R1423 VPB.n1272 VPB.n1269 1.794
R1424 VPB.n1501 VPB.n1498 1.794
R1425 VPB.n330 VPB.n327 1.435
R1426 VPB.n393 VPB.n390 1.435
R1427 VPB.n622 VPB.n619 1.435
R1428 VPB.n851 VPB.n848 1.435
R1429 VPB.n1016 VPB.n1013 1.435
R1430 VPB.n1245 VPB.n1242 1.435
R1431 VPB.n1474 VPB.n1471 1.435
R1432 VPB.n163 VPB.n156 1.402
R1433 VPB.n163 VPB.n157 1.402
R1434 VPB.n163 VPB.n161 1.402
R1435 VPB.n163 VPB.n162 1.402
R1436 VPB.n460 VPB.n457 1.076
R1437 VPB.n543 VPB.n540 1.076
R1438 VPB.n689 VPB.n686 1.076
R1439 VPB.n772 VPB.n769 1.076
R1440 VPB.n123 VPB.n120 1.076
R1441 VPB.n937 VPB.n934 1.076
R1442 VPB.n1083 VPB.n1080 1.076
R1443 VPB.n1166 VPB.n1163 1.076
R1444 VPB.n1312 VPB.n1309 1.076
R1445 VPB.n1395 VPB.n1392 1.076
R1446 VPB.n1541 VPB.n1538 1.076
R1447 VPB.n48 VPB.n45 1.076
R1448 VPB.n164 VPB.n163 0.735
R1449 VPB.n163 VPB.n153 0.735
R1450 VPB.n499 VPB.n496 0.717
R1451 VPB.n582 VPB.n579 0.717
R1452 VPB.n728 VPB.n725 0.717
R1453 VPB.n811 VPB.n808 0.717
R1454 VPB.n893 VPB.n890 0.717
R1455 VPB.n976 VPB.n973 0.717
R1456 VPB.n1122 VPB.n1119 0.717
R1457 VPB.n1205 VPB.n1202 0.717
R1458 VPB.n1351 VPB.n1348 0.717
R1459 VPB.n1434 VPB.n1431 0.717
R1460 VPB.n1580 VPB.n1577 0.717
R1461 VPB.n78 VPB.n77 0.717
R1462 VPB.n207 VPB.n206 0.387
R1463 VPB.n207 VPB.n202 0.387
R1464 VPB.n207 VPB.n197 0.387
R1465 VPB.n208 VPB.n207 0.387
R1466 VPB.n262 VPB.n261 0.387
R1467 VPB.n262 VPB.n257 0.387
R1468 VPB.n262 VPB.n252 0.387
R1469 VPB.n263 VPB.n262 0.387
R1470 VPB.n317 VPB.n316 0.387
R1471 VPB.n317 VPB.n312 0.387
R1472 VPB.n317 VPB.n307 0.387
R1473 VPB.n318 VPB.n317 0.387
R1474 VPB.n380 VPB.n379 0.387
R1475 VPB.n380 VPB.n375 0.387
R1476 VPB.n380 VPB.n370 0.387
R1477 VPB.n381 VPB.n380 0.387
R1478 VPB.n443 VPB.n442 0.387
R1479 VPB.n443 VPB.n438 0.387
R1480 VPB.n443 VPB.n433 0.387
R1481 VPB.n444 VPB.n443 0.387
R1482 VPB.n526 VPB.n525 0.387
R1483 VPB.n526 VPB.n521 0.387
R1484 VPB.n526 VPB.n516 0.387
R1485 VPB.n527 VPB.n526 0.387
R1486 VPB.n609 VPB.n608 0.387
R1487 VPB.n609 VPB.n604 0.387
R1488 VPB.n609 VPB.n599 0.387
R1489 VPB.n610 VPB.n609 0.387
R1490 VPB.n672 VPB.n671 0.387
R1491 VPB.n672 VPB.n667 0.387
R1492 VPB.n672 VPB.n662 0.387
R1493 VPB.n673 VPB.n672 0.387
R1494 VPB.n755 VPB.n754 0.387
R1495 VPB.n755 VPB.n750 0.387
R1496 VPB.n755 VPB.n745 0.387
R1497 VPB.n756 VPB.n755 0.387
R1498 VPB.n838 VPB.n837 0.387
R1499 VPB.n838 VPB.n833 0.387
R1500 VPB.n838 VPB.n828 0.387
R1501 VPB.n839 VPB.n838 0.387
R1502 VPB.n101 VPB.n100 0.387
R1503 VPB.n101 VPB.n96 0.387
R1504 VPB.n101 VPB.n91 0.387
R1505 VPB.n102 VPB.n101 0.387
R1506 VPB.n920 VPB.n919 0.387
R1507 VPB.n920 VPB.n915 0.387
R1508 VPB.n920 VPB.n910 0.387
R1509 VPB.n921 VPB.n920 0.387
R1510 VPB.n1003 VPB.n1002 0.387
R1511 VPB.n1003 VPB.n998 0.387
R1512 VPB.n1003 VPB.n993 0.387
R1513 VPB.n1004 VPB.n1003 0.387
R1514 VPB.n1066 VPB.n1065 0.387
R1515 VPB.n1066 VPB.n1061 0.387
R1516 VPB.n1066 VPB.n1056 0.387
R1517 VPB.n1067 VPB.n1066 0.387
R1518 VPB.n1149 VPB.n1148 0.387
R1519 VPB.n1149 VPB.n1144 0.387
R1520 VPB.n1149 VPB.n1139 0.387
R1521 VPB.n1150 VPB.n1149 0.387
R1522 VPB.n1232 VPB.n1231 0.387
R1523 VPB.n1232 VPB.n1227 0.387
R1524 VPB.n1232 VPB.n1222 0.387
R1525 VPB.n1233 VPB.n1232 0.387
R1526 VPB.n1295 VPB.n1294 0.387
R1527 VPB.n1295 VPB.n1290 0.387
R1528 VPB.n1295 VPB.n1285 0.387
R1529 VPB.n1296 VPB.n1295 0.387
R1530 VPB.n1378 VPB.n1377 0.387
R1531 VPB.n1378 VPB.n1373 0.387
R1532 VPB.n1378 VPB.n1368 0.387
R1533 VPB.n1379 VPB.n1378 0.387
R1534 VPB.n1461 VPB.n1460 0.387
R1535 VPB.n1461 VPB.n1456 0.387
R1536 VPB.n1461 VPB.n1451 0.387
R1537 VPB.n1462 VPB.n1461 0.387
R1538 VPB.n1524 VPB.n1523 0.387
R1539 VPB.n1524 VPB.n1519 0.387
R1540 VPB.n1524 VPB.n1514 0.387
R1541 VPB.n1525 VPB.n1524 0.387
R1542 VPB.n33 VPB.n32 0.387
R1543 VPB.n33 VPB.n28 0.387
R1544 VPB.n33 VPB.n23 0.387
R1545 VPB.n34 VPB.n33 0.387
R1546 VPB.n1609 VPB.n13 0.387
R1547 VPB.n1609 VPB.n9 0.387
R1548 VPB.n1609 VPB.n4 0.387
R1549 VPB.n1609 VPB.n1608 0.387
R1550 VPB.n216 VPB.n189 0.272
R1551 VPB.n271 VPB.n244 0.272
R1552 VPB.n326 VPB.n299 0.272
R1553 VPB.n389 VPB.n362 0.272
R1554 VPB.n452 VPB.n425 0.272
R1555 VPB.n535 VPB.n508 0.272
R1556 VPB.n618 VPB.n591 0.272
R1557 VPB.n681 VPB.n654 0.272
R1558 VPB.n764 VPB.n737 0.272
R1559 VPB.n847 VPB.n820 0.272
R1560 VPB.n877 VPB.n876 0.272
R1561 VPB.n929 VPB.n902 0.272
R1562 VPB.n1012 VPB.n985 0.272
R1563 VPB.n1075 VPB.n1048 0.272
R1564 VPB.n1158 VPB.n1131 0.272
R1565 VPB.n1241 VPB.n1214 0.272
R1566 VPB.n1304 VPB.n1277 0.272
R1567 VPB.n1387 VPB.n1360 0.272
R1568 VPB.n1470 VPB.n1443 0.272
R1569 VPB.n1533 VPB.n1506 0.272
R1570 VPB.n1590 VPB.n1589 0.272
R1571 VPB.n1601 VPB 0.198
R1572 VPB.n179 VPB.n175 0.136
R1573 VPB.n185 VPB.n179 0.136
R1574 VPB.n189 VPB.n185 0.136
R1575 VPB.n220 VPB.n216 0.136
R1576 VPB.n224 VPB.n220 0.136
R1577 VPB.n228 VPB.n224 0.136
R1578 VPB.n232 VPB.n228 0.136
R1579 VPB.n236 VPB.n232 0.136
R1580 VPB.n240 VPB.n236 0.136
R1581 VPB.n244 VPB.n240 0.136
R1582 VPB.n275 VPB.n271 0.136
R1583 VPB.n279 VPB.n275 0.136
R1584 VPB.n283 VPB.n279 0.136
R1585 VPB.n287 VPB.n283 0.136
R1586 VPB.n291 VPB.n287 0.136
R1587 VPB.n295 VPB.n291 0.136
R1588 VPB.n299 VPB.n295 0.136
R1589 VPB.n331 VPB.n326 0.136
R1590 VPB.n336 VPB.n331 0.136
R1591 VPB.n343 VPB.n336 0.136
R1592 VPB.n348 VPB.n343 0.136
R1593 VPB.n353 VPB.n348 0.136
R1594 VPB.n358 VPB.n353 0.136
R1595 VPB.n362 VPB.n358 0.136
R1596 VPB.n394 VPB.n389 0.136
R1597 VPB.n399 VPB.n394 0.136
R1598 VPB.n406 VPB.n399 0.136
R1599 VPB.n411 VPB.n406 0.136
R1600 VPB.n416 VPB.n411 0.136
R1601 VPB.n421 VPB.n416 0.136
R1602 VPB.n425 VPB.n421 0.136
R1603 VPB.n456 VPB.n452 0.136
R1604 VPB.n461 VPB.n456 0.136
R1605 VPB.n466 VPB.n461 0.136
R1606 VPB.n473 VPB.n466 0.136
R1607 VPB.n478 VPB.n473 0.136
R1608 VPB.n483 VPB.n478 0.136
R1609 VPB.n490 VPB.n483 0.136
R1610 VPB.n495 VPB.n490 0.136
R1611 VPB.n500 VPB.n495 0.136
R1612 VPB.n504 VPB.n500 0.136
R1613 VPB.n508 VPB.n504 0.136
R1614 VPB.n539 VPB.n535 0.136
R1615 VPB.n544 VPB.n539 0.136
R1616 VPB.n549 VPB.n544 0.136
R1617 VPB.n556 VPB.n549 0.136
R1618 VPB.n561 VPB.n556 0.136
R1619 VPB.n566 VPB.n561 0.136
R1620 VPB.n573 VPB.n566 0.136
R1621 VPB.n578 VPB.n573 0.136
R1622 VPB.n583 VPB.n578 0.136
R1623 VPB.n587 VPB.n583 0.136
R1624 VPB.n591 VPB.n587 0.136
R1625 VPB.n623 VPB.n618 0.136
R1626 VPB.n628 VPB.n623 0.136
R1627 VPB.n635 VPB.n628 0.136
R1628 VPB.n640 VPB.n635 0.136
R1629 VPB.n645 VPB.n640 0.136
R1630 VPB.n650 VPB.n645 0.136
R1631 VPB.n654 VPB.n650 0.136
R1632 VPB.n685 VPB.n681 0.136
R1633 VPB.n690 VPB.n685 0.136
R1634 VPB.n695 VPB.n690 0.136
R1635 VPB.n702 VPB.n695 0.136
R1636 VPB.n707 VPB.n702 0.136
R1637 VPB.n712 VPB.n707 0.136
R1638 VPB.n719 VPB.n712 0.136
R1639 VPB.n724 VPB.n719 0.136
R1640 VPB.n729 VPB.n724 0.136
R1641 VPB.n733 VPB.n729 0.136
R1642 VPB.n737 VPB.n733 0.136
R1643 VPB.n768 VPB.n764 0.136
R1644 VPB.n773 VPB.n768 0.136
R1645 VPB.n778 VPB.n773 0.136
R1646 VPB.n785 VPB.n778 0.136
R1647 VPB.n790 VPB.n785 0.136
R1648 VPB.n795 VPB.n790 0.136
R1649 VPB.n802 VPB.n795 0.136
R1650 VPB.n807 VPB.n802 0.136
R1651 VPB.n812 VPB.n807 0.136
R1652 VPB.n816 VPB.n812 0.136
R1653 VPB.n820 VPB.n816 0.136
R1654 VPB.n852 VPB.n847 0.136
R1655 VPB.n857 VPB.n852 0.136
R1656 VPB.n864 VPB.n857 0.136
R1657 VPB.n869 VPB.n864 0.136
R1658 VPB.n874 VPB.n869 0.136
R1659 VPB.n875 VPB.n874 0.136
R1660 VPB.n876 VPB.n875 0.136
R1661 VPB.n878 VPB.n877 0.136
R1662 VPB.n879 VPB.n878 0.136
R1663 VPB.n880 VPB.n879 0.136
R1664 VPB.n881 VPB.n880 0.136
R1665 VPB.n882 VPB.n881 0.136
R1666 VPB.n883 VPB.n882 0.136
R1667 VPB.n884 VPB.n883 0.136
R1668 VPB.n885 VPB.n884 0.136
R1669 VPB.n898 VPB.n894 0.136
R1670 VPB.n902 VPB.n898 0.136
R1671 VPB.n933 VPB.n929 0.136
R1672 VPB.n938 VPB.n933 0.136
R1673 VPB.n943 VPB.n938 0.136
R1674 VPB.n950 VPB.n943 0.136
R1675 VPB.n955 VPB.n950 0.136
R1676 VPB.n960 VPB.n955 0.136
R1677 VPB.n967 VPB.n960 0.136
R1678 VPB.n972 VPB.n967 0.136
R1679 VPB.n977 VPB.n972 0.136
R1680 VPB.n981 VPB.n977 0.136
R1681 VPB.n985 VPB.n981 0.136
R1682 VPB.n1017 VPB.n1012 0.136
R1683 VPB.n1022 VPB.n1017 0.136
R1684 VPB.n1029 VPB.n1022 0.136
R1685 VPB.n1034 VPB.n1029 0.136
R1686 VPB.n1039 VPB.n1034 0.136
R1687 VPB.n1044 VPB.n1039 0.136
R1688 VPB.n1048 VPB.n1044 0.136
R1689 VPB.n1079 VPB.n1075 0.136
R1690 VPB.n1084 VPB.n1079 0.136
R1691 VPB.n1089 VPB.n1084 0.136
R1692 VPB.n1096 VPB.n1089 0.136
R1693 VPB.n1101 VPB.n1096 0.136
R1694 VPB.n1106 VPB.n1101 0.136
R1695 VPB.n1113 VPB.n1106 0.136
R1696 VPB.n1118 VPB.n1113 0.136
R1697 VPB.n1123 VPB.n1118 0.136
R1698 VPB.n1127 VPB.n1123 0.136
R1699 VPB.n1131 VPB.n1127 0.136
R1700 VPB.n1162 VPB.n1158 0.136
R1701 VPB.n1167 VPB.n1162 0.136
R1702 VPB.n1172 VPB.n1167 0.136
R1703 VPB.n1179 VPB.n1172 0.136
R1704 VPB.n1184 VPB.n1179 0.136
R1705 VPB.n1189 VPB.n1184 0.136
R1706 VPB.n1196 VPB.n1189 0.136
R1707 VPB.n1201 VPB.n1196 0.136
R1708 VPB.n1206 VPB.n1201 0.136
R1709 VPB.n1210 VPB.n1206 0.136
R1710 VPB.n1214 VPB.n1210 0.136
R1711 VPB.n1246 VPB.n1241 0.136
R1712 VPB.n1251 VPB.n1246 0.136
R1713 VPB.n1258 VPB.n1251 0.136
R1714 VPB.n1263 VPB.n1258 0.136
R1715 VPB.n1268 VPB.n1263 0.136
R1716 VPB.n1273 VPB.n1268 0.136
R1717 VPB.n1277 VPB.n1273 0.136
R1718 VPB.n1308 VPB.n1304 0.136
R1719 VPB.n1313 VPB.n1308 0.136
R1720 VPB.n1318 VPB.n1313 0.136
R1721 VPB.n1325 VPB.n1318 0.136
R1722 VPB.n1330 VPB.n1325 0.136
R1723 VPB.n1335 VPB.n1330 0.136
R1724 VPB.n1342 VPB.n1335 0.136
R1725 VPB.n1347 VPB.n1342 0.136
R1726 VPB.n1352 VPB.n1347 0.136
R1727 VPB.n1356 VPB.n1352 0.136
R1728 VPB.n1360 VPB.n1356 0.136
R1729 VPB.n1391 VPB.n1387 0.136
R1730 VPB.n1396 VPB.n1391 0.136
R1731 VPB.n1401 VPB.n1396 0.136
R1732 VPB.n1408 VPB.n1401 0.136
R1733 VPB.n1413 VPB.n1408 0.136
R1734 VPB.n1418 VPB.n1413 0.136
R1735 VPB.n1425 VPB.n1418 0.136
R1736 VPB.n1430 VPB.n1425 0.136
R1737 VPB.n1435 VPB.n1430 0.136
R1738 VPB.n1439 VPB.n1435 0.136
R1739 VPB.n1443 VPB.n1439 0.136
R1740 VPB.n1475 VPB.n1470 0.136
R1741 VPB.n1480 VPB.n1475 0.136
R1742 VPB.n1487 VPB.n1480 0.136
R1743 VPB.n1492 VPB.n1487 0.136
R1744 VPB.n1497 VPB.n1492 0.136
R1745 VPB.n1502 VPB.n1497 0.136
R1746 VPB.n1506 VPB.n1502 0.136
R1747 VPB.n1537 VPB.n1533 0.136
R1748 VPB.n1542 VPB.n1537 0.136
R1749 VPB.n1547 VPB.n1542 0.136
R1750 VPB.n1554 VPB.n1547 0.136
R1751 VPB.n1559 VPB.n1554 0.136
R1752 VPB.n1564 VPB.n1559 0.136
R1753 VPB.n1571 VPB.n1564 0.136
R1754 VPB.n1576 VPB.n1571 0.136
R1755 VPB.n1581 VPB.n1576 0.136
R1756 VPB.n1585 VPB.n1581 0.136
R1757 VPB.n1589 VPB.n1585 0.136
R1758 VPB.n1591 VPB.n1590 0.136
R1759 VPB.n1592 VPB.n1591 0.136
R1760 VPB.n1593 VPB.n1592 0.136
R1761 VPB.n1594 VPB.n1593 0.136
R1762 VPB.n1595 VPB.n1594 0.136
R1763 VPB.n1596 VPB.n1595 0.136
R1764 VPB.n1597 VPB.n1596 0.136
R1765 VPB.n1598 VPB.n1597 0.136
R1766 VPB.n1599 VPB.n1598 0.136
R1767 VPB.n1600 VPB.n1599 0.136
R1768 VPB.n1601 VPB.n1600 0.136
R1769 VPB.n885 VPB 0.068
R1770 VPB.n894 VPB 0.068
R1771 a_14511_943.n2 a_14511_943.t6 475.572
R1772 a_14511_943.n1 a_14511_943.t7 469.145
R1773 a_14511_943.n6 a_14511_943.t8 454.685
R1774 a_14511_943.n6 a_14511_943.t13 428.979
R1775 a_14511_943.n2 a_14511_943.t10 384.527
R1776 a_14511_943.n1 a_14511_943.t9 384.527
R1777 a_14511_943.n3 a_14511_943.t12 277.772
R1778 a_14511_943.n5 a_14511_943.t11 251.219
R1779 a_14511_943.n7 a_14511_943.t5 248.006
R1780 a_14511_943.n13 a_14511_943.n12 220.639
R1781 a_14511_943.n4 a_14511_943.n3 156.851
R1782 a_14511_943.n14 a_14511_943.n13 135.994
R1783 a_14511_943.n7 a_14511_943.n6 81.941
R1784 a_14511_943.n8 a_14511_943.n7 78.947
R1785 a_14511_943.n8 a_14511_943.n5 77.859
R1786 a_14511_943.n15 a_14511_943.n14 76.001
R1787 a_14511_943.n13 a_14511_943.n8 76
R1788 a_14511_943.n3 a_14511_943.n2 67.889
R1789 a_14511_943.n4 a_14511_943.n1 66.88
R1790 a_14511_943.n12 a_14511_943.n11 30
R1791 a_14511_943.n5 a_14511_943.n4 26.552
R1792 a_14511_943.n10 a_14511_943.n9 24.383
R1793 a_14511_943.n12 a_14511_943.n10 23.684
R1794 a_14511_943.n0 a_14511_943.t2 14.282
R1795 a_14511_943.n0 a_14511_943.t1 14.282
R1796 a_14511_943.n15 a_14511_943.t3 14.282
R1797 a_14511_943.t4 a_14511_943.n15 14.282
R1798 a_14511_943.n14 a_14511_943.n0 12.85
R1799 a_9331_943.n9 a_9331_943.t19 512.525
R1800 a_9331_943.n4 a_9331_943.t32 512.525
R1801 a_9331_943.n12 a_9331_943.t4 480.392
R1802 a_9331_943.n5 a_9331_943.t34 477.179
R1803 a_9331_943.n24 a_9331_943.t28 454.685
R1804 a_9331_943.n33 a_9331_943.t33 454.685
R1805 a_9331_943.n24 a_9331_943.t26 428.979
R1806 a_9331_943.n33 a_9331_943.t21 428.979
R1807 a_9331_943.n5 a_9331_943.t30 406.485
R1808 a_9331_943.n12 a_9331_943.t6 403.272
R1809 a_9331_943.n9 a_9331_943.t27 371.139
R1810 a_9331_943.n4 a_9331_943.t23 371.139
R1811 a_9331_943.n6 a_9331_943.t31 346.633
R1812 a_9331_943.n10 a_9331_943.t20 271.162
R1813 a_9331_943.n13 a_9331_943.t29 266.974
R1814 a_9331_943.n8 a_9331_943.t24 260.547
R1815 a_9331_943.n25 a_9331_943.t22 221.453
R1816 a_9331_943.n34 a_9331_943.t25 221.453
R1817 a_9331_943.n32 a_9331_943.n31 209.609
R1818 a_9331_943.n23 a_9331_943.n22 196.598
R1819 a_9331_943.n42 a_9331_943.n40 194.086
R1820 a_9331_943.n23 a_9331_943.n18 180.846
R1821 a_9331_943.n10 a_9331_943.n9 172.76
R1822 a_9331_943.n32 a_9331_943.n28 162.547
R1823 a_9331_943.n40 a_9331_943.n3 162.547
R1824 a_9331_943.n7 a_9331_943.n6 154.675
R1825 a_9331_943.n13 a_9331_943.n12 108.494
R1826 a_9331_943.n25 a_9331_943.n24 108.494
R1827 a_9331_943.n34 a_9331_943.n33 108.494
R1828 a_9331_943.n7 a_9331_943.n4 89.615
R1829 a_9331_943.n11 a_9331_943.n8 85.204
R1830 a_9331_943.n8 a_9331_943.n7 79.658
R1831 a_9331_943.n17 a_9331_943.n16 79.232
R1832 a_9331_943.n35 a_9331_943.n34 78.947
R1833 a_9331_943.n3 a_9331_943.n2 76.002
R1834 a_9331_943.n28 a_9331_943.n27 76.002
R1835 a_9331_943.n35 a_9331_943.n32 76
R1836 a_9331_943.n36 a_9331_943.n25 76
R1837 a_9331_943.n37 a_9331_943.n23 76
R1838 a_9331_943.n38 a_9331_943.n13 76
R1839 a_9331_943.n11 a_9331_943.n10 76
R1840 a_9331_943.n40 a_9331_943.n39 76
R1841 a_9331_943.n18 a_9331_943.n17 63.152
R1842 a_9331_943.n22 a_9331_943.n21 30
R1843 a_9331_943.n42 a_9331_943.n41 30
R1844 a_9331_943.n6 a_9331_943.n5 29.194
R1845 a_9331_943.n20 a_9331_943.n19 24.383
R1846 a_9331_943.n43 a_9331_943.n0 24.383
R1847 a_9331_943.n22 a_9331_943.n20 23.684
R1848 a_9331_943.n43 a_9331_943.n42 23.684
R1849 a_9331_943.n31 a_9331_943.n29 22.578
R1850 a_9331_943.n18 a_9331_943.n14 16.08
R1851 a_9331_943.n17 a_9331_943.n15 16.08
R1852 a_9331_943.n14 a_9331_943.t17 14.282
R1853 a_9331_943.n14 a_9331_943.t16 14.282
R1854 a_9331_943.n15 a_9331_943.t2 14.282
R1855 a_9331_943.n15 a_9331_943.t3 14.282
R1856 a_9331_943.n16 a_9331_943.t12 14.282
R1857 a_9331_943.n16 a_9331_943.t14 14.282
R1858 a_9331_943.n26 a_9331_943.t0 14.282
R1859 a_9331_943.n26 a_9331_943.t15 14.282
R1860 a_9331_943.n27 a_9331_943.t11 14.282
R1861 a_9331_943.n27 a_9331_943.t1 14.282
R1862 a_9331_943.n1 a_9331_943.t9 14.282
R1863 a_9331_943.n1 a_9331_943.t8 14.282
R1864 a_9331_943.n2 a_9331_943.t5 14.282
R1865 a_9331_943.n2 a_9331_943.t7 14.282
R1866 a_9331_943.n28 a_9331_943.n26 12.85
R1867 a_9331_943.n3 a_9331_943.n1 12.85
R1868 a_9331_943.n31 a_9331_943.n30 8.58
R1869 a_9331_943.n37 a_9331_943.n36 4.035
R1870 a_9331_943.n36 a_9331_943.n35 2.947
R1871 a_9331_943.n38 a_9331_943.n37 1.315
R1872 a_9331_943.n39 a_9331_943.n11 1.315
R1873 a_9331_943.n39 a_9331_943.n38 1.043
R1874 a_5327_159.n10 a_5327_159.t10 512.525
R1875 a_5327_159.n8 a_5327_159.t15 472.359
R1876 a_5327_159.n6 a_5327_159.t12 472.359
R1877 a_5327_159.n8 a_5327_159.t11 384.527
R1878 a_5327_159.n6 a_5327_159.t8 384.527
R1879 a_5327_159.n10 a_5327_159.t13 371.139
R1880 a_5327_159.n11 a_5327_159.t14 324.268
R1881 a_5327_159.n9 a_5327_159.t9 277.772
R1882 a_5327_159.n7 a_5327_159.t7 277.772
R1883 a_5327_159.n16 a_5327_159.n14 249.704
R1884 a_5327_159.n14 a_5327_159.n5 127.74
R1885 a_5327_159.n11 a_5327_159.n10 119.654
R1886 a_5327_159.n12 a_5327_159.n11 83.572
R1887 a_5327_159.n13 a_5327_159.n7 81.396
R1888 a_5327_159.n4 a_5327_159.n3 79.232
R1889 a_5327_159.n12 a_5327_159.n9 76
R1890 a_5327_159.n14 a_5327_159.n13 76
R1891 a_5327_159.n9 a_5327_159.n8 67.001
R1892 a_5327_159.n7 a_5327_159.n6 67.001
R1893 a_5327_159.n5 a_5327_159.n4 63.152
R1894 a_5327_159.n16 a_5327_159.n15 30
R1895 a_5327_159.n17 a_5327_159.n0 24.383
R1896 a_5327_159.n17 a_5327_159.n16 23.684
R1897 a_5327_159.n5 a_5327_159.n1 16.08
R1898 a_5327_159.n4 a_5327_159.n2 16.08
R1899 a_5327_159.n1 a_5327_159.t3 14.282
R1900 a_5327_159.n1 a_5327_159.t4 14.282
R1901 a_5327_159.n2 a_5327_159.t1 14.282
R1902 a_5327_159.n2 a_5327_159.t2 14.282
R1903 a_5327_159.n3 a_5327_159.t0 14.282
R1904 a_5327_159.n3 a_5327_159.t6 14.282
R1905 a_5327_159.n13 a_5327_159.n12 4.035
R1906 a_9806_73.n10 a_9806_73.n9 93.333
R1907 a_9806_73.n2 a_9806_73.n1 41.622
R1908 a_9806_73.n13 a_9806_73.n12 26.667
R1909 a_9806_73.n6 a_9806_73.n5 24.977
R1910 a_9806_73.t0 a_9806_73.n2 21.209
R1911 a_9806_73.t0 a_9806_73.n3 11.595
R1912 a_9806_73.t1 a_9806_73.n8 8.137
R1913 a_9806_73.t0 a_9806_73.n0 6.109
R1914 a_9806_73.t1 a_9806_73.n7 4.864
R1915 a_9806_73.t0 a_9806_73.n4 3.871
R1916 a_9806_73.t0 a_9806_73.n13 2.535
R1917 a_9806_73.n13 a_9806_73.t1 1.145
R1918 a_9806_73.n7 a_9806_73.n6 1.13
R1919 a_9806_73.t1 a_9806_73.n11 0.804
R1920 a_9806_73.n11 a_9806_73.n10 0.136
R1921 a_6233_75.n4 a_6233_75.n3 19.724
R1922 a_6233_75.t0 a_6233_75.n5 11.595
R1923 a_6233_75.t0 a_6233_75.n4 9.207
R1924 a_6233_75.n2 a_6233_75.n0 8.543
R1925 a_6233_75.t0 a_6233_75.n2 3.034
R1926 a_6233_75.n2 a_6233_75.n1 0.443
R1927 a_6514_182.n12 a_6514_182.n10 82.852
R1928 a_6514_182.n13 a_6514_182.n0 49.6
R1929 a_6514_182.t1 a_6514_182.n2 46.91
R1930 a_6514_182.n7 a_6514_182.n5 34.805
R1931 a_6514_182.n7 a_6514_182.n6 32.622
R1932 a_6514_182.n10 a_6514_182.t1 32.416
R1933 a_6514_182.n12 a_6514_182.n11 27.2
R1934 a_6514_182.n13 a_6514_182.n12 22.4
R1935 a_6514_182.n9 a_6514_182.n7 19.017
R1936 a_6514_182.n2 a_6514_182.n1 17.006
R1937 a_6514_182.n5 a_6514_182.n4 7.5
R1938 a_6514_182.n9 a_6514_182.n8 7.5
R1939 a_6514_182.t1 a_6514_182.n3 7.04
R1940 a_6514_182.n10 a_6514_182.n9 1.435
R1941 a_5779_943.n5 a_5779_943.t10 480.392
R1942 a_5779_943.n7 a_5779_943.t7 454.685
R1943 a_5779_943.n7 a_5779_943.t9 428.979
R1944 a_5779_943.n5 a_5779_943.t8 403.272
R1945 a_5779_943.n6 a_5779_943.t12 266.974
R1946 a_5779_943.n8 a_5779_943.t11 221.453
R1947 a_5779_943.n12 a_5779_943.n10 203.12
R1948 a_5779_943.n10 a_5779_943.n4 180.846
R1949 a_5779_943.n8 a_5779_943.n7 108.494
R1950 a_5779_943.n6 a_5779_943.n5 108.494
R1951 a_5779_943.n9 a_5779_943.n8 80.035
R1952 a_5779_943.n3 a_5779_943.n2 79.232
R1953 a_5779_943.n9 a_5779_943.n6 77.315
R1954 a_5779_943.n10 a_5779_943.n9 76
R1955 a_5779_943.n4 a_5779_943.n3 63.152
R1956 a_5779_943.n4 a_5779_943.n0 16.08
R1957 a_5779_943.n3 a_5779_943.n1 16.08
R1958 a_5779_943.n12 a_5779_943.n11 15.218
R1959 a_5779_943.n0 a_5779_943.t5 14.282
R1960 a_5779_943.n0 a_5779_943.t4 14.282
R1961 a_5779_943.n1 a_5779_943.t3 14.282
R1962 a_5779_943.n1 a_5779_943.t2 14.282
R1963 a_5779_943.n2 a_5779_943.t0 14.282
R1964 a_5779_943.n2 a_5779_943.t1 14.282
R1965 a_5779_943.n13 a_5779_943.n12 12.014
R1966 a_5457_1004.n8 a_5457_1004.t8 512.525
R1967 a_5457_1004.n6 a_5457_1004.t7 512.525
R1968 a_5457_1004.n8 a_5457_1004.t10 371.139
R1969 a_5457_1004.n6 a_5457_1004.t9 371.139
R1970 a_5457_1004.n9 a_5457_1004.t12 297.715
R1971 a_5457_1004.n7 a_5457_1004.t11 297.715
R1972 a_5457_1004.n13 a_5457_1004.n11 223.151
R1973 a_5457_1004.n11 a_5457_1004.n5 154.293
R1974 a_5457_1004.n9 a_5457_1004.n8 146.207
R1975 a_5457_1004.n7 a_5457_1004.n6 146.207
R1976 a_5457_1004.n10 a_5457_1004.n7 85.476
R1977 a_5457_1004.n4 a_5457_1004.n3 79.232
R1978 a_5457_1004.n11 a_5457_1004.n10 77.315
R1979 a_5457_1004.n10 a_5457_1004.n9 76
R1980 a_5457_1004.n5 a_5457_1004.n4 63.152
R1981 a_5457_1004.n13 a_5457_1004.n12 30
R1982 a_5457_1004.n14 a_5457_1004.n0 24.383
R1983 a_5457_1004.n14 a_5457_1004.n13 23.684
R1984 a_5457_1004.n5 a_5457_1004.n1 16.08
R1985 a_5457_1004.n4 a_5457_1004.n2 16.08
R1986 a_5457_1004.n1 a_5457_1004.t4 14.282
R1987 a_5457_1004.n1 a_5457_1004.t5 14.282
R1988 a_5457_1004.n2 a_5457_1004.t3 14.282
R1989 a_5457_1004.n2 a_5457_1004.t2 14.282
R1990 a_5457_1004.n3 a_5457_1004.t1 14.282
R1991 a_5457_1004.n3 a_5457_1004.t0 14.282
R1992 a_147_159.n17 a_147_159.t14 512.525
R1993 a_147_159.n2 a_147_159.t23 480.392
R1994 a_147_159.n15 a_147_159.t17 472.359
R1995 a_147_159.n0 a_147_159.t25 472.359
R1996 a_147_159.n2 a_147_159.t16 403.272
R1997 a_147_159.n15 a_147_159.t22 384.527
R1998 a_147_159.n0 a_147_159.t18 384.527
R1999 a_147_159.n17 a_147_159.t19 371.139
R2000 a_147_159.n18 a_147_159.t24 324.268
R2001 a_147_159.n3 a_147_159.t15 320.08
R2002 a_147_159.n16 a_147_159.t21 277.772
R2003 a_147_159.n1 a_147_159.t20 277.772
R2004 a_147_159.n13 a_147_159.n12 265.227
R2005 a_147_159.n25 a_147_159.n24 249.704
R2006 a_147_159.n13 a_147_159.n9 127.74
R2007 a_147_159.n29 a_147_159.n25 127.74
R2008 a_147_159.n18 a_147_159.n17 119.654
R2009 a_147_159.n19 a_147_159.n18 83.572
R2010 a_147_159.n8 a_147_159.n7 79.232
R2011 a_147_159.n28 a_147_159.n27 79.232
R2012 a_147_159.n4 a_147_159.n1 76.499
R2013 a_147_159.n19 a_147_159.n16 76
R2014 a_147_159.n4 a_147_159.n3 76
R2015 a_147_159.n14 a_147_159.n13 76
R2016 a_147_159.n25 a_147_159.n20 76
R2017 a_147_159.n16 a_147_159.n15 67.001
R2018 a_147_159.n1 a_147_159.n0 67.001
R2019 a_147_159.n9 a_147_159.n8 63.152
R2020 a_147_159.n29 a_147_159.n28 63.152
R2021 a_147_159.n3 a_147_159.n2 55.388
R2022 a_147_159.n24 a_147_159.n23 30
R2023 a_147_159.n22 a_147_159.n21 24.383
R2024 a_147_159.n24 a_147_159.n22 23.684
R2025 a_147_159.n12 a_147_159.n11 22.578
R2026 a_147_159.n28 a_147_159.n26 16.08
R2027 a_147_159.n9 a_147_159.n5 16.08
R2028 a_147_159.n8 a_147_159.n6 16.08
R2029 a_147_159.n30 a_147_159.n29 16.078
R2030 a_147_159.n26 a_147_159.t6 14.282
R2031 a_147_159.n26 a_147_159.t7 14.282
R2032 a_147_159.n27 a_147_159.t4 14.282
R2033 a_147_159.n27 a_147_159.t5 14.282
R2034 a_147_159.n5 a_147_159.t0 14.282
R2035 a_147_159.n5 a_147_159.t8 14.282
R2036 a_147_159.n6 a_147_159.t11 14.282
R2037 a_147_159.n6 a_147_159.t10 14.282
R2038 a_147_159.n7 a_147_159.t1 14.282
R2039 a_147_159.n7 a_147_159.t2 14.282
R2040 a_147_159.n30 a_147_159.t9 14.282
R2041 a_147_159.t12 a_147_159.n30 14.282
R2042 a_147_159.n12 a_147_159.n10 8.58
R2043 a_147_159.n20 a_147_159.n19 4.035
R2044 a_147_159.n20 a_147_159.n14 3.491
R2045 a_147_159.n14 a_147_159.n4 1.315
R2046 a_277_1004.n7 a_277_1004.t10 512.525
R2047 a_277_1004.n5 a_277_1004.t8 512.525
R2048 a_277_1004.n7 a_277_1004.t12 371.139
R2049 a_277_1004.n5 a_277_1004.t11 371.139
R2050 a_277_1004.n8 a_277_1004.t9 297.715
R2051 a_277_1004.n6 a_277_1004.t7 297.715
R2052 a_277_1004.n12 a_277_1004.n10 229.673
R2053 a_277_1004.n10 a_277_1004.n4 154.293
R2054 a_277_1004.n8 a_277_1004.n7 146.207
R2055 a_277_1004.n6 a_277_1004.n5 146.207
R2056 a_277_1004.n9 a_277_1004.n6 85.476
R2057 a_277_1004.n3 a_277_1004.n2 79.232
R2058 a_277_1004.n10 a_277_1004.n9 77.315
R2059 a_277_1004.n9 a_277_1004.n8 76
R2060 a_277_1004.n4 a_277_1004.n3 63.152
R2061 a_277_1004.n4 a_277_1004.n0 16.08
R2062 a_277_1004.n3 a_277_1004.n1 16.08
R2063 a_277_1004.n12 a_277_1004.n11 15.218
R2064 a_277_1004.n0 a_277_1004.t4 14.282
R2065 a_277_1004.n0 a_277_1004.t0 14.282
R2066 a_277_1004.n1 a_277_1004.t3 14.282
R2067 a_277_1004.n1 a_277_1004.t2 14.282
R2068 a_277_1004.n2 a_277_1004.t6 14.282
R2069 a_277_1004.n2 a_277_1004.t5 14.282
R2070 a_277_1004.n13 a_277_1004.n12 12.014
R2071 a_4151_943.n2 a_4151_943.t13 512.525
R2072 a_4151_943.n1 a_4151_943.t10 512.525
R2073 a_4151_943.n6 a_4151_943.t7 454.685
R2074 a_4151_943.n6 a_4151_943.t11 428.979
R2075 a_4151_943.n2 a_4151_943.t8 371.139
R2076 a_4151_943.n1 a_4151_943.t5 371.139
R2077 a_4151_943.n3 a_4151_943.n2 258.98
R2078 a_4151_943.n5 a_4151_943.n1 195.827
R2079 a_4151_943.n14 a_4151_943.n13 189.099
R2080 a_4151_943.n7 a_4151_943.t12 183.653
R2081 a_4151_943.n3 a_4151_943.t9 176.995
R2082 a_4151_943.n4 a_4151_943.t6 170.569
R2083 a_4151_943.n13 a_4151_943.n12 167.533
R2084 a_4151_943.n4 a_4151_943.n3 153.043
R2085 a_4151_943.n7 a_4151_943.n6 135.047
R2086 a_4151_943.n8 a_4151_943.n5 118.94
R2087 a_4151_943.n8 a_4151_943.n7 78.947
R2088 a_4151_943.n15 a_4151_943.n14 76.001
R2089 a_4151_943.n13 a_4151_943.n8 76
R2090 a_4151_943.n5 a_4151_943.n4 63.152
R2091 a_4151_943.n12 a_4151_943.n11 30
R2092 a_4151_943.n10 a_4151_943.n9 24.383
R2093 a_4151_943.n12 a_4151_943.n10 23.684
R2094 a_4151_943.n0 a_4151_943.t0 14.282
R2095 a_4151_943.n0 a_4151_943.t2 14.282
R2096 a_4151_943.n15 a_4151_943.t1 14.282
R2097 a_4151_943.t3 a_4151_943.n15 14.282
R2098 a_4151_943.n14 a_4151_943.n0 12.85
R2099 a_16421_1005.n4 a_16421_1005.n3 196.002
R2100 a_16421_1005.t0 a_16421_1005.n5 89.556
R2101 a_16421_1005.n3 a_16421_1005.n2 75.271
R2102 a_16421_1005.n5 a_16421_1005.n4 75.214
R2103 a_16421_1005.n3 a_16421_1005.n1 36.52
R2104 a_16421_1005.n4 a_16421_1005.t6 14.338
R2105 a_16421_1005.n1 a_16421_1005.t7 14.282
R2106 a_16421_1005.n1 a_16421_1005.t4 14.282
R2107 a_16421_1005.n2 a_16421_1005.t2 14.282
R2108 a_16421_1005.n2 a_16421_1005.t3 14.282
R2109 a_16421_1005.n0 a_16421_1005.t1 14.282
R2110 a_16421_1005.n0 a_16421_1005.t5 14.282
R2111 a_16421_1005.n5 a_16421_1005.n0 12.119
R2112 a_15757_1005.n4 a_15757_1005.n3 195.987
R2113 a_15757_1005.n2 a_15757_1005.t7 89.553
R2114 a_15757_1005.n4 a_15757_1005.n0 75.271
R2115 a_15757_1005.n3 a_15757_1005.n2 75.214
R2116 a_15757_1005.n5 a_15757_1005.n4 36.517
R2117 a_15757_1005.n3 a_15757_1005.t5 14.338
R2118 a_15757_1005.n1 a_15757_1005.t6 14.282
R2119 a_15757_1005.n1 a_15757_1005.t4 14.282
R2120 a_15757_1005.n0 a_15757_1005.t2 14.282
R2121 a_15757_1005.n0 a_15757_1005.t3 14.282
R2122 a_15757_1005.t1 a_15757_1005.n5 14.282
R2123 a_15757_1005.n5 a_15757_1005.t0 14.282
R2124 a_15757_1005.n2 a_15757_1005.n1 12.119
R2125 a_10637_1004.n8 a_10637_1004.t12 512.525
R2126 a_10637_1004.n6 a_10637_1004.t11 512.525
R2127 a_10637_1004.n8 a_10637_1004.t8 371.139
R2128 a_10637_1004.n6 a_10637_1004.t7 371.139
R2129 a_10637_1004.n9 a_10637_1004.t10 297.715
R2130 a_10637_1004.n7 a_10637_1004.t9 297.715
R2131 a_10637_1004.n13 a_10637_1004.n11 223.151
R2132 a_10637_1004.n11 a_10637_1004.n5 154.293
R2133 a_10637_1004.n9 a_10637_1004.n8 146.207
R2134 a_10637_1004.n7 a_10637_1004.n6 146.207
R2135 a_10637_1004.n10 a_10637_1004.n7 85.476
R2136 a_10637_1004.n4 a_10637_1004.n3 79.232
R2137 a_10637_1004.n11 a_10637_1004.n10 77.315
R2138 a_10637_1004.n10 a_10637_1004.n9 76
R2139 a_10637_1004.n5 a_10637_1004.n4 63.152
R2140 a_10637_1004.n13 a_10637_1004.n12 30
R2141 a_10637_1004.n14 a_10637_1004.n0 24.383
R2142 a_10637_1004.n14 a_10637_1004.n13 23.684
R2143 a_10637_1004.n5 a_10637_1004.n1 16.08
R2144 a_10637_1004.n4 a_10637_1004.n2 16.08
R2145 a_10637_1004.n1 a_10637_1004.t2 14.282
R2146 a_10637_1004.n1 a_10637_1004.t1 14.282
R2147 a_10637_1004.n2 a_10637_1004.t6 14.282
R2148 a_10637_1004.n2 a_10637_1004.t5 14.282
R2149 a_10637_1004.n3 a_10637_1004.t4 14.282
R2150 a_10637_1004.n3 a_10637_1004.t3 14.282
R2151 a_14284_182.n9 a_14284_182.n7 82.852
R2152 a_14284_182.n3 a_14284_182.n1 44.628
R2153 a_14284_182.t0 a_14284_182.n9 32.417
R2154 a_14284_182.n7 a_14284_182.n6 27.2
R2155 a_14284_182.n5 a_14284_182.n4 23.498
R2156 a_14284_182.n3 a_14284_182.n2 23.284
R2157 a_14284_182.n7 a_14284_182.n5 22.4
R2158 a_14284_182.t0 a_14284_182.n11 20.241
R2159 a_14284_182.n11 a_14284_182.n10 13.494
R2160 a_14284_182.t0 a_14284_182.n0 8.137
R2161 a_14284_182.t0 a_14284_182.n3 5.727
R2162 a_14284_182.n9 a_14284_182.n8 1.435
R2163 a_13041_75.t0 a_13041_75.n3 117.777
R2164 a_13041_75.n6 a_13041_75.n5 45.444
R2165 a_13041_75.t0 a_13041_75.n6 21.213
R2166 a_13041_75.t0 a_13041_75.n4 11.595
R2167 a_13041_75.n2 a_13041_75.n0 8.543
R2168 a_13041_75.t0 a_13041_75.n2 3.034
R2169 a_13041_75.n2 a_13041_75.n1 0.443
R2170 VNB VNB.n1451 300.778
R2171 VNB.n170 VNB.n169 199.897
R2172 VNB.n229 VNB.n228 199.897
R2173 VNB.n288 VNB.n287 199.897
R2174 VNB.n347 VNB.n346 199.897
R2175 VNB.n406 VNB.n405 199.897
R2176 VNB.n481 VNB.n480 199.897
R2177 VNB.n549 VNB.n548 199.897
R2178 VNB.n608 VNB.n607 199.897
R2179 VNB.n683 VNB.n682 199.897
R2180 VNB.n758 VNB.n757 199.897
R2181 VNB.n74 VNB.n73 199.897
R2182 VNB.n837 VNB.n836 199.897
R2183 VNB.n905 VNB.n904 199.897
R2184 VNB.n964 VNB.n963 199.897
R2185 VNB.n1032 VNB.n1031 199.897
R2186 VNB.n1107 VNB.n1106 199.897
R2187 VNB.n1166 VNB.n1165 199.897
R2188 VNB.n1241 VNB.n1240 199.897
R2189 VNB.n1309 VNB.n1308 199.897
R2190 VNB.n1361 VNB.n1360 199.897
R2191 VNB.n18 VNB.n17 199.897
R2192 VNB.n238 VNB.n236 154.509
R2193 VNB.n179 VNB.n177 154.509
R2194 VNB.n356 VNB.n354 154.509
R2195 VNB.n297 VNB.n295 154.509
R2196 VNB.n490 VNB.n488 154.509
R2197 VNB.n415 VNB.n413 154.509
R2198 VNB.n617 VNB.n615 154.509
R2199 VNB.n558 VNB.n556 154.509
R2200 VNB.n767 VNB.n765 154.509
R2201 VNB.n692 VNB.n690 154.509
R2202 VNB.n846 VNB.n844 154.509
R2203 VNB.n89 VNB.n87 154.509
R2204 VNB.n973 VNB.n971 154.509
R2205 VNB.n914 VNB.n912 154.509
R2206 VNB.n1116 VNB.n1114 154.509
R2207 VNB.n1041 VNB.n1039 154.509
R2208 VNB.n1250 VNB.n1248 154.509
R2209 VNB.n1175 VNB.n1173 154.509
R2210 VNB.n1370 VNB.n1368 154.509
R2211 VNB.n1318 VNB.n1316 154.509
R2212 VNB.n27 VNB.n25 154.509
R2213 VNB.n447 VNB.n446 147.75
R2214 VNB.n649 VNB.n648 147.75
R2215 VNB.n724 VNB.n723 147.75
R2216 VNB.n804 VNB.n803 147.75
R2217 VNB.n1073 VNB.n1072 147.75
R2218 VNB.n1207 VNB.n1206 147.75
R2219 VNB.n1402 VNB.n1401 147.75
R2220 VNB.n51 VNB.n50 147.75
R2221 VNB.n195 VNB.n194 121.366
R2222 VNB.n254 VNB.n253 121.366
R2223 VNB.n313 VNB.n312 121.366
R2224 VNB.n372 VNB.n371 121.366
R2225 VNB.n459 VNB.n456 121.366
R2226 VNB.n574 VNB.n573 121.366
R2227 VNB.n661 VNB.n658 121.366
R2228 VNB.n736 VNB.n733 121.366
R2229 VNB.n815 VNB.n812 121.366
R2230 VNB.n930 VNB.n929 121.366
R2231 VNB.n1085 VNB.n1082 121.366
R2232 VNB.n1132 VNB.n1131 121.366
R2233 VNB.n1219 VNB.n1216 121.366
R2234 VNB.n1414 VNB.n1411 121.366
R2235 VNB.n56 VNB.n54 121.366
R2236 VNB.n526 VNB.n525 85.559
R2237 VNB.n882 VNB.n881 85.559
R2238 VNB.n1009 VNB.n1008 85.559
R2239 VNB.n1286 VNB.n1285 85.559
R2240 VNB.n787 VNB.n786 84.842
R2241 VNB.n1338 VNB.n1337 84.842
R2242 VNB.n138 VNB.n129 76.136
R2243 VNB.n138 VNB.n137 76
R2244 VNB.n1438 VNB.n1437 76
R2245 VNB.n1425 VNB.n1424 76
R2246 VNB.n1421 VNB.n1420 76
R2247 VNB.n1417 VNB.n1416 76
R2248 VNB.n1405 VNB.n1404 76
R2249 VNB.n1400 VNB.n1399 76
R2250 VNB.n1396 VNB.n1395 76
R2251 VNB.n1392 VNB.n1391 76
R2252 VNB.n1388 VNB.n1387 76
R2253 VNB.n1384 VNB.n1383 76
R2254 VNB.n1380 VNB.n1379 76
R2255 VNB.n1376 VNB.n1375 76
R2256 VNB.n1372 VNB.n1371 76
R2257 VNB.n1350 VNB.n1349 76
R2258 VNB.n1346 VNB.n1345 76
R2259 VNB.n1342 VNB.n1341 76
R2260 VNB.n1336 VNB.n1335 76
R2261 VNB.n1332 VNB.n1331 76
R2262 VNB.n1328 VNB.n1327 76
R2263 VNB.n1324 VNB.n1323 76
R2264 VNB.n1320 VNB.n1319 76
R2265 VNB.n1298 VNB.n1297 76
R2266 VNB.n1294 VNB.n1293 76
R2267 VNB.n1290 VNB.n1289 76
R2268 VNB.n1284 VNB.n1283 76
R2269 VNB.n1280 VNB.n1279 76
R2270 VNB.n1276 VNB.n1275 76
R2271 VNB.n1272 VNB.n1271 76
R2272 VNB.n1268 VNB.n1267 76
R2273 VNB.n1264 VNB.n1263 76
R2274 VNB.n1260 VNB.n1259 76
R2275 VNB.n1256 VNB.n1255 76
R2276 VNB.n1252 VNB.n1251 76
R2277 VNB.n1230 VNB.n1229 76
R2278 VNB.n1226 VNB.n1225 76
R2279 VNB.n1222 VNB.n1221 76
R2280 VNB.n1210 VNB.n1209 76
R2281 VNB.n1205 VNB.n1204 76
R2282 VNB.n1201 VNB.n1200 76
R2283 VNB.n1197 VNB.n1196 76
R2284 VNB.n1193 VNB.n1192 76
R2285 VNB.n1189 VNB.n1188 76
R2286 VNB.n1185 VNB.n1184 76
R2287 VNB.n1181 VNB.n1180 76
R2288 VNB.n1177 VNB.n1176 76
R2289 VNB.n1155 VNB.n1154 76
R2290 VNB.n1151 VNB.n1150 76
R2291 VNB.n1147 VNB.n1146 76
R2292 VNB.n1136 VNB.n1135 76
R2293 VNB.n1130 VNB.n1129 76
R2294 VNB.n1126 VNB.n1125 76
R2295 VNB.n1122 VNB.n1121 76
R2296 VNB.n1118 VNB.n1117 76
R2297 VNB.n1096 VNB.n1095 76
R2298 VNB.n1092 VNB.n1091 76
R2299 VNB.n1088 VNB.n1087 76
R2300 VNB.n1076 VNB.n1075 76
R2301 VNB.n1071 VNB.n1070 76
R2302 VNB.n1067 VNB.n1066 76
R2303 VNB.n1063 VNB.n1062 76
R2304 VNB.n1059 VNB.n1058 76
R2305 VNB.n1055 VNB.n1054 76
R2306 VNB.n1051 VNB.n1050 76
R2307 VNB.n1047 VNB.n1046 76
R2308 VNB.n1043 VNB.n1042 76
R2309 VNB.n1021 VNB.n1020 76
R2310 VNB.n1017 VNB.n1016 76
R2311 VNB.n1013 VNB.n1012 76
R2312 VNB.n1007 VNB.n1006 76
R2313 VNB.n1003 VNB.n1002 76
R2314 VNB.n999 VNB.n998 76
R2315 VNB.n995 VNB.n994 76
R2316 VNB.n991 VNB.n990 76
R2317 VNB.n987 VNB.n986 76
R2318 VNB.n983 VNB.n982 76
R2319 VNB.n979 VNB.n978 76
R2320 VNB.n975 VNB.n974 76
R2321 VNB.n953 VNB.n952 76
R2322 VNB.n949 VNB.n948 76
R2323 VNB.n945 VNB.n944 76
R2324 VNB.n934 VNB.n933 76
R2325 VNB.n928 VNB.n927 76
R2326 VNB.n924 VNB.n923 76
R2327 VNB.n920 VNB.n919 76
R2328 VNB.n916 VNB.n915 76
R2329 VNB.n894 VNB.n893 76
R2330 VNB.n890 VNB.n889 76
R2331 VNB.n886 VNB.n885 76
R2332 VNB.n880 VNB.n879 76
R2333 VNB.n876 VNB.n875 76
R2334 VNB.n872 VNB.n871 76
R2335 VNB.n868 VNB.n867 76
R2336 VNB.n864 VNB.n863 76
R2337 VNB.n860 VNB.n859 76
R2338 VNB.n856 VNB.n855 76
R2339 VNB.n852 VNB.n851 76
R2340 VNB.n848 VNB.n847 76
R2341 VNB.n826 VNB.n825 76
R2342 VNB.n822 VNB.n821 76
R2343 VNB.n818 VNB.n817 76
R2344 VNB.n806 VNB.n802 76
R2345 VNB.n791 VNB.n790 76
R2346 VNB.n785 VNB.n784 76
R2347 VNB.n781 VNB.n780 76
R2348 VNB.n777 VNB.n776 76
R2349 VNB.n773 VNB.n772 76
R2350 VNB.n769 VNB.n768 76
R2351 VNB.n747 VNB.n746 76
R2352 VNB.n743 VNB.n742 76
R2353 VNB.n739 VNB.n738 76
R2354 VNB.n727 VNB.n726 76
R2355 VNB.n722 VNB.n721 76
R2356 VNB.n718 VNB.n717 76
R2357 VNB.n714 VNB.n713 76
R2358 VNB.n710 VNB.n709 76
R2359 VNB.n706 VNB.n705 76
R2360 VNB.n702 VNB.n701 76
R2361 VNB.n698 VNB.n697 76
R2362 VNB.n694 VNB.n693 76
R2363 VNB.n672 VNB.n671 76
R2364 VNB.n668 VNB.n667 76
R2365 VNB.n664 VNB.n663 76
R2366 VNB.n652 VNB.n651 76
R2367 VNB.n647 VNB.n646 76
R2368 VNB.n643 VNB.n642 76
R2369 VNB.n639 VNB.n638 76
R2370 VNB.n635 VNB.n634 76
R2371 VNB.n631 VNB.n630 76
R2372 VNB.n627 VNB.n626 76
R2373 VNB.n623 VNB.n622 76
R2374 VNB.n619 VNB.n618 76
R2375 VNB.n597 VNB.n596 76
R2376 VNB.n593 VNB.n592 76
R2377 VNB.n589 VNB.n588 76
R2378 VNB.n578 VNB.n577 76
R2379 VNB.n572 VNB.n571 76
R2380 VNB.n568 VNB.n567 76
R2381 VNB.n564 VNB.n563 76
R2382 VNB.n560 VNB.n559 76
R2383 VNB.n538 VNB.n537 76
R2384 VNB.n534 VNB.n533 76
R2385 VNB.n530 VNB.n529 76
R2386 VNB.n524 VNB.n523 76
R2387 VNB.n520 VNB.n519 76
R2388 VNB.n516 VNB.n515 76
R2389 VNB.n512 VNB.n511 76
R2390 VNB.n508 VNB.n507 76
R2391 VNB.n504 VNB.n503 76
R2392 VNB.n500 VNB.n499 76
R2393 VNB.n496 VNB.n495 76
R2394 VNB.n492 VNB.n491 76
R2395 VNB.n470 VNB.n469 76
R2396 VNB.n466 VNB.n465 76
R2397 VNB.n462 VNB.n461 76
R2398 VNB.n450 VNB.n449 76
R2399 VNB.n445 VNB.n444 76
R2400 VNB.n441 VNB.n440 76
R2401 VNB.n437 VNB.n436 76
R2402 VNB.n433 VNB.n432 76
R2403 VNB.n429 VNB.n428 76
R2404 VNB.n425 VNB.n424 76
R2405 VNB.n421 VNB.n420 76
R2406 VNB.n417 VNB.n416 76
R2407 VNB.n395 VNB.n394 76
R2408 VNB.n391 VNB.n390 76
R2409 VNB.n387 VNB.n386 76
R2410 VNB.n376 VNB.n375 76
R2411 VNB.n370 VNB.n369 76
R2412 VNB.n366 VNB.n365 76
R2413 VNB.n362 VNB.n361 76
R2414 VNB.n358 VNB.n357 76
R2415 VNB.n336 VNB.n335 76
R2416 VNB.n332 VNB.n331 76
R2417 VNB.n328 VNB.n327 76
R2418 VNB.n317 VNB.n316 76
R2419 VNB.n311 VNB.n310 76
R2420 VNB.n307 VNB.n306 76
R2421 VNB.n303 VNB.n302 76
R2422 VNB.n299 VNB.n298 76
R2423 VNB.n277 VNB.n276 76
R2424 VNB.n273 VNB.n272 76
R2425 VNB.n269 VNB.n268 76
R2426 VNB.n258 VNB.n257 76
R2427 VNB.n252 VNB.n251 76
R2428 VNB.n248 VNB.n247 76
R2429 VNB.n244 VNB.n243 76
R2430 VNB.n240 VNB.n239 76
R2431 VNB.n218 VNB.n217 76
R2432 VNB.n214 VNB.n213 76
R2433 VNB.n210 VNB.n209 76
R2434 VNB.n199 VNB.n198 76
R2435 VNB.n193 VNB.n192 76
R2436 VNB.n189 VNB.n188 76
R2437 VNB.n185 VNB.n184 76
R2438 VNB.n181 VNB.n180 76
R2439 VNB.n159 VNB.n158 76
R2440 VNB.n155 VNB.n154 76
R2441 VNB.n147 VNB.n146 76
R2442 VNB.n61 VNB.n60 73.875
R2443 VNB.n455 VNB.n454 64.552
R2444 VNB.n657 VNB.n656 64.552
R2445 VNB.n732 VNB.n731 64.552
R2446 VNB.n811 VNB.n810 64.552
R2447 VNB.n1081 VNB.n1080 64.552
R2448 VNB.n1215 VNB.n1214 64.552
R2449 VNB.n1410 VNB.n1409 64.552
R2450 VNB.n59 VNB.n7 64.552
R2451 VNB.n204 VNB.n203 63.835
R2452 VNB.n263 VNB.n262 63.835
R2453 VNB.n322 VNB.n321 63.835
R2454 VNB.n381 VNB.n380 63.835
R2455 VNB.n583 VNB.n582 63.835
R2456 VNB.n939 VNB.n938 63.835
R2457 VNB.n1141 VNB.n1140 63.835
R2458 VNB.n145 VNB.n144 49.896
R2459 VNB.n528 VNB.n527 41.971
R2460 VNB.n884 VNB.n883 41.971
R2461 VNB.n1011 VNB.n1010 41.971
R2462 VNB.n1288 VNB.n1287 41.971
R2463 VNB.n196 VNB.n195 36.937
R2464 VNB.n255 VNB.n254 36.937
R2465 VNB.n314 VNB.n313 36.937
R2466 VNB.n373 VNB.n372 36.937
R2467 VNB.n459 VNB.n458 36.937
R2468 VNB.n575 VNB.n574 36.937
R2469 VNB.n661 VNB.n660 36.937
R2470 VNB.n736 VNB.n735 36.937
R2471 VNB.n815 VNB.n814 36.937
R2472 VNB.n931 VNB.n930 36.937
R2473 VNB.n1085 VNB.n1084 36.937
R2474 VNB.n1133 VNB.n1132 36.937
R2475 VNB.n1219 VNB.n1218 36.937
R2476 VNB.n1414 VNB.n1413 36.937
R2477 VNB.n56 VNB.n55 36.937
R2478 VNB.n789 VNB.n788 36.678
R2479 VNB.n1340 VNB.n1339 36.678
R2480 VNB.n133 VNB.n132 35.01
R2481 VNB.n458 VNB.n457 29.844
R2482 VNB.n660 VNB.n659 29.844
R2483 VNB.n735 VNB.n734 29.844
R2484 VNB.n814 VNB.n813 29.844
R2485 VNB.n1084 VNB.n1083 29.844
R2486 VNB.n1218 VNB.n1217 29.844
R2487 VNB.n1413 VNB.n1412 29.844
R2488 VNB.n131 VNB.n130 29.127
R2489 VNB.n203 VNB.n202 28.421
R2490 VNB.n262 VNB.n261 28.421
R2491 VNB.n321 VNB.n320 28.421
R2492 VNB.n380 VNB.n379 28.421
R2493 VNB.n454 VNB.n453 28.421
R2494 VNB.n582 VNB.n581 28.421
R2495 VNB.n656 VNB.n655 28.421
R2496 VNB.n731 VNB.n730 28.421
R2497 VNB.n810 VNB.n809 28.421
R2498 VNB.n938 VNB.n937 28.421
R2499 VNB.n1080 VNB.n1079 28.421
R2500 VNB.n1140 VNB.n1139 28.421
R2501 VNB.n1214 VNB.n1213 28.421
R2502 VNB.n1409 VNB.n1408 28.421
R2503 VNB.n7 VNB.n6 28.421
R2504 VNB.n207 VNB.n206 27.855
R2505 VNB.n266 VNB.n265 27.855
R2506 VNB.n325 VNB.n324 27.855
R2507 VNB.n384 VNB.n383 27.855
R2508 VNB.n586 VNB.n585 27.855
R2509 VNB.n942 VNB.n941 27.855
R2510 VNB.n1144 VNB.n1143 27.855
R2511 VNB.n203 VNB.n201 25.263
R2512 VNB.n262 VNB.n260 25.263
R2513 VNB.n321 VNB.n319 25.263
R2514 VNB.n380 VNB.n378 25.263
R2515 VNB.n454 VNB.n452 25.263
R2516 VNB.n582 VNB.n580 25.263
R2517 VNB.n656 VNB.n654 25.263
R2518 VNB.n731 VNB.n729 25.263
R2519 VNB.n810 VNB.n808 25.263
R2520 VNB.n938 VNB.n936 25.263
R2521 VNB.n1080 VNB.n1078 25.263
R2522 VNB.n1140 VNB.n1138 25.263
R2523 VNB.n1214 VNB.n1212 25.263
R2524 VNB.n1409 VNB.n1407 25.263
R2525 VNB.n7 VNB.n5 25.263
R2526 VNB.n201 VNB.n200 24.383
R2527 VNB.n260 VNB.n259 24.383
R2528 VNB.n319 VNB.n318 24.383
R2529 VNB.n378 VNB.n377 24.383
R2530 VNB.n452 VNB.n451 24.383
R2531 VNB.n580 VNB.n579 24.383
R2532 VNB.n654 VNB.n653 24.383
R2533 VNB.n729 VNB.n728 24.383
R2534 VNB.n808 VNB.n807 24.383
R2535 VNB.n936 VNB.n935 24.383
R2536 VNB.n1078 VNB.n1077 24.383
R2537 VNB.n1138 VNB.n1137 24.383
R2538 VNB.n1212 VNB.n1211 24.383
R2539 VNB.n1407 VNB.n1406 24.383
R2540 VNB.n5 VNB.n4 24.383
R2541 VNB.n141 VNB.t10 20.794
R2542 VNB.n129 VNB.n126 20.452
R2543 VNB.n1439 VNB.n1438 20.452
R2544 VNB.n134 VNB.n133 20.094
R2545 VNB.n143 VNB.n142 20.094
R2546 VNB.n151 VNB.n150 20.094
R2547 VNB.n133 VNB.n131 19.017
R2548 VNB.n208 VNB.n207 16.721
R2549 VNB.n267 VNB.n266 16.721
R2550 VNB.n326 VNB.n325 16.721
R2551 VNB.n385 VNB.n384 16.721
R2552 VNB.n587 VNB.n586 16.721
R2553 VNB.n943 VNB.n942 16.721
R2554 VNB.n1145 VNB.n1144 16.721
R2555 VNB.n137 VNB.n136 13.653
R2556 VNB.n136 VNB.n135 13.653
R2557 VNB.n146 VNB.n145 13.653
R2558 VNB.n154 VNB.n153 13.653
R2559 VNB.n153 VNB.n152 13.653
R2560 VNB.n158 VNB.n157 13.653
R2561 VNB.n157 VNB.n156 13.653
R2562 VNB.n180 VNB.n179 13.653
R2563 VNB.n179 VNB.n178 13.653
R2564 VNB.n184 VNB.n183 13.653
R2565 VNB.n183 VNB.n182 13.653
R2566 VNB.n188 VNB.n187 13.653
R2567 VNB.n187 VNB.n186 13.653
R2568 VNB.n192 VNB.n191 13.653
R2569 VNB.n191 VNB.n190 13.653
R2570 VNB.n198 VNB.n197 13.653
R2571 VNB.n197 VNB.n196 13.653
R2572 VNB.n209 VNB.n208 13.653
R2573 VNB.n213 VNB.n212 13.653
R2574 VNB.n212 VNB.n211 13.653
R2575 VNB.n217 VNB.n216 13.653
R2576 VNB.n216 VNB.n215 13.653
R2577 VNB.n239 VNB.n238 13.653
R2578 VNB.n238 VNB.n237 13.653
R2579 VNB.n243 VNB.n242 13.653
R2580 VNB.n242 VNB.n241 13.653
R2581 VNB.n247 VNB.n246 13.653
R2582 VNB.n246 VNB.n245 13.653
R2583 VNB.n251 VNB.n250 13.653
R2584 VNB.n250 VNB.n249 13.653
R2585 VNB.n257 VNB.n256 13.653
R2586 VNB.n256 VNB.n255 13.653
R2587 VNB.n268 VNB.n267 13.653
R2588 VNB.n272 VNB.n271 13.653
R2589 VNB.n271 VNB.n270 13.653
R2590 VNB.n276 VNB.n275 13.653
R2591 VNB.n275 VNB.n274 13.653
R2592 VNB.n298 VNB.n297 13.653
R2593 VNB.n297 VNB.n296 13.653
R2594 VNB.n302 VNB.n301 13.653
R2595 VNB.n301 VNB.n300 13.653
R2596 VNB.n306 VNB.n305 13.653
R2597 VNB.n305 VNB.n304 13.653
R2598 VNB.n310 VNB.n309 13.653
R2599 VNB.n309 VNB.n308 13.653
R2600 VNB.n316 VNB.n315 13.653
R2601 VNB.n315 VNB.n314 13.653
R2602 VNB.n327 VNB.n326 13.653
R2603 VNB.n331 VNB.n330 13.653
R2604 VNB.n330 VNB.n329 13.653
R2605 VNB.n335 VNB.n334 13.653
R2606 VNB.n334 VNB.n333 13.653
R2607 VNB.n357 VNB.n356 13.653
R2608 VNB.n356 VNB.n355 13.653
R2609 VNB.n361 VNB.n360 13.653
R2610 VNB.n360 VNB.n359 13.653
R2611 VNB.n365 VNB.n364 13.653
R2612 VNB.n364 VNB.n363 13.653
R2613 VNB.n369 VNB.n368 13.653
R2614 VNB.n368 VNB.n367 13.653
R2615 VNB.n375 VNB.n374 13.653
R2616 VNB.n374 VNB.n373 13.653
R2617 VNB.n386 VNB.n385 13.653
R2618 VNB.n390 VNB.n389 13.653
R2619 VNB.n389 VNB.n388 13.653
R2620 VNB.n394 VNB.n393 13.653
R2621 VNB.n393 VNB.n392 13.653
R2622 VNB.n416 VNB.n415 13.653
R2623 VNB.n415 VNB.n414 13.653
R2624 VNB.n420 VNB.n419 13.653
R2625 VNB.n419 VNB.n418 13.653
R2626 VNB.n424 VNB.n423 13.653
R2627 VNB.n423 VNB.n422 13.653
R2628 VNB.n428 VNB.n427 13.653
R2629 VNB.n427 VNB.n426 13.653
R2630 VNB.n432 VNB.n431 13.653
R2631 VNB.n431 VNB.n430 13.653
R2632 VNB.n436 VNB.n435 13.653
R2633 VNB.n435 VNB.n434 13.653
R2634 VNB.n440 VNB.n439 13.653
R2635 VNB.n439 VNB.n438 13.653
R2636 VNB.n444 VNB.n443 13.653
R2637 VNB.n443 VNB.n442 13.653
R2638 VNB.n449 VNB.n448 13.653
R2639 VNB.n448 VNB.n447 13.653
R2640 VNB.n461 VNB.n460 13.653
R2641 VNB.n460 VNB.n459 13.653
R2642 VNB.n465 VNB.n464 13.653
R2643 VNB.n464 VNB.n463 13.653
R2644 VNB.n469 VNB.n468 13.653
R2645 VNB.n468 VNB.n467 13.653
R2646 VNB.n491 VNB.n490 13.653
R2647 VNB.n490 VNB.n489 13.653
R2648 VNB.n495 VNB.n494 13.653
R2649 VNB.n494 VNB.n493 13.653
R2650 VNB.n499 VNB.n498 13.653
R2651 VNB.n498 VNB.n497 13.653
R2652 VNB.n503 VNB.n502 13.653
R2653 VNB.n502 VNB.n501 13.653
R2654 VNB.n507 VNB.n506 13.653
R2655 VNB.n506 VNB.n505 13.653
R2656 VNB.n511 VNB.n510 13.653
R2657 VNB.n510 VNB.n509 13.653
R2658 VNB.n515 VNB.n514 13.653
R2659 VNB.n514 VNB.n513 13.653
R2660 VNB.n519 VNB.n518 13.653
R2661 VNB.n518 VNB.n517 13.653
R2662 VNB.n523 VNB.n522 13.653
R2663 VNB.n522 VNB.n521 13.653
R2664 VNB.n529 VNB.n528 13.653
R2665 VNB.n533 VNB.n532 13.653
R2666 VNB.n532 VNB.n531 13.653
R2667 VNB.n537 VNB.n536 13.653
R2668 VNB.n536 VNB.n535 13.653
R2669 VNB.n559 VNB.n558 13.653
R2670 VNB.n558 VNB.n557 13.653
R2671 VNB.n563 VNB.n562 13.653
R2672 VNB.n562 VNB.n561 13.653
R2673 VNB.n567 VNB.n566 13.653
R2674 VNB.n566 VNB.n565 13.653
R2675 VNB.n571 VNB.n570 13.653
R2676 VNB.n570 VNB.n569 13.653
R2677 VNB.n577 VNB.n576 13.653
R2678 VNB.n576 VNB.n575 13.653
R2679 VNB.n588 VNB.n587 13.653
R2680 VNB.n592 VNB.n591 13.653
R2681 VNB.n591 VNB.n590 13.653
R2682 VNB.n596 VNB.n595 13.653
R2683 VNB.n595 VNB.n594 13.653
R2684 VNB.n618 VNB.n617 13.653
R2685 VNB.n617 VNB.n616 13.653
R2686 VNB.n622 VNB.n621 13.653
R2687 VNB.n621 VNB.n620 13.653
R2688 VNB.n626 VNB.n625 13.653
R2689 VNB.n625 VNB.n624 13.653
R2690 VNB.n630 VNB.n629 13.653
R2691 VNB.n629 VNB.n628 13.653
R2692 VNB.n634 VNB.n633 13.653
R2693 VNB.n633 VNB.n632 13.653
R2694 VNB.n638 VNB.n637 13.653
R2695 VNB.n637 VNB.n636 13.653
R2696 VNB.n642 VNB.n641 13.653
R2697 VNB.n641 VNB.n640 13.653
R2698 VNB.n646 VNB.n645 13.653
R2699 VNB.n645 VNB.n644 13.653
R2700 VNB.n651 VNB.n650 13.653
R2701 VNB.n650 VNB.n649 13.653
R2702 VNB.n663 VNB.n662 13.653
R2703 VNB.n662 VNB.n661 13.653
R2704 VNB.n667 VNB.n666 13.653
R2705 VNB.n666 VNB.n665 13.653
R2706 VNB.n671 VNB.n670 13.653
R2707 VNB.n670 VNB.n669 13.653
R2708 VNB.n693 VNB.n692 13.653
R2709 VNB.n692 VNB.n691 13.653
R2710 VNB.n697 VNB.n696 13.653
R2711 VNB.n696 VNB.n695 13.653
R2712 VNB.n701 VNB.n700 13.653
R2713 VNB.n700 VNB.n699 13.653
R2714 VNB.n705 VNB.n704 13.653
R2715 VNB.n704 VNB.n703 13.653
R2716 VNB.n709 VNB.n708 13.653
R2717 VNB.n708 VNB.n707 13.653
R2718 VNB.n713 VNB.n712 13.653
R2719 VNB.n712 VNB.n711 13.653
R2720 VNB.n717 VNB.n716 13.653
R2721 VNB.n716 VNB.n715 13.653
R2722 VNB.n721 VNB.n720 13.653
R2723 VNB.n720 VNB.n719 13.653
R2724 VNB.n726 VNB.n725 13.653
R2725 VNB.n725 VNB.n724 13.653
R2726 VNB.n738 VNB.n737 13.653
R2727 VNB.n737 VNB.n736 13.653
R2728 VNB.n742 VNB.n741 13.653
R2729 VNB.n741 VNB.n740 13.653
R2730 VNB.n746 VNB.n745 13.653
R2731 VNB.n745 VNB.n744 13.653
R2732 VNB.n768 VNB.n767 13.653
R2733 VNB.n767 VNB.n766 13.653
R2734 VNB.n772 VNB.n771 13.653
R2735 VNB.n771 VNB.n770 13.653
R2736 VNB.n776 VNB.n775 13.653
R2737 VNB.n775 VNB.n774 13.653
R2738 VNB.n780 VNB.n779 13.653
R2739 VNB.n779 VNB.n778 13.653
R2740 VNB.n784 VNB.n783 13.653
R2741 VNB.n783 VNB.n782 13.653
R2742 VNB.n790 VNB.n789 13.653
R2743 VNB.n82 VNB.n81 13.653
R2744 VNB.n81 VNB.n80 13.653
R2745 VNB.n85 VNB.n84 13.653
R2746 VNB.n84 VNB.n83 13.653
R2747 VNB.n90 VNB.n89 13.653
R2748 VNB.n89 VNB.n88 13.653
R2749 VNB.n93 VNB.n92 13.653
R2750 VNB.n92 VNB.n91 13.653
R2751 VNB.n96 VNB.n95 13.653
R2752 VNB.n95 VNB.n94 13.653
R2753 VNB.n99 VNB.n98 13.653
R2754 VNB.n98 VNB.n97 13.653
R2755 VNB.n102 VNB.n101 13.653
R2756 VNB.n101 VNB.n100 13.653
R2757 VNB.n105 VNB.n104 13.653
R2758 VNB.n104 VNB.n103 13.653
R2759 VNB.n108 VNB.n107 13.653
R2760 VNB.n107 VNB.n106 13.653
R2761 VNB.n111 VNB.n110 13.653
R2762 VNB.n110 VNB.n109 13.653
R2763 VNB.n806 VNB.n805 13.653
R2764 VNB.n805 VNB.n804 13.653
R2765 VNB.n817 VNB.n816 13.653
R2766 VNB.n816 VNB.n815 13.653
R2767 VNB.n821 VNB.n820 13.653
R2768 VNB.n820 VNB.n819 13.653
R2769 VNB.n825 VNB.n824 13.653
R2770 VNB.n824 VNB.n823 13.653
R2771 VNB.n847 VNB.n846 13.653
R2772 VNB.n846 VNB.n845 13.653
R2773 VNB.n851 VNB.n850 13.653
R2774 VNB.n850 VNB.n849 13.653
R2775 VNB.n855 VNB.n854 13.653
R2776 VNB.n854 VNB.n853 13.653
R2777 VNB.n859 VNB.n858 13.653
R2778 VNB.n858 VNB.n857 13.653
R2779 VNB.n863 VNB.n862 13.653
R2780 VNB.n862 VNB.n861 13.653
R2781 VNB.n867 VNB.n866 13.653
R2782 VNB.n866 VNB.n865 13.653
R2783 VNB.n871 VNB.n870 13.653
R2784 VNB.n870 VNB.n869 13.653
R2785 VNB.n875 VNB.n874 13.653
R2786 VNB.n874 VNB.n873 13.653
R2787 VNB.n879 VNB.n878 13.653
R2788 VNB.n878 VNB.n877 13.653
R2789 VNB.n885 VNB.n884 13.653
R2790 VNB.n889 VNB.n888 13.653
R2791 VNB.n888 VNB.n887 13.653
R2792 VNB.n893 VNB.n892 13.653
R2793 VNB.n892 VNB.n891 13.653
R2794 VNB.n915 VNB.n914 13.653
R2795 VNB.n914 VNB.n913 13.653
R2796 VNB.n919 VNB.n918 13.653
R2797 VNB.n918 VNB.n917 13.653
R2798 VNB.n923 VNB.n922 13.653
R2799 VNB.n922 VNB.n921 13.653
R2800 VNB.n927 VNB.n926 13.653
R2801 VNB.n926 VNB.n925 13.653
R2802 VNB.n933 VNB.n932 13.653
R2803 VNB.n932 VNB.n931 13.653
R2804 VNB.n944 VNB.n943 13.653
R2805 VNB.n948 VNB.n947 13.653
R2806 VNB.n947 VNB.n946 13.653
R2807 VNB.n952 VNB.n951 13.653
R2808 VNB.n951 VNB.n950 13.653
R2809 VNB.n974 VNB.n973 13.653
R2810 VNB.n973 VNB.n972 13.653
R2811 VNB.n978 VNB.n977 13.653
R2812 VNB.n977 VNB.n976 13.653
R2813 VNB.n982 VNB.n981 13.653
R2814 VNB.n981 VNB.n980 13.653
R2815 VNB.n986 VNB.n985 13.653
R2816 VNB.n985 VNB.n984 13.653
R2817 VNB.n990 VNB.n989 13.653
R2818 VNB.n989 VNB.n988 13.653
R2819 VNB.n994 VNB.n993 13.653
R2820 VNB.n993 VNB.n992 13.653
R2821 VNB.n998 VNB.n997 13.653
R2822 VNB.n997 VNB.n996 13.653
R2823 VNB.n1002 VNB.n1001 13.653
R2824 VNB.n1001 VNB.n1000 13.653
R2825 VNB.n1006 VNB.n1005 13.653
R2826 VNB.n1005 VNB.n1004 13.653
R2827 VNB.n1012 VNB.n1011 13.653
R2828 VNB.n1016 VNB.n1015 13.653
R2829 VNB.n1015 VNB.n1014 13.653
R2830 VNB.n1020 VNB.n1019 13.653
R2831 VNB.n1019 VNB.n1018 13.653
R2832 VNB.n1042 VNB.n1041 13.653
R2833 VNB.n1041 VNB.n1040 13.653
R2834 VNB.n1046 VNB.n1045 13.653
R2835 VNB.n1045 VNB.n1044 13.653
R2836 VNB.n1050 VNB.n1049 13.653
R2837 VNB.n1049 VNB.n1048 13.653
R2838 VNB.n1054 VNB.n1053 13.653
R2839 VNB.n1053 VNB.n1052 13.653
R2840 VNB.n1058 VNB.n1057 13.653
R2841 VNB.n1057 VNB.n1056 13.653
R2842 VNB.n1062 VNB.n1061 13.653
R2843 VNB.n1061 VNB.n1060 13.653
R2844 VNB.n1066 VNB.n1065 13.653
R2845 VNB.n1065 VNB.n1064 13.653
R2846 VNB.n1070 VNB.n1069 13.653
R2847 VNB.n1069 VNB.n1068 13.653
R2848 VNB.n1075 VNB.n1074 13.653
R2849 VNB.n1074 VNB.n1073 13.653
R2850 VNB.n1087 VNB.n1086 13.653
R2851 VNB.n1086 VNB.n1085 13.653
R2852 VNB.n1091 VNB.n1090 13.653
R2853 VNB.n1090 VNB.n1089 13.653
R2854 VNB.n1095 VNB.n1094 13.653
R2855 VNB.n1094 VNB.n1093 13.653
R2856 VNB.n1117 VNB.n1116 13.653
R2857 VNB.n1116 VNB.n1115 13.653
R2858 VNB.n1121 VNB.n1120 13.653
R2859 VNB.n1120 VNB.n1119 13.653
R2860 VNB.n1125 VNB.n1124 13.653
R2861 VNB.n1124 VNB.n1123 13.653
R2862 VNB.n1129 VNB.n1128 13.653
R2863 VNB.n1128 VNB.n1127 13.653
R2864 VNB.n1135 VNB.n1134 13.653
R2865 VNB.n1134 VNB.n1133 13.653
R2866 VNB.n1146 VNB.n1145 13.653
R2867 VNB.n1150 VNB.n1149 13.653
R2868 VNB.n1149 VNB.n1148 13.653
R2869 VNB.n1154 VNB.n1153 13.653
R2870 VNB.n1153 VNB.n1152 13.653
R2871 VNB.n1176 VNB.n1175 13.653
R2872 VNB.n1175 VNB.n1174 13.653
R2873 VNB.n1180 VNB.n1179 13.653
R2874 VNB.n1179 VNB.n1178 13.653
R2875 VNB.n1184 VNB.n1183 13.653
R2876 VNB.n1183 VNB.n1182 13.653
R2877 VNB.n1188 VNB.n1187 13.653
R2878 VNB.n1187 VNB.n1186 13.653
R2879 VNB.n1192 VNB.n1191 13.653
R2880 VNB.n1191 VNB.n1190 13.653
R2881 VNB.n1196 VNB.n1195 13.653
R2882 VNB.n1195 VNB.n1194 13.653
R2883 VNB.n1200 VNB.n1199 13.653
R2884 VNB.n1199 VNB.n1198 13.653
R2885 VNB.n1204 VNB.n1203 13.653
R2886 VNB.n1203 VNB.n1202 13.653
R2887 VNB.n1209 VNB.n1208 13.653
R2888 VNB.n1208 VNB.n1207 13.653
R2889 VNB.n1221 VNB.n1220 13.653
R2890 VNB.n1220 VNB.n1219 13.653
R2891 VNB.n1225 VNB.n1224 13.653
R2892 VNB.n1224 VNB.n1223 13.653
R2893 VNB.n1229 VNB.n1228 13.653
R2894 VNB.n1228 VNB.n1227 13.653
R2895 VNB.n1251 VNB.n1250 13.653
R2896 VNB.n1250 VNB.n1249 13.653
R2897 VNB.n1255 VNB.n1254 13.653
R2898 VNB.n1254 VNB.n1253 13.653
R2899 VNB.n1259 VNB.n1258 13.653
R2900 VNB.n1258 VNB.n1257 13.653
R2901 VNB.n1263 VNB.n1262 13.653
R2902 VNB.n1262 VNB.n1261 13.653
R2903 VNB.n1267 VNB.n1266 13.653
R2904 VNB.n1266 VNB.n1265 13.653
R2905 VNB.n1271 VNB.n1270 13.653
R2906 VNB.n1270 VNB.n1269 13.653
R2907 VNB.n1275 VNB.n1274 13.653
R2908 VNB.n1274 VNB.n1273 13.653
R2909 VNB.n1279 VNB.n1278 13.653
R2910 VNB.n1278 VNB.n1277 13.653
R2911 VNB.n1283 VNB.n1282 13.653
R2912 VNB.n1282 VNB.n1281 13.653
R2913 VNB.n1289 VNB.n1288 13.653
R2914 VNB.n1293 VNB.n1292 13.653
R2915 VNB.n1292 VNB.n1291 13.653
R2916 VNB.n1297 VNB.n1296 13.653
R2917 VNB.n1296 VNB.n1295 13.653
R2918 VNB.n1319 VNB.n1318 13.653
R2919 VNB.n1318 VNB.n1317 13.653
R2920 VNB.n1323 VNB.n1322 13.653
R2921 VNB.n1322 VNB.n1321 13.653
R2922 VNB.n1327 VNB.n1326 13.653
R2923 VNB.n1326 VNB.n1325 13.653
R2924 VNB.n1331 VNB.n1330 13.653
R2925 VNB.n1330 VNB.n1329 13.653
R2926 VNB.n1335 VNB.n1334 13.653
R2927 VNB.n1334 VNB.n1333 13.653
R2928 VNB.n1341 VNB.n1340 13.653
R2929 VNB.n1345 VNB.n1344 13.653
R2930 VNB.n1344 VNB.n1343 13.653
R2931 VNB.n1349 VNB.n1348 13.653
R2932 VNB.n1348 VNB.n1347 13.653
R2933 VNB.n1371 VNB.n1370 13.653
R2934 VNB.n1370 VNB.n1369 13.653
R2935 VNB.n1375 VNB.n1374 13.653
R2936 VNB.n1374 VNB.n1373 13.653
R2937 VNB.n1379 VNB.n1378 13.653
R2938 VNB.n1378 VNB.n1377 13.653
R2939 VNB.n1383 VNB.n1382 13.653
R2940 VNB.n1382 VNB.n1381 13.653
R2941 VNB.n1387 VNB.n1386 13.653
R2942 VNB.n1386 VNB.n1385 13.653
R2943 VNB.n1391 VNB.n1390 13.653
R2944 VNB.n1390 VNB.n1389 13.653
R2945 VNB.n1395 VNB.n1394 13.653
R2946 VNB.n1394 VNB.n1393 13.653
R2947 VNB.n1399 VNB.n1398 13.653
R2948 VNB.n1398 VNB.n1397 13.653
R2949 VNB.n1404 VNB.n1403 13.653
R2950 VNB.n1403 VNB.n1402 13.653
R2951 VNB.n1416 VNB.n1415 13.653
R2952 VNB.n1415 VNB.n1414 13.653
R2953 VNB.n1420 VNB.n1419 13.653
R2954 VNB.n1419 VNB.n1418 13.653
R2955 VNB.n1424 VNB.n1423 13.653
R2956 VNB.n1423 VNB.n1422 13.653
R2957 VNB.n28 VNB.n27 13.653
R2958 VNB.n27 VNB.n26 13.653
R2959 VNB.n31 VNB.n30 13.653
R2960 VNB.n30 VNB.n29 13.653
R2961 VNB.n34 VNB.n33 13.653
R2962 VNB.n33 VNB.n32 13.653
R2963 VNB.n37 VNB.n36 13.653
R2964 VNB.n36 VNB.n35 13.653
R2965 VNB.n40 VNB.n39 13.653
R2966 VNB.n39 VNB.n38 13.653
R2967 VNB.n43 VNB.n42 13.653
R2968 VNB.n42 VNB.n41 13.653
R2969 VNB.n46 VNB.n45 13.653
R2970 VNB.n45 VNB.n44 13.653
R2971 VNB.n49 VNB.n48 13.653
R2972 VNB.n48 VNB.n47 13.653
R2973 VNB.n53 VNB.n52 13.653
R2974 VNB.n52 VNB.n51 13.653
R2975 VNB.n58 VNB.n57 13.653
R2976 VNB.n57 VNB.n56 13.653
R2977 VNB.n63 VNB.n62 13.653
R2978 VNB.n62 VNB.n61 13.653
R2979 VNB.n1438 VNB.n0 13.653
R2980 VNB VNB.n0 13.653
R2981 VNB.n129 VNB.n128 13.653
R2982 VNB.n128 VNB.n127 13.653
R2983 VNB.n1446 VNB.n1443 13.577
R2984 VNB.n114 VNB.n112 13.276
R2985 VNB.n126 VNB.n114 13.276
R2986 VNB.n162 VNB.n160 13.276
R2987 VNB.n175 VNB.n162 13.276
R2988 VNB.n221 VNB.n219 13.276
R2989 VNB.n234 VNB.n221 13.276
R2990 VNB.n280 VNB.n278 13.276
R2991 VNB.n293 VNB.n280 13.276
R2992 VNB.n339 VNB.n337 13.276
R2993 VNB.n352 VNB.n339 13.276
R2994 VNB.n398 VNB.n396 13.276
R2995 VNB.n411 VNB.n398 13.276
R2996 VNB.n473 VNB.n471 13.276
R2997 VNB.n486 VNB.n473 13.276
R2998 VNB.n541 VNB.n539 13.276
R2999 VNB.n554 VNB.n541 13.276
R3000 VNB.n600 VNB.n598 13.276
R3001 VNB.n613 VNB.n600 13.276
R3002 VNB.n675 VNB.n673 13.276
R3003 VNB.n688 VNB.n675 13.276
R3004 VNB.n750 VNB.n748 13.276
R3005 VNB.n763 VNB.n750 13.276
R3006 VNB.n66 VNB.n64 13.276
R3007 VNB.n79 VNB.n66 13.276
R3008 VNB.n829 VNB.n827 13.276
R3009 VNB.n842 VNB.n829 13.276
R3010 VNB.n897 VNB.n895 13.276
R3011 VNB.n910 VNB.n897 13.276
R3012 VNB.n956 VNB.n954 13.276
R3013 VNB.n969 VNB.n956 13.276
R3014 VNB.n1024 VNB.n1022 13.276
R3015 VNB.n1037 VNB.n1024 13.276
R3016 VNB.n1099 VNB.n1097 13.276
R3017 VNB.n1112 VNB.n1099 13.276
R3018 VNB.n1158 VNB.n1156 13.276
R3019 VNB.n1171 VNB.n1158 13.276
R3020 VNB.n1233 VNB.n1231 13.276
R3021 VNB.n1246 VNB.n1233 13.276
R3022 VNB.n1301 VNB.n1299 13.276
R3023 VNB.n1314 VNB.n1301 13.276
R3024 VNB.n1353 VNB.n1351 13.276
R3025 VNB.n1366 VNB.n1353 13.276
R3026 VNB.n10 VNB.n8 13.276
R3027 VNB.n23 VNB.n10 13.276
R3028 VNB.n180 VNB.n176 13.276
R3029 VNB.n239 VNB.n235 13.276
R3030 VNB.n298 VNB.n294 13.276
R3031 VNB.n357 VNB.n353 13.276
R3032 VNB.n416 VNB.n412 13.276
R3033 VNB.n491 VNB.n487 13.276
R3034 VNB.n559 VNB.n555 13.276
R3035 VNB.n618 VNB.n614 13.276
R3036 VNB.n693 VNB.n689 13.276
R3037 VNB.n768 VNB.n764 13.276
R3038 VNB.n85 VNB.n82 13.276
R3039 VNB.n86 VNB.n85 13.276
R3040 VNB.n90 VNB.n86 13.276
R3041 VNB.n93 VNB.n90 13.276
R3042 VNB.n96 VNB.n93 13.276
R3043 VNB.n99 VNB.n96 13.276
R3044 VNB.n102 VNB.n99 13.276
R3045 VNB.n105 VNB.n102 13.276
R3046 VNB.n108 VNB.n105 13.276
R3047 VNB.n111 VNB.n108 13.276
R3048 VNB.n806 VNB.n111 13.276
R3049 VNB.n817 VNB.n806 13.276
R3050 VNB.n847 VNB.n843 13.276
R3051 VNB.n915 VNB.n911 13.276
R3052 VNB.n974 VNB.n970 13.276
R3053 VNB.n1042 VNB.n1038 13.276
R3054 VNB.n1117 VNB.n1113 13.276
R3055 VNB.n1176 VNB.n1172 13.276
R3056 VNB.n1251 VNB.n1247 13.276
R3057 VNB.n1319 VNB.n1315 13.276
R3058 VNB.n1371 VNB.n1367 13.276
R3059 VNB.n28 VNB.n24 13.276
R3060 VNB.n31 VNB.n28 13.276
R3061 VNB.n34 VNB.n31 13.276
R3062 VNB.n37 VNB.n34 13.276
R3063 VNB.n40 VNB.n37 13.276
R3064 VNB.n43 VNB.n40 13.276
R3065 VNB.n46 VNB.n43 13.276
R3066 VNB.n49 VNB.n46 13.276
R3067 VNB.n53 VNB.n49 13.276
R3068 VNB.n58 VNB.n53 13.276
R3069 VNB.n1438 VNB.n63 13.276
R3070 VNB.n3 VNB.n1 13.276
R3071 VNB.n1439 VNB.n3 13.276
R3072 VNB.n150 VNB.n149 12.837
R3073 VNB.n63 VNB.n59 12.02
R3074 VNB.n149 VNB.n148 7.566
R3075 VNB.n1448 VNB.n1447 7.5
R3076 VNB.n168 VNB.n167 7.5
R3077 VNB.n164 VNB.n163 7.5
R3078 VNB.n162 VNB.n161 7.5
R3079 VNB.n175 VNB.n174 7.5
R3080 VNB.n227 VNB.n226 7.5
R3081 VNB.n223 VNB.n222 7.5
R3082 VNB.n221 VNB.n220 7.5
R3083 VNB.n234 VNB.n233 7.5
R3084 VNB.n286 VNB.n285 7.5
R3085 VNB.n282 VNB.n281 7.5
R3086 VNB.n280 VNB.n279 7.5
R3087 VNB.n293 VNB.n292 7.5
R3088 VNB.n345 VNB.n344 7.5
R3089 VNB.n341 VNB.n340 7.5
R3090 VNB.n339 VNB.n338 7.5
R3091 VNB.n352 VNB.n351 7.5
R3092 VNB.n404 VNB.n403 7.5
R3093 VNB.n400 VNB.n399 7.5
R3094 VNB.n398 VNB.n397 7.5
R3095 VNB.n411 VNB.n410 7.5
R3096 VNB.n479 VNB.n478 7.5
R3097 VNB.n475 VNB.n474 7.5
R3098 VNB.n473 VNB.n472 7.5
R3099 VNB.n486 VNB.n485 7.5
R3100 VNB.n547 VNB.n546 7.5
R3101 VNB.n543 VNB.n542 7.5
R3102 VNB.n541 VNB.n540 7.5
R3103 VNB.n554 VNB.n553 7.5
R3104 VNB.n606 VNB.n605 7.5
R3105 VNB.n602 VNB.n601 7.5
R3106 VNB.n600 VNB.n599 7.5
R3107 VNB.n613 VNB.n612 7.5
R3108 VNB.n681 VNB.n680 7.5
R3109 VNB.n677 VNB.n676 7.5
R3110 VNB.n675 VNB.n674 7.5
R3111 VNB.n688 VNB.n687 7.5
R3112 VNB.n756 VNB.n755 7.5
R3113 VNB.n752 VNB.n751 7.5
R3114 VNB.n750 VNB.n749 7.5
R3115 VNB.n763 VNB.n762 7.5
R3116 VNB.n72 VNB.n71 7.5
R3117 VNB.n68 VNB.n67 7.5
R3118 VNB.n66 VNB.n65 7.5
R3119 VNB.n79 VNB.n78 7.5
R3120 VNB.n835 VNB.n834 7.5
R3121 VNB.n831 VNB.n830 7.5
R3122 VNB.n829 VNB.n828 7.5
R3123 VNB.n842 VNB.n841 7.5
R3124 VNB.n903 VNB.n902 7.5
R3125 VNB.n899 VNB.n898 7.5
R3126 VNB.n897 VNB.n896 7.5
R3127 VNB.n910 VNB.n909 7.5
R3128 VNB.n962 VNB.n961 7.5
R3129 VNB.n958 VNB.n957 7.5
R3130 VNB.n956 VNB.n955 7.5
R3131 VNB.n969 VNB.n968 7.5
R3132 VNB.n1030 VNB.n1029 7.5
R3133 VNB.n1026 VNB.n1025 7.5
R3134 VNB.n1024 VNB.n1023 7.5
R3135 VNB.n1037 VNB.n1036 7.5
R3136 VNB.n1105 VNB.n1104 7.5
R3137 VNB.n1101 VNB.n1100 7.5
R3138 VNB.n1099 VNB.n1098 7.5
R3139 VNB.n1112 VNB.n1111 7.5
R3140 VNB.n1164 VNB.n1163 7.5
R3141 VNB.n1160 VNB.n1159 7.5
R3142 VNB.n1158 VNB.n1157 7.5
R3143 VNB.n1171 VNB.n1170 7.5
R3144 VNB.n1239 VNB.n1238 7.5
R3145 VNB.n1235 VNB.n1234 7.5
R3146 VNB.n1233 VNB.n1232 7.5
R3147 VNB.n1246 VNB.n1245 7.5
R3148 VNB.n1307 VNB.n1306 7.5
R3149 VNB.n1303 VNB.n1302 7.5
R3150 VNB.n1301 VNB.n1300 7.5
R3151 VNB.n1314 VNB.n1313 7.5
R3152 VNB.n1359 VNB.n1358 7.5
R3153 VNB.n1355 VNB.n1354 7.5
R3154 VNB.n1353 VNB.n1352 7.5
R3155 VNB.n1366 VNB.n1365 7.5
R3156 VNB.n16 VNB.n15 7.5
R3157 VNB.n12 VNB.n11 7.5
R3158 VNB.n10 VNB.n9 7.5
R3159 VNB.n23 VNB.n22 7.5
R3160 VNB.n1440 VNB.n1439 7.5
R3161 VNB.n3 VNB.n2 7.5
R3162 VNB.n1445 VNB.n1444 7.5
R3163 VNB.n120 VNB.n119 7.5
R3164 VNB.n116 VNB.n115 7.5
R3165 VNB.n114 VNB.n113 7.5
R3166 VNB.n126 VNB.n125 7.5
R3167 VNB.n176 VNB.n175 7.176
R3168 VNB.n235 VNB.n234 7.176
R3169 VNB.n294 VNB.n293 7.176
R3170 VNB.n353 VNB.n352 7.176
R3171 VNB.n412 VNB.n411 7.176
R3172 VNB.n487 VNB.n486 7.176
R3173 VNB.n555 VNB.n554 7.176
R3174 VNB.n614 VNB.n613 7.176
R3175 VNB.n689 VNB.n688 7.176
R3176 VNB.n764 VNB.n763 7.176
R3177 VNB.n86 VNB.n79 7.176
R3178 VNB.n843 VNB.n842 7.176
R3179 VNB.n911 VNB.n910 7.176
R3180 VNB.n970 VNB.n969 7.176
R3181 VNB.n1038 VNB.n1037 7.176
R3182 VNB.n1113 VNB.n1112 7.176
R3183 VNB.n1172 VNB.n1171 7.176
R3184 VNB.n1247 VNB.n1246 7.176
R3185 VNB.n1315 VNB.n1314 7.176
R3186 VNB.n1367 VNB.n1366 7.176
R3187 VNB.n24 VNB.n23 7.176
R3188 VNB.n1450 VNB.n1448 7.011
R3189 VNB.n171 VNB.n168 7.011
R3190 VNB.n166 VNB.n164 7.011
R3191 VNB.n230 VNB.n227 7.011
R3192 VNB.n225 VNB.n223 7.011
R3193 VNB.n289 VNB.n286 7.011
R3194 VNB.n284 VNB.n282 7.011
R3195 VNB.n348 VNB.n345 7.011
R3196 VNB.n343 VNB.n341 7.011
R3197 VNB.n407 VNB.n404 7.011
R3198 VNB.n402 VNB.n400 7.011
R3199 VNB.n482 VNB.n479 7.011
R3200 VNB.n477 VNB.n475 7.011
R3201 VNB.n550 VNB.n547 7.011
R3202 VNB.n545 VNB.n543 7.011
R3203 VNB.n609 VNB.n606 7.011
R3204 VNB.n604 VNB.n602 7.011
R3205 VNB.n684 VNB.n681 7.011
R3206 VNB.n679 VNB.n677 7.011
R3207 VNB.n759 VNB.n756 7.011
R3208 VNB.n754 VNB.n752 7.011
R3209 VNB.n75 VNB.n72 7.011
R3210 VNB.n70 VNB.n68 7.011
R3211 VNB.n838 VNB.n835 7.011
R3212 VNB.n833 VNB.n831 7.011
R3213 VNB.n906 VNB.n903 7.011
R3214 VNB.n901 VNB.n899 7.011
R3215 VNB.n965 VNB.n962 7.011
R3216 VNB.n960 VNB.n958 7.011
R3217 VNB.n1033 VNB.n1030 7.011
R3218 VNB.n1028 VNB.n1026 7.011
R3219 VNB.n1108 VNB.n1105 7.011
R3220 VNB.n1103 VNB.n1101 7.011
R3221 VNB.n1167 VNB.n1164 7.011
R3222 VNB.n1162 VNB.n1160 7.011
R3223 VNB.n1242 VNB.n1239 7.011
R3224 VNB.n1237 VNB.n1235 7.011
R3225 VNB.n1310 VNB.n1307 7.011
R3226 VNB.n1305 VNB.n1303 7.011
R3227 VNB.n1362 VNB.n1359 7.011
R3228 VNB.n1357 VNB.n1355 7.011
R3229 VNB.n19 VNB.n16 7.011
R3230 VNB.n14 VNB.n12 7.011
R3231 VNB.n122 VNB.n120 7.011
R3232 VNB.n118 VNB.n116 7.011
R3233 VNB.n174 VNB.n173 7.01
R3234 VNB.n166 VNB.n165 7.01
R3235 VNB.n171 VNB.n170 7.01
R3236 VNB.n233 VNB.n232 7.01
R3237 VNB.n225 VNB.n224 7.01
R3238 VNB.n230 VNB.n229 7.01
R3239 VNB.n292 VNB.n291 7.01
R3240 VNB.n284 VNB.n283 7.01
R3241 VNB.n289 VNB.n288 7.01
R3242 VNB.n351 VNB.n350 7.01
R3243 VNB.n343 VNB.n342 7.01
R3244 VNB.n348 VNB.n347 7.01
R3245 VNB.n410 VNB.n409 7.01
R3246 VNB.n402 VNB.n401 7.01
R3247 VNB.n407 VNB.n406 7.01
R3248 VNB.n485 VNB.n484 7.01
R3249 VNB.n477 VNB.n476 7.01
R3250 VNB.n482 VNB.n481 7.01
R3251 VNB.n553 VNB.n552 7.01
R3252 VNB.n545 VNB.n544 7.01
R3253 VNB.n550 VNB.n549 7.01
R3254 VNB.n612 VNB.n611 7.01
R3255 VNB.n604 VNB.n603 7.01
R3256 VNB.n609 VNB.n608 7.01
R3257 VNB.n687 VNB.n686 7.01
R3258 VNB.n679 VNB.n678 7.01
R3259 VNB.n684 VNB.n683 7.01
R3260 VNB.n762 VNB.n761 7.01
R3261 VNB.n754 VNB.n753 7.01
R3262 VNB.n759 VNB.n758 7.01
R3263 VNB.n78 VNB.n77 7.01
R3264 VNB.n70 VNB.n69 7.01
R3265 VNB.n75 VNB.n74 7.01
R3266 VNB.n841 VNB.n840 7.01
R3267 VNB.n833 VNB.n832 7.01
R3268 VNB.n838 VNB.n837 7.01
R3269 VNB.n909 VNB.n908 7.01
R3270 VNB.n901 VNB.n900 7.01
R3271 VNB.n906 VNB.n905 7.01
R3272 VNB.n968 VNB.n967 7.01
R3273 VNB.n960 VNB.n959 7.01
R3274 VNB.n965 VNB.n964 7.01
R3275 VNB.n1036 VNB.n1035 7.01
R3276 VNB.n1028 VNB.n1027 7.01
R3277 VNB.n1033 VNB.n1032 7.01
R3278 VNB.n1111 VNB.n1110 7.01
R3279 VNB.n1103 VNB.n1102 7.01
R3280 VNB.n1108 VNB.n1107 7.01
R3281 VNB.n1170 VNB.n1169 7.01
R3282 VNB.n1162 VNB.n1161 7.01
R3283 VNB.n1167 VNB.n1166 7.01
R3284 VNB.n1245 VNB.n1244 7.01
R3285 VNB.n1237 VNB.n1236 7.01
R3286 VNB.n1242 VNB.n1241 7.01
R3287 VNB.n1313 VNB.n1312 7.01
R3288 VNB.n1305 VNB.n1304 7.01
R3289 VNB.n1310 VNB.n1309 7.01
R3290 VNB.n1365 VNB.n1364 7.01
R3291 VNB.n1357 VNB.n1356 7.01
R3292 VNB.n1362 VNB.n1361 7.01
R3293 VNB.n22 VNB.n21 7.01
R3294 VNB.n14 VNB.n13 7.01
R3295 VNB.n19 VNB.n18 7.01
R3296 VNB.n125 VNB.n124 7.01
R3297 VNB.n118 VNB.n117 7.01
R3298 VNB.n122 VNB.n121 7.01
R3299 VNB.n1450 VNB.n1449 7.01
R3300 VNB.n1446 VNB.n1445 6.788
R3301 VNB.n1441 VNB.n1440 6.788
R3302 VNB.n140 VNB.n139 4.551
R3303 VNB.n137 VNB.n134 4.305
R3304 VNB.n154 VNB.n151 3.947
R3305 VNB.n209 VNB.n204 2.511
R3306 VNB.n268 VNB.n263 2.511
R3307 VNB.n327 VNB.n322 2.511
R3308 VNB.n386 VNB.n381 2.511
R3309 VNB.n588 VNB.n583 2.511
R3310 VNB.n790 VNB.n787 2.511
R3311 VNB.n944 VNB.n939 2.511
R3312 VNB.n1146 VNB.n1141 2.511
R3313 VNB.n1341 VNB.n1338 2.511
R3314 VNB.t10 VNB.n140 2.238
R3315 VNB.n207 VNB.n205 1.99
R3316 VNB.n266 VNB.n264 1.99
R3317 VNB.n325 VNB.n323 1.99
R3318 VNB.n384 VNB.n382 1.99
R3319 VNB.n586 VNB.n584 1.99
R3320 VNB.n942 VNB.n940 1.99
R3321 VNB.n1144 VNB.n1142 1.99
R3322 VNB.n461 VNB.n455 1.255
R3323 VNB.n529 VNB.n526 1.255
R3324 VNB.n663 VNB.n657 1.255
R3325 VNB.n738 VNB.n732 1.255
R3326 VNB.n817 VNB.n811 1.255
R3327 VNB.n885 VNB.n882 1.255
R3328 VNB.n1012 VNB.n1009 1.255
R3329 VNB.n1087 VNB.n1081 1.255
R3330 VNB.n1221 VNB.n1215 1.255
R3331 VNB.n1289 VNB.n1286 1.255
R3332 VNB.n1416 VNB.n1410 1.255
R3333 VNB.n59 VNB.n58 1.255
R3334 VNB.n1451 VNB.n1442 0.921
R3335 VNB.n1451 VNB.n1446 0.476
R3336 VNB.n1451 VNB.n1441 0.475
R3337 VNB.n142 VNB.n141 0.358
R3338 VNB.n181 VNB.n159 0.272
R3339 VNB.n240 VNB.n218 0.272
R3340 VNB.n299 VNB.n277 0.272
R3341 VNB.n358 VNB.n336 0.272
R3342 VNB.n417 VNB.n395 0.272
R3343 VNB.n492 VNB.n470 0.272
R3344 VNB.n560 VNB.n538 0.272
R3345 VNB.n619 VNB.n597 0.272
R3346 VNB.n694 VNB.n672 0.272
R3347 VNB.n769 VNB.n747 0.272
R3348 VNB.n794 VNB.n793 0.272
R3349 VNB.n848 VNB.n826 0.272
R3350 VNB.n916 VNB.n894 0.272
R3351 VNB.n975 VNB.n953 0.272
R3352 VNB.n1043 VNB.n1021 0.272
R3353 VNB.n1118 VNB.n1096 0.272
R3354 VNB.n1177 VNB.n1155 0.272
R3355 VNB.n1252 VNB.n1230 0.272
R3356 VNB.n1320 VNB.n1298 0.272
R3357 VNB.n1372 VNB.n1350 0.272
R3358 VNB.n1426 VNB.n1425 0.272
R3359 VNB.n172 VNB.n166 0.246
R3360 VNB.n173 VNB.n172 0.246
R3361 VNB.n172 VNB.n171 0.246
R3362 VNB.n231 VNB.n225 0.246
R3363 VNB.n232 VNB.n231 0.246
R3364 VNB.n231 VNB.n230 0.246
R3365 VNB.n290 VNB.n284 0.246
R3366 VNB.n291 VNB.n290 0.246
R3367 VNB.n290 VNB.n289 0.246
R3368 VNB.n349 VNB.n343 0.246
R3369 VNB.n350 VNB.n349 0.246
R3370 VNB.n349 VNB.n348 0.246
R3371 VNB.n408 VNB.n402 0.246
R3372 VNB.n409 VNB.n408 0.246
R3373 VNB.n408 VNB.n407 0.246
R3374 VNB.n483 VNB.n477 0.246
R3375 VNB.n484 VNB.n483 0.246
R3376 VNB.n483 VNB.n482 0.246
R3377 VNB.n551 VNB.n545 0.246
R3378 VNB.n552 VNB.n551 0.246
R3379 VNB.n551 VNB.n550 0.246
R3380 VNB.n610 VNB.n604 0.246
R3381 VNB.n611 VNB.n610 0.246
R3382 VNB.n610 VNB.n609 0.246
R3383 VNB.n685 VNB.n679 0.246
R3384 VNB.n686 VNB.n685 0.246
R3385 VNB.n685 VNB.n684 0.246
R3386 VNB.n760 VNB.n754 0.246
R3387 VNB.n761 VNB.n760 0.246
R3388 VNB.n760 VNB.n759 0.246
R3389 VNB.n76 VNB.n70 0.246
R3390 VNB.n77 VNB.n76 0.246
R3391 VNB.n76 VNB.n75 0.246
R3392 VNB.n839 VNB.n833 0.246
R3393 VNB.n840 VNB.n839 0.246
R3394 VNB.n839 VNB.n838 0.246
R3395 VNB.n907 VNB.n901 0.246
R3396 VNB.n908 VNB.n907 0.246
R3397 VNB.n907 VNB.n906 0.246
R3398 VNB.n966 VNB.n960 0.246
R3399 VNB.n967 VNB.n966 0.246
R3400 VNB.n966 VNB.n965 0.246
R3401 VNB.n1034 VNB.n1028 0.246
R3402 VNB.n1035 VNB.n1034 0.246
R3403 VNB.n1034 VNB.n1033 0.246
R3404 VNB.n1109 VNB.n1103 0.246
R3405 VNB.n1110 VNB.n1109 0.246
R3406 VNB.n1109 VNB.n1108 0.246
R3407 VNB.n1168 VNB.n1162 0.246
R3408 VNB.n1169 VNB.n1168 0.246
R3409 VNB.n1168 VNB.n1167 0.246
R3410 VNB.n1243 VNB.n1237 0.246
R3411 VNB.n1244 VNB.n1243 0.246
R3412 VNB.n1243 VNB.n1242 0.246
R3413 VNB.n1311 VNB.n1305 0.246
R3414 VNB.n1312 VNB.n1311 0.246
R3415 VNB.n1311 VNB.n1310 0.246
R3416 VNB.n1363 VNB.n1357 0.246
R3417 VNB.n1364 VNB.n1363 0.246
R3418 VNB.n1363 VNB.n1362 0.246
R3419 VNB.n20 VNB.n14 0.246
R3420 VNB.n21 VNB.n20 0.246
R3421 VNB.n20 VNB.n19 0.246
R3422 VNB.n123 VNB.n118 0.246
R3423 VNB.n124 VNB.n123 0.246
R3424 VNB.n123 VNB.n122 0.246
R3425 VNB.n1451 VNB.n1450 0.246
R3426 VNB.n1437 VNB 0.198
R3427 VNB.n146 VNB.n143 0.179
R3428 VNB.n147 VNB.n138 0.136
R3429 VNB.n155 VNB.n147 0.136
R3430 VNB.n159 VNB.n155 0.136
R3431 VNB.n185 VNB.n181 0.136
R3432 VNB.n189 VNB.n185 0.136
R3433 VNB.n193 VNB.n189 0.136
R3434 VNB.n199 VNB.n193 0.136
R3435 VNB.n210 VNB.n199 0.136
R3436 VNB.n214 VNB.n210 0.136
R3437 VNB.n218 VNB.n214 0.136
R3438 VNB.n244 VNB.n240 0.136
R3439 VNB.n248 VNB.n244 0.136
R3440 VNB.n252 VNB.n248 0.136
R3441 VNB.n258 VNB.n252 0.136
R3442 VNB.n269 VNB.n258 0.136
R3443 VNB.n273 VNB.n269 0.136
R3444 VNB.n277 VNB.n273 0.136
R3445 VNB.n303 VNB.n299 0.136
R3446 VNB.n307 VNB.n303 0.136
R3447 VNB.n311 VNB.n307 0.136
R3448 VNB.n317 VNB.n311 0.136
R3449 VNB.n328 VNB.n317 0.136
R3450 VNB.n332 VNB.n328 0.136
R3451 VNB.n336 VNB.n332 0.136
R3452 VNB.n362 VNB.n358 0.136
R3453 VNB.n366 VNB.n362 0.136
R3454 VNB.n370 VNB.n366 0.136
R3455 VNB.n376 VNB.n370 0.136
R3456 VNB.n387 VNB.n376 0.136
R3457 VNB.n391 VNB.n387 0.136
R3458 VNB.n395 VNB.n391 0.136
R3459 VNB.n421 VNB.n417 0.136
R3460 VNB.n425 VNB.n421 0.136
R3461 VNB.n429 VNB.n425 0.136
R3462 VNB.n433 VNB.n429 0.136
R3463 VNB.n437 VNB.n433 0.136
R3464 VNB.n441 VNB.n437 0.136
R3465 VNB.n445 VNB.n441 0.136
R3466 VNB.n450 VNB.n445 0.136
R3467 VNB.n462 VNB.n450 0.136
R3468 VNB.n466 VNB.n462 0.136
R3469 VNB.n470 VNB.n466 0.136
R3470 VNB.n496 VNB.n492 0.136
R3471 VNB.n500 VNB.n496 0.136
R3472 VNB.n504 VNB.n500 0.136
R3473 VNB.n508 VNB.n504 0.136
R3474 VNB.n512 VNB.n508 0.136
R3475 VNB.n516 VNB.n512 0.136
R3476 VNB.n520 VNB.n516 0.136
R3477 VNB.n524 VNB.n520 0.136
R3478 VNB.n530 VNB.n524 0.136
R3479 VNB.n534 VNB.n530 0.136
R3480 VNB.n538 VNB.n534 0.136
R3481 VNB.n564 VNB.n560 0.136
R3482 VNB.n568 VNB.n564 0.136
R3483 VNB.n572 VNB.n568 0.136
R3484 VNB.n578 VNB.n572 0.136
R3485 VNB.n589 VNB.n578 0.136
R3486 VNB.n593 VNB.n589 0.136
R3487 VNB.n597 VNB.n593 0.136
R3488 VNB.n623 VNB.n619 0.136
R3489 VNB.n627 VNB.n623 0.136
R3490 VNB.n631 VNB.n627 0.136
R3491 VNB.n635 VNB.n631 0.136
R3492 VNB.n639 VNB.n635 0.136
R3493 VNB.n643 VNB.n639 0.136
R3494 VNB.n647 VNB.n643 0.136
R3495 VNB.n652 VNB.n647 0.136
R3496 VNB.n664 VNB.n652 0.136
R3497 VNB.n668 VNB.n664 0.136
R3498 VNB.n672 VNB.n668 0.136
R3499 VNB.n698 VNB.n694 0.136
R3500 VNB.n702 VNB.n698 0.136
R3501 VNB.n706 VNB.n702 0.136
R3502 VNB.n710 VNB.n706 0.136
R3503 VNB.n714 VNB.n710 0.136
R3504 VNB.n718 VNB.n714 0.136
R3505 VNB.n722 VNB.n718 0.136
R3506 VNB.n727 VNB.n722 0.136
R3507 VNB.n739 VNB.n727 0.136
R3508 VNB.n743 VNB.n739 0.136
R3509 VNB.n747 VNB.n743 0.136
R3510 VNB.n773 VNB.n769 0.136
R3511 VNB.n777 VNB.n773 0.136
R3512 VNB.n781 VNB.n777 0.136
R3513 VNB.n785 VNB.n781 0.136
R3514 VNB.n791 VNB.n785 0.136
R3515 VNB.n792 VNB.n791 0.136
R3516 VNB.n793 VNB.n792 0.136
R3517 VNB.n795 VNB.n794 0.136
R3518 VNB.n796 VNB.n795 0.136
R3519 VNB.n797 VNB.n796 0.136
R3520 VNB.n798 VNB.n797 0.136
R3521 VNB.n799 VNB.n798 0.136
R3522 VNB.n800 VNB.n799 0.136
R3523 VNB.n801 VNB.n800 0.136
R3524 VNB.n802 VNB.n801 0.136
R3525 VNB.n822 VNB.n818 0.136
R3526 VNB.n826 VNB.n822 0.136
R3527 VNB.n852 VNB.n848 0.136
R3528 VNB.n856 VNB.n852 0.136
R3529 VNB.n860 VNB.n856 0.136
R3530 VNB.n864 VNB.n860 0.136
R3531 VNB.n868 VNB.n864 0.136
R3532 VNB.n872 VNB.n868 0.136
R3533 VNB.n876 VNB.n872 0.136
R3534 VNB.n880 VNB.n876 0.136
R3535 VNB.n886 VNB.n880 0.136
R3536 VNB.n890 VNB.n886 0.136
R3537 VNB.n894 VNB.n890 0.136
R3538 VNB.n920 VNB.n916 0.136
R3539 VNB.n924 VNB.n920 0.136
R3540 VNB.n928 VNB.n924 0.136
R3541 VNB.n934 VNB.n928 0.136
R3542 VNB.n945 VNB.n934 0.136
R3543 VNB.n949 VNB.n945 0.136
R3544 VNB.n953 VNB.n949 0.136
R3545 VNB.n979 VNB.n975 0.136
R3546 VNB.n983 VNB.n979 0.136
R3547 VNB.n987 VNB.n983 0.136
R3548 VNB.n991 VNB.n987 0.136
R3549 VNB.n995 VNB.n991 0.136
R3550 VNB.n999 VNB.n995 0.136
R3551 VNB.n1003 VNB.n999 0.136
R3552 VNB.n1007 VNB.n1003 0.136
R3553 VNB.n1013 VNB.n1007 0.136
R3554 VNB.n1017 VNB.n1013 0.136
R3555 VNB.n1021 VNB.n1017 0.136
R3556 VNB.n1047 VNB.n1043 0.136
R3557 VNB.n1051 VNB.n1047 0.136
R3558 VNB.n1055 VNB.n1051 0.136
R3559 VNB.n1059 VNB.n1055 0.136
R3560 VNB.n1063 VNB.n1059 0.136
R3561 VNB.n1067 VNB.n1063 0.136
R3562 VNB.n1071 VNB.n1067 0.136
R3563 VNB.n1076 VNB.n1071 0.136
R3564 VNB.n1088 VNB.n1076 0.136
R3565 VNB.n1092 VNB.n1088 0.136
R3566 VNB.n1096 VNB.n1092 0.136
R3567 VNB.n1122 VNB.n1118 0.136
R3568 VNB.n1126 VNB.n1122 0.136
R3569 VNB.n1130 VNB.n1126 0.136
R3570 VNB.n1136 VNB.n1130 0.136
R3571 VNB.n1147 VNB.n1136 0.136
R3572 VNB.n1151 VNB.n1147 0.136
R3573 VNB.n1155 VNB.n1151 0.136
R3574 VNB.n1181 VNB.n1177 0.136
R3575 VNB.n1185 VNB.n1181 0.136
R3576 VNB.n1189 VNB.n1185 0.136
R3577 VNB.n1193 VNB.n1189 0.136
R3578 VNB.n1197 VNB.n1193 0.136
R3579 VNB.n1201 VNB.n1197 0.136
R3580 VNB.n1205 VNB.n1201 0.136
R3581 VNB.n1210 VNB.n1205 0.136
R3582 VNB.n1222 VNB.n1210 0.136
R3583 VNB.n1226 VNB.n1222 0.136
R3584 VNB.n1230 VNB.n1226 0.136
R3585 VNB.n1256 VNB.n1252 0.136
R3586 VNB.n1260 VNB.n1256 0.136
R3587 VNB.n1264 VNB.n1260 0.136
R3588 VNB.n1268 VNB.n1264 0.136
R3589 VNB.n1272 VNB.n1268 0.136
R3590 VNB.n1276 VNB.n1272 0.136
R3591 VNB.n1280 VNB.n1276 0.136
R3592 VNB.n1284 VNB.n1280 0.136
R3593 VNB.n1290 VNB.n1284 0.136
R3594 VNB.n1294 VNB.n1290 0.136
R3595 VNB.n1298 VNB.n1294 0.136
R3596 VNB.n1324 VNB.n1320 0.136
R3597 VNB.n1328 VNB.n1324 0.136
R3598 VNB.n1332 VNB.n1328 0.136
R3599 VNB.n1336 VNB.n1332 0.136
R3600 VNB.n1342 VNB.n1336 0.136
R3601 VNB.n1346 VNB.n1342 0.136
R3602 VNB.n1350 VNB.n1346 0.136
R3603 VNB.n1376 VNB.n1372 0.136
R3604 VNB.n1380 VNB.n1376 0.136
R3605 VNB.n1384 VNB.n1380 0.136
R3606 VNB.n1388 VNB.n1384 0.136
R3607 VNB.n1392 VNB.n1388 0.136
R3608 VNB.n1396 VNB.n1392 0.136
R3609 VNB.n1400 VNB.n1396 0.136
R3610 VNB.n1405 VNB.n1400 0.136
R3611 VNB.n1417 VNB.n1405 0.136
R3612 VNB.n1421 VNB.n1417 0.136
R3613 VNB.n1425 VNB.n1421 0.136
R3614 VNB.n1427 VNB.n1426 0.136
R3615 VNB.n1428 VNB.n1427 0.136
R3616 VNB.n1429 VNB.n1428 0.136
R3617 VNB.n1430 VNB.n1429 0.136
R3618 VNB.n1431 VNB.n1430 0.136
R3619 VNB.n1432 VNB.n1431 0.136
R3620 VNB.n1433 VNB.n1432 0.136
R3621 VNB.n1434 VNB.n1433 0.136
R3622 VNB.n1435 VNB.n1434 0.136
R3623 VNB.n1436 VNB.n1435 0.136
R3624 VNB.n1437 VNB.n1436 0.136
R3625 VNB.n802 VNB 0.068
R3626 VNB.n818 VNB 0.068
R3627 a_599_943.n6 a_599_943.t7 480.392
R3628 a_599_943.n8 a_599_943.t11 454.685
R3629 a_599_943.n8 a_599_943.t9 428.979
R3630 a_599_943.n6 a_599_943.t10 403.272
R3631 a_599_943.n7 a_599_943.t8 266.974
R3632 a_599_943.n9 a_599_943.t12 221.453
R3633 a_599_943.n13 a_599_943.n11 196.598
R3634 a_599_943.n11 a_599_943.n5 180.846
R3635 a_599_943.n9 a_599_943.n8 108.494
R3636 a_599_943.n7 a_599_943.n6 108.494
R3637 a_599_943.n10 a_599_943.n9 80.035
R3638 a_599_943.n4 a_599_943.n3 79.232
R3639 a_599_943.n10 a_599_943.n7 77.315
R3640 a_599_943.n11 a_599_943.n10 76
R3641 a_599_943.n5 a_599_943.n4 63.152
R3642 a_599_943.n13 a_599_943.n12 30
R3643 a_599_943.n14 a_599_943.n0 24.383
R3644 a_599_943.n14 a_599_943.n13 23.684
R3645 a_599_943.n5 a_599_943.n1 16.08
R3646 a_599_943.n4 a_599_943.n2 16.08
R3647 a_599_943.n1 a_599_943.t4 14.282
R3648 a_599_943.n1 a_599_943.t5 14.282
R3649 a_599_943.n2 a_599_943.t0 14.282
R3650 a_599_943.n2 a_599_943.t1 14.282
R3651 a_599_943.n3 a_599_943.t3 14.282
R3652 a_599_943.n3 a_599_943.t2 14.282
R3653 a_15932_181.n4 a_15932_181.t8 512.525
R3654 a_15932_181.n4 a_15932_181.t9 371.139
R3655 a_15932_181.n5 a_15932_181.t7 273.368
R3656 a_15932_181.n16 a_15932_181.n6 226.775
R3657 a_15932_181.n6 a_15932_181.n5 153.043
R3658 a_15932_181.n6 a_15932_181.n3 110.158
R3659 a_15932_181.n5 a_15932_181.n4 105.194
R3660 a_15932_181.n15 a_15932_181.n14 98.501
R3661 a_15932_181.n15 a_15932_181.n10 96.417
R3662 a_15932_181.n16 a_15932_181.n15 78.403
R3663 a_15932_181.n3 a_15932_181.n2 75.271
R3664 a_15932_181.n19 a_15932_181.n0 55.263
R3665 a_15932_181.n10 a_15932_181.n9 30
R3666 a_15932_181.n14 a_15932_181.n13 30
R3667 a_15932_181.n18 a_15932_181.n17 30
R3668 a_15932_181.n19 a_15932_181.n18 25.263
R3669 a_15932_181.n8 a_15932_181.n7 24.383
R3670 a_15932_181.n12 a_15932_181.n11 24.383
R3671 a_15932_181.n10 a_15932_181.n8 23.684
R3672 a_15932_181.n14 a_15932_181.n12 23.684
R3673 a_15932_181.n18 a_15932_181.n16 20.417
R3674 a_15932_181.n1 a_15932_181.t3 14.282
R3675 a_15932_181.n1 a_15932_181.t2 14.282
R3676 a_15932_181.n2 a_15932_181.t5 14.282
R3677 a_15932_181.n2 a_15932_181.t6 14.282
R3678 a_15932_181.n3 a_15932_181.n1 12.119
R3679 a_3643_75.n4 a_3643_75.n3 19.724
R3680 a_3643_75.t0 a_3643_75.n5 11.595
R3681 a_3643_75.t0 a_3643_75.n4 9.207
R3682 a_3643_75.n2 a_3643_75.n0 8.543
R3683 a_3643_75.t0 a_3643_75.n2 3.034
R3684 a_3643_75.n2 a_3643_75.n1 0.443
R3685 a_91_75.n1 a_91_75.n0 25.576
R3686 a_91_75.n3 a_91_75.n2 9.111
R3687 a_91_75.n7 a_91_75.n5 7.859
R3688 a_91_75.t0 a_91_75.n7 3.034
R3689 a_91_75.n5 a_91_75.n3 1.964
R3690 a_91_75.n5 a_91_75.n4 1.964
R3691 a_91_75.t0 a_91_75.n1 1.871
R3692 a_91_75.n7 a_91_75.n6 0.443
R3693 a_372_182.n8 a_372_182.n6 96.467
R3694 a_372_182.n3 a_372_182.n1 44.628
R3695 a_372_182.t0 a_372_182.n8 32.417
R3696 a_372_182.n3 a_372_182.n2 23.284
R3697 a_372_182.n6 a_372_182.n5 22.349
R3698 a_372_182.t0 a_372_182.n10 20.241
R3699 a_372_182.n10 a_372_182.n9 13.494
R3700 a_372_182.n6 a_372_182.n4 8.443
R3701 a_372_182.t0 a_372_182.n0 8.137
R3702 a_372_182.t0 a_372_182.n3 5.727
R3703 a_372_182.n8 a_372_182.n7 1.435
R3704 a_5271_75.n4 a_5271_75.n3 19.724
R3705 a_5271_75.t0 a_5271_75.n5 11.595
R3706 a_5271_75.t0 a_5271_75.n4 9.207
R3707 a_5271_75.n2 a_5271_75.n0 8.543
R3708 a_5271_75.t0 a_5271_75.n2 3.034
R3709 a_5271_75.n2 a_5271_75.n1 0.443
R3710 a_5552_182.n10 a_5552_182.n8 82.852
R3711 a_5552_182.n11 a_5552_182.n0 49.6
R3712 a_5552_182.n7 a_5552_182.n6 32.833
R3713 a_5552_182.n8 a_5552_182.t1 32.416
R3714 a_5552_182.n10 a_5552_182.n9 27.2
R3715 a_5552_182.n3 a_5552_182.n2 23.284
R3716 a_5552_182.n11 a_5552_182.n10 22.4
R3717 a_5552_182.n7 a_5552_182.n4 19.017
R3718 a_5552_182.n6 a_5552_182.n5 13.494
R3719 a_5552_182.t1 a_5552_182.n1 7.04
R3720 a_5552_182.t1 a_5552_182.n3 5.727
R3721 a_5552_182.n8 a_5552_182.n7 1.435
R3722 a_16318_73.n2 a_16318_73.n0 34.602
R3723 a_16318_73.n2 a_16318_73.n1 2.138
R3724 a_16318_73.t0 a_16318_73.n2 0.069
R3725 a_2141_1004.n4 a_2141_1004.t6 512.525
R3726 a_2141_1004.n4 a_2141_1004.t7 371.139
R3727 a_2141_1004.n5 a_2141_1004.t5 271.162
R3728 a_2141_1004.n8 a_2141_1004.n6 194.086
R3729 a_2141_1004.n5 a_2141_1004.n4 172.76
R3730 a_2141_1004.n6 a_2141_1004.n3 162.547
R3731 a_2141_1004.n6 a_2141_1004.n5 153.315
R3732 a_2141_1004.n3 a_2141_1004.n2 76.002
R3733 a_2141_1004.n8 a_2141_1004.n7 30
R3734 a_2141_1004.n9 a_2141_1004.n0 24.383
R3735 a_2141_1004.n9 a_2141_1004.n8 23.684
R3736 a_2141_1004.n1 a_2141_1004.t3 14.282
R3737 a_2141_1004.n1 a_2141_1004.t2 14.282
R3738 a_2141_1004.n2 a_2141_1004.t1 14.282
R3739 a_2141_1004.n2 a_2141_1004.t0 14.282
R3740 a_2141_1004.n3 a_2141_1004.n1 12.85
R3741 a_9009_1004.n6 a_9009_1004.t8 480.392
R3742 a_9009_1004.n6 a_9009_1004.t7 403.272
R3743 a_9009_1004.n7 a_9009_1004.t9 293.527
R3744 a_9009_1004.n10 a_9009_1004.n8 223.151
R3745 a_9009_1004.n8 a_9009_1004.n5 154.293
R3746 a_9009_1004.n8 a_9009_1004.n7 153.315
R3747 a_9009_1004.n7 a_9009_1004.n6 81.941
R3748 a_9009_1004.n4 a_9009_1004.n3 79.232
R3749 a_9009_1004.n5 a_9009_1004.n4 63.152
R3750 a_9009_1004.n10 a_9009_1004.n9 30
R3751 a_9009_1004.n11 a_9009_1004.n0 24.383
R3752 a_9009_1004.n11 a_9009_1004.n10 23.684
R3753 a_9009_1004.n5 a_9009_1004.n1 16.08
R3754 a_9009_1004.n4 a_9009_1004.n2 16.08
R3755 a_9009_1004.n1 a_9009_1004.t1 14.282
R3756 a_9009_1004.n1 a_9009_1004.t0 14.282
R3757 a_9009_1004.n2 a_9009_1004.t6 14.282
R3758 a_9009_1004.n2 a_9009_1004.t5 14.282
R3759 a_9009_1004.n3 a_9009_1004.t4 14.282
R3760 a_9009_1004.n3 a_9009_1004.t3 14.282
R3761 a_4626_73.n12 a_4626_73.n11 26.811
R3762 a_4626_73.n6 a_4626_73.n5 24.977
R3763 a_4626_73.n2 a_4626_73.n1 24.877
R3764 a_4626_73.t0 a_4626_73.n2 12.677
R3765 a_4626_73.t0 a_4626_73.n3 11.595
R3766 a_4626_73.t1 a_4626_73.n8 8.137
R3767 a_4626_73.t0 a_4626_73.n4 7.273
R3768 a_4626_73.t0 a_4626_73.n0 6.109
R3769 a_4626_73.t1 a_4626_73.n7 4.864
R3770 a_4626_73.t0 a_4626_73.n12 2.074
R3771 a_4626_73.n7 a_4626_73.n6 1.13
R3772 a_4626_73.n12 a_4626_73.t1 0.937
R3773 a_4626_73.t1 a_4626_73.n10 0.804
R3774 a_4626_73.n10 a_4626_73.n9 0.136
R3775 a_2036_73.n12 a_2036_73.n11 26.811
R3776 a_2036_73.n6 a_2036_73.n5 24.977
R3777 a_2036_73.n2 a_2036_73.n1 24.877
R3778 a_2036_73.t0 a_2036_73.n2 12.677
R3779 a_2036_73.t0 a_2036_73.n3 11.595
R3780 a_2036_73.t1 a_2036_73.n8 8.137
R3781 a_2036_73.t0 a_2036_73.n4 7.273
R3782 a_2036_73.t0 a_2036_73.n0 6.109
R3783 a_2036_73.t1 a_2036_73.n7 4.864
R3784 a_2036_73.t0 a_2036_73.n12 2.074
R3785 a_2036_73.n7 a_2036_73.n6 1.13
R3786 a_2036_73.n12 a_2036_73.t1 0.937
R3787 a_2036_73.t1 a_2036_73.n10 0.804
R3788 a_2036_73.n10 a_2036_73.n9 0.136
R3789 a_14003_75.n5 a_14003_75.n4 19.724
R3790 a_14003_75.t0 a_14003_75.n3 11.595
R3791 a_14003_75.t0 a_14003_75.n5 9.207
R3792 a_14003_75.n2 a_14003_75.n1 2.455
R3793 a_14003_75.n2 a_14003_75.n0 1.32
R3794 a_14003_75.t0 a_14003_75.n2 0.246
R3795 a_2681_75.n4 a_2681_75.n3 19.724
R3796 a_2681_75.t0 a_2681_75.n5 11.595
R3797 a_2681_75.t0 a_2681_75.n4 9.207
R3798 a_2681_75.n2 a_2681_75.n0 8.543
R3799 a_2681_75.t0 a_2681_75.n2 3.034
R3800 a_2681_75.n2 a_2681_75.n1 0.443
R3801 a_1334_182.n10 a_1334_182.n8 82.852
R3802 a_1334_182.n7 a_1334_182.n6 32.833
R3803 a_1334_182.n8 a_1334_182.t1 32.416
R3804 a_1334_182.n10 a_1334_182.n9 27.2
R3805 a_1334_182.n11 a_1334_182.n0 23.498
R3806 a_1334_182.n3 a_1334_182.n2 23.284
R3807 a_1334_182.n11 a_1334_182.n10 22.4
R3808 a_1334_182.n7 a_1334_182.n4 19.017
R3809 a_1334_182.n6 a_1334_182.n5 13.494
R3810 a_1334_182.t1 a_1334_182.n1 7.04
R3811 a_1334_182.t1 a_1334_182.n3 5.727
R3812 a_1334_182.n8 a_1334_182.n7 1.435
R3813 a_10732_182.n9 a_10732_182.n7 82.852
R3814 a_10732_182.n3 a_10732_182.n1 44.628
R3815 a_10732_182.t0 a_10732_182.n9 32.417
R3816 a_10732_182.n7 a_10732_182.n6 27.2
R3817 a_10732_182.n5 a_10732_182.n4 23.498
R3818 a_10732_182.n3 a_10732_182.n2 23.284
R3819 a_10732_182.n7 a_10732_182.n5 22.4
R3820 a_10732_182.t0 a_10732_182.n11 20.241
R3821 a_10732_182.n11 a_10732_182.n10 13.494
R3822 a_10732_182.t0 a_10732_182.n0 8.137
R3823 a_10732_182.t0 a_10732_182.n3 5.727
R3824 a_10732_182.n9 a_10732_182.n8 1.435
R3825 a_13322_182.n10 a_13322_182.n8 82.852
R3826 a_13322_182.n11 a_13322_182.n0 49.6
R3827 a_13322_182.n7 a_13322_182.n6 32.833
R3828 a_13322_182.n8 a_13322_182.t1 32.416
R3829 a_13322_182.n10 a_13322_182.n9 27.2
R3830 a_13322_182.n3 a_13322_182.n2 23.284
R3831 a_13322_182.n11 a_13322_182.n10 22.4
R3832 a_13322_182.n7 a_13322_182.n4 19.017
R3833 a_13322_182.n6 a_13322_182.n5 13.494
R3834 a_13322_182.t1 a_13322_182.n1 7.04
R3835 a_13322_182.t1 a_13322_182.n3 5.727
R3836 a_13322_182.n8 a_13322_182.n7 1.435
R3837 a_17723_182.n2 a_17723_182.n0 362.371
R3838 a_17723_182.n2 a_17723_182.n1 15.218
R3839 a_17723_182.n0 a_17723_182.t1 14.282
R3840 a_17723_182.n0 a_17723_182.t0 14.282
R3841 a_17723_182.n3 a_17723_182.n2 12.014
R3842 a_3924_182.n8 a_3924_182.n6 96.467
R3843 a_3924_182.n3 a_3924_182.n1 44.628
R3844 a_3924_182.t0 a_3924_182.n8 32.417
R3845 a_3924_182.n3 a_3924_182.n2 23.284
R3846 a_3924_182.n6 a_3924_182.n5 22.349
R3847 a_3924_182.t0 a_3924_182.n10 20.241
R3848 a_3924_182.n10 a_3924_182.n9 13.494
R3849 a_3924_182.n6 a_3924_182.n4 8.443
R3850 a_3924_182.t0 a_3924_182.n0 8.137
R3851 a_3924_182.t0 a_3924_182.n3 5.727
R3852 a_3924_182.n8 a_3924_182.n7 1.435
R3853 a_7216_73.t0 a_7216_73.n1 34.62
R3854 a_7216_73.t0 a_7216_73.n0 8.137
R3855 a_7216_73.t0 a_7216_73.n2 4.69
R3856 a_7321_1004.n3 a_7321_1004.t5 512.525
R3857 a_7321_1004.n3 a_7321_1004.t6 371.139
R3858 a_7321_1004.n4 a_7321_1004.t7 271.162
R3859 a_7321_1004.n7 a_7321_1004.n5 200.608
R3860 a_7321_1004.n4 a_7321_1004.n3 172.76
R3861 a_7321_1004.n5 a_7321_1004.n2 162.547
R3862 a_7321_1004.n5 a_7321_1004.n4 153.315
R3863 a_7321_1004.n2 a_7321_1004.n1 76.002
R3864 a_7321_1004.n7 a_7321_1004.n6 15.218
R3865 a_7321_1004.n0 a_7321_1004.t0 14.282
R3866 a_7321_1004.n0 a_7321_1004.t1 14.282
R3867 a_7321_1004.n1 a_7321_1004.t3 14.282
R3868 a_7321_1004.n1 a_7321_1004.t4 14.282
R3869 a_7321_1004.n2 a_7321_1004.n0 12.85
R3870 a_7321_1004.n8 a_7321_1004.n7 12.014
R3871 a_15652_73.n1 a_15652_73.n0 32.249
R3872 a_15652_73.t0 a_15652_73.n5 7.911
R3873 a_15652_73.n4 a_15652_73.n2 4.032
R3874 a_15652_73.n4 a_15652_73.n3 3.644
R3875 a_15652_73.t0 a_15652_73.n1 2.534
R3876 a_15652_73.t0 a_15652_73.n4 1.099
R3877 a_14986_73.t0 a_14986_73.n1 34.62
R3878 a_14986_73.t0 a_14986_73.n0 8.137
R3879 a_14986_73.t0 a_14986_73.n2 4.69
R3880 a_11694_182.n10 a_11694_182.n8 82.852
R3881 a_11694_182.n7 a_11694_182.n6 32.833
R3882 a_11694_182.n8 a_11694_182.t1 32.416
R3883 a_11694_182.n10 a_11694_182.n9 27.2
R3884 a_11694_182.n11 a_11694_182.n0 23.498
R3885 a_11694_182.n3 a_11694_182.n2 23.284
R3886 a_11694_182.n11 a_11694_182.n10 22.4
R3887 a_11694_182.n7 a_11694_182.n4 19.017
R3888 a_11694_182.n6 a_11694_182.n5 13.494
R3889 a_11694_182.t1 a_11694_182.n1 7.04
R3890 a_11694_182.t1 a_11694_182.n3 5.727
R3891 a_11694_182.n8 a_11694_182.n7 1.435
R3892 a_9104_182.n9 a_9104_182.n7 82.852
R3893 a_9104_182.n3 a_9104_182.n1 44.628
R3894 a_9104_182.t0 a_9104_182.n9 32.417
R3895 a_9104_182.n7 a_9104_182.n6 27.2
R3896 a_9104_182.n5 a_9104_182.n4 23.498
R3897 a_9104_182.n3 a_9104_182.n2 23.284
R3898 a_9104_182.n7 a_9104_182.n5 22.4
R3899 a_9104_182.t0 a_9104_182.n11 20.241
R3900 a_9104_182.n11 a_9104_182.n10 13.494
R3901 a_9104_182.t0 a_9104_182.n0 8.137
R3902 a_9104_182.t0 a_9104_182.n3 5.727
R3903 a_9104_182.n9 a_9104_182.n8 1.435
R3904 a_1053_75.n1 a_1053_75.n0 25.576
R3905 a_1053_75.n3 a_1053_75.n2 9.111
R3906 a_1053_75.n7 a_1053_75.n6 2.455
R3907 a_1053_75.n5 a_1053_75.n3 1.964
R3908 a_1053_75.n5 a_1053_75.n4 1.964
R3909 a_1053_75.t0 a_1053_75.n1 1.871
R3910 a_1053_75.n7 a_1053_75.n5 0.636
R3911 a_1053_75.t0 a_1053_75.n7 0.246
R3912 a_2962_182.n10 a_2962_182.n8 82.852
R3913 a_2962_182.n11 a_2962_182.n0 49.6
R3914 a_2962_182.n7 a_2962_182.n6 32.833
R3915 a_2962_182.n8 a_2962_182.t1 32.416
R3916 a_2962_182.n10 a_2962_182.n9 27.2
R3917 a_2962_182.n3 a_2962_182.n2 23.284
R3918 a_2962_182.n11 a_2962_182.n10 22.4
R3919 a_2962_182.n7 a_2962_182.n4 19.017
R3920 a_2962_182.n6 a_2962_182.n5 13.494
R3921 a_2962_182.t1 a_2962_182.n1 7.04
R3922 a_2962_182.t1 a_2962_182.n3 5.727
R3923 a_2962_182.n8 a_2962_182.n7 1.435
R3924 a_16984_73.t0 a_16984_73.n1 34.62
R3925 a_16984_73.t0 a_16984_73.n0 8.137
R3926 a_16984_73.t0 a_16984_73.n2 4.69
R3927 a_11413_75.n5 a_11413_75.n4 19.724
R3928 a_11413_75.t0 a_11413_75.n3 11.595
R3929 a_11413_75.t0 a_11413_75.n5 9.207
R3930 a_11413_75.n2 a_11413_75.n1 2.455
R3931 a_11413_75.n2 a_11413_75.n0 1.32
R3932 a_11413_75.t0 a_11413_75.n2 0.246
R3933 a_8142_182.n10 a_8142_182.n8 82.852
R3934 a_8142_182.n7 a_8142_182.n6 32.833
R3935 a_8142_182.n8 a_8142_182.t1 32.416
R3936 a_8142_182.n10 a_8142_182.n9 27.2
R3937 a_8142_182.n11 a_8142_182.n0 23.498
R3938 a_8142_182.n3 a_8142_182.n2 23.284
R3939 a_8142_182.n11 a_8142_182.n10 22.4
R3940 a_8142_182.n7 a_8142_182.n4 19.017
R3941 a_8142_182.n6 a_8142_182.n5 13.494
R3942 a_8142_182.t1 a_8142_182.n1 7.04
R3943 a_8142_182.t1 a_8142_182.n3 5.727
R3944 a_8142_182.n8 a_8142_182.n7 1.435
R3945 a_12396_73.n12 a_12396_73.n11 26.811
R3946 a_12396_73.n6 a_12396_73.n5 24.977
R3947 a_12396_73.n2 a_12396_73.n1 24.877
R3948 a_12396_73.t0 a_12396_73.n2 12.677
R3949 a_12396_73.t0 a_12396_73.n3 11.595
R3950 a_12396_73.t1 a_12396_73.n8 8.137
R3951 a_12396_73.t0 a_12396_73.n4 7.273
R3952 a_12396_73.t0 a_12396_73.n0 6.109
R3953 a_12396_73.t1 a_12396_73.n7 4.864
R3954 a_12396_73.t0 a_12396_73.n12 2.074
R3955 a_12396_73.n7 a_12396_73.n6 1.13
R3956 a_12396_73.n12 a_12396_73.t1 0.937
R3957 a_12396_73.t1 a_12396_73.n10 0.804
R3958 a_12396_73.n10 a_12396_73.n9 0.136
R3959 a_10451_75.n5 a_10451_75.n4 19.724
R3960 a_10451_75.t0 a_10451_75.n3 11.595
R3961 a_10451_75.t0 a_10451_75.n5 9.207
R3962 a_10451_75.n2 a_10451_75.n1 2.455
R3963 a_10451_75.n2 a_10451_75.n0 1.32
R3964 a_10451_75.t0 a_10451_75.n2 0.246
R3965 a_8823_75.n5 a_8823_75.n4 19.724
R3966 a_8823_75.t0 a_8823_75.n3 11.595
R3967 a_8823_75.t0 a_8823_75.n5 9.207
R3968 a_8823_75.n2 a_8823_75.n1 2.455
R3969 a_8823_75.n2 a_8823_75.n0 1.32
R3970 a_8823_75.t0 a_8823_75.n2 0.246
R3971 a_7861_75.n1 a_7861_75.n0 25.576
R3972 a_7861_75.n3 a_7861_75.n2 9.111
R3973 a_7861_75.n7 a_7861_75.n6 2.455
R3974 a_7861_75.n5 a_7861_75.n3 1.964
R3975 a_7861_75.n5 a_7861_75.n4 1.964
R3976 a_7861_75.t0 a_7861_75.n1 1.871
R3977 a_7861_75.n7 a_7861_75.n5 0.636
R3978 a_7861_75.t0 a_7861_75.n7 0.246
C6 VPB VNB 66.83fF
C7 a_7861_75.n0 VNB 0.09fF
C8 a_7861_75.n1 VNB 0.10fF
C9 a_7861_75.n2 VNB 0.05fF
C10 a_7861_75.n3 VNB 0.03fF
C11 a_7861_75.n4 VNB 0.04fF
C12 a_7861_75.n5 VNB 0.03fF
C13 a_7861_75.n6 VNB 0.04fF
C14 a_8823_75.n0 VNB 0.10fF
C15 a_8823_75.n1 VNB 0.04fF
C16 a_8823_75.n2 VNB 0.03fF
C17 a_8823_75.n3 VNB 0.07fF
C18 a_8823_75.n4 VNB 0.08fF
C19 a_8823_75.n5 VNB 0.06fF
C20 a_10451_75.n0 VNB 0.10fF
C21 a_10451_75.n1 VNB 0.04fF
C22 a_10451_75.n2 VNB 0.03fF
C23 a_10451_75.n3 VNB 0.07fF
C24 a_10451_75.n4 VNB 0.08fF
C25 a_10451_75.n5 VNB 0.06fF
C26 a_12396_73.n0 VNB 0.02fF
C27 a_12396_73.n1 VNB 0.10fF
C28 a_12396_73.n2 VNB 0.06fF
C29 a_12396_73.n3 VNB 0.06fF
C30 a_12396_73.n4 VNB 0.00fF
C31 a_12396_73.n5 VNB 0.04fF
C32 a_12396_73.n6 VNB 0.05fF
C33 a_12396_73.n7 VNB 0.02fF
C34 a_12396_73.n8 VNB 0.05fF
C35 a_12396_73.n9 VNB 0.08fF
C36 a_12396_73.n10 VNB 0.17fF
C37 a_12396_73.t1 VNB 0.23fF
C38 a_12396_73.n11 VNB 0.09fF
C39 a_12396_73.n12 VNB 0.00fF
C40 a_8142_182.n0 VNB 0.02fF
C41 a_8142_182.n1 VNB 0.09fF
C42 a_8142_182.n2 VNB 0.13fF
C43 a_8142_182.n3 VNB 0.11fF
C44 a_8142_182.t1 VNB 0.30fF
C45 a_8142_182.n4 VNB 0.09fF
C46 a_8142_182.n5 VNB 0.06fF
C47 a_8142_182.n6 VNB 0.01fF
C48 a_8142_182.n7 VNB 0.03fF
C49 a_8142_182.n8 VNB 0.11fF
C50 a_8142_182.n9 VNB 0.02fF
C51 a_8142_182.n10 VNB 0.05fF
C52 a_8142_182.n11 VNB 0.03fF
C53 a_11413_75.n0 VNB 0.10fF
C54 a_11413_75.n1 VNB 0.04fF
C55 a_11413_75.n2 VNB 0.03fF
C56 a_11413_75.n3 VNB 0.07fF
C57 a_11413_75.n4 VNB 0.08fF
C58 a_11413_75.n5 VNB 0.06fF
C59 a_16984_73.n0 VNB 0.06fF
C60 a_16984_73.n1 VNB 0.13fF
C61 a_16984_73.n2 VNB 0.04fF
C62 a_2962_182.n0 VNB 0.02fF
C63 a_2962_182.n1 VNB 0.09fF
C64 a_2962_182.n2 VNB 0.13fF
C65 a_2962_182.n3 VNB 0.11fF
C66 a_2962_182.t1 VNB 0.30fF
C67 a_2962_182.n4 VNB 0.09fF
C68 a_2962_182.n5 VNB 0.06fF
C69 a_2962_182.n6 VNB 0.01fF
C70 a_2962_182.n7 VNB 0.03fF
C71 a_2962_182.n8 VNB 0.11fF
C72 a_2962_182.n9 VNB 0.02fF
C73 a_2962_182.n10 VNB 0.05fF
C74 a_2962_182.n11 VNB 0.02fF
C75 a_1053_75.n0 VNB 0.09fF
C76 a_1053_75.n1 VNB 0.10fF
C77 a_1053_75.n2 VNB 0.05fF
C78 a_1053_75.n3 VNB 0.03fF
C79 a_1053_75.n4 VNB 0.04fF
C80 a_1053_75.n5 VNB 0.03fF
C81 a_1053_75.n6 VNB 0.04fF
C82 a_9104_182.n0 VNB 0.07fF
C83 a_9104_182.n1 VNB 0.09fF
C84 a_9104_182.n2 VNB 0.13fF
C85 a_9104_182.n3 VNB 0.11fF
C86 a_9104_182.n4 VNB 0.02fF
C87 a_9104_182.n5 VNB 0.03fF
C88 a_9104_182.n6 VNB 0.02fF
C89 a_9104_182.n7 VNB 0.05fF
C90 a_9104_182.n8 VNB 0.03fF
C91 a_9104_182.n9 VNB 0.11fF
C92 a_9104_182.n10 VNB 0.06fF
C93 a_9104_182.n11 VNB 0.01fF
C94 a_9104_182.t0 VNB 0.33fF
C95 a_11694_182.n0 VNB 0.02fF
C96 a_11694_182.n1 VNB 0.09fF
C97 a_11694_182.n2 VNB 0.13fF
C98 a_11694_182.n3 VNB 0.11fF
C99 a_11694_182.t1 VNB 0.30fF
C100 a_11694_182.n4 VNB 0.09fF
C101 a_11694_182.n5 VNB 0.06fF
C102 a_11694_182.n6 VNB 0.01fF
C103 a_11694_182.n7 VNB 0.03fF
C104 a_11694_182.n8 VNB 0.11fF
C105 a_11694_182.n9 VNB 0.02fF
C106 a_11694_182.n10 VNB 0.05fF
C107 a_11694_182.n11 VNB 0.03fF
C108 a_14986_73.n0 VNB 0.05fF
C109 a_14986_73.n1 VNB 0.12fF
C110 a_14986_73.n2 VNB 0.04fF
C111 a_15652_73.n0 VNB 0.11fF
C112 a_15652_73.n1 VNB 0.09fF
C113 a_15652_73.n2 VNB 0.08fF
C114 a_15652_73.n3 VNB 0.02fF
C115 a_15652_73.n4 VNB 0.01fF
C116 a_15652_73.n5 VNB 0.06fF
C117 a_7321_1004.n0 VNB 0.61fF
C118 a_7321_1004.n1 VNB 0.72fF
C119 a_7321_1004.n2 VNB 0.36fF
C120 a_7321_1004.n3 VNB 0.40fF
C121 a_7321_1004.n4 VNB 0.74fF
C122 a_7321_1004.n5 VNB 0.69fF
C123 a_7321_1004.n6 VNB 0.10fF
C124 a_7321_1004.n7 VNB 0.31fF
C125 a_7321_1004.n8 VNB 0.05fF
C126 a_7216_73.n0 VNB 0.05fF
C127 a_7216_73.n1 VNB 0.12fF
C128 a_7216_73.n2 VNB 0.04fF
C129 a_3924_182.n0 VNB 0.07fF
C130 a_3924_182.n1 VNB 0.09fF
C131 a_3924_182.n2 VNB 0.13fF
C132 a_3924_182.n3 VNB 0.11fF
C133 a_3924_182.n4 VNB 0.02fF
C134 a_3924_182.n5 VNB 0.03fF
C135 a_3924_182.n6 VNB 0.06fF
C136 a_3924_182.n7 VNB 0.03fF
C137 a_3924_182.n8 VNB 0.12fF
C138 a_3924_182.n9 VNB 0.06fF
C139 a_3924_182.n10 VNB 0.01fF
C140 a_3924_182.t0 VNB 0.33fF
C141 a_17723_182.n0 VNB 1.03fF
C142 a_17723_182.n1 VNB 0.09fF
C143 a_17723_182.n2 VNB 0.49fF
C144 a_17723_182.n3 VNB 0.05fF
C145 a_13322_182.n0 VNB 0.02fF
C146 a_13322_182.n1 VNB 0.09fF
C147 a_13322_182.n2 VNB 0.13fF
C148 a_13322_182.n3 VNB 0.11fF
C149 a_13322_182.t1 VNB 0.30fF
C150 a_13322_182.n4 VNB 0.09fF
C151 a_13322_182.n5 VNB 0.06fF
C152 a_13322_182.n6 VNB 0.01fF
C153 a_13322_182.n7 VNB 0.03fF
C154 a_13322_182.n8 VNB 0.11fF
C155 a_13322_182.n9 VNB 0.02fF
C156 a_13322_182.n10 VNB 0.05fF
C157 a_13322_182.n11 VNB 0.02fF
C158 a_10732_182.n0 VNB 0.07fF
C159 a_10732_182.n1 VNB 0.09fF
C160 a_10732_182.n2 VNB 0.13fF
C161 a_10732_182.n3 VNB 0.11fF
C162 a_10732_182.n4 VNB 0.02fF
C163 a_10732_182.n5 VNB 0.03fF
C164 a_10732_182.n6 VNB 0.02fF
C165 a_10732_182.n7 VNB 0.05fF
C166 a_10732_182.n8 VNB 0.03fF
C167 a_10732_182.n9 VNB 0.11fF
C168 a_10732_182.n10 VNB 0.06fF
C169 a_10732_182.n11 VNB 0.01fF
C170 a_10732_182.t0 VNB 0.33fF
C171 a_1334_182.n0 VNB 0.02fF
C172 a_1334_182.n1 VNB 0.09fF
C173 a_1334_182.n2 VNB 0.13fF
C174 a_1334_182.n3 VNB 0.11fF
C175 a_1334_182.t1 VNB 0.30fF
C176 a_1334_182.n4 VNB 0.09fF
C177 a_1334_182.n5 VNB 0.06fF
C178 a_1334_182.n6 VNB 0.01fF
C179 a_1334_182.n7 VNB 0.03fF
C180 a_1334_182.n8 VNB 0.11fF
C181 a_1334_182.n9 VNB 0.02fF
C182 a_1334_182.n10 VNB 0.05fF
C183 a_1334_182.n11 VNB 0.03fF
C184 a_2681_75.n0 VNB 0.20fF
C185 a_2681_75.n1 VNB 0.04fF
C186 a_2681_75.n2 VNB 0.01fF
C187 a_2681_75.n3 VNB 0.08fF
C188 a_2681_75.n4 VNB 0.06fF
C189 a_2681_75.n5 VNB 0.07fF
C190 a_14003_75.n0 VNB 0.10fF
C191 a_14003_75.n1 VNB 0.04fF
C192 a_14003_75.n2 VNB 0.03fF
C193 a_14003_75.n3 VNB 0.07fF
C194 a_14003_75.n4 VNB 0.08fF
C195 a_14003_75.n5 VNB 0.06fF
C196 a_2036_73.n0 VNB 0.02fF
C197 a_2036_73.n1 VNB 0.10fF
C198 a_2036_73.n2 VNB 0.06fF
C199 a_2036_73.n3 VNB 0.06fF
C200 a_2036_73.n4 VNB 0.00fF
C201 a_2036_73.n5 VNB 0.04fF
C202 a_2036_73.n6 VNB 0.05fF
C203 a_2036_73.n7 VNB 0.02fF
C204 a_2036_73.n8 VNB 0.05fF
C205 a_2036_73.n9 VNB 0.08fF
C206 a_2036_73.n10 VNB 0.17fF
C207 a_2036_73.t1 VNB 0.23fF
C208 a_2036_73.n11 VNB 0.09fF
C209 a_2036_73.n12 VNB 0.00fF
C210 a_4626_73.n0 VNB 0.02fF
C211 a_4626_73.n1 VNB 0.10fF
C212 a_4626_73.n2 VNB 0.06fF
C213 a_4626_73.n3 VNB 0.06fF
C214 a_4626_73.n4 VNB 0.00fF
C215 a_4626_73.n5 VNB 0.04fF
C216 a_4626_73.n6 VNB 0.05fF
C217 a_4626_73.n7 VNB 0.02fF
C218 a_4626_73.n8 VNB 0.05fF
C219 a_4626_73.n9 VNB 0.08fF
C220 a_4626_73.n10 VNB 0.17fF
C221 a_4626_73.t1 VNB 0.23fF
C222 a_4626_73.n11 VNB 0.09fF
C223 a_4626_73.n12 VNB 0.00fF
C224 a_9009_1004.n0 VNB 0.04fF
C225 a_9009_1004.n1 VNB 0.56fF
C226 a_9009_1004.n2 VNB 0.56fF
C227 a_9009_1004.n3 VNB 0.66fF
C228 a_9009_1004.n4 VNB 0.21fF
C229 a_9009_1004.n5 VNB 0.30fF
C230 a_9009_1004.n6 VNB 0.37fF
C231 a_9009_1004.n7 VNB 0.59fF
C232 a_9009_1004.n8 VNB 0.65fF
C233 a_9009_1004.n9 VNB 0.04fF
C234 a_9009_1004.n10 VNB 0.33fF
C235 a_9009_1004.n11 VNB 0.06fF
C236 a_2141_1004.n0 VNB 0.04fF
C237 a_2141_1004.n1 VNB 0.55fF
C238 a_2141_1004.n2 VNB 0.65fF
C239 a_2141_1004.n3 VNB 0.33fF
C240 a_2141_1004.n4 VNB 0.36fF
C241 a_2141_1004.n5 VNB 0.67fF
C242 a_2141_1004.n6 VNB 0.62fF
C243 a_2141_1004.n7 VNB 0.04fF
C244 a_2141_1004.n8 VNB 0.29fF
C245 a_2141_1004.n9 VNB 0.06fF
C246 a_16318_73.n0 VNB 0.13fF
C247 a_16318_73.n1 VNB 0.13fF
C248 a_16318_73.n2 VNB 0.14fF
C249 a_5552_182.n0 VNB 0.02fF
C250 a_5552_182.n1 VNB 0.09fF
C251 a_5552_182.n2 VNB 0.13fF
C252 a_5552_182.n3 VNB 0.11fF
C253 a_5552_182.t1 VNB 0.30fF
C254 a_5552_182.n4 VNB 0.09fF
C255 a_5552_182.n5 VNB 0.06fF
C256 a_5552_182.n6 VNB 0.01fF
C257 a_5552_182.n7 VNB 0.03fF
C258 a_5552_182.n8 VNB 0.11fF
C259 a_5552_182.n9 VNB 0.02fF
C260 a_5552_182.n10 VNB 0.05fF
C261 a_5552_182.n11 VNB 0.02fF
C262 a_5271_75.n0 VNB 0.20fF
C263 a_5271_75.n1 VNB 0.04fF
C264 a_5271_75.n2 VNB 0.01fF
C265 a_5271_75.n3 VNB 0.08fF
C266 a_5271_75.n4 VNB 0.06fF
C267 a_5271_75.n5 VNB 0.07fF
C268 a_372_182.n0 VNB 0.07fF
C269 a_372_182.n1 VNB 0.09fF
C270 a_372_182.n2 VNB 0.13fF
C271 a_372_182.n3 VNB 0.11fF
C272 a_372_182.n4 VNB 0.02fF
C273 a_372_182.n5 VNB 0.03fF
C274 a_372_182.n6 VNB 0.06fF
C275 a_372_182.n7 VNB 0.03fF
C276 a_372_182.n8 VNB 0.12fF
C277 a_372_182.n9 VNB 0.06fF
C278 a_372_182.n10 VNB 0.01fF
C279 a_372_182.t0 VNB 0.33fF
C280 a_91_75.n0 VNB 0.09fF
C281 a_91_75.n1 VNB 0.09fF
C282 a_91_75.n2 VNB 0.04fF
C283 a_91_75.n3 VNB 0.03fF
C284 a_91_75.n4 VNB 0.04fF
C285 a_91_75.n5 VNB 0.11fF
C286 a_91_75.n6 VNB 0.04fF
C287 a_3643_75.n0 VNB 0.20fF
C288 a_3643_75.n1 VNB 0.04fF
C289 a_3643_75.n2 VNB 0.01fF
C290 a_3643_75.n3 VNB 0.08fF
C291 a_3643_75.n4 VNB 0.06fF
C292 a_3643_75.n5 VNB 0.07fF
C293 a_15932_181.n0 VNB 0.04fF
C294 a_15932_181.n1 VNB 0.38fF
C295 a_15932_181.n2 VNB 0.47fF
C296 a_15932_181.n3 VNB 0.22fF
C297 a_15932_181.n4 VNB 0.24fF
C298 a_15932_181.t7 VNB 0.49fF
C299 a_15932_181.n5 VNB 0.49fF
C300 a_15932_181.n6 VNB 0.46fF
C301 a_15932_181.n7 VNB 0.03fF
C302 a_15932_181.n8 VNB 0.05fF
C303 a_15932_181.n9 VNB 0.03fF
C304 a_15932_181.n10 VNB 0.09fF
C305 a_15932_181.n11 VNB 0.03fF
C306 a_15932_181.n12 VNB 0.05fF
C307 a_15932_181.n13 VNB 0.03fF
C308 a_15932_181.n14 VNB 0.09fF
C309 a_15932_181.n15 VNB 0.98fF
C310 a_15932_181.n16 VNB 0.27fF
C311 a_15932_181.n17 VNB 0.03fF
C312 a_15932_181.n18 VNB 0.05fF
C313 a_15932_181.n19 VNB 0.04fF
C314 a_599_943.n0 VNB 0.04fF
C315 a_599_943.n1 VNB 0.59fF
C316 a_599_943.n2 VNB 0.59fF
C317 a_599_943.n3 VNB 0.69fF
C318 a_599_943.n4 VNB 0.22fF
C319 a_599_943.n5 VNB 0.35fF
C320 a_599_943.n6 VNB 0.43fF
C321 a_599_943.n7 VNB 0.42fF
C322 a_599_943.n8 VNB 0.43fF
C323 a_599_943.t12 VNB 0.57fF
C324 a_599_943.n9 VNB 0.42fF
C325 a_599_943.n10 VNB 1.37fF
C326 a_599_943.n11 VNB 0.49fF
C327 a_599_943.n12 VNB 0.04fF
C328 a_599_943.n13 VNB 0.31fF
C329 a_599_943.n14 VNB 0.06fF
C330 a_13041_75.n0 VNB 0.20fF
C331 a_13041_75.n1 VNB 0.04fF
C332 a_13041_75.n2 VNB 0.01fF
C333 a_13041_75.n3 VNB 0.03fF
C334 a_13041_75.n4 VNB 0.05fF
C335 a_13041_75.n5 VNB 0.09fF
C336 a_13041_75.n6 VNB 0.07fF
C337 a_14284_182.n0 VNB 0.07fF
C338 a_14284_182.n1 VNB 0.09fF
C339 a_14284_182.n2 VNB 0.13fF
C340 a_14284_182.n3 VNB 0.11fF
C341 a_14284_182.n4 VNB 0.02fF
C342 a_14284_182.n5 VNB 0.03fF
C343 a_14284_182.n6 VNB 0.02fF
C344 a_14284_182.n7 VNB 0.05fF
C345 a_14284_182.n8 VNB 0.03fF
C346 a_14284_182.n9 VNB 0.11fF
C347 a_14284_182.n10 VNB 0.06fF
C348 a_14284_182.n11 VNB 0.01fF
C349 a_14284_182.t0 VNB 0.33fF
C350 a_10637_1004.n0 VNB 0.07fF
C351 a_10637_1004.n1 VNB 0.91fF
C352 a_10637_1004.n2 VNB 0.91fF
C353 a_10637_1004.n3 VNB 1.07fF
C354 a_10637_1004.n4 VNB 0.34fF
C355 a_10637_1004.n5 VNB 0.49fF
C356 a_10637_1004.n6 VNB 0.54fF
C357 a_10637_1004.n7 VNB 1.00fF
C358 a_10637_1004.n8 VNB 0.54fF
C359 a_10637_1004.n9 VNB 0.80fF
C360 a_10637_1004.n10 VNB 4.00fF
C361 a_10637_1004.n11 VNB 0.76fF
C362 a_10637_1004.n12 VNB 0.06fF
C363 a_10637_1004.n13 VNB 0.53fF
C364 a_10637_1004.n14 VNB 0.09fF
C365 a_15757_1005.n0 VNB 0.40fF
C366 a_15757_1005.n1 VNB 0.32fF
C367 a_15757_1005.n2 VNB 0.23fF
C368 a_15757_1005.n3 VNB 0.62fF
C369 a_15757_1005.n4 VNB 0.28fF
C370 a_15757_1005.n5 VNB 0.36fF
C371 a_16421_1005.n0 VNB 0.29fF
C372 a_16421_1005.n1 VNB 0.28fF
C373 a_16421_1005.n2 VNB 0.36fF
C374 a_16421_1005.n3 VNB 0.25fF
C375 a_16421_1005.n4 VNB 0.57fF
C376 a_16421_1005.n5 VNB 0.20fF
C377 a_4151_943.n0 VNB 1.21fF
C378 a_4151_943.n1 VNB 0.90fF
C379 a_4151_943.n2 VNB 1.06fF
C380 a_4151_943.n3 VNB 1.32fF
C381 a_4151_943.t6 VNB 1.00fF
C382 a_4151_943.n4 VNB 0.79fF
C383 a_4151_943.n5 VNB 4.66fF
C384 a_4151_943.n6 VNB 0.96fF
C385 a_4151_943.t12 VNB 1.12fF
C386 a_4151_943.n7 VNB 0.83fF
C387 a_4151_943.n8 VNB 19.51fF
C388 a_4151_943.n9 VNB 0.09fF
C389 a_4151_943.n10 VNB 0.12fF
C390 a_4151_943.n11 VNB 0.08fF
C391 a_4151_943.n12 VNB 0.57fF
C392 a_4151_943.n13 VNB 0.96fF
C393 a_4151_943.n14 VNB 0.80fF
C394 a_4151_943.n15 VNB 1.44fF
C395 a_277_1004.n0 VNB 0.79fF
C396 a_277_1004.n1 VNB 0.79fF
C397 a_277_1004.n2 VNB 0.93fF
C398 a_277_1004.n3 VNB 0.29fF
C399 a_277_1004.n4 VNB 0.42fF
C400 a_277_1004.n5 VNB 0.47fF
C401 a_277_1004.n6 VNB 0.87fF
C402 a_277_1004.n7 VNB 0.47fF
C403 a_277_1004.n8 VNB 0.70fF
C404 a_277_1004.n9 VNB 3.48fF
C405 a_277_1004.n10 VNB 0.67fF
C406 a_277_1004.n11 VNB 0.12fF
C407 a_277_1004.n12 VNB 0.45fF
C408 a_277_1004.n13 VNB 0.07fF
C409 a_147_159.n0 VNB 0.37fF
C410 a_147_159.t20 VNB 0.73fF
C411 a_147_159.n1 VNB 0.48fF
C412 a_147_159.n2 VNB 0.42fF
C413 a_147_159.n3 VNB 0.50fF
C414 a_147_159.n4 VNB 0.40fF
C415 a_147_159.n5 VNB 0.69fF
C416 a_147_159.n6 VNB 0.69fF
C417 a_147_159.n7 VNB 0.81fF
C418 a_147_159.n8 VNB 0.25fF
C419 a_147_159.n9 VNB 0.33fF
C420 a_147_159.n10 VNB 0.05fF
C421 a_147_159.n11 VNB 0.07fF
C422 a_147_159.n12 VNB 0.45fF
C423 a_147_159.n13 VNB 0.60fF
C424 a_147_159.n14 VNB 0.71fF
C425 a_147_159.n15 VNB 0.37fF
C426 a_147_159.t21 VNB 0.73fF
C427 a_147_159.n16 VNB 0.48fF
C428 a_147_159.n17 VNB 0.37fF
C429 a_147_159.n18 VNB 0.71fF
C430 a_147_159.n19 VNB 2.70fF
C431 a_147_159.n20 VNB 1.10fF
C432 a_147_159.n21 VNB 0.05fF
C433 a_147_159.n22 VNB 0.07fF
C434 a_147_159.n23 VNB 0.04fF
C435 a_147_159.n24 VNB 0.44fF
C436 a_147_159.n25 VNB 0.57fF
C437 a_147_159.n26 VNB 0.69fF
C438 a_147_159.n27 VNB 0.81fF
C439 a_147_159.n28 VNB 0.25fF
C440 a_147_159.n29 VNB 0.33fF
C441 a_147_159.n30 VNB 0.69fF
C442 a_5457_1004.n0 VNB 0.07fF
C443 a_5457_1004.n1 VNB 0.88fF
C444 a_5457_1004.n2 VNB 0.88fF
C445 a_5457_1004.n3 VNB 1.04fF
C446 a_5457_1004.n4 VNB 0.33fF
C447 a_5457_1004.n5 VNB 0.47fF
C448 a_5457_1004.n6 VNB 0.52fF
C449 a_5457_1004.n7 VNB 0.98fF
C450 a_5457_1004.n8 VNB 0.52fF
C451 a_5457_1004.n9 VNB 0.78fF
C452 a_5457_1004.n10 VNB 3.88fF
C453 a_5457_1004.n11 VNB 0.73fF
C454 a_5457_1004.n12 VNB 0.06fF
C455 a_5457_1004.n13 VNB 0.52fF
C456 a_5457_1004.n14 VNB 0.09fF
C457 a_5779_943.n0 VNB 0.74fF
C458 a_5779_943.n1 VNB 0.74fF
C459 a_5779_943.n2 VNB 0.87fF
C460 a_5779_943.n3 VNB 0.27fF
C461 a_5779_943.n4 VNB 0.44fF
C462 a_5779_943.n5 VNB 0.54fF
C463 a_5779_943.n6 VNB 0.53fF
C464 a_5779_943.n7 VNB 0.54fF
C465 a_5779_943.t11 VNB 0.71fF
C466 a_5779_943.n8 VNB 0.53fF
C467 a_5779_943.n9 VNB 1.72fF
C468 a_5779_943.n10 VNB 0.63fF
C469 a_5779_943.n11 VNB 0.11fF
C470 a_5779_943.n12 VNB 0.38fF
C471 a_5779_943.n13 VNB 0.06fF
C472 a_6514_182.n0 VNB 0.02fF
C473 a_6514_182.n1 VNB 0.07fF
C474 a_6514_182.n2 VNB 0.13fF
C475 a_6514_182.n3 VNB 0.09fF
C476 a_6514_182.t1 VNB 0.25fF
C477 a_6514_182.n4 VNB 0.05fF
C478 a_6514_182.n5 VNB 0.06fF
C479 a_6514_182.n6 VNB 0.07fF
C480 a_6514_182.n7 VNB 0.07fF
C481 a_6514_182.n8 VNB 0.03fF
C482 a_6514_182.n9 VNB 0.01fF
C483 a_6514_182.n10 VNB 0.11fF
C484 a_6514_182.n11 VNB 0.02fF
C485 a_6514_182.n12 VNB 0.05fF
C486 a_6514_182.n13 VNB 0.02fF
C487 a_6233_75.n0 VNB 0.20fF
C488 a_6233_75.n1 VNB 0.04fF
C489 a_6233_75.n2 VNB 0.01fF
C490 a_6233_75.n3 VNB 0.08fF
C491 a_6233_75.n4 VNB 0.06fF
C492 a_6233_75.n5 VNB 0.07fF
C493 a_9806_73.n0 VNB 0.02fF
C494 a_9806_73.n1 VNB 0.10fF
C495 a_9806_73.n2 VNB 0.07fF
C496 a_9806_73.n3 VNB 0.05fF
C497 a_9806_73.n4 VNB 0.00fF
C498 a_9806_73.n5 VNB 0.04fF
C499 a_9806_73.n6 VNB 0.05fF
C500 a_9806_73.n7 VNB 0.02fF
C501 a_9806_73.n8 VNB 0.05fF
C502 a_9806_73.n9 VNB 0.02fF
C503 a_9806_73.n10 VNB 0.08fF
C504 a_9806_73.n11 VNB 0.17fF
C505 a_9806_73.t1 VNB 0.23fF
C506 a_9806_73.n12 VNB 0.09fF
C507 a_9806_73.n13 VNB 0.00fF
C508 a_5327_159.n0 VNB 0.07fF
C509 a_5327_159.n1 VNB 0.94fF
C510 a_5327_159.n2 VNB 0.94fF
C511 a_5327_159.n3 VNB 1.11fF
C512 a_5327_159.n4 VNB 0.35fF
C513 a_5327_159.n5 VNB 0.45fF
C514 a_5327_159.n6 VNB 0.51fF
C515 a_5327_159.t7 VNB 1.00fF
C516 a_5327_159.n7 VNB 0.73fF
C517 a_5327_159.n8 VNB 0.51fF
C518 a_5327_159.t9 VNB 1.00fF
C519 a_5327_159.n9 VNB 0.66fF
C520 a_5327_159.n10 VNB 0.50fF
C521 a_5327_159.n11 VNB 0.97fF
C522 a_5327_159.n12 VNB 3.69fF
C523 a_5327_159.n13 VNB 2.91fF
C524 a_5327_159.n14 VNB 0.78fF
C525 a_5327_159.n15 VNB 0.06fF
C526 a_5327_159.n16 VNB 0.60fF
C527 a_5327_159.n17 VNB 0.09fF
C528 a_9331_943.n0 VNB 0.06fF
C529 a_9331_943.n1 VNB 0.78fF
C530 a_9331_943.n2 VNB 0.92fF
C531 a_9331_943.n3 VNB 0.47fF
C532 a_9331_943.n4 VNB 0.38fF
C533 a_9331_943.n5 VNB 0.43fF
C534 a_9331_943.n6 VNB 1.07fF
C535 a_9331_943.n7 VNB 0.79fF
C536 a_9331_943.n8 VNB 0.67fF
C537 a_9331_943.n9 VNB 0.51fF
C538 a_9331_943.n10 VNB 0.69fF
C539 a_9331_943.n11 VNB 3.13fF
C540 a_9331_943.n12 VNB 0.57fF
C541 a_9331_943.n13 VNB 0.56fF
C542 a_9331_943.n14 VNB 0.79fF
C543 a_9331_943.n15 VNB 0.79fF
C544 a_9331_943.n16 VNB 0.93fF
C545 a_9331_943.n17 VNB 0.29fF
C546 a_9331_943.n18 VNB 0.47fF
C547 a_9331_943.n19 VNB 0.06fF
C548 a_9331_943.n20 VNB 0.08fF
C549 a_9331_943.n21 VNB 0.05fF
C550 a_9331_943.n22 VNB 0.41fF
C551 a_9331_943.n23 VNB 0.65fF
C552 a_9331_943.n24 VNB 0.57fF
C553 a_9331_943.t22 VNB 0.76fF
C554 a_9331_943.n25 VNB 0.53fF
C555 a_9331_943.n26 VNB 0.78fF
C556 a_9331_943.n27 VNB 0.92fF
C557 a_9331_943.n28 VNB 0.47fF
C558 a_9331_943.n29 VNB 0.10fF
C559 a_9331_943.n30 VNB 0.04fF
C560 a_9331_943.n31 VNB 0.42fF
C561 a_9331_943.n32 VNB 0.65fF
C562 a_9331_943.n33 VNB 0.57fF
C563 a_9331_943.t25 VNB 0.76fF
C564 a_9331_943.n34 VNB 0.55fF
C565 a_9331_943.n35 VNB 1.50fF
C566 a_9331_943.n36 VNB 1.17fF
C567 a_9331_943.n37 VNB 0.91fF
C568 a_9331_943.n38 VNB 0.42fF
C569 a_9331_943.n39 VNB 0.42fF
C570 a_9331_943.n40 VNB 0.61fF
C571 a_9331_943.n41 VNB 0.05fF
C572 a_9331_943.n42 VNB 0.41fF
C573 a_9331_943.n43 VNB 0.08fF
C574 a_14511_943.n0 VNB 0.59fF
C575 a_14511_943.n1 VNB 0.32fF
C576 a_14511_943.n2 VNB 0.36fF
C577 a_14511_943.t12 VNB 0.64fF
C578 a_14511_943.n3 VNB 1.08fF
C579 a_14511_943.n4 VNB 0.76fF
C580 a_14511_943.t11 VNB 0.61fF
C581 a_14511_943.n5 VNB 0.34fF
C582 a_14511_943.n6 VNB 0.40fF
C583 a_14511_943.t5 VNB 0.61fF
C584 a_14511_943.n7 VNB 0.42fF
C585 a_14511_943.n8 VNB 1.27fF
C586 a_14511_943.n9 VNB 0.05fF
C587 a_14511_943.n10 VNB 0.06fF
C588 a_14511_943.n11 VNB 0.04fF
C589 a_14511_943.n12 VNB 0.35fF
C590 a_14511_943.n13 VNB 0.47fF
C591 a_14511_943.n14 VNB 0.32fF
C592 a_14511_943.n15 VNB 0.70fF
C593 VPB.n0 VNB 0.03fF
C594 VPB.n1 VNB 0.04fF
C595 VPB.n2 VNB 0.02fF
C596 VPB.n3 VNB 0.19fF
C597 VPB.n5 VNB 0.02fF
C598 VPB.n6 VNB 0.02fF
C599 VPB.n7 VNB 0.02fF
C600 VPB.n8 VNB 0.02fF
C601 VPB.n10 VNB 0.02fF
C602 VPB.n11 VNB 0.02fF
C603 VPB.n12 VNB 0.02fF
C604 VPB.n14 VNB 0.10fF
C605 VPB.n15 VNB 0.10fF
C606 VPB.n16 VNB 0.02fF
C607 VPB.n17 VNB 0.02fF
C608 VPB.n18 VNB 0.02fF
C609 VPB.n19 VNB 0.04fF
C610 VPB.n20 VNB 0.02fF
C611 VPB.n21 VNB 0.29fF
C612 VPB.n22 VNB 0.04fF
C613 VPB.n24 VNB 0.02fF
C614 VPB.n25 VNB 0.02fF
C615 VPB.n26 VNB 0.02fF
C616 VPB.n27 VNB 0.02fF
C617 VPB.n29 VNB 0.02fF
C618 VPB.n30 VNB 0.02fF
C619 VPB.n31 VNB 0.02fF
C620 VPB.n33 VNB 0.28fF
C621 VPB.n35 VNB 0.03fF
C622 VPB.n36 VNB 0.02fF
C623 VPB.n37 VNB 0.03fF
C624 VPB.n38 VNB 0.03fF
C625 VPB.n39 VNB 0.28fF
C626 VPB.n40 VNB 0.01fF
C627 VPB.n41 VNB 0.02fF
C628 VPB.n42 VNB 0.28fF
C629 VPB.n43 VNB 0.02fF
C630 VPB.n44 VNB 0.02fF
C631 VPB.n45 VNB 0.05fF
C632 VPB.n46 VNB 0.21fF
C633 VPB.n47 VNB 0.02fF
C634 VPB.n48 VNB 0.01fF
C635 VPB.n49 VNB 0.14fF
C636 VPB.n50 VNB 0.16fF
C637 VPB.n51 VNB 0.02fF
C638 VPB.n52 VNB 0.02fF
C639 VPB.n53 VNB 0.14fF
C640 VPB.n54 VNB 0.16fF
C641 VPB.n55 VNB 0.02fF
C642 VPB.n56 VNB 0.02fF
C643 VPB.n57 VNB 0.02fF
C644 VPB.n58 VNB 0.14fF
C645 VPB.n59 VNB 0.15fF
C646 VPB.n60 VNB 0.02fF
C647 VPB.n61 VNB 0.02fF
C648 VPB.n62 VNB 0.14fF
C649 VPB.n63 VNB 0.15fF
C650 VPB.n64 VNB 0.02fF
C651 VPB.n65 VNB 0.02fF
C652 VPB.n66 VNB 0.02fF
C653 VPB.n67 VNB 0.14fF
C654 VPB.n68 VNB 0.16fF
C655 VPB.n69 VNB 0.02fF
C656 VPB.n70 VNB 0.02fF
C657 VPB.n71 VNB 0.14fF
C658 VPB.n72 VNB 0.16fF
C659 VPB.n73 VNB 0.02fF
C660 VPB.n74 VNB 0.02fF
C661 VPB.n75 VNB 0.21fF
C662 VPB.n76 VNB 0.02fF
C663 VPB.n77 VNB 0.01fF
C664 VPB.n78 VNB 0.06fF
C665 VPB.n79 VNB 0.28fF
C666 VPB.n80 VNB 0.02fF
C667 VPB.n81 VNB 0.02fF
C668 VPB.n82 VNB 0.10fF
C669 VPB.n83 VNB 0.10fF
C670 VPB.n84 VNB 0.02fF
C671 VPB.n85 VNB 0.02fF
C672 VPB.n86 VNB 0.02fF
C673 VPB.n87 VNB 0.04fF
C674 VPB.n88 VNB 0.02fF
C675 VPB.n89 VNB 0.24fF
C676 VPB.n90 VNB 0.04fF
C677 VPB.n92 VNB 0.02fF
C678 VPB.n93 VNB 0.02fF
C679 VPB.n94 VNB 0.02fF
C680 VPB.n95 VNB 0.02fF
C681 VPB.n97 VNB 0.02fF
C682 VPB.n98 VNB 0.02fF
C683 VPB.n99 VNB 0.02fF
C684 VPB.n101 VNB 0.28fF
C685 VPB.n103 VNB 0.03fF
C686 VPB.n104 VNB 0.02fF
C687 VPB.n105 VNB 0.06fF
C688 VPB.n106 VNB 0.24fF
C689 VPB.n107 VNB 0.02fF
C690 VPB.n108 VNB 0.01fF
C691 VPB.n109 VNB 0.28fF
C692 VPB.n110 VNB 0.01fF
C693 VPB.n111 VNB 0.02fF
C694 VPB.n112 VNB 0.03fF
C695 VPB.n113 VNB 0.03fF
C696 VPB.n114 VNB 0.28fF
C697 VPB.n115 VNB 0.01fF
C698 VPB.n116 VNB 0.02fF
C699 VPB.n117 VNB 0.28fF
C700 VPB.n118 VNB 0.02fF
C701 VPB.n119 VNB 0.02fF
C702 VPB.n120 VNB 0.05fF
C703 VPB.n121 VNB 0.21fF
C704 VPB.n122 VNB 0.02fF
C705 VPB.n123 VNB 0.01fF
C706 VPB.n124 VNB 0.14fF
C707 VPB.n125 VNB 0.16fF
C708 VPB.n126 VNB 0.02fF
C709 VPB.n127 VNB 0.02fF
C710 VPB.n128 VNB 0.14fF
C711 VPB.n129 VNB 0.16fF
C712 VPB.n130 VNB 0.02fF
C713 VPB.n131 VNB 0.02fF
C714 VPB.n132 VNB 0.02fF
C715 VPB.n133 VNB 0.14fF
C716 VPB.n134 VNB 0.15fF
C717 VPB.n135 VNB 0.02fF
C718 VPB.n136 VNB 0.02fF
C719 VPB.n137 VNB 0.14fF
C720 VPB.n138 VNB 0.15fF
C721 VPB.n139 VNB 0.02fF
C722 VPB.n140 VNB 0.02fF
C723 VPB.n141 VNB 0.02fF
C724 VPB.n142 VNB 0.14fF
C725 VPB.n143 VNB 0.16fF
C726 VPB.n144 VNB 0.02fF
C727 VPB.n145 VNB 0.02fF
C728 VPB.n146 VNB 0.02fF
C729 VPB.n147 VNB 0.02fF
C730 VPB.n148 VNB 0.02fF
C731 VPB.n149 VNB 0.11fF
C732 VPB.n150 VNB 0.03fF
C733 VPB.n151 VNB 0.02fF
C734 VPB.n152 VNB 0.05fF
C735 VPB.n153 VNB 0.01fF
C736 VPB.n154 VNB 0.02fF
C737 VPB.n155 VNB 0.02fF
C738 VPB.n158 VNB 0.02fF
C739 VPB.n159 VNB 0.02fF
C740 VPB.n160 VNB 0.02fF
C741 VPB.n163 VNB 0.46fF
C742 VPB.n165 VNB 0.04fF
C743 VPB.n166 VNB 0.04fF
C744 VPB.n167 VNB 0.28fF
C745 VPB.n168 VNB 0.03fF
C746 VPB.n169 VNB 0.03fF
C747 VPB.n170 VNB 0.06fF
C748 VPB.n171 VNB 0.14fF
C749 VPB.n172 VNB 0.19fF
C750 VPB.n173 VNB 0.02fF
C751 VPB.n174 VNB 0.01fF
C752 VPB.n175 VNB 0.07fF
C753 VPB.n176 VNB 0.16fF
C754 VPB.n177 VNB 0.02fF
C755 VPB.n178 VNB 0.02fF
C756 VPB.n179 VNB 0.02fF
C757 VPB.n180 VNB 0.06fF
C758 VPB.n181 VNB 0.14fF
C759 VPB.n182 VNB 0.20fF
C760 VPB.n183 VNB 0.02fF
C761 VPB.n184 VNB 0.01fF
C762 VPB.n185 VNB 0.02fF
C763 VPB.n186 VNB 0.28fF
C764 VPB.n187 VNB 0.01fF
C765 VPB.n188 VNB 0.02fF
C766 VPB.n189 VNB 0.04fF
C767 VPB.n190 VNB 0.02fF
C768 VPB.n191 VNB 0.02fF
C769 VPB.n192 VNB 0.02fF
C770 VPB.n193 VNB 0.04fF
C771 VPB.n194 VNB 0.02fF
C772 VPB.n195 VNB 0.17fF
C773 VPB.n196 VNB 0.04fF
C774 VPB.n198 VNB 0.02fF
C775 VPB.n199 VNB 0.02fF
C776 VPB.n200 VNB 0.02fF
C777 VPB.n201 VNB 0.02fF
C778 VPB.n203 VNB 0.02fF
C779 VPB.n204 VNB 0.02fF
C780 VPB.n205 VNB 0.02fF
C781 VPB.n207 VNB 0.28fF
C782 VPB.n209 VNB 0.03fF
C783 VPB.n210 VNB 0.02fF
C784 VPB.n211 VNB 0.03fF
C785 VPB.n212 VNB 0.03fF
C786 VPB.n213 VNB 0.28fF
C787 VPB.n214 VNB 0.01fF
C788 VPB.n215 VNB 0.02fF
C789 VPB.n216 VNB 0.04fF
C790 VPB.n217 VNB 0.28fF
C791 VPB.n218 VNB 0.02fF
C792 VPB.n219 VNB 0.02fF
C793 VPB.n220 VNB 0.02fF
C794 VPB.n221 VNB 0.28fF
C795 VPB.n222 VNB 0.02fF
C796 VPB.n223 VNB 0.02fF
C797 VPB.n224 VNB 0.02fF
C798 VPB.n225 VNB 0.28fF
C799 VPB.n226 VNB 0.02fF
C800 VPB.n227 VNB 0.02fF
C801 VPB.n228 VNB 0.02fF
C802 VPB.n229 VNB 0.28fF
C803 VPB.n230 VNB 0.02fF
C804 VPB.n231 VNB 0.02fF
C805 VPB.n232 VNB 0.02fF
C806 VPB.n233 VNB 0.28fF
C807 VPB.n234 VNB 0.02fF
C808 VPB.n235 VNB 0.02fF
C809 VPB.n236 VNB 0.02fF
C810 VPB.n237 VNB 0.28fF
C811 VPB.n238 VNB 0.02fF
C812 VPB.n239 VNB 0.02fF
C813 VPB.n240 VNB 0.02fF
C814 VPB.n241 VNB 0.28fF
C815 VPB.n242 VNB 0.01fF
C816 VPB.n243 VNB 0.02fF
C817 VPB.n244 VNB 0.04fF
C818 VPB.n245 VNB 0.02fF
C819 VPB.n246 VNB 0.02fF
C820 VPB.n247 VNB 0.02fF
C821 VPB.n248 VNB 0.04fF
C822 VPB.n249 VNB 0.02fF
C823 VPB.n250 VNB 0.20fF
C824 VPB.n251 VNB 0.04fF
C825 VPB.n253 VNB 0.02fF
C826 VPB.n254 VNB 0.02fF
C827 VPB.n255 VNB 0.02fF
C828 VPB.n256 VNB 0.02fF
C829 VPB.n258 VNB 0.02fF
C830 VPB.n259 VNB 0.02fF
C831 VPB.n260 VNB 0.02fF
C832 VPB.n262 VNB 0.28fF
C833 VPB.n264 VNB 0.03fF
C834 VPB.n265 VNB 0.02fF
C835 VPB.n266 VNB 0.03fF
C836 VPB.n267 VNB 0.03fF
C837 VPB.n268 VNB 0.28fF
C838 VPB.n269 VNB 0.01fF
C839 VPB.n270 VNB 0.02fF
C840 VPB.n271 VNB 0.04fF
C841 VPB.n272 VNB 0.28fF
C842 VPB.n273 VNB 0.02fF
C843 VPB.n274 VNB 0.02fF
C844 VPB.n275 VNB 0.02fF
C845 VPB.n276 VNB 0.28fF
C846 VPB.n277 VNB 0.02fF
C847 VPB.n278 VNB 0.02fF
C848 VPB.n279 VNB 0.02fF
C849 VPB.n280 VNB 0.28fF
C850 VPB.n281 VNB 0.02fF
C851 VPB.n282 VNB 0.02fF
C852 VPB.n283 VNB 0.02fF
C853 VPB.n284 VNB 0.28fF
C854 VPB.n285 VNB 0.02fF
C855 VPB.n286 VNB 0.02fF
C856 VPB.n287 VNB 0.02fF
C857 VPB.n288 VNB 0.28fF
C858 VPB.n289 VNB 0.02fF
C859 VPB.n290 VNB 0.02fF
C860 VPB.n291 VNB 0.02fF
C861 VPB.n292 VNB 0.28fF
C862 VPB.n293 VNB 0.02fF
C863 VPB.n294 VNB 0.02fF
C864 VPB.n295 VNB 0.02fF
C865 VPB.n296 VNB 0.28fF
C866 VPB.n297 VNB 0.01fF
C867 VPB.n298 VNB 0.02fF
C868 VPB.n299 VNB 0.04fF
C869 VPB.n300 VNB 0.02fF
C870 VPB.n301 VNB 0.02fF
C871 VPB.n302 VNB 0.02fF
C872 VPB.n303 VNB 0.04fF
C873 VPB.n304 VNB 0.02fF
C874 VPB.n305 VNB 0.20fF
C875 VPB.n306 VNB 0.04fF
C876 VPB.n308 VNB 0.02fF
C877 VPB.n309 VNB 0.02fF
C878 VPB.n310 VNB 0.02fF
C879 VPB.n311 VNB 0.02fF
C880 VPB.n313 VNB 0.02fF
C881 VPB.n314 VNB 0.02fF
C882 VPB.n315 VNB 0.02fF
C883 VPB.n317 VNB 0.28fF
C884 VPB.n319 VNB 0.03fF
C885 VPB.n320 VNB 0.02fF
C886 VPB.n321 VNB 0.03fF
C887 VPB.n322 VNB 0.03fF
C888 VPB.n323 VNB 0.28fF
C889 VPB.n324 VNB 0.01fF
C890 VPB.n325 VNB 0.02fF
C891 VPB.n326 VNB 0.04fF
C892 VPB.n327 VNB 0.06fF
C893 VPB.n328 VNB 0.23fF
C894 VPB.n329 VNB 0.02fF
C895 VPB.n330 VNB 0.01fF
C896 VPB.n331 VNB 0.02fF
C897 VPB.n332 VNB 0.14fF
C898 VPB.n333 VNB 0.16fF
C899 VPB.n334 VNB 0.02fF
C900 VPB.n335 VNB 0.02fF
C901 VPB.n336 VNB 0.02fF
C902 VPB.n337 VNB 0.10fF
C903 VPB.n338 VNB 0.02fF
C904 VPB.n339 VNB 0.14fF
C905 VPB.n340 VNB 0.15fF
C906 VPB.n341 VNB 0.02fF
C907 VPB.n342 VNB 0.02fF
C908 VPB.n343 VNB 0.02fF
C909 VPB.n344 VNB 0.14fF
C910 VPB.n345 VNB 0.15fF
C911 VPB.n346 VNB 0.02fF
C912 VPB.n347 VNB 0.02fF
C913 VPB.n348 VNB 0.02fF
C914 VPB.n349 VNB 0.14fF
C915 VPB.n350 VNB 0.16fF
C916 VPB.n351 VNB 0.02fF
C917 VPB.n352 VNB 0.02fF
C918 VPB.n353 VNB 0.02fF
C919 VPB.n354 VNB 0.06fF
C920 VPB.n355 VNB 0.24fF
C921 VPB.n356 VNB 0.02fF
C922 VPB.n357 VNB 0.01fF
C923 VPB.n358 VNB 0.02fF
C924 VPB.n359 VNB 0.28fF
C925 VPB.n360 VNB 0.01fF
C926 VPB.n361 VNB 0.02fF
C927 VPB.n362 VNB 0.04fF
C928 VPB.n363 VNB 0.02fF
C929 VPB.n364 VNB 0.02fF
C930 VPB.n365 VNB 0.02fF
C931 VPB.n366 VNB 0.04fF
C932 VPB.n367 VNB 0.02fF
C933 VPB.n368 VNB 0.20fF
C934 VPB.n369 VNB 0.04fF
C935 VPB.n371 VNB 0.02fF
C936 VPB.n372 VNB 0.02fF
C937 VPB.n373 VNB 0.02fF
C938 VPB.n374 VNB 0.02fF
C939 VPB.n376 VNB 0.02fF
C940 VPB.n377 VNB 0.02fF
C941 VPB.n378 VNB 0.02fF
C942 VPB.n380 VNB 0.28fF
C943 VPB.n382 VNB 0.03fF
C944 VPB.n383 VNB 0.02fF
C945 VPB.n384 VNB 0.03fF
C946 VPB.n385 VNB 0.03fF
C947 VPB.n386 VNB 0.28fF
C948 VPB.n387 VNB 0.01fF
C949 VPB.n388 VNB 0.02fF
C950 VPB.n389 VNB 0.04fF
C951 VPB.n390 VNB 0.05fF
C952 VPB.n391 VNB 0.23fF
C953 VPB.n392 VNB 0.02fF
C954 VPB.n393 VNB 0.01fF
C955 VPB.n394 VNB 0.02fF
C956 VPB.n395 VNB 0.14fF
C957 VPB.n396 VNB 0.16fF
C958 VPB.n397 VNB 0.02fF
C959 VPB.n398 VNB 0.02fF
C960 VPB.n399 VNB 0.02fF
C961 VPB.n400 VNB 0.10fF
C962 VPB.n401 VNB 0.02fF
C963 VPB.n402 VNB 0.14fF
C964 VPB.n403 VNB 0.15fF
C965 VPB.n404 VNB 0.02fF
C966 VPB.n405 VNB 0.02fF
C967 VPB.n406 VNB 0.02fF
C968 VPB.n407 VNB 0.14fF
C969 VPB.n408 VNB 0.15fF
C970 VPB.n409 VNB 0.02fF
C971 VPB.n410 VNB 0.02fF
C972 VPB.n411 VNB 0.02fF
C973 VPB.n412 VNB 0.14fF
C974 VPB.n413 VNB 0.16fF
C975 VPB.n414 VNB 0.02fF
C976 VPB.n415 VNB 0.02fF
C977 VPB.n416 VNB 0.02fF
C978 VPB.n417 VNB 0.06fF
C979 VPB.n418 VNB 0.24fF
C980 VPB.n419 VNB 0.02fF
C981 VPB.n420 VNB 0.01fF
C982 VPB.n421 VNB 0.02fF
C983 VPB.n422 VNB 0.28fF
C984 VPB.n423 VNB 0.01fF
C985 VPB.n424 VNB 0.02fF
C986 VPB.n425 VNB 0.04fF
C987 VPB.n426 VNB 0.02fF
C988 VPB.n427 VNB 0.02fF
C989 VPB.n428 VNB 0.02fF
C990 VPB.n429 VNB 0.04fF
C991 VPB.n430 VNB 0.02fF
C992 VPB.n431 VNB 0.24fF
C993 VPB.n432 VNB 0.04fF
C994 VPB.n434 VNB 0.02fF
C995 VPB.n435 VNB 0.02fF
C996 VPB.n436 VNB 0.02fF
C997 VPB.n437 VNB 0.02fF
C998 VPB.n439 VNB 0.02fF
C999 VPB.n440 VNB 0.02fF
C1000 VPB.n441 VNB 0.02fF
C1001 VPB.n443 VNB 0.28fF
C1002 VPB.n445 VNB 0.03fF
C1003 VPB.n446 VNB 0.02fF
C1004 VPB.n447 VNB 0.03fF
C1005 VPB.n448 VNB 0.03fF
C1006 VPB.n449 VNB 0.28fF
C1007 VPB.n450 VNB 0.01fF
C1008 VPB.n451 VNB 0.02fF
C1009 VPB.n452 VNB 0.04fF
C1010 VPB.n453 VNB 0.28fF
C1011 VPB.n454 VNB 0.02fF
C1012 VPB.n455 VNB 0.02fF
C1013 VPB.n456 VNB 0.02fF
C1014 VPB.n457 VNB 0.05fF
C1015 VPB.n458 VNB 0.21fF
C1016 VPB.n459 VNB 0.02fF
C1017 VPB.n460 VNB 0.01fF
C1018 VPB.n461 VNB 0.02fF
C1019 VPB.n462 VNB 0.14fF
C1020 VPB.n463 VNB 0.16fF
C1021 VPB.n464 VNB 0.02fF
C1022 VPB.n465 VNB 0.02fF
C1023 VPB.n466 VNB 0.02fF
C1024 VPB.n467 VNB 0.10fF
C1025 VPB.n468 VNB 0.02fF
C1026 VPB.n469 VNB 0.14fF
C1027 VPB.n470 VNB 0.16fF
C1028 VPB.n471 VNB 0.02fF
C1029 VPB.n472 VNB 0.02fF
C1030 VPB.n473 VNB 0.02fF
C1031 VPB.n474 VNB 0.14fF
C1032 VPB.n475 VNB 0.15fF
C1033 VPB.n476 VNB 0.02fF
C1034 VPB.n477 VNB 0.02fF
C1035 VPB.n478 VNB 0.02fF
C1036 VPB.n479 VNB 0.14fF
C1037 VPB.n480 VNB 0.15fF
C1038 VPB.n481 VNB 0.02fF
C1039 VPB.n482 VNB 0.02fF
C1040 VPB.n483 VNB 0.02fF
C1041 VPB.n484 VNB 0.10fF
C1042 VPB.n485 VNB 0.02fF
C1043 VPB.n486 VNB 0.14fF
C1044 VPB.n487 VNB 0.16fF
C1045 VPB.n488 VNB 0.02fF
C1046 VPB.n489 VNB 0.02fF
C1047 VPB.n490 VNB 0.02fF
C1048 VPB.n491 VNB 0.14fF
C1049 VPB.n492 VNB 0.16fF
C1050 VPB.n493 VNB 0.02fF
C1051 VPB.n494 VNB 0.02fF
C1052 VPB.n495 VNB 0.02fF
C1053 VPB.n496 VNB 0.06fF
C1054 VPB.n497 VNB 0.21fF
C1055 VPB.n498 VNB 0.02fF
C1056 VPB.n499 VNB 0.01fF
C1057 VPB.n500 VNB 0.02fF
C1058 VPB.n501 VNB 0.28fF
C1059 VPB.n502 VNB 0.02fF
C1060 VPB.n503 VNB 0.02fF
C1061 VPB.n504 VNB 0.02fF
C1062 VPB.n505 VNB 0.28fF
C1063 VPB.n506 VNB 0.01fF
C1064 VPB.n507 VNB 0.02fF
C1065 VPB.n508 VNB 0.04fF
C1066 VPB.n509 VNB 0.02fF
C1067 VPB.n510 VNB 0.02fF
C1068 VPB.n511 VNB 0.02fF
C1069 VPB.n512 VNB 0.04fF
C1070 VPB.n513 VNB 0.02fF
C1071 VPB.n514 VNB 0.29fF
C1072 VPB.n515 VNB 0.04fF
C1073 VPB.n517 VNB 0.02fF
C1074 VPB.n518 VNB 0.02fF
C1075 VPB.n519 VNB 0.02fF
C1076 VPB.n520 VNB 0.02fF
C1077 VPB.n522 VNB 0.02fF
C1078 VPB.n523 VNB 0.02fF
C1079 VPB.n524 VNB 0.02fF
C1080 VPB.n526 VNB 0.28fF
C1081 VPB.n528 VNB 0.03fF
C1082 VPB.n529 VNB 0.02fF
C1083 VPB.n530 VNB 0.03fF
C1084 VPB.n531 VNB 0.03fF
C1085 VPB.n532 VNB 0.28fF
C1086 VPB.n533 VNB 0.01fF
C1087 VPB.n534 VNB 0.02fF
C1088 VPB.n535 VNB 0.04fF
C1089 VPB.n536 VNB 0.28fF
C1090 VPB.n537 VNB 0.02fF
C1091 VPB.n538 VNB 0.02fF
C1092 VPB.n539 VNB 0.02fF
C1093 VPB.n540 VNB 0.05fF
C1094 VPB.n541 VNB 0.21fF
C1095 VPB.n542 VNB 0.02fF
C1096 VPB.n543 VNB 0.01fF
C1097 VPB.n544 VNB 0.02fF
C1098 VPB.n545 VNB 0.14fF
C1099 VPB.n546 VNB 0.16fF
C1100 VPB.n547 VNB 0.02fF
C1101 VPB.n548 VNB 0.02fF
C1102 VPB.n549 VNB 0.02fF
C1103 VPB.n550 VNB 0.10fF
C1104 VPB.n551 VNB 0.02fF
C1105 VPB.n552 VNB 0.14fF
C1106 VPB.n553 VNB 0.16fF
C1107 VPB.n554 VNB 0.02fF
C1108 VPB.n555 VNB 0.02fF
C1109 VPB.n556 VNB 0.02fF
C1110 VPB.n557 VNB 0.14fF
C1111 VPB.n558 VNB 0.15fF
C1112 VPB.n559 VNB 0.02fF
C1113 VPB.n560 VNB 0.02fF
C1114 VPB.n561 VNB 0.02fF
C1115 VPB.n562 VNB 0.14fF
C1116 VPB.n563 VNB 0.15fF
C1117 VPB.n564 VNB 0.02fF
C1118 VPB.n565 VNB 0.02fF
C1119 VPB.n566 VNB 0.02fF
C1120 VPB.n567 VNB 0.10fF
C1121 VPB.n568 VNB 0.02fF
C1122 VPB.n569 VNB 0.14fF
C1123 VPB.n570 VNB 0.16fF
C1124 VPB.n571 VNB 0.02fF
C1125 VPB.n572 VNB 0.02fF
C1126 VPB.n573 VNB 0.02fF
C1127 VPB.n574 VNB 0.14fF
C1128 VPB.n575 VNB 0.16fF
C1129 VPB.n576 VNB 0.02fF
C1130 VPB.n577 VNB 0.02fF
C1131 VPB.n578 VNB 0.02fF
C1132 VPB.n579 VNB 0.06fF
C1133 VPB.n580 VNB 0.21fF
C1134 VPB.n581 VNB 0.02fF
C1135 VPB.n582 VNB 0.01fF
C1136 VPB.n583 VNB 0.02fF
C1137 VPB.n584 VNB 0.28fF
C1138 VPB.n585 VNB 0.02fF
C1139 VPB.n586 VNB 0.02fF
C1140 VPB.n587 VNB 0.02fF
C1141 VPB.n588 VNB 0.28fF
C1142 VPB.n589 VNB 0.01fF
C1143 VPB.n590 VNB 0.02fF
C1144 VPB.n591 VNB 0.04fF
C1145 VPB.n592 VNB 0.02fF
C1146 VPB.n593 VNB 0.02fF
C1147 VPB.n594 VNB 0.02fF
C1148 VPB.n595 VNB 0.04fF
C1149 VPB.n596 VNB 0.02fF
C1150 VPB.n597 VNB 0.24fF
C1151 VPB.n598 VNB 0.04fF
C1152 VPB.n600 VNB 0.02fF
C1153 VPB.n601 VNB 0.02fF
C1154 VPB.n602 VNB 0.02fF
C1155 VPB.n603 VNB 0.02fF
C1156 VPB.n605 VNB 0.02fF
C1157 VPB.n606 VNB 0.02fF
C1158 VPB.n607 VNB 0.02fF
C1159 VPB.n609 VNB 0.28fF
C1160 VPB.n611 VNB 0.03fF
C1161 VPB.n612 VNB 0.02fF
C1162 VPB.n613 VNB 0.03fF
C1163 VPB.n614 VNB 0.03fF
C1164 VPB.n615 VNB 0.28fF
C1165 VPB.n616 VNB 0.01fF
C1166 VPB.n617 VNB 0.02fF
C1167 VPB.n618 VNB 0.04fF
C1168 VPB.n619 VNB 0.05fF
C1169 VPB.n620 VNB 0.23fF
C1170 VPB.n621 VNB 0.02fF
C1171 VPB.n622 VNB 0.01fF
C1172 VPB.n623 VNB 0.02fF
C1173 VPB.n624 VNB 0.14fF
C1174 VPB.n625 VNB 0.16fF
C1175 VPB.n626 VNB 0.02fF
C1176 VPB.n627 VNB 0.02fF
C1177 VPB.n628 VNB 0.02fF
C1178 VPB.n629 VNB 0.10fF
C1179 VPB.n630 VNB 0.02fF
C1180 VPB.n631 VNB 0.14fF
C1181 VPB.n632 VNB 0.15fF
C1182 VPB.n633 VNB 0.02fF
C1183 VPB.n634 VNB 0.02fF
C1184 VPB.n635 VNB 0.02fF
C1185 VPB.n636 VNB 0.14fF
C1186 VPB.n637 VNB 0.15fF
C1187 VPB.n638 VNB 0.02fF
C1188 VPB.n639 VNB 0.02fF
C1189 VPB.n640 VNB 0.02fF
C1190 VPB.n641 VNB 0.14fF
C1191 VPB.n642 VNB 0.16fF
C1192 VPB.n643 VNB 0.02fF
C1193 VPB.n644 VNB 0.02fF
C1194 VPB.n645 VNB 0.02fF
C1195 VPB.n646 VNB 0.06fF
C1196 VPB.n647 VNB 0.24fF
C1197 VPB.n648 VNB 0.02fF
C1198 VPB.n649 VNB 0.01fF
C1199 VPB.n650 VNB 0.02fF
C1200 VPB.n651 VNB 0.28fF
C1201 VPB.n652 VNB 0.01fF
C1202 VPB.n653 VNB 0.02fF
C1203 VPB.n654 VNB 0.04fF
C1204 VPB.n655 VNB 0.02fF
C1205 VPB.n656 VNB 0.02fF
C1206 VPB.n657 VNB 0.02fF
C1207 VPB.n658 VNB 0.04fF
C1208 VPB.n659 VNB 0.02fF
C1209 VPB.n660 VNB 0.24fF
C1210 VPB.n661 VNB 0.04fF
C1211 VPB.n663 VNB 0.02fF
C1212 VPB.n664 VNB 0.02fF
C1213 VPB.n665 VNB 0.02fF
C1214 VPB.n666 VNB 0.02fF
C1215 VPB.n668 VNB 0.02fF
C1216 VPB.n669 VNB 0.02fF
C1217 VPB.n670 VNB 0.02fF
C1218 VPB.n672 VNB 0.28fF
C1219 VPB.n674 VNB 0.03fF
C1220 VPB.n675 VNB 0.02fF
C1221 VPB.n676 VNB 0.03fF
C1222 VPB.n677 VNB 0.03fF
C1223 VPB.n678 VNB 0.28fF
C1224 VPB.n679 VNB 0.01fF
C1225 VPB.n680 VNB 0.02fF
C1226 VPB.n681 VNB 0.04fF
C1227 VPB.n682 VNB 0.28fF
C1228 VPB.n683 VNB 0.02fF
C1229 VPB.n684 VNB 0.02fF
C1230 VPB.n685 VNB 0.02fF
C1231 VPB.n686 VNB 0.05fF
C1232 VPB.n687 VNB 0.21fF
C1233 VPB.n688 VNB 0.02fF
C1234 VPB.n689 VNB 0.01fF
C1235 VPB.n690 VNB 0.02fF
C1236 VPB.n691 VNB 0.14fF
C1237 VPB.n692 VNB 0.16fF
C1238 VPB.n693 VNB 0.02fF
C1239 VPB.n694 VNB 0.02fF
C1240 VPB.n695 VNB 0.02fF
C1241 VPB.n696 VNB 0.10fF
C1242 VPB.n697 VNB 0.02fF
C1243 VPB.n698 VNB 0.14fF
C1244 VPB.n699 VNB 0.16fF
C1245 VPB.n700 VNB 0.02fF
C1246 VPB.n701 VNB 0.02fF
C1247 VPB.n702 VNB 0.02fF
C1248 VPB.n703 VNB 0.14fF
C1249 VPB.n704 VNB 0.15fF
C1250 VPB.n705 VNB 0.02fF
C1251 VPB.n706 VNB 0.02fF
C1252 VPB.n707 VNB 0.02fF
C1253 VPB.n708 VNB 0.14fF
C1254 VPB.n709 VNB 0.15fF
C1255 VPB.n710 VNB 0.02fF
C1256 VPB.n711 VNB 0.02fF
C1257 VPB.n712 VNB 0.02fF
C1258 VPB.n713 VNB 0.10fF
C1259 VPB.n714 VNB 0.02fF
C1260 VPB.n715 VNB 0.14fF
C1261 VPB.n716 VNB 0.16fF
C1262 VPB.n717 VNB 0.02fF
C1263 VPB.n718 VNB 0.02fF
C1264 VPB.n719 VNB 0.02fF
C1265 VPB.n720 VNB 0.14fF
C1266 VPB.n721 VNB 0.16fF
C1267 VPB.n722 VNB 0.02fF
C1268 VPB.n723 VNB 0.02fF
C1269 VPB.n724 VNB 0.02fF
C1270 VPB.n725 VNB 0.06fF
C1271 VPB.n726 VNB 0.21fF
C1272 VPB.n727 VNB 0.02fF
C1273 VPB.n728 VNB 0.01fF
C1274 VPB.n729 VNB 0.02fF
C1275 VPB.n730 VNB 0.28fF
C1276 VPB.n731 VNB 0.02fF
C1277 VPB.n732 VNB 0.02fF
C1278 VPB.n733 VNB 0.02fF
C1279 VPB.n734 VNB 0.28fF
C1280 VPB.n735 VNB 0.01fF
C1281 VPB.n736 VNB 0.02fF
C1282 VPB.n737 VNB 0.04fF
C1283 VPB.n738 VNB 0.02fF
C1284 VPB.n739 VNB 0.02fF
C1285 VPB.n740 VNB 0.02fF
C1286 VPB.n741 VNB 0.04fF
C1287 VPB.n742 VNB 0.02fF
C1288 VPB.n743 VNB 0.29fF
C1289 VPB.n744 VNB 0.04fF
C1290 VPB.n746 VNB 0.02fF
C1291 VPB.n747 VNB 0.02fF
C1292 VPB.n748 VNB 0.02fF
C1293 VPB.n749 VNB 0.02fF
C1294 VPB.n751 VNB 0.02fF
C1295 VPB.n752 VNB 0.02fF
C1296 VPB.n753 VNB 0.02fF
C1297 VPB.n755 VNB 0.28fF
C1298 VPB.n757 VNB 0.03fF
C1299 VPB.n758 VNB 0.02fF
C1300 VPB.n759 VNB 0.03fF
C1301 VPB.n760 VNB 0.03fF
C1302 VPB.n761 VNB 0.28fF
C1303 VPB.n762 VNB 0.01fF
C1304 VPB.n763 VNB 0.02fF
C1305 VPB.n764 VNB 0.04fF
C1306 VPB.n765 VNB 0.28fF
C1307 VPB.n766 VNB 0.02fF
C1308 VPB.n767 VNB 0.02fF
C1309 VPB.n768 VNB 0.02fF
C1310 VPB.n769 VNB 0.05fF
C1311 VPB.n770 VNB 0.21fF
C1312 VPB.n771 VNB 0.02fF
C1313 VPB.n772 VNB 0.01fF
C1314 VPB.n773 VNB 0.02fF
C1315 VPB.n774 VNB 0.14fF
C1316 VPB.n775 VNB 0.16fF
C1317 VPB.n776 VNB 0.02fF
C1318 VPB.n777 VNB 0.02fF
C1319 VPB.n778 VNB 0.02fF
C1320 VPB.n779 VNB 0.10fF
C1321 VPB.n780 VNB 0.02fF
C1322 VPB.n781 VNB 0.14fF
C1323 VPB.n782 VNB 0.16fF
C1324 VPB.n783 VNB 0.02fF
C1325 VPB.n784 VNB 0.02fF
C1326 VPB.n785 VNB 0.02fF
C1327 VPB.n786 VNB 0.14fF
C1328 VPB.n787 VNB 0.15fF
C1329 VPB.n788 VNB 0.02fF
C1330 VPB.n789 VNB 0.02fF
C1331 VPB.n790 VNB 0.02fF
C1332 VPB.n791 VNB 0.14fF
C1333 VPB.n792 VNB 0.15fF
C1334 VPB.n793 VNB 0.02fF
C1335 VPB.n794 VNB 0.02fF
C1336 VPB.n795 VNB 0.02fF
C1337 VPB.n796 VNB 0.10fF
C1338 VPB.n797 VNB 0.02fF
C1339 VPB.n798 VNB 0.14fF
C1340 VPB.n799 VNB 0.16fF
C1341 VPB.n800 VNB 0.02fF
C1342 VPB.n801 VNB 0.02fF
C1343 VPB.n802 VNB 0.02fF
C1344 VPB.n803 VNB 0.14fF
C1345 VPB.n804 VNB 0.16fF
C1346 VPB.n805 VNB 0.02fF
C1347 VPB.n806 VNB 0.02fF
C1348 VPB.n807 VNB 0.02fF
C1349 VPB.n808 VNB 0.06fF
C1350 VPB.n809 VNB 0.21fF
C1351 VPB.n810 VNB 0.02fF
C1352 VPB.n811 VNB 0.01fF
C1353 VPB.n812 VNB 0.02fF
C1354 VPB.n813 VNB 0.28fF
C1355 VPB.n814 VNB 0.02fF
C1356 VPB.n815 VNB 0.02fF
C1357 VPB.n816 VNB 0.02fF
C1358 VPB.n817 VNB 0.28fF
C1359 VPB.n818 VNB 0.01fF
C1360 VPB.n819 VNB 0.02fF
C1361 VPB.n820 VNB 0.04fF
C1362 VPB.n821 VNB 0.02fF
C1363 VPB.n822 VNB 0.02fF
C1364 VPB.n823 VNB 0.02fF
C1365 VPB.n824 VNB 0.04fF
C1366 VPB.n825 VNB 0.02fF
C1367 VPB.n826 VNB 0.24fF
C1368 VPB.n827 VNB 0.04fF
C1369 VPB.n829 VNB 0.02fF
C1370 VPB.n830 VNB 0.02fF
C1371 VPB.n831 VNB 0.02fF
C1372 VPB.n832 VNB 0.02fF
C1373 VPB.n834 VNB 0.02fF
C1374 VPB.n835 VNB 0.02fF
C1375 VPB.n836 VNB 0.02fF
C1376 VPB.n838 VNB 0.28fF
C1377 VPB.n840 VNB 0.03fF
C1378 VPB.n841 VNB 0.02fF
C1379 VPB.n842 VNB 0.03fF
C1380 VPB.n843 VNB 0.03fF
C1381 VPB.n844 VNB 0.28fF
C1382 VPB.n845 VNB 0.01fF
C1383 VPB.n846 VNB 0.02fF
C1384 VPB.n847 VNB 0.04fF
C1385 VPB.n848 VNB 0.05fF
C1386 VPB.n849 VNB 0.23fF
C1387 VPB.n850 VNB 0.02fF
C1388 VPB.n851 VNB 0.01fF
C1389 VPB.n852 VNB 0.02fF
C1390 VPB.n853 VNB 0.14fF
C1391 VPB.n854 VNB 0.16fF
C1392 VPB.n855 VNB 0.02fF
C1393 VPB.n856 VNB 0.02fF
C1394 VPB.n857 VNB 0.02fF
C1395 VPB.n858 VNB 0.10fF
C1396 VPB.n859 VNB 0.02fF
C1397 VPB.n860 VNB 0.14fF
C1398 VPB.n861 VNB 0.15fF
C1399 VPB.n862 VNB 0.02fF
C1400 VPB.n863 VNB 0.02fF
C1401 VPB.n864 VNB 0.02fF
C1402 VPB.n865 VNB 0.14fF
C1403 VPB.n866 VNB 0.15fF
C1404 VPB.n867 VNB 0.02fF
C1405 VPB.n868 VNB 0.02fF
C1406 VPB.n869 VNB 0.02fF
C1407 VPB.n870 VNB 0.14fF
C1408 VPB.n871 VNB 0.16fF
C1409 VPB.n872 VNB 0.02fF
C1410 VPB.n873 VNB 0.02fF
C1411 VPB.n874 VNB 0.02fF
C1412 VPB.n875 VNB 0.02fF
C1413 VPB.n876 VNB 0.04fF
C1414 VPB.n877 VNB 0.04fF
C1415 VPB.n878 VNB 0.02fF
C1416 VPB.n879 VNB 0.02fF
C1417 VPB.n880 VNB 0.02fF
C1418 VPB.n881 VNB 0.02fF
C1419 VPB.n882 VNB 0.02fF
C1420 VPB.n883 VNB 0.02fF
C1421 VPB.n884 VNB 0.02fF
C1422 VPB.n885 VNB 0.02fF
C1423 VPB.n886 VNB 0.14fF
C1424 VPB.n887 VNB 0.16fF
C1425 VPB.n888 VNB 0.02fF
C1426 VPB.n889 VNB 0.02fF
C1427 VPB.n890 VNB 0.06fF
C1428 VPB.n891 VNB 0.21fF
C1429 VPB.n892 VNB 0.02fF
C1430 VPB.n893 VNB 0.01fF
C1431 VPB.n894 VNB 0.02fF
C1432 VPB.n895 VNB 0.28fF
C1433 VPB.n896 VNB 0.02fF
C1434 VPB.n897 VNB 0.02fF
C1435 VPB.n898 VNB 0.02fF
C1436 VPB.n899 VNB 0.28fF
C1437 VPB.n900 VNB 0.01fF
C1438 VPB.n901 VNB 0.02fF
C1439 VPB.n902 VNB 0.04fF
C1440 VPB.n903 VNB 0.02fF
C1441 VPB.n904 VNB 0.02fF
C1442 VPB.n905 VNB 0.02fF
C1443 VPB.n906 VNB 0.04fF
C1444 VPB.n907 VNB 0.02fF
C1445 VPB.n908 VNB 0.29fF
C1446 VPB.n909 VNB 0.04fF
C1447 VPB.n911 VNB 0.02fF
C1448 VPB.n912 VNB 0.02fF
C1449 VPB.n913 VNB 0.02fF
C1450 VPB.n914 VNB 0.02fF
C1451 VPB.n916 VNB 0.02fF
C1452 VPB.n917 VNB 0.02fF
C1453 VPB.n918 VNB 0.02fF
C1454 VPB.n920 VNB 0.28fF
C1455 VPB.n922 VNB 0.03fF
C1456 VPB.n923 VNB 0.02fF
C1457 VPB.n924 VNB 0.03fF
C1458 VPB.n925 VNB 0.03fF
C1459 VPB.n926 VNB 0.28fF
C1460 VPB.n927 VNB 0.01fF
C1461 VPB.n928 VNB 0.02fF
C1462 VPB.n929 VNB 0.04fF
C1463 VPB.n930 VNB 0.28fF
C1464 VPB.n931 VNB 0.02fF
C1465 VPB.n932 VNB 0.02fF
C1466 VPB.n933 VNB 0.02fF
C1467 VPB.n934 VNB 0.05fF
C1468 VPB.n935 VNB 0.21fF
C1469 VPB.n936 VNB 0.02fF
C1470 VPB.n937 VNB 0.01fF
C1471 VPB.n938 VNB 0.02fF
C1472 VPB.n939 VNB 0.14fF
C1473 VPB.n940 VNB 0.16fF
C1474 VPB.n941 VNB 0.02fF
C1475 VPB.n942 VNB 0.02fF
C1476 VPB.n943 VNB 0.02fF
C1477 VPB.n944 VNB 0.10fF
C1478 VPB.n945 VNB 0.02fF
C1479 VPB.n946 VNB 0.14fF
C1480 VPB.n947 VNB 0.16fF
C1481 VPB.n948 VNB 0.02fF
C1482 VPB.n949 VNB 0.02fF
C1483 VPB.n950 VNB 0.02fF
C1484 VPB.n951 VNB 0.14fF
C1485 VPB.n952 VNB 0.15fF
C1486 VPB.n953 VNB 0.02fF
C1487 VPB.n954 VNB 0.02fF
C1488 VPB.n955 VNB 0.02fF
C1489 VPB.n956 VNB 0.14fF
C1490 VPB.n957 VNB 0.15fF
C1491 VPB.n958 VNB 0.02fF
C1492 VPB.n959 VNB 0.02fF
C1493 VPB.n960 VNB 0.02fF
C1494 VPB.n961 VNB 0.10fF
C1495 VPB.n962 VNB 0.02fF
C1496 VPB.n963 VNB 0.14fF
C1497 VPB.n964 VNB 0.16fF
C1498 VPB.n965 VNB 0.02fF
C1499 VPB.n966 VNB 0.02fF
C1500 VPB.n967 VNB 0.02fF
C1501 VPB.n968 VNB 0.14fF
C1502 VPB.n969 VNB 0.16fF
C1503 VPB.n970 VNB 0.02fF
C1504 VPB.n971 VNB 0.02fF
C1505 VPB.n972 VNB 0.02fF
C1506 VPB.n973 VNB 0.06fF
C1507 VPB.n974 VNB 0.21fF
C1508 VPB.n975 VNB 0.02fF
C1509 VPB.n976 VNB 0.01fF
C1510 VPB.n977 VNB 0.02fF
C1511 VPB.n978 VNB 0.28fF
C1512 VPB.n979 VNB 0.02fF
C1513 VPB.n980 VNB 0.02fF
C1514 VPB.n981 VNB 0.02fF
C1515 VPB.n982 VNB 0.28fF
C1516 VPB.n983 VNB 0.01fF
C1517 VPB.n984 VNB 0.02fF
C1518 VPB.n985 VNB 0.04fF
C1519 VPB.n986 VNB 0.02fF
C1520 VPB.n987 VNB 0.02fF
C1521 VPB.n988 VNB 0.02fF
C1522 VPB.n989 VNB 0.04fF
C1523 VPB.n990 VNB 0.02fF
C1524 VPB.n991 VNB 0.24fF
C1525 VPB.n992 VNB 0.04fF
C1526 VPB.n994 VNB 0.02fF
C1527 VPB.n995 VNB 0.02fF
C1528 VPB.n996 VNB 0.02fF
C1529 VPB.n997 VNB 0.02fF
C1530 VPB.n999 VNB 0.02fF
C1531 VPB.n1000 VNB 0.02fF
C1532 VPB.n1001 VNB 0.02fF
C1533 VPB.n1003 VNB 0.28fF
C1534 VPB.n1005 VNB 0.03fF
C1535 VPB.n1006 VNB 0.02fF
C1536 VPB.n1007 VNB 0.03fF
C1537 VPB.n1008 VNB 0.03fF
C1538 VPB.n1009 VNB 0.28fF
C1539 VPB.n1010 VNB 0.01fF
C1540 VPB.n1011 VNB 0.02fF
C1541 VPB.n1012 VNB 0.04fF
C1542 VPB.n1013 VNB 0.05fF
C1543 VPB.n1014 VNB 0.23fF
C1544 VPB.n1015 VNB 0.02fF
C1545 VPB.n1016 VNB 0.01fF
C1546 VPB.n1017 VNB 0.02fF
C1547 VPB.n1018 VNB 0.14fF
C1548 VPB.n1019 VNB 0.16fF
C1549 VPB.n1020 VNB 0.02fF
C1550 VPB.n1021 VNB 0.02fF
C1551 VPB.n1022 VNB 0.02fF
C1552 VPB.n1023 VNB 0.10fF
C1553 VPB.n1024 VNB 0.02fF
C1554 VPB.n1025 VNB 0.14fF
C1555 VPB.n1026 VNB 0.15fF
C1556 VPB.n1027 VNB 0.02fF
C1557 VPB.n1028 VNB 0.02fF
C1558 VPB.n1029 VNB 0.02fF
C1559 VPB.n1030 VNB 0.14fF
C1560 VPB.n1031 VNB 0.15fF
C1561 VPB.n1032 VNB 0.02fF
C1562 VPB.n1033 VNB 0.02fF
C1563 VPB.n1034 VNB 0.02fF
C1564 VPB.n1035 VNB 0.14fF
C1565 VPB.n1036 VNB 0.16fF
C1566 VPB.n1037 VNB 0.02fF
C1567 VPB.n1038 VNB 0.02fF
C1568 VPB.n1039 VNB 0.02fF
C1569 VPB.n1040 VNB 0.06fF
C1570 VPB.n1041 VNB 0.24fF
C1571 VPB.n1042 VNB 0.02fF
C1572 VPB.n1043 VNB 0.01fF
C1573 VPB.n1044 VNB 0.02fF
C1574 VPB.n1045 VNB 0.28fF
C1575 VPB.n1046 VNB 0.01fF
C1576 VPB.n1047 VNB 0.02fF
C1577 VPB.n1048 VNB 0.04fF
C1578 VPB.n1049 VNB 0.02fF
C1579 VPB.n1050 VNB 0.02fF
C1580 VPB.n1051 VNB 0.02fF
C1581 VPB.n1052 VNB 0.04fF
C1582 VPB.n1053 VNB 0.02fF
C1583 VPB.n1054 VNB 0.24fF
C1584 VPB.n1055 VNB 0.04fF
C1585 VPB.n1057 VNB 0.02fF
C1586 VPB.n1058 VNB 0.02fF
C1587 VPB.n1059 VNB 0.02fF
C1588 VPB.n1060 VNB 0.02fF
C1589 VPB.n1062 VNB 0.02fF
C1590 VPB.n1063 VNB 0.02fF
C1591 VPB.n1064 VNB 0.02fF
C1592 VPB.n1066 VNB 0.28fF
C1593 VPB.n1068 VNB 0.03fF
C1594 VPB.n1069 VNB 0.02fF
C1595 VPB.n1070 VNB 0.03fF
C1596 VPB.n1071 VNB 0.03fF
C1597 VPB.n1072 VNB 0.28fF
C1598 VPB.n1073 VNB 0.01fF
C1599 VPB.n1074 VNB 0.02fF
C1600 VPB.n1075 VNB 0.04fF
C1601 VPB.n1076 VNB 0.28fF
C1602 VPB.n1077 VNB 0.02fF
C1603 VPB.n1078 VNB 0.02fF
C1604 VPB.n1079 VNB 0.02fF
C1605 VPB.n1080 VNB 0.05fF
C1606 VPB.n1081 VNB 0.21fF
C1607 VPB.n1082 VNB 0.02fF
C1608 VPB.n1083 VNB 0.01fF
C1609 VPB.n1084 VNB 0.02fF
C1610 VPB.n1085 VNB 0.14fF
C1611 VPB.n1086 VNB 0.16fF
C1612 VPB.n1087 VNB 0.02fF
C1613 VPB.n1088 VNB 0.02fF
C1614 VPB.n1089 VNB 0.02fF
C1615 VPB.n1090 VNB 0.10fF
C1616 VPB.n1091 VNB 0.02fF
C1617 VPB.n1092 VNB 0.14fF
C1618 VPB.n1093 VNB 0.16fF
C1619 VPB.n1094 VNB 0.02fF
C1620 VPB.n1095 VNB 0.02fF
C1621 VPB.n1096 VNB 0.02fF
C1622 VPB.n1097 VNB 0.14fF
C1623 VPB.n1098 VNB 0.15fF
C1624 VPB.n1099 VNB 0.02fF
C1625 VPB.n1100 VNB 0.02fF
C1626 VPB.n1101 VNB 0.02fF
C1627 VPB.n1102 VNB 0.14fF
C1628 VPB.n1103 VNB 0.15fF
C1629 VPB.n1104 VNB 0.02fF
C1630 VPB.n1105 VNB 0.02fF
C1631 VPB.n1106 VNB 0.02fF
C1632 VPB.n1107 VNB 0.10fF
C1633 VPB.n1108 VNB 0.02fF
C1634 VPB.n1109 VNB 0.14fF
C1635 VPB.n1110 VNB 0.16fF
C1636 VPB.n1111 VNB 0.02fF
C1637 VPB.n1112 VNB 0.02fF
C1638 VPB.n1113 VNB 0.02fF
C1639 VPB.n1114 VNB 0.14fF
C1640 VPB.n1115 VNB 0.16fF
C1641 VPB.n1116 VNB 0.02fF
C1642 VPB.n1117 VNB 0.02fF
C1643 VPB.n1118 VNB 0.02fF
C1644 VPB.n1119 VNB 0.06fF
C1645 VPB.n1120 VNB 0.21fF
C1646 VPB.n1121 VNB 0.02fF
C1647 VPB.n1122 VNB 0.01fF
C1648 VPB.n1123 VNB 0.02fF
C1649 VPB.n1124 VNB 0.28fF
C1650 VPB.n1125 VNB 0.02fF
C1651 VPB.n1126 VNB 0.02fF
C1652 VPB.n1127 VNB 0.02fF
C1653 VPB.n1128 VNB 0.28fF
C1654 VPB.n1129 VNB 0.01fF
C1655 VPB.n1130 VNB 0.02fF
C1656 VPB.n1131 VNB 0.04fF
C1657 VPB.n1132 VNB 0.02fF
C1658 VPB.n1133 VNB 0.02fF
C1659 VPB.n1134 VNB 0.02fF
C1660 VPB.n1135 VNB 0.04fF
C1661 VPB.n1136 VNB 0.02fF
C1662 VPB.n1137 VNB 0.29fF
C1663 VPB.n1138 VNB 0.04fF
C1664 VPB.n1140 VNB 0.02fF
C1665 VPB.n1141 VNB 0.02fF
C1666 VPB.n1142 VNB 0.02fF
C1667 VPB.n1143 VNB 0.02fF
C1668 VPB.n1145 VNB 0.02fF
C1669 VPB.n1146 VNB 0.02fF
C1670 VPB.n1147 VNB 0.02fF
C1671 VPB.n1149 VNB 0.28fF
C1672 VPB.n1151 VNB 0.03fF
C1673 VPB.n1152 VNB 0.02fF
C1674 VPB.n1153 VNB 0.03fF
C1675 VPB.n1154 VNB 0.03fF
C1676 VPB.n1155 VNB 0.28fF
C1677 VPB.n1156 VNB 0.01fF
C1678 VPB.n1157 VNB 0.02fF
C1679 VPB.n1158 VNB 0.04fF
C1680 VPB.n1159 VNB 0.28fF
C1681 VPB.n1160 VNB 0.02fF
C1682 VPB.n1161 VNB 0.02fF
C1683 VPB.n1162 VNB 0.02fF
C1684 VPB.n1163 VNB 0.05fF
C1685 VPB.n1164 VNB 0.21fF
C1686 VPB.n1165 VNB 0.02fF
C1687 VPB.n1166 VNB 0.01fF
C1688 VPB.n1167 VNB 0.02fF
C1689 VPB.n1168 VNB 0.14fF
C1690 VPB.n1169 VNB 0.16fF
C1691 VPB.n1170 VNB 0.02fF
C1692 VPB.n1171 VNB 0.02fF
C1693 VPB.n1172 VNB 0.02fF
C1694 VPB.n1173 VNB 0.10fF
C1695 VPB.n1174 VNB 0.02fF
C1696 VPB.n1175 VNB 0.14fF
C1697 VPB.n1176 VNB 0.16fF
C1698 VPB.n1177 VNB 0.02fF
C1699 VPB.n1178 VNB 0.02fF
C1700 VPB.n1179 VNB 0.02fF
C1701 VPB.n1180 VNB 0.14fF
C1702 VPB.n1181 VNB 0.15fF
C1703 VPB.n1182 VNB 0.02fF
C1704 VPB.n1183 VNB 0.02fF
C1705 VPB.n1184 VNB 0.02fF
C1706 VPB.n1185 VNB 0.14fF
C1707 VPB.n1186 VNB 0.15fF
C1708 VPB.n1187 VNB 0.02fF
C1709 VPB.n1188 VNB 0.02fF
C1710 VPB.n1189 VNB 0.02fF
C1711 VPB.n1190 VNB 0.10fF
C1712 VPB.n1191 VNB 0.02fF
C1713 VPB.n1192 VNB 0.14fF
C1714 VPB.n1193 VNB 0.16fF
C1715 VPB.n1194 VNB 0.02fF
C1716 VPB.n1195 VNB 0.02fF
C1717 VPB.n1196 VNB 0.02fF
C1718 VPB.n1197 VNB 0.14fF
C1719 VPB.n1198 VNB 0.16fF
C1720 VPB.n1199 VNB 0.02fF
C1721 VPB.n1200 VNB 0.02fF
C1722 VPB.n1201 VNB 0.02fF
C1723 VPB.n1202 VNB 0.06fF
C1724 VPB.n1203 VNB 0.21fF
C1725 VPB.n1204 VNB 0.02fF
C1726 VPB.n1205 VNB 0.01fF
C1727 VPB.n1206 VNB 0.02fF
C1728 VPB.n1207 VNB 0.28fF
C1729 VPB.n1208 VNB 0.02fF
C1730 VPB.n1209 VNB 0.02fF
C1731 VPB.n1210 VNB 0.02fF
C1732 VPB.n1211 VNB 0.28fF
C1733 VPB.n1212 VNB 0.01fF
C1734 VPB.n1213 VNB 0.02fF
C1735 VPB.n1214 VNB 0.04fF
C1736 VPB.n1215 VNB 0.02fF
C1737 VPB.n1216 VNB 0.02fF
C1738 VPB.n1217 VNB 0.02fF
C1739 VPB.n1218 VNB 0.04fF
C1740 VPB.n1219 VNB 0.02fF
C1741 VPB.n1220 VNB 0.24fF
C1742 VPB.n1221 VNB 0.04fF
C1743 VPB.n1223 VNB 0.02fF
C1744 VPB.n1224 VNB 0.02fF
C1745 VPB.n1225 VNB 0.02fF
C1746 VPB.n1226 VNB 0.02fF
C1747 VPB.n1228 VNB 0.02fF
C1748 VPB.n1229 VNB 0.02fF
C1749 VPB.n1230 VNB 0.02fF
C1750 VPB.n1232 VNB 0.28fF
C1751 VPB.n1234 VNB 0.03fF
C1752 VPB.n1235 VNB 0.02fF
C1753 VPB.n1236 VNB 0.03fF
C1754 VPB.n1237 VNB 0.03fF
C1755 VPB.n1238 VNB 0.28fF
C1756 VPB.n1239 VNB 0.01fF
C1757 VPB.n1240 VNB 0.02fF
C1758 VPB.n1241 VNB 0.04fF
C1759 VPB.n1242 VNB 0.05fF
C1760 VPB.n1243 VNB 0.23fF
C1761 VPB.n1244 VNB 0.02fF
C1762 VPB.n1245 VNB 0.01fF
C1763 VPB.n1246 VNB 0.02fF
C1764 VPB.n1247 VNB 0.14fF
C1765 VPB.n1248 VNB 0.16fF
C1766 VPB.n1249 VNB 0.02fF
C1767 VPB.n1250 VNB 0.02fF
C1768 VPB.n1251 VNB 0.02fF
C1769 VPB.n1252 VNB 0.10fF
C1770 VPB.n1253 VNB 0.02fF
C1771 VPB.n1254 VNB 0.14fF
C1772 VPB.n1255 VNB 0.15fF
C1773 VPB.n1256 VNB 0.02fF
C1774 VPB.n1257 VNB 0.02fF
C1775 VPB.n1258 VNB 0.02fF
C1776 VPB.n1259 VNB 0.14fF
C1777 VPB.n1260 VNB 0.15fF
C1778 VPB.n1261 VNB 0.02fF
C1779 VPB.n1262 VNB 0.02fF
C1780 VPB.n1263 VNB 0.02fF
C1781 VPB.n1264 VNB 0.14fF
C1782 VPB.n1265 VNB 0.16fF
C1783 VPB.n1266 VNB 0.02fF
C1784 VPB.n1267 VNB 0.02fF
C1785 VPB.n1268 VNB 0.02fF
C1786 VPB.n1269 VNB 0.06fF
C1787 VPB.n1270 VNB 0.24fF
C1788 VPB.n1271 VNB 0.02fF
C1789 VPB.n1272 VNB 0.01fF
C1790 VPB.n1273 VNB 0.02fF
C1791 VPB.n1274 VNB 0.28fF
C1792 VPB.n1275 VNB 0.01fF
C1793 VPB.n1276 VNB 0.02fF
C1794 VPB.n1277 VNB 0.04fF
C1795 VPB.n1278 VNB 0.02fF
C1796 VPB.n1279 VNB 0.02fF
C1797 VPB.n1280 VNB 0.02fF
C1798 VPB.n1281 VNB 0.04fF
C1799 VPB.n1282 VNB 0.02fF
C1800 VPB.n1283 VNB 0.24fF
C1801 VPB.n1284 VNB 0.04fF
C1802 VPB.n1286 VNB 0.02fF
C1803 VPB.n1287 VNB 0.02fF
C1804 VPB.n1288 VNB 0.02fF
C1805 VPB.n1289 VNB 0.02fF
C1806 VPB.n1291 VNB 0.02fF
C1807 VPB.n1292 VNB 0.02fF
C1808 VPB.n1293 VNB 0.02fF
C1809 VPB.n1295 VNB 0.28fF
C1810 VPB.n1297 VNB 0.03fF
C1811 VPB.n1298 VNB 0.02fF
C1812 VPB.n1299 VNB 0.03fF
C1813 VPB.n1300 VNB 0.03fF
C1814 VPB.n1301 VNB 0.28fF
C1815 VPB.n1302 VNB 0.01fF
C1816 VPB.n1303 VNB 0.02fF
C1817 VPB.n1304 VNB 0.04fF
C1818 VPB.n1305 VNB 0.28fF
C1819 VPB.n1306 VNB 0.02fF
C1820 VPB.n1307 VNB 0.02fF
C1821 VPB.n1308 VNB 0.02fF
C1822 VPB.n1309 VNB 0.05fF
C1823 VPB.n1310 VNB 0.21fF
C1824 VPB.n1311 VNB 0.02fF
C1825 VPB.n1312 VNB 0.01fF
C1826 VPB.n1313 VNB 0.02fF
C1827 VPB.n1314 VNB 0.14fF
C1828 VPB.n1315 VNB 0.16fF
C1829 VPB.n1316 VNB 0.02fF
C1830 VPB.n1317 VNB 0.02fF
C1831 VPB.n1318 VNB 0.02fF
C1832 VPB.n1319 VNB 0.10fF
C1833 VPB.n1320 VNB 0.02fF
C1834 VPB.n1321 VNB 0.14fF
C1835 VPB.n1322 VNB 0.16fF
C1836 VPB.n1323 VNB 0.02fF
C1837 VPB.n1324 VNB 0.02fF
C1838 VPB.n1325 VNB 0.02fF
C1839 VPB.n1326 VNB 0.14fF
C1840 VPB.n1327 VNB 0.15fF
C1841 VPB.n1328 VNB 0.02fF
C1842 VPB.n1329 VNB 0.02fF
C1843 VPB.n1330 VNB 0.02fF
C1844 VPB.n1331 VNB 0.14fF
C1845 VPB.n1332 VNB 0.15fF
C1846 VPB.n1333 VNB 0.02fF
C1847 VPB.n1334 VNB 0.02fF
C1848 VPB.n1335 VNB 0.02fF
C1849 VPB.n1336 VNB 0.10fF
C1850 VPB.n1337 VNB 0.02fF
C1851 VPB.n1338 VNB 0.14fF
C1852 VPB.n1339 VNB 0.16fF
C1853 VPB.n1340 VNB 0.02fF
C1854 VPB.n1341 VNB 0.02fF
C1855 VPB.n1342 VNB 0.02fF
C1856 VPB.n1343 VNB 0.14fF
C1857 VPB.n1344 VNB 0.16fF
C1858 VPB.n1345 VNB 0.02fF
C1859 VPB.n1346 VNB 0.02fF
C1860 VPB.n1347 VNB 0.02fF
C1861 VPB.n1348 VNB 0.06fF
C1862 VPB.n1349 VNB 0.21fF
C1863 VPB.n1350 VNB 0.02fF
C1864 VPB.n1351 VNB 0.01fF
C1865 VPB.n1352 VNB 0.02fF
C1866 VPB.n1353 VNB 0.28fF
C1867 VPB.n1354 VNB 0.02fF
C1868 VPB.n1355 VNB 0.02fF
C1869 VPB.n1356 VNB 0.02fF
C1870 VPB.n1357 VNB 0.28fF
C1871 VPB.n1358 VNB 0.01fF
C1872 VPB.n1359 VNB 0.02fF
C1873 VPB.n1360 VNB 0.04fF
C1874 VPB.n1361 VNB 0.02fF
C1875 VPB.n1362 VNB 0.02fF
C1876 VPB.n1363 VNB 0.02fF
C1877 VPB.n1364 VNB 0.04fF
C1878 VPB.n1365 VNB 0.02fF
C1879 VPB.n1366 VNB 0.29fF
C1880 VPB.n1367 VNB 0.04fF
C1881 VPB.n1369 VNB 0.02fF
C1882 VPB.n1370 VNB 0.02fF
C1883 VPB.n1371 VNB 0.02fF
C1884 VPB.n1372 VNB 0.02fF
C1885 VPB.n1374 VNB 0.02fF
C1886 VPB.n1375 VNB 0.02fF
C1887 VPB.n1376 VNB 0.02fF
C1888 VPB.n1378 VNB 0.28fF
C1889 VPB.n1380 VNB 0.03fF
C1890 VPB.n1381 VNB 0.02fF
C1891 VPB.n1382 VNB 0.03fF
C1892 VPB.n1383 VNB 0.03fF
C1893 VPB.n1384 VNB 0.28fF
C1894 VPB.n1385 VNB 0.01fF
C1895 VPB.n1386 VNB 0.02fF
C1896 VPB.n1387 VNB 0.04fF
C1897 VPB.n1388 VNB 0.28fF
C1898 VPB.n1389 VNB 0.02fF
C1899 VPB.n1390 VNB 0.02fF
C1900 VPB.n1391 VNB 0.02fF
C1901 VPB.n1392 VNB 0.05fF
C1902 VPB.n1393 VNB 0.21fF
C1903 VPB.n1394 VNB 0.02fF
C1904 VPB.n1395 VNB 0.01fF
C1905 VPB.n1396 VNB 0.02fF
C1906 VPB.n1397 VNB 0.14fF
C1907 VPB.n1398 VNB 0.16fF
C1908 VPB.n1399 VNB 0.02fF
C1909 VPB.n1400 VNB 0.02fF
C1910 VPB.n1401 VNB 0.02fF
C1911 VPB.n1402 VNB 0.10fF
C1912 VPB.n1403 VNB 0.02fF
C1913 VPB.n1404 VNB 0.14fF
C1914 VPB.n1405 VNB 0.16fF
C1915 VPB.n1406 VNB 0.02fF
C1916 VPB.n1407 VNB 0.02fF
C1917 VPB.n1408 VNB 0.02fF
C1918 VPB.n1409 VNB 0.14fF
C1919 VPB.n1410 VNB 0.15fF
C1920 VPB.n1411 VNB 0.02fF
C1921 VPB.n1412 VNB 0.02fF
C1922 VPB.n1413 VNB 0.02fF
C1923 VPB.n1414 VNB 0.14fF
C1924 VPB.n1415 VNB 0.15fF
C1925 VPB.n1416 VNB 0.02fF
C1926 VPB.n1417 VNB 0.02fF
C1927 VPB.n1418 VNB 0.02fF
C1928 VPB.n1419 VNB 0.10fF
C1929 VPB.n1420 VNB 0.02fF
C1930 VPB.n1421 VNB 0.14fF
C1931 VPB.n1422 VNB 0.16fF
C1932 VPB.n1423 VNB 0.02fF
C1933 VPB.n1424 VNB 0.02fF
C1934 VPB.n1425 VNB 0.02fF
C1935 VPB.n1426 VNB 0.14fF
C1936 VPB.n1427 VNB 0.16fF
C1937 VPB.n1428 VNB 0.02fF
C1938 VPB.n1429 VNB 0.02fF
C1939 VPB.n1430 VNB 0.02fF
C1940 VPB.n1431 VNB 0.06fF
C1941 VPB.n1432 VNB 0.21fF
C1942 VPB.n1433 VNB 0.02fF
C1943 VPB.n1434 VNB 0.01fF
C1944 VPB.n1435 VNB 0.02fF
C1945 VPB.n1436 VNB 0.28fF
C1946 VPB.n1437 VNB 0.02fF
C1947 VPB.n1438 VNB 0.02fF
C1948 VPB.n1439 VNB 0.02fF
C1949 VPB.n1440 VNB 0.28fF
C1950 VPB.n1441 VNB 0.01fF
C1951 VPB.n1442 VNB 0.02fF
C1952 VPB.n1443 VNB 0.04fF
C1953 VPB.n1444 VNB 0.02fF
C1954 VPB.n1445 VNB 0.02fF
C1955 VPB.n1446 VNB 0.02fF
C1956 VPB.n1447 VNB 0.04fF
C1957 VPB.n1448 VNB 0.02fF
C1958 VPB.n1449 VNB 0.24fF
C1959 VPB.n1450 VNB 0.04fF
C1960 VPB.n1452 VNB 0.02fF
C1961 VPB.n1453 VNB 0.02fF
C1962 VPB.n1454 VNB 0.02fF
C1963 VPB.n1455 VNB 0.02fF
C1964 VPB.n1457 VNB 0.02fF
C1965 VPB.n1458 VNB 0.02fF
C1966 VPB.n1459 VNB 0.02fF
C1967 VPB.n1461 VNB 0.28fF
C1968 VPB.n1463 VNB 0.03fF
C1969 VPB.n1464 VNB 0.02fF
C1970 VPB.n1465 VNB 0.03fF
C1971 VPB.n1466 VNB 0.03fF
C1972 VPB.n1467 VNB 0.28fF
C1973 VPB.n1468 VNB 0.01fF
C1974 VPB.n1469 VNB 0.02fF
C1975 VPB.n1470 VNB 0.04fF
C1976 VPB.n1471 VNB 0.05fF
C1977 VPB.n1472 VNB 0.23fF
C1978 VPB.n1473 VNB 0.02fF
C1979 VPB.n1474 VNB 0.01fF
C1980 VPB.n1475 VNB 0.02fF
C1981 VPB.n1476 VNB 0.14fF
C1982 VPB.n1477 VNB 0.16fF
C1983 VPB.n1478 VNB 0.02fF
C1984 VPB.n1479 VNB 0.02fF
C1985 VPB.n1480 VNB 0.02fF
C1986 VPB.n1481 VNB 0.10fF
C1987 VPB.n1482 VNB 0.02fF
C1988 VPB.n1483 VNB 0.14fF
C1989 VPB.n1484 VNB 0.15fF
C1990 VPB.n1485 VNB 0.02fF
C1991 VPB.n1486 VNB 0.02fF
C1992 VPB.n1487 VNB 0.02fF
C1993 VPB.n1488 VNB 0.14fF
C1994 VPB.n1489 VNB 0.15fF
C1995 VPB.n1490 VNB 0.02fF
C1996 VPB.n1491 VNB 0.02fF
C1997 VPB.n1492 VNB 0.02fF
C1998 VPB.n1493 VNB 0.14fF
C1999 VPB.n1494 VNB 0.16fF
C2000 VPB.n1495 VNB 0.02fF
C2001 VPB.n1496 VNB 0.02fF
C2002 VPB.n1497 VNB 0.02fF
C2003 VPB.n1498 VNB 0.06fF
C2004 VPB.n1499 VNB 0.24fF
C2005 VPB.n1500 VNB 0.02fF
C2006 VPB.n1501 VNB 0.01fF
C2007 VPB.n1502 VNB 0.02fF
C2008 VPB.n1503 VNB 0.28fF
C2009 VPB.n1504 VNB 0.01fF
C2010 VPB.n1505 VNB 0.02fF
C2011 VPB.n1506 VNB 0.04fF
C2012 VPB.n1507 VNB 0.02fF
C2013 VPB.n1508 VNB 0.02fF
C2014 VPB.n1509 VNB 0.02fF
C2015 VPB.n1510 VNB 0.04fF
C2016 VPB.n1511 VNB 0.02fF
C2017 VPB.n1512 VNB 0.24fF
C2018 VPB.n1513 VNB 0.04fF
C2019 VPB.n1515 VNB 0.02fF
C2020 VPB.n1516 VNB 0.02fF
C2021 VPB.n1517 VNB 0.02fF
C2022 VPB.n1518 VNB 0.02fF
C2023 VPB.n1520 VNB 0.02fF
C2024 VPB.n1521 VNB 0.02fF
C2025 VPB.n1522 VNB 0.02fF
C2026 VPB.n1524 VNB 0.28fF
C2027 VPB.n1526 VNB 0.03fF
C2028 VPB.n1527 VNB 0.02fF
C2029 VPB.n1528 VNB 0.03fF
C2030 VPB.n1529 VNB 0.03fF
C2031 VPB.n1530 VNB 0.28fF
C2032 VPB.n1531 VNB 0.01fF
C2033 VPB.n1532 VNB 0.02fF
C2034 VPB.n1533 VNB 0.04fF
C2035 VPB.n1534 VNB 0.28fF
C2036 VPB.n1535 VNB 0.02fF
C2037 VPB.n1536 VNB 0.02fF
C2038 VPB.n1537 VNB 0.02fF
C2039 VPB.n1538 VNB 0.05fF
C2040 VPB.n1539 VNB 0.21fF
C2041 VPB.n1540 VNB 0.02fF
C2042 VPB.n1541 VNB 0.01fF
C2043 VPB.n1542 VNB 0.02fF
C2044 VPB.n1543 VNB 0.14fF
C2045 VPB.n1544 VNB 0.16fF
C2046 VPB.n1545 VNB 0.02fF
C2047 VPB.n1546 VNB 0.02fF
C2048 VPB.n1547 VNB 0.02fF
C2049 VPB.n1548 VNB 0.10fF
C2050 VPB.n1549 VNB 0.02fF
C2051 VPB.n1550 VNB 0.14fF
C2052 VPB.n1551 VNB 0.16fF
C2053 VPB.n1552 VNB 0.02fF
C2054 VPB.n1553 VNB 0.02fF
C2055 VPB.n1554 VNB 0.02fF
C2056 VPB.n1555 VNB 0.14fF
C2057 VPB.n1556 VNB 0.15fF
C2058 VPB.n1557 VNB 0.02fF
C2059 VPB.n1558 VNB 0.02fF
C2060 VPB.n1559 VNB 0.02fF
C2061 VPB.n1560 VNB 0.14fF
C2062 VPB.n1561 VNB 0.15fF
C2063 VPB.n1562 VNB 0.02fF
C2064 VPB.n1563 VNB 0.02fF
C2065 VPB.n1564 VNB 0.02fF
C2066 VPB.n1565 VNB 0.10fF
C2067 VPB.n1566 VNB 0.02fF
C2068 VPB.n1567 VNB 0.14fF
C2069 VPB.n1568 VNB 0.16fF
C2070 VPB.n1569 VNB 0.02fF
C2071 VPB.n1570 VNB 0.02fF
C2072 VPB.n1571 VNB 0.02fF
C2073 VPB.n1572 VNB 0.14fF
C2074 VPB.n1573 VNB 0.16fF
C2075 VPB.n1574 VNB 0.02fF
C2076 VPB.n1575 VNB 0.02fF
C2077 VPB.n1576 VNB 0.02fF
C2078 VPB.n1577 VNB 0.06fF
C2079 VPB.n1578 VNB 0.21fF
C2080 VPB.n1579 VNB 0.02fF
C2081 VPB.n1580 VNB 0.01fF
C2082 VPB.n1581 VNB 0.02fF
C2083 VPB.n1582 VNB 0.28fF
C2084 VPB.n1583 VNB 0.02fF
C2085 VPB.n1584 VNB 0.02fF
C2086 VPB.n1585 VNB 0.02fF
C2087 VPB.n1586 VNB 0.28fF
C2088 VPB.n1587 VNB 0.01fF
C2089 VPB.n1588 VNB 0.02fF
C2090 VPB.n1589 VNB 0.04fF
C2091 VPB.n1590 VNB 0.04fF
C2092 VPB.n1591 VNB 0.02fF
C2093 VPB.n1592 VNB 0.02fF
C2094 VPB.n1593 VNB 0.02fF
C2095 VPB.n1594 VNB 0.02fF
C2096 VPB.n1595 VNB 0.02fF
C2097 VPB.n1596 VNB 0.02fF
C2098 VPB.n1597 VNB 0.02fF
C2099 VPB.n1598 VNB 0.02fF
C2100 VPB.n1599 VNB 0.02fF
C2101 VPB.n1600 VNB 0.02fF
C2102 VPB.n1601 VNB 0.03fF
C2103 VPB.n1602 VNB 0.04fF
C2104 VPB.n1603 VNB 0.02fF
C2105 VPB.n1604 VNB 0.02fF
C2106 VPB.n1605 VNB 0.02fF
C2107 VPB.n1606 VNB 0.04fF
C2108 VPB.n1607 VNB 0.04fF
C2109 VPB.n1609 VNB 0.43fF
C2110 a_10507_159.n0 VNB 0.05fF
C2111 a_10507_159.n1 VNB 0.72fF
C2112 a_10507_159.n2 VNB 0.72fF
C2113 a_10507_159.n3 VNB 0.84fF
C2114 a_10507_159.n4 VNB 0.26fF
C2115 a_10507_159.n5 VNB 0.34fF
C2116 a_10507_159.n6 VNB 0.38fF
C2117 a_10507_159.t22 VNB 0.76fF
C2118 a_10507_159.n7 VNB 0.50fF
C2119 a_10507_159.n8 VNB 0.43fF
C2120 a_10507_159.n9 VNB 0.52fF
C2121 a_10507_159.n10 VNB 0.41fF
C2122 a_10507_159.n11 VNB 0.72fF
C2123 a_10507_159.n12 VNB 0.72fF
C2124 a_10507_159.n13 VNB 0.84fF
C2125 a_10507_159.n14 VNB 0.26fF
C2126 a_10507_159.n15 VNB 0.34fF
C2127 a_10507_159.n16 VNB 0.05fF
C2128 a_10507_159.n17 VNB 0.07fF
C2129 a_10507_159.n18 VNB 0.05fF
C2130 a_10507_159.n19 VNB 0.46fF
C2131 a_10507_159.n20 VNB 0.59fF
C2132 a_10507_159.n21 VNB 0.38fF
C2133 a_10507_159.t25 VNB 0.76fF
C2134 a_10507_159.n22 VNB 0.50fF
C2135 a_10507_159.n23 VNB 0.38fF
C2136 a_10507_159.n24 VNB 0.74fF
C2137 a_10507_159.n25 VNB 2.80fF
C2138 a_10507_159.n26 VNB 1.14fF
C2139 a_10507_159.n27 VNB 0.74fF
C2140 a_10507_159.n28 VNB 0.59fF
C2141 a_10507_159.n29 VNB 0.06fF
C2142 a_10507_159.n30 VNB 0.46fF
C2143 a_10507_159.n31 VNB 0.06fF
.ends
