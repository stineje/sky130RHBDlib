magic
tech sky130A
magscale 1 2
timestamp 1647326732
<< nwell >>
rect 52 -435 352 37
<< pmos >>
rect 144 -399 174 1
rect 232 -399 262 1
<< pdiff >>
rect 88 -107 144 1
rect 88 -141 98 -107
rect 132 -141 144 -107
rect 88 -175 144 -141
rect 88 -209 98 -175
rect 132 -209 144 -175
rect 88 -243 144 -209
rect 88 -277 98 -243
rect 132 -277 144 -243
rect 88 -399 144 -277
rect 174 -107 232 1
rect 174 -141 186 -107
rect 220 -141 232 -107
rect 174 -175 232 -141
rect 174 -209 186 -175
rect 220 -209 232 -175
rect 174 -243 232 -209
rect 174 -277 186 -243
rect 220 -277 232 -243
rect 174 -399 232 -277
rect 262 -107 316 1
rect 262 -141 274 -107
rect 308 -141 316 -107
rect 262 -175 316 -141
rect 262 -209 274 -175
rect 308 -209 316 -175
rect 262 -243 316 -209
rect 262 -277 274 -243
rect 308 -277 316 -243
rect 262 -399 316 -277
<< pdiffc >>
rect 98 -141 132 -107
rect 98 -209 132 -175
rect 98 -277 132 -243
rect 186 -141 220 -107
rect 186 -209 220 -175
rect 186 -277 220 -243
rect 274 -141 308 -107
rect 274 -209 308 -175
rect 274 -277 308 -243
<< poly >>
rect 144 1 174 27
rect 232 1 262 27
rect 144 -430 174 -399
rect 232 -430 262 -399
rect 144 -460 262 -430
<< locali >>
rect 98 -107 132 -91
rect 98 -175 132 -141
rect 98 -243 132 -209
rect 98 -293 132 -277
rect 186 -107 220 -91
rect 186 -175 220 -141
rect 186 -243 220 -209
rect 186 -293 220 -277
rect 274 -107 308 -91
rect 274 -175 308 -141
rect 274 -243 308 -209
rect 274 -293 308 -277
<< end >>
