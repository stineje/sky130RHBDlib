magic
tech sky130A
magscale 1 2
timestamp 1652393950
<< nwell >>
rect 87 1529 579 1550
rect 753 1529 1245 1550
rect 1419 1529 1911 1550
rect 84 1508 582 1529
rect 34 1503 582 1508
rect 750 1504 1248 1529
rect 1416 1505 1914 1529
rect 34 1456 580 1503
rect 752 1460 1246 1504
rect 1418 1502 1914 1505
rect 1418 1463 1912 1502
rect 750 1456 1246 1460
rect 34 1446 582 1456
rect 84 786 582 1446
rect 750 786 1248 1456
rect 1416 1455 1912 1463
rect 1416 786 1914 1455
<< pwell >>
rect -34 -34 2032 544
<< pdiffc >>
rect 141 1331 175 1365
rect 229 1331 263 1365
rect 317 1331 351 1365
rect 405 1331 439 1365
rect 493 1331 527 1365
rect 805 1331 839 1365
rect 981 1331 1015 1365
rect 1157 1331 1191 1365
rect 1473 1331 1507 1365
rect 1649 1331 1683 1365
rect 1825 1331 1859 1365
rect 141 1059 175 1093
rect 229 1059 263 1093
rect 493 1059 527 1093
rect 893 1059 927 1093
rect 1561 1059 1595 1093
rect 1737 1059 1771 1093
<< psubdiff >>
rect 34 482 632 544
rect 700 482 1298 544
rect 1366 482 1964 544
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 632 17
rect 34 -34 632 -17
rect 700 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1298 17
rect 700 -34 1298 -17
rect 1366 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1964 17
rect 1366 -34 1964 -17
<< nsubdiff >>
rect 34 1497 632 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 632 1497
rect 700 1497 1298 1514
rect 700 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1298 1497
rect 1366 1497 1964 1514
rect 1366 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1964 1497
rect 1946 1459 1964 1463
rect 34 822 635 884
rect 697 822 1301 884
rect 1363 822 1964 884
<< psubdiffcont >>
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
<< poly >>
rect 175 944 187 974
rect 1145 944 1157 974
rect 1507 944 1519 974
rect 168 375 198 413
rect 362 381 392 383
rect 834 375 864 413
rect 1134 382 1164 413
rect 1500 375 1530 413
rect 1694 382 1724 383
<< locali >>
rect 34 1497 632 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 632 1497
rect 34 1446 632 1463
rect 700 1497 1298 1514
rect 700 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1298 1497
rect 700 1446 1298 1463
rect 1366 1497 1964 1514
rect 1366 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1964 1497
rect 1366 1446 1964 1463
rect 141 1365 175 1446
rect 141 1313 175 1331
rect 229 1365 265 1399
rect 317 1365 351 1446
rect 229 1313 263 1331
rect 317 1313 351 1331
rect 405 1365 439 1399
rect 405 1313 439 1331
rect 493 1365 527 1446
rect 493 1313 527 1331
rect 805 1365 1191 1399
rect 805 1313 839 1331
rect 981 1313 1015 1331
rect 1157 1313 1191 1331
rect 1473 1365 1859 1399
rect 1473 1313 1507 1331
rect 1649 1313 1683 1331
rect 1825 1313 1859 1331
rect 141 1093 175 1111
rect 141 1025 175 1059
rect 229 1093 263 1111
rect 405 1075 439 1111
rect 493 1093 527 1111
rect 805 1075 839 1127
rect 893 1093 927 1111
rect 229 1025 405 1059
rect 493 1025 527 1059
rect 1069 1075 1103 1111
rect 1157 1075 1191 1111
rect 1473 1075 1507 1111
rect 1561 1093 1595 1111
rect 1737 1093 1771 1127
rect 805 1023 839 1054
rect 893 1025 1103 1059
rect 1473 1025 1507 1038
rect 1561 1025 1867 1059
rect 131 433 165 942
rect 353 908 361 942
rect 353 439 387 908
rect 353 433 357 439
rect 871 430 905 908
rect 1167 433 1201 942
rect 1463 423 1497 908
rect 1685 433 1719 974
rect 1833 346 1867 1025
rect 1745 312 1867 346
rect 1745 269 1779 312
rect 219 34 253 159
rect 885 34 919 159
rect 1551 34 1585 159
rect 34 17 632 34
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 632 17
rect 34 -34 632 -17
rect 700 17 1298 34
rect 700 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1298 17
rect 700 -34 1298 -17
rect 1366 17 1964 34
rect 1366 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1964 17
rect 1366 -34 1964 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
<< metal1 >>
rect 34 1497 632 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 632 1497
rect 34 1446 632 1463
rect 700 1497 1298 1514
rect 700 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1298 1497
rect 700 1446 1298 1463
rect 1366 1497 1964 1514
rect 1366 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1964 1497
rect 1366 1446 1964 1463
rect 475 1025 799 1059
rect 1135 1025 1466 1059
rect 166 871 905 905
rect 389 797 1690 831
rect 1201 399 1453 433
rect 449 219 1744 253
rect 34 17 632 34
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 632 17
rect 34 -34 632 -17
rect 700 17 1298 34
rect 700 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1298 17
rect 700 -34 1298 -17
rect 1366 17 1964 34
rect 1366 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1964 17
rect 1366 -34 1964 -17
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 148 0 1 888
box -53 -33 29 33
use pmos2_1  pmos2_1_0
timestamp 1647326732
transform 1 0 43 0 1 1404
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 149 -1 0 942
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_5
timestamp 1648060378
transform 0 1 149 -1 0 417
box -32 -28 34 26
use nmos_bottom  nmos_bottom_0
timestamp 1651256857
transform -1 0 360 0 1 73
box 0 0 248 302
use diff_ring_side  diff_ring_side_1
timestamp 1652319726
transform 1 0 0 0 1 0
box -87 -34 87 1550
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 370 0 1 814
box -53 -33 29 33
use pmos2_1  pmos2_1_1
timestamp 1647326732
transform 1 0 219 0 1 1404
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 379 -1 0 942
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 422 0 1 1042
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 -1 369 1 0 415
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 430 0 1 236
box -53 -33 29 33
use nmos_top  nmos_top_0
timestamp 1651256841
transform -1 0 552 0 1 73
box 0 0 246 308
use pmos2_1  pmos2_1_3
timestamp 1647326732
transform -1 0 1113 0 1 1404
box 52 -460 352 37
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 822 0 -1 1042
box -53 -33 29 33
use nmos_bottom  nmos_bottom_1
timestamp 1651256857
transform -1 0 1026 0 1 73
box 0 0 248 302
use diff_ring_side  diff_ring_side_2
timestamp 1652319726
transform 1 0 666 0 1 0
box -87 -34 87 1550
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 888 0 1 888
box -53 -33 29 33
use pmos2_1  pmos2_1_2
timestamp 1647326732
transform -1 0 1289 0 1 1404
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_7
timestamp 1648060378
transform 0 -1 887 -1 0 942
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 1086 0 -1 1042
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_4
timestamp 1648060378
transform 0 -1 887 -1 0 417
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 1096 0 1 236
box -53 -33 29 33
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1651256895
transform 1 0 972 0 1 73
box 0 0 248 309
use poly_li1_contact  poly_li1_contact_6
timestamp 1648060378
transform 0 -1 1183 -1 0 942
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 1184 0 1 416
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 -1 1183 -1 0 417
box -32 -28 34 26
use diff_ring_side  diff_ring_side_3
timestamp 1652319726
transform 1 0 1332 0 1 0
box -87 -34 87 1550
use poly_li1_contact  poly_li1_contact_10
timestamp 1648060378
transform 0 -1 1479 -1 0 417
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform 1 0 1480 0 1 416
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 1762 0 1 236
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_11
timestamp 1648060378
transform 0 -1 1701 -1 0 417
box -32 -28 34 26
use nmos_bottom  nmos_bottom_2
timestamp 1651256857
transform -1 0 1692 0 1 73
box 0 0 248 302
use nmos_top_trim2  nmos_top_trim2_2
timestamp 1651256905
transform -1 0 1886 0 1 73
box 0 0 248 309
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform 1 0 1702 0 1 814
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_8
timestamp 1648060378
transform 0 1 1481 -1 0 942
box -32 -28 34 26
use pmos2_1  pmos2_1_4
timestamp 1647326732
transform 1 0 1375 0 1 1404
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_9
timestamp 1648060378
transform 0 1 1707 -1 0 942
box -32 -28 34 26
use pmos2_1  pmos2_1_5
timestamp 1647326732
transform 1 0 1551 0 1 1404
box 52 -460 352 37
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform 1 0 1490 0 1 1042
box -53 -33 29 33
use diff_ring_side  diff_ring_side_0
timestamp 1652319726
transform 1 0 1998 0 1 0
box -87 -34 87 1550
<< end >>
