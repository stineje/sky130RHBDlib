* SPICE3 file created from VOTER3X1.ext - technology: sky130A

.subckt VOTER3X1 Y A B C VPB VNB
M1000 a_217_1005.t1 A VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VNB B a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=1.6781p pd=12.81u as=0p ps=0u
M1002 VNB a_1027_944# a_1444_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_217_1005.t6 a_1027_944# a_881_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_392_181.t5 a_1027_944# a_881_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_392_181.t1 A a_881_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t3 B a_217_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_881_1005.t6 a_1027_944# a_217_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t5 a_392_181.t7 a_2183_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPB.t1 A a_217_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_881_1005.t3 B a_217_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_881_1005.t4 a_1027_944# a_392_181.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_2183_182.t0 a_392_181.t9 VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_217_1005.t2 B VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_217_1005.t4 B a_881_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VNB B a_778_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_881_1005.t0 A a_392_181.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB A 0.48fF
C1 B VPB 0.40fF
C2 a_1027_944# VPB 0.18fF
C3 B A 0.93fF
C4 a_1027_944# A 0.30fF
C5 a_1027_944# B 0.15fF
R0 VPB VPB.n143 122.382
R1 VPB.n121 VPB.n119 94.117
R2 VPB.n207 VPB.n205 94.117
R3 VPB.n67 VPB.n65 91.036
R4 VPB.n29 VPB.n23 76.136
R5 VPB.n29 VPB.n28 76
R6 VPB.n33 VPB.n32 76
R7 VPB.n39 VPB.n38 76
R8 VPB.n43 VPB.n42 76
R9 VPB.n69 VPB.n68 76
R10 VPB.n73 VPB.n72 76
R11 VPB.n77 VPB.n76 76
R12 VPB.n81 VPB.n80 76
R13 VPB.n85 VPB.n84 76
R14 VPB.n89 VPB.n88 76
R15 VPB.n93 VPB.n92 76
R16 VPB.n97 VPB.n96 76
R17 VPB.n123 VPB.n122 76
R18 VPB.n233 VPB.n232 76
R19 VPB.n229 VPB.n228 76
R20 VPB.n225 VPB.n224 76
R21 VPB.n221 VPB.n220 76
R22 VPB.n217 VPB.n216 76
R23 VPB.n213 VPB.n212 76
R24 VPB.n209 VPB.n208 76
R25 VPB.n183 VPB.n182 76
R26 VPB.n179 VPB.n178 76
R27 VPB.n174 VPB.n173 76
R28 VPB.n169 VPB.n168 76
R29 VPB.n162 VPB.n161 76
R30 VPB.n157 VPB.n156 76
R31 VPB.n152 VPB.n151 76
R32 VPB.n147 VPB.n146 76
R33 VPB.n35 VPB.n34 68.979
R34 VPB.n26 VPB.n25 64.528
R35 VPB.n188 VPB.n187 61.764
R36 VPB.n102 VPB.n101 61.764
R37 VPB.n48 VPB.n47 61.764
R38 VPB.n148 VPB.t4 55.465
R39 VPB.n175 VPB.t1 55.465
R40 VPB.n37 VPB.t0 55.106
R41 VPB.n24 VPB.t5 55.106
R42 VPB.n171 VPB.n170 48.952
R43 VPB.n154 VPB.n153 44.502
R44 VPB.n164 VPB.n163 41.183
R45 VPB.n146 VPB.n127 20.452
R46 VPB.n23 VPB.n20 20.452
R47 VPB.n166 VPB.n165 17.801
R48 VPB.n163 VPB.t2 14.282
R49 VPB.n163 VPB.t3 14.282
R50 VPB.n23 VPB.n22 13.653
R51 VPB.n22 VPB.n21 13.653
R52 VPB.n28 VPB.n27 13.653
R53 VPB.n27 VPB.n26 13.653
R54 VPB.n32 VPB.n31 13.653
R55 VPB.n31 VPB.n30 13.653
R56 VPB.n38 VPB.n36 13.653
R57 VPB.n36 VPB.n35 13.653
R58 VPB.n42 VPB.n41 13.653
R59 VPB.n41 VPB.n40 13.653
R60 VPB.n68 VPB.n67 13.653
R61 VPB.n67 VPB.n66 13.653
R62 VPB.n72 VPB.n71 13.653
R63 VPB.n71 VPB.n70 13.653
R64 VPB.n76 VPB.n75 13.653
R65 VPB.n75 VPB.n74 13.653
R66 VPB.n80 VPB.n79 13.653
R67 VPB.n79 VPB.n78 13.653
R68 VPB.n84 VPB.n83 13.653
R69 VPB.n83 VPB.n82 13.653
R70 VPB.n88 VPB.n87 13.653
R71 VPB.n87 VPB.n86 13.653
R72 VPB.n92 VPB.n91 13.653
R73 VPB.n91 VPB.n90 13.653
R74 VPB.n96 VPB.n95 13.653
R75 VPB.n95 VPB.n94 13.653
R76 VPB.n122 VPB.n121 13.653
R77 VPB.n121 VPB.n120 13.653
R78 VPB.n232 VPB.n231 13.653
R79 VPB.n231 VPB.n230 13.653
R80 VPB.n228 VPB.n227 13.653
R81 VPB.n227 VPB.n226 13.653
R82 VPB.n224 VPB.n223 13.653
R83 VPB.n223 VPB.n222 13.653
R84 VPB.n220 VPB.n219 13.653
R85 VPB.n219 VPB.n218 13.653
R86 VPB.n216 VPB.n215 13.653
R87 VPB.n215 VPB.n214 13.653
R88 VPB.n212 VPB.n211 13.653
R89 VPB.n211 VPB.n210 13.653
R90 VPB.n208 VPB.n207 13.653
R91 VPB.n207 VPB.n206 13.653
R92 VPB.n182 VPB.n181 13.653
R93 VPB.n181 VPB.n180 13.653
R94 VPB.n178 VPB.n177 13.653
R95 VPB.n177 VPB.n176 13.653
R96 VPB.n173 VPB.n172 13.653
R97 VPB.n172 VPB.n171 13.653
R98 VPB.n168 VPB.n167 13.653
R99 VPB.n167 VPB.n166 13.653
R100 VPB.n161 VPB.n160 13.653
R101 VPB.n160 VPB.n159 13.653
R102 VPB.n156 VPB.n155 13.653
R103 VPB.n155 VPB.n154 13.653
R104 VPB.n151 VPB.n150 13.653
R105 VPB.n150 VPB.n149 13.653
R106 VPB.n146 VPB.n145 13.653
R107 VPB.n145 VPB.n144 13.653
R108 VPB.n159 VPB.n158 13.35
R109 VPB.n63 VPB.n46 13.276
R110 VPB.n46 VPB.n44 13.276
R111 VPB.n117 VPB.n100 13.276
R112 VPB.n100 VPB.n98 13.276
R113 VPB.n203 VPB.n186 13.276
R114 VPB.n186 VPB.n184 13.276
R115 VPB.n127 VPB.n126 13.276
R116 VPB.n126 VPB.n124 13.276
R117 VPB.n20 VPB.n19 13.276
R118 VPB.n19 VPB.n17 13.276
R119 VPB.n68 VPB.n64 13.276
R120 VPB.n122 VPB.n118 13.276
R121 VPB.n208 VPB.n204 13.276
R122 VPB.n4 VPB.n2 12.796
R123 VPB.n4 VPB.n3 12.564
R124 VPB.n13 VPB.n12 12.198
R125 VPB.n11 VPB.n10 12.198
R126 VPB.n8 VPB.n7 12.198
R127 VPB.n126 VPB.n125 7.5
R128 VPB.n132 VPB.n131 7.5
R129 VPB.n135 VPB.n134 7.5
R130 VPB.n137 VPB.n136 7.5
R131 VPB.n140 VPB.n139 7.5
R132 VPB.n128 VPB.n127 7.5
R133 VPB.n186 VPB.n185 7.5
R134 VPB.n198 VPB.n197 7.5
R135 VPB.n192 VPB.n191 7.5
R136 VPB.n194 VPB.n193 7.5
R137 VPB.n200 VPB.n190 7.5
R138 VPB.n200 VPB.n188 7.5
R139 VPB.n203 VPB.n202 7.5
R140 VPB.n100 VPB.n99 7.5
R141 VPB.n112 VPB.n111 7.5
R142 VPB.n106 VPB.n105 7.5
R143 VPB.n108 VPB.n107 7.5
R144 VPB.n114 VPB.n104 7.5
R145 VPB.n114 VPB.n102 7.5
R146 VPB.n117 VPB.n116 7.5
R147 VPB.n46 VPB.n45 7.5
R148 VPB.n58 VPB.n57 7.5
R149 VPB.n52 VPB.n51 7.5
R150 VPB.n54 VPB.n53 7.5
R151 VPB.n60 VPB.n50 7.5
R152 VPB.n60 VPB.n48 7.5
R153 VPB.n63 VPB.n62 7.5
R154 VPB.n20 VPB.n16 7.5
R155 VPB.n2 VPB.n1 7.5
R156 VPB.n7 VPB.n6 7.5
R157 VPB.n10 VPB.n9 7.5
R158 VPB.n19 VPB.n18 7.5
R159 VPB.n14 VPB.n0 7.5
R160 VPB.n64 VPB.n63 7.176
R161 VPB.n118 VPB.n117 7.176
R162 VPB.n204 VPB.n203 7.176
R163 VPB.n199 VPB.n196 6.729
R164 VPB.n195 VPB.n192 6.729
R165 VPB.n113 VPB.n110 6.729
R166 VPB.n109 VPB.n106 6.729
R167 VPB.n59 VPB.n56 6.729
R168 VPB.n55 VPB.n52 6.729
R169 VPB.n195 VPB.n194 6.728
R170 VPB.n199 VPB.n198 6.728
R171 VPB.n202 VPB.n201 6.728
R172 VPB.n109 VPB.n108 6.728
R173 VPB.n113 VPB.n112 6.728
R174 VPB.n116 VPB.n115 6.728
R175 VPB.n55 VPB.n54 6.728
R176 VPB.n59 VPB.n58 6.728
R177 VPB.n62 VPB.n61 6.728
R178 VPB.n129 VPB.n128 6.728
R179 VPB.n133 VPB.n130 6.728
R180 VPB.n138 VPB.n135 6.728
R181 VPB.n142 VPB.n140 6.728
R182 VPB.n142 VPB.n141 6.728
R183 VPB.n138 VPB.n137 6.728
R184 VPB.n133 VPB.n132 6.728
R185 VPB.n168 VPB.n164 6.458
R186 VPB.n16 VPB.n15 6.398
R187 VPB.n190 VPB.n189 6.166
R188 VPB.n104 VPB.n103 6.166
R189 VPB.n50 VPB.n49 6.166
R190 VPB.n144 VPB 4.45
R191 VPB.n28 VPB.n24 2.691
R192 VPB.n38 VPB.n37 2.332
R193 VPB.n151 VPB.n148 1.794
R194 VPB.n178 VPB.n175 1.435
R195 VPB.n14 VPB.n5 1.402
R196 VPB.n14 VPB.n8 1.402
R197 VPB.n14 VPB.n11 1.402
R198 VPB.n14 VPB.n13 1.402
R199 VPB.n15 VPB.n14 0.735
R200 VPB.n14 VPB.n4 0.735
R201 VPB.n200 VPB.n199 0.387
R202 VPB.n200 VPB.n195 0.387
R203 VPB.n201 VPB.n200 0.387
R204 VPB.n114 VPB.n113 0.387
R205 VPB.n114 VPB.n109 0.387
R206 VPB.n115 VPB.n114 0.387
R207 VPB.n60 VPB.n59 0.387
R208 VPB.n60 VPB.n55 0.387
R209 VPB.n61 VPB.n60 0.387
R210 VPB.n143 VPB.n142 0.387
R211 VPB.n143 VPB.n138 0.387
R212 VPB.n143 VPB.n133 0.387
R213 VPB.n143 VPB.n129 0.387
R214 VPB.n69 VPB.n43 0.272
R215 VPB.n123 VPB.n97 0.272
R216 VPB.n209 VPB.n183 0.272
R217 VPB.n147 VPB 0.198
R218 VPB.n33 VPB.n29 0.136
R219 VPB.n39 VPB.n33 0.136
R220 VPB.n43 VPB.n39 0.136
R221 VPB.n73 VPB.n69 0.136
R222 VPB.n77 VPB.n73 0.136
R223 VPB.n81 VPB.n77 0.136
R224 VPB.n85 VPB.n81 0.136
R225 VPB.n89 VPB.n85 0.136
R226 VPB.n93 VPB.n89 0.136
R227 VPB.n97 VPB.n93 0.136
R228 VPB.n233 VPB.n229 0.136
R229 VPB.n229 VPB.n225 0.136
R230 VPB.n225 VPB.n221 0.136
R231 VPB.n221 VPB.n217 0.136
R232 VPB.n217 VPB.n213 0.136
R233 VPB.n213 VPB.n209 0.136
R234 VPB.n183 VPB.n179 0.136
R235 VPB.n179 VPB.n174 0.136
R236 VPB.n174 VPB.n169 0.136
R237 VPB.n169 VPB.n162 0.136
R238 VPB.n162 VPB.n157 0.136
R239 VPB.n157 VPB.n152 0.136
R240 VPB.n152 VPB.n147 0.136
R241 VPB VPB.n123 0.068
R242 VPB VPB.n233 0.068
R243 a_217_1005.n4 a_217_1005.n3 195.987
R244 a_217_1005.n2 a_217_1005.t6 89.553
R245 a_217_1005.n4 a_217_1005.n0 75.271
R246 a_217_1005.n3 a_217_1005.n2 75.214
R247 a_217_1005.n5 a_217_1005.n4 36.517
R248 a_217_1005.n3 a_217_1005.t5 14.338
R249 a_217_1005.n1 a_217_1005.t7 14.282
R250 a_217_1005.n1 a_217_1005.t4 14.282
R251 a_217_1005.n0 a_217_1005.t3 14.282
R252 a_217_1005.n0 a_217_1005.t2 14.282
R253 a_217_1005.n5 a_217_1005.t0 14.282
R254 a_217_1005.t1 a_217_1005.n5 14.282
R255 a_217_1005.n2 a_217_1005.n1 12.119
R256 a_881_1005.n4 a_881_1005.n3 196.002
R257 a_881_1005.n2 a_881_1005.t0 89.553
R258 a_881_1005.n5 a_881_1005.n4 75.27
R259 a_881_1005.n3 a_881_1005.n2 75.214
R260 a_881_1005.n4 a_881_1005.n0 36.52
R261 a_881_1005.n3 a_881_1005.t5 14.338
R262 a_881_1005.n0 a_881_1005.t7 14.282
R263 a_881_1005.n0 a_881_1005.t6 14.282
R264 a_881_1005.n1 a_881_1005.t1 14.282
R265 a_881_1005.n1 a_881_1005.t4 14.282
R266 a_881_1005.n5 a_881_1005.t2 14.282
R267 a_881_1005.t3 a_881_1005.n5 14.282
R268 a_881_1005.n2 a_881_1005.n1 12.119
R269 a_392_181.n4 a_392_181.t7 512.525
R270 a_392_181.n4 a_392_181.t9 371.139
R271 a_392_181.n5 a_392_181.t8 273.368
R272 a_392_181.n16 a_392_181.n6 226.775
R273 a_392_181.n6 a_392_181.n5 153.043
R274 a_392_181.n6 a_392_181.n3 110.158
R275 a_392_181.n5 a_392_181.n4 105.194
R276 a_392_181.n15 a_392_181.n14 98.501
R277 a_392_181.n15 a_392_181.n10 96.417
R278 a_392_181.n16 a_392_181.n15 78.403
R279 a_392_181.n3 a_392_181.n2 75.271
R280 a_392_181.n19 a_392_181.n0 55.263
R281 a_392_181.n10 a_392_181.n9 30
R282 a_392_181.n14 a_392_181.n13 30
R283 a_392_181.n18 a_392_181.n17 30
R284 a_392_181.n19 a_392_181.n18 25.263
R285 a_392_181.n8 a_392_181.n7 24.383
R286 a_392_181.n12 a_392_181.n11 24.383
R287 a_392_181.n10 a_392_181.n8 23.684
R288 a_392_181.n14 a_392_181.n12 23.684
R289 a_392_181.n18 a_392_181.n16 20.417
R290 a_392_181.n1 a_392_181.t0 14.282
R291 a_392_181.n1 a_392_181.t1 14.282
R292 a_392_181.n2 a_392_181.t4 14.282
R293 a_392_181.n2 a_392_181.t5 14.282
R294 a_392_181.n3 a_392_181.n1 12.119
R295 a_1444_73.t0 a_1444_73.n1 93.333
R296 a_1444_73.n4 a_1444_73.n2 55.07
R297 a_1444_73.t0 a_1444_73.n0 8.137
R298 a_1444_73.n4 a_1444_73.n3 4.619
R299 a_1444_73.t0 a_1444_73.n4 0.071
R300 a_112_73.t0 a_112_73.n0 93.333
R301 a_112_73.n2 a_112_73.n1 51.404
R302 a_112_73.t0 a_112_73.n6 7.911
R303 a_112_73.t0 a_112_73.n2 4.039
R304 a_112_73.n5 a_112_73.n3 4.032
R305 a_112_73.n5 a_112_73.n4 3.644
R306 a_112_73.t0 a_112_73.n5 1.099
R307 a_778_73.t0 a_778_73.n0 93.333
R308 a_778_73.n3 a_778_73.n1 55.048
R309 a_778_73.n3 a_778_73.n2 2.097
R310 a_778_73.t0 a_778_73.n3 0.11
R311 a_2183_182.n3 a_2183_182.n1 355.848
R312 a_2183_182.n3 a_2183_182.n2 30
R313 a_2183_182.n4 a_2183_182.n0 24.383
R314 a_2183_182.n4 a_2183_182.n3 23.684
R315 a_2183_182.n1 a_2183_182.t1 14.282
R316 a_2183_182.n1 a_2183_182.t0 14.282
R317 VNB VNB.n218 300.778
R318 VNB.n83 VNB.n82 199.897
R319 VNB.n66 VNB.n65 199.897
R320 VNB.n15 VNB.n14 199.897
R321 VNB.n176 VNB.n174 154.509
R322 VNB.n99 VNB.n97 154.509
R323 VNB.n35 VNB.n33 154.509
R324 VNB.n113 VNB.n72 84.842
R325 VNB.n22 VNB.n21 84.842
R326 VNB.n49 VNB.n4 84.842
R327 VNB.n150 VNB.n141 76.136
R328 VNB.n150 VNB.n149 76
R329 VNB.n205 VNB.n204 76
R330 VNB.n193 VNB.n192 76
R331 VNB.n189 VNB.n188 76
R332 VNB.n185 VNB.n184 76
R333 VNB.n181 VNB.n180 76
R334 VNB.n177 VNB.n173 76
R335 VNB.n163 VNB.n162 76
R336 VNB.n159 VNB.n158 76
R337 VNB.n157 VNB.n156 49.896
R338 VNB.n115 VNB.n114 36.678
R339 VNB.n24 VNB.n23 36.678
R340 VNB.n51 VNB.n50 36.678
R341 VNB.n145 VNB.n144 35.01
R342 VNB.n143 VNB.n142 29.127
R343 VNB.n153 VNB.t2 20.794
R344 VNB.n141 VNB.n138 20.452
R345 VNB.n206 VNB.n205 20.452
R346 VNB.n146 VNB.n145 20.094
R347 VNB.n155 VNB.n154 20.094
R348 VNB.n92 VNB.n91 20.094
R349 VNB.n145 VNB.n143 19.017
R350 VNB.n149 VNB.n148 13.653
R351 VNB.n148 VNB.n147 13.653
R352 VNB.n158 VNB.n157 13.653
R353 VNB.n162 VNB.n161 13.653
R354 VNB.n161 VNB.n160 13.653
R355 VNB.n95 VNB.n94 13.653
R356 VNB.n94 VNB.n93 13.653
R357 VNB.n100 VNB.n99 13.653
R358 VNB.n99 VNB.n98 13.653
R359 VNB.n103 VNB.n102 13.653
R360 VNB.n102 VNB.n101 13.653
R361 VNB.n106 VNB.n105 13.653
R362 VNB.n105 VNB.n104 13.653
R363 VNB.n109 VNB.n108 13.653
R364 VNB.n108 VNB.n107 13.653
R365 VNB.n112 VNB.n111 13.653
R366 VNB.n111 VNB.n110 13.653
R367 VNB.n116 VNB.n115 13.653
R368 VNB.n119 VNB.n118 13.653
R369 VNB.n118 VNB.n117 13.653
R370 VNB.n122 VNB.n121 13.653
R371 VNB.n121 VNB.n120 13.653
R372 VNB.n177 VNB.n176 13.653
R373 VNB.n176 VNB.n175 13.653
R374 VNB.n180 VNB.n179 13.653
R375 VNB.n179 VNB.n178 13.653
R376 VNB.n184 VNB.n183 13.653
R377 VNB.n183 VNB.n182 13.653
R378 VNB.n188 VNB.n187 13.653
R379 VNB.n187 VNB.n186 13.653
R380 VNB.n192 VNB.n191 13.653
R381 VNB.n191 VNB.n190 13.653
R382 VNB.n25 VNB.n24 13.653
R383 VNB.n28 VNB.n27 13.653
R384 VNB.n27 VNB.n26 13.653
R385 VNB.n31 VNB.n30 13.653
R386 VNB.n30 VNB.n29 13.653
R387 VNB.n36 VNB.n35 13.653
R388 VNB.n35 VNB.n34 13.653
R389 VNB.n39 VNB.n38 13.653
R390 VNB.n38 VNB.n37 13.653
R391 VNB.n42 VNB.n41 13.653
R392 VNB.n41 VNB.n40 13.653
R393 VNB.n45 VNB.n44 13.653
R394 VNB.n44 VNB.n43 13.653
R395 VNB.n48 VNB.n47 13.653
R396 VNB.n47 VNB.n46 13.653
R397 VNB.n52 VNB.n51 13.653
R398 VNB.n55 VNB.n54 13.653
R399 VNB.n54 VNB.n53 13.653
R400 VNB.n205 VNB.n0 13.653
R401 VNB VNB.n0 13.653
R402 VNB.n141 VNB.n140 13.653
R403 VNB.n140 VNB.n139 13.653
R404 VNB.n213 VNB.n210 13.577
R405 VNB.n126 VNB.n124 13.276
R406 VNB.n138 VNB.n126 13.276
R407 VNB.n75 VNB.n73 13.276
R408 VNB.n88 VNB.n75 13.276
R409 VNB.n58 VNB.n56 13.276
R410 VNB.n71 VNB.n58 13.276
R411 VNB.n7 VNB.n5 13.276
R412 VNB.n20 VNB.n7 13.276
R413 VNB.n96 VNB.n95 13.276
R414 VNB.n100 VNB.n96 13.276
R415 VNB.n103 VNB.n100 13.276
R416 VNB.n106 VNB.n103 13.276
R417 VNB.n109 VNB.n106 13.276
R418 VNB.n112 VNB.n109 13.276
R419 VNB.n119 VNB.n116 13.276
R420 VNB.n122 VNB.n119 13.276
R421 VNB.n123 VNB.n122 13.276
R422 VNB.n177 VNB.n123 13.276
R423 VNB.n180 VNB.n177 13.276
R424 VNB.n28 VNB.n25 13.276
R425 VNB.n31 VNB.n28 13.276
R426 VNB.n32 VNB.n31 13.276
R427 VNB.n36 VNB.n32 13.276
R428 VNB.n39 VNB.n36 13.276
R429 VNB.n42 VNB.n39 13.276
R430 VNB.n45 VNB.n42 13.276
R431 VNB.n48 VNB.n45 13.276
R432 VNB.n55 VNB.n52 13.276
R433 VNB.n205 VNB.n55 13.276
R434 VNB.n3 VNB.n1 13.276
R435 VNB.n206 VNB.n3 13.276
R436 VNB.n91 VNB.n90 12.837
R437 VNB.n113 VNB.n112 10.764
R438 VNB.n49 VNB.n48 10.764
R439 VNB.n95 VNB.n92 9.329
R440 VNB.n90 VNB.n89 7.566
R441 VNB.n215 VNB.n214 7.5
R442 VNB.n81 VNB.n80 7.5
R443 VNB.n77 VNB.n76 7.5
R444 VNB.n75 VNB.n74 7.5
R445 VNB.n88 VNB.n87 7.5
R446 VNB.n64 VNB.n63 7.5
R447 VNB.n60 VNB.n59 7.5
R448 VNB.n58 VNB.n57 7.5
R449 VNB.n71 VNB.n70 7.5
R450 VNB.n13 VNB.n12 7.5
R451 VNB.n9 VNB.n8 7.5
R452 VNB.n7 VNB.n6 7.5
R453 VNB.n20 VNB.n19 7.5
R454 VNB.n207 VNB.n206 7.5
R455 VNB.n3 VNB.n2 7.5
R456 VNB.n212 VNB.n211 7.5
R457 VNB.n132 VNB.n131 7.5
R458 VNB.n128 VNB.n127 7.5
R459 VNB.n126 VNB.n125 7.5
R460 VNB.n138 VNB.n137 7.5
R461 VNB.n96 VNB.n88 7.176
R462 VNB.n123 VNB.n71 7.176
R463 VNB.n32 VNB.n20 7.176
R464 VNB.n217 VNB.n215 7.011
R465 VNB.n84 VNB.n81 7.011
R466 VNB.n79 VNB.n77 7.011
R467 VNB.n67 VNB.n64 7.011
R468 VNB.n62 VNB.n60 7.011
R469 VNB.n16 VNB.n13 7.011
R470 VNB.n11 VNB.n9 7.011
R471 VNB.n134 VNB.n132 7.011
R472 VNB.n130 VNB.n128 7.011
R473 VNB.n87 VNB.n86 7.01
R474 VNB.n79 VNB.n78 7.01
R475 VNB.n84 VNB.n83 7.01
R476 VNB.n70 VNB.n69 7.01
R477 VNB.n62 VNB.n61 7.01
R478 VNB.n67 VNB.n66 7.01
R479 VNB.n19 VNB.n18 7.01
R480 VNB.n11 VNB.n10 7.01
R481 VNB.n16 VNB.n15 7.01
R482 VNB.n137 VNB.n136 7.01
R483 VNB.n130 VNB.n129 7.01
R484 VNB.n134 VNB.n133 7.01
R485 VNB.n217 VNB.n216 7.01
R486 VNB.n213 VNB.n212 6.788
R487 VNB.n208 VNB.n207 6.788
R488 VNB.n152 VNB.n151 4.551
R489 VNB.n149 VNB.n146 4.305
R490 VNB.n116 VNB.n113 2.511
R491 VNB.n25 VNB.n22 2.511
R492 VNB.n52 VNB.n49 2.511
R493 VNB.t2 VNB.n152 2.238
R494 VNB.n218 VNB.n209 0.921
R495 VNB.n218 VNB.n213 0.476
R496 VNB.n218 VNB.n208 0.475
R497 VNB.n154 VNB.n153 0.358
R498 VNB.n165 VNB.n164 0.272
R499 VNB.n173 VNB.n172 0.272
R500 VNB.n197 VNB.n196 0.272
R501 VNB.n85 VNB.n79 0.246
R502 VNB.n86 VNB.n85 0.246
R503 VNB.n85 VNB.n84 0.246
R504 VNB.n68 VNB.n62 0.246
R505 VNB.n69 VNB.n68 0.246
R506 VNB.n68 VNB.n67 0.246
R507 VNB.n17 VNB.n11 0.246
R508 VNB.n18 VNB.n17 0.246
R509 VNB.n17 VNB.n16 0.246
R510 VNB.n135 VNB.n130 0.246
R511 VNB.n136 VNB.n135 0.246
R512 VNB.n135 VNB.n134 0.246
R513 VNB.n218 VNB.n217 0.246
R514 VNB.n204 VNB 0.198
R515 VNB.n158 VNB.n155 0.179
R516 VNB.n159 VNB.n150 0.136
R517 VNB.n163 VNB.n159 0.136
R518 VNB.n164 VNB.n163 0.136
R519 VNB.n166 VNB.n165 0.136
R520 VNB.n167 VNB.n166 0.136
R521 VNB.n168 VNB.n167 0.136
R522 VNB.n169 VNB.n168 0.136
R523 VNB.n170 VNB.n169 0.136
R524 VNB.n171 VNB.n170 0.136
R525 VNB.n172 VNB.n171 0.136
R526 VNB.n185 VNB.n181 0.136
R527 VNB.n189 VNB.n185 0.136
R528 VNB.n193 VNB.n189 0.136
R529 VNB.n194 VNB.n193 0.136
R530 VNB.n195 VNB.n194 0.136
R531 VNB.n196 VNB.n195 0.136
R532 VNB.n198 VNB.n197 0.136
R533 VNB.n199 VNB.n198 0.136
R534 VNB.n200 VNB.n199 0.136
R535 VNB.n201 VNB.n200 0.136
R536 VNB.n202 VNB.n201 0.136
R537 VNB.n203 VNB.n202 0.136
R538 VNB.n204 VNB.n203 0.136
R539 VNB.n173 VNB 0.068
R540 VNB.n181 VNB 0.068
C6 VPB VNB 10.25fF
C7 a_2183_182.n0 VNB 0.04fF
C8 a_2183_182.n1 VNB 1.02fF
C9 a_2183_182.n2 VNB 0.04fF
C10 a_2183_182.n3 VNB 0.50fF
C11 a_2183_182.n4 VNB 0.06fF
C12 a_778_73.n0 VNB 0.02fF
C13 a_778_73.n1 VNB 0.13fF
C14 a_778_73.n2 VNB 0.12fF
C15 a_778_73.n3 VNB 0.14fF
C16 a_112_73.n0 VNB 0.02fF
C17 a_112_73.n1 VNB 0.10fF
C18 a_112_73.n2 VNB 0.09fF
C19 a_112_73.n3 VNB 0.07fF
C20 a_112_73.n4 VNB 0.02fF
C21 a_112_73.n5 VNB 0.01fF
C22 a_112_73.n6 VNB 0.06fF
C23 a_1444_73.n0 VNB 0.06fF
C24 a_1444_73.n1 VNB 0.03fF
C25 a_1444_73.n2 VNB 0.13fF
C26 a_1444_73.n3 VNB 0.04fF
C27 a_1444_73.n4 VNB 0.18fF
C28 a_392_181.n0 VNB 0.04fF
C29 a_392_181.n1 VNB 0.38fF
C30 a_392_181.n2 VNB 0.46fF
C31 a_392_181.n3 VNB 0.21fF
C32 a_392_181.n4 VNB 0.24fF
C33 a_392_181.t8 VNB 0.48fF
C34 a_392_181.n5 VNB 0.48fF
C35 a_392_181.n6 VNB 0.45fF
C36 a_392_181.n7 VNB 0.03fF
C37 a_392_181.n8 VNB 0.04fF
C38 a_392_181.n9 VNB 0.03fF
C39 a_392_181.n10 VNB 0.08fF
C40 a_392_181.n11 VNB 0.03fF
C41 a_392_181.n12 VNB 0.04fF
C42 a_392_181.n13 VNB 0.03fF
C43 a_392_181.n14 VNB 0.09fF
C44 a_392_181.n15 VNB 0.96fF
C45 a_392_181.n16 VNB 0.26fF
C46 a_392_181.n17 VNB 0.03fF
C47 a_392_181.n18 VNB 0.05fF
C48 a_392_181.n19 VNB 0.04fF
C49 a_881_1005.n0 VNB 0.28fF
C50 a_881_1005.n1 VNB 0.29fF
C51 a_881_1005.n2 VNB 0.20fF
C52 a_881_1005.n3 VNB 0.57fF
C53 a_881_1005.n4 VNB 0.25fF
C54 a_881_1005.n5 VNB 0.36fF
C55 a_217_1005.n0 VNB 0.40fF
C56 a_217_1005.n1 VNB 0.32fF
C57 a_217_1005.n2 VNB 0.23fF
C58 a_217_1005.n3 VNB 0.61fF
C59 a_217_1005.n4 VNB 0.27fF
C60 a_217_1005.n5 VNB 0.36fF
C61 VPB.n0 VNB 0.10fF
C62 VPB.n1 VNB 0.03fF
C63 VPB.n2 VNB 0.02fF
C64 VPB.n3 VNB 0.05fF
C65 VPB.n4 VNB 0.01fF
C66 VPB.n6 VNB 0.02fF
C67 VPB.n7 VNB 0.02fF
C68 VPB.n9 VNB 0.02fF
C69 VPB.n10 VNB 0.02fF
C70 VPB.n12 VNB 0.02fF
C71 VPB.n14 VNB 0.45fF
C72 VPB.n16 VNB 0.04fF
C73 VPB.n17 VNB 0.02fF
C74 VPB.n18 VNB 0.02fF
C75 VPB.n19 VNB 0.02fF
C76 VPB.n20 VNB 0.04fF
C77 VPB.n21 VNB 0.27fF
C78 VPB.n22 VNB 0.03fF
C79 VPB.n23 VNB 0.03fF
C80 VPB.n24 VNB 0.06fF
C81 VPB.n25 VNB 0.13fF
C82 VPB.n26 VNB 0.19fF
C83 VPB.n27 VNB 0.02fF
C84 VPB.n28 VNB 0.01fF
C85 VPB.n29 VNB 0.07fF
C86 VPB.n30 VNB 0.16fF
C87 VPB.n31 VNB 0.02fF
C88 VPB.n32 VNB 0.02fF
C89 VPB.n33 VNB 0.02fF
C90 VPB.n34 VNB 0.13fF
C91 VPB.n35 VNB 0.19fF
C92 VPB.n36 VNB 0.02fF
C93 VPB.n37 VNB 0.06fF
C94 VPB.n38 VNB 0.01fF
C95 VPB.n39 VNB 0.02fF
C96 VPB.n40 VNB 0.27fF
C97 VPB.n41 VNB 0.01fF
C98 VPB.n42 VNB 0.02fF
C99 VPB.n43 VNB 0.04fF
C100 VPB.n44 VNB 0.02fF
C101 VPB.n45 VNB 0.02fF
C102 VPB.n46 VNB 0.02fF
C103 VPB.n47 VNB 0.16fF
C104 VPB.n48 VNB 0.04fF
C105 VPB.n49 VNB 0.03fF
C106 VPB.n50 VNB 0.02fF
C107 VPB.n51 VNB 0.02fF
C108 VPB.n52 VNB 0.02fF
C109 VPB.n53 VNB 0.03fF
C110 VPB.n54 VNB 0.02fF
C111 VPB.n56 VNB 0.02fF
C112 VPB.n57 VNB 0.02fF
C113 VPB.n58 VNB 0.02fF
C114 VPB.n60 VNB 0.27fF
C115 VPB.n62 VNB 0.02fF
C116 VPB.n63 VNB 0.02fF
C117 VPB.n64 VNB 0.03fF
C118 VPB.n65 VNB 0.03fF
C119 VPB.n66 VNB 0.27fF
C120 VPB.n67 VNB 0.01fF
C121 VPB.n68 VNB 0.02fF
C122 VPB.n69 VNB 0.04fF
C123 VPB.n70 VNB 0.27fF
C124 VPB.n71 VNB 0.02fF
C125 VPB.n72 VNB 0.02fF
C126 VPB.n73 VNB 0.02fF
C127 VPB.n74 VNB 0.27fF
C128 VPB.n75 VNB 0.02fF
C129 VPB.n76 VNB 0.02fF
C130 VPB.n77 VNB 0.02fF
C131 VPB.n78 VNB 0.27fF
C132 VPB.n79 VNB 0.02fF
C133 VPB.n80 VNB 0.02fF
C134 VPB.n81 VNB 0.02fF
C135 VPB.n82 VNB 0.27fF
C136 VPB.n83 VNB 0.02fF
C137 VPB.n84 VNB 0.02fF
C138 VPB.n85 VNB 0.02fF
C139 VPB.n86 VNB 0.27fF
C140 VPB.n87 VNB 0.02fF
C141 VPB.n88 VNB 0.02fF
C142 VPB.n89 VNB 0.02fF
C143 VPB.n90 VNB 0.27fF
C144 VPB.n91 VNB 0.02fF
C145 VPB.n92 VNB 0.02fF
C146 VPB.n93 VNB 0.02fF
C147 VPB.n94 VNB 0.27fF
C148 VPB.n95 VNB 0.01fF
C149 VPB.n96 VNB 0.02fF
C150 VPB.n97 VNB 0.04fF
C151 VPB.n98 VNB 0.02fF
C152 VPB.n99 VNB 0.02fF
C153 VPB.n100 VNB 0.02fF
C154 VPB.n101 VNB 0.19fF
C155 VPB.n102 VNB 0.04fF
C156 VPB.n103 VNB 0.03fF
C157 VPB.n104 VNB 0.02fF
C158 VPB.n105 VNB 0.02fF
C159 VPB.n106 VNB 0.02fF
C160 VPB.n107 VNB 0.03fF
C161 VPB.n108 VNB 0.02fF
C162 VPB.n110 VNB 0.02fF
C163 VPB.n111 VNB 0.02fF
C164 VPB.n112 VNB 0.02fF
C165 VPB.n114 VNB 0.27fF
C166 VPB.n116 VNB 0.03fF
C167 VPB.n117 VNB 0.02fF
C168 VPB.n118 VNB 0.03fF
C169 VPB.n119 VNB 0.03fF
C170 VPB.n120 VNB 0.27fF
C171 VPB.n121 VNB 0.01fF
C172 VPB.n122 VNB 0.02fF
C173 VPB.n123 VNB 0.03fF
C174 VPB.n124 VNB 0.02fF
C175 VPB.n125 VNB 0.02fF
C176 VPB.n126 VNB 0.02fF
C177 VPB.n127 VNB 0.04fF
C178 VPB.n128 VNB 0.04fF
C179 VPB.n130 VNB 0.02fF
C180 VPB.n131 VNB 0.02fF
C181 VPB.n132 VNB 0.02fF
C182 VPB.n134 VNB 0.02fF
C183 VPB.n135 VNB 0.02fF
C184 VPB.n136 VNB 0.02fF
C185 VPB.n137 VNB 0.02fF
C186 VPB.n139 VNB 0.04fF
C187 VPB.n140 VNB 0.02fF
C188 VPB.n141 VNB 0.14fF
C189 VPB.n143 VNB 0.42fF
C190 VPB.n144 VNB 0.14fF
C191 VPB.n145 VNB 0.03fF
C192 VPB.n146 VNB 0.03fF
C193 VPB.n147 VNB 0.03fF
C194 VPB.n148 VNB 0.06fF
C195 VPB.n149 VNB 0.23fF
C196 VPB.n150 VNB 0.02fF
C197 VPB.n151 VNB 0.01fF
C198 VPB.n152 VNB 0.02fF
C199 VPB.n153 VNB 0.13fF
C200 VPB.n154 VNB 0.16fF
C201 VPB.n155 VNB 0.02fF
C202 VPB.n156 VNB 0.02fF
C203 VPB.n157 VNB 0.02fF
C204 VPB.n158 VNB 0.13fF
C205 VPB.n159 VNB 0.15fF
C206 VPB.n160 VNB 0.02fF
C207 VPB.n161 VNB 0.02fF
C208 VPB.n162 VNB 0.02fF
C209 VPB.n163 VNB 0.10fF
C210 VPB.n164 VNB 0.02fF
C211 VPB.n165 VNB 0.13fF
C212 VPB.n166 VNB 0.15fF
C213 VPB.n167 VNB 0.02fF
C214 VPB.n168 VNB 0.02fF
C215 VPB.n169 VNB 0.02fF
C216 VPB.n170 VNB 0.13fF
C217 VPB.n171 VNB 0.16fF
C218 VPB.n172 VNB 0.02fF
C219 VPB.n173 VNB 0.02fF
C220 VPB.n174 VNB 0.02fF
C221 VPB.n175 VNB 0.06fF
C222 VPB.n176 VNB 0.23fF
C223 VPB.n177 VNB 0.02fF
C224 VPB.n178 VNB 0.01fF
C225 VPB.n179 VNB 0.02fF
C226 VPB.n180 VNB 0.27fF
C227 VPB.n181 VNB 0.01fF
C228 VPB.n182 VNB 0.02fF
C229 VPB.n183 VNB 0.04fF
C230 VPB.n184 VNB 0.02fF
C231 VPB.n185 VNB 0.02fF
C232 VPB.n186 VNB 0.02fF
C233 VPB.n187 VNB 0.20fF
C234 VPB.n188 VNB 0.04fF
C235 VPB.n189 VNB 0.03fF
C236 VPB.n190 VNB 0.02fF
C237 VPB.n191 VNB 0.02fF
C238 VPB.n192 VNB 0.02fF
C239 VPB.n193 VNB 0.03fF
C240 VPB.n194 VNB 0.02fF
C241 VPB.n196 VNB 0.02fF
C242 VPB.n197 VNB 0.02fF
C243 VPB.n198 VNB 0.02fF
C244 VPB.n200 VNB 0.27fF
C245 VPB.n202 VNB 0.03fF
C246 VPB.n203 VNB 0.02fF
C247 VPB.n204 VNB 0.03fF
C248 VPB.n205 VNB 0.03fF
C249 VPB.n206 VNB 0.27fF
C250 VPB.n207 VNB 0.01fF
C251 VPB.n208 VNB 0.02fF
C252 VPB.n209 VNB 0.04fF
C253 VPB.n210 VNB 0.27fF
C254 VPB.n211 VNB 0.02fF
C255 VPB.n212 VNB 0.02fF
C256 VPB.n213 VNB 0.02fF
C257 VPB.n214 VNB 0.27fF
C258 VPB.n215 VNB 0.02fF
C259 VPB.n216 VNB 0.02fF
C260 VPB.n217 VNB 0.02fF
C261 VPB.n218 VNB 0.27fF
C262 VPB.n219 VNB 0.02fF
C263 VPB.n220 VNB 0.02fF
C264 VPB.n221 VNB 0.02fF
C265 VPB.n222 VNB 0.27fF
C266 VPB.n223 VNB 0.02fF
C267 VPB.n224 VNB 0.02fF
C268 VPB.n225 VNB 0.02fF
C269 VPB.n226 VNB 0.27fF
C270 VPB.n227 VNB 0.02fF
C271 VPB.n228 VNB 0.02fF
C272 VPB.n229 VNB 0.02fF
C273 VPB.n230 VNB 0.27fF
C274 VPB.n231 VNB 0.02fF
C275 VPB.n232 VNB 0.02fF
C276 VPB.n233 VNB 0.02fF
.ends
