// File: HA.spi.pex
// Created: Tue Oct 15 15:49:12 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_HA\%GND ( 1 29 33 36 41 49 52 57 61 83 87 90 95 99 107 115 121 127 \
 132 137 141 154 166 178 180 183 188 195 196 197 198 199 200 )
c249 ( 200 0 ) capacitor c=0.0583152f //x=14.925 //y=0.37
c250 ( 199 0 ) capacitor c=0.0210151f //x=12.09 //y=0.87
c251 ( 198 0 ) capacitor c=0.0210151f //x=8.76 //y=0.87
c252 ( 197 0 ) capacitor c=0.0572847f //x=6.045 //y=0.37
c253 ( 196 0 ) capacitor c=0.0578714f //x=3.825 //y=0.37
c254 ( 195 0 ) capacitor c=0.0208198f //x=0.99 //y=0.865
c255 ( 188 0 ) capacitor c=0.229233f //x=16.02 //y=0
c256 ( 183 0 ) capacitor c=0.103612f //x=14.43 //y=0
c257 ( 182 0 ) capacitor c=0.0044012f //x=12.21 //y=0
c258 ( 180 0 ) capacitor c=0.104587f //x=11.1 //y=0
c259 ( 179 0 ) capacitor c=0.0044012f //x=8.95 //y=0
c260 ( 178 0 ) capacitor c=0.102385f //x=7.77 //y=0
c261 ( 166 0 ) capacitor c=0.0972387f //x=5.55 //y=0
c262 ( 154 0 ) capacitor c=0.10149f //x=3.33 //y=0
c263 ( 153 0 ) capacitor c=0.00440095f //x=1.18 //y=0
c264 ( 144 0 ) capacitor c=0.00592191f //x=16.02 //y=0.45
c265 ( 141 0 ) capacitor c=0.00644318f //x=15.935 //y=0.535
c266 ( 140 0 ) capacitor c=0.00479856f //x=15.535 //y=0.45
c267 ( 137 0 ) capacitor c=0.00531808f //x=15.45 //y=0.535
c268 ( 132 0 ) capacitor c=0.00587411f //x=15.05 //y=0.45
c269 ( 127 0 ) capacitor c=0.0160123f //x=14.965 //y=0
c270 ( 121 0 ) capacitor c=0.0720515f //x=14.26 //y=0
c271 ( 115 0 ) capacitor c=0.0389232f //x=12.195 //y=0
c272 ( 107 0 ) capacitor c=0.072035f //x=10.93 //y=0
c273 ( 99 0 ) capacitor c=0.0389232f //x=8.865 //y=0
c274 ( 96 0 ) capacitor c=0.0360673f //x=7.235 //y=0
c275 ( 95 0 ) capacitor c=0.0160123f //x=7.6 //y=0
c276 ( 90 0 ) capacitor c=0.00587411f //x=7.15 //y=0.45
c277 ( 87 0 ) capacitor c=0.00531771f //x=7.065 //y=0.535
c278 ( 86 0 ) capacitor c=0.00479856f //x=6.665 //y=0.45
c279 ( 83 0 ) capacitor c=0.00643449f //x=6.58 //y=0.535
c280 ( 78 0 ) capacitor c=0.00592191f //x=6.18 //y=0.45
c281 ( 73 0 ) capacitor c=0.0190475f //x=6.095 //y=0
c282 ( 70 0 ) capacitor c=0.0360689f //x=5.015 //y=0
c283 ( 69 0 ) capacitor c=0.0184787f //x=5.38 //y=0
c284 ( 64 0 ) capacitor c=0.00583665f //x=4.93 //y=0.45
c285 ( 61 0 ) capacitor c=0.00536917f //x=4.845 //y=0.535
c286 ( 60 0 ) capacitor c=0.00479856f //x=4.445 //y=0.45
c287 ( 57 0 ) capacitor c=0.00640467f //x=4.36 //y=0.535
c288 ( 52 0 ) capacitor c=0.00588377f //x=3.96 //y=0.45
c289 ( 49 0 ) capacitor c=0.0164879f //x=3.875 //y=0
c290 ( 41 0 ) capacitor c=0.0720403f //x=3.16 //y=0
c291 ( 36 0 ) capacitor c=0.179504f //x=0.74 //y=0
c292 ( 33 0 ) capacitor c=0.0426751f //x=1.095 //y=0
c293 ( 29 0 ) capacitor c=0.566732f //x=15.91 //y=0
r294 (  187 188 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=15.91 //y=0 //x2=16.02 //y2=0
r295 (  185 187 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=15.535 //y=0 //x2=15.91 //y2=0
r296 (  184 185 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.05 //y=0 //x2=15.535 //y2=0
r297 (  170 171 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=7.03 //y=0 //x2=7.15 //y2=0
r298 (  168 170 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=6.665 //y=0 //x2=7.03 //y2=0
r299 (  167 168 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.18 //y=0 //x2=6.665 //y2=0
r300 (  158 159 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.445 //y=0 //x2=4.93 //y2=0
r301 (  157 158 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=4.44 //y=0 //x2=4.445 //y2=0
r302 (  155 157 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=3.96 //y=0 //x2=4.44 //y2=0
r303 (  145 200 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.02 //y=0.62 //x2=16.02 //y2=0.535
r304 (  145 200 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=16.02 //y=0.62 //x2=16.02 //y2=1.225
r305 (  144 200 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.02 //y=0.45 //x2=16.02 //y2=0.535
r306 (  143 188 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.02 //y=0.17 //x2=16.02 //y2=0
r307 (  143 144 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=16.02 //y=0.17 //x2=16.02 //y2=0.45
r308 (  142 200 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.62 //y=0.535 //x2=15.535 //y2=0.535
r309 (  141 200 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.935 //y=0.535 //x2=16.02 //y2=0.535
r310 (  141 142 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=15.935 //y=0.535 //x2=15.62 //y2=0.535
r311 (  140 200 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.535 //y=0.45 //x2=15.535 //y2=0.535
r312 (  139 185 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.535 //y=0.17 //x2=15.535 //y2=0
r313 (  139 140 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=15.535 //y=0.17 //x2=15.535 //y2=0.45
r314 (  138 200 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.135 //y=0.535 //x2=15.05 //y2=0.535
r315 (  137 200 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.45 //y=0.535 //x2=15.535 //y2=0.535
r316 (  137 138 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=15.45 //y=0.535 //x2=15.135 //y2=0.535
r317 (  133 200 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.05 //y=0.62 //x2=15.05 //y2=0.535
r318 (  133 200 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=15.05 //y=0.62 //x2=15.05 //y2=1.225
r319 (  132 200 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.05 //y=0.45 //x2=15.05 //y2=0.535
r320 (  131 184 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.05 //y=0.17 //x2=15.05 //y2=0
r321 (  131 132 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=15.05 //y=0.17 //x2=15.05 //y2=0.45
r322 (  128 183 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=14.43 //y2=0
r323 (  128 130 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=14.8 //y2=0
r324 (  127 184 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.965 //y=0 //x2=15.05 //y2=0
r325 (  127 130 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=14.965 //y=0 //x2=14.8 //y2=0
r326 (  122 182 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.365 //y=0 //x2=12.28 //y2=0
r327 (  122 124 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=12.365 //y=0 //x2=13.32 //y2=0
r328 (  121 183 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=14.43 //y2=0
r329 (  121 124 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=13.32 //y2=0
r330 (  117 182 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.28 //y=0.17 //x2=12.28 //y2=0
r331 (  117 199 ) resistor r=54.0749 //w=0.187 //l=0.79 //layer=li \
 //thickness=0.1 //x=12.28 //y=0.17 //x2=12.28 //y2=0.96
r332 (  116 180 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.27 //y=0 //x2=11.1 //y2=0
r333 (  115 182 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.195 //y=0 //x2=12.28 //y2=0
r334 (  115 116 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=12.195 //y=0 //x2=11.27 //y2=0
r335 (  110 112 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=9.62 //y=0 //x2=10.73 //y2=0
r336 (  108 179 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.035 //y=0 //x2=8.95 //y2=0
r337 (  108 110 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=9.035 //y=0 //x2=9.62 //y2=0
r338 (  107 180 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.93 //y=0 //x2=11.1 //y2=0
r339 (  107 112 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=10.93 //y=0 //x2=10.73 //y2=0
r340 (  103 179 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.95 //y=0.17 //x2=8.95 //y2=0
r341 (  103 198 ) resistor r=54.0749 //w=0.187 //l=0.79 //layer=li \
 //thickness=0.1 //x=8.95 //y=0.17 //x2=8.95 //y2=0.96
r342 (  100 178 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.94 //y=0 //x2=7.77 //y2=0
r343 (  100 102 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=7.94 //y=0 //x2=8.51 //y2=0
r344 (  99 179 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.865 //y=0 //x2=8.95 //y2=0
r345 (  99 102 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=8.865 //y=0 //x2=8.51 //y2=0
r346 (  96 171 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.235 //y=0 //x2=7.15 //y2=0
r347 (  95 178 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.6 //y=0 //x2=7.77 //y2=0
r348 (  95 96 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=7.6 //y=0 //x2=7.235 //y2=0
r349 (  91 197 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.62 //x2=7.15 //y2=0.535
r350 (  91 197 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.62 //x2=7.15 //y2=1.225
r351 (  90 197 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.45 //x2=7.15 //y2=0.535
r352 (  89 171 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.17 //x2=7.15 //y2=0
r353 (  89 90 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=7.15 //y=0.17 //x2=7.15 //y2=0.45
r354 (  88 197 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.75 //y=0.535 //x2=6.665 //y2=0.535
r355 (  87 197 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.065 //y=0.535 //x2=7.15 //y2=0.535
r356 (  87 88 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=7.065 //y=0.535 //x2=6.75 //y2=0.535
r357 (  86 197 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.665 //y=0.45 //x2=6.665 //y2=0.535
r358 (  85 168 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.665 //y=0.17 //x2=6.665 //y2=0
r359 (  85 86 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=6.665 //y=0.17 //x2=6.665 //y2=0.45
r360 (  84 197 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.265 //y=0.535 //x2=6.18 //y2=0.535
r361 (  83 197 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.58 //y=0.535 //x2=6.665 //y2=0.535
r362 (  83 84 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=6.58 //y=0.535 //x2=6.265 //y2=0.535
r363 (  79 197 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.62 //x2=6.18 //y2=0.535
r364 (  79 197 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.62 //x2=6.18 //y2=1.225
r365 (  78 197 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.45 //x2=6.18 //y2=0.535
r366 (  77 167 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.17 //x2=6.18 //y2=0
r367 (  77 78 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=6.18 //y=0.17 //x2=6.18 //y2=0.45
r368 (  74 166 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.55 //y2=0
r369 (  74 76 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.92 //y2=0
r370 (  73 167 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.095 //y=0 //x2=6.18 //y2=0
r371 (  73 76 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=6.095 //y=0 //x2=5.92 //y2=0
r372 (  70 159 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.015 //y=0 //x2=4.93 //y2=0
r373 (  69 166 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=5.55 //y2=0
r374 (  69 70 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=5.015 //y2=0
r375 (  65 196 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.62 //x2=4.93 //y2=0.535
r376 (  65 196 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.62 //x2=4.93 //y2=1.225
r377 (  64 196 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.45 //x2=4.93 //y2=0.535
r378 (  63 159 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.17 //x2=4.93 //y2=0
r379 (  63 64 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.17 //x2=4.93 //y2=0.45
r380 (  62 196 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.53 //y=0.535 //x2=4.445 //y2=0.535
r381 (  61 196 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.845 //y=0.535 //x2=4.93 //y2=0.535
r382 (  61 62 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.845 //y=0.535 //x2=4.53 //y2=0.535
r383 (  60 196 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.45 //x2=4.445 //y2=0.535
r384 (  59 158 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.17 //x2=4.445 //y2=0
r385 (  59 60 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.17 //x2=4.445 //y2=0.45
r386 (  58 196 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.045 //y=0.535 //x2=3.96 //y2=0.535
r387 (  57 196 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.36 //y=0.535 //x2=4.445 //y2=0.535
r388 (  57 58 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.36 //y=0.535 //x2=4.045 //y2=0.535
r389 (  53 196 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.62 //x2=3.96 //y2=0.535
r390 (  53 196 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.62 //x2=3.96 //y2=1.225
r391 (  52 196 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.45 //x2=3.96 //y2=0.535
r392 (  51 155 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.17 //x2=3.96 //y2=0
r393 (  51 52 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.17 //x2=3.96 //y2=0.45
r394 (  50 154 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=0 //x2=3.33 //y2=0
r395 (  49 155 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.875 //y=0 //x2=3.96 //y2=0
r396 (  49 50 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=3.875 //y=0 //x2=3.5 //y2=0
r397 (  44 46 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r398 (  42 153 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.18 //y2=0
r399 (  42 44 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.85 //y2=0
r400 (  41 154 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=3.33 //y2=0
r401 (  41 46 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r402 (  37 153 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r403 (  37 195 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.955
r404 (  33 153 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=1.18 //y2=0
r405 (  33 36 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=0.74 //y2=0
r406 (  29 187 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.91 //y=0 //x2=15.91 //y2=0
r407 (  27 130 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.8 //y=0 //x2=14.8 //y2=0
r408 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.8 //y=0 //x2=15.91 //y2=0
r409 (  25 124 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.32 //y=0 //x2=13.32 //y2=0
r410 (  25 27 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=13.32 //y=0 //x2=14.8 //y2=0
r411 (  23 182 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.21 //y=0 //x2=12.21 //y2=0
r412 (  23 25 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=0 //x2=13.32 //y2=0
r413 (  21 112 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=0 //x2=10.73 //y2=0
r414 (  21 23 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=0 //x2=12.21 //y2=0
r415 (  19 110 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=0 //x2=9.62 //y2=0
r416 (  19 21 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.62 //y=0 //x2=10.73 //y2=0
r417 (  17 102 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.51 //y=0 //x2=8.51 //y2=0
r418 (  17 19 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.51 //y=0 //x2=9.62 //y2=0
r419 (  14 170 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=0 //x2=7.03 //y2=0
r420 (  12 76 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=0 //x2=5.92 //y2=0
r421 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=0 //x2=7.03 //y2=0
r422 (  10 157 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r423 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.92 //y2=0
r424 (  8 46 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r425 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r426 (  6 44 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r427 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r428 (  3 36 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r429 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r430 (  1 17 ) resistor r=0.0768272 //w=0.301 //l=0.185 //layer=m1 \
 //thickness=0.36 //x=8.325 //y=0 //x2=8.51 //y2=0
r431 (  1 14 ) resistor r=0.537791 //w=0.301 //l=1.295 //layer=m1 \
 //thickness=0.36 //x=8.325 //y=0 //x2=7.03 //y2=0
ends PM_HA\%GND

subckt PM_HA\%VDD ( 1 29 41 49 59 65 73 83 87 97 105 109 117 125 133 139 149 \
 162 165 168 172 174 176 179 180 181 182 183 184 185 186 187 188 189 190 )
c238 ( 190 0 ) capacitor c=0.0420685f //x=15.83 //y=5.02
c239 ( 189 0 ) capacitor c=0.0433633f //x=14.97 //y=5.02
c240 ( 188 0 ) capacitor c=0.0266033f //x=12.185 //y=5.02
c241 ( 187 0 ) capacitor c=0.0265042f //x=8.855 //y=5.02
c242 ( 186 0 ) capacitor c=0.0432963f //x=6.96 //y=5.02
c243 ( 185 0 ) capacitor c=0.0420333f //x=6.09 //y=5.02
c244 ( 184 0 ) capacitor c=0.0432963f //x=4.74 //y=5.02
c245 ( 183 0 ) capacitor c=0.0422219f //x=3.87 //y=5.02
c246 ( 182 0 ) capacitor c=0.0381505f //x=2.405 //y=5.02
c247 ( 181 0 ) capacitor c=0.0240879f //x=1.525 //y=5.02
c248 ( 180 0 ) capacitor c=0.053196f //x=0.655 //y=5.02
c249 ( 179 0 ) capacitor c=0.232571f //x=15.91 //y=7.4
c250 ( 177 0 ) capacitor c=0.00591168f //x=15.095 //y=7.4
c251 ( 176 0 ) capacitor c=0.105702f //x=14.43 //y=7.4
c252 ( 175 0 ) capacitor c=0.00591168f //x=12.33 //y=7.4
c253 ( 174 0 ) capacitor c=0.110106f //x=11.1 //y=7.4
c254 ( 173 0 ) capacitor c=0.00591168f //x=9 //y=7.4
c255 ( 172 0 ) capacitor c=0.110701f //x=7.77 //y=7.4
c256 ( 171 0 ) capacitor c=0.00591168f //x=7.03 //y=7.4
c257 ( 169 0 ) capacitor c=0.00591168f //x=6.225 //y=7.4
c258 ( 168 0 ) capacitor c=0.1056f //x=5.55 //y=7.4
c259 ( 167 0 ) capacitor c=0.00591168f //x=4.885 //y=7.4
c260 ( 166 0 ) capacitor c=0.00591168f //x=4.005 //y=7.4
c261 ( 165 0 ) capacitor c=0.108116f //x=3.33 //y=7.4
c262 ( 164 0 ) capacitor c=0.00591168f //x=2.55 //y=7.4
c263 ( 163 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c264 ( 162 0 ) capacitor c=0.248183f //x=0.74 //y=7.4
c265 ( 149 0 ) capacitor c=0.0289356f //x=15.89 //y=7.4
c266 ( 139 0 ) capacitor c=0.0181526f //x=15.01 //y=7.4
c267 ( 133 0 ) capacitor c=0.0747638f //x=14.26 //y=7.4
c268 ( 125 0 ) capacitor c=0.0428656f //x=12.245 //y=7.4
c269 ( 117 0 ) capacitor c=0.0750963f //x=10.93 //y=7.4
c270 ( 109 0 ) capacitor c=0.042884f //x=8.915 //y=7.4
c271 ( 105 0 ) capacitor c=0.0181526f //x=7.6 //y=7.4
c272 ( 97 0 ) capacitor c=0.0291066f //x=7.02 //y=7.4
c273 ( 87 0 ) capacitor c=0.0186283f //x=6.14 //y=7.4
c274 ( 83 0 ) capacitor c=0.0181526f //x=5.38 //y=7.4
c275 ( 73 0 ) capacitor c=0.0289624f //x=4.8 //y=7.4
c276 ( 65 0 ) capacitor c=0.0186283f //x=3.92 //y=7.4
c277 ( 59 0 ) capacitor c=0.0236224f //x=3.16 //y=7.4
c278 ( 49 0 ) capacitor c=0.0288639f //x=2.465 //y=7.4
c279 ( 41 0 ) capacitor c=0.028955f //x=1.585 //y=7.4
c280 ( 29 0 ) capacitor c=0.581105f //x=15.91 //y=7.4
r281 (  151 179 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.975 //y=7.23 //x2=15.975 //y2=7.4
r282 (  151 190 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=15.975 //y=7.23 //x2=15.975 //y2=6.405
r283 (  150 177 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.18 //y=7.4 //x2=15.095 //y2=7.4
r284 (  149 179 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.89 //y=7.4 //x2=15.975 //y2=7.4
r285 (  149 150 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=15.89 //y=7.4 //x2=15.18 //y2=7.4
r286 (  143 177 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.095 //y=7.23 //x2=15.095 //y2=7.4
r287 (  143 189 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=15.095 //y=7.23 //x2=15.095 //y2=6.405
r288 (  140 176 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=14.43 //y2=7.4
r289 (  140 142 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=14.8 //y2=7.4
r290 (  139 177 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.01 //y=7.4 //x2=15.095 //y2=7.4
r291 (  139 142 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=15.01 //y=7.4 //x2=14.8 //y2=7.4
r292 (  134 175 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.415 //y=7.4 //x2=12.33 //y2=7.4
r293 (  134 136 ) resistor r=32.4482 //w=0.357 //l=0.905 //layer=li \
 //thickness=0.1 //x=12.415 //y=7.4 //x2=13.32 //y2=7.4
r294 (  133 176 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=14.43 //y2=7.4
r295 (  133 136 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=13.32 //y2=7.4
r296 (  129 175 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.33 //y=7.23 //x2=12.33 //y2=7.4
r297 (  129 188 ) resistor r=80.4278 //w=0.187 //l=1.175 //layer=li \
 //thickness=0.1 //x=12.33 //y=7.23 //x2=12.33 //y2=6.055
r298 (  126 174 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.27 //y=7.4 //x2=11.1 //y2=7.4
r299 (  126 128 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=11.27 //y=7.4 //x2=12.21 //y2=7.4
r300 (  125 175 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.245 //y=7.4 //x2=12.33 //y2=7.4
r301 (  125 128 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=12.245 //y=7.4 //x2=12.21 //y2=7.4
r302 (  120 122 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=9.62 //y=7.4 //x2=10.73 //y2=7.4
r303 (  118 173 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.085 //y=7.4 //x2=9 //y2=7.4
r304 (  118 120 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=9.085 //y=7.4 //x2=9.62 //y2=7.4
r305 (  117 174 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.93 //y=7.4 //x2=11.1 //y2=7.4
r306 (  117 122 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=10.93 //y=7.4 //x2=10.73 //y2=7.4
r307 (  113 173 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9 //y=7.23 //x2=9 //y2=7.4
r308 (  113 187 ) resistor r=80.4278 //w=0.187 //l=1.175 //layer=li \
 //thickness=0.1 //x=9 //y=7.23 //x2=9 //y2=6.055
r309 (  110 172 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.94 //y=7.4 //x2=7.77 //y2=7.4
r310 (  110 112 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=7.94 //y=7.4 //x2=8.51 //y2=7.4
r311 (  109 173 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.915 //y=7.4 //x2=9 //y2=7.4
r312 (  109 112 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=8.915 //y=7.4 //x2=8.51 //y2=7.4
r313 (  106 171 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.19 //y=7.4 //x2=7.105 //y2=7.4
r314 (  105 172 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.6 //y=7.4 //x2=7.77 //y2=7.4
r315 (  105 106 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=7.6 //y=7.4 //x2=7.19 //y2=7.4
r316 (  99 171 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.105 //y=7.23 //x2=7.105 //y2=7.4
r317 (  99 186 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=7.105 //y=7.23 //x2=7.105 //y2=6.405
r318 (  98 169 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.31 //y=7.4 //x2=6.225 //y2=7.4
r319 (  97 171 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.02 //y=7.4 //x2=7.105 //y2=7.4
r320 (  97 98 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.02 //y=7.4 //x2=6.31 //y2=7.4
r321 (  91 169 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.225 //y=7.23 //x2=6.225 //y2=7.4
r322 (  91 185 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=6.225 //y=7.23 //x2=6.225 //y2=6.405
r323 (  88 168 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.55 //y2=7.4
r324 (  88 90 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.92 //y2=7.4
r325 (  87 169 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.14 //y=7.4 //x2=6.225 //y2=7.4
r326 (  87 90 ) resistor r=7.88796 //w=0.357 //l=0.22 //layer=li \
 //thickness=0.1 //x=6.14 //y=7.4 //x2=5.92 //y2=7.4
r327 (  84 167 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.97 //y=7.4 //x2=4.885 //y2=7.4
r328 (  83 168 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=5.55 //y2=7.4
r329 (  83 84 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=4.97 //y2=7.4
r330 (  77 167 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.885 //y=7.23 //x2=4.885 //y2=7.4
r331 (  77 184 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.885 //y=7.23 //x2=4.885 //y2=6.405
r332 (  74 166 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.09 //y=7.4 //x2=4.005 //y2=7.4
r333 (  74 76 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li \
 //thickness=0.1 //x=4.09 //y=7.4 //x2=4.44 //y2=7.4
r334 (  73 167 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.8 //y=7.4 //x2=4.885 //y2=7.4
r335 (  73 76 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=4.8 //y=7.4 //x2=4.44 //y2=7.4
r336 (  67 166 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.005 //y=7.23 //x2=4.005 //y2=7.4
r337 (  67 183 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.005 //y=7.23 //x2=4.005 //y2=6.405
r338 (  66 165 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r339 (  65 166 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.92 //y=7.4 //x2=4.005 //y2=7.4
r340 (  65 66 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=3.92 //y=7.4 //x2=3.5 //y2=7.4
r341 (  60 164 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.55 //y2=7.4
r342 (  60 62 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.96 //y2=7.4
r343 (  59 165 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r344 (  59 62 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r345 (  53 164 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r346 (  53 182 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.745
r347 (  50 163 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r348 (  50 52 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r349 (  49 164 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r350 (  49 52 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r351 (  43 163 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r352 (  43 181 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.745
r353 (  42 162 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r354 (  41 163 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r355 (  41 42 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r356 (  35 162 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r357 (  35 180 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.405
r358 (  29 179 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.91 //y=7.4 //x2=15.91 //y2=7.4
r359 (  27 142 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.8 //y=7.4 //x2=14.8 //y2=7.4
r360 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.8 //y=7.4 //x2=15.91 //y2=7.4
r361 (  25 136 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.32 //y=7.4 //x2=13.32 //y2=7.4
r362 (  25 27 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=13.32 //y=7.4 //x2=14.8 //y2=7.4
r363 (  23 128 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.21 //y=7.4 //x2=12.21 //y2=7.4
r364 (  23 25 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=7.4 //x2=13.32 //y2=7.4
r365 (  21 122 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=7.4 //x2=10.73 //y2=7.4
r366 (  21 23 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=7.4 //x2=12.21 //y2=7.4
r367 (  19 120 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=7.4 //x2=9.62 //y2=7.4
r368 (  19 21 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.62 //y=7.4 //x2=10.73 //y2=7.4
r369 (  17 112 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.51 //y=7.4 //x2=8.51 //y2=7.4
r370 (  17 19 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.51 //y=7.4 //x2=9.62 //y2=7.4
r371 (  14 171 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=7.4 //x2=7.03 //y2=7.4
r372 (  12 90 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=7.4 //x2=5.92 //y2=7.4
r373 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=7.4 //x2=7.03 //y2=7.4
r374 (  10 76 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r375 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.92 //y2=7.4
r376 (  8 62 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r377 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r378 (  6 52 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r379 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r380 (  3 162 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r381 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r382 (  1 17 ) resistor r=0.0768272 //w=0.301 //l=0.185 //layer=m1 \
 //thickness=0.36 //x=8.325 //y=7.4 //x2=8.51 //y2=7.4
r383 (  1 14 ) resistor r=0.537791 //w=0.301 //l=1.295 //layer=m1 \
 //thickness=0.36 //x=8.325 //y=7.4 //x2=7.03 //y2=7.4
ends PM_HA\%VDD

subckt PM_HA\%noxref_3 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 52 \
 53 54 56 62 63 65 73 75 76 )
c142 ( 76 0 ) capacitor c=0.0220291f //x=1.965 //y=5.02
c143 ( 75 0 ) capacitor c=0.0217503f //x=1.085 //y=5.02
c144 ( 73 0 ) capacitor c=0.0084702f //x=1.96 //y=0.905
c145 ( 65 0 ) capacitor c=0.0528806f //x=4.07 //y=2.085
c146 ( 63 0 ) capacitor c=0.0435629f //x=4.71 //y=1.255
c147 ( 62 0 ) capacitor c=0.0200386f //x=4.71 //y=0.91
c148 ( 56 0 ) capacitor c=0.0152946f //x=4.555 //y=1.41
c149 ( 54 0 ) capacitor c=0.0157804f //x=4.555 //y=0.755
c150 ( 53 0 ) capacitor c=0.0490829f //x=4.3 //y=4.79
c151 ( 52 0 ) capacitor c=0.0304104f //x=4.59 //y=4.79
c152 ( 48 0 ) capacitor c=0.0290017f //x=4.18 //y=1.92
c153 ( 47 0 ) capacitor c=0.0250027f //x=4.18 //y=1.565
c154 ( 46 0 ) capacitor c=0.0234316f //x=4.18 //y=1.255
c155 ( 45 0 ) capacitor c=0.0200596f //x=4.18 //y=0.91
c156 ( 44 0 ) capacitor c=0.154218f //x=4.665 //y=6.02
c157 ( 43 0 ) capacitor c=0.154243f //x=4.225 //y=6.02
c158 ( 41 0 ) capacitor c=0.0023043f //x=2.11 //y=5.2
c159 ( 34 0 ) capacitor c=0.0891812f //x=4.07 //y=2.085
c160 ( 32 0 ) capacitor c=0.107172f //x=2.59 //y=3.33
c161 ( 28 0 ) capacitor c=0.00525782f //x=2.235 //y=1.655
c162 ( 27 0 ) capacitor c=0.0139525f //x=2.505 //y=1.655
c163 ( 25 0 ) capacitor c=0.0141863f //x=2.505 //y=5.2
c164 ( 14 0 ) capacitor c=0.00260571f //x=1.315 //y=5.2
c165 ( 13 0 ) capacitor c=0.0149571f //x=2.025 //y=5.2
c166 ( 2 0 ) capacitor c=0.0136218f //x=2.705 //y=3.33
c167 ( 1 0 ) capacitor c=0.0547127f //x=3.955 //y=3.33
r168 (  65 66 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.07 //y=2.085 //x2=4.18 //y2=2.085
r169 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.71 //y=1.255 //x2=4.67 //y2=1.41
r170 (  62 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.71 //y=0.91 //x2=4.67 //y2=0.755
r171 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.71 //y=0.91 //x2=4.71 //y2=1.255
r172 (  57 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.335 //y=1.41 //x2=4.22 //y2=1.41
r173 (  56 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.555 //y=1.41 //x2=4.67 //y2=1.41
r174 (  55 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.335 //y=0.755 //x2=4.22 //y2=0.755
r175 (  54 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.555 //y=0.755 //x2=4.67 //y2=0.755
r176 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.555 //y=0.755 //x2=4.335 //y2=0.755
r177 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.59 //y=4.79 //x2=4.665 //y2=4.865
r178 (  52 53 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=4.59 //y=4.79 //x2=4.3 //y2=4.79
r179 (  49 53 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.225 //y=4.865 //x2=4.3 //y2=4.79
r180 (  49 68 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=4.225 //y=4.865 //x2=4.07 //y2=4.7
r181 (  48 66 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.92 //x2=4.18 //y2=2.085
r182 (  47 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.565 //x2=4.22 //y2=1.41
r183 (  47 48 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.565 //x2=4.18 //y2=1.92
r184 (  46 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.255 //x2=4.22 //y2=1.41
r185 (  45 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=0.91 //x2=4.22 //y2=0.755
r186 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.18 //y=0.91 //x2=4.18 //y2=1.255
r187 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.665 //y=6.02 //x2=4.665 //y2=4.865
r188 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.225 //y=6.02 //x2=4.225 //y2=4.865
r189 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.445 //y=1.41 //x2=4.555 //y2=1.41
r190 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.445 //y=1.41 //x2=4.335 //y2=1.41
r191 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=4.7 //x2=4.07 //y2=4.7
r192 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=3.33 //x2=4.07 //y2=4.7
r193 (  34 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=2.085 //x2=4.07 //y2=2.085
r194 (  34 37 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=4.07 //y=2.085 //x2=4.07 //y2=3.33
r195 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.115 //x2=2.59 //y2=3.33
r196 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=3.33
r197 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r198 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r199 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.195 //y=5.2 //x2=2.11 //y2=5.2
r200 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.59 //y2=5.115
r201 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.195 //y2=5.2
r202 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.235 //y2=1.655
r203 (  21 73 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r204 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.2
r205 (  15 76 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.725
r206 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=2.11 //y2=5.2
r207 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=1.315 //y2=5.2
r208 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.315 //y2=5.2
r209 (  7 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.23 //y2=5.725
r210 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.33 //x2=4.07 //y2=3.33
r211 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=3.33 //x2=2.59 //y2=3.33
r212 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=3.33 //x2=2.59 //y2=3.33
r213 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.955 //y=3.33 //x2=4.07 //y2=3.33
r214 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=3.955 //y=3.33 //x2=2.705 //y2=3.33
ends PM_HA\%noxref_3

subckt PM_HA\%A ( 1 2 3 4 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 27 40 \
 52 62 63 64 65 66 67 68 69 70 71 72 73 74 78 80 83 84 88 89 90 91 95 96 97 99 \
 105 106 107 108 109 110 114 116 119 120 130 134 148 )
c234 ( 148 0 ) capacitor c=0.0615343f //x=8.88 //y=4.7
c235 ( 134 0 ) capacitor c=0.0537799f //x=6.29 //y=2.085
c236 ( 130 0 ) capacitor c=0.0598647f //x=1.11 //y=4.7
c237 ( 120 0 ) capacitor c=0.0318948f //x=9.215 //y=1.215
c238 ( 119 0 ) capacitor c=0.0187407f //x=9.215 //y=0.87
c239 ( 116 0 ) capacitor c=0.0141798f //x=9.06 //y=1.37
c240 ( 114 0 ) capacitor c=0.0149852f //x=9.06 //y=0.715
c241 ( 110 0 ) capacitor c=0.0836807f //x=8.685 //y=1.92
c242 ( 109 0 ) capacitor c=0.0229722f //x=8.685 //y=1.525
c243 ( 108 0 ) capacitor c=0.0234352f //x=8.685 //y=1.215
c244 ( 107 0 ) capacitor c=0.0199366f //x=8.685 //y=0.87
c245 ( 106 0 ) capacitor c=0.0435629f //x=6.93 //y=1.255
c246 ( 105 0 ) capacitor c=0.0200386f //x=6.93 //y=0.91
c247 ( 99 0 ) capacitor c=0.0152946f //x=6.775 //y=1.41
c248 ( 97 0 ) capacitor c=0.0157804f //x=6.775 //y=0.755
c249 ( 96 0 ) capacitor c=0.0490957f //x=6.52 //y=4.79
c250 ( 95 0 ) capacitor c=0.0303096f //x=6.81 //y=4.79
c251 ( 91 0 ) capacitor c=0.0290017f //x=6.4 //y=1.92
c252 ( 90 0 ) capacitor c=0.0250027f //x=6.4 //y=1.565
c253 ( 89 0 ) capacitor c=0.0234316f //x=6.4 //y=1.255
c254 ( 88 0 ) capacitor c=0.0200596f //x=6.4 //y=0.91
c255 ( 84 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c256 ( 83 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c257 ( 80 0 ) capacitor c=0.0141798f //x=1.29 //y=1.365
c258 ( 78 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c259 ( 74 0 ) capacitor c=0.0860049f //x=0.915 //y=1.915
c260 ( 73 0 ) capacitor c=0.0229722f //x=0.915 //y=1.52
c261 ( 72 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c262 ( 71 0 ) capacitor c=0.0199343f //x=0.915 //y=0.865
c263 ( 70 0 ) capacitor c=0.110797f //x=9.22 //y=6.02
c264 ( 69 0 ) capacitor c=0.154322f //x=8.78 //y=6.02
c265 ( 68 0 ) capacitor c=0.154218f //x=6.885 //y=6.02
c266 ( 67 0 ) capacitor c=0.154243f //x=6.445 //y=6.02
c267 ( 66 0 ) capacitor c=0.110275f //x=1.45 //y=6.02
c268 ( 65 0 ) capacitor c=0.154305f //x=1.01 //y=6.02
c269 ( 52 0 ) capacitor c=0.100543f //x=8.88 //y=2.085
c270 ( 40 0 ) capacitor c=0.0908218f //x=6.29 //y=2.085
c271 ( 27 0 ) capacitor c=0.112176f //x=1.11 //y=2.08
c272 ( 4 0 ) capacitor c=0.00595795f //x=6.405 //y=4.07
c273 ( 3 0 ) capacitor c=0.0693107f //x=8.765 //y=4.07
c274 ( 2 0 ) capacitor c=0.0159773f //x=1.225 //y=4.07
c275 ( 1 0 ) capacitor c=0.130577f //x=6.175 //y=4.07
r276 (  146 148 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=8.78 //y=4.7 //x2=8.88 //y2=4.7
r277 (  134 135 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.29 //y=2.085 //x2=6.4 //y2=2.085
r278 (  128 130 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.7 //x2=1.11 //y2=4.7
r279 (  121 148 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=9.22 //y=4.865 //x2=8.88 //y2=4.7
r280 (  120 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.215 //x2=9.175 //y2=1.37
r281 (  119 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.215 //y=0.87 //x2=9.175 //y2=0.715
r282 (  119 120 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.215 //y=0.87 //x2=9.215 //y2=1.215
r283 (  117 145 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.84 //y=1.37 //x2=8.725 //y2=1.37
r284 (  116 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.06 //y=1.37 //x2=9.175 //y2=1.37
r285 (  115 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.84 //y=0.715 //x2=8.725 //y2=0.715
r286 (  114 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.06 //y=0.715 //x2=9.175 //y2=0.715
r287 (  114 115 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=9.06 //y=0.715 //x2=8.84 //y2=0.715
r288 (  111 146 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.78 //y=4.865 //x2=8.78 //y2=4.7
r289 (  110 143 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=8.685 //y=1.92 //x2=8.88 //y2=2.085
r290 (  109 145 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.685 //y=1.525 //x2=8.725 //y2=1.37
r291 (  109 110 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=8.685 //y=1.525 //x2=8.685 //y2=1.92
r292 (  108 145 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.685 //y=1.215 //x2=8.725 //y2=1.37
r293 (  107 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.685 //y=0.87 //x2=8.725 //y2=0.715
r294 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.685 //y=0.87 //x2=8.685 //y2=1.215
r295 (  106 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.93 //y=1.255 //x2=6.89 //y2=1.41
r296 (  105 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.93 //y=0.91 //x2=6.89 //y2=0.755
r297 (  105 106 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.93 //y=0.91 //x2=6.93 //y2=1.255
r298 (  100 139 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.555 //y=1.41 //x2=6.44 //y2=1.41
r299 (  99 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.775 //y=1.41 //x2=6.89 //y2=1.41
r300 (  98 138 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.555 //y=0.755 //x2=6.44 //y2=0.755
r301 (  97 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.775 //y=0.755 //x2=6.89 //y2=0.755
r302 (  97 98 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.775 //y=0.755 //x2=6.555 //y2=0.755
r303 (  95 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.81 //y=4.79 //x2=6.885 //y2=4.865
r304 (  95 96 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=6.81 //y=4.79 //x2=6.52 //y2=4.79
r305 (  92 96 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.445 //y=4.865 //x2=6.52 //y2=4.79
r306 (  92 137 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=6.445 //y=4.865 //x2=6.29 //y2=4.7
r307 (  91 135 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.4 //y=1.92 //x2=6.4 //y2=2.085
r308 (  90 139 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.4 //y=1.565 //x2=6.44 //y2=1.41
r309 (  90 91 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=6.4 //y=1.565 //x2=6.4 //y2=1.92
r310 (  89 139 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.4 //y=1.255 //x2=6.44 //y2=1.41
r311 (  88 138 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.4 //y=0.91 //x2=6.44 //y2=0.755
r312 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.4 //y=0.91 //x2=6.4 //y2=1.255
r313 (  85 130 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=1.45 //y=4.865 //x2=1.11 //y2=4.7
r314 (  84 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r315 (  83 131 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r316 (  83 84 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r317 (  81 127 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r318 (  80 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r319 (  79 126 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r320 (  78 131 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r321 (  78 79 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r322 (  75 128 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.865 //x2=1.01 //y2=4.7
r323 (  74 125 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r324 (  73 127 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r325 (  73 74 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r326 (  72 127 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r327 (  71 126 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r328 (  71 72 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r329 (  70 121 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.22 //y=6.02 //x2=9.22 //y2=4.865
r330 (  69 111 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.78 //y=6.02 //x2=8.78 //y2=4.865
r331 (  68 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.885 //y=6.02 //x2=6.885 //y2=4.865
r332 (  67 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.445 //y=6.02 //x2=6.445 //y2=4.865
r333 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.02 //x2=1.45 //y2=4.865
r334 (  65 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.02 //x2=1.01 //y2=4.865
r335 (  64 116 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.37 //x2=9.06 //y2=1.37
r336 (  64 117 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.37 //x2=8.84 //y2=1.37
r337 (  63 99 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.665 //y=1.41 //x2=6.775 //y2=1.41
r338 (  63 100 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.665 //y=1.41 //x2=6.555 //y2=1.41
r339 (  62 80 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r340 (  62 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r341 (  60 148 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.88 //y=4.7 //x2=8.88 //y2=4.7
r342 (  52 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.88 //y=2.085 //x2=8.88 //y2=2.085
r343 (  49 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.29 //y=4.7 //x2=6.29 //y2=4.7
r344 (  40 134 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.29 //y=2.085 //x2=6.29 //y2=2.085
r345 (  37 130 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r346 (  27 125 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r347 (  25 60 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=8.88 //y=4.44 //x2=8.88 //y2=4.7
r348 (  24 25 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=8.88 //y=4.07 //x2=8.88 //y2=4.44
r349 (  23 24 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=8.88 //y=3.33 //x2=8.88 //y2=4.07
r350 (  22 23 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=8.88 //y=2.96 //x2=8.88 //y2=3.33
r351 (  22 52 ) resistor r=59.893 //w=0.187 //l=0.875 //layer=li \
 //thickness=0.1 //x=8.88 //y=2.96 //x2=8.88 //y2=2.085
r352 (  21 49 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=6.29 //y=4.44 //x2=6.29 //y2=4.7
r353 (  20 21 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=6.29 //y=4.07 //x2=6.29 //y2=4.44
r354 (  19 20 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=6.29 //y=3.33 //x2=6.29 //y2=4.07
r355 (  18 19 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=6.29 //y=2.96 //x2=6.29 //y2=3.33
r356 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=6.29 //y=2.59 //x2=6.29 //y2=2.96
r357 (  17 40 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=6.29 //y=2.59 //x2=6.29 //y2=2.085
r358 (  16 37 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.44 //x2=1.11 //y2=4.7
r359 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r360 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r361 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r362 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r363 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r364 (  11 27 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.59 //x2=1.11 //y2=2.08
r365 (  10 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.88 //y=4.07 //x2=8.88 //y2=4.07
r366 (  8 20 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.29 //y=4.07 //x2=6.29 //y2=4.07
r367 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.07
r368 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.405 //y=4.07 //x2=6.29 //y2=4.07
r369 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=4.07 //x2=8.88 //y2=4.07
r370 (  3 4 ) resistor r=2.25191 //w=0.131 //l=2.36 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=4.07 //x2=6.405 //y2=4.07
r371 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=4.07 //x2=1.11 //y2=4.07
r372 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.175 //y=4.07 //x2=6.29 //y2=4.07
r373 (  1 2 ) resistor r=4.72328 //w=0.131 //l=4.95 //layer=m1 \
 //thickness=0.36 //x=6.175 //y=4.07 //x2=1.225 //y2=4.07
ends PM_HA\%A

subckt PM_HA\%B ( 1 2 3 4 5 6 7 8 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 \
 38 39 41 57 69 84 85 86 87 88 89 90 91 92 93 94 95 100 102 104 110 111 112 \
 113 114 115 116 118 121 122 129 130 134 135 136 138 141 144 145 146 147 149 \
 150 153 169 174 )
c313 ( 174 0 ) capacitor c=0.051138f //x=15.8 //y=2.085
c314 ( 169 0 ) capacitor c=0.0606568f //x=12.21 //y=4.7
c315 ( 153 0 ) capacitor c=0.0331552f //x=1.88 //y=4.7
c316 ( 150 0 ) capacitor c=0.0279499f //x=1.85 //y=1.915
c317 ( 149 0 ) capacitor c=0.0437302f //x=1.85 //y=2.08
c318 ( 147 0 ) capacitor c=0.0290017f //x=15.8 //y=1.92
c319 ( 146 0 ) capacitor c=0.0250171f //x=15.8 //y=1.565
c320 ( 145 0 ) capacitor c=0.0234316f //x=15.8 //y=1.255
c321 ( 144 0 ) capacitor c=0.0200712f //x=15.8 //y=0.91
c322 ( 141 0 ) capacitor c=0.0488625f //x=15.755 //y=4.865
c323 ( 138 0 ) capacitor c=0.0152946f //x=15.645 //y=1.41
c324 ( 136 0 ) capacitor c=0.0157804f //x=15.645 //y=0.755
c325 ( 135 0 ) capacitor c=0.0129718f //x=15.39 //y=4.79
c326 ( 134 0 ) capacitor c=0.0172687f //x=15.68 //y=4.79
c327 ( 130 0 ) capacitor c=0.0435512f //x=15.27 //y=1.255
c328 ( 129 0 ) capacitor c=0.0200269f //x=15.27 //y=0.91
c329 ( 122 0 ) capacitor c=0.0417768f //x=10.185 //y=1.255
c330 ( 121 0 ) capacitor c=0.0192208f //x=10.185 //y=0.91
c331 ( 118 0 ) capacitor c=0.0124204f //x=10.03 //y=1.41
c332 ( 116 0 ) capacitor c=0.0157803f //x=10.03 //y=0.755
c333 ( 115 0 ) capacitor c=0.0903325f //x=9.655 //y=1.92
c334 ( 114 0 ) capacitor c=0.0194674f //x=9.655 //y=1.565
c335 ( 113 0 ) capacitor c=0.0168481f //x=9.655 //y=1.255
c336 ( 112 0 ) capacitor c=0.0174345f //x=9.655 //y=0.91
c337 ( 111 0 ) capacitor c=0.0429696f //x=2.415 //y=1.25
c338 ( 110 0 ) capacitor c=0.0192208f //x=2.415 //y=0.905
c339 ( 104 0 ) capacitor c=0.0158629f //x=2.26 //y=1.405
c340 ( 102 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c341 ( 100 0 ) capacitor c=0.0300505f //x=2.255 //y=4.79
c342 ( 95 0 ) capacitor c=0.0205163f //x=1.885 //y=1.56
c343 ( 94 0 ) capacitor c=0.0168481f //x=1.885 //y=1.25
c344 ( 93 0 ) capacitor c=0.0174783f //x=1.885 //y=0.905
c345 ( 92 0 ) capacitor c=0.154243f //x=15.755 //y=6.02
c346 ( 91 0 ) capacitor c=0.154218f //x=15.315 //y=6.02
c347 ( 90 0 ) capacitor c=0.110797f //x=12.55 //y=6.02
c348 ( 89 0 ) capacitor c=0.154322f //x=12.11 //y=6.02
c349 ( 88 0 ) capacitor c=0.15358f //x=2.33 //y=6.02
c350 ( 87 0 ) capacitor c=0.110281f //x=1.89 //y=6.02
c351 ( 69 0 ) capacitor c=0.106666f //x=15.91 //y=2.085
c352 ( 57 0 ) capacitor c=0.0306114f //x=9.99 //y=2.085
c353 ( 41 0 ) capacitor c=0.0765209f //x=1.85 //y=2.08
c354 ( 39 0 ) capacitor c=0.00453889f //x=1.85 //y=4.535
c355 ( 32 0 ) capacitor c=0.0151539f //x=12.21 //y=4.44
c356 ( 28 0 ) capacitor c=0.0375706f //x=9.62 //y=3.7
c357 ( 8 0 ) capacitor c=0.00543706f //x=12.325 //y=4.44
c358 ( 7 0 ) capacitor c=0.093123f //x=15.795 //y=4.44
c359 ( 6 0 ) capacitor c=0.0154186f //x=10.105 //y=2.96
c360 ( 5 0 ) capacitor c=0.130205f //x=15.795 //y=2.96
c361 ( 4 0 ) capacitor c=0.0156999f //x=9.735 //y=4.44
c362 ( 3 0 ) capacitor c=0.0540768f //x=12.095 //y=4.44
c363 ( 2 0 ) capacitor c=0.0160493f //x=1.965 //y=3.7
c364 ( 1 0 ) capacitor c=0.186881f //x=9.505 //y=3.7
r365 (  174 176 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.8 //y=2.085 //x2=15.91 //y2=2.085
r366 (  167 169 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=12.11 //y=4.7 //x2=12.21 //y2=4.7
r367 (  155 156 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.79 //x2=1.88 //y2=4.865
r368 (  153 155 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.7 //x2=1.88 //y2=4.79
r369 (  149 150 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r370 (  147 174 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=15.8 //y=1.92 //x2=15.8 //y2=2.085
r371 (  146 173 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.8 //y=1.565 //x2=15.76 //y2=1.41
r372 (  146 147 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=15.8 //y=1.565 //x2=15.8 //y2=1.92
r373 (  145 173 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.8 //y=1.255 //x2=15.76 //y2=1.41
r374 (  144 172 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.8 //y=0.91 //x2=15.76 //y2=0.755
r375 (  144 145 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.8 //y=0.91 //x2=15.8 //y2=1.255
r376 (  141 178 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=15.755 //y=4.865 //x2=15.91 //y2=4.7
r377 (  139 171 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.425 //y=1.41 //x2=15.31 //y2=1.41
r378 (  138 173 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.645 //y=1.41 //x2=15.76 //y2=1.41
r379 (  137 170 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.425 //y=0.755 //x2=15.31 //y2=0.755
r380 (  136 172 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.645 //y=0.755 //x2=15.76 //y2=0.755
r381 (  136 137 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.645 //y=0.755 //x2=15.425 //y2=0.755
r382 (  134 141 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.68 //y=4.79 //x2=15.755 //y2=4.865
r383 (  134 135 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=15.68 //y=4.79 //x2=15.39 //y2=4.79
r384 (  131 135 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.315 //y=4.865 //x2=15.39 //y2=4.79
r385 (  130 171 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.27 //y=1.255 //x2=15.31 //y2=1.41
r386 (  129 170 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.27 //y=0.91 //x2=15.31 //y2=0.755
r387 (  129 130 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.27 //y=0.91 //x2=15.27 //y2=1.255
r388 (  126 169 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=12.55 //y=4.865 //x2=12.21 //y2=4.7
r389 (  123 167 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=12.11 //y=4.865 //x2=12.11 //y2=4.7
r390 (  122 166 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.185 //y=1.255 //x2=10.145 //y2=1.41
r391 (  121 165 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.185 //y=0.91 //x2=10.145 //y2=0.755
r392 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.185 //y=0.91 //x2=10.185 //y2=1.255
r393 (  119 162 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.81 //y=1.41 //x2=9.695 //y2=1.41
r394 (  118 166 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.03 //y=1.41 //x2=10.145 //y2=1.41
r395 (  117 161 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.81 //y=0.755 //x2=9.695 //y2=0.755
r396 (  116 165 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.03 //y=0.755 //x2=10.145 //y2=0.755
r397 (  116 117 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.03 //y=0.755 //x2=9.81 //y2=0.755
r398 (  115 164 ) resistor r=67.2792 //w=0.24 //l=0.438891 //layer=ply \
 //thickness=0.18 //x=9.655 //y=1.92 //x2=9.99 //y2=2.16
r399 (  114 162 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.655 //y=1.565 //x2=9.695 //y2=1.41
r400 (  114 115 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=9.655 //y=1.565 //x2=9.655 //y2=1.92
r401 (  113 162 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.655 //y=1.255 //x2=9.695 //y2=1.41
r402 (  112 161 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.655 //y=0.91 //x2=9.695 //y2=0.755
r403 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.655 //y=0.91 //x2=9.655 //y2=1.255
r404 (  111 160 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r405 (  110 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r406 (  110 111 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r407 (  105 158 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r408 (  104 160 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r409 (  103 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r410 (  102 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r411 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r412 (  101 155 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.015 //y=4.79 //x2=1.88 //y2=4.79
r413 (  100 107 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.33 //y2=4.865
r414 (  100 101 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.015 //y2=4.79
r415 (  95 158 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r416 (  95 150 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r417 (  94 158 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r418 (  93 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r419 (  93 94 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r420 (  92 141 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.755 //y=6.02 //x2=15.755 //y2=4.865
r421 (  91 131 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.315 //y=6.02 //x2=15.315 //y2=4.865
r422 (  90 126 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.55 //y=6.02 //x2=12.55 //y2=4.865
r423 (  89 123 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.11 //y=6.02 //x2=12.11 //y2=4.865
r424 (  88 107 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.02 //x2=2.33 //y2=4.865
r425 (  87 156 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.02 //x2=1.89 //y2=4.865
r426 (  86 138 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.535 //y=1.41 //x2=15.645 //y2=1.41
r427 (  86 139 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.535 //y=1.41 //x2=15.425 //y2=1.41
r428 (  85 118 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.92 //y=1.41 //x2=10.03 //y2=1.41
r429 (  85 119 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.92 //y=1.41 //x2=9.81 //y2=1.41
r430 (  84 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r431 (  84 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r432 (  83 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.88 //y=4.7 //x2=1.88 //y2=4.7
r433 (  80 178 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.91 //y=4.7 //x2=15.91 //y2=4.7
r434 (  69 176 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.91 //y=2.085 //x2=15.91 //y2=2.085
r435 (  66 169 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.21 //y=4.7 //x2=12.21 //y2=4.7
r436 (  57 164 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.99 //y=2.085 //x2=9.99 //y2=2.085
r437 (  41 149 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r438 (  39 83 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.865 //y2=4.7
r439 (  38 80 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=15.91 //y=4.44 //x2=15.91 //y2=4.7
r440 (  37 38 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.91 //y=4.07 //x2=15.91 //y2=4.44
r441 (  36 37 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.91 //y=3.7 //x2=15.91 //y2=4.07
r442 (  35 36 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.91 //y=3.33 //x2=15.91 //y2=3.7
r443 (  34 35 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.91 //y=2.96 //x2=15.91 //y2=3.33
r444 (  33 34 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.91 //y=2.59 //x2=15.91 //y2=2.96
r445 (  33 69 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=15.91 //y=2.59 //x2=15.91 //y2=2.085
r446 (  32 66 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=12.21 //y=4.44 //x2=12.21 //y2=4.7
r447 (  31 57 ) resistor r=59.893 //w=0.187 //l=0.875 //layer=li \
 //thickness=0.1 //x=9.99 //y=2.96 //x2=9.99 //y2=2.085
r448 (  29 30 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=9.62 //y=4.07 //x2=9.62 //y2=4.44
r449 (  28 29 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=9.62 //y=3.7 //x2=9.62 //y2=4.07
r450 (  27 39 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.44 //x2=1.85 //y2=4.535
r451 (  26 27 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=1.85 //y=3.7 //x2=1.85 //y2=4.44
r452 (  25 26 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.85 //y=3.33 //x2=1.85 //y2=3.7
r453 (  24 25 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.96 //x2=1.85 //y2=3.33
r454 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.59 //x2=1.85 //y2=2.96
r455 (  23 41 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.59 //x2=1.85 //y2=2.08
r456 (  22 38 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.91 //y=4.44 //x2=15.91 //y2=4.44
r457 (  20 34 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.91 //y=2.96 //x2=15.91 //y2=2.96
r458 (  18 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.21 //y=4.44 //x2=12.21 //y2=4.44
r459 (  16 31 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.99 //y=2.96 //x2=9.99 //y2=2.96
r460 (  14 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.62 //y=3.7 //x2=9.62 //y2=3.7
r461 (  12 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.62 //y=4.44 //x2=9.62 //y2=4.44
r462 (  10 26 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.85 //y=3.7 //x2=1.85 //y2=3.7
r463 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.325 //y=4.44 //x2=12.21 //y2=4.44
r464 (  7 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=4.44 //x2=15.91 //y2=4.44
r465 (  7 8 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=4.44 //x2=12.325 //y2=4.44
r466 (  6 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.105 //y=2.96 //x2=9.99 //y2=2.96
r467 (  5 20 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=2.96 //x2=15.91 //y2=2.96
r468 (  5 6 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=2.96 //x2=10.105 //y2=2.96
r469 (  4 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.735 //y=4.44 //x2=9.62 //y2=4.44
r470 (  3 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.095 //y=4.44 //x2=12.21 //y2=4.44
r471 (  3 4 ) resistor r=2.25191 //w=0.131 //l=2.36 //layer=m1 \
 //thickness=0.36 //x=12.095 //y=4.44 //x2=9.735 //y2=4.44
r472 (  2 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.965 //y=3.7 //x2=1.85 //y2=3.7
r473 (  1 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=3.7 //x2=9.62 //y2=3.7
r474 (  1 2 ) resistor r=7.19466 //w=0.131 //l=7.54 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=3.7 //x2=1.965 //y2=3.7
ends PM_HA\%B

subckt PM_HA\%noxref_6 ( 1 2 17 18 19 20 24 26 33 34 35 36 37 38 39 43 45 51 \
 52 60 62 64 )
c175 ( 64 0 ) capacitor c=0.0288629f //x=6.52 //y=5.02
c176 ( 62 0 ) capacitor c=0.0173218f //x=6.475 //y=0.91
c177 ( 60 0 ) capacitor c=0.058481f //x=13.32 //y=4.7
c178 ( 52 0 ) capacitor c=0.0417768f //x=13.515 //y=1.255
c179 ( 51 0 ) capacitor c=0.0192208f //x=13.515 //y=0.91
c180 ( 45 0 ) capacitor c=0.0124204f //x=13.36 //y=1.41
c181 ( 43 0 ) capacitor c=0.0157803f //x=13.36 //y=0.755
c182 ( 39 0 ) capacitor c=0.0903287f //x=12.985 //y=1.92
c183 ( 38 0 ) capacitor c=0.0194674f //x=12.985 //y=1.565
c184 ( 37 0 ) capacitor c=0.0168481f //x=12.985 //y=1.255
c185 ( 36 0 ) capacitor c=0.0174345f //x=12.985 //y=0.91
c186 ( 35 0 ) capacitor c=0.153255f //x=13.43 //y=6.02
c187 ( 34 0 ) capacitor c=0.110227f //x=12.99 //y=6.02
c188 ( 26 0 ) capacitor c=0.0737449f //x=13.32 //y=2.085
c189 ( 24 0 ) capacitor c=0.0836439f //x=7.03 //y=2.59
c190 ( 20 0 ) capacitor c=0.00417404f //x=6.75 //y=4.58
c191 ( 19 0 ) capacitor c=0.0118459f //x=6.945 //y=4.58
c192 ( 18 0 ) capacitor c=0.00612032f //x=6.745 //y=2.08
c193 ( 17 0 ) capacitor c=0.0133843f //x=6.945 //y=2.08
c194 ( 2 0 ) capacitor c=0.0160697f //x=7.145 //y=2.59
c195 ( 1 0 ) capacitor c=0.16891f //x=13.205 //y=2.59
r196 (  60 61 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.32 //y=4.7 //x2=13.43 //y2=4.7
r197 (  52 58 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.515 //y=1.255 //x2=13.475 //y2=1.41
r198 (  51 57 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.515 //y=0.91 //x2=13.475 //y2=0.755
r199 (  51 52 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.515 //y=0.91 //x2=13.515 //y2=1.255
r200 (  48 61 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=13.43 //y=4.865 //x2=13.43 //y2=4.7
r201 (  46 54 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.14 //y=1.41 //x2=13.025 //y2=1.41
r202 (  45 58 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.36 //y=1.41 //x2=13.475 //y2=1.41
r203 (  44 53 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.14 //y=0.755 //x2=13.025 //y2=0.755
r204 (  43 57 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.36 //y=0.755 //x2=13.475 //y2=0.755
r205 (  43 44 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=13.36 //y=0.755 //x2=13.14 //y2=0.755
r206 (  40 60 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=12.99 //y=4.865 //x2=13.32 //y2=4.7
r207 (  39 56 ) resistor r=67.2792 //w=0.24 //l=0.438891 //layer=ply \
 //thickness=0.18 //x=12.985 //y=1.92 //x2=13.32 //y2=2.16
r208 (  38 54 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.985 //y=1.565 //x2=13.025 //y2=1.41
r209 (  38 39 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=12.985 //y=1.565 //x2=12.985 //y2=1.92
r210 (  37 54 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.985 //y=1.255 //x2=13.025 //y2=1.41
r211 (  36 53 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.985 //y=0.91 //x2=13.025 //y2=0.755
r212 (  36 37 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.985 //y=0.91 //x2=12.985 //y2=1.255
r213 (  35 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.43 //y=6.02 //x2=13.43 //y2=4.865
r214 (  34 40 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.99 //y=6.02 //x2=12.99 //y2=4.865
r215 (  33 45 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.25 //y=1.41 //x2=13.36 //y2=1.41
r216 (  33 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.25 //y=1.41 //x2=13.14 //y2=1.41
r217 (  31 60 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=13.32 //y=4.7 //x2=13.32 //y2=4.7
r218 (  29 31 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=13.32 //y=2.59 //x2=13.32 //y2=4.7
r219 (  26 56 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=13.32 //y=2.085 //x2=13.32 //y2=2.085
r220 (  26 29 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=13.32 //y=2.085 //x2=13.32 //y2=2.59
r221 (  22 24 ) resistor r=130.396 //w=0.187 //l=1.905 //layer=li \
 //thickness=0.1 //x=7.03 //y=4.495 //x2=7.03 //y2=2.59
r222 (  21 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.165 //x2=7.03 //y2=2.59
r223 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.945 //y=4.58 //x2=7.03 //y2=4.495
r224 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=6.945 //y=4.58 //x2=6.75 //y2=4.58
r225 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.945 //y=2.08 //x2=7.03 //y2=2.165
r226 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=6.945 //y=2.08 //x2=6.745 //y2=2.08
r227 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.665 //y=4.665 //x2=6.75 //y2=4.58
r228 (  11 64 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=6.665 //y=4.665 //x2=6.665 //y2=5.725
r229 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.66 //y=1.995 //x2=6.745 //y2=2.08
r230 (  7 62 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=6.66 //y=1.995 //x2=6.66 //y2=1.005
r231 (  6 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=13.32 //y=2.59 //x2=13.32 //y2=2.59
r232 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.03 //y=2.59 //x2=7.03 //y2=2.59
r233 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.145 //y=2.59 //x2=7.03 //y2=2.59
r234 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.205 //y=2.59 //x2=13.32 //y2=2.59
r235 (  1 2 ) resistor r=5.78244 //w=0.131 //l=6.06 //layer=m1 \
 //thickness=0.36 //x=13.205 //y=2.59 //x2=7.145 //y2=2.59
ends PM_HA\%noxref_6

subckt PM_HA\%SUM ( 1 2 7 8 9 10 11 12 13 14 25 26 27 28 46 47 48 49 57 58 61 \
 62 )
c152 ( 62 0 ) capacitor c=0.0159588f //x=13.065 //y=5.02
c153 ( 61 0 ) capacitor c=0.0159588f //x=9.735 //y=5.02
c154 ( 58 0 ) capacitor c=0.00827922f //x=13.06 //y=0.91
c155 ( 57 0 ) capacitor c=0.00846882f //x=9.73 //y=0.91
c156 ( 49 0 ) capacitor c=0.00178322f //x=13.335 //y=1.655
c157 ( 48 0 ) capacitor c=0.0112025f //x=13.605 //y=1.655
c158 ( 47 0 ) capacitor c=0.00235465f //x=13.295 //y=5.205
c159 ( 46 0 ) capacitor c=0.0121398f //x=13.605 //y=5.205
c160 ( 28 0 ) capacitor c=0.00178606f //x=10.005 //y=1.655
c161 ( 27 0 ) capacitor c=0.0109582f //x=10.275 //y=1.655
c162 ( 26 0 ) capacitor c=0.00235465f //x=9.965 //y=5.205
c163 ( 25 0 ) capacitor c=0.0119514f //x=10.275 //y=5.205
c164 ( 11 0 ) capacitor c=0.0892717f //x=13.69 //y=2.22
c165 ( 7 0 ) capacitor c=0.101908f //x=10.36 //y=2.22
c166 ( 2 0 ) capacitor c=0.0058186f //x=10.475 //y=3.7
c167 ( 1 0 ) capacitor c=0.0664888f //x=13.575 //y=3.7
r168 (  48 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.655 //x2=13.69 //y2=1.74
r169 (  48 49 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.655 //x2=13.335 //y2=1.655
r170 (  46 51 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.205 //x2=13.69 //y2=5.12
r171 (  46 47 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.205 //x2=13.295 //y2=5.205
r172 (  42 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.25 //y=1.57 //x2=13.335 //y2=1.655
r173 (  42 58 ) resistor r=38.6738 //w=0.187 //l=0.565 //layer=li \
 //thickness=0.1 //x=13.25 //y=1.57 //x2=13.25 //y2=1.005
r174 (  36 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.21 //y=5.29 //x2=13.295 //y2=5.205
r175 (  36 62 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=13.21 //y=5.29 //x2=13.21 //y2=5.715
r176 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.275 //y=1.655 //x2=10.36 //y2=1.74
r177 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=10.275 //y=1.655 //x2=10.005 //y2=1.655
r178 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.275 //y=5.205 //x2=10.36 //y2=5.12
r179 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=10.275 //y=5.205 //x2=9.965 //y2=5.205
r180 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.92 //y=1.57 //x2=10.005 //y2=1.655
r181 (  21 57 ) resistor r=38.6738 //w=0.187 //l=0.565 //layer=li \
 //thickness=0.1 //x=9.92 //y=1.57 //x2=9.92 //y2=1.005
r182 (  15 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.88 //y=5.29 //x2=9.965 //y2=5.205
r183 (  15 61 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=9.88 //y=5.29 //x2=9.88 //y2=5.715
r184 (  14 51 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=13.69 //y=4.81 //x2=13.69 //y2=5.12
r185 (  13 14 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=13.69 //y=3.7 //x2=13.69 //y2=4.81
r186 (  12 13 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=13.69 //y=2.59 //x2=13.69 //y2=3.7
r187 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=13.69 //y=2.22 //x2=13.69 //y2=2.59
r188 (  11 50 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li \
 //thickness=0.1 //x=13.69 //y=2.22 //x2=13.69 //y2=1.74
r189 (  10 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=10.36 //y=4.81 //x2=10.36 //y2=5.12
r190 (  9 10 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=10.36 //y=3.7 //x2=10.36 //y2=4.81
r191 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=10.36 //y=3.33 //x2=10.36 //y2=3.7
r192 (  7 8 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li //thickness=0.1 \
 //x=10.36 //y=2.22 //x2=10.36 //y2=3.33
r193 (  7 29 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.22 //x2=10.36 //y2=1.74
r194 (  6 13 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=13.69 //y=3.7 //x2=13.69 //y2=3.7
r195 (  4 9 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=3.7 //x2=10.36 //y2=3.7
r196 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.475 //y=3.7 //x2=10.36 //y2=3.7
r197 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.575 //y=3.7 //x2=13.69 //y2=3.7
r198 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=13.575 //y=3.7 //x2=10.475 //y2=3.7
ends PM_HA\%SUM

subckt PM_HA\%noxref_8 ( 1 2 3 4 14 20 28 31 32 33 34 45 46 47 54 55 56 57 58 \
 60 63 64 66 74 76 )
c164 ( 76 0 ) capacitor c=0.028734f //x=15.39 //y=5.02
c165 ( 74 0 ) capacitor c=0.0173218f //x=15.345 //y=0.91
c166 ( 66 0 ) capacitor c=0.0576608f //x=9.99 //y=4.7
c167 ( 64 0 ) capacitor c=0.0318948f //x=12.545 //y=1.215
c168 ( 63 0 ) capacitor c=0.0187407f //x=12.545 //y=0.87
c169 ( 60 0 ) capacitor c=0.0141798f //x=12.39 //y=1.37
c170 ( 58 0 ) capacitor c=0.0149852f //x=12.39 //y=0.715
c171 ( 57 0 ) capacitor c=0.0836807f //x=12.015 //y=1.92
c172 ( 56 0 ) capacitor c=0.0229722f //x=12.015 //y=1.525
c173 ( 55 0 ) capacitor c=0.0234352f //x=12.015 //y=1.215
c174 ( 54 0 ) capacitor c=0.0199366f //x=12.015 //y=0.87
c175 ( 47 0 ) capacitor c=0.153255f //x=10.1 //y=6.02
c176 ( 46 0 ) capacitor c=0.110227f //x=9.66 //y=6.02
c177 ( 34 0 ) capacitor c=0.00670488f //x=15.255 //y=4.58
c178 ( 33 0 ) capacitor c=0.0137356f //x=15.45 //y=4.58
c179 ( 32 0 ) capacitor c=0.00580686f //x=15.255 //y=2.08
c180 ( 31 0 ) capacitor c=0.0128831f //x=15.455 //y=2.08
c181 ( 28 0 ) capacitor c=0.0775792f //x=15.17 //y=3.33
c182 ( 20 0 ) capacitor c=0.0551449f //x=12.21 //y=2.085
c183 ( 14 0 ) capacitor c=0.016943f //x=9.99 //y=4.07
c184 ( 4 0 ) capacitor c=0.0126928f //x=12.325 //y=3.33
c185 ( 3 0 ) capacitor c=0.0544915f //x=15.055 //y=3.33
c186 ( 2 0 ) capacitor c=0.00882264f //x=10.105 //y=4.07
c187 ( 1 0 ) capacitor c=0.0848617f //x=15.055 //y=4.07
r188 (  66 67 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.99 //y=4.7 //x2=10.1 //y2=4.7
r189 (  64 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.545 //y=1.215 //x2=12.505 //y2=1.37
r190 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.545 //y=0.87 //x2=12.505 //y2=0.715
r191 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.545 //y=0.87 //x2=12.545 //y2=1.215
r192 (  61 71 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.17 //y=1.37 //x2=12.055 //y2=1.37
r193 (  60 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.39 //y=1.37 //x2=12.505 //y2=1.37
r194 (  59 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.17 //y=0.715 //x2=12.055 //y2=0.715
r195 (  58 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.39 //y=0.715 //x2=12.505 //y2=0.715
r196 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=12.39 //y=0.715 //x2=12.17 //y2=0.715
r197 (  57 69 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=12.015 //y=1.92 //x2=12.21 //y2=2.085
r198 (  56 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.015 //y=1.525 //x2=12.055 //y2=1.37
r199 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=12.015 //y=1.525 //x2=12.015 //y2=1.92
r200 (  55 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.015 //y=1.215 //x2=12.055 //y2=1.37
r201 (  54 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.015 //y=0.87 //x2=12.055 //y2=0.715
r202 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.015 //y=0.87 //x2=12.015 //y2=1.215
r203 (  51 67 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=10.1 //y=4.865 //x2=10.1 //y2=4.7
r204 (  48 66 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=9.66 //y=4.865 //x2=9.99 //y2=4.7
r205 (  47 51 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.1 //y=6.02 //x2=10.1 //y2=4.865
r206 (  46 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.66 //y=6.02 //x2=9.66 //y2=4.865
r207 (  45 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.28 //y=1.37 //x2=12.39 //y2=1.37
r208 (  45 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.28 //y=1.37 //x2=12.17 //y2=1.37
r209 (  41 74 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=15.54 //y=1.995 //x2=15.54 //y2=1.005
r210 (  35 76 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=15.535 //y=4.665 //x2=15.535 //y2=5.725
r211 (  33 35 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.45 //y=4.58 //x2=15.535 //y2=4.665
r212 (  33 34 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=15.45 //y=4.58 //x2=15.255 //y2=4.58
r213 (  31 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.455 //y=2.08 //x2=15.54 //y2=1.995
r214 (  31 32 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=15.455 //y=2.08 //x2=15.255 //y2=2.08
r215 (  28 30 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=15.17 //y=3.33 //x2=15.17 //y2=4.07
r216 (  26 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.17 //y=4.495 //x2=15.255 //y2=4.58
r217 (  26 30 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=15.17 //y=4.495 //x2=15.17 //y2=4.07
r218 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.17 //y=2.165 //x2=15.255 //y2=2.08
r219 (  25 28 ) resistor r=79.7433 //w=0.187 //l=1.165 //layer=li \
 //thickness=0.1 //x=15.17 //y=2.165 //x2=15.17 //y2=3.33
r220 (  20 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.21 //y=2.085 //x2=12.21 //y2=2.085
r221 (  20 23 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=12.21 //y=2.085 //x2=12.21 //y2=3.33
r222 (  17 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.99 //y=4.7 //x2=9.99 //y2=4.7
r223 (  14 17 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=9.99 //y=4.07 //x2=9.99 //y2=4.7
r224 (  12 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.17 //y=4.07 //x2=15.17 //y2=4.07
r225 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.17 //y=3.33 //x2=15.17 //y2=3.33
r226 (  8 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.21 //y=3.33 //x2=12.21 //y2=3.33
r227 (  6 14 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.99 //y=4.07 //x2=9.99 //y2=4.07
r228 (  4 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.325 //y=3.33 //x2=12.21 //y2=3.33
r229 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.055 //y=3.33 //x2=15.17 //y2=3.33
r230 (  3 4 ) resistor r=2.60496 //w=0.131 //l=2.73 //layer=m1 \
 //thickness=0.36 //x=15.055 //y=3.33 //x2=12.325 //y2=3.33
r231 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.105 //y=4.07 //x2=9.99 //y2=4.07
r232 (  1 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.055 //y=4.07 //x2=15.17 //y2=4.07
r233 (  1 2 ) resistor r=4.72328 //w=0.131 //l=4.95 //layer=m1 \
 //thickness=0.36 //x=15.055 //y=4.07 //x2=10.105 //y2=4.07
ends PM_HA\%noxref_8

subckt PM_HA\%noxref_9 ( 1 5 9 10 13 17 29 )
c55 ( 29 0 ) capacitor c=0.0633899f //x=0.56 //y=0.365
c56 ( 17 0 ) capacitor c=0.00722223f //x=2.635 //y=0.615
c57 ( 13 0 ) capacitor c=0.0150745f //x=2.55 //y=0.53
c58 ( 10 0 ) capacitor c=0.00705906f //x=1.665 //y=1.495
c59 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c60 ( 5 0 ) capacitor c=0.0218843f //x=1.58 //y=1.58
c61 ( 1 0 ) capacitor c=0.0113547f //x=0.695 //y=1.495
r62 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r63 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r64 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r65 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=2.15 //y2=0.53
r66 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r67 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.15 //y2=0.53
r68 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r69 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r70 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r71 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r72 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r73 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r74 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r75 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r76 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r77 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_HA\%noxref_9

subckt PM_HA\%COUT ( 1 2 3 4 5 16 17 18 19 27 29 )
c55 ( 29 0 ) capacitor c=0.028734f //x=4.3 //y=5.02
c56 ( 27 0 ) capacitor c=0.0173218f //x=4.255 //y=0.91
c57 ( 19 0 ) capacitor c=0.00417404f //x=4.53 //y=4.58
c58 ( 18 0 ) capacitor c=0.0118896f //x=4.725 //y=4.58
c59 ( 17 0 ) capacitor c=0.00612032f //x=4.525 //y=2.08
c60 ( 16 0 ) capacitor c=0.0138937f //x=4.725 //y=2.08
c61 ( 1 0 ) capacitor c=0.0826122f //x=4.81 //y=2.22
r62 (  18 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=4.58 //x2=4.81 //y2=4.495
r63 (  18 19 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=4.725 //y=4.58 //x2=4.53 //y2=4.58
r64 (  16 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=2.08 //x2=4.81 //y2=2.165
r65 (  16 17 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=4.725 //y=2.08 //x2=4.525 //y2=2.08
r66 (  10 19 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.445 //y=4.665 //x2=4.53 //y2=4.58
r67 (  10 29 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=4.445 //y=4.665 //x2=4.445 //y2=5.725
r68 (  6 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.44 //y=1.995 //x2=4.525 //y2=2.08
r69 (  6 27 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=4.44 //y=1.995 //x2=4.44 //y2=1.005
r70 (  5 21 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=4.81 //y=4.44 //x2=4.81 //y2=4.495
r71 (  4 5 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li //thickness=0.1 \
 //x=4.81 //y=3.33 //x2=4.81 //y2=4.44
r72 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.81 //y=2.96 //x2=4.81 //y2=3.33
r73 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.81 //y=2.59 //x2=4.81 //y2=2.96
r74 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.81 //y=2.22 //x2=4.81 //y2=2.59
r75 (  1 20 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=4.81 //y=2.22 //x2=4.81 //y2=2.165
ends PM_HA\%COUT

subckt PM_HA\%noxref_11 ( 7 8 15 16 23 24 25 )
c44 ( 25 0 ) capacitor c=0.0305804f //x=10.175 //y=5.02
c45 ( 24 0 ) capacitor c=0.0185379f //x=9.295 //y=5.02
c46 ( 23 0 ) capacitor c=0.0384176f //x=8.425 //y=5.02
c47 ( 16 0 ) capacitor c=0.00194711f //x=9.525 //y=6.905
c48 ( 15 0 ) capacitor c=0.0132608f //x=10.235 //y=6.905
c49 ( 8 0 ) capacitor c=0.00644339f //x=8.645 //y=5.205
c50 ( 7 0 ) capacitor c=0.0195248f //x=9.355 //y=5.205
r51 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.32 //y=6.82 //x2=10.32 //y2=6.735
r52 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.235 //y=6.905 //x2=10.32 //y2=6.82
r53 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.235 //y=6.905 //x2=9.525 //y2=6.905
r54 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.44 //y=6.82 //x2=9.525 //y2=6.905
r55 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=9.44 //y=6.82 //x2=9.44 //y2=6.395
r56 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=9.44 //y=5.29 //x2=9.44 //y2=5.715
r57 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.355 //y=5.205 //x2=9.44 //y2=5.29
r58 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=9.355 //y=5.205 //x2=8.645 //y2=5.205
r59 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.56 //y=5.29 //x2=8.645 //y2=5.205
r60 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=8.56 //y=5.29 //x2=8.56 //y2=5.715
ends PM_HA\%noxref_11

subckt PM_HA\%noxref_12 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.0632228f //x=8.33 //y=0.37
c54 ( 17 0 ) capacitor c=0.00723243f //x=10.405 //y=0.62
c55 ( 13 0 ) capacitor c=0.0150659f //x=10.32 //y=0.535
c56 ( 10 0 ) capacitor c=0.00656687f //x=9.435 //y=1.5
c57 ( 9 0 ) capacitor c=0.00677124f //x=9.435 //y=0.62
c58 ( 5 0 ) capacitor c=0.0181169f //x=9.35 //y=1.585
c59 ( 1 0 ) capacitor c=0.0076549f //x=8.465 //y=1.5
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=10.405 //y=0.62 //x2=10.405 //y2=0.495
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=10.405 //y=0.62 //x2=10.405 //y2=0.885
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.52 //y=0.535 //x2=9.435 //y2=0.495
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.52 //y=0.535 //x2=9.92 //y2=0.535
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.32 //y=0.535 //x2=10.405 //y2=0.495
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.32 //y=0.535 //x2=9.92 //y2=0.535
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.435 //y=1.5 //x2=9.435 //y2=1.625
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.435 //y=1.5 //x2=9.435 //y2=0.885
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.435 //y=0.62 //x2=9.435 //y2=0.495
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=9.435 //y=0.62 //x2=9.435 //y2=0.885
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.55 //y=1.585 //x2=8.465 //y2=1.625
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.55 //y=1.585 //x2=8.95 //y2=1.585
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.35 //y=1.585 //x2=9.435 //y2=1.625
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.35 //y=1.585 //x2=8.95 //y2=1.585
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.465 //y=1.5 //x2=8.465 //y2=1.625
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.465 //y=1.5 //x2=8.465 //y2=0.885
ends PM_HA\%noxref_12

subckt PM_HA\%noxref_13 ( 7 8 15 16 23 24 25 )
c43 ( 25 0 ) capacitor c=0.0305804f //x=13.505 //y=5.02
c44 ( 24 0 ) capacitor c=0.0185379f //x=12.625 //y=5.02
c45 ( 23 0 ) capacitor c=0.0384176f //x=11.755 //y=5.02
c46 ( 16 0 ) capacitor c=0.00194711f //x=12.855 //y=6.905
c47 ( 15 0 ) capacitor c=0.0133643f //x=13.565 //y=6.905
c48 ( 8 0 ) capacitor c=0.00598116f //x=11.975 //y=5.205
c49 ( 7 0 ) capacitor c=0.0182615f //x=12.685 //y=5.205
r50 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.65 //y=6.82 //x2=13.65 //y2=6.735
r51 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.565 //y=6.905 //x2=13.65 //y2=6.82
r52 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=13.565 //y=6.905 //x2=12.855 //y2=6.905
r53 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.77 //y=6.82 //x2=12.855 //y2=6.905
r54 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=12.77 //y=6.82 //x2=12.77 //y2=6.395
r55 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=12.77 //y=5.29 //x2=12.77 //y2=5.715
r56 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.685 //y=5.205 //x2=12.77 //y2=5.29
r57 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=12.685 //y=5.205 //x2=11.975 //y2=5.205
r58 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.89 //y=5.29 //x2=11.975 //y2=5.205
r59 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=11.89 //y=5.29 //x2=11.89 //y2=5.715
ends PM_HA\%noxref_13

subckt PM_HA\%noxref_14 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.063541f //x=11.66 //y=0.37
c54 ( 17 0 ) capacitor c=0.00723243f //x=13.735 //y=0.62
c55 ( 13 0 ) capacitor c=0.0153645f //x=13.65 //y=0.535
c56 ( 10 0 ) capacitor c=0.00656687f //x=12.765 //y=1.5
c57 ( 9 0 ) capacitor c=0.00677124f //x=12.765 //y=0.62
c58 ( 5 0 ) capacitor c=0.0181169f //x=12.68 //y=1.585
c59 ( 1 0 ) capacitor c=0.0076549f //x=11.795 //y=1.5
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=13.735 //y=0.62 //x2=13.735 //y2=0.495
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=13.735 //y=0.62 //x2=13.735 //y2=0.885
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.85 //y=0.535 //x2=12.765 //y2=0.495
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.85 //y=0.535 //x2=13.25 //y2=0.535
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.65 //y=0.535 //x2=13.735 //y2=0.495
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.65 //y=0.535 //x2=13.25 //y2=0.535
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=12.765 //y=1.5 //x2=12.765 //y2=1.625
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=12.765 //y=1.5 //x2=12.765 //y2=0.885
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=12.765 //y=0.62 //x2=12.765 //y2=0.495
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=12.765 //y=0.62 //x2=12.765 //y2=0.885
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.88 //y=1.585 //x2=11.795 //y2=1.625
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.88 //y=1.585 //x2=12.28 //y2=1.585
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.68 //y=1.585 //x2=12.765 //y2=1.625
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.68 //y=1.585 //x2=12.28 //y2=1.585
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.795 //y=1.5 //x2=11.795 //y2=1.625
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=11.795 //y=1.5 //x2=11.795 //y2=0.885
ends PM_HA\%noxref_14

