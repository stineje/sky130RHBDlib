magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 157 187 203
rect 1 21 781 157
rect 84 -17 118 21
<< scnmos >>
rect 79 47 109 177
rect 188 47 218 131
rect 284 47 314 131
rect 409 47 439 131
rect 505 47 535 131
rect 673 47 703 131
<< scpmoshvt >>
rect 79 297 109 497
rect 188 374 218 458
rect 291 374 321 458
rect 505 374 535 458
rect 577 374 607 458
rect 673 374 703 458
<< ndiff >>
rect 27 112 79 177
rect 27 78 35 112
rect 69 78 79 112
rect 27 47 79 78
rect 109 131 161 177
rect 109 93 188 131
rect 109 59 119 93
rect 153 59 188 93
rect 109 47 188 59
rect 218 47 284 131
rect 314 108 409 131
rect 314 74 326 108
rect 360 74 409 108
rect 314 47 409 74
rect 439 47 505 131
rect 535 108 673 131
rect 535 74 561 108
rect 595 74 629 108
rect 663 74 673 108
rect 535 47 673 74
rect 703 108 755 131
rect 703 74 713 108
rect 747 74 755 108
rect 703 47 755 74
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 161 497
rect 109 451 119 485
rect 153 458 161 485
rect 153 451 188 458
rect 109 417 188 451
rect 109 383 119 417
rect 153 383 188 417
rect 109 374 188 383
rect 218 374 291 458
rect 321 425 505 458
rect 321 391 355 425
rect 389 391 430 425
rect 464 391 505 425
rect 321 374 505 391
rect 535 374 577 458
rect 607 425 673 458
rect 607 391 627 425
rect 661 391 673 425
rect 607 374 673 391
rect 703 425 759 458
rect 703 391 713 425
rect 747 391 759 425
rect 703 374 759 391
rect 109 349 161 374
rect 109 315 119 349
rect 153 315 161 349
rect 109 297 161 315
<< ndiffc >>
rect 35 78 69 112
rect 119 59 153 93
rect 326 74 360 108
rect 561 74 595 108
rect 629 74 663 108
rect 713 74 747 108
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 355 391 389 425
rect 430 391 464 425
rect 627 391 661 425
rect 713 391 747 425
rect 119 315 153 349
<< poly >>
rect 79 497 109 523
rect 188 458 218 484
rect 291 458 321 484
rect 505 458 535 484
rect 577 458 607 484
rect 673 458 703 484
rect 79 265 109 297
rect 188 265 218 374
rect 291 359 321 374
rect 291 329 439 359
rect 505 342 535 374
rect 76 249 130 265
rect 76 215 86 249
rect 120 215 130 249
rect 76 199 130 215
rect 172 249 226 265
rect 172 215 182 249
rect 216 215 226 249
rect 409 229 439 329
rect 481 326 535 342
rect 481 292 491 326
rect 525 292 535 326
rect 481 276 535 292
rect 172 199 226 215
rect 284 213 367 229
rect 79 177 109 199
rect 188 131 218 199
rect 284 179 323 213
rect 357 179 367 213
rect 284 163 367 179
rect 409 213 463 229
rect 577 223 607 374
rect 673 342 703 374
rect 649 326 703 342
rect 649 292 659 326
rect 693 292 703 326
rect 649 276 703 292
rect 409 179 419 213
rect 453 179 463 213
rect 565 213 631 223
rect 565 199 581 213
rect 409 163 463 179
rect 505 179 581 199
rect 615 179 631 213
rect 505 169 631 179
rect 284 131 314 163
rect 409 131 439 163
rect 505 131 535 169
rect 673 131 703 276
rect 79 21 109 47
rect 188 21 218 47
rect 284 21 314 47
rect 409 21 439 47
rect 505 21 535 47
rect 673 21 703 47
<< polycont >>
rect 86 215 120 249
rect 182 215 216 249
rect 491 292 525 326
rect 323 179 357 213
rect 659 292 693 326
rect 419 179 453 213
rect 581 179 615 213
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 485 85 493
rect 18 451 35 485
rect 69 451 85 485
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 18 315 35 349
rect 69 315 85 349
rect 18 299 85 315
rect 119 485 153 527
rect 119 417 153 451
rect 119 349 153 383
rect 119 299 153 315
rect 187 459 593 493
rect 18 165 52 299
rect 187 265 221 459
rect 86 249 137 265
rect 120 215 137 249
rect 86 199 137 215
rect 182 249 221 265
rect 216 215 221 249
rect 182 199 221 215
rect 255 391 355 425
rect 389 391 430 425
rect 464 391 480 425
rect 103 165 137 199
rect 255 165 289 391
rect 18 112 69 165
rect 103 131 289 165
rect 323 326 525 357
rect 323 323 491 326
rect 323 213 357 323
rect 487 292 491 323
rect 323 163 357 179
rect 398 213 453 283
rect 398 179 419 213
rect 18 78 35 112
rect 254 124 289 131
rect 254 108 360 124
rect 18 51 69 78
rect 103 93 169 97
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 254 74 326 108
rect 254 51 360 74
rect 398 51 453 179
rect 487 51 525 292
rect 559 326 593 459
rect 627 425 661 527
rect 627 375 661 391
rect 708 425 811 457
rect 708 391 713 425
rect 747 391 811 425
rect 708 375 811 391
rect 559 292 659 326
rect 693 292 709 326
rect 559 288 709 292
rect 743 213 811 375
rect 565 179 581 213
rect 615 179 811 213
rect 561 108 663 124
rect 595 74 629 108
rect 561 17 663 74
rect 707 108 756 179
rect 707 74 713 108
rect 747 74 756 108
rect 707 58 756 74
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 674 289 708 323 0 FreeSans 250 0 0 0 S
port 3 nsew signal input
flabel locali s 582 289 616 323 0 FreeSans 250 0 0 0 S
port 3 nsew signal input
flabel locali s 490 153 524 187 0 FreeSans 250 0 0 0 A1
port 2 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 250 0 0 0 A1
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 250 0 0 0 A0
port 1 nsew signal input
flabel locali s 30 85 64 119 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
flabel locali s 30 357 64 391 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
flabel locali s 30 425 64 459 0 FreeSans 250 0 0 0 X
port 8 nsew signal output
flabel nwell s 74 527 108 561 0 FreeSans 250 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 84 -17 118 17 0 FreeSans 250 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 mux2_1
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 1684336
string GDS_START 1677508
string path 0.000 0.000 20.700 0.000 
<< end >>
