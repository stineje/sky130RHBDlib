VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO TMRDFFRNQNX1
  CLASS CORE ;
  FOREIGN TMRDFFRNQNX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 87.690 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.734950 ;
    PORT
      LAYER li1 ;
        RECT 85.505 5.295 85.675 6.565 ;
        RECT 86.385 5.295 86.555 6.565 ;
        RECT 85.505 5.125 87.035 5.295 ;
        RECT 86.865 1.730 87.035 5.125 ;
        RECT 86.425 1.560 87.035 1.730 ;
        RECT 79.765 1.170 79.935 1.345 ;
        RECT 79.760 1.015 79.935 1.170 ;
        RECT 79.760 0.835 79.930 1.015 ;
        RECT 83.095 0.835 83.265 1.345 ;
        RECT 86.425 0.835 86.595 1.560 ;
      LAYER mcon ;
        RECT 79.765 1.095 79.935 1.265 ;
        RECT 83.095 1.095 83.265 1.265 ;
        RECT 86.425 1.095 86.595 1.265 ;
      LAYER met1 ;
        RECT 79.735 1.265 79.965 1.295 ;
        RECT 83.065 1.265 83.295 1.295 ;
        RECT 86.395 1.265 86.625 1.295 ;
        RECT 79.705 1.095 86.655 1.265 ;
        RECT 79.735 1.065 79.965 1.095 ;
        RECT 83.065 1.065 83.295 1.095 ;
        RECT 86.395 1.065 86.625 1.095 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.044550 ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.915 7.115 4.865 ;
        RECT 32.845 1.915 33.015 4.865 ;
        RECT 58.745 1.915 58.915 4.865 ;
      LAYER mcon ;
        RECT 6.945 2.505 7.115 2.675 ;
        RECT 32.845 2.505 33.015 2.675 ;
        RECT 58.745 2.505 58.915 2.675 ;
      LAYER met1 ;
        RECT 6.915 2.675 7.145 2.705 ;
        RECT 32.815 2.675 33.045 2.705 ;
        RECT 58.715 2.675 58.945 2.705 ;
        RECT 6.885 2.505 59.095 2.675 ;
        RECT 6.915 2.475 7.145 2.505 ;
        RECT 32.815 2.475 33.045 2.505 ;
        RECT 58.715 2.475 58.945 2.505 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.089100 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
        RECT 15.085 1.915 15.255 4.865 ;
        RECT 28.035 1.915 28.205 4.865 ;
        RECT 40.985 1.915 41.155 4.865 ;
        RECT 53.935 1.915 54.105 4.865 ;
        RECT 66.885 1.915 67.055 4.865 ;
      LAYER mcon ;
        RECT 2.135 4.355 2.305 4.525 ;
        RECT 15.085 4.355 15.255 4.525 ;
        RECT 28.035 4.355 28.205 4.525 ;
        RECT 40.985 4.355 41.155 4.525 ;
        RECT 53.935 4.355 54.105 4.525 ;
        RECT 66.885 4.355 67.055 4.525 ;
      LAYER met1 ;
        RECT 2.105 4.525 2.335 4.555 ;
        RECT 15.055 4.525 15.285 4.555 ;
        RECT 28.005 4.525 28.235 4.555 ;
        RECT 40.955 4.525 41.185 4.555 ;
        RECT 53.905 4.525 54.135 4.555 ;
        RECT 66.855 4.525 67.085 4.555 ;
        RECT 2.075 4.355 67.115 4.525 ;
        RECT 2.105 4.325 2.335 4.355 ;
        RECT 15.055 4.325 15.285 4.355 ;
        RECT 28.005 4.325 28.235 4.355 ;
        RECT 40.955 4.325 41.185 4.355 ;
        RECT 53.905 4.325 54.135 4.355 ;
        RECT 66.855 4.325 67.085 4.355 ;
    END
  END CLK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.208050 ;
    PORT
      LAYER li1 ;
        RECT 8.055 1.915 8.225 4.865 ;
        RECT 16.195 1.915 16.365 4.865 ;
        RECT 19.895 1.915 20.065 4.865 ;
        RECT 33.955 1.915 34.125 4.865 ;
        RECT 42.095 1.915 42.265 4.865 ;
        RECT 45.795 1.915 45.965 4.865 ;
        RECT 59.855 1.915 60.025 4.865 ;
        RECT 67.995 1.915 68.165 4.865 ;
        RECT 71.695 1.915 71.865 4.865 ;
      LAYER mcon ;
        RECT 8.055 2.135 8.225 2.305 ;
        RECT 16.195 2.135 16.365 2.305 ;
        RECT 19.895 2.135 20.065 2.305 ;
        RECT 33.955 2.135 34.125 2.305 ;
        RECT 42.095 2.135 42.265 2.305 ;
        RECT 45.795 2.135 45.965 2.305 ;
        RECT 59.855 2.135 60.025 2.305 ;
        RECT 67.995 2.135 68.165 2.305 ;
        RECT 71.695 2.135 71.865 2.305 ;
      LAYER met1 ;
        RECT 8.025 2.305 8.255 2.335 ;
        RECT 16.165 2.305 16.395 2.335 ;
        RECT 19.865 2.305 20.095 2.335 ;
        RECT 33.925 2.305 34.155 2.335 ;
        RECT 42.065 2.305 42.295 2.335 ;
        RECT 45.765 2.305 45.995 2.335 ;
        RECT 59.825 2.305 60.055 2.335 ;
        RECT 67.965 2.305 68.195 2.335 ;
        RECT 71.665 2.305 71.895 2.335 ;
        RECT 7.995 2.135 71.925 2.305 ;
        RECT 8.025 2.105 8.255 2.135 ;
        RECT 16.165 2.105 16.395 2.135 ;
        RECT 19.865 2.105 20.095 2.135 ;
        RECT 33.925 2.105 34.155 2.135 ;
        RECT 42.065 2.105 42.295 2.135 ;
        RECT 45.765 2.105 45.995 2.135 ;
        RECT 59.825 2.105 60.055 2.135 ;
        RECT 67.965 2.105 68.195 2.135 ;
        RECT 71.665 2.105 71.895 2.135 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 88.125 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 87.860 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.815 5.215 5.985 7.230 ;
        RECT 6.695 5.555 6.865 7.230 ;
        RECT 7.575 5.555 7.745 7.230 ;
        RECT 8.455 5.555 8.625 7.230 ;
        RECT 9.450 4.110 9.790 7.230 ;
        RECT 10.325 5.135 10.495 7.230 ;
        RECT 11.205 5.555 11.375 7.230 ;
        RECT 12.085 5.555 12.255 7.230 ;
        RECT 12.780 4.110 13.120 7.230 ;
        RECT 13.955 5.215 14.125 7.230 ;
        RECT 14.835 5.555 15.005 7.230 ;
        RECT 15.715 5.555 15.885 7.230 ;
        RECT 16.595 5.555 16.765 7.230 ;
        RECT 17.590 4.110 17.930 7.230 ;
        RECT 18.765 5.215 18.935 7.230 ;
        RECT 19.645 5.555 19.815 7.230 ;
        RECT 20.525 5.555 20.695 7.230 ;
        RECT 21.405 5.555 21.575 7.230 ;
        RECT 22.400 4.110 22.740 7.230 ;
        RECT 23.275 5.135 23.445 7.230 ;
        RECT 24.155 5.555 24.325 7.230 ;
        RECT 25.035 5.555 25.205 7.230 ;
        RECT 25.730 4.110 26.070 7.230 ;
        RECT 26.905 5.215 27.075 7.230 ;
        RECT 27.785 5.555 27.955 7.230 ;
        RECT 28.665 5.555 28.835 7.230 ;
        RECT 29.545 5.555 29.715 7.230 ;
        RECT 30.540 4.110 30.880 7.230 ;
        RECT 31.715 5.215 31.885 7.230 ;
        RECT 32.595 5.555 32.765 7.230 ;
        RECT 33.475 5.555 33.645 7.230 ;
        RECT 34.355 5.555 34.525 7.230 ;
        RECT 35.350 4.110 35.690 7.230 ;
        RECT 36.225 5.135 36.395 7.230 ;
        RECT 37.105 5.555 37.275 7.230 ;
        RECT 37.985 5.555 38.155 7.230 ;
        RECT 38.680 4.110 39.020 7.230 ;
        RECT 39.855 5.215 40.025 7.230 ;
        RECT 40.735 5.555 40.905 7.230 ;
        RECT 41.615 5.555 41.785 7.230 ;
        RECT 42.495 5.555 42.665 7.230 ;
        RECT 43.490 4.110 43.830 7.230 ;
        RECT 44.665 5.215 44.835 7.230 ;
        RECT 45.545 5.555 45.715 7.230 ;
        RECT 46.425 5.555 46.595 7.230 ;
        RECT 47.305 5.555 47.475 7.230 ;
        RECT 48.300 4.110 48.640 7.230 ;
        RECT 49.175 5.135 49.345 7.230 ;
        RECT 50.055 5.555 50.225 7.230 ;
        RECT 50.935 5.555 51.105 7.230 ;
        RECT 51.630 4.110 51.970 7.230 ;
        RECT 52.805 5.215 52.975 7.230 ;
        RECT 53.685 5.555 53.855 7.230 ;
        RECT 54.565 5.555 54.735 7.230 ;
        RECT 55.445 5.555 55.615 7.230 ;
        RECT 56.440 4.110 56.780 7.230 ;
        RECT 57.615 5.215 57.785 7.230 ;
        RECT 58.495 5.555 58.665 7.230 ;
        RECT 59.375 5.555 59.545 7.230 ;
        RECT 60.255 5.555 60.425 7.230 ;
        RECT 61.250 4.110 61.590 7.230 ;
        RECT 62.125 5.135 62.295 7.230 ;
        RECT 63.005 5.555 63.175 7.230 ;
        RECT 63.885 5.555 64.055 7.230 ;
        RECT 64.580 4.110 64.920 7.230 ;
        RECT 65.755 5.215 65.925 7.230 ;
        RECT 66.635 5.555 66.805 7.230 ;
        RECT 67.515 5.555 67.685 7.230 ;
        RECT 68.395 5.555 68.565 7.230 ;
        RECT 69.390 4.110 69.730 7.230 ;
        RECT 70.565 5.215 70.735 7.230 ;
        RECT 71.445 5.555 71.615 7.230 ;
        RECT 72.325 5.555 72.495 7.230 ;
        RECT 73.205 5.555 73.375 7.230 ;
        RECT 74.200 4.110 74.540 7.230 ;
        RECT 75.075 5.135 75.245 7.230 ;
        RECT 75.955 5.555 76.125 7.230 ;
        RECT 76.835 5.555 77.005 7.230 ;
        RECT 77.530 4.110 77.870 7.230 ;
        RECT 78.405 5.125 78.575 7.230 ;
        RECT 79.285 5.555 79.455 7.230 ;
        RECT 80.165 5.125 80.335 7.230 ;
        RECT 80.860 4.110 81.200 7.230 ;
        RECT 84.190 4.110 84.530 7.230 ;
        RECT 87.520 4.110 87.860 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.015 7.315 11.185 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 13.235 7.315 13.405 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.565 7.315 16.735 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
        RECT 19.895 7.315 20.065 7.485 ;
        RECT 20.265 7.315 20.435 7.485 ;
        RECT 20.635 7.315 20.805 7.485 ;
        RECT 21.005 7.315 21.175 7.485 ;
        RECT 21.375 7.315 21.545 7.485 ;
        RECT 21.745 7.315 21.915 7.485 ;
        RECT 22.115 7.315 22.285 7.485 ;
        RECT 22.855 7.315 23.025 7.485 ;
        RECT 23.225 7.315 23.395 7.485 ;
        RECT 23.595 7.315 23.765 7.485 ;
        RECT 23.965 7.315 24.135 7.485 ;
        RECT 24.335 7.315 24.505 7.485 ;
        RECT 24.705 7.315 24.875 7.485 ;
        RECT 25.075 7.315 25.245 7.485 ;
        RECT 25.445 7.315 25.615 7.485 ;
        RECT 26.185 7.315 26.355 7.485 ;
        RECT 26.555 7.315 26.725 7.485 ;
        RECT 26.925 7.315 27.095 7.485 ;
        RECT 27.295 7.315 27.465 7.485 ;
        RECT 27.665 7.315 27.835 7.485 ;
        RECT 28.035 7.315 28.205 7.485 ;
        RECT 28.405 7.315 28.575 7.485 ;
        RECT 28.775 7.315 28.945 7.485 ;
        RECT 29.145 7.315 29.315 7.485 ;
        RECT 29.515 7.315 29.685 7.485 ;
        RECT 29.885 7.315 30.055 7.485 ;
        RECT 30.255 7.315 30.425 7.485 ;
        RECT 30.995 7.315 31.165 7.485 ;
        RECT 31.365 7.315 31.535 7.485 ;
        RECT 31.735 7.315 31.905 7.485 ;
        RECT 32.105 7.315 32.275 7.485 ;
        RECT 32.475 7.315 32.645 7.485 ;
        RECT 32.845 7.315 33.015 7.485 ;
        RECT 33.215 7.315 33.385 7.485 ;
        RECT 33.585 7.315 33.755 7.485 ;
        RECT 33.955 7.315 34.125 7.485 ;
        RECT 34.325 7.315 34.495 7.485 ;
        RECT 34.695 7.315 34.865 7.485 ;
        RECT 35.065 7.315 35.235 7.485 ;
        RECT 35.805 7.315 35.975 7.485 ;
        RECT 36.175 7.315 36.345 7.485 ;
        RECT 36.545 7.315 36.715 7.485 ;
        RECT 36.915 7.315 37.085 7.485 ;
        RECT 37.285 7.315 37.455 7.485 ;
        RECT 37.655 7.315 37.825 7.485 ;
        RECT 38.025 7.315 38.195 7.485 ;
        RECT 38.395 7.315 38.565 7.485 ;
        RECT 39.135 7.315 39.305 7.485 ;
        RECT 39.505 7.315 39.675 7.485 ;
        RECT 39.875 7.315 40.045 7.485 ;
        RECT 40.245 7.315 40.415 7.485 ;
        RECT 40.615 7.315 40.785 7.485 ;
        RECT 40.985 7.315 41.155 7.485 ;
        RECT 41.355 7.315 41.525 7.485 ;
        RECT 41.725 7.315 41.895 7.485 ;
        RECT 42.095 7.315 42.265 7.485 ;
        RECT 42.465 7.315 42.635 7.485 ;
        RECT 42.835 7.315 43.005 7.485 ;
        RECT 43.205 7.315 43.375 7.485 ;
        RECT 43.945 7.315 44.115 7.485 ;
        RECT 44.315 7.315 44.485 7.485 ;
        RECT 44.685 7.315 44.855 7.485 ;
        RECT 45.055 7.315 45.225 7.485 ;
        RECT 45.425 7.315 45.595 7.485 ;
        RECT 45.795 7.315 45.965 7.485 ;
        RECT 46.165 7.315 46.335 7.485 ;
        RECT 46.535 7.315 46.705 7.485 ;
        RECT 46.905 7.315 47.075 7.485 ;
        RECT 47.275 7.315 47.445 7.485 ;
        RECT 47.645 7.315 47.815 7.485 ;
        RECT 48.015 7.315 48.185 7.485 ;
        RECT 48.755 7.315 48.925 7.485 ;
        RECT 49.125 7.315 49.295 7.485 ;
        RECT 49.495 7.315 49.665 7.485 ;
        RECT 49.865 7.315 50.035 7.485 ;
        RECT 50.235 7.315 50.405 7.485 ;
        RECT 50.605 7.315 50.775 7.485 ;
        RECT 50.975 7.315 51.145 7.485 ;
        RECT 51.345 7.315 51.515 7.485 ;
        RECT 52.085 7.315 52.255 7.485 ;
        RECT 52.455 7.315 52.625 7.485 ;
        RECT 52.825 7.315 52.995 7.485 ;
        RECT 53.195 7.315 53.365 7.485 ;
        RECT 53.565 7.315 53.735 7.485 ;
        RECT 53.935 7.315 54.105 7.485 ;
        RECT 54.305 7.315 54.475 7.485 ;
        RECT 54.675 7.315 54.845 7.485 ;
        RECT 55.045 7.315 55.215 7.485 ;
        RECT 55.415 7.315 55.585 7.485 ;
        RECT 55.785 7.315 55.955 7.485 ;
        RECT 56.155 7.315 56.325 7.485 ;
        RECT 56.895 7.315 57.065 7.485 ;
        RECT 57.265 7.315 57.435 7.485 ;
        RECT 57.635 7.315 57.805 7.485 ;
        RECT 58.005 7.315 58.175 7.485 ;
        RECT 58.375 7.315 58.545 7.485 ;
        RECT 58.745 7.315 58.915 7.485 ;
        RECT 59.115 7.315 59.285 7.485 ;
        RECT 59.485 7.315 59.655 7.485 ;
        RECT 59.855 7.315 60.025 7.485 ;
        RECT 60.225 7.315 60.395 7.485 ;
        RECT 60.595 7.315 60.765 7.485 ;
        RECT 60.965 7.315 61.135 7.485 ;
        RECT 61.705 7.315 61.875 7.485 ;
        RECT 62.075 7.315 62.245 7.485 ;
        RECT 62.445 7.315 62.615 7.485 ;
        RECT 62.815 7.315 62.985 7.485 ;
        RECT 63.185 7.315 63.355 7.485 ;
        RECT 63.555 7.315 63.725 7.485 ;
        RECT 63.925 7.315 64.095 7.485 ;
        RECT 64.295 7.315 64.465 7.485 ;
        RECT 65.035 7.315 65.205 7.485 ;
        RECT 65.405 7.315 65.575 7.485 ;
        RECT 65.775 7.315 65.945 7.485 ;
        RECT 66.145 7.315 66.315 7.485 ;
        RECT 66.515 7.315 66.685 7.485 ;
        RECT 66.885 7.315 67.055 7.485 ;
        RECT 67.255 7.315 67.425 7.485 ;
        RECT 67.625 7.315 67.795 7.485 ;
        RECT 67.995 7.315 68.165 7.485 ;
        RECT 68.365 7.315 68.535 7.485 ;
        RECT 68.735 7.315 68.905 7.485 ;
        RECT 69.105 7.315 69.275 7.485 ;
        RECT 69.845 7.315 70.015 7.485 ;
        RECT 70.215 7.315 70.385 7.485 ;
        RECT 70.585 7.315 70.755 7.485 ;
        RECT 70.955 7.315 71.125 7.485 ;
        RECT 71.325 7.315 71.495 7.485 ;
        RECT 71.695 7.315 71.865 7.485 ;
        RECT 72.065 7.315 72.235 7.485 ;
        RECT 72.435 7.315 72.605 7.485 ;
        RECT 72.805 7.315 72.975 7.485 ;
        RECT 73.175 7.315 73.345 7.485 ;
        RECT 73.545 7.315 73.715 7.485 ;
        RECT 73.915 7.315 74.085 7.485 ;
        RECT 74.655 7.315 74.825 7.485 ;
        RECT 75.025 7.315 75.195 7.485 ;
        RECT 75.395 7.315 75.565 7.485 ;
        RECT 75.765 7.315 75.935 7.485 ;
        RECT 76.135 7.315 76.305 7.485 ;
        RECT 76.505 7.315 76.675 7.485 ;
        RECT 76.875 7.315 77.045 7.485 ;
        RECT 77.245 7.315 77.415 7.485 ;
        RECT 77.985 7.315 78.155 7.485 ;
        RECT 78.355 7.315 78.525 7.485 ;
        RECT 78.725 7.315 78.895 7.485 ;
        RECT 79.095 7.315 79.265 7.485 ;
        RECT 79.465 7.315 79.635 7.485 ;
        RECT 79.835 7.315 80.005 7.485 ;
        RECT 80.205 7.315 80.375 7.485 ;
        RECT 80.575 7.315 80.745 7.485 ;
        RECT 81.315 7.315 81.485 7.485 ;
        RECT 81.685 7.315 81.855 7.485 ;
        RECT 82.055 7.315 82.225 7.485 ;
        RECT 82.425 7.315 82.595 7.485 ;
        RECT 82.795 7.315 82.965 7.485 ;
        RECT 83.165 7.315 83.335 7.485 ;
        RECT 83.535 7.315 83.705 7.485 ;
        RECT 83.905 7.315 84.075 7.485 ;
        RECT 84.645 7.315 84.815 7.485 ;
        RECT 85.015 7.315 85.185 7.485 ;
        RECT 85.385 7.315 85.555 7.485 ;
        RECT 85.755 7.315 85.925 7.485 ;
        RECT 86.125 7.315 86.295 7.485 ;
        RECT 86.495 7.315 86.665 7.485 ;
        RECT 86.865 7.315 87.035 7.485 ;
        RECT 87.235 7.315 87.405 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 87.860 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 87.860 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.800 0.170 5.970 1.130 ;
        RECT 9.450 0.170 9.790 2.720 ;
        RECT 10.715 0.170 10.885 1.120 ;
        RECT 12.780 0.170 13.120 2.720 ;
        RECT 13.940 0.170 14.110 1.130 ;
        RECT 17.590 0.170 17.930 2.720 ;
        RECT 18.750 0.170 18.920 1.130 ;
        RECT 22.400 0.170 22.740 2.720 ;
        RECT 23.665 0.170 23.835 1.120 ;
        RECT 25.730 0.170 26.070 2.720 ;
        RECT 26.890 0.170 27.060 1.130 ;
        RECT 30.540 0.170 30.880 2.720 ;
        RECT 31.700 0.170 31.870 1.130 ;
        RECT 35.350 0.170 35.690 2.720 ;
        RECT 36.615 0.170 36.785 1.120 ;
        RECT 38.680 0.170 39.020 2.720 ;
        RECT 39.840 0.170 40.010 1.130 ;
        RECT 43.490 0.170 43.830 2.720 ;
        RECT 44.650 0.170 44.820 1.130 ;
        RECT 48.300 0.170 48.640 2.720 ;
        RECT 49.565 0.170 49.735 1.120 ;
        RECT 51.630 0.170 51.970 2.720 ;
        RECT 52.790 0.170 52.960 1.130 ;
        RECT 56.440 0.170 56.780 2.720 ;
        RECT 57.600 0.170 57.770 1.130 ;
        RECT 61.250 0.170 61.590 2.720 ;
        RECT 62.515 0.170 62.685 1.120 ;
        RECT 64.580 0.170 64.920 2.720 ;
        RECT 65.740 0.170 65.910 1.130 ;
        RECT 69.390 0.170 69.730 2.720 ;
        RECT 70.550 0.170 70.720 1.130 ;
        RECT 74.200 0.170 74.540 2.720 ;
        RECT 75.465 0.170 75.635 1.120 ;
        RECT 77.530 0.170 77.870 2.720 ;
        RECT 78.795 0.170 78.965 1.120 ;
        RECT 80.860 0.170 81.200 2.720 ;
        RECT 82.125 0.170 82.295 1.120 ;
        RECT 84.190 0.170 84.530 2.720 ;
        RECT 85.455 0.170 85.625 1.120 ;
        RECT 87.520 0.170 87.860 2.720 ;
        RECT -0.170 -0.170 87.860 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.015 -0.085 11.185 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 13.235 -0.085 13.405 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.565 -0.085 16.735 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
        RECT 19.895 -0.085 20.065 0.085 ;
        RECT 20.265 -0.085 20.435 0.085 ;
        RECT 20.635 -0.085 20.805 0.085 ;
        RECT 21.005 -0.085 21.175 0.085 ;
        RECT 21.375 -0.085 21.545 0.085 ;
        RECT 21.745 -0.085 21.915 0.085 ;
        RECT 22.115 -0.085 22.285 0.085 ;
        RECT 22.855 -0.085 23.025 0.085 ;
        RECT 23.225 -0.085 23.395 0.085 ;
        RECT 23.595 -0.085 23.765 0.085 ;
        RECT 23.965 -0.085 24.135 0.085 ;
        RECT 24.335 -0.085 24.505 0.085 ;
        RECT 24.705 -0.085 24.875 0.085 ;
        RECT 25.075 -0.085 25.245 0.085 ;
        RECT 25.445 -0.085 25.615 0.085 ;
        RECT 26.185 -0.085 26.355 0.085 ;
        RECT 26.555 -0.085 26.725 0.085 ;
        RECT 26.925 -0.085 27.095 0.085 ;
        RECT 27.295 -0.085 27.465 0.085 ;
        RECT 27.665 -0.085 27.835 0.085 ;
        RECT 28.035 -0.085 28.205 0.085 ;
        RECT 28.405 -0.085 28.575 0.085 ;
        RECT 28.775 -0.085 28.945 0.085 ;
        RECT 29.145 -0.085 29.315 0.085 ;
        RECT 29.515 -0.085 29.685 0.085 ;
        RECT 29.885 -0.085 30.055 0.085 ;
        RECT 30.255 -0.085 30.425 0.085 ;
        RECT 30.995 -0.085 31.165 0.085 ;
        RECT 31.365 -0.085 31.535 0.085 ;
        RECT 31.735 -0.085 31.905 0.085 ;
        RECT 32.105 -0.085 32.275 0.085 ;
        RECT 32.475 -0.085 32.645 0.085 ;
        RECT 32.845 -0.085 33.015 0.085 ;
        RECT 33.215 -0.085 33.385 0.085 ;
        RECT 33.585 -0.085 33.755 0.085 ;
        RECT 33.955 -0.085 34.125 0.085 ;
        RECT 34.325 -0.085 34.495 0.085 ;
        RECT 34.695 -0.085 34.865 0.085 ;
        RECT 35.065 -0.085 35.235 0.085 ;
        RECT 35.805 -0.085 35.975 0.085 ;
        RECT 36.175 -0.085 36.345 0.085 ;
        RECT 36.545 -0.085 36.715 0.085 ;
        RECT 36.915 -0.085 37.085 0.085 ;
        RECT 37.285 -0.085 37.455 0.085 ;
        RECT 37.655 -0.085 37.825 0.085 ;
        RECT 38.025 -0.085 38.195 0.085 ;
        RECT 38.395 -0.085 38.565 0.085 ;
        RECT 39.135 -0.085 39.305 0.085 ;
        RECT 39.505 -0.085 39.675 0.085 ;
        RECT 39.875 -0.085 40.045 0.085 ;
        RECT 40.245 -0.085 40.415 0.085 ;
        RECT 40.615 -0.085 40.785 0.085 ;
        RECT 40.985 -0.085 41.155 0.085 ;
        RECT 41.355 -0.085 41.525 0.085 ;
        RECT 41.725 -0.085 41.895 0.085 ;
        RECT 42.095 -0.085 42.265 0.085 ;
        RECT 42.465 -0.085 42.635 0.085 ;
        RECT 42.835 -0.085 43.005 0.085 ;
        RECT 43.205 -0.085 43.375 0.085 ;
        RECT 43.945 -0.085 44.115 0.085 ;
        RECT 44.315 -0.085 44.485 0.085 ;
        RECT 44.685 -0.085 44.855 0.085 ;
        RECT 45.055 -0.085 45.225 0.085 ;
        RECT 45.425 -0.085 45.595 0.085 ;
        RECT 45.795 -0.085 45.965 0.085 ;
        RECT 46.165 -0.085 46.335 0.085 ;
        RECT 46.535 -0.085 46.705 0.085 ;
        RECT 46.905 -0.085 47.075 0.085 ;
        RECT 47.275 -0.085 47.445 0.085 ;
        RECT 47.645 -0.085 47.815 0.085 ;
        RECT 48.015 -0.085 48.185 0.085 ;
        RECT 48.755 -0.085 48.925 0.085 ;
        RECT 49.125 -0.085 49.295 0.085 ;
        RECT 49.495 -0.085 49.665 0.085 ;
        RECT 49.865 -0.085 50.035 0.085 ;
        RECT 50.235 -0.085 50.405 0.085 ;
        RECT 50.605 -0.085 50.775 0.085 ;
        RECT 50.975 -0.085 51.145 0.085 ;
        RECT 51.345 -0.085 51.515 0.085 ;
        RECT 52.085 -0.085 52.255 0.085 ;
        RECT 52.455 -0.085 52.625 0.085 ;
        RECT 52.825 -0.085 52.995 0.085 ;
        RECT 53.195 -0.085 53.365 0.085 ;
        RECT 53.565 -0.085 53.735 0.085 ;
        RECT 53.935 -0.085 54.105 0.085 ;
        RECT 54.305 -0.085 54.475 0.085 ;
        RECT 54.675 -0.085 54.845 0.085 ;
        RECT 55.045 -0.085 55.215 0.085 ;
        RECT 55.415 -0.085 55.585 0.085 ;
        RECT 55.785 -0.085 55.955 0.085 ;
        RECT 56.155 -0.085 56.325 0.085 ;
        RECT 56.895 -0.085 57.065 0.085 ;
        RECT 57.265 -0.085 57.435 0.085 ;
        RECT 57.635 -0.085 57.805 0.085 ;
        RECT 58.005 -0.085 58.175 0.085 ;
        RECT 58.375 -0.085 58.545 0.085 ;
        RECT 58.745 -0.085 58.915 0.085 ;
        RECT 59.115 -0.085 59.285 0.085 ;
        RECT 59.485 -0.085 59.655 0.085 ;
        RECT 59.855 -0.085 60.025 0.085 ;
        RECT 60.225 -0.085 60.395 0.085 ;
        RECT 60.595 -0.085 60.765 0.085 ;
        RECT 60.965 -0.085 61.135 0.085 ;
        RECT 61.705 -0.085 61.875 0.085 ;
        RECT 62.075 -0.085 62.245 0.085 ;
        RECT 62.445 -0.085 62.615 0.085 ;
        RECT 62.815 -0.085 62.985 0.085 ;
        RECT 63.185 -0.085 63.355 0.085 ;
        RECT 63.555 -0.085 63.725 0.085 ;
        RECT 63.925 -0.085 64.095 0.085 ;
        RECT 64.295 -0.085 64.465 0.085 ;
        RECT 65.035 -0.085 65.205 0.085 ;
        RECT 65.405 -0.085 65.575 0.085 ;
        RECT 65.775 -0.085 65.945 0.085 ;
        RECT 66.145 -0.085 66.315 0.085 ;
        RECT 66.515 -0.085 66.685 0.085 ;
        RECT 66.885 -0.085 67.055 0.085 ;
        RECT 67.255 -0.085 67.425 0.085 ;
        RECT 67.625 -0.085 67.795 0.085 ;
        RECT 67.995 -0.085 68.165 0.085 ;
        RECT 68.365 -0.085 68.535 0.085 ;
        RECT 68.735 -0.085 68.905 0.085 ;
        RECT 69.105 -0.085 69.275 0.085 ;
        RECT 69.845 -0.085 70.015 0.085 ;
        RECT 70.215 -0.085 70.385 0.085 ;
        RECT 70.585 -0.085 70.755 0.085 ;
        RECT 70.955 -0.085 71.125 0.085 ;
        RECT 71.325 -0.085 71.495 0.085 ;
        RECT 71.695 -0.085 71.865 0.085 ;
        RECT 72.065 -0.085 72.235 0.085 ;
        RECT 72.435 -0.085 72.605 0.085 ;
        RECT 72.805 -0.085 72.975 0.085 ;
        RECT 73.175 -0.085 73.345 0.085 ;
        RECT 73.545 -0.085 73.715 0.085 ;
        RECT 73.915 -0.085 74.085 0.085 ;
        RECT 74.655 -0.085 74.825 0.085 ;
        RECT 75.025 -0.085 75.195 0.085 ;
        RECT 75.395 -0.085 75.565 0.085 ;
        RECT 75.765 -0.085 75.935 0.085 ;
        RECT 76.135 -0.085 76.305 0.085 ;
        RECT 76.505 -0.085 76.675 0.085 ;
        RECT 76.875 -0.085 77.045 0.085 ;
        RECT 77.245 -0.085 77.415 0.085 ;
        RECT 77.985 -0.085 78.155 0.085 ;
        RECT 78.355 -0.085 78.525 0.085 ;
        RECT 78.725 -0.085 78.895 0.085 ;
        RECT 79.095 -0.085 79.265 0.085 ;
        RECT 79.465 -0.085 79.635 0.085 ;
        RECT 79.835 -0.085 80.005 0.085 ;
        RECT 80.205 -0.085 80.375 0.085 ;
        RECT 80.575 -0.085 80.745 0.085 ;
        RECT 81.315 -0.085 81.485 0.085 ;
        RECT 81.685 -0.085 81.855 0.085 ;
        RECT 82.055 -0.085 82.225 0.085 ;
        RECT 82.425 -0.085 82.595 0.085 ;
        RECT 82.795 -0.085 82.965 0.085 ;
        RECT 83.165 -0.085 83.335 0.085 ;
        RECT 83.535 -0.085 83.705 0.085 ;
        RECT 83.905 -0.085 84.075 0.085 ;
        RECT 84.645 -0.085 84.815 0.085 ;
        RECT 85.015 -0.085 85.185 0.085 ;
        RECT 85.385 -0.085 85.555 0.085 ;
        RECT 85.755 -0.085 85.925 0.085 ;
        RECT 86.125 -0.085 86.295 0.085 ;
        RECT 86.495 -0.085 86.665 0.085 ;
        RECT 86.865 -0.085 87.035 0.085 ;
        RECT 87.235 -0.085 87.405 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 87.860 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 6.255 5.240 6.425 7.020 ;
        RECT 7.135 5.240 7.305 7.020 ;
        RECT 8.015 5.240 8.185 7.020 ;
        RECT 10.765 5.285 10.935 7.020 ;
        RECT 11.645 5.285 11.815 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 6.255 5.070 8.965 5.240 ;
        RECT 10.765 5.115 12.295 5.285 ;
        RECT 1.025 1.915 1.195 4.865 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.835 1.915 6.005 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 5.315 1.675 5.485 1.755 ;
        RECT 6.285 1.675 6.455 1.755 ;
        RECT 7.255 1.675 7.425 1.755 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 5.315 1.505 7.425 1.675 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
        RECT 5.315 0.375 5.485 1.505 ;
        RECT 6.285 0.625 6.455 1.505 ;
        RECT 7.255 1.425 7.425 1.505 ;
        RECT 6.775 1.080 6.945 1.160 ;
        RECT 7.825 1.080 7.995 1.755 ;
        RECT 8.795 1.750 8.965 5.070 ;
        RECT 10.645 1.915 10.815 4.865 ;
        RECT 11.415 4.710 11.585 4.865 ;
        RECT 11.385 4.535 11.585 4.710 ;
        RECT 11.385 1.915 11.555 4.535 ;
        RECT 6.775 0.910 7.995 1.080 ;
        RECT 6.775 0.830 6.945 0.910 ;
        RECT 7.255 0.625 7.425 0.705 ;
        RECT 6.285 0.455 7.425 0.625 ;
        RECT 6.285 0.375 6.455 0.455 ;
        RECT 7.255 0.375 7.425 0.455 ;
        RECT 7.825 0.625 7.995 0.910 ;
        RECT 8.310 1.580 8.965 1.750 ;
        RECT 10.230 1.665 10.400 1.745 ;
        RECT 11.200 1.665 11.370 1.745 ;
        RECT 12.125 1.740 12.295 5.115 ;
        RECT 14.395 5.240 14.565 7.020 ;
        RECT 15.275 5.240 15.445 7.020 ;
        RECT 16.155 5.240 16.325 7.020 ;
        RECT 19.205 5.240 19.375 7.020 ;
        RECT 20.085 5.240 20.255 7.020 ;
        RECT 20.965 5.240 21.135 7.020 ;
        RECT 23.715 5.285 23.885 7.020 ;
        RECT 24.595 5.285 24.765 7.020 ;
        RECT 14.395 5.070 17.105 5.240 ;
        RECT 19.205 5.070 21.915 5.240 ;
        RECT 23.715 5.115 25.245 5.285 ;
        RECT 13.975 1.915 14.145 4.865 ;
        RECT 8.310 0.845 8.480 1.580 ;
        RECT 10.230 1.495 11.370 1.665 ;
        RECT 8.795 0.625 8.965 1.395 ;
        RECT 7.825 0.455 8.965 0.625 ;
        RECT 7.825 0.375 7.995 0.455 ;
        RECT 8.795 0.375 8.965 0.455 ;
        RECT 10.230 0.365 10.400 1.495 ;
        RECT 11.200 0.615 11.370 1.495 ;
        RECT 11.685 1.570 12.295 1.740 ;
        RECT 13.455 1.675 13.625 1.755 ;
        RECT 14.425 1.675 14.595 1.755 ;
        RECT 15.395 1.675 15.565 1.755 ;
        RECT 11.685 0.835 11.855 1.570 ;
        RECT 13.455 1.505 15.565 1.675 ;
        RECT 12.170 0.615 12.340 1.385 ;
        RECT 11.200 0.445 12.340 0.615 ;
        RECT 11.200 0.365 11.370 0.445 ;
        RECT 12.170 0.365 12.340 0.445 ;
        RECT 13.455 0.375 13.625 1.505 ;
        RECT 14.425 0.625 14.595 1.505 ;
        RECT 15.395 1.425 15.565 1.505 ;
        RECT 14.915 1.080 15.085 1.160 ;
        RECT 15.965 1.080 16.135 1.755 ;
        RECT 16.935 1.750 17.105 5.070 ;
        RECT 18.785 1.915 18.955 4.865 ;
        RECT 21.005 1.915 21.175 4.865 ;
        RECT 14.915 0.910 16.135 1.080 ;
        RECT 14.915 0.830 15.085 0.910 ;
        RECT 15.395 0.625 15.565 0.705 ;
        RECT 14.425 0.455 15.565 0.625 ;
        RECT 14.425 0.375 14.595 0.455 ;
        RECT 15.395 0.375 15.565 0.455 ;
        RECT 15.965 0.625 16.135 0.910 ;
        RECT 16.450 1.580 17.105 1.750 ;
        RECT 18.265 1.675 18.435 1.755 ;
        RECT 19.235 1.675 19.405 1.755 ;
        RECT 20.205 1.675 20.375 1.755 ;
        RECT 16.450 0.845 16.620 1.580 ;
        RECT 18.265 1.505 20.375 1.675 ;
        RECT 16.935 0.625 17.105 1.395 ;
        RECT 15.965 0.455 17.105 0.625 ;
        RECT 15.965 0.375 16.135 0.455 ;
        RECT 16.935 0.375 17.105 0.455 ;
        RECT 18.265 0.375 18.435 1.505 ;
        RECT 19.235 0.625 19.405 1.505 ;
        RECT 20.205 1.425 20.375 1.505 ;
        RECT 19.725 1.080 19.895 1.160 ;
        RECT 20.775 1.080 20.945 1.755 ;
        RECT 21.745 1.750 21.915 5.070 ;
        RECT 23.595 1.915 23.765 4.865 ;
        RECT 24.365 4.710 24.535 4.865 ;
        RECT 24.335 4.535 24.535 4.710 ;
        RECT 24.335 1.915 24.505 4.535 ;
        RECT 19.725 0.910 20.945 1.080 ;
        RECT 19.725 0.830 19.895 0.910 ;
        RECT 20.205 0.625 20.375 0.705 ;
        RECT 19.235 0.455 20.375 0.625 ;
        RECT 19.235 0.375 19.405 0.455 ;
        RECT 20.205 0.375 20.375 0.455 ;
        RECT 20.775 0.625 20.945 0.910 ;
        RECT 21.260 1.580 21.915 1.750 ;
        RECT 23.180 1.665 23.350 1.745 ;
        RECT 24.150 1.665 24.320 1.745 ;
        RECT 25.075 1.740 25.245 5.115 ;
        RECT 27.345 5.240 27.515 7.020 ;
        RECT 28.225 5.240 28.395 7.020 ;
        RECT 29.105 5.240 29.275 7.020 ;
        RECT 32.155 5.240 32.325 7.020 ;
        RECT 33.035 5.240 33.205 7.020 ;
        RECT 33.915 5.240 34.085 7.020 ;
        RECT 36.665 5.285 36.835 7.020 ;
        RECT 37.545 5.285 37.715 7.020 ;
        RECT 27.345 5.070 30.055 5.240 ;
        RECT 32.155 5.070 34.865 5.240 ;
        RECT 36.665 5.115 38.195 5.285 ;
        RECT 26.925 1.915 27.095 4.865 ;
        RECT 29.145 1.915 29.315 4.865 ;
        RECT 21.260 0.845 21.430 1.580 ;
        RECT 23.180 1.495 24.320 1.665 ;
        RECT 21.745 0.625 21.915 1.395 ;
        RECT 20.775 0.455 21.915 0.625 ;
        RECT 20.775 0.375 20.945 0.455 ;
        RECT 21.745 0.375 21.915 0.455 ;
        RECT 23.180 0.365 23.350 1.495 ;
        RECT 24.150 0.615 24.320 1.495 ;
        RECT 24.635 1.570 25.245 1.740 ;
        RECT 26.405 1.675 26.575 1.755 ;
        RECT 27.375 1.675 27.545 1.755 ;
        RECT 28.345 1.675 28.515 1.755 ;
        RECT 24.635 0.835 24.805 1.570 ;
        RECT 26.405 1.505 28.515 1.675 ;
        RECT 25.120 0.615 25.290 1.385 ;
        RECT 24.150 0.445 25.290 0.615 ;
        RECT 24.150 0.365 24.320 0.445 ;
        RECT 25.120 0.365 25.290 0.445 ;
        RECT 26.405 0.375 26.575 1.505 ;
        RECT 27.375 0.625 27.545 1.505 ;
        RECT 28.345 1.425 28.515 1.505 ;
        RECT 27.865 1.080 28.035 1.160 ;
        RECT 28.915 1.080 29.085 1.755 ;
        RECT 29.885 1.750 30.055 5.070 ;
        RECT 31.735 1.915 31.905 4.865 ;
        RECT 27.865 0.910 29.085 1.080 ;
        RECT 27.865 0.830 28.035 0.910 ;
        RECT 28.345 0.625 28.515 0.705 ;
        RECT 27.375 0.455 28.515 0.625 ;
        RECT 27.375 0.375 27.545 0.455 ;
        RECT 28.345 0.375 28.515 0.455 ;
        RECT 28.915 0.625 29.085 0.910 ;
        RECT 29.400 1.580 30.055 1.750 ;
        RECT 31.215 1.675 31.385 1.755 ;
        RECT 32.185 1.675 32.355 1.755 ;
        RECT 33.155 1.675 33.325 1.755 ;
        RECT 29.400 0.845 29.570 1.580 ;
        RECT 31.215 1.505 33.325 1.675 ;
        RECT 29.885 0.625 30.055 1.395 ;
        RECT 28.915 0.455 30.055 0.625 ;
        RECT 28.915 0.375 29.085 0.455 ;
        RECT 29.885 0.375 30.055 0.455 ;
        RECT 31.215 0.375 31.385 1.505 ;
        RECT 32.185 0.625 32.355 1.505 ;
        RECT 33.155 1.425 33.325 1.505 ;
        RECT 32.675 1.080 32.845 1.160 ;
        RECT 33.725 1.080 33.895 1.755 ;
        RECT 34.695 1.750 34.865 5.070 ;
        RECT 36.545 1.915 36.715 4.865 ;
        RECT 37.315 4.710 37.485 4.865 ;
        RECT 37.285 4.535 37.485 4.710 ;
        RECT 37.285 1.915 37.455 4.535 ;
        RECT 32.675 0.910 33.895 1.080 ;
        RECT 32.675 0.830 32.845 0.910 ;
        RECT 33.155 0.625 33.325 0.705 ;
        RECT 32.185 0.455 33.325 0.625 ;
        RECT 32.185 0.375 32.355 0.455 ;
        RECT 33.155 0.375 33.325 0.455 ;
        RECT 33.725 0.625 33.895 0.910 ;
        RECT 34.210 1.580 34.865 1.750 ;
        RECT 36.130 1.665 36.300 1.745 ;
        RECT 37.100 1.665 37.270 1.745 ;
        RECT 38.025 1.740 38.195 5.115 ;
        RECT 40.295 5.240 40.465 7.020 ;
        RECT 41.175 5.240 41.345 7.020 ;
        RECT 42.055 5.240 42.225 7.020 ;
        RECT 45.105 5.240 45.275 7.020 ;
        RECT 45.985 5.240 46.155 7.020 ;
        RECT 46.865 5.240 47.035 7.020 ;
        RECT 49.615 5.285 49.785 7.020 ;
        RECT 50.495 5.285 50.665 7.020 ;
        RECT 40.295 5.070 43.005 5.240 ;
        RECT 45.105 5.070 47.815 5.240 ;
        RECT 49.615 5.115 51.145 5.285 ;
        RECT 39.875 1.915 40.045 4.865 ;
        RECT 34.210 0.845 34.380 1.580 ;
        RECT 36.130 1.495 37.270 1.665 ;
        RECT 34.695 0.625 34.865 1.395 ;
        RECT 33.725 0.455 34.865 0.625 ;
        RECT 33.725 0.375 33.895 0.455 ;
        RECT 34.695 0.375 34.865 0.455 ;
        RECT 36.130 0.365 36.300 1.495 ;
        RECT 37.100 0.615 37.270 1.495 ;
        RECT 37.585 1.570 38.195 1.740 ;
        RECT 39.355 1.675 39.525 1.755 ;
        RECT 40.325 1.675 40.495 1.755 ;
        RECT 41.295 1.675 41.465 1.755 ;
        RECT 37.585 0.835 37.755 1.570 ;
        RECT 39.355 1.505 41.465 1.675 ;
        RECT 38.070 0.615 38.240 1.385 ;
        RECT 37.100 0.445 38.240 0.615 ;
        RECT 37.100 0.365 37.270 0.445 ;
        RECT 38.070 0.365 38.240 0.445 ;
        RECT 39.355 0.375 39.525 1.505 ;
        RECT 40.325 0.625 40.495 1.505 ;
        RECT 41.295 1.425 41.465 1.505 ;
        RECT 40.815 1.080 40.985 1.160 ;
        RECT 41.865 1.080 42.035 1.755 ;
        RECT 42.835 1.750 43.005 5.070 ;
        RECT 44.685 1.915 44.855 4.865 ;
        RECT 46.905 1.915 47.075 4.865 ;
        RECT 40.815 0.910 42.035 1.080 ;
        RECT 40.815 0.830 40.985 0.910 ;
        RECT 41.295 0.625 41.465 0.705 ;
        RECT 40.325 0.455 41.465 0.625 ;
        RECT 40.325 0.375 40.495 0.455 ;
        RECT 41.295 0.375 41.465 0.455 ;
        RECT 41.865 0.625 42.035 0.910 ;
        RECT 42.350 1.580 43.005 1.750 ;
        RECT 44.165 1.675 44.335 1.755 ;
        RECT 45.135 1.675 45.305 1.755 ;
        RECT 46.105 1.675 46.275 1.755 ;
        RECT 42.350 0.845 42.520 1.580 ;
        RECT 44.165 1.505 46.275 1.675 ;
        RECT 42.835 0.625 43.005 1.395 ;
        RECT 41.865 0.455 43.005 0.625 ;
        RECT 41.865 0.375 42.035 0.455 ;
        RECT 42.835 0.375 43.005 0.455 ;
        RECT 44.165 0.375 44.335 1.505 ;
        RECT 45.135 0.625 45.305 1.505 ;
        RECT 46.105 1.425 46.275 1.505 ;
        RECT 45.625 1.080 45.795 1.160 ;
        RECT 46.675 1.080 46.845 1.755 ;
        RECT 47.645 1.750 47.815 5.070 ;
        RECT 49.495 1.915 49.665 4.865 ;
        RECT 50.265 4.710 50.435 4.865 ;
        RECT 50.235 4.535 50.435 4.710 ;
        RECT 50.235 1.915 50.405 4.535 ;
        RECT 45.625 0.910 46.845 1.080 ;
        RECT 45.625 0.830 45.795 0.910 ;
        RECT 46.105 0.625 46.275 0.705 ;
        RECT 45.135 0.455 46.275 0.625 ;
        RECT 45.135 0.375 45.305 0.455 ;
        RECT 46.105 0.375 46.275 0.455 ;
        RECT 46.675 0.625 46.845 0.910 ;
        RECT 47.160 1.580 47.815 1.750 ;
        RECT 49.080 1.665 49.250 1.745 ;
        RECT 50.050 1.665 50.220 1.745 ;
        RECT 50.975 1.740 51.145 5.115 ;
        RECT 53.245 5.240 53.415 7.020 ;
        RECT 54.125 5.240 54.295 7.020 ;
        RECT 55.005 5.240 55.175 7.020 ;
        RECT 58.055 5.240 58.225 7.020 ;
        RECT 58.935 5.240 59.105 7.020 ;
        RECT 59.815 5.240 59.985 7.020 ;
        RECT 62.565 5.285 62.735 7.020 ;
        RECT 63.445 5.285 63.615 7.020 ;
        RECT 53.245 5.070 55.955 5.240 ;
        RECT 58.055 5.070 60.765 5.240 ;
        RECT 62.565 5.115 64.095 5.285 ;
        RECT 52.825 1.915 52.995 4.865 ;
        RECT 55.045 1.915 55.215 4.865 ;
        RECT 47.160 0.845 47.330 1.580 ;
        RECT 49.080 1.495 50.220 1.665 ;
        RECT 47.645 0.625 47.815 1.395 ;
        RECT 46.675 0.455 47.815 0.625 ;
        RECT 46.675 0.375 46.845 0.455 ;
        RECT 47.645 0.375 47.815 0.455 ;
        RECT 49.080 0.365 49.250 1.495 ;
        RECT 50.050 0.615 50.220 1.495 ;
        RECT 50.535 1.570 51.145 1.740 ;
        RECT 52.305 1.675 52.475 1.755 ;
        RECT 53.275 1.675 53.445 1.755 ;
        RECT 54.245 1.675 54.415 1.755 ;
        RECT 50.535 0.835 50.705 1.570 ;
        RECT 52.305 1.505 54.415 1.675 ;
        RECT 51.020 0.615 51.190 1.385 ;
        RECT 50.050 0.445 51.190 0.615 ;
        RECT 50.050 0.365 50.220 0.445 ;
        RECT 51.020 0.365 51.190 0.445 ;
        RECT 52.305 0.375 52.475 1.505 ;
        RECT 53.275 0.625 53.445 1.505 ;
        RECT 54.245 1.425 54.415 1.505 ;
        RECT 53.765 1.080 53.935 1.160 ;
        RECT 54.815 1.080 54.985 1.755 ;
        RECT 55.785 1.750 55.955 5.070 ;
        RECT 57.635 1.915 57.805 4.865 ;
        RECT 53.765 0.910 54.985 1.080 ;
        RECT 53.765 0.830 53.935 0.910 ;
        RECT 54.245 0.625 54.415 0.705 ;
        RECT 53.275 0.455 54.415 0.625 ;
        RECT 53.275 0.375 53.445 0.455 ;
        RECT 54.245 0.375 54.415 0.455 ;
        RECT 54.815 0.625 54.985 0.910 ;
        RECT 55.300 1.580 55.955 1.750 ;
        RECT 57.115 1.675 57.285 1.755 ;
        RECT 58.085 1.675 58.255 1.755 ;
        RECT 59.055 1.675 59.225 1.755 ;
        RECT 55.300 0.845 55.470 1.580 ;
        RECT 57.115 1.505 59.225 1.675 ;
        RECT 55.785 0.625 55.955 1.395 ;
        RECT 54.815 0.455 55.955 0.625 ;
        RECT 54.815 0.375 54.985 0.455 ;
        RECT 55.785 0.375 55.955 0.455 ;
        RECT 57.115 0.375 57.285 1.505 ;
        RECT 58.085 0.625 58.255 1.505 ;
        RECT 59.055 1.425 59.225 1.505 ;
        RECT 58.575 1.080 58.745 1.160 ;
        RECT 59.625 1.080 59.795 1.755 ;
        RECT 60.595 1.750 60.765 5.070 ;
        RECT 62.445 1.915 62.615 4.865 ;
        RECT 63.215 4.710 63.385 4.865 ;
        RECT 63.185 4.535 63.385 4.710 ;
        RECT 63.185 1.915 63.355 4.535 ;
        RECT 58.575 0.910 59.795 1.080 ;
        RECT 58.575 0.830 58.745 0.910 ;
        RECT 59.055 0.625 59.225 0.705 ;
        RECT 58.085 0.455 59.225 0.625 ;
        RECT 58.085 0.375 58.255 0.455 ;
        RECT 59.055 0.375 59.225 0.455 ;
        RECT 59.625 0.625 59.795 0.910 ;
        RECT 60.110 1.580 60.765 1.750 ;
        RECT 62.030 1.665 62.200 1.745 ;
        RECT 63.000 1.665 63.170 1.745 ;
        RECT 63.925 1.740 64.095 5.115 ;
        RECT 66.195 5.240 66.365 7.020 ;
        RECT 67.075 5.240 67.245 7.020 ;
        RECT 67.955 5.240 68.125 7.020 ;
        RECT 71.005 5.240 71.175 7.020 ;
        RECT 71.885 5.240 72.055 7.020 ;
        RECT 72.765 5.240 72.935 7.020 ;
        RECT 75.515 5.285 75.685 7.020 ;
        RECT 76.395 5.285 76.565 7.020 ;
        RECT 78.845 6.825 79.025 6.995 ;
        RECT 78.845 5.295 79.015 6.825 ;
        RECT 79.725 5.295 79.895 6.995 ;
        RECT 66.195 5.070 68.905 5.240 ;
        RECT 71.005 5.070 73.715 5.240 ;
        RECT 75.515 5.115 77.045 5.285 ;
        RECT 78.845 5.125 79.895 5.295 ;
        RECT 65.775 1.915 65.945 4.865 ;
        RECT 60.110 0.845 60.280 1.580 ;
        RECT 62.030 1.495 63.170 1.665 ;
        RECT 60.595 0.625 60.765 1.395 ;
        RECT 59.625 0.455 60.765 0.625 ;
        RECT 59.625 0.375 59.795 0.455 ;
        RECT 60.595 0.375 60.765 0.455 ;
        RECT 62.030 0.365 62.200 1.495 ;
        RECT 63.000 0.615 63.170 1.495 ;
        RECT 63.485 1.570 64.095 1.740 ;
        RECT 65.255 1.675 65.425 1.755 ;
        RECT 66.225 1.675 66.395 1.755 ;
        RECT 67.195 1.675 67.365 1.755 ;
        RECT 63.485 0.835 63.655 1.570 ;
        RECT 65.255 1.505 67.365 1.675 ;
        RECT 63.970 0.615 64.140 1.385 ;
        RECT 63.000 0.445 64.140 0.615 ;
        RECT 63.000 0.365 63.170 0.445 ;
        RECT 63.970 0.365 64.140 0.445 ;
        RECT 65.255 0.375 65.425 1.505 ;
        RECT 66.225 0.625 66.395 1.505 ;
        RECT 67.195 1.425 67.365 1.505 ;
        RECT 66.715 1.080 66.885 1.160 ;
        RECT 67.765 1.080 67.935 1.755 ;
        RECT 68.735 1.750 68.905 5.070 ;
        RECT 70.585 1.915 70.755 4.865 ;
        RECT 72.805 1.915 72.975 4.865 ;
        RECT 66.715 0.910 67.935 1.080 ;
        RECT 66.715 0.830 66.885 0.910 ;
        RECT 67.195 0.625 67.365 0.705 ;
        RECT 66.225 0.455 67.365 0.625 ;
        RECT 66.225 0.375 66.395 0.455 ;
        RECT 67.195 0.375 67.365 0.455 ;
        RECT 67.765 0.625 67.935 0.910 ;
        RECT 68.250 1.580 68.905 1.750 ;
        RECT 70.065 1.675 70.235 1.755 ;
        RECT 71.035 1.675 71.205 1.755 ;
        RECT 72.005 1.675 72.175 1.755 ;
        RECT 68.250 0.845 68.420 1.580 ;
        RECT 70.065 1.505 72.175 1.675 ;
        RECT 68.735 0.625 68.905 1.395 ;
        RECT 67.765 0.455 68.905 0.625 ;
        RECT 67.765 0.375 67.935 0.455 ;
        RECT 68.735 0.375 68.905 0.455 ;
        RECT 70.065 0.375 70.235 1.505 ;
        RECT 71.035 0.625 71.205 1.505 ;
        RECT 72.005 1.425 72.175 1.505 ;
        RECT 71.525 1.080 71.695 1.160 ;
        RECT 72.575 1.080 72.745 1.755 ;
        RECT 73.545 1.750 73.715 5.070 ;
        RECT 75.395 1.915 75.565 4.865 ;
        RECT 76.165 4.710 76.335 4.865 ;
        RECT 76.135 4.535 76.335 4.710 ;
        RECT 76.135 1.915 76.305 4.535 ;
        RECT 71.525 0.910 72.745 1.080 ;
        RECT 71.525 0.830 71.695 0.910 ;
        RECT 72.005 0.625 72.175 0.705 ;
        RECT 71.035 0.455 72.175 0.625 ;
        RECT 71.035 0.375 71.205 0.455 ;
        RECT 72.005 0.375 72.175 0.455 ;
        RECT 72.575 0.625 72.745 0.910 ;
        RECT 73.060 1.580 73.715 1.750 ;
        RECT 74.980 1.665 75.150 1.745 ;
        RECT 75.950 1.665 76.120 1.745 ;
        RECT 76.875 1.740 77.045 5.115 ;
        RECT 79.725 5.045 79.895 5.125 ;
        RECT 81.725 6.825 83.655 6.995 ;
        RECT 81.725 5.045 81.895 6.825 ;
        RECT 82.165 5.295 82.335 6.565 ;
        RECT 82.605 5.555 82.775 6.825 ;
        RECT 83.045 5.295 83.215 6.565 ;
        RECT 83.485 5.375 83.655 6.825 ;
        RECT 85.065 6.825 86.995 6.995 ;
        RECT 82.165 5.125 83.215 5.295 ;
        RECT 83.045 5.045 83.215 5.125 ;
        RECT 85.065 5.045 85.235 6.825 ;
        RECT 85.945 5.555 86.115 6.825 ;
        RECT 86.825 5.555 86.995 6.825 ;
        RECT 78.355 1.915 78.525 4.870 ;
        RECT 79.505 4.710 79.675 4.870 ;
        RECT 79.465 4.540 79.675 4.710 ;
        RECT 79.465 1.915 79.635 4.540 ;
        RECT 82.055 1.915 82.225 4.870 ;
        RECT 83.535 1.915 83.705 4.870 ;
        RECT 85.015 1.915 85.185 4.870 ;
        RECT 86.125 4.540 86.315 4.870 ;
        RECT 86.125 1.915 86.295 4.540 ;
        RECT 73.060 0.845 73.230 1.580 ;
        RECT 74.980 1.495 76.120 1.665 ;
        RECT 73.545 0.625 73.715 1.395 ;
        RECT 72.575 0.455 73.715 0.625 ;
        RECT 72.575 0.375 72.745 0.455 ;
        RECT 73.545 0.375 73.715 0.455 ;
        RECT 74.980 0.365 75.150 1.495 ;
        RECT 75.950 0.615 76.120 1.495 ;
        RECT 76.435 1.570 77.045 1.740 ;
        RECT 78.310 1.665 78.480 1.745 ;
        RECT 79.280 1.665 79.450 1.745 ;
        RECT 76.435 0.835 76.605 1.570 ;
        RECT 78.310 1.495 79.450 1.665 ;
        RECT 76.920 0.615 77.090 1.385 ;
        RECT 75.950 0.445 77.090 0.615 ;
        RECT 75.950 0.365 76.120 0.445 ;
        RECT 76.920 0.365 77.090 0.445 ;
        RECT 78.310 0.365 78.480 1.495 ;
        RECT 79.280 0.615 79.450 1.495 ;
        RECT 80.250 0.615 80.420 1.745 ;
        RECT 79.280 0.445 80.420 0.615 ;
        RECT 79.280 0.365 79.450 0.445 ;
        RECT 80.250 0.365 80.420 0.445 ;
        RECT 81.640 1.665 81.810 1.745 ;
        RECT 82.610 1.665 82.780 1.745 ;
        RECT 81.640 1.495 82.780 1.665 ;
        RECT 81.640 0.365 81.810 1.495 ;
        RECT 82.610 0.615 82.780 1.495 ;
        RECT 83.580 0.615 83.750 1.745 ;
        RECT 82.610 0.445 83.750 0.615 ;
        RECT 82.610 0.365 82.780 0.445 ;
        RECT 83.580 0.365 83.750 0.445 ;
        RECT 84.970 1.665 85.140 1.745 ;
        RECT 85.940 1.665 86.110 1.745 ;
        RECT 84.970 1.495 86.110 1.665 ;
        RECT 84.970 0.365 85.140 1.495 ;
        RECT 85.940 0.615 86.110 1.495 ;
        RECT 86.910 0.615 87.080 1.390 ;
        RECT 85.940 0.445 87.080 0.615 ;
        RECT 85.940 0.365 86.110 0.445 ;
        RECT 86.910 0.365 87.080 0.445 ;
      LAYER mcon ;
        RECT 1.025 3.985 1.195 4.155 ;
        RECT 3.245 3.245 3.415 3.415 ;
        RECT 3.985 3.615 4.155 3.785 ;
        RECT 5.835 3.615 6.005 3.785 ;
        RECT 8.795 3.245 8.965 3.415 ;
        RECT 10.645 3.245 10.815 3.415 ;
        RECT 11.385 3.985 11.555 4.155 ;
        RECT 12.125 3.245 12.295 3.415 ;
        RECT 13.975 3.245 14.145 3.415 ;
        RECT 16.935 3.985 17.105 4.155 ;
        RECT 18.785 3.615 18.955 3.785 ;
        RECT 21.005 2.875 21.175 3.045 ;
        RECT 21.745 3.985 21.915 4.155 ;
        RECT 23.595 3.985 23.765 4.155 ;
        RECT 24.335 3.985 24.505 4.155 ;
        RECT 25.075 2.875 25.245 3.045 ;
        RECT 26.925 3.985 27.095 4.155 ;
        RECT 29.145 3.245 29.315 3.415 ;
        RECT 29.885 3.615 30.055 3.785 ;
        RECT 31.735 3.615 31.905 3.785 ;
        RECT 34.695 3.245 34.865 3.415 ;
        RECT 36.545 3.245 36.715 3.415 ;
        RECT 37.285 3.985 37.455 4.155 ;
        RECT 38.025 3.245 38.195 3.415 ;
        RECT 39.875 3.245 40.045 3.415 ;
        RECT 42.835 3.985 43.005 4.155 ;
        RECT 44.685 3.615 44.855 3.785 ;
        RECT 46.905 3.245 47.075 3.415 ;
        RECT 47.645 3.615 47.815 3.785 ;
        RECT 49.495 3.615 49.665 3.785 ;
        RECT 50.235 3.985 50.405 4.155 ;
        RECT 50.975 3.245 51.145 3.415 ;
        RECT 52.825 3.985 52.995 4.155 ;
        RECT 55.045 3.245 55.215 3.415 ;
        RECT 55.785 3.615 55.955 3.785 ;
        RECT 57.635 3.615 57.805 3.785 ;
        RECT 60.595 3.245 60.765 3.415 ;
        RECT 62.445 3.245 62.615 3.415 ;
        RECT 63.185 3.985 63.355 4.155 ;
        RECT 79.725 5.125 79.895 5.295 ;
        RECT 63.925 3.245 64.095 3.415 ;
        RECT 65.775 3.245 65.945 3.415 ;
        RECT 68.735 3.985 68.905 4.155 ;
        RECT 70.585 3.615 70.755 3.785 ;
        RECT 72.805 3.615 72.975 3.785 ;
        RECT 73.545 3.985 73.715 4.155 ;
        RECT 75.395 3.985 75.565 4.155 ;
        RECT 76.135 3.985 76.305 4.155 ;
        RECT 81.725 5.125 81.895 5.295 ;
        RECT 83.045 5.125 83.215 5.295 ;
        RECT 85.065 5.125 85.235 5.295 ;
        RECT 76.875 3.615 77.045 3.785 ;
        RECT 78.355 4.355 78.525 4.525 ;
        RECT 78.355 3.245 78.525 3.415 ;
        RECT 79.465 3.985 79.635 4.155 ;
        RECT 79.465 3.615 79.635 3.785 ;
        RECT 82.055 4.355 82.225 4.525 ;
        RECT 83.535 2.875 83.705 3.045 ;
        RECT 83.535 1.995 83.705 2.165 ;
        RECT 85.015 1.995 85.185 2.165 ;
        RECT 86.125 3.985 86.295 4.155 ;
      LAYER met1 ;
        RECT 79.695 5.295 79.925 5.325 ;
        RECT 81.695 5.295 81.925 5.325 ;
        RECT 83.015 5.295 83.245 5.325 ;
        RECT 85.035 5.295 85.265 5.325 ;
        RECT 79.665 5.125 81.955 5.295 ;
        RECT 82.985 5.125 85.295 5.295 ;
        RECT 79.695 5.095 79.925 5.125 ;
        RECT 81.695 5.095 81.925 5.125 ;
        RECT 83.015 5.095 83.245 5.125 ;
        RECT 85.035 5.095 85.265 5.125 ;
        RECT 78.325 4.525 78.555 4.555 ;
        RECT 82.025 4.525 82.255 4.555 ;
        RECT 78.295 4.355 82.285 4.525 ;
        RECT 78.325 4.325 78.555 4.355 ;
        RECT 82.025 4.325 82.255 4.355 ;
        RECT 0.995 4.155 1.225 4.185 ;
        RECT 11.355 4.155 11.585 4.185 ;
        RECT 16.905 4.155 17.135 4.185 ;
        RECT 21.715 4.155 21.945 4.185 ;
        RECT 23.565 4.155 23.795 4.185 ;
        RECT 24.305 4.155 24.535 4.185 ;
        RECT 26.895 4.155 27.125 4.185 ;
        RECT 37.255 4.155 37.485 4.185 ;
        RECT 42.805 4.155 43.035 4.185 ;
        RECT 50.205 4.155 50.435 4.185 ;
        RECT 52.795 4.155 53.025 4.185 ;
        RECT 63.155 4.155 63.385 4.185 ;
        RECT 68.705 4.155 68.935 4.185 ;
        RECT 73.515 4.155 73.745 4.185 ;
        RECT 75.365 4.155 75.595 4.185 ;
        RECT 76.105 4.155 76.335 4.185 ;
        RECT 79.435 4.155 79.665 4.185 ;
        RECT 86.095 4.155 86.325 4.185 ;
        RECT 0.965 3.985 24.565 4.155 ;
        RECT 26.865 3.985 50.465 4.155 ;
        RECT 52.765 3.985 76.365 4.155 ;
        RECT 79.405 3.985 86.355 4.155 ;
        RECT 0.995 3.955 1.225 3.985 ;
        RECT 11.355 3.955 11.585 3.985 ;
        RECT 16.905 3.955 17.135 3.985 ;
        RECT 21.715 3.955 21.945 3.985 ;
        RECT 23.565 3.955 23.795 3.985 ;
        RECT 24.305 3.955 24.535 3.985 ;
        RECT 26.895 3.955 27.125 3.985 ;
        RECT 37.255 3.955 37.485 3.985 ;
        RECT 42.805 3.955 43.035 3.985 ;
        RECT 50.205 3.955 50.435 3.985 ;
        RECT 52.795 3.955 53.025 3.985 ;
        RECT 63.155 3.955 63.385 3.985 ;
        RECT 68.705 3.955 68.935 3.985 ;
        RECT 73.515 3.955 73.745 3.985 ;
        RECT 75.365 3.955 75.595 3.985 ;
        RECT 76.105 3.955 76.335 3.985 ;
        RECT 79.435 3.955 79.665 3.985 ;
        RECT 86.095 3.955 86.325 3.985 ;
        RECT 3.955 3.785 4.185 3.815 ;
        RECT 5.805 3.785 6.035 3.815 ;
        RECT 18.755 3.785 18.985 3.815 ;
        RECT 29.855 3.785 30.085 3.815 ;
        RECT 31.705 3.785 31.935 3.815 ;
        RECT 44.655 3.785 44.885 3.815 ;
        RECT 47.615 3.785 47.845 3.815 ;
        RECT 49.465 3.785 49.695 3.815 ;
        RECT 55.755 3.785 55.985 3.815 ;
        RECT 57.605 3.785 57.835 3.815 ;
        RECT 70.555 3.785 70.785 3.815 ;
        RECT 72.775 3.785 73.005 3.815 ;
        RECT 76.845 3.785 77.075 3.815 ;
        RECT 79.435 3.785 79.665 3.815 ;
        RECT 3.925 3.615 19.015 3.785 ;
        RECT 29.825 3.615 44.915 3.785 ;
        RECT 47.585 3.615 49.725 3.785 ;
        RECT 55.725 3.615 70.815 3.785 ;
        RECT 72.745 3.615 79.695 3.785 ;
        RECT 3.955 3.585 4.185 3.615 ;
        RECT 5.805 3.585 6.035 3.615 ;
        RECT 18.755 3.585 18.985 3.615 ;
        RECT 29.855 3.585 30.085 3.615 ;
        RECT 31.705 3.585 31.935 3.615 ;
        RECT 44.655 3.585 44.885 3.615 ;
        RECT 47.615 3.585 47.845 3.615 ;
        RECT 49.465 3.585 49.695 3.615 ;
        RECT 55.755 3.585 55.985 3.615 ;
        RECT 57.605 3.585 57.835 3.615 ;
        RECT 70.555 3.585 70.785 3.615 ;
        RECT 72.775 3.585 73.005 3.615 ;
        RECT 76.845 3.585 77.075 3.615 ;
        RECT 79.435 3.585 79.665 3.615 ;
        RECT 3.215 3.415 3.445 3.445 ;
        RECT 8.765 3.415 8.995 3.445 ;
        RECT 10.615 3.415 10.845 3.445 ;
        RECT 12.095 3.415 12.325 3.445 ;
        RECT 13.945 3.415 14.175 3.445 ;
        RECT 29.115 3.415 29.345 3.445 ;
        RECT 34.665 3.415 34.895 3.445 ;
        RECT 36.515 3.415 36.745 3.445 ;
        RECT 37.995 3.415 38.225 3.445 ;
        RECT 39.845 3.415 40.075 3.445 ;
        RECT 46.875 3.415 47.105 3.445 ;
        RECT 50.945 3.415 51.175 3.445 ;
        RECT 55.015 3.415 55.245 3.445 ;
        RECT 60.565 3.415 60.795 3.445 ;
        RECT 62.415 3.415 62.645 3.445 ;
        RECT 63.895 3.415 64.125 3.445 ;
        RECT 65.745 3.415 65.975 3.445 ;
        RECT 78.325 3.415 78.555 3.445 ;
        RECT 3.185 3.245 10.875 3.415 ;
        RECT 12.065 3.245 14.205 3.415 ;
        RECT 29.085 3.245 36.775 3.415 ;
        RECT 37.965 3.245 40.105 3.415 ;
        RECT 46.845 3.245 78.585 3.415 ;
        RECT 3.215 3.215 3.445 3.245 ;
        RECT 8.765 3.215 8.995 3.245 ;
        RECT 10.615 3.215 10.845 3.245 ;
        RECT 12.095 3.215 12.325 3.245 ;
        RECT 13.945 3.215 14.175 3.245 ;
        RECT 29.115 3.215 29.345 3.245 ;
        RECT 34.665 3.215 34.895 3.245 ;
        RECT 36.515 3.215 36.745 3.245 ;
        RECT 37.995 3.215 38.225 3.245 ;
        RECT 39.845 3.215 40.075 3.245 ;
        RECT 46.875 3.215 47.105 3.245 ;
        RECT 50.945 3.215 51.175 3.245 ;
        RECT 55.015 3.215 55.245 3.245 ;
        RECT 60.565 3.215 60.795 3.245 ;
        RECT 62.415 3.215 62.645 3.245 ;
        RECT 63.895 3.215 64.125 3.245 ;
        RECT 65.745 3.215 65.975 3.245 ;
        RECT 78.325 3.215 78.555 3.245 ;
        RECT 20.975 3.045 21.205 3.075 ;
        RECT 25.045 3.045 25.275 3.075 ;
        RECT 83.505 3.045 83.735 3.075 ;
        RECT 20.945 2.875 83.765 3.045 ;
        RECT 20.975 2.845 21.205 2.875 ;
        RECT 25.045 2.845 25.275 2.875 ;
        RECT 83.505 2.845 83.735 2.875 ;
        RECT 83.505 2.165 83.735 2.195 ;
        RECT 84.985 2.165 85.215 2.195 ;
        RECT 83.475 1.995 85.245 2.165 ;
        RECT 83.505 1.965 83.735 1.995 ;
        RECT 84.985 1.965 85.215 1.995 ;
  END
END TMRDFFRNQNX1
END LIBRARY

