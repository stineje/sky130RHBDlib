* SPICE3 file created from TMRDFFSNQNX1.ext - technology: sky130A

.subckt TMRDFFSNQNX1 D CLK SN QN VNB VPB
M1000 VPB.t48 CLK a_5227_383.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_15533_1005.t5 a_3473_1004.t5 a_15044_181.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VNB D a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=3.7611p pd=32.97u as=0p ps=0u
M1003 a_3599_383.t6 SN VPB.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VNB a_343_383.t11 a_3368_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1005 VNB a_9985_1004.t8 a_11487_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t42 CLK a_11033_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t1 a_8357_1004.t5 a_8483_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_5227_383.t1 CLK VPB.t47 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_14869_1005.t5 a_3473_1004.t6 a_15533_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t39 D a_217_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPB.t4 a_1265_943.t5 a_1905_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t37 D a_5101_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_9985_1004.t3 a_10111_383.t7 VPB.t72 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPB.t85 a_5101_1004.t5 a_6789_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_15533_1005.t1 a_8357_1004.t6 a_15044_181.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_6789_1004.t5 a_6149_943.t6 VPB.t89 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t13 a_11033_943.t6 a_11673_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_3599_383.t1 a_1265_943.t6 VPB.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_13241_1004.t4 a_10111_383.t9 VPB.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VNB D a_9880_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1905_1004.t4 a_217_1004.t6 VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t93 a_11673_1004.t7 a_11033_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_14869_1005.t7 a_13241_1004.t5 a_15533_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPB.t59 a_343_383.t7 a_217_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPB.t30 a_5227_383.t7 a_5101_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_11673_1004.t2 a_11033_943.t7 VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPB.t68 a_217_1004.t7 a_343_383.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPB.t40 a_13241_1004.t7 a_13367_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_3473_1004.t2 a_3599_383.t7 VPB.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_10111_383.t3 CLK VPB.t46 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 VNB a_217_1004.t10 a_757_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_5227_383.t5 a_6149_943.t7 VPB.t91 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPB.t64 a_11033_943.t9 a_10111_383.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_13241_1004.t2 a_13367_383.t7 VPB.t63 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPB.t33 a_5227_383.t9 a_8357_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 VNB a_1905_1004.t7 a_2702_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_6149_943.t3 CLK VPB.t52 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_14869_1005.t0 a_13241_1004.t9 VPB.t53 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VNB a_10111_383.t10 a_13136_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_13367_383.t0 a_13241_1004.t10 VPB.t57 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPB.t92 a_6149_943.t8 a_8483_383.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VNB a_5227_383.t8 a_8252_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1043 VNB a_8357_1004.t13 a_8897_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPB.t26 a_8357_1004.t7 a_14869_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 VPB.t49 CLK a_343_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_3473_1004.t4 a_343_383.t9 VPB.t86 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPB.t5 a_1905_1004.t8 a_1265_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_8483_383.t3 SN VPB.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPB.t83 SN a_13367_383.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_10111_383.t0 a_9985_1004.t5 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_15533_1005.t6 a_13241_1004.t11 a_14869_1005.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 VPB.t15 a_10111_383.t11 a_9985_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 VNB a_13241_1004.t8 a_14764_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1054 VPB.t79 SN a_11673_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_6149_943.t1 a_6789_1004.t7 VPB.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 VPB.t58 a_3473_1004.t9 a_3599_383.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 VPB.t3 a_1265_943.t8 a_3599_383.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 VNB a_217_1004.t5 a_1719_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1059 VPB.t0 a_1265_943.t9 a_343_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 a_8483_383.t0 a_8357_1004.t9 VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 VPB.t16 a_11033_943.t10 a_13367_383.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 VPB.t65 a_5101_1004.t8 a_5227_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_15533_1005.t2 a_3473_1004.t11 a_14869_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_8483_383.t4 a_6149_943.t9 VPB.t87 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 a_217_1004.t0 D VPB.t38 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 VPB.t34 D a_9985_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_1905_1004.t0 a_1265_943.t10 VPB.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_6789_1004.t0 a_5101_1004.t9 VPB.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 VPB.t10 a_9985_1004.t7 a_11673_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_15044_181.t0 a_8357_1004.t10 a_15533_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 VPB.t76 SN a_3599_383.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 VPB.t78 SN a_6789_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 VNB a_6789_1004.t8 a_7586_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1074 VNB a_3473_1004.t10 a_16096_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1075 VNB D a_4996_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1076 a_11033_943.t3 a_11673_1004.t8 VPB.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 VNB a_13241_1004.t6 a_13781_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1078 a_1905_1004.t6 SN VPB.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 a_5101_1004.t0 a_5227_383.t10 VPB.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_217_1004.t3 a_343_383.t10 VPB.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 VNB a_5101_1004.t6 a_5641_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1082 a_6789_1004.t1 SN VPB.t77 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_15044_181.t6 a_3473_1004.t12 a_15533_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 VPB.t24 a_9985_1004.t9 a_10111_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 VPB.t8 a_8483_383.t8 a_8357_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_343_383.t5 a_217_1004.t8 VPB.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 VPB.t88 a_6149_943.t11 a_6789_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 VPB.t69 a_10111_383.t12 a_13241_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_10111_383.t4 a_11033_943.t11 VPB.t70 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 a_8357_1004.t3 a_5227_383.t11 VPB.t32 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 VPB.t67 a_217_1004.t9 a_1905_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 VPB.t27 a_6789_1004.t9 a_6149_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_11033_943.t1 CLK VPB.t41 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_5101_1004.t3 D VPB.t36 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 a_343_383.t0 CLK VPB.t50 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 a_14869_1005.t2 a_8357_1004.t11 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 VNB a_5101_1004.t7 a_6603_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_9985_1004.t0 D VPB.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 a_13367_383.t5 SN VPB.t81 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_1265_943.t1 a_1905_1004.t9 VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 VPB.t9 a_3599_383.t9 a_3473_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 VNB a_3473_1004.t8 a_4013_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1103 VPB.t45 CLK a_10111_383.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_11673_1004.t5 SN VPB.t82 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 VPB.t44 CLK a_1265_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VPB.t90 a_6149_943.t12 a_5227_383.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 VPB.t55 a_13367_383.t9 a_13241_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 VNB a_11673_1004.t9 a_12470_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1109 a_8357_1004.t2 a_8483_383.t9 VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_3599_383.t3 a_3473_1004.t13 VPB.t54 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 VPB.t51 CLK a_6149_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1112 VPB.t61 a_13241_1004.t13 a_14869_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 VNB a_9985_1004.t6 a_10525_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1114 VNB a_13241_1004.t12 a_15430_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1115 a_343_383.t2 a_1265_943.t13 VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 VPB.t60 a_343_383.t12 a_3473_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_5227_383.t0 a_5101_1004.t10 VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_13367_383.t3 a_11033_943.t13 VPB.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 VPB.t80 SN a_8483_383.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 a_1265_943.t2 CLK VPB.t43 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 VPB.t74 SN a_1905_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 a_11673_1004.t0 a_9985_1004.t10 VPB.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 D VPB 0.24fF
C1 CLK VPB 3.26fF
C2 SN VPB 0.30fF
C3 D CLK 1.75fF
C4 D SN 3.39fF
C5 CLK SN 0.41fF
R0 a_6149_943.n6 a_6149_943.t6 454.685
R1 a_6149_943.n8 a_6149_943.t7 454.685
R2 a_6149_943.n4 a_6149_943.t9 454.685
R3 a_6149_943.n6 a_6149_943.t11 428.979
R4 a_6149_943.n8 a_6149_943.t12 428.979
R5 a_6149_943.n4 a_6149_943.t8 428.979
R6 a_6149_943.n7 a_6149_943.t5 248.006
R7 a_6149_943.n9 a_6149_943.t13 248.006
R8 a_6149_943.n5 a_6149_943.t10 248.006
R9 a_6149_943.n14 a_6149_943.n12 220.639
R10 a_6149_943.n12 a_6149_943.n3 135.994
R11 a_6149_943.n7 a_6149_943.n6 81.941
R12 a_6149_943.n9 a_6149_943.n8 81.941
R13 a_6149_943.n5 a_6149_943.n4 81.941
R14 a_6149_943.n11 a_6149_943.n5 81.396
R15 a_6149_943.n10 a_6149_943.n9 79.491
R16 a_6149_943.n3 a_6149_943.n2 76.002
R17 a_6149_943.n10 a_6149_943.n7 76
R18 a_6149_943.n12 a_6149_943.n11 76
R19 a_6149_943.n14 a_6149_943.n13 30
R20 a_6149_943.n15 a_6149_943.n0 24.383
R21 a_6149_943.n15 a_6149_943.n14 23.684
R22 a_6149_943.n1 a_6149_943.t2 14.282
R23 a_6149_943.n1 a_6149_943.t3 14.282
R24 a_6149_943.n2 a_6149_943.t0 14.282
R25 a_6149_943.n2 a_6149_943.t1 14.282
R26 a_6149_943.n3 a_6149_943.n1 12.85
R27 a_6149_943.n11 a_6149_943.n10 2.947
R28 a_6884_182.n12 a_6884_182.n10 82.852
R29 a_6884_182.t1 a_6884_182.n2 46.91
R30 a_6884_182.n7 a_6884_182.n5 34.805
R31 a_6884_182.n7 a_6884_182.n6 32.622
R32 a_6884_182.n10 a_6884_182.t1 32.416
R33 a_6884_182.n12 a_6884_182.n11 27.2
R34 a_6884_182.n13 a_6884_182.n0 23.498
R35 a_6884_182.n13 a_6884_182.n12 22.4
R36 a_6884_182.n9 a_6884_182.n7 19.017
R37 a_6884_182.n2 a_6884_182.n1 17.006
R38 a_6884_182.n5 a_6884_182.n4 7.5
R39 a_6884_182.n9 a_6884_182.n8 7.5
R40 a_6884_182.t1 a_6884_182.n3 7.04
R41 a_6884_182.n10 a_6884_182.n9 1.435
R42 a_6789_1004.n5 a_6789_1004.t9 480.392
R43 a_6789_1004.n5 a_6789_1004.t7 403.272
R44 a_6789_1004.n7 a_6789_1004.n4 233.952
R45 a_6789_1004.n6 a_6789_1004.t8 213.869
R46 a_6789_1004.n6 a_6789_1004.n5 161.6
R47 a_6789_1004.n7 a_6789_1004.n6 153.315
R48 a_6789_1004.n9 a_6789_1004.n7 150.014
R49 a_6789_1004.n3 a_6789_1004.n2 79.232
R50 a_6789_1004.n4 a_6789_1004.n3 63.152
R51 a_6789_1004.n4 a_6789_1004.n0 16.08
R52 a_6789_1004.n3 a_6789_1004.n1 16.08
R53 a_6789_1004.n9 a_6789_1004.n8 15.218
R54 a_6789_1004.n0 a_6789_1004.t4 14.282
R55 a_6789_1004.n0 a_6789_1004.t5 14.282
R56 a_6789_1004.n1 a_6789_1004.t2 14.282
R57 a_6789_1004.n1 a_6789_1004.t1 14.282
R58 a_6789_1004.n2 a_6789_1004.t3 14.282
R59 a_6789_1004.n2 a_6789_1004.t0 14.282
R60 a_6789_1004.n10 a_6789_1004.n9 12.014
R61 a_5227_383.n6 a_5227_383.t9 480.392
R62 a_5227_383.n8 a_5227_383.t7 472.359
R63 a_5227_383.n6 a_5227_383.t11 403.272
R64 a_5227_383.n8 a_5227_383.t10 384.527
R65 a_5227_383.n7 a_5227_383.t8 320.08
R66 a_5227_383.n9 a_5227_383.t12 277.772
R67 a_5227_383.n13 a_5227_383.n11 249.364
R68 a_5227_383.n11 a_5227_383.n5 127.401
R69 a_5227_383.n10 a_5227_383.n7 83.304
R70 a_5227_383.n10 a_5227_383.n9 80.032
R71 a_5227_383.n4 a_5227_383.n3 79.232
R72 a_5227_383.n11 a_5227_383.n10 76
R73 a_5227_383.n9 a_5227_383.n8 67.001
R74 a_5227_383.n5 a_5227_383.n4 63.152
R75 a_5227_383.n7 a_5227_383.n6 55.388
R76 a_5227_383.n13 a_5227_383.n12 30
R77 a_5227_383.n14 a_5227_383.n0 24.383
R78 a_5227_383.n14 a_5227_383.n13 23.684
R79 a_5227_383.n5 a_5227_383.n1 16.08
R80 a_5227_383.n4 a_5227_383.n2 16.08
R81 a_5227_383.n1 a_5227_383.t4 14.282
R82 a_5227_383.n1 a_5227_383.t5 14.282
R83 a_5227_383.n2 a_5227_383.t2 14.282
R84 a_5227_383.n2 a_5227_383.t1 14.282
R85 a_5227_383.n3 a_5227_383.t3 14.282
R86 a_5227_383.n3 a_5227_383.t0 14.282
R87 VPB VPB.n1501 126.832
R88 VPB.n39 VPB.n37 94.117
R89 VPB.n1428 VPB.n1426 94.117
R90 VPB.n1345 VPB.n1343 94.117
R91 VPB.n1282 VPB.n1280 94.117
R92 VPB.n1219 VPB.n1217 94.117
R93 VPB.n1136 VPB.n1134 94.117
R94 VPB.n1073 VPB.n1071 94.117
R95 VPB.n990 VPB.n988 94.117
R96 VPB.n907 VPB.n905 94.117
R97 VPB.n844 VPB.n842 94.117
R98 VPB.n781 VPB.n779 94.117
R99 VPB.n698 VPB.n696 94.117
R100 VPB.n635 VPB.n633 94.117
R101 VPB.n552 VPB.n550 94.117
R102 VPB.n469 VPB.n467 94.117
R103 VPB.n406 VPB.n404 94.117
R104 VPB.n343 VPB.n341 94.117
R105 VPB.n260 VPB.n258 94.117
R106 VPB.n197 VPB.n195 94.117
R107 VPB.n142 VPB.n140 94.117
R108 VPB.n273 VPB.n272 80.104
R109 VPB.n482 VPB.n481 80.104
R110 VPB.n565 VPB.n564 80.104
R111 VPB.n711 VPB.n710 80.104
R112 VPB.n920 VPB.n919 80.104
R113 VPB.n1003 VPB.n1002 80.104
R114 VPB.n1149 VPB.n1148 80.104
R115 VPB.n1358 VPB.n1357 80.104
R116 VPB.n1441 VPB.n1440 80.104
R117 VPB.n105 VPB.n104 76
R118 VPB.n109 VPB.n108 76
R119 VPB.n113 VPB.n112 76
R120 VPB.n117 VPB.n116 76
R121 VPB.n144 VPB.n143 76
R122 VPB.n148 VPB.n147 76
R123 VPB.n152 VPB.n151 76
R124 VPB.n156 VPB.n155 76
R125 VPB.n160 VPB.n159 76
R126 VPB.n164 VPB.n163 76
R127 VPB.n168 VPB.n167 76
R128 VPB.n172 VPB.n171 76
R129 VPB.n199 VPB.n198 76
R130 VPB.n204 VPB.n203 76
R131 VPB.n209 VPB.n208 76
R132 VPB.n216 VPB.n215 76
R133 VPB.n221 VPB.n220 76
R134 VPB.n226 VPB.n225 76
R135 VPB.n231 VPB.n230 76
R136 VPB.n235 VPB.n234 76
R137 VPB.n262 VPB.n261 76
R138 VPB.n266 VPB.n265 76
R139 VPB.n271 VPB.n270 76
R140 VPB.n276 VPB.n275 76
R141 VPB.n283 VPB.n282 76
R142 VPB.n288 VPB.n287 76
R143 VPB.n293 VPB.n292 76
R144 VPB.n300 VPB.n299 76
R145 VPB.n305 VPB.n304 76
R146 VPB.n310 VPB.n309 76
R147 VPB.n314 VPB.n313 76
R148 VPB.n318 VPB.n317 76
R149 VPB.n345 VPB.n344 76
R150 VPB.n350 VPB.n349 76
R151 VPB.n355 VPB.n354 76
R152 VPB.n362 VPB.n361 76
R153 VPB.n367 VPB.n366 76
R154 VPB.n372 VPB.n371 76
R155 VPB.n377 VPB.n376 76
R156 VPB.n381 VPB.n380 76
R157 VPB.n408 VPB.n407 76
R158 VPB.n413 VPB.n412 76
R159 VPB.n418 VPB.n417 76
R160 VPB.n425 VPB.n424 76
R161 VPB.n430 VPB.n429 76
R162 VPB.n435 VPB.n434 76
R163 VPB.n440 VPB.n439 76
R164 VPB.n444 VPB.n443 76
R165 VPB.n471 VPB.n470 76
R166 VPB.n475 VPB.n474 76
R167 VPB.n480 VPB.n479 76
R168 VPB.n485 VPB.n484 76
R169 VPB.n492 VPB.n491 76
R170 VPB.n497 VPB.n496 76
R171 VPB.n502 VPB.n501 76
R172 VPB.n509 VPB.n508 76
R173 VPB.n514 VPB.n513 76
R174 VPB.n519 VPB.n518 76
R175 VPB.n523 VPB.n522 76
R176 VPB.n527 VPB.n526 76
R177 VPB.n554 VPB.n553 76
R178 VPB.n558 VPB.n557 76
R179 VPB.n563 VPB.n562 76
R180 VPB.n568 VPB.n567 76
R181 VPB.n575 VPB.n574 76
R182 VPB.n580 VPB.n579 76
R183 VPB.n585 VPB.n584 76
R184 VPB.n592 VPB.n591 76
R185 VPB.n597 VPB.n596 76
R186 VPB.n602 VPB.n601 76
R187 VPB.n606 VPB.n605 76
R188 VPB.n610 VPB.n609 76
R189 VPB.n637 VPB.n636 76
R190 VPB.n642 VPB.n641 76
R191 VPB.n647 VPB.n646 76
R192 VPB.n654 VPB.n653 76
R193 VPB.n659 VPB.n658 76
R194 VPB.n664 VPB.n663 76
R195 VPB.n669 VPB.n668 76
R196 VPB.n673 VPB.n672 76
R197 VPB.n700 VPB.n699 76
R198 VPB.n704 VPB.n703 76
R199 VPB.n709 VPB.n708 76
R200 VPB.n714 VPB.n713 76
R201 VPB.n721 VPB.n720 76
R202 VPB.n726 VPB.n725 76
R203 VPB.n731 VPB.n730 76
R204 VPB.n738 VPB.n737 76
R205 VPB.n743 VPB.n742 76
R206 VPB.n748 VPB.n747 76
R207 VPB.n752 VPB.n751 76
R208 VPB.n756 VPB.n755 76
R209 VPB.n783 VPB.n782 76
R210 VPB.n788 VPB.n787 76
R211 VPB.n793 VPB.n792 76
R212 VPB.n800 VPB.n799 76
R213 VPB.n805 VPB.n804 76
R214 VPB.n810 VPB.n809 76
R215 VPB.n815 VPB.n814 76
R216 VPB.n819 VPB.n818 76
R217 VPB.n846 VPB.n845 76
R218 VPB.n851 VPB.n850 76
R219 VPB.n856 VPB.n855 76
R220 VPB.n863 VPB.n862 76
R221 VPB.n868 VPB.n867 76
R222 VPB.n873 VPB.n872 76
R223 VPB.n878 VPB.n877 76
R224 VPB.n882 VPB.n881 76
R225 VPB.n909 VPB.n908 76
R226 VPB.n913 VPB.n912 76
R227 VPB.n918 VPB.n917 76
R228 VPB.n923 VPB.n922 76
R229 VPB.n930 VPB.n929 76
R230 VPB.n935 VPB.n934 76
R231 VPB.n940 VPB.n939 76
R232 VPB.n947 VPB.n946 76
R233 VPB.n952 VPB.n951 76
R234 VPB.n957 VPB.n956 76
R235 VPB.n961 VPB.n960 76
R236 VPB.n965 VPB.n964 76
R237 VPB.n992 VPB.n991 76
R238 VPB.n996 VPB.n995 76
R239 VPB.n1001 VPB.n1000 76
R240 VPB.n1006 VPB.n1005 76
R241 VPB.n1013 VPB.n1012 76
R242 VPB.n1018 VPB.n1017 76
R243 VPB.n1023 VPB.n1022 76
R244 VPB.n1030 VPB.n1029 76
R245 VPB.n1035 VPB.n1034 76
R246 VPB.n1040 VPB.n1039 76
R247 VPB.n1044 VPB.n1043 76
R248 VPB.n1048 VPB.n1047 76
R249 VPB.n1075 VPB.n1074 76
R250 VPB.n1080 VPB.n1079 76
R251 VPB.n1085 VPB.n1084 76
R252 VPB.n1092 VPB.n1091 76
R253 VPB.n1097 VPB.n1096 76
R254 VPB.n1102 VPB.n1101 76
R255 VPB.n1107 VPB.n1106 76
R256 VPB.n1111 VPB.n1110 76
R257 VPB.n1138 VPB.n1137 76
R258 VPB.n1142 VPB.n1141 76
R259 VPB.n1147 VPB.n1146 76
R260 VPB.n1152 VPB.n1151 76
R261 VPB.n1159 VPB.n1158 76
R262 VPB.n1164 VPB.n1163 76
R263 VPB.n1169 VPB.n1168 76
R264 VPB.n1176 VPB.n1175 76
R265 VPB.n1181 VPB.n1180 76
R266 VPB.n1186 VPB.n1185 76
R267 VPB.n1190 VPB.n1189 76
R268 VPB.n1194 VPB.n1193 76
R269 VPB.n1221 VPB.n1220 76
R270 VPB.n1226 VPB.n1225 76
R271 VPB.n1231 VPB.n1230 76
R272 VPB.n1238 VPB.n1237 76
R273 VPB.n1243 VPB.n1242 76
R274 VPB.n1248 VPB.n1247 76
R275 VPB.n1253 VPB.n1252 76
R276 VPB.n1257 VPB.n1256 76
R277 VPB.n1284 VPB.n1283 76
R278 VPB.n1289 VPB.n1288 76
R279 VPB.n1294 VPB.n1293 76
R280 VPB.n1301 VPB.n1300 76
R281 VPB.n1306 VPB.n1305 76
R282 VPB.n1311 VPB.n1310 76
R283 VPB.n1316 VPB.n1315 76
R284 VPB.n1320 VPB.n1319 76
R285 VPB.n1347 VPB.n1346 76
R286 VPB.n1351 VPB.n1350 76
R287 VPB.n1356 VPB.n1355 76
R288 VPB.n1361 VPB.n1360 76
R289 VPB.n1368 VPB.n1367 76
R290 VPB.n1373 VPB.n1372 76
R291 VPB.n1378 VPB.n1377 76
R292 VPB.n1385 VPB.n1384 76
R293 VPB.n1390 VPB.n1389 76
R294 VPB.n1395 VPB.n1394 76
R295 VPB.n1399 VPB.n1398 76
R296 VPB.n1403 VPB.n1402 76
R297 VPB.n1430 VPB.n1429 76
R298 VPB.n1434 VPB.n1433 76
R299 VPB.n1439 VPB.n1438 76
R300 VPB.n1444 VPB.n1443 76
R301 VPB.n1451 VPB.n1450 76
R302 VPB.n1456 VPB.n1455 76
R303 VPB.n1461 VPB.n1460 76
R304 VPB.n1468 VPB.n1467 76
R305 VPB.n1473 VPB.n1472 76
R306 VPB.n1478 VPB.n1477 76
R307 VPB.n1482 VPB.n1481 76
R308 VPB.n1486 VPB.n1485 76
R309 VPB.n302 VPB.n301 75.654
R310 VPB.n511 VPB.n510 75.654
R311 VPB.n594 VPB.n593 75.654
R312 VPB.n740 VPB.n739 75.654
R313 VPB.n949 VPB.n948 75.654
R314 VPB.n1032 VPB.n1031 75.654
R315 VPB.n1178 VPB.n1177 75.654
R316 VPB.n1387 VPB.n1386 75.654
R317 VPB.n1470 VPB.n1469 75.654
R318 VPB.n21 VPB.n20 61.764
R319 VPB.n1410 VPB.n1409 61.764
R320 VPB.n1327 VPB.n1326 61.764
R321 VPB.n1264 VPB.n1263 61.764
R322 VPB.n1201 VPB.n1200 61.764
R323 VPB.n1118 VPB.n1117 61.764
R324 VPB.n1055 VPB.n1054 61.764
R325 VPB.n972 VPB.n971 61.764
R326 VPB.n889 VPB.n888 61.764
R327 VPB.n826 VPB.n825 61.764
R328 VPB.n763 VPB.n762 61.764
R329 VPB.n680 VPB.n679 61.764
R330 VPB.n617 VPB.n616 61.764
R331 VPB.n534 VPB.n533 61.764
R332 VPB.n451 VPB.n450 61.764
R333 VPB.n388 VPB.n387 61.764
R334 VPB.n325 VPB.n324 61.764
R335 VPB.n242 VPB.n241 61.764
R336 VPB.n179 VPB.n178 61.764
R337 VPB.n124 VPB.n123 61.764
R338 VPB.n227 VPB.t53 55.465
R339 VPB.n200 VPB.t26 55.465
R340 VPB.n62 VPB.t38 55.106
R341 VPB.n1474 VPB.t71 55.106
R342 VPB.n1391 VPB.t14 55.106
R343 VPB.n1312 VPB.t11 55.106
R344 VPB.n1249 VPB.t86 55.106
R345 VPB.n1182 VPB.t54 55.106
R346 VPB.n1103 VPB.t36 55.106
R347 VPB.n1036 VPB.t2 55.106
R348 VPB.n953 VPB.t66 55.106
R349 VPB.n874 VPB.t28 55.106
R350 VPB.n811 VPB.t32 55.106
R351 VPB.n744 VPB.t7 55.106
R352 VPB.n665 VPB.t35 55.106
R353 VPB.n598 VPB.t6 55.106
R354 VPB.n515 VPB.t25 55.106
R355 VPB.n436 VPB.t56 55.106
R356 VPB.n373 VPB.t23 55.106
R357 VPB.n306 VPB.t57 55.106
R358 VPB.n44 VPB.t59 55.106
R359 VPB.n1435 VPB.t0 55.106
R360 VPB.n1352 VPB.t4 55.106
R361 VPB.n1285 VPB.t44 55.106
R362 VPB.n1222 VPB.t9 55.106
R363 VPB.n1143 VPB.t3 55.106
R364 VPB.n1076 VPB.t30 55.106
R365 VPB.n997 VPB.t90 55.106
R366 VPB.n914 VPB.t88 55.106
R367 VPB.n847 VPB.t51 55.106
R368 VPB.n784 VPB.t8 55.106
R369 VPB.n705 VPB.t92 55.106
R370 VPB.n638 VPB.t15 55.106
R371 VPB.n559 VPB.t64 55.106
R372 VPB.n476 VPB.t13 55.106
R373 VPB.n409 VPB.t42 55.106
R374 VPB.n346 VPB.t55 55.106
R375 VPB.n267 VPB.t16 55.106
R376 VPB.n206 VPB.n205 48.952
R377 VPB.n280 VPB.n279 48.952
R378 VPB.n352 VPB.n351 48.952
R379 VPB.n415 VPB.n414 48.952
R380 VPB.n489 VPB.n488 48.952
R381 VPB.n572 VPB.n571 48.952
R382 VPB.n644 VPB.n643 48.952
R383 VPB.n718 VPB.n717 48.952
R384 VPB.n790 VPB.n789 48.952
R385 VPB.n853 VPB.n852 48.952
R386 VPB.n927 VPB.n926 48.952
R387 VPB.n1010 VPB.n1009 48.952
R388 VPB.n1082 VPB.n1081 48.952
R389 VPB.n1156 VPB.n1155 48.952
R390 VPB.n1228 VPB.n1227 48.952
R391 VPB.n1291 VPB.n1290 48.952
R392 VPB.n1365 VPB.n1364 48.952
R393 VPB.n1448 VPB.n1447 48.952
R394 VPB.n46 VPB.n45 48.952
R395 VPB.n223 VPB.n222 44.502
R396 VPB.n297 VPB.n296 44.502
R397 VPB.n369 VPB.n368 44.502
R398 VPB.n432 VPB.n431 44.502
R399 VPB.n506 VPB.n505 44.502
R400 VPB.n589 VPB.n588 44.502
R401 VPB.n661 VPB.n660 44.502
R402 VPB.n735 VPB.n734 44.502
R403 VPB.n807 VPB.n806 44.502
R404 VPB.n870 VPB.n869 44.502
R405 VPB.n944 VPB.n943 44.502
R406 VPB.n1027 VPB.n1026 44.502
R407 VPB.n1099 VPB.n1098 44.502
R408 VPB.n1173 VPB.n1172 44.502
R409 VPB.n1245 VPB.n1244 44.502
R410 VPB.n1308 VPB.n1307 44.502
R411 VPB.n1382 VPB.n1381 44.502
R412 VPB.n1465 VPB.n1464 44.502
R413 VPB.n59 VPB.n58 44.502
R414 VPB.n211 VPB.n210 41.183
R415 VPB.n53 VPB.n14 40.824
R416 VPB.n1463 VPB.n1462 40.824
R417 VPB.n1446 VPB.n1445 40.824
R418 VPB.n1380 VPB.n1379 40.824
R419 VPB.n1363 VPB.n1362 40.824
R420 VPB.n1296 VPB.n1295 40.824
R421 VPB.n1233 VPB.n1232 40.824
R422 VPB.n1171 VPB.n1170 40.824
R423 VPB.n1154 VPB.n1153 40.824
R424 VPB.n1087 VPB.n1086 40.824
R425 VPB.n1025 VPB.n1024 40.824
R426 VPB.n1008 VPB.n1007 40.824
R427 VPB.n942 VPB.n941 40.824
R428 VPB.n925 VPB.n924 40.824
R429 VPB.n858 VPB.n857 40.824
R430 VPB.n795 VPB.n794 40.824
R431 VPB.n733 VPB.n732 40.824
R432 VPB.n716 VPB.n715 40.824
R433 VPB.n649 VPB.n648 40.824
R434 VPB.n587 VPB.n586 40.824
R435 VPB.n570 VPB.n569 40.824
R436 VPB.n504 VPB.n503 40.824
R437 VPB.n487 VPB.n486 40.824
R438 VPB.n420 VPB.n419 40.824
R439 VPB.n357 VPB.n356 40.824
R440 VPB.n295 VPB.n294 40.824
R441 VPB.n278 VPB.n277 40.824
R442 VPB.n100 VPB.n99 35.118
R443 VPB.n1493 VPB.n1492 35.118
R444 VPB.n1498 VPB.n1494 20.452
R445 VPB.n89 VPB.n86 20.452
R446 VPB.n213 VPB.n212 17.801
R447 VPB.n285 VPB.n284 17.801
R448 VPB.n359 VPB.n358 17.801
R449 VPB.n422 VPB.n421 17.801
R450 VPB.n494 VPB.n493 17.801
R451 VPB.n577 VPB.n576 17.801
R452 VPB.n651 VPB.n650 17.801
R453 VPB.n723 VPB.n722 17.801
R454 VPB.n797 VPB.n796 17.801
R455 VPB.n860 VPB.n859 17.801
R456 VPB.n932 VPB.n931 17.801
R457 VPB.n1015 VPB.n1014 17.801
R458 VPB.n1089 VPB.n1088 17.801
R459 VPB.n1161 VPB.n1160 17.801
R460 VPB.n1235 VPB.n1234 17.801
R461 VPB.n1298 VPB.n1297 17.801
R462 VPB.n1370 VPB.n1369 17.801
R463 VPB.n1453 VPB.n1452 17.801
R464 VPB.n50 VPB.n49 17.801
R465 VPB.n14 VPB.t62 14.282
R466 VPB.n14 VPB.t39 14.282
R467 VPB.n1462 VPB.t50 14.282
R468 VPB.n1462 VPB.t68 14.282
R469 VPB.n1445 VPB.t20 14.282
R470 VPB.n1445 VPB.t49 14.282
R471 VPB.n1379 VPB.t75 14.282
R472 VPB.n1379 VPB.t67 14.282
R473 VPB.n1362 VPB.t22 14.282
R474 VPB.n1362 VPB.t74 14.282
R475 VPB.n1295 VPB.t43 14.282
R476 VPB.n1295 VPB.t5 14.282
R477 VPB.n1232 VPB.t29 14.282
R478 VPB.n1232 VPB.t60 14.282
R479 VPB.n1170 VPB.t73 14.282
R480 VPB.n1170 VPB.t58 14.282
R481 VPB.n1153 VPB.t21 14.282
R482 VPB.n1153 VPB.t76 14.282
R483 VPB.n1086 VPB.t31 14.282
R484 VPB.n1086 VPB.t37 14.282
R485 VPB.n1024 VPB.t47 14.282
R486 VPB.n1024 VPB.t65 14.282
R487 VPB.n1007 VPB.t91 14.282
R488 VPB.n1007 VPB.t48 14.282
R489 VPB.n941 VPB.t77 14.282
R490 VPB.n941 VPB.t85 14.282
R491 VPB.n924 VPB.t89 14.282
R492 VPB.n924 VPB.t78 14.282
R493 VPB.n857 VPB.t52 14.282
R494 VPB.n857 VPB.t27 14.282
R495 VPB.n794 VPB.t17 14.282
R496 VPB.n794 VPB.t33 14.282
R497 VPB.n732 VPB.t84 14.282
R498 VPB.n732 VPB.t1 14.282
R499 VPB.n715 VPB.t87 14.282
R500 VPB.n715 VPB.t80 14.282
R501 VPB.n648 VPB.t72 14.282
R502 VPB.n648 VPB.t34 14.282
R503 VPB.n586 VPB.t46 14.282
R504 VPB.n586 VPB.t24 14.282
R505 VPB.n569 VPB.t70 14.282
R506 VPB.n569 VPB.t45 14.282
R507 VPB.n503 VPB.t82 14.282
R508 VPB.n503 VPB.t10 14.282
R509 VPB.n486 VPB.t18 14.282
R510 VPB.n486 VPB.t79 14.282
R511 VPB.n419 VPB.t41 14.282
R512 VPB.n419 VPB.t93 14.282
R513 VPB.n356 VPB.t63 14.282
R514 VPB.n356 VPB.t69 14.282
R515 VPB.n294 VPB.t81 14.282
R516 VPB.n294 VPB.t40 14.282
R517 VPB.n277 VPB.t19 14.282
R518 VPB.n277 VPB.t83 14.282
R519 VPB.n210 VPB.t12 14.282
R520 VPB.n210 VPB.t61 14.282
R521 VPB.n89 VPB.n88 13.653
R522 VPB.n88 VPB.n87 13.653
R523 VPB.n98 VPB.n97 13.653
R524 VPB.n97 VPB.n96 13.653
R525 VPB.n95 VPB.n94 13.653
R526 VPB.n94 VPB.n93 13.653
R527 VPB.n92 VPB.n91 13.653
R528 VPB.n91 VPB.n90 13.653
R529 VPB.n104 VPB.n103 13.653
R530 VPB.n103 VPB.n102 13.653
R531 VPB.n108 VPB.n107 13.653
R532 VPB.n107 VPB.n106 13.653
R533 VPB.n112 VPB.n111 13.653
R534 VPB.n111 VPB.n110 13.653
R535 VPB.n116 VPB.n115 13.653
R536 VPB.n115 VPB.n114 13.653
R537 VPB.n143 VPB.n142 13.653
R538 VPB.n142 VPB.n141 13.653
R539 VPB.n147 VPB.n146 13.653
R540 VPB.n146 VPB.n145 13.653
R541 VPB.n151 VPB.n150 13.653
R542 VPB.n150 VPB.n149 13.653
R543 VPB.n155 VPB.n154 13.653
R544 VPB.n154 VPB.n153 13.653
R545 VPB.n159 VPB.n158 13.653
R546 VPB.n158 VPB.n157 13.653
R547 VPB.n163 VPB.n162 13.653
R548 VPB.n162 VPB.n161 13.653
R549 VPB.n167 VPB.n166 13.653
R550 VPB.n166 VPB.n165 13.653
R551 VPB.n171 VPB.n170 13.653
R552 VPB.n170 VPB.n169 13.653
R553 VPB.n198 VPB.n197 13.653
R554 VPB.n197 VPB.n196 13.653
R555 VPB.n203 VPB.n202 13.653
R556 VPB.n202 VPB.n201 13.653
R557 VPB.n208 VPB.n207 13.653
R558 VPB.n207 VPB.n206 13.653
R559 VPB.n215 VPB.n214 13.653
R560 VPB.n214 VPB.n213 13.653
R561 VPB.n220 VPB.n219 13.653
R562 VPB.n219 VPB.n218 13.653
R563 VPB.n225 VPB.n224 13.653
R564 VPB.n224 VPB.n223 13.653
R565 VPB.n230 VPB.n229 13.653
R566 VPB.n229 VPB.n228 13.653
R567 VPB.n234 VPB.n233 13.653
R568 VPB.n233 VPB.n232 13.653
R569 VPB.n261 VPB.n260 13.653
R570 VPB.n260 VPB.n259 13.653
R571 VPB.n265 VPB.n264 13.653
R572 VPB.n264 VPB.n263 13.653
R573 VPB.n270 VPB.n269 13.653
R574 VPB.n269 VPB.n268 13.653
R575 VPB.n275 VPB.n274 13.653
R576 VPB.n274 VPB.n273 13.653
R577 VPB.n282 VPB.n281 13.653
R578 VPB.n281 VPB.n280 13.653
R579 VPB.n287 VPB.n286 13.653
R580 VPB.n286 VPB.n285 13.653
R581 VPB.n292 VPB.n291 13.653
R582 VPB.n291 VPB.n290 13.653
R583 VPB.n299 VPB.n298 13.653
R584 VPB.n298 VPB.n297 13.653
R585 VPB.n304 VPB.n303 13.653
R586 VPB.n303 VPB.n302 13.653
R587 VPB.n309 VPB.n308 13.653
R588 VPB.n308 VPB.n307 13.653
R589 VPB.n313 VPB.n312 13.653
R590 VPB.n312 VPB.n311 13.653
R591 VPB.n317 VPB.n316 13.653
R592 VPB.n316 VPB.n315 13.653
R593 VPB.n344 VPB.n343 13.653
R594 VPB.n343 VPB.n342 13.653
R595 VPB.n349 VPB.n348 13.653
R596 VPB.n348 VPB.n347 13.653
R597 VPB.n354 VPB.n353 13.653
R598 VPB.n353 VPB.n352 13.653
R599 VPB.n361 VPB.n360 13.653
R600 VPB.n360 VPB.n359 13.653
R601 VPB.n366 VPB.n365 13.653
R602 VPB.n365 VPB.n364 13.653
R603 VPB.n371 VPB.n370 13.653
R604 VPB.n370 VPB.n369 13.653
R605 VPB.n376 VPB.n375 13.653
R606 VPB.n375 VPB.n374 13.653
R607 VPB.n380 VPB.n379 13.653
R608 VPB.n379 VPB.n378 13.653
R609 VPB.n407 VPB.n406 13.653
R610 VPB.n406 VPB.n405 13.653
R611 VPB.n412 VPB.n411 13.653
R612 VPB.n411 VPB.n410 13.653
R613 VPB.n417 VPB.n416 13.653
R614 VPB.n416 VPB.n415 13.653
R615 VPB.n424 VPB.n423 13.653
R616 VPB.n423 VPB.n422 13.653
R617 VPB.n429 VPB.n428 13.653
R618 VPB.n428 VPB.n427 13.653
R619 VPB.n434 VPB.n433 13.653
R620 VPB.n433 VPB.n432 13.653
R621 VPB.n439 VPB.n438 13.653
R622 VPB.n438 VPB.n437 13.653
R623 VPB.n443 VPB.n442 13.653
R624 VPB.n442 VPB.n441 13.653
R625 VPB.n470 VPB.n469 13.653
R626 VPB.n469 VPB.n468 13.653
R627 VPB.n474 VPB.n473 13.653
R628 VPB.n473 VPB.n472 13.653
R629 VPB.n479 VPB.n478 13.653
R630 VPB.n478 VPB.n477 13.653
R631 VPB.n484 VPB.n483 13.653
R632 VPB.n483 VPB.n482 13.653
R633 VPB.n491 VPB.n490 13.653
R634 VPB.n490 VPB.n489 13.653
R635 VPB.n496 VPB.n495 13.653
R636 VPB.n495 VPB.n494 13.653
R637 VPB.n501 VPB.n500 13.653
R638 VPB.n500 VPB.n499 13.653
R639 VPB.n508 VPB.n507 13.653
R640 VPB.n507 VPB.n506 13.653
R641 VPB.n513 VPB.n512 13.653
R642 VPB.n512 VPB.n511 13.653
R643 VPB.n518 VPB.n517 13.653
R644 VPB.n517 VPB.n516 13.653
R645 VPB.n522 VPB.n521 13.653
R646 VPB.n521 VPB.n520 13.653
R647 VPB.n526 VPB.n525 13.653
R648 VPB.n525 VPB.n524 13.653
R649 VPB.n553 VPB.n552 13.653
R650 VPB.n552 VPB.n551 13.653
R651 VPB.n557 VPB.n556 13.653
R652 VPB.n556 VPB.n555 13.653
R653 VPB.n562 VPB.n561 13.653
R654 VPB.n561 VPB.n560 13.653
R655 VPB.n567 VPB.n566 13.653
R656 VPB.n566 VPB.n565 13.653
R657 VPB.n574 VPB.n573 13.653
R658 VPB.n573 VPB.n572 13.653
R659 VPB.n579 VPB.n578 13.653
R660 VPB.n578 VPB.n577 13.653
R661 VPB.n584 VPB.n583 13.653
R662 VPB.n583 VPB.n582 13.653
R663 VPB.n591 VPB.n590 13.653
R664 VPB.n590 VPB.n589 13.653
R665 VPB.n596 VPB.n595 13.653
R666 VPB.n595 VPB.n594 13.653
R667 VPB.n601 VPB.n600 13.653
R668 VPB.n600 VPB.n599 13.653
R669 VPB.n605 VPB.n604 13.653
R670 VPB.n604 VPB.n603 13.653
R671 VPB.n609 VPB.n608 13.653
R672 VPB.n608 VPB.n607 13.653
R673 VPB.n636 VPB.n635 13.653
R674 VPB.n635 VPB.n634 13.653
R675 VPB.n641 VPB.n640 13.653
R676 VPB.n640 VPB.n639 13.653
R677 VPB.n646 VPB.n645 13.653
R678 VPB.n645 VPB.n644 13.653
R679 VPB.n653 VPB.n652 13.653
R680 VPB.n652 VPB.n651 13.653
R681 VPB.n658 VPB.n657 13.653
R682 VPB.n657 VPB.n656 13.653
R683 VPB.n663 VPB.n662 13.653
R684 VPB.n662 VPB.n661 13.653
R685 VPB.n668 VPB.n667 13.653
R686 VPB.n667 VPB.n666 13.653
R687 VPB.n672 VPB.n671 13.653
R688 VPB.n671 VPB.n670 13.653
R689 VPB.n699 VPB.n698 13.653
R690 VPB.n698 VPB.n697 13.653
R691 VPB.n703 VPB.n702 13.653
R692 VPB.n702 VPB.n701 13.653
R693 VPB.n708 VPB.n707 13.653
R694 VPB.n707 VPB.n706 13.653
R695 VPB.n713 VPB.n712 13.653
R696 VPB.n712 VPB.n711 13.653
R697 VPB.n720 VPB.n719 13.653
R698 VPB.n719 VPB.n718 13.653
R699 VPB.n725 VPB.n724 13.653
R700 VPB.n724 VPB.n723 13.653
R701 VPB.n730 VPB.n729 13.653
R702 VPB.n729 VPB.n728 13.653
R703 VPB.n737 VPB.n736 13.653
R704 VPB.n736 VPB.n735 13.653
R705 VPB.n742 VPB.n741 13.653
R706 VPB.n741 VPB.n740 13.653
R707 VPB.n747 VPB.n746 13.653
R708 VPB.n746 VPB.n745 13.653
R709 VPB.n751 VPB.n750 13.653
R710 VPB.n750 VPB.n749 13.653
R711 VPB.n755 VPB.n754 13.653
R712 VPB.n754 VPB.n753 13.653
R713 VPB.n782 VPB.n781 13.653
R714 VPB.n781 VPB.n780 13.653
R715 VPB.n787 VPB.n786 13.653
R716 VPB.n786 VPB.n785 13.653
R717 VPB.n792 VPB.n791 13.653
R718 VPB.n791 VPB.n790 13.653
R719 VPB.n799 VPB.n798 13.653
R720 VPB.n798 VPB.n797 13.653
R721 VPB.n804 VPB.n803 13.653
R722 VPB.n803 VPB.n802 13.653
R723 VPB.n809 VPB.n808 13.653
R724 VPB.n808 VPB.n807 13.653
R725 VPB.n814 VPB.n813 13.653
R726 VPB.n813 VPB.n812 13.653
R727 VPB.n818 VPB.n817 13.653
R728 VPB.n817 VPB.n816 13.653
R729 VPB.n845 VPB.n844 13.653
R730 VPB.n844 VPB.n843 13.653
R731 VPB.n850 VPB.n849 13.653
R732 VPB.n849 VPB.n848 13.653
R733 VPB.n855 VPB.n854 13.653
R734 VPB.n854 VPB.n853 13.653
R735 VPB.n862 VPB.n861 13.653
R736 VPB.n861 VPB.n860 13.653
R737 VPB.n867 VPB.n866 13.653
R738 VPB.n866 VPB.n865 13.653
R739 VPB.n872 VPB.n871 13.653
R740 VPB.n871 VPB.n870 13.653
R741 VPB.n877 VPB.n876 13.653
R742 VPB.n876 VPB.n875 13.653
R743 VPB.n881 VPB.n880 13.653
R744 VPB.n880 VPB.n879 13.653
R745 VPB.n908 VPB.n907 13.653
R746 VPB.n907 VPB.n906 13.653
R747 VPB.n912 VPB.n911 13.653
R748 VPB.n911 VPB.n910 13.653
R749 VPB.n917 VPB.n916 13.653
R750 VPB.n916 VPB.n915 13.653
R751 VPB.n922 VPB.n921 13.653
R752 VPB.n921 VPB.n920 13.653
R753 VPB.n929 VPB.n928 13.653
R754 VPB.n928 VPB.n927 13.653
R755 VPB.n934 VPB.n933 13.653
R756 VPB.n933 VPB.n932 13.653
R757 VPB.n939 VPB.n938 13.653
R758 VPB.n938 VPB.n937 13.653
R759 VPB.n946 VPB.n945 13.653
R760 VPB.n945 VPB.n944 13.653
R761 VPB.n951 VPB.n950 13.653
R762 VPB.n950 VPB.n949 13.653
R763 VPB.n956 VPB.n955 13.653
R764 VPB.n955 VPB.n954 13.653
R765 VPB.n960 VPB.n959 13.653
R766 VPB.n959 VPB.n958 13.653
R767 VPB.n964 VPB.n963 13.653
R768 VPB.n963 VPB.n962 13.653
R769 VPB.n991 VPB.n990 13.653
R770 VPB.n990 VPB.n989 13.653
R771 VPB.n995 VPB.n994 13.653
R772 VPB.n994 VPB.n993 13.653
R773 VPB.n1000 VPB.n999 13.653
R774 VPB.n999 VPB.n998 13.653
R775 VPB.n1005 VPB.n1004 13.653
R776 VPB.n1004 VPB.n1003 13.653
R777 VPB.n1012 VPB.n1011 13.653
R778 VPB.n1011 VPB.n1010 13.653
R779 VPB.n1017 VPB.n1016 13.653
R780 VPB.n1016 VPB.n1015 13.653
R781 VPB.n1022 VPB.n1021 13.653
R782 VPB.n1021 VPB.n1020 13.653
R783 VPB.n1029 VPB.n1028 13.653
R784 VPB.n1028 VPB.n1027 13.653
R785 VPB.n1034 VPB.n1033 13.653
R786 VPB.n1033 VPB.n1032 13.653
R787 VPB.n1039 VPB.n1038 13.653
R788 VPB.n1038 VPB.n1037 13.653
R789 VPB.n1043 VPB.n1042 13.653
R790 VPB.n1042 VPB.n1041 13.653
R791 VPB.n1047 VPB.n1046 13.653
R792 VPB.n1046 VPB.n1045 13.653
R793 VPB.n1074 VPB.n1073 13.653
R794 VPB.n1073 VPB.n1072 13.653
R795 VPB.n1079 VPB.n1078 13.653
R796 VPB.n1078 VPB.n1077 13.653
R797 VPB.n1084 VPB.n1083 13.653
R798 VPB.n1083 VPB.n1082 13.653
R799 VPB.n1091 VPB.n1090 13.653
R800 VPB.n1090 VPB.n1089 13.653
R801 VPB.n1096 VPB.n1095 13.653
R802 VPB.n1095 VPB.n1094 13.653
R803 VPB.n1101 VPB.n1100 13.653
R804 VPB.n1100 VPB.n1099 13.653
R805 VPB.n1106 VPB.n1105 13.653
R806 VPB.n1105 VPB.n1104 13.653
R807 VPB.n1110 VPB.n1109 13.653
R808 VPB.n1109 VPB.n1108 13.653
R809 VPB.n1137 VPB.n1136 13.653
R810 VPB.n1136 VPB.n1135 13.653
R811 VPB.n1141 VPB.n1140 13.653
R812 VPB.n1140 VPB.n1139 13.653
R813 VPB.n1146 VPB.n1145 13.653
R814 VPB.n1145 VPB.n1144 13.653
R815 VPB.n1151 VPB.n1150 13.653
R816 VPB.n1150 VPB.n1149 13.653
R817 VPB.n1158 VPB.n1157 13.653
R818 VPB.n1157 VPB.n1156 13.653
R819 VPB.n1163 VPB.n1162 13.653
R820 VPB.n1162 VPB.n1161 13.653
R821 VPB.n1168 VPB.n1167 13.653
R822 VPB.n1167 VPB.n1166 13.653
R823 VPB.n1175 VPB.n1174 13.653
R824 VPB.n1174 VPB.n1173 13.653
R825 VPB.n1180 VPB.n1179 13.653
R826 VPB.n1179 VPB.n1178 13.653
R827 VPB.n1185 VPB.n1184 13.653
R828 VPB.n1184 VPB.n1183 13.653
R829 VPB.n1189 VPB.n1188 13.653
R830 VPB.n1188 VPB.n1187 13.653
R831 VPB.n1193 VPB.n1192 13.653
R832 VPB.n1192 VPB.n1191 13.653
R833 VPB.n1220 VPB.n1219 13.653
R834 VPB.n1219 VPB.n1218 13.653
R835 VPB.n1225 VPB.n1224 13.653
R836 VPB.n1224 VPB.n1223 13.653
R837 VPB.n1230 VPB.n1229 13.653
R838 VPB.n1229 VPB.n1228 13.653
R839 VPB.n1237 VPB.n1236 13.653
R840 VPB.n1236 VPB.n1235 13.653
R841 VPB.n1242 VPB.n1241 13.653
R842 VPB.n1241 VPB.n1240 13.653
R843 VPB.n1247 VPB.n1246 13.653
R844 VPB.n1246 VPB.n1245 13.653
R845 VPB.n1252 VPB.n1251 13.653
R846 VPB.n1251 VPB.n1250 13.653
R847 VPB.n1256 VPB.n1255 13.653
R848 VPB.n1255 VPB.n1254 13.653
R849 VPB.n1283 VPB.n1282 13.653
R850 VPB.n1282 VPB.n1281 13.653
R851 VPB.n1288 VPB.n1287 13.653
R852 VPB.n1287 VPB.n1286 13.653
R853 VPB.n1293 VPB.n1292 13.653
R854 VPB.n1292 VPB.n1291 13.653
R855 VPB.n1300 VPB.n1299 13.653
R856 VPB.n1299 VPB.n1298 13.653
R857 VPB.n1305 VPB.n1304 13.653
R858 VPB.n1304 VPB.n1303 13.653
R859 VPB.n1310 VPB.n1309 13.653
R860 VPB.n1309 VPB.n1308 13.653
R861 VPB.n1315 VPB.n1314 13.653
R862 VPB.n1314 VPB.n1313 13.653
R863 VPB.n1319 VPB.n1318 13.653
R864 VPB.n1318 VPB.n1317 13.653
R865 VPB.n1346 VPB.n1345 13.653
R866 VPB.n1345 VPB.n1344 13.653
R867 VPB.n1350 VPB.n1349 13.653
R868 VPB.n1349 VPB.n1348 13.653
R869 VPB.n1355 VPB.n1354 13.653
R870 VPB.n1354 VPB.n1353 13.653
R871 VPB.n1360 VPB.n1359 13.653
R872 VPB.n1359 VPB.n1358 13.653
R873 VPB.n1367 VPB.n1366 13.653
R874 VPB.n1366 VPB.n1365 13.653
R875 VPB.n1372 VPB.n1371 13.653
R876 VPB.n1371 VPB.n1370 13.653
R877 VPB.n1377 VPB.n1376 13.653
R878 VPB.n1376 VPB.n1375 13.653
R879 VPB.n1384 VPB.n1383 13.653
R880 VPB.n1383 VPB.n1382 13.653
R881 VPB.n1389 VPB.n1388 13.653
R882 VPB.n1388 VPB.n1387 13.653
R883 VPB.n1394 VPB.n1393 13.653
R884 VPB.n1393 VPB.n1392 13.653
R885 VPB.n1398 VPB.n1397 13.653
R886 VPB.n1397 VPB.n1396 13.653
R887 VPB.n1402 VPB.n1401 13.653
R888 VPB.n1401 VPB.n1400 13.653
R889 VPB.n1429 VPB.n1428 13.653
R890 VPB.n1428 VPB.n1427 13.653
R891 VPB.n1433 VPB.n1432 13.653
R892 VPB.n1432 VPB.n1431 13.653
R893 VPB.n1438 VPB.n1437 13.653
R894 VPB.n1437 VPB.n1436 13.653
R895 VPB.n1443 VPB.n1442 13.653
R896 VPB.n1442 VPB.n1441 13.653
R897 VPB.n1450 VPB.n1449 13.653
R898 VPB.n1449 VPB.n1448 13.653
R899 VPB.n1455 VPB.n1454 13.653
R900 VPB.n1454 VPB.n1453 13.653
R901 VPB.n1460 VPB.n1459 13.653
R902 VPB.n1459 VPB.n1458 13.653
R903 VPB.n1467 VPB.n1466 13.653
R904 VPB.n1466 VPB.n1465 13.653
R905 VPB.n1472 VPB.n1471 13.653
R906 VPB.n1471 VPB.n1470 13.653
R907 VPB.n1477 VPB.n1476 13.653
R908 VPB.n1476 VPB.n1475 13.653
R909 VPB.n1481 VPB.n1480 13.653
R910 VPB.n1480 VPB.n1479 13.653
R911 VPB.n1485 VPB.n1484 13.653
R912 VPB.n1484 VPB.n1483 13.653
R913 VPB.n40 VPB.n39 13.653
R914 VPB.n39 VPB.n38 13.653
R915 VPB.n43 VPB.n42 13.653
R916 VPB.n42 VPB.n41 13.653
R917 VPB.n48 VPB.n47 13.653
R918 VPB.n47 VPB.n46 13.653
R919 VPB.n52 VPB.n51 13.653
R920 VPB.n51 VPB.n50 13.653
R921 VPB.n57 VPB.n56 13.653
R922 VPB.n56 VPB.n55 13.653
R923 VPB.n61 VPB.n60 13.653
R924 VPB.n60 VPB.n59 13.653
R925 VPB.n65 VPB.n64 13.653
R926 VPB.n64 VPB.n63 13.653
R927 VPB.n1494 VPB.n0 13.653
R928 VPB VPB.n0 13.653
R929 VPB.n218 VPB.n217 13.35
R930 VPB.n290 VPB.n289 13.35
R931 VPB.n364 VPB.n363 13.35
R932 VPB.n427 VPB.n426 13.35
R933 VPB.n499 VPB.n498 13.35
R934 VPB.n582 VPB.n581 13.35
R935 VPB.n656 VPB.n655 13.35
R936 VPB.n728 VPB.n727 13.35
R937 VPB.n802 VPB.n801 13.35
R938 VPB.n865 VPB.n864 13.35
R939 VPB.n937 VPB.n936 13.35
R940 VPB.n1020 VPB.n1019 13.35
R941 VPB.n1094 VPB.n1093 13.35
R942 VPB.n1166 VPB.n1165 13.35
R943 VPB.n1240 VPB.n1239 13.35
R944 VPB.n1303 VPB.n1302 13.35
R945 VPB.n1375 VPB.n1374 13.35
R946 VPB.n1458 VPB.n1457 13.35
R947 VPB.n55 VPB.n54 13.35
R948 VPB.n1498 VPB.n1497 13.276
R949 VPB.n1497 VPB.n1495 13.276
R950 VPB.n35 VPB.n17 13.276
R951 VPB.n17 VPB.n15 13.276
R952 VPB.n1424 VPB.n1406 13.276
R953 VPB.n1406 VPB.n1404 13.276
R954 VPB.n1341 VPB.n1323 13.276
R955 VPB.n1323 VPB.n1321 13.276
R956 VPB.n1278 VPB.n1260 13.276
R957 VPB.n1260 VPB.n1258 13.276
R958 VPB.n1215 VPB.n1197 13.276
R959 VPB.n1197 VPB.n1195 13.276
R960 VPB.n1132 VPB.n1114 13.276
R961 VPB.n1114 VPB.n1112 13.276
R962 VPB.n1069 VPB.n1051 13.276
R963 VPB.n1051 VPB.n1049 13.276
R964 VPB.n986 VPB.n968 13.276
R965 VPB.n968 VPB.n966 13.276
R966 VPB.n903 VPB.n885 13.276
R967 VPB.n885 VPB.n883 13.276
R968 VPB.n840 VPB.n822 13.276
R969 VPB.n822 VPB.n820 13.276
R970 VPB.n777 VPB.n759 13.276
R971 VPB.n759 VPB.n757 13.276
R972 VPB.n694 VPB.n676 13.276
R973 VPB.n676 VPB.n674 13.276
R974 VPB.n631 VPB.n613 13.276
R975 VPB.n613 VPB.n611 13.276
R976 VPB.n548 VPB.n530 13.276
R977 VPB.n530 VPB.n528 13.276
R978 VPB.n465 VPB.n447 13.276
R979 VPB.n447 VPB.n445 13.276
R980 VPB.n402 VPB.n384 13.276
R981 VPB.n384 VPB.n382 13.276
R982 VPB.n339 VPB.n321 13.276
R983 VPB.n321 VPB.n319 13.276
R984 VPB.n256 VPB.n238 13.276
R985 VPB.n238 VPB.n236 13.276
R986 VPB.n193 VPB.n175 13.276
R987 VPB.n175 VPB.n173 13.276
R988 VPB.n138 VPB.n120 13.276
R989 VPB.n120 VPB.n118 13.276
R990 VPB.n98 VPB.n95 13.276
R991 VPB.n95 VPB.n92 13.276
R992 VPB.n143 VPB.n139 13.276
R993 VPB.n198 VPB.n194 13.276
R994 VPB.n261 VPB.n257 13.276
R995 VPB.n344 VPB.n340 13.276
R996 VPB.n407 VPB.n403 13.276
R997 VPB.n470 VPB.n466 13.276
R998 VPB.n553 VPB.n549 13.276
R999 VPB.n636 VPB.n632 13.276
R1000 VPB.n699 VPB.n695 13.276
R1001 VPB.n782 VPB.n778 13.276
R1002 VPB.n845 VPB.n841 13.276
R1003 VPB.n908 VPB.n904 13.276
R1004 VPB.n991 VPB.n987 13.276
R1005 VPB.n1074 VPB.n1070 13.276
R1006 VPB.n1137 VPB.n1133 13.276
R1007 VPB.n1220 VPB.n1216 13.276
R1008 VPB.n1283 VPB.n1279 13.276
R1009 VPB.n1346 VPB.n1342 13.276
R1010 VPB.n1429 VPB.n1425 13.276
R1011 VPB.n40 VPB.n36 13.276
R1012 VPB.n43 VPB.n40 13.276
R1013 VPB.n52 VPB.n48 13.276
R1014 VPB.n61 VPB.n57 13.276
R1015 VPB.n86 VPB.n68 13.276
R1016 VPB.n68 VPB.n66 13.276
R1017 VPB.n73 VPB.n71 12.796
R1018 VPB.n73 VPB.n72 12.564
R1019 VPB.n82 VPB.n81 12.198
R1020 VPB.n79 VPB.n78 12.198
R1021 VPB.n79 VPB.n76 12.198
R1022 VPB.n48 VPB.n44 11.841
R1023 VPB.n62 VPB.n61 11.482
R1024 VPB.n86 VPB.n85 7.5
R1025 VPB.n71 VPB.n70 7.5
R1026 VPB.n78 VPB.n77 7.5
R1027 VPB.n76 VPB.n75 7.5
R1028 VPB.n68 VPB.n67 7.5
R1029 VPB.n83 VPB.n69 7.5
R1030 VPB.n120 VPB.n119 7.5
R1031 VPB.n133 VPB.n132 7.5
R1032 VPB.n127 VPB.n126 7.5
R1033 VPB.n129 VPB.n128 7.5
R1034 VPB.n122 VPB.n121 7.5
R1035 VPB.n138 VPB.n137 7.5
R1036 VPB.n175 VPB.n174 7.5
R1037 VPB.n188 VPB.n187 7.5
R1038 VPB.n182 VPB.n181 7.5
R1039 VPB.n184 VPB.n183 7.5
R1040 VPB.n177 VPB.n176 7.5
R1041 VPB.n193 VPB.n192 7.5
R1042 VPB.n238 VPB.n237 7.5
R1043 VPB.n251 VPB.n250 7.5
R1044 VPB.n245 VPB.n244 7.5
R1045 VPB.n247 VPB.n246 7.5
R1046 VPB.n240 VPB.n239 7.5
R1047 VPB.n256 VPB.n255 7.5
R1048 VPB.n321 VPB.n320 7.5
R1049 VPB.n334 VPB.n333 7.5
R1050 VPB.n328 VPB.n327 7.5
R1051 VPB.n330 VPB.n329 7.5
R1052 VPB.n323 VPB.n322 7.5
R1053 VPB.n339 VPB.n338 7.5
R1054 VPB.n384 VPB.n383 7.5
R1055 VPB.n397 VPB.n396 7.5
R1056 VPB.n391 VPB.n390 7.5
R1057 VPB.n393 VPB.n392 7.5
R1058 VPB.n386 VPB.n385 7.5
R1059 VPB.n402 VPB.n401 7.5
R1060 VPB.n447 VPB.n446 7.5
R1061 VPB.n460 VPB.n459 7.5
R1062 VPB.n454 VPB.n453 7.5
R1063 VPB.n456 VPB.n455 7.5
R1064 VPB.n449 VPB.n448 7.5
R1065 VPB.n465 VPB.n464 7.5
R1066 VPB.n530 VPB.n529 7.5
R1067 VPB.n543 VPB.n542 7.5
R1068 VPB.n537 VPB.n536 7.5
R1069 VPB.n539 VPB.n538 7.5
R1070 VPB.n532 VPB.n531 7.5
R1071 VPB.n548 VPB.n547 7.5
R1072 VPB.n613 VPB.n612 7.5
R1073 VPB.n626 VPB.n625 7.5
R1074 VPB.n620 VPB.n619 7.5
R1075 VPB.n622 VPB.n621 7.5
R1076 VPB.n615 VPB.n614 7.5
R1077 VPB.n631 VPB.n630 7.5
R1078 VPB.n676 VPB.n675 7.5
R1079 VPB.n689 VPB.n688 7.5
R1080 VPB.n683 VPB.n682 7.5
R1081 VPB.n685 VPB.n684 7.5
R1082 VPB.n678 VPB.n677 7.5
R1083 VPB.n694 VPB.n693 7.5
R1084 VPB.n759 VPB.n758 7.5
R1085 VPB.n772 VPB.n771 7.5
R1086 VPB.n766 VPB.n765 7.5
R1087 VPB.n768 VPB.n767 7.5
R1088 VPB.n761 VPB.n760 7.5
R1089 VPB.n777 VPB.n776 7.5
R1090 VPB.n822 VPB.n821 7.5
R1091 VPB.n835 VPB.n834 7.5
R1092 VPB.n829 VPB.n828 7.5
R1093 VPB.n831 VPB.n830 7.5
R1094 VPB.n824 VPB.n823 7.5
R1095 VPB.n840 VPB.n839 7.5
R1096 VPB.n885 VPB.n884 7.5
R1097 VPB.n898 VPB.n897 7.5
R1098 VPB.n892 VPB.n891 7.5
R1099 VPB.n894 VPB.n893 7.5
R1100 VPB.n887 VPB.n886 7.5
R1101 VPB.n903 VPB.n902 7.5
R1102 VPB.n968 VPB.n967 7.5
R1103 VPB.n981 VPB.n980 7.5
R1104 VPB.n975 VPB.n974 7.5
R1105 VPB.n977 VPB.n976 7.5
R1106 VPB.n970 VPB.n969 7.5
R1107 VPB.n986 VPB.n985 7.5
R1108 VPB.n1051 VPB.n1050 7.5
R1109 VPB.n1064 VPB.n1063 7.5
R1110 VPB.n1058 VPB.n1057 7.5
R1111 VPB.n1060 VPB.n1059 7.5
R1112 VPB.n1053 VPB.n1052 7.5
R1113 VPB.n1069 VPB.n1068 7.5
R1114 VPB.n1114 VPB.n1113 7.5
R1115 VPB.n1127 VPB.n1126 7.5
R1116 VPB.n1121 VPB.n1120 7.5
R1117 VPB.n1123 VPB.n1122 7.5
R1118 VPB.n1116 VPB.n1115 7.5
R1119 VPB.n1132 VPB.n1131 7.5
R1120 VPB.n1197 VPB.n1196 7.5
R1121 VPB.n1210 VPB.n1209 7.5
R1122 VPB.n1204 VPB.n1203 7.5
R1123 VPB.n1206 VPB.n1205 7.5
R1124 VPB.n1199 VPB.n1198 7.5
R1125 VPB.n1215 VPB.n1214 7.5
R1126 VPB.n1260 VPB.n1259 7.5
R1127 VPB.n1273 VPB.n1272 7.5
R1128 VPB.n1267 VPB.n1266 7.5
R1129 VPB.n1269 VPB.n1268 7.5
R1130 VPB.n1262 VPB.n1261 7.5
R1131 VPB.n1278 VPB.n1277 7.5
R1132 VPB.n1323 VPB.n1322 7.5
R1133 VPB.n1336 VPB.n1335 7.5
R1134 VPB.n1330 VPB.n1329 7.5
R1135 VPB.n1332 VPB.n1331 7.5
R1136 VPB.n1325 VPB.n1324 7.5
R1137 VPB.n1341 VPB.n1340 7.5
R1138 VPB.n1406 VPB.n1405 7.5
R1139 VPB.n1419 VPB.n1418 7.5
R1140 VPB.n1413 VPB.n1412 7.5
R1141 VPB.n1415 VPB.n1414 7.5
R1142 VPB.n1408 VPB.n1407 7.5
R1143 VPB.n1424 VPB.n1423 7.5
R1144 VPB.n17 VPB.n16 7.5
R1145 VPB.n30 VPB.n29 7.5
R1146 VPB.n24 VPB.n23 7.5
R1147 VPB.n26 VPB.n25 7.5
R1148 VPB.n19 VPB.n18 7.5
R1149 VPB.n35 VPB.n34 7.5
R1150 VPB.n1497 VPB.n1496 7.5
R1151 VPB.n12 VPB.n11 7.5
R1152 VPB.n6 VPB.n5 7.5
R1153 VPB.n8 VPB.n7 7.5
R1154 VPB.n2 VPB.n1 7.5
R1155 VPB.n1499 VPB.n1498 7.5
R1156 VPB.n36 VPB.n35 7.176
R1157 VPB.n1425 VPB.n1424 7.176
R1158 VPB.n1342 VPB.n1341 7.176
R1159 VPB.n1279 VPB.n1278 7.176
R1160 VPB.n1216 VPB.n1215 7.176
R1161 VPB.n1133 VPB.n1132 7.176
R1162 VPB.n1070 VPB.n1069 7.176
R1163 VPB.n987 VPB.n986 7.176
R1164 VPB.n904 VPB.n903 7.176
R1165 VPB.n841 VPB.n840 7.176
R1166 VPB.n778 VPB.n777 7.176
R1167 VPB.n695 VPB.n694 7.176
R1168 VPB.n632 VPB.n631 7.176
R1169 VPB.n549 VPB.n548 7.176
R1170 VPB.n466 VPB.n465 7.176
R1171 VPB.n403 VPB.n402 7.176
R1172 VPB.n340 VPB.n339 7.176
R1173 VPB.n257 VPB.n256 7.176
R1174 VPB.n194 VPB.n193 7.176
R1175 VPB.n139 VPB.n138 7.176
R1176 VPB.n57 VPB.n53 6.817
R1177 VPB.n134 VPB.n131 6.729
R1178 VPB.n130 VPB.n127 6.729
R1179 VPB.n125 VPB.n122 6.729
R1180 VPB.n189 VPB.n186 6.729
R1181 VPB.n185 VPB.n182 6.729
R1182 VPB.n180 VPB.n177 6.729
R1183 VPB.n252 VPB.n249 6.729
R1184 VPB.n248 VPB.n245 6.729
R1185 VPB.n243 VPB.n240 6.729
R1186 VPB.n335 VPB.n332 6.729
R1187 VPB.n331 VPB.n328 6.729
R1188 VPB.n326 VPB.n323 6.729
R1189 VPB.n398 VPB.n395 6.729
R1190 VPB.n394 VPB.n391 6.729
R1191 VPB.n389 VPB.n386 6.729
R1192 VPB.n461 VPB.n458 6.729
R1193 VPB.n457 VPB.n454 6.729
R1194 VPB.n452 VPB.n449 6.729
R1195 VPB.n544 VPB.n541 6.729
R1196 VPB.n540 VPB.n537 6.729
R1197 VPB.n535 VPB.n532 6.729
R1198 VPB.n627 VPB.n624 6.729
R1199 VPB.n623 VPB.n620 6.729
R1200 VPB.n618 VPB.n615 6.729
R1201 VPB.n690 VPB.n687 6.729
R1202 VPB.n686 VPB.n683 6.729
R1203 VPB.n681 VPB.n678 6.729
R1204 VPB.n773 VPB.n770 6.729
R1205 VPB.n769 VPB.n766 6.729
R1206 VPB.n764 VPB.n761 6.729
R1207 VPB.n836 VPB.n833 6.729
R1208 VPB.n832 VPB.n829 6.729
R1209 VPB.n827 VPB.n824 6.729
R1210 VPB.n899 VPB.n896 6.729
R1211 VPB.n895 VPB.n892 6.729
R1212 VPB.n890 VPB.n887 6.729
R1213 VPB.n982 VPB.n979 6.729
R1214 VPB.n978 VPB.n975 6.729
R1215 VPB.n973 VPB.n970 6.729
R1216 VPB.n1065 VPB.n1062 6.729
R1217 VPB.n1061 VPB.n1058 6.729
R1218 VPB.n1056 VPB.n1053 6.729
R1219 VPB.n1128 VPB.n1125 6.729
R1220 VPB.n1124 VPB.n1121 6.729
R1221 VPB.n1119 VPB.n1116 6.729
R1222 VPB.n1211 VPB.n1208 6.729
R1223 VPB.n1207 VPB.n1204 6.729
R1224 VPB.n1202 VPB.n1199 6.729
R1225 VPB.n1274 VPB.n1271 6.729
R1226 VPB.n1270 VPB.n1267 6.729
R1227 VPB.n1265 VPB.n1262 6.729
R1228 VPB.n1337 VPB.n1334 6.729
R1229 VPB.n1333 VPB.n1330 6.729
R1230 VPB.n1328 VPB.n1325 6.729
R1231 VPB.n1420 VPB.n1417 6.729
R1232 VPB.n1416 VPB.n1413 6.729
R1233 VPB.n1411 VPB.n1408 6.729
R1234 VPB.n31 VPB.n28 6.729
R1235 VPB.n27 VPB.n24 6.729
R1236 VPB.n22 VPB.n19 6.729
R1237 VPB.n13 VPB.n10 6.729
R1238 VPB.n9 VPB.n6 6.729
R1239 VPB.n4 VPB.n2 6.729
R1240 VPB.n125 VPB.n124 6.728
R1241 VPB.n130 VPB.n129 6.728
R1242 VPB.n134 VPB.n133 6.728
R1243 VPB.n137 VPB.n136 6.728
R1244 VPB.n180 VPB.n179 6.728
R1245 VPB.n185 VPB.n184 6.728
R1246 VPB.n189 VPB.n188 6.728
R1247 VPB.n192 VPB.n191 6.728
R1248 VPB.n243 VPB.n242 6.728
R1249 VPB.n248 VPB.n247 6.728
R1250 VPB.n252 VPB.n251 6.728
R1251 VPB.n255 VPB.n254 6.728
R1252 VPB.n326 VPB.n325 6.728
R1253 VPB.n331 VPB.n330 6.728
R1254 VPB.n335 VPB.n334 6.728
R1255 VPB.n338 VPB.n337 6.728
R1256 VPB.n389 VPB.n388 6.728
R1257 VPB.n394 VPB.n393 6.728
R1258 VPB.n398 VPB.n397 6.728
R1259 VPB.n401 VPB.n400 6.728
R1260 VPB.n452 VPB.n451 6.728
R1261 VPB.n457 VPB.n456 6.728
R1262 VPB.n461 VPB.n460 6.728
R1263 VPB.n464 VPB.n463 6.728
R1264 VPB.n535 VPB.n534 6.728
R1265 VPB.n540 VPB.n539 6.728
R1266 VPB.n544 VPB.n543 6.728
R1267 VPB.n547 VPB.n546 6.728
R1268 VPB.n618 VPB.n617 6.728
R1269 VPB.n623 VPB.n622 6.728
R1270 VPB.n627 VPB.n626 6.728
R1271 VPB.n630 VPB.n629 6.728
R1272 VPB.n681 VPB.n680 6.728
R1273 VPB.n686 VPB.n685 6.728
R1274 VPB.n690 VPB.n689 6.728
R1275 VPB.n693 VPB.n692 6.728
R1276 VPB.n764 VPB.n763 6.728
R1277 VPB.n769 VPB.n768 6.728
R1278 VPB.n773 VPB.n772 6.728
R1279 VPB.n776 VPB.n775 6.728
R1280 VPB.n827 VPB.n826 6.728
R1281 VPB.n832 VPB.n831 6.728
R1282 VPB.n836 VPB.n835 6.728
R1283 VPB.n839 VPB.n838 6.728
R1284 VPB.n890 VPB.n889 6.728
R1285 VPB.n895 VPB.n894 6.728
R1286 VPB.n899 VPB.n898 6.728
R1287 VPB.n902 VPB.n901 6.728
R1288 VPB.n973 VPB.n972 6.728
R1289 VPB.n978 VPB.n977 6.728
R1290 VPB.n982 VPB.n981 6.728
R1291 VPB.n985 VPB.n984 6.728
R1292 VPB.n1056 VPB.n1055 6.728
R1293 VPB.n1061 VPB.n1060 6.728
R1294 VPB.n1065 VPB.n1064 6.728
R1295 VPB.n1068 VPB.n1067 6.728
R1296 VPB.n1119 VPB.n1118 6.728
R1297 VPB.n1124 VPB.n1123 6.728
R1298 VPB.n1128 VPB.n1127 6.728
R1299 VPB.n1131 VPB.n1130 6.728
R1300 VPB.n1202 VPB.n1201 6.728
R1301 VPB.n1207 VPB.n1206 6.728
R1302 VPB.n1211 VPB.n1210 6.728
R1303 VPB.n1214 VPB.n1213 6.728
R1304 VPB.n1265 VPB.n1264 6.728
R1305 VPB.n1270 VPB.n1269 6.728
R1306 VPB.n1274 VPB.n1273 6.728
R1307 VPB.n1277 VPB.n1276 6.728
R1308 VPB.n1328 VPB.n1327 6.728
R1309 VPB.n1333 VPB.n1332 6.728
R1310 VPB.n1337 VPB.n1336 6.728
R1311 VPB.n1340 VPB.n1339 6.728
R1312 VPB.n1411 VPB.n1410 6.728
R1313 VPB.n1416 VPB.n1415 6.728
R1314 VPB.n1420 VPB.n1419 6.728
R1315 VPB.n1423 VPB.n1422 6.728
R1316 VPB.n22 VPB.n21 6.728
R1317 VPB.n27 VPB.n26 6.728
R1318 VPB.n31 VPB.n30 6.728
R1319 VPB.n34 VPB.n33 6.728
R1320 VPB.n4 VPB.n3 6.728
R1321 VPB.n9 VPB.n8 6.728
R1322 VPB.n13 VPB.n12 6.728
R1323 VPB.n1500 VPB.n1499 6.728
R1324 VPB.n215 VPB.n211 6.458
R1325 VPB.n361 VPB.n357 6.458
R1326 VPB.n424 VPB.n420 6.458
R1327 VPB.n653 VPB.n649 6.458
R1328 VPB.n799 VPB.n795 6.458
R1329 VPB.n862 VPB.n858 6.458
R1330 VPB.n1091 VPB.n1087 6.458
R1331 VPB.n1237 VPB.n1233 6.458
R1332 VPB.n1300 VPB.n1296 6.458
R1333 VPB.n53 VPB.n52 6.458
R1334 VPB.n85 VPB.n84 6.398
R1335 VPB.n99 VPB.n89 6.112
R1336 VPB.n1494 VPB.n1493 6.111
R1337 VPB.n99 VPB.n98 6.101
R1338 VPB.n1493 VPB.n65 6.1
R1339 VPB.n299 VPB.n295 4.305
R1340 VPB.n508 VPB.n504 4.305
R1341 VPB.n591 VPB.n587 4.305
R1342 VPB.n737 VPB.n733 4.305
R1343 VPB.n946 VPB.n942 4.305
R1344 VPB.n1029 VPB.n1025 4.305
R1345 VPB.n1175 VPB.n1171 4.305
R1346 VPB.n1384 VPB.n1380 4.305
R1347 VPB.n1467 VPB.n1463 4.305
R1348 VPB.n282 VPB.n278 3.947
R1349 VPB.n491 VPB.n487 3.947
R1350 VPB.n574 VPB.n570 3.947
R1351 VPB.n720 VPB.n716 3.947
R1352 VPB.n929 VPB.n925 3.947
R1353 VPB.n1012 VPB.n1008 3.947
R1354 VPB.n1158 VPB.n1154 3.947
R1355 VPB.n1367 VPB.n1363 3.947
R1356 VPB.n1450 VPB.n1446 3.947
R1357 VPB.n230 VPB.n227 1.794
R1358 VPB.n376 VPB.n373 1.794
R1359 VPB.n439 VPB.n436 1.794
R1360 VPB.n668 VPB.n665 1.794
R1361 VPB.n814 VPB.n811 1.794
R1362 VPB.n877 VPB.n874 1.794
R1363 VPB.n1106 VPB.n1103 1.794
R1364 VPB.n1252 VPB.n1249 1.794
R1365 VPB.n1315 VPB.n1312 1.794
R1366 VPB.n65 VPB.n62 1.794
R1367 VPB.n203 VPB.n200 1.435
R1368 VPB.n349 VPB.n346 1.435
R1369 VPB.n412 VPB.n409 1.435
R1370 VPB.n641 VPB.n638 1.435
R1371 VPB.n787 VPB.n784 1.435
R1372 VPB.n850 VPB.n847 1.435
R1373 VPB.n1079 VPB.n1076 1.435
R1374 VPB.n1225 VPB.n1222 1.435
R1375 VPB.n1288 VPB.n1285 1.435
R1376 VPB.n44 VPB.n43 1.435
R1377 VPB.n83 VPB.n74 1.402
R1378 VPB.n83 VPB.n79 1.402
R1379 VPB.n83 VPB.n80 1.402
R1380 VPB.n83 VPB.n82 1.402
R1381 VPB.n270 VPB.n267 1.076
R1382 VPB.n479 VPB.n476 1.076
R1383 VPB.n562 VPB.n559 1.076
R1384 VPB.n708 VPB.n705 1.076
R1385 VPB.n917 VPB.n914 1.076
R1386 VPB.n1000 VPB.n997 1.076
R1387 VPB.n1146 VPB.n1143 1.076
R1388 VPB.n1355 VPB.n1352 1.076
R1389 VPB.n1438 VPB.n1435 1.076
R1390 VPB.n84 VPB.n83 0.735
R1391 VPB.n83 VPB.n73 0.735
R1392 VPB.n309 VPB.n306 0.717
R1393 VPB.n518 VPB.n515 0.717
R1394 VPB.n601 VPB.n598 0.717
R1395 VPB.n747 VPB.n744 0.717
R1396 VPB.n956 VPB.n953 0.717
R1397 VPB.n1039 VPB.n1036 0.717
R1398 VPB.n1185 VPB.n1182 0.717
R1399 VPB.n1394 VPB.n1391 0.717
R1400 VPB.n1477 VPB.n1474 0.717
R1401 VPB.n135 VPB.n134 0.387
R1402 VPB.n135 VPB.n130 0.387
R1403 VPB.n135 VPB.n125 0.387
R1404 VPB.n136 VPB.n135 0.387
R1405 VPB.n190 VPB.n189 0.387
R1406 VPB.n190 VPB.n185 0.387
R1407 VPB.n190 VPB.n180 0.387
R1408 VPB.n191 VPB.n190 0.387
R1409 VPB.n253 VPB.n252 0.387
R1410 VPB.n253 VPB.n248 0.387
R1411 VPB.n253 VPB.n243 0.387
R1412 VPB.n254 VPB.n253 0.387
R1413 VPB.n336 VPB.n335 0.387
R1414 VPB.n336 VPB.n331 0.387
R1415 VPB.n336 VPB.n326 0.387
R1416 VPB.n337 VPB.n336 0.387
R1417 VPB.n399 VPB.n398 0.387
R1418 VPB.n399 VPB.n394 0.387
R1419 VPB.n399 VPB.n389 0.387
R1420 VPB.n400 VPB.n399 0.387
R1421 VPB.n462 VPB.n461 0.387
R1422 VPB.n462 VPB.n457 0.387
R1423 VPB.n462 VPB.n452 0.387
R1424 VPB.n463 VPB.n462 0.387
R1425 VPB.n545 VPB.n544 0.387
R1426 VPB.n545 VPB.n540 0.387
R1427 VPB.n545 VPB.n535 0.387
R1428 VPB.n546 VPB.n545 0.387
R1429 VPB.n628 VPB.n627 0.387
R1430 VPB.n628 VPB.n623 0.387
R1431 VPB.n628 VPB.n618 0.387
R1432 VPB.n629 VPB.n628 0.387
R1433 VPB.n691 VPB.n690 0.387
R1434 VPB.n691 VPB.n686 0.387
R1435 VPB.n691 VPB.n681 0.387
R1436 VPB.n692 VPB.n691 0.387
R1437 VPB.n774 VPB.n773 0.387
R1438 VPB.n774 VPB.n769 0.387
R1439 VPB.n774 VPB.n764 0.387
R1440 VPB.n775 VPB.n774 0.387
R1441 VPB.n837 VPB.n836 0.387
R1442 VPB.n837 VPB.n832 0.387
R1443 VPB.n837 VPB.n827 0.387
R1444 VPB.n838 VPB.n837 0.387
R1445 VPB.n900 VPB.n899 0.387
R1446 VPB.n900 VPB.n895 0.387
R1447 VPB.n900 VPB.n890 0.387
R1448 VPB.n901 VPB.n900 0.387
R1449 VPB.n983 VPB.n982 0.387
R1450 VPB.n983 VPB.n978 0.387
R1451 VPB.n983 VPB.n973 0.387
R1452 VPB.n984 VPB.n983 0.387
R1453 VPB.n1066 VPB.n1065 0.387
R1454 VPB.n1066 VPB.n1061 0.387
R1455 VPB.n1066 VPB.n1056 0.387
R1456 VPB.n1067 VPB.n1066 0.387
R1457 VPB.n1129 VPB.n1128 0.387
R1458 VPB.n1129 VPB.n1124 0.387
R1459 VPB.n1129 VPB.n1119 0.387
R1460 VPB.n1130 VPB.n1129 0.387
R1461 VPB.n1212 VPB.n1211 0.387
R1462 VPB.n1212 VPB.n1207 0.387
R1463 VPB.n1212 VPB.n1202 0.387
R1464 VPB.n1213 VPB.n1212 0.387
R1465 VPB.n1275 VPB.n1274 0.387
R1466 VPB.n1275 VPB.n1270 0.387
R1467 VPB.n1275 VPB.n1265 0.387
R1468 VPB.n1276 VPB.n1275 0.387
R1469 VPB.n1338 VPB.n1337 0.387
R1470 VPB.n1338 VPB.n1333 0.387
R1471 VPB.n1338 VPB.n1328 0.387
R1472 VPB.n1339 VPB.n1338 0.387
R1473 VPB.n1421 VPB.n1420 0.387
R1474 VPB.n1421 VPB.n1416 0.387
R1475 VPB.n1421 VPB.n1411 0.387
R1476 VPB.n1422 VPB.n1421 0.387
R1477 VPB.n32 VPB.n31 0.387
R1478 VPB.n32 VPB.n27 0.387
R1479 VPB.n32 VPB.n22 0.387
R1480 VPB.n33 VPB.n32 0.387
R1481 VPB.n1501 VPB.n13 0.387
R1482 VPB.n1501 VPB.n9 0.387
R1483 VPB.n1501 VPB.n4 0.387
R1484 VPB.n1501 VPB.n1500 0.387
R1485 VPB.n144 VPB.n117 0.272
R1486 VPB.n199 VPB.n172 0.272
R1487 VPB.n262 VPB.n235 0.272
R1488 VPB.n345 VPB.n318 0.272
R1489 VPB.n408 VPB.n381 0.272
R1490 VPB.n471 VPB.n444 0.272
R1491 VPB.n554 VPB.n527 0.272
R1492 VPB.n637 VPB.n610 0.272
R1493 VPB.n700 VPB.n673 0.272
R1494 VPB.n783 VPB.n756 0.272
R1495 VPB.n846 VPB.n819 0.272
R1496 VPB.n909 VPB.n882 0.272
R1497 VPB.n992 VPB.n965 0.272
R1498 VPB.n1075 VPB.n1048 0.272
R1499 VPB.n1138 VPB.n1111 0.272
R1500 VPB.n1221 VPB.n1194 0.272
R1501 VPB.n1284 VPB.n1257 0.272
R1502 VPB.n1347 VPB.n1320 0.272
R1503 VPB.n1430 VPB.n1403 0.272
R1504 VPB.n1487 VPB.n1486 0.272
R1505 VPB.n101 VPB.n100 0.136
R1506 VPB.n105 VPB.n101 0.136
R1507 VPB.n109 VPB.n105 0.136
R1508 VPB.n113 VPB.n109 0.136
R1509 VPB.n117 VPB.n113 0.136
R1510 VPB.n148 VPB.n144 0.136
R1511 VPB.n152 VPB.n148 0.136
R1512 VPB.n156 VPB.n152 0.136
R1513 VPB.n160 VPB.n156 0.136
R1514 VPB.n164 VPB.n160 0.136
R1515 VPB.n168 VPB.n164 0.136
R1516 VPB.n172 VPB.n168 0.136
R1517 VPB.n204 VPB.n199 0.136
R1518 VPB.n209 VPB.n204 0.136
R1519 VPB.n216 VPB.n209 0.136
R1520 VPB.n221 VPB.n216 0.136
R1521 VPB.n226 VPB.n221 0.136
R1522 VPB.n231 VPB.n226 0.136
R1523 VPB.n235 VPB.n231 0.136
R1524 VPB.n266 VPB.n262 0.136
R1525 VPB.n271 VPB.n266 0.136
R1526 VPB.n276 VPB.n271 0.136
R1527 VPB.n283 VPB.n276 0.136
R1528 VPB.n288 VPB.n283 0.136
R1529 VPB.n293 VPB.n288 0.136
R1530 VPB.n300 VPB.n293 0.136
R1531 VPB.n305 VPB.n300 0.136
R1532 VPB.n310 VPB.n305 0.136
R1533 VPB.n314 VPB.n310 0.136
R1534 VPB.n318 VPB.n314 0.136
R1535 VPB.n350 VPB.n345 0.136
R1536 VPB.n355 VPB.n350 0.136
R1537 VPB.n362 VPB.n355 0.136
R1538 VPB.n367 VPB.n362 0.136
R1539 VPB.n372 VPB.n367 0.136
R1540 VPB.n377 VPB.n372 0.136
R1541 VPB.n381 VPB.n377 0.136
R1542 VPB.n413 VPB.n408 0.136
R1543 VPB.n418 VPB.n413 0.136
R1544 VPB.n425 VPB.n418 0.136
R1545 VPB.n430 VPB.n425 0.136
R1546 VPB.n435 VPB.n430 0.136
R1547 VPB.n440 VPB.n435 0.136
R1548 VPB.n444 VPB.n440 0.136
R1549 VPB.n475 VPB.n471 0.136
R1550 VPB.n480 VPB.n475 0.136
R1551 VPB.n485 VPB.n480 0.136
R1552 VPB.n492 VPB.n485 0.136
R1553 VPB.n497 VPB.n492 0.136
R1554 VPB.n502 VPB.n497 0.136
R1555 VPB.n509 VPB.n502 0.136
R1556 VPB.n514 VPB.n509 0.136
R1557 VPB.n519 VPB.n514 0.136
R1558 VPB.n523 VPB.n519 0.136
R1559 VPB.n527 VPB.n523 0.136
R1560 VPB.n558 VPB.n554 0.136
R1561 VPB.n563 VPB.n558 0.136
R1562 VPB.n568 VPB.n563 0.136
R1563 VPB.n575 VPB.n568 0.136
R1564 VPB.n580 VPB.n575 0.136
R1565 VPB.n585 VPB.n580 0.136
R1566 VPB.n592 VPB.n585 0.136
R1567 VPB.n597 VPB.n592 0.136
R1568 VPB.n602 VPB.n597 0.136
R1569 VPB.n606 VPB.n602 0.136
R1570 VPB.n610 VPB.n606 0.136
R1571 VPB.n642 VPB.n637 0.136
R1572 VPB.n647 VPB.n642 0.136
R1573 VPB.n654 VPB.n647 0.136
R1574 VPB.n659 VPB.n654 0.136
R1575 VPB.n664 VPB.n659 0.136
R1576 VPB.n669 VPB.n664 0.136
R1577 VPB.n673 VPB.n669 0.136
R1578 VPB.n704 VPB.n700 0.136
R1579 VPB.n709 VPB.n704 0.136
R1580 VPB.n714 VPB.n709 0.136
R1581 VPB.n721 VPB.n714 0.136
R1582 VPB.n726 VPB.n721 0.136
R1583 VPB.n731 VPB.n726 0.136
R1584 VPB.n738 VPB.n731 0.136
R1585 VPB.n743 VPB.n738 0.136
R1586 VPB.n748 VPB.n743 0.136
R1587 VPB.n752 VPB.n748 0.136
R1588 VPB.n756 VPB.n752 0.136
R1589 VPB.n788 VPB.n783 0.136
R1590 VPB.n793 VPB.n788 0.136
R1591 VPB.n800 VPB.n793 0.136
R1592 VPB.n805 VPB.n800 0.136
R1593 VPB.n810 VPB.n805 0.136
R1594 VPB.n815 VPB.n810 0.136
R1595 VPB.n819 VPB.n815 0.136
R1596 VPB.n851 VPB.n846 0.136
R1597 VPB.n856 VPB.n851 0.136
R1598 VPB.n863 VPB.n856 0.136
R1599 VPB.n868 VPB.n863 0.136
R1600 VPB.n873 VPB.n868 0.136
R1601 VPB.n878 VPB.n873 0.136
R1602 VPB.n882 VPB.n878 0.136
R1603 VPB.n913 VPB.n909 0.136
R1604 VPB.n918 VPB.n913 0.136
R1605 VPB.n923 VPB.n918 0.136
R1606 VPB.n930 VPB.n923 0.136
R1607 VPB.n935 VPB.n930 0.136
R1608 VPB.n940 VPB.n935 0.136
R1609 VPB.n947 VPB.n940 0.136
R1610 VPB.n952 VPB.n947 0.136
R1611 VPB.n957 VPB.n952 0.136
R1612 VPB.n961 VPB.n957 0.136
R1613 VPB.n965 VPB.n961 0.136
R1614 VPB.n996 VPB.n992 0.136
R1615 VPB.n1001 VPB.n996 0.136
R1616 VPB.n1006 VPB.n1001 0.136
R1617 VPB.n1013 VPB.n1006 0.136
R1618 VPB.n1018 VPB.n1013 0.136
R1619 VPB.n1023 VPB.n1018 0.136
R1620 VPB.n1030 VPB.n1023 0.136
R1621 VPB.n1035 VPB.n1030 0.136
R1622 VPB.n1040 VPB.n1035 0.136
R1623 VPB.n1044 VPB.n1040 0.136
R1624 VPB.n1048 VPB.n1044 0.136
R1625 VPB.n1080 VPB.n1075 0.136
R1626 VPB.n1085 VPB.n1080 0.136
R1627 VPB.n1092 VPB.n1085 0.136
R1628 VPB.n1097 VPB.n1092 0.136
R1629 VPB.n1102 VPB.n1097 0.136
R1630 VPB.n1107 VPB.n1102 0.136
R1631 VPB.n1111 VPB.n1107 0.136
R1632 VPB.n1142 VPB.n1138 0.136
R1633 VPB.n1147 VPB.n1142 0.136
R1634 VPB.n1152 VPB.n1147 0.136
R1635 VPB.n1159 VPB.n1152 0.136
R1636 VPB.n1164 VPB.n1159 0.136
R1637 VPB.n1169 VPB.n1164 0.136
R1638 VPB.n1176 VPB.n1169 0.136
R1639 VPB.n1181 VPB.n1176 0.136
R1640 VPB.n1186 VPB.n1181 0.136
R1641 VPB.n1190 VPB.n1186 0.136
R1642 VPB.n1194 VPB.n1190 0.136
R1643 VPB.n1226 VPB.n1221 0.136
R1644 VPB.n1231 VPB.n1226 0.136
R1645 VPB.n1238 VPB.n1231 0.136
R1646 VPB.n1243 VPB.n1238 0.136
R1647 VPB.n1248 VPB.n1243 0.136
R1648 VPB.n1253 VPB.n1248 0.136
R1649 VPB.n1257 VPB.n1253 0.136
R1650 VPB.n1289 VPB.n1284 0.136
R1651 VPB.n1294 VPB.n1289 0.136
R1652 VPB.n1301 VPB.n1294 0.136
R1653 VPB.n1306 VPB.n1301 0.136
R1654 VPB.n1311 VPB.n1306 0.136
R1655 VPB.n1316 VPB.n1311 0.136
R1656 VPB.n1320 VPB.n1316 0.136
R1657 VPB.n1351 VPB.n1347 0.136
R1658 VPB.n1356 VPB.n1351 0.136
R1659 VPB.n1361 VPB.n1356 0.136
R1660 VPB.n1368 VPB.n1361 0.136
R1661 VPB.n1373 VPB.n1368 0.136
R1662 VPB.n1378 VPB.n1373 0.136
R1663 VPB.n1385 VPB.n1378 0.136
R1664 VPB.n1390 VPB.n1385 0.136
R1665 VPB.n1395 VPB.n1390 0.136
R1666 VPB.n1399 VPB.n1395 0.136
R1667 VPB.n1403 VPB.n1399 0.136
R1668 VPB.n1434 VPB.n1430 0.136
R1669 VPB.n1439 VPB.n1434 0.136
R1670 VPB.n1444 VPB.n1439 0.136
R1671 VPB.n1451 VPB.n1444 0.136
R1672 VPB.n1456 VPB.n1451 0.136
R1673 VPB.n1461 VPB.n1456 0.136
R1674 VPB.n1468 VPB.n1461 0.136
R1675 VPB.n1473 VPB.n1468 0.136
R1676 VPB.n1478 VPB.n1473 0.136
R1677 VPB.n1482 VPB.n1478 0.136
R1678 VPB.n1486 VPB.n1482 0.136
R1679 VPB.n1488 VPB.n1487 0.136
R1680 VPB.n1489 VPB.n1488 0.136
R1681 VPB.n1490 VPB.n1489 0.136
R1682 VPB.n1491 VPB.n1490 0.136
R1683 VPB.n1492 VPB.n1491 0.136
R1684 a_3473_1004.n8 a_3473_1004.t9 512.525
R1685 a_3473_1004.n4 a_3473_1004.t5 512.525
R1686 a_3473_1004.n3 a_3473_1004.t11 512.525
R1687 a_3473_1004.n8 a_3473_1004.t13 371.139
R1688 a_3473_1004.n4 a_3473_1004.t12 371.139
R1689 a_3473_1004.n3 a_3473_1004.t6 371.139
R1690 a_3473_1004.n9 a_3473_1004.t8 266.342
R1691 a_3473_1004.n5 a_3473_1004.n4 258.98
R1692 a_3473_1004.n13 a_3473_1004.n11 200.608
R1693 a_3473_1004.n5 a_3473_1004.t10 176.995
R1694 a_3473_1004.n9 a_3473_1004.n8 172.76
R1695 a_3473_1004.n6 a_3473_1004.t7 170.569
R1696 a_3473_1004.n7 a_3473_1004.n3 169.274
R1697 a_3473_1004.n11 a_3473_1004.n2 162.547
R1698 a_3473_1004.n6 a_3473_1004.n5 153.043
R1699 a_3473_1004.n10 a_3473_1004.n7 118.94
R1700 a_3473_1004.n7 a_3473_1004.n6 89.705
R1701 a_3473_1004.n11 a_3473_1004.n10 77.315
R1702 a_3473_1004.n2 a_3473_1004.n1 76.002
R1703 a_3473_1004.n10 a_3473_1004.n9 76
R1704 a_3473_1004.n13 a_3473_1004.n12 15.218
R1705 a_3473_1004.n0 a_3473_1004.t1 14.282
R1706 a_3473_1004.n0 a_3473_1004.t2 14.282
R1707 a_3473_1004.n1 a_3473_1004.t3 14.282
R1708 a_3473_1004.n1 a_3473_1004.t4 14.282
R1709 a_3473_1004.n2 a_3473_1004.n0 12.85
R1710 a_3473_1004.n14 a_3473_1004.n13 12.014
R1711 a_15044_181.n11 a_15044_181.n2 336.934
R1712 a_15044_181.n10 a_15044_181.n9 114.024
R1713 a_15044_181.n10 a_15044_181.n6 96.417
R1714 a_15044_181.n11 a_15044_181.n10 78.403
R1715 a_15044_181.n2 a_15044_181.n1 75.271
R1716 a_15044_181.n6 a_15044_181.n5 30
R1717 a_15044_181.n13 a_15044_181.n11 27.275
R1718 a_15044_181.n4 a_15044_181.n3 24.383
R1719 a_15044_181.n6 a_15044_181.n4 23.684
R1720 a_15044_181.n9 a_15044_181.n8 22.578
R1721 a_15044_181.n13 a_15044_181.n12 15.001
R1722 a_15044_181.n0 a_15044_181.t1 14.282
R1723 a_15044_181.n0 a_15044_181.t0 14.282
R1724 a_15044_181.n1 a_15044_181.t4 14.282
R1725 a_15044_181.n1 a_15044_181.t6 14.282
R1726 a_15044_181.n14 a_15044_181.n13 12.632
R1727 a_15044_181.n2 a_15044_181.n0 12.119
R1728 a_15044_181.n9 a_15044_181.n7 8.58
R1729 a_15533_1005.n3 a_15533_1005.n2 196.002
R1730 a_15533_1005.n4 a_15533_1005.t1 89.553
R1731 a_15533_1005.n2 a_15533_1005.n1 75.271
R1732 a_15533_1005.n4 a_15533_1005.n3 75.214
R1733 a_15533_1005.n2 a_15533_1005.n0 36.52
R1734 a_15533_1005.n3 a_15533_1005.t4 14.338
R1735 a_15533_1005.n0 a_15533_1005.t3 14.282
R1736 a_15533_1005.n0 a_15533_1005.t2 14.282
R1737 a_15533_1005.n1 a_15533_1005.t7 14.282
R1738 a_15533_1005.n1 a_15533_1005.t6 14.282
R1739 a_15533_1005.n5 a_15533_1005.t0 14.282
R1740 a_15533_1005.t5 a_15533_1005.n5 14.282
R1741 a_15533_1005.n5 a_15533_1005.n4 12.122
R1742 a_3599_383.n6 a_3599_383.t9 472.359
R1743 a_3599_383.n6 a_3599_383.t7 384.527
R1744 a_3599_383.n7 a_3599_383.t8 277.772
R1745 a_3599_383.n10 a_3599_383.n8 249.704
R1746 a_3599_383.n8 a_3599_383.n7 156.035
R1747 a_3599_383.n8 a_3599_383.n5 127.74
R1748 a_3599_383.n4 a_3599_383.n3 79.232
R1749 a_3599_383.n7 a_3599_383.n6 67.001
R1750 a_3599_383.n5 a_3599_383.n4 63.152
R1751 a_3599_383.n11 a_3599_383.n0 55.263
R1752 a_3599_383.n10 a_3599_383.n9 30
R1753 a_3599_383.n11 a_3599_383.n10 23.684
R1754 a_3599_383.n5 a_3599_383.n1 16.08
R1755 a_3599_383.n4 a_3599_383.n2 16.08
R1756 a_3599_383.n1 a_3599_383.t0 14.282
R1757 a_3599_383.n1 a_3599_383.t1 14.282
R1758 a_3599_383.n2 a_3599_383.t5 14.282
R1759 a_3599_383.n2 a_3599_383.t6 14.282
R1760 a_3599_383.n3 a_3599_383.t4 14.282
R1761 a_3599_383.n3 a_3599_383.t3 14.282
R1762 a_11033_943.n6 a_11033_943.t7 454.685
R1763 a_11033_943.n8 a_11033_943.t11 454.685
R1764 a_11033_943.n4 a_11033_943.t13 454.685
R1765 a_11033_943.n6 a_11033_943.t6 428.979
R1766 a_11033_943.n8 a_11033_943.t9 428.979
R1767 a_11033_943.n4 a_11033_943.t10 428.979
R1768 a_11033_943.n7 a_11033_943.t8 248.006
R1769 a_11033_943.n9 a_11033_943.t5 248.006
R1770 a_11033_943.n5 a_11033_943.t12 248.006
R1771 a_11033_943.n14 a_11033_943.n12 220.639
R1772 a_11033_943.n12 a_11033_943.n3 135.994
R1773 a_11033_943.n7 a_11033_943.n6 81.941
R1774 a_11033_943.n9 a_11033_943.n8 81.941
R1775 a_11033_943.n5 a_11033_943.n4 81.941
R1776 a_11033_943.n11 a_11033_943.n5 81.396
R1777 a_11033_943.n10 a_11033_943.n9 79.491
R1778 a_11033_943.n3 a_11033_943.n2 76.002
R1779 a_11033_943.n10 a_11033_943.n7 76
R1780 a_11033_943.n12 a_11033_943.n11 76
R1781 a_11033_943.n14 a_11033_943.n13 30
R1782 a_11033_943.n15 a_11033_943.n0 24.383
R1783 a_11033_943.n15 a_11033_943.n14 23.684
R1784 a_11033_943.n1 a_11033_943.t2 14.282
R1785 a_11033_943.n1 a_11033_943.t1 14.282
R1786 a_11033_943.n2 a_11033_943.t4 14.282
R1787 a_11033_943.n2 a_11033_943.t3 14.282
R1788 a_11033_943.n3 a_11033_943.n1 12.85
R1789 a_11033_943.n11 a_11033_943.n10 2.947
R1790 a_8357_1004.n8 a_8357_1004.t5 512.525
R1791 a_8357_1004.n4 a_8357_1004.t6 475.572
R1792 a_8357_1004.n3 a_8357_1004.t7 469.145
R1793 a_8357_1004.n4 a_8357_1004.t10 384.527
R1794 a_8357_1004.n3 a_8357_1004.t11 384.527
R1795 a_8357_1004.n8 a_8357_1004.t9 371.139
R1796 a_8357_1004.n5 a_8357_1004.t12 277.772
R1797 a_8357_1004.n9 a_8357_1004.n8 225.866
R1798 a_8357_1004.n9 a_8357_1004.t13 218.057
R1799 a_8357_1004.n11 a_8357_1004.n2 215.652
R1800 a_8357_1004.n7 a_8357_1004.t8 198.113
R1801 a_8357_1004.n6 a_8357_1004.n5 156.851
R1802 a_8357_1004.n13 a_8357_1004.n11 147.503
R1803 a_8357_1004.n10 a_8357_1004.n7 98.138
R1804 a_8357_1004.n7 a_8357_1004.n6 79.658
R1805 a_8357_1004.n11 a_8357_1004.n10 77.315
R1806 a_8357_1004.n2 a_8357_1004.n1 76.002
R1807 a_8357_1004.n10 a_8357_1004.n9 76
R1808 a_8357_1004.n5 a_8357_1004.n4 67.889
R1809 a_8357_1004.n6 a_8357_1004.n3 66.88
R1810 a_8357_1004.n13 a_8357_1004.n12 15.218
R1811 a_8357_1004.n0 a_8357_1004.t0 14.282
R1812 a_8357_1004.n0 a_8357_1004.t2 14.282
R1813 a_8357_1004.n1 a_8357_1004.t4 14.282
R1814 a_8357_1004.n1 a_8357_1004.t3 14.282
R1815 a_8357_1004.n2 a_8357_1004.n0 12.85
R1816 a_8357_1004.n14 a_8357_1004.n13 12.014
R1817 a_8483_383.n6 a_8483_383.t8 472.359
R1818 a_8483_383.n6 a_8483_383.t9 384.527
R1819 a_8483_383.n7 a_8483_383.t7 277.772
R1820 a_8483_383.n10 a_8483_383.n8 249.704
R1821 a_8483_383.n8 a_8483_383.n7 156.035
R1822 a_8483_383.n8 a_8483_383.n5 127.74
R1823 a_8483_383.n4 a_8483_383.n3 79.232
R1824 a_8483_383.n7 a_8483_383.n6 67.001
R1825 a_8483_383.n5 a_8483_383.n4 63.152
R1826 a_8483_383.n10 a_8483_383.n9 30
R1827 a_8483_383.n11 a_8483_383.n0 24.383
R1828 a_8483_383.n11 a_8483_383.n10 23.684
R1829 a_8483_383.n5 a_8483_383.n1 16.08
R1830 a_8483_383.n4 a_8483_383.n2 16.08
R1831 a_8483_383.n1 a_8483_383.t5 14.282
R1832 a_8483_383.n1 a_8483_383.t4 14.282
R1833 a_8483_383.n2 a_8483_383.t2 14.282
R1834 a_8483_383.n2 a_8483_383.t3 14.282
R1835 a_8483_383.n3 a_8483_383.t1 14.282
R1836 a_8483_383.n3 a_8483_383.t0 14.282
R1837 a_9880_73.t0 a_9880_73.n1 93.333
R1838 a_9880_73.n4 a_9880_73.n2 55.07
R1839 a_9880_73.t0 a_9880_73.n0 8.137
R1840 a_9880_73.n4 a_9880_73.n3 4.619
R1841 a_9880_73.t0 a_9880_73.n4 0.071
R1842 VNB VNB.n1315 300.778
R1843 VNB.n117 VNB.n116 199.897
R1844 VNB.n176 VNB.n175 199.897
R1845 VNB.n228 VNB.n227 199.897
R1846 VNB.n303 VNB.n302 199.897
R1847 VNB.n355 VNB.n354 199.897
R1848 VNB.n414 VNB.n413 199.897
R1849 VNB.n482 VNB.n481 199.897
R1850 VNB.n550 VNB.n549 199.897
R1851 VNB.n602 VNB.n601 199.897
R1852 VNB.n677 VNB.n676 199.897
R1853 VNB.n736 VNB.n735 199.897
R1854 VNB.n795 VNB.n794 199.897
R1855 VNB.n863 VNB.n862 199.897
R1856 VNB.n931 VNB.n930 199.897
R1857 VNB.n990 VNB.n989 199.897
R1858 VNB.n1065 VNB.n1064 199.897
R1859 VNB.n1117 VNB.n1116 199.897
R1860 VNB.n1169 VNB.n1168 199.897
R1861 VNB.n1237 VNB.n1236 199.897
R1862 VNB.n18 VNB.n17 199.897
R1863 VNB.n126 VNB.n124 154.509
R1864 VNB.n237 VNB.n235 154.509
R1865 VNB.n185 VNB.n183 154.509
R1866 VNB.n364 VNB.n362 154.509
R1867 VNB.n312 VNB.n310 154.509
R1868 VNB.n491 VNB.n489 154.509
R1869 VNB.n423 VNB.n421 154.509
R1870 VNB.n611 VNB.n609 154.509
R1871 VNB.n559 VNB.n557 154.509
R1872 VNB.n745 VNB.n743 154.509
R1873 VNB.n686 VNB.n684 154.509
R1874 VNB.n872 VNB.n870 154.509
R1875 VNB.n804 VNB.n802 154.509
R1876 VNB.n999 VNB.n997 154.509
R1877 VNB.n940 VNB.n938 154.509
R1878 VNB.n1126 VNB.n1124 154.509
R1879 VNB.n1074 VNB.n1072 154.509
R1880 VNB.n1246 VNB.n1244 154.509
R1881 VNB.n1178 VNB.n1176 154.509
R1882 VNB.n27 VNB.n25 154.509
R1883 VNB.n269 VNB.n268 147.75
R1884 VNB.n643 VNB.n642 147.75
R1885 VNB.n1031 VNB.n1030 147.75
R1886 VNB.n83 VNB.n82 121.366
R1887 VNB.n142 VNB.n141 121.366
R1888 VNB.n281 VNB.n278 121.366
R1889 VNB.n380 VNB.n379 121.366
R1890 VNB.n655 VNB.n652 121.366
R1891 VNB.n702 VNB.n701 121.366
R1892 VNB.n761 VNB.n760 121.366
R1893 VNB.n956 VNB.n955 121.366
R1894 VNB.n1043 VNB.n1040 121.366
R1895 VNB.n39 VNB.n38 121.366
R1896 VNB.n459 VNB.n458 85.559
R1897 VNB.n527 VNB.n526 85.559
R1898 VNB.n840 VNB.n839 85.559
R1899 VNB.n908 VNB.n907 85.559
R1900 VNB.n1214 VNB.n1213 85.559
R1901 VNB.n1282 VNB.n1281 85.559
R1902 VNB.n205 VNB.n204 84.842
R1903 VNB.n332 VNB.n331 84.842
R1904 VNB.n579 VNB.n578 84.842
R1905 VNB.n1094 VNB.n1093 84.842
R1906 VNB.n1146 VNB.n1145 84.842
R1907 VNB.n1294 VNB.n1293 76
R1908 VNB.n1290 VNB.n1289 76
R1909 VNB.n1286 VNB.n1285 76
R1910 VNB.n1280 VNB.n1279 76
R1911 VNB.n1276 VNB.n1275 76
R1912 VNB.n1272 VNB.n1271 76
R1913 VNB.n1268 VNB.n1267 76
R1914 VNB.n1264 VNB.n1263 76
R1915 VNB.n1260 VNB.n1259 76
R1916 VNB.n1256 VNB.n1255 76
R1917 VNB.n1252 VNB.n1251 76
R1918 VNB.n1248 VNB.n1247 76
R1919 VNB.n1226 VNB.n1225 76
R1920 VNB.n1222 VNB.n1221 76
R1921 VNB.n1218 VNB.n1217 76
R1922 VNB.n1212 VNB.n1211 76
R1923 VNB.n1208 VNB.n1207 76
R1924 VNB.n1204 VNB.n1203 76
R1925 VNB.n1200 VNB.n1199 76
R1926 VNB.n1196 VNB.n1195 76
R1927 VNB.n1192 VNB.n1191 76
R1928 VNB.n1188 VNB.n1187 76
R1929 VNB.n1184 VNB.n1183 76
R1930 VNB.n1180 VNB.n1179 76
R1931 VNB.n1158 VNB.n1157 76
R1932 VNB.n1154 VNB.n1153 76
R1933 VNB.n1150 VNB.n1149 76
R1934 VNB.n1144 VNB.n1143 76
R1935 VNB.n1140 VNB.n1139 76
R1936 VNB.n1136 VNB.n1135 76
R1937 VNB.n1132 VNB.n1131 76
R1938 VNB.n1128 VNB.n1127 76
R1939 VNB.n1106 VNB.n1105 76
R1940 VNB.n1102 VNB.n1101 76
R1941 VNB.n1098 VNB.n1097 76
R1942 VNB.n1092 VNB.n1091 76
R1943 VNB.n1088 VNB.n1087 76
R1944 VNB.n1084 VNB.n1083 76
R1945 VNB.n1080 VNB.n1079 76
R1946 VNB.n1076 VNB.n1075 76
R1947 VNB.n1054 VNB.n1053 76
R1948 VNB.n1050 VNB.n1049 76
R1949 VNB.n1046 VNB.n1045 76
R1950 VNB.n1034 VNB.n1033 76
R1951 VNB.n1029 VNB.n1028 76
R1952 VNB.n1025 VNB.n1024 76
R1953 VNB.n1021 VNB.n1020 76
R1954 VNB.n1017 VNB.n1016 76
R1955 VNB.n1013 VNB.n1012 76
R1956 VNB.n1009 VNB.n1008 76
R1957 VNB.n1005 VNB.n1004 76
R1958 VNB.n1001 VNB.n1000 76
R1959 VNB.n979 VNB.n978 76
R1960 VNB.n975 VNB.n974 76
R1961 VNB.n971 VNB.n970 76
R1962 VNB.n960 VNB.n959 76
R1963 VNB.n954 VNB.n953 76
R1964 VNB.n950 VNB.n949 76
R1965 VNB.n946 VNB.n945 76
R1966 VNB.n942 VNB.n941 76
R1967 VNB.n920 VNB.n919 76
R1968 VNB.n916 VNB.n915 76
R1969 VNB.n912 VNB.n911 76
R1970 VNB.n906 VNB.n905 76
R1971 VNB.n902 VNB.n901 76
R1972 VNB.n898 VNB.n897 76
R1973 VNB.n894 VNB.n893 76
R1974 VNB.n890 VNB.n889 76
R1975 VNB.n886 VNB.n885 76
R1976 VNB.n882 VNB.n881 76
R1977 VNB.n878 VNB.n877 76
R1978 VNB.n874 VNB.n873 76
R1979 VNB.n852 VNB.n851 76
R1980 VNB.n848 VNB.n847 76
R1981 VNB.n844 VNB.n843 76
R1982 VNB.n838 VNB.n837 76
R1983 VNB.n834 VNB.n833 76
R1984 VNB.n830 VNB.n829 76
R1985 VNB.n826 VNB.n825 76
R1986 VNB.n822 VNB.n821 76
R1987 VNB.n818 VNB.n817 76
R1988 VNB.n814 VNB.n813 76
R1989 VNB.n810 VNB.n809 76
R1990 VNB.n806 VNB.n805 76
R1991 VNB.n784 VNB.n783 76
R1992 VNB.n780 VNB.n779 76
R1993 VNB.n776 VNB.n775 76
R1994 VNB.n765 VNB.n764 76
R1995 VNB.n759 VNB.n758 76
R1996 VNB.n755 VNB.n754 76
R1997 VNB.n751 VNB.n750 76
R1998 VNB.n747 VNB.n746 76
R1999 VNB.n725 VNB.n724 76
R2000 VNB.n721 VNB.n720 76
R2001 VNB.n717 VNB.n716 76
R2002 VNB.n706 VNB.n705 76
R2003 VNB.n700 VNB.n699 76
R2004 VNB.n696 VNB.n695 76
R2005 VNB.n692 VNB.n691 76
R2006 VNB.n688 VNB.n687 76
R2007 VNB.n666 VNB.n665 76
R2008 VNB.n662 VNB.n661 76
R2009 VNB.n658 VNB.n657 76
R2010 VNB.n646 VNB.n645 76
R2011 VNB.n641 VNB.n640 76
R2012 VNB.n637 VNB.n636 76
R2013 VNB.n633 VNB.n632 76
R2014 VNB.n629 VNB.n628 76
R2015 VNB.n625 VNB.n624 76
R2016 VNB.n621 VNB.n620 76
R2017 VNB.n617 VNB.n616 76
R2018 VNB.n613 VNB.n612 76
R2019 VNB.n591 VNB.n590 76
R2020 VNB.n587 VNB.n586 76
R2021 VNB.n583 VNB.n582 76
R2022 VNB.n577 VNB.n576 76
R2023 VNB.n573 VNB.n572 76
R2024 VNB.n569 VNB.n568 76
R2025 VNB.n565 VNB.n564 76
R2026 VNB.n561 VNB.n560 76
R2027 VNB.n539 VNB.n538 76
R2028 VNB.n535 VNB.n534 76
R2029 VNB.n531 VNB.n530 76
R2030 VNB.n525 VNB.n524 76
R2031 VNB.n521 VNB.n520 76
R2032 VNB.n517 VNB.n516 76
R2033 VNB.n513 VNB.n512 76
R2034 VNB.n509 VNB.n508 76
R2035 VNB.n505 VNB.n504 76
R2036 VNB.n501 VNB.n500 76
R2037 VNB.n497 VNB.n496 76
R2038 VNB.n493 VNB.n492 76
R2039 VNB.n471 VNB.n470 76
R2040 VNB.n467 VNB.n466 76
R2041 VNB.n463 VNB.n462 76
R2042 VNB.n457 VNB.n456 76
R2043 VNB.n453 VNB.n452 76
R2044 VNB.n449 VNB.n448 76
R2045 VNB.n445 VNB.n444 76
R2046 VNB.n441 VNB.n440 76
R2047 VNB.n437 VNB.n436 76
R2048 VNB.n433 VNB.n432 76
R2049 VNB.n429 VNB.n428 76
R2050 VNB.n425 VNB.n424 76
R2051 VNB.n403 VNB.n402 76
R2052 VNB.n399 VNB.n398 76
R2053 VNB.n395 VNB.n394 76
R2054 VNB.n384 VNB.n383 76
R2055 VNB.n378 VNB.n377 76
R2056 VNB.n374 VNB.n373 76
R2057 VNB.n370 VNB.n369 76
R2058 VNB.n366 VNB.n365 76
R2059 VNB.n344 VNB.n343 76
R2060 VNB.n340 VNB.n339 76
R2061 VNB.n336 VNB.n335 76
R2062 VNB.n330 VNB.n329 76
R2063 VNB.n326 VNB.n325 76
R2064 VNB.n322 VNB.n321 76
R2065 VNB.n318 VNB.n317 76
R2066 VNB.n314 VNB.n313 76
R2067 VNB.n292 VNB.n291 76
R2068 VNB.n288 VNB.n287 76
R2069 VNB.n284 VNB.n283 76
R2070 VNB.n272 VNB.n271 76
R2071 VNB.n267 VNB.n266 76
R2072 VNB.n263 VNB.n262 76
R2073 VNB.n259 VNB.n258 76
R2074 VNB.n255 VNB.n254 76
R2075 VNB.n251 VNB.n250 76
R2076 VNB.n247 VNB.n246 76
R2077 VNB.n243 VNB.n242 76
R2078 VNB.n239 VNB.n238 76
R2079 VNB.n217 VNB.n216 76
R2080 VNB.n213 VNB.n212 76
R2081 VNB.n209 VNB.n208 76
R2082 VNB.n203 VNB.n202 76
R2083 VNB.n199 VNB.n198 76
R2084 VNB.n195 VNB.n194 76
R2085 VNB.n191 VNB.n190 76
R2086 VNB.n187 VNB.n186 76
R2087 VNB.n165 VNB.n164 76
R2088 VNB.n161 VNB.n160 76
R2089 VNB.n157 VNB.n156 76
R2090 VNB.n146 VNB.n145 76
R2091 VNB.n140 VNB.n139 76
R2092 VNB.n136 VNB.n135 76
R2093 VNB.n132 VNB.n131 76
R2094 VNB.n128 VNB.n127 76
R2095 VNB.n106 VNB.n105 76
R2096 VNB.n102 VNB.n101 76
R2097 VNB.n98 VNB.n97 76
R2098 VNB.n87 VNB.n86 76
R2099 VNB.n277 VNB.n276 64.552
R2100 VNB.n651 VNB.n650 64.552
R2101 VNB.n1039 VNB.n1038 64.552
R2102 VNB.n92 VNB.n91 63.835
R2103 VNB.n151 VNB.n150 63.835
R2104 VNB.n389 VNB.n388 63.835
R2105 VNB.n711 VNB.n710 63.835
R2106 VNB.n770 VNB.n769 63.835
R2107 VNB.n965 VNB.n964 63.835
R2108 VNB.n43 VNB.n7 63.835
R2109 VNB.n461 VNB.n460 41.971
R2110 VNB.n529 VNB.n528 41.971
R2111 VNB.n842 VNB.n841 41.971
R2112 VNB.n910 VNB.n909 41.971
R2113 VNB.n1216 VNB.n1215 41.971
R2114 VNB.n1284 VNB.n1283 41.971
R2115 VNB.n84 VNB.n83 36.937
R2116 VNB.n143 VNB.n142 36.937
R2117 VNB.n281 VNB.n280 36.937
R2118 VNB.n381 VNB.n380 36.937
R2119 VNB.n655 VNB.n654 36.937
R2120 VNB.n703 VNB.n702 36.937
R2121 VNB.n762 VNB.n761 36.937
R2122 VNB.n957 VNB.n956 36.937
R2123 VNB.n1043 VNB.n1042 36.937
R2124 VNB.n40 VNB.n39 36.937
R2125 VNB.n207 VNB.n206 36.678
R2126 VNB.n334 VNB.n333 36.678
R2127 VNB.n581 VNB.n580 36.678
R2128 VNB.n1096 VNB.n1095 36.678
R2129 VNB.n1148 VNB.n1147 36.678
R2130 VNB.n80 VNB.n79 35.118
R2131 VNB.n1301 VNB.n1300 35.118
R2132 VNB.n280 VNB.n279 29.844
R2133 VNB.n654 VNB.n653 29.844
R2134 VNB.n1042 VNB.n1041 29.844
R2135 VNB.n91 VNB.n90 28.421
R2136 VNB.n150 VNB.n149 28.421
R2137 VNB.n276 VNB.n275 28.421
R2138 VNB.n388 VNB.n387 28.421
R2139 VNB.n650 VNB.n649 28.421
R2140 VNB.n710 VNB.n709 28.421
R2141 VNB.n769 VNB.n768 28.421
R2142 VNB.n964 VNB.n963 28.421
R2143 VNB.n1038 VNB.n1037 28.421
R2144 VNB.n7 VNB.n6 28.421
R2145 VNB.n95 VNB.n94 27.855
R2146 VNB.n154 VNB.n153 27.855
R2147 VNB.n392 VNB.n391 27.855
R2148 VNB.n714 VNB.n713 27.855
R2149 VNB.n773 VNB.n772 27.855
R2150 VNB.n968 VNB.n967 27.855
R2151 VNB.n46 VNB.n45 27.855
R2152 VNB.n91 VNB.n89 25.263
R2153 VNB.n150 VNB.n148 25.263
R2154 VNB.n276 VNB.n274 25.263
R2155 VNB.n388 VNB.n386 25.263
R2156 VNB.n650 VNB.n648 25.263
R2157 VNB.n710 VNB.n708 25.263
R2158 VNB.n769 VNB.n767 25.263
R2159 VNB.n964 VNB.n962 25.263
R2160 VNB.n1038 VNB.n1036 25.263
R2161 VNB.n7 VNB.n5 25.263
R2162 VNB.n89 VNB.n88 24.383
R2163 VNB.n148 VNB.n147 24.383
R2164 VNB.n274 VNB.n273 24.383
R2165 VNB.n386 VNB.n385 24.383
R2166 VNB.n648 VNB.n647 24.383
R2167 VNB.n708 VNB.n707 24.383
R2168 VNB.n767 VNB.n766 24.383
R2169 VNB.n962 VNB.n961 24.383
R2170 VNB.n1036 VNB.n1035 24.383
R2171 VNB.n5 VNB.n4 24.383
R2172 VNB.n69 VNB.n66 20.452
R2173 VNB.n1303 VNB.n1302 20.452
R2174 VNB.n96 VNB.n95 16.721
R2175 VNB.n155 VNB.n154 16.721
R2176 VNB.n393 VNB.n392 16.721
R2177 VNB.n715 VNB.n714 16.721
R2178 VNB.n774 VNB.n773 16.721
R2179 VNB.n969 VNB.n968 16.721
R2180 VNB.n47 VNB.n46 16.721
R2181 VNB.n78 VNB.n77 13.653
R2182 VNB.n77 VNB.n76 13.653
R2183 VNB.n75 VNB.n74 13.653
R2184 VNB.n74 VNB.n73 13.653
R2185 VNB.n72 VNB.n71 13.653
R2186 VNB.n71 VNB.n70 13.653
R2187 VNB.n86 VNB.n85 13.653
R2188 VNB.n85 VNB.n84 13.653
R2189 VNB.n97 VNB.n96 13.653
R2190 VNB.n101 VNB.n100 13.653
R2191 VNB.n100 VNB.n99 13.653
R2192 VNB.n105 VNB.n104 13.653
R2193 VNB.n104 VNB.n103 13.653
R2194 VNB.n127 VNB.n126 13.653
R2195 VNB.n126 VNB.n125 13.653
R2196 VNB.n131 VNB.n130 13.653
R2197 VNB.n130 VNB.n129 13.653
R2198 VNB.n135 VNB.n134 13.653
R2199 VNB.n134 VNB.n133 13.653
R2200 VNB.n139 VNB.n138 13.653
R2201 VNB.n138 VNB.n137 13.653
R2202 VNB.n145 VNB.n144 13.653
R2203 VNB.n144 VNB.n143 13.653
R2204 VNB.n156 VNB.n155 13.653
R2205 VNB.n160 VNB.n159 13.653
R2206 VNB.n159 VNB.n158 13.653
R2207 VNB.n164 VNB.n163 13.653
R2208 VNB.n163 VNB.n162 13.653
R2209 VNB.n186 VNB.n185 13.653
R2210 VNB.n185 VNB.n184 13.653
R2211 VNB.n190 VNB.n189 13.653
R2212 VNB.n189 VNB.n188 13.653
R2213 VNB.n194 VNB.n193 13.653
R2214 VNB.n193 VNB.n192 13.653
R2215 VNB.n198 VNB.n197 13.653
R2216 VNB.n197 VNB.n196 13.653
R2217 VNB.n202 VNB.n201 13.653
R2218 VNB.n201 VNB.n200 13.653
R2219 VNB.n208 VNB.n207 13.653
R2220 VNB.n212 VNB.n211 13.653
R2221 VNB.n211 VNB.n210 13.653
R2222 VNB.n216 VNB.n215 13.653
R2223 VNB.n215 VNB.n214 13.653
R2224 VNB.n238 VNB.n237 13.653
R2225 VNB.n237 VNB.n236 13.653
R2226 VNB.n242 VNB.n241 13.653
R2227 VNB.n241 VNB.n240 13.653
R2228 VNB.n246 VNB.n245 13.653
R2229 VNB.n245 VNB.n244 13.653
R2230 VNB.n250 VNB.n249 13.653
R2231 VNB.n249 VNB.n248 13.653
R2232 VNB.n254 VNB.n253 13.653
R2233 VNB.n253 VNB.n252 13.653
R2234 VNB.n258 VNB.n257 13.653
R2235 VNB.n257 VNB.n256 13.653
R2236 VNB.n262 VNB.n261 13.653
R2237 VNB.n261 VNB.n260 13.653
R2238 VNB.n266 VNB.n265 13.653
R2239 VNB.n265 VNB.n264 13.653
R2240 VNB.n271 VNB.n270 13.653
R2241 VNB.n270 VNB.n269 13.653
R2242 VNB.n283 VNB.n282 13.653
R2243 VNB.n282 VNB.n281 13.653
R2244 VNB.n287 VNB.n286 13.653
R2245 VNB.n286 VNB.n285 13.653
R2246 VNB.n291 VNB.n290 13.653
R2247 VNB.n290 VNB.n289 13.653
R2248 VNB.n313 VNB.n312 13.653
R2249 VNB.n312 VNB.n311 13.653
R2250 VNB.n317 VNB.n316 13.653
R2251 VNB.n316 VNB.n315 13.653
R2252 VNB.n321 VNB.n320 13.653
R2253 VNB.n320 VNB.n319 13.653
R2254 VNB.n325 VNB.n324 13.653
R2255 VNB.n324 VNB.n323 13.653
R2256 VNB.n329 VNB.n328 13.653
R2257 VNB.n328 VNB.n327 13.653
R2258 VNB.n335 VNB.n334 13.653
R2259 VNB.n339 VNB.n338 13.653
R2260 VNB.n338 VNB.n337 13.653
R2261 VNB.n343 VNB.n342 13.653
R2262 VNB.n342 VNB.n341 13.653
R2263 VNB.n365 VNB.n364 13.653
R2264 VNB.n364 VNB.n363 13.653
R2265 VNB.n369 VNB.n368 13.653
R2266 VNB.n368 VNB.n367 13.653
R2267 VNB.n373 VNB.n372 13.653
R2268 VNB.n372 VNB.n371 13.653
R2269 VNB.n377 VNB.n376 13.653
R2270 VNB.n376 VNB.n375 13.653
R2271 VNB.n383 VNB.n382 13.653
R2272 VNB.n382 VNB.n381 13.653
R2273 VNB.n394 VNB.n393 13.653
R2274 VNB.n398 VNB.n397 13.653
R2275 VNB.n397 VNB.n396 13.653
R2276 VNB.n402 VNB.n401 13.653
R2277 VNB.n401 VNB.n400 13.653
R2278 VNB.n424 VNB.n423 13.653
R2279 VNB.n423 VNB.n422 13.653
R2280 VNB.n428 VNB.n427 13.653
R2281 VNB.n427 VNB.n426 13.653
R2282 VNB.n432 VNB.n431 13.653
R2283 VNB.n431 VNB.n430 13.653
R2284 VNB.n436 VNB.n435 13.653
R2285 VNB.n435 VNB.n434 13.653
R2286 VNB.n440 VNB.n439 13.653
R2287 VNB.n439 VNB.n438 13.653
R2288 VNB.n444 VNB.n443 13.653
R2289 VNB.n443 VNB.n442 13.653
R2290 VNB.n448 VNB.n447 13.653
R2291 VNB.n447 VNB.n446 13.653
R2292 VNB.n452 VNB.n451 13.653
R2293 VNB.n451 VNB.n450 13.653
R2294 VNB.n456 VNB.n455 13.653
R2295 VNB.n455 VNB.n454 13.653
R2296 VNB.n462 VNB.n461 13.653
R2297 VNB.n466 VNB.n465 13.653
R2298 VNB.n465 VNB.n464 13.653
R2299 VNB.n470 VNB.n469 13.653
R2300 VNB.n469 VNB.n468 13.653
R2301 VNB.n492 VNB.n491 13.653
R2302 VNB.n491 VNB.n490 13.653
R2303 VNB.n496 VNB.n495 13.653
R2304 VNB.n495 VNB.n494 13.653
R2305 VNB.n500 VNB.n499 13.653
R2306 VNB.n499 VNB.n498 13.653
R2307 VNB.n504 VNB.n503 13.653
R2308 VNB.n503 VNB.n502 13.653
R2309 VNB.n508 VNB.n507 13.653
R2310 VNB.n507 VNB.n506 13.653
R2311 VNB.n512 VNB.n511 13.653
R2312 VNB.n511 VNB.n510 13.653
R2313 VNB.n516 VNB.n515 13.653
R2314 VNB.n515 VNB.n514 13.653
R2315 VNB.n520 VNB.n519 13.653
R2316 VNB.n519 VNB.n518 13.653
R2317 VNB.n524 VNB.n523 13.653
R2318 VNB.n523 VNB.n522 13.653
R2319 VNB.n530 VNB.n529 13.653
R2320 VNB.n534 VNB.n533 13.653
R2321 VNB.n533 VNB.n532 13.653
R2322 VNB.n538 VNB.n537 13.653
R2323 VNB.n537 VNB.n536 13.653
R2324 VNB.n560 VNB.n559 13.653
R2325 VNB.n559 VNB.n558 13.653
R2326 VNB.n564 VNB.n563 13.653
R2327 VNB.n563 VNB.n562 13.653
R2328 VNB.n568 VNB.n567 13.653
R2329 VNB.n567 VNB.n566 13.653
R2330 VNB.n572 VNB.n571 13.653
R2331 VNB.n571 VNB.n570 13.653
R2332 VNB.n576 VNB.n575 13.653
R2333 VNB.n575 VNB.n574 13.653
R2334 VNB.n582 VNB.n581 13.653
R2335 VNB.n586 VNB.n585 13.653
R2336 VNB.n585 VNB.n584 13.653
R2337 VNB.n590 VNB.n589 13.653
R2338 VNB.n589 VNB.n588 13.653
R2339 VNB.n612 VNB.n611 13.653
R2340 VNB.n611 VNB.n610 13.653
R2341 VNB.n616 VNB.n615 13.653
R2342 VNB.n615 VNB.n614 13.653
R2343 VNB.n620 VNB.n619 13.653
R2344 VNB.n619 VNB.n618 13.653
R2345 VNB.n624 VNB.n623 13.653
R2346 VNB.n623 VNB.n622 13.653
R2347 VNB.n628 VNB.n627 13.653
R2348 VNB.n627 VNB.n626 13.653
R2349 VNB.n632 VNB.n631 13.653
R2350 VNB.n631 VNB.n630 13.653
R2351 VNB.n636 VNB.n635 13.653
R2352 VNB.n635 VNB.n634 13.653
R2353 VNB.n640 VNB.n639 13.653
R2354 VNB.n639 VNB.n638 13.653
R2355 VNB.n645 VNB.n644 13.653
R2356 VNB.n644 VNB.n643 13.653
R2357 VNB.n657 VNB.n656 13.653
R2358 VNB.n656 VNB.n655 13.653
R2359 VNB.n661 VNB.n660 13.653
R2360 VNB.n660 VNB.n659 13.653
R2361 VNB.n665 VNB.n664 13.653
R2362 VNB.n664 VNB.n663 13.653
R2363 VNB.n687 VNB.n686 13.653
R2364 VNB.n686 VNB.n685 13.653
R2365 VNB.n691 VNB.n690 13.653
R2366 VNB.n690 VNB.n689 13.653
R2367 VNB.n695 VNB.n694 13.653
R2368 VNB.n694 VNB.n693 13.653
R2369 VNB.n699 VNB.n698 13.653
R2370 VNB.n698 VNB.n697 13.653
R2371 VNB.n705 VNB.n704 13.653
R2372 VNB.n704 VNB.n703 13.653
R2373 VNB.n716 VNB.n715 13.653
R2374 VNB.n720 VNB.n719 13.653
R2375 VNB.n719 VNB.n718 13.653
R2376 VNB.n724 VNB.n723 13.653
R2377 VNB.n723 VNB.n722 13.653
R2378 VNB.n746 VNB.n745 13.653
R2379 VNB.n745 VNB.n744 13.653
R2380 VNB.n750 VNB.n749 13.653
R2381 VNB.n749 VNB.n748 13.653
R2382 VNB.n754 VNB.n753 13.653
R2383 VNB.n753 VNB.n752 13.653
R2384 VNB.n758 VNB.n757 13.653
R2385 VNB.n757 VNB.n756 13.653
R2386 VNB.n764 VNB.n763 13.653
R2387 VNB.n763 VNB.n762 13.653
R2388 VNB.n775 VNB.n774 13.653
R2389 VNB.n779 VNB.n778 13.653
R2390 VNB.n778 VNB.n777 13.653
R2391 VNB.n783 VNB.n782 13.653
R2392 VNB.n782 VNB.n781 13.653
R2393 VNB.n805 VNB.n804 13.653
R2394 VNB.n804 VNB.n803 13.653
R2395 VNB.n809 VNB.n808 13.653
R2396 VNB.n808 VNB.n807 13.653
R2397 VNB.n813 VNB.n812 13.653
R2398 VNB.n812 VNB.n811 13.653
R2399 VNB.n817 VNB.n816 13.653
R2400 VNB.n816 VNB.n815 13.653
R2401 VNB.n821 VNB.n820 13.653
R2402 VNB.n820 VNB.n819 13.653
R2403 VNB.n825 VNB.n824 13.653
R2404 VNB.n824 VNB.n823 13.653
R2405 VNB.n829 VNB.n828 13.653
R2406 VNB.n828 VNB.n827 13.653
R2407 VNB.n833 VNB.n832 13.653
R2408 VNB.n832 VNB.n831 13.653
R2409 VNB.n837 VNB.n836 13.653
R2410 VNB.n836 VNB.n835 13.653
R2411 VNB.n843 VNB.n842 13.653
R2412 VNB.n847 VNB.n846 13.653
R2413 VNB.n846 VNB.n845 13.653
R2414 VNB.n851 VNB.n850 13.653
R2415 VNB.n850 VNB.n849 13.653
R2416 VNB.n873 VNB.n872 13.653
R2417 VNB.n872 VNB.n871 13.653
R2418 VNB.n877 VNB.n876 13.653
R2419 VNB.n876 VNB.n875 13.653
R2420 VNB.n881 VNB.n880 13.653
R2421 VNB.n880 VNB.n879 13.653
R2422 VNB.n885 VNB.n884 13.653
R2423 VNB.n884 VNB.n883 13.653
R2424 VNB.n889 VNB.n888 13.653
R2425 VNB.n888 VNB.n887 13.653
R2426 VNB.n893 VNB.n892 13.653
R2427 VNB.n892 VNB.n891 13.653
R2428 VNB.n897 VNB.n896 13.653
R2429 VNB.n896 VNB.n895 13.653
R2430 VNB.n901 VNB.n900 13.653
R2431 VNB.n900 VNB.n899 13.653
R2432 VNB.n905 VNB.n904 13.653
R2433 VNB.n904 VNB.n903 13.653
R2434 VNB.n911 VNB.n910 13.653
R2435 VNB.n915 VNB.n914 13.653
R2436 VNB.n914 VNB.n913 13.653
R2437 VNB.n919 VNB.n918 13.653
R2438 VNB.n918 VNB.n917 13.653
R2439 VNB.n941 VNB.n940 13.653
R2440 VNB.n940 VNB.n939 13.653
R2441 VNB.n945 VNB.n944 13.653
R2442 VNB.n944 VNB.n943 13.653
R2443 VNB.n949 VNB.n948 13.653
R2444 VNB.n948 VNB.n947 13.653
R2445 VNB.n953 VNB.n952 13.653
R2446 VNB.n952 VNB.n951 13.653
R2447 VNB.n959 VNB.n958 13.653
R2448 VNB.n958 VNB.n957 13.653
R2449 VNB.n970 VNB.n969 13.653
R2450 VNB.n974 VNB.n973 13.653
R2451 VNB.n973 VNB.n972 13.653
R2452 VNB.n978 VNB.n977 13.653
R2453 VNB.n977 VNB.n976 13.653
R2454 VNB.n1000 VNB.n999 13.653
R2455 VNB.n999 VNB.n998 13.653
R2456 VNB.n1004 VNB.n1003 13.653
R2457 VNB.n1003 VNB.n1002 13.653
R2458 VNB.n1008 VNB.n1007 13.653
R2459 VNB.n1007 VNB.n1006 13.653
R2460 VNB.n1012 VNB.n1011 13.653
R2461 VNB.n1011 VNB.n1010 13.653
R2462 VNB.n1016 VNB.n1015 13.653
R2463 VNB.n1015 VNB.n1014 13.653
R2464 VNB.n1020 VNB.n1019 13.653
R2465 VNB.n1019 VNB.n1018 13.653
R2466 VNB.n1024 VNB.n1023 13.653
R2467 VNB.n1023 VNB.n1022 13.653
R2468 VNB.n1028 VNB.n1027 13.653
R2469 VNB.n1027 VNB.n1026 13.653
R2470 VNB.n1033 VNB.n1032 13.653
R2471 VNB.n1032 VNB.n1031 13.653
R2472 VNB.n1045 VNB.n1044 13.653
R2473 VNB.n1044 VNB.n1043 13.653
R2474 VNB.n1049 VNB.n1048 13.653
R2475 VNB.n1048 VNB.n1047 13.653
R2476 VNB.n1053 VNB.n1052 13.653
R2477 VNB.n1052 VNB.n1051 13.653
R2478 VNB.n1075 VNB.n1074 13.653
R2479 VNB.n1074 VNB.n1073 13.653
R2480 VNB.n1079 VNB.n1078 13.653
R2481 VNB.n1078 VNB.n1077 13.653
R2482 VNB.n1083 VNB.n1082 13.653
R2483 VNB.n1082 VNB.n1081 13.653
R2484 VNB.n1087 VNB.n1086 13.653
R2485 VNB.n1086 VNB.n1085 13.653
R2486 VNB.n1091 VNB.n1090 13.653
R2487 VNB.n1090 VNB.n1089 13.653
R2488 VNB.n1097 VNB.n1096 13.653
R2489 VNB.n1101 VNB.n1100 13.653
R2490 VNB.n1100 VNB.n1099 13.653
R2491 VNB.n1105 VNB.n1104 13.653
R2492 VNB.n1104 VNB.n1103 13.653
R2493 VNB.n1127 VNB.n1126 13.653
R2494 VNB.n1126 VNB.n1125 13.653
R2495 VNB.n1131 VNB.n1130 13.653
R2496 VNB.n1130 VNB.n1129 13.653
R2497 VNB.n1135 VNB.n1134 13.653
R2498 VNB.n1134 VNB.n1133 13.653
R2499 VNB.n1139 VNB.n1138 13.653
R2500 VNB.n1138 VNB.n1137 13.653
R2501 VNB.n1143 VNB.n1142 13.653
R2502 VNB.n1142 VNB.n1141 13.653
R2503 VNB.n1149 VNB.n1148 13.653
R2504 VNB.n1153 VNB.n1152 13.653
R2505 VNB.n1152 VNB.n1151 13.653
R2506 VNB.n1157 VNB.n1156 13.653
R2507 VNB.n1156 VNB.n1155 13.653
R2508 VNB.n1179 VNB.n1178 13.653
R2509 VNB.n1178 VNB.n1177 13.653
R2510 VNB.n1183 VNB.n1182 13.653
R2511 VNB.n1182 VNB.n1181 13.653
R2512 VNB.n1187 VNB.n1186 13.653
R2513 VNB.n1186 VNB.n1185 13.653
R2514 VNB.n1191 VNB.n1190 13.653
R2515 VNB.n1190 VNB.n1189 13.653
R2516 VNB.n1195 VNB.n1194 13.653
R2517 VNB.n1194 VNB.n1193 13.653
R2518 VNB.n1199 VNB.n1198 13.653
R2519 VNB.n1198 VNB.n1197 13.653
R2520 VNB.n1203 VNB.n1202 13.653
R2521 VNB.n1202 VNB.n1201 13.653
R2522 VNB.n1207 VNB.n1206 13.653
R2523 VNB.n1206 VNB.n1205 13.653
R2524 VNB.n1211 VNB.n1210 13.653
R2525 VNB.n1210 VNB.n1209 13.653
R2526 VNB.n1217 VNB.n1216 13.653
R2527 VNB.n1221 VNB.n1220 13.653
R2528 VNB.n1220 VNB.n1219 13.653
R2529 VNB.n1225 VNB.n1224 13.653
R2530 VNB.n1224 VNB.n1223 13.653
R2531 VNB.n1247 VNB.n1246 13.653
R2532 VNB.n1246 VNB.n1245 13.653
R2533 VNB.n1251 VNB.n1250 13.653
R2534 VNB.n1250 VNB.n1249 13.653
R2535 VNB.n1255 VNB.n1254 13.653
R2536 VNB.n1254 VNB.n1253 13.653
R2537 VNB.n1259 VNB.n1258 13.653
R2538 VNB.n1258 VNB.n1257 13.653
R2539 VNB.n1263 VNB.n1262 13.653
R2540 VNB.n1262 VNB.n1261 13.653
R2541 VNB.n1267 VNB.n1266 13.653
R2542 VNB.n1266 VNB.n1265 13.653
R2543 VNB.n1271 VNB.n1270 13.653
R2544 VNB.n1270 VNB.n1269 13.653
R2545 VNB.n1275 VNB.n1274 13.653
R2546 VNB.n1274 VNB.n1273 13.653
R2547 VNB.n1279 VNB.n1278 13.653
R2548 VNB.n1278 VNB.n1277 13.653
R2549 VNB.n1285 VNB.n1284 13.653
R2550 VNB.n1289 VNB.n1288 13.653
R2551 VNB.n1288 VNB.n1287 13.653
R2552 VNB.n1293 VNB.n1292 13.653
R2553 VNB.n1292 VNB.n1291 13.653
R2554 VNB.n28 VNB.n27 13.653
R2555 VNB.n27 VNB.n26 13.653
R2556 VNB.n31 VNB.n30 13.653
R2557 VNB.n30 VNB.n29 13.653
R2558 VNB.n34 VNB.n33 13.653
R2559 VNB.n33 VNB.n32 13.653
R2560 VNB.n37 VNB.n36 13.653
R2561 VNB.n36 VNB.n35 13.653
R2562 VNB.n42 VNB.n41 13.653
R2563 VNB.n41 VNB.n40 13.653
R2564 VNB.n48 VNB.n47 13.653
R2565 VNB.n51 VNB.n50 13.653
R2566 VNB.n50 VNB.n49 13.653
R2567 VNB.n1302 VNB.n0 13.653
R2568 VNB VNB.n0 13.653
R2569 VNB.n69 VNB.n68 13.653
R2570 VNB.n68 VNB.n67 13.653
R2571 VNB.n1310 VNB.n1307 13.577
R2572 VNB.n54 VNB.n52 13.276
R2573 VNB.n66 VNB.n54 13.276
R2574 VNB.n109 VNB.n107 13.276
R2575 VNB.n122 VNB.n109 13.276
R2576 VNB.n168 VNB.n166 13.276
R2577 VNB.n181 VNB.n168 13.276
R2578 VNB.n220 VNB.n218 13.276
R2579 VNB.n233 VNB.n220 13.276
R2580 VNB.n295 VNB.n293 13.276
R2581 VNB.n308 VNB.n295 13.276
R2582 VNB.n347 VNB.n345 13.276
R2583 VNB.n360 VNB.n347 13.276
R2584 VNB.n406 VNB.n404 13.276
R2585 VNB.n419 VNB.n406 13.276
R2586 VNB.n474 VNB.n472 13.276
R2587 VNB.n487 VNB.n474 13.276
R2588 VNB.n542 VNB.n540 13.276
R2589 VNB.n555 VNB.n542 13.276
R2590 VNB.n594 VNB.n592 13.276
R2591 VNB.n607 VNB.n594 13.276
R2592 VNB.n669 VNB.n667 13.276
R2593 VNB.n682 VNB.n669 13.276
R2594 VNB.n728 VNB.n726 13.276
R2595 VNB.n741 VNB.n728 13.276
R2596 VNB.n787 VNB.n785 13.276
R2597 VNB.n800 VNB.n787 13.276
R2598 VNB.n855 VNB.n853 13.276
R2599 VNB.n868 VNB.n855 13.276
R2600 VNB.n923 VNB.n921 13.276
R2601 VNB.n936 VNB.n923 13.276
R2602 VNB.n982 VNB.n980 13.276
R2603 VNB.n995 VNB.n982 13.276
R2604 VNB.n1057 VNB.n1055 13.276
R2605 VNB.n1070 VNB.n1057 13.276
R2606 VNB.n1109 VNB.n1107 13.276
R2607 VNB.n1122 VNB.n1109 13.276
R2608 VNB.n1161 VNB.n1159 13.276
R2609 VNB.n1174 VNB.n1161 13.276
R2610 VNB.n1229 VNB.n1227 13.276
R2611 VNB.n1242 VNB.n1229 13.276
R2612 VNB.n10 VNB.n8 13.276
R2613 VNB.n23 VNB.n10 13.276
R2614 VNB.n78 VNB.n75 13.276
R2615 VNB.n75 VNB.n72 13.276
R2616 VNB.n127 VNB.n123 13.276
R2617 VNB.n186 VNB.n182 13.276
R2618 VNB.n238 VNB.n234 13.276
R2619 VNB.n313 VNB.n309 13.276
R2620 VNB.n365 VNB.n361 13.276
R2621 VNB.n424 VNB.n420 13.276
R2622 VNB.n492 VNB.n488 13.276
R2623 VNB.n560 VNB.n556 13.276
R2624 VNB.n612 VNB.n608 13.276
R2625 VNB.n687 VNB.n683 13.276
R2626 VNB.n746 VNB.n742 13.276
R2627 VNB.n805 VNB.n801 13.276
R2628 VNB.n873 VNB.n869 13.276
R2629 VNB.n941 VNB.n937 13.276
R2630 VNB.n1000 VNB.n996 13.276
R2631 VNB.n1075 VNB.n1071 13.276
R2632 VNB.n1127 VNB.n1123 13.276
R2633 VNB.n1179 VNB.n1175 13.276
R2634 VNB.n1247 VNB.n1243 13.276
R2635 VNB.n28 VNB.n24 13.276
R2636 VNB.n31 VNB.n28 13.276
R2637 VNB.n34 VNB.n31 13.276
R2638 VNB.n37 VNB.n34 13.276
R2639 VNB.n42 VNB.n37 13.276
R2640 VNB.n51 VNB.n48 13.276
R2641 VNB.n3 VNB.n1 13.276
R2642 VNB.n1303 VNB.n3 13.276
R2643 VNB.n43 VNB.n42 10.764
R2644 VNB.n1312 VNB.n1311 7.5
R2645 VNB.n115 VNB.n114 7.5
R2646 VNB.n111 VNB.n110 7.5
R2647 VNB.n109 VNB.n108 7.5
R2648 VNB.n122 VNB.n121 7.5
R2649 VNB.n174 VNB.n173 7.5
R2650 VNB.n170 VNB.n169 7.5
R2651 VNB.n168 VNB.n167 7.5
R2652 VNB.n181 VNB.n180 7.5
R2653 VNB.n226 VNB.n225 7.5
R2654 VNB.n222 VNB.n221 7.5
R2655 VNB.n220 VNB.n219 7.5
R2656 VNB.n233 VNB.n232 7.5
R2657 VNB.n301 VNB.n300 7.5
R2658 VNB.n297 VNB.n296 7.5
R2659 VNB.n295 VNB.n294 7.5
R2660 VNB.n308 VNB.n307 7.5
R2661 VNB.n353 VNB.n352 7.5
R2662 VNB.n349 VNB.n348 7.5
R2663 VNB.n347 VNB.n346 7.5
R2664 VNB.n360 VNB.n359 7.5
R2665 VNB.n412 VNB.n411 7.5
R2666 VNB.n408 VNB.n407 7.5
R2667 VNB.n406 VNB.n405 7.5
R2668 VNB.n419 VNB.n418 7.5
R2669 VNB.n480 VNB.n479 7.5
R2670 VNB.n476 VNB.n475 7.5
R2671 VNB.n474 VNB.n473 7.5
R2672 VNB.n487 VNB.n486 7.5
R2673 VNB.n548 VNB.n547 7.5
R2674 VNB.n544 VNB.n543 7.5
R2675 VNB.n542 VNB.n541 7.5
R2676 VNB.n555 VNB.n554 7.5
R2677 VNB.n600 VNB.n599 7.5
R2678 VNB.n596 VNB.n595 7.5
R2679 VNB.n594 VNB.n593 7.5
R2680 VNB.n607 VNB.n606 7.5
R2681 VNB.n675 VNB.n674 7.5
R2682 VNB.n671 VNB.n670 7.5
R2683 VNB.n669 VNB.n668 7.5
R2684 VNB.n682 VNB.n681 7.5
R2685 VNB.n734 VNB.n733 7.5
R2686 VNB.n730 VNB.n729 7.5
R2687 VNB.n728 VNB.n727 7.5
R2688 VNB.n741 VNB.n740 7.5
R2689 VNB.n793 VNB.n792 7.5
R2690 VNB.n789 VNB.n788 7.5
R2691 VNB.n787 VNB.n786 7.5
R2692 VNB.n800 VNB.n799 7.5
R2693 VNB.n861 VNB.n860 7.5
R2694 VNB.n857 VNB.n856 7.5
R2695 VNB.n855 VNB.n854 7.5
R2696 VNB.n868 VNB.n867 7.5
R2697 VNB.n929 VNB.n928 7.5
R2698 VNB.n925 VNB.n924 7.5
R2699 VNB.n923 VNB.n922 7.5
R2700 VNB.n936 VNB.n935 7.5
R2701 VNB.n988 VNB.n987 7.5
R2702 VNB.n984 VNB.n983 7.5
R2703 VNB.n982 VNB.n981 7.5
R2704 VNB.n995 VNB.n994 7.5
R2705 VNB.n1063 VNB.n1062 7.5
R2706 VNB.n1059 VNB.n1058 7.5
R2707 VNB.n1057 VNB.n1056 7.5
R2708 VNB.n1070 VNB.n1069 7.5
R2709 VNB.n1115 VNB.n1114 7.5
R2710 VNB.n1111 VNB.n1110 7.5
R2711 VNB.n1109 VNB.n1108 7.5
R2712 VNB.n1122 VNB.n1121 7.5
R2713 VNB.n1167 VNB.n1166 7.5
R2714 VNB.n1163 VNB.n1162 7.5
R2715 VNB.n1161 VNB.n1160 7.5
R2716 VNB.n1174 VNB.n1173 7.5
R2717 VNB.n1235 VNB.n1234 7.5
R2718 VNB.n1231 VNB.n1230 7.5
R2719 VNB.n1229 VNB.n1228 7.5
R2720 VNB.n1242 VNB.n1241 7.5
R2721 VNB.n16 VNB.n15 7.5
R2722 VNB.n12 VNB.n11 7.5
R2723 VNB.n10 VNB.n9 7.5
R2724 VNB.n23 VNB.n22 7.5
R2725 VNB.n1304 VNB.n1303 7.5
R2726 VNB.n3 VNB.n2 7.5
R2727 VNB.n1309 VNB.n1308 7.5
R2728 VNB.n60 VNB.n59 7.5
R2729 VNB.n56 VNB.n55 7.5
R2730 VNB.n54 VNB.n53 7.5
R2731 VNB.n66 VNB.n65 7.5
R2732 VNB.n123 VNB.n122 7.176
R2733 VNB.n182 VNB.n181 7.176
R2734 VNB.n234 VNB.n233 7.176
R2735 VNB.n309 VNB.n308 7.176
R2736 VNB.n361 VNB.n360 7.176
R2737 VNB.n420 VNB.n419 7.176
R2738 VNB.n488 VNB.n487 7.176
R2739 VNB.n556 VNB.n555 7.176
R2740 VNB.n608 VNB.n607 7.176
R2741 VNB.n683 VNB.n682 7.176
R2742 VNB.n742 VNB.n741 7.176
R2743 VNB.n801 VNB.n800 7.176
R2744 VNB.n869 VNB.n868 7.176
R2745 VNB.n937 VNB.n936 7.176
R2746 VNB.n996 VNB.n995 7.176
R2747 VNB.n1071 VNB.n1070 7.176
R2748 VNB.n1123 VNB.n1122 7.176
R2749 VNB.n1175 VNB.n1174 7.176
R2750 VNB.n1243 VNB.n1242 7.176
R2751 VNB.n24 VNB.n23 7.176
R2752 VNB.n1314 VNB.n1312 7.011
R2753 VNB.n118 VNB.n115 7.011
R2754 VNB.n113 VNB.n111 7.011
R2755 VNB.n177 VNB.n174 7.011
R2756 VNB.n172 VNB.n170 7.011
R2757 VNB.n229 VNB.n226 7.011
R2758 VNB.n224 VNB.n222 7.011
R2759 VNB.n304 VNB.n301 7.011
R2760 VNB.n299 VNB.n297 7.011
R2761 VNB.n356 VNB.n353 7.011
R2762 VNB.n351 VNB.n349 7.011
R2763 VNB.n415 VNB.n412 7.011
R2764 VNB.n410 VNB.n408 7.011
R2765 VNB.n483 VNB.n480 7.011
R2766 VNB.n478 VNB.n476 7.011
R2767 VNB.n551 VNB.n548 7.011
R2768 VNB.n546 VNB.n544 7.011
R2769 VNB.n603 VNB.n600 7.011
R2770 VNB.n598 VNB.n596 7.011
R2771 VNB.n678 VNB.n675 7.011
R2772 VNB.n673 VNB.n671 7.011
R2773 VNB.n737 VNB.n734 7.011
R2774 VNB.n732 VNB.n730 7.011
R2775 VNB.n796 VNB.n793 7.011
R2776 VNB.n791 VNB.n789 7.011
R2777 VNB.n864 VNB.n861 7.011
R2778 VNB.n859 VNB.n857 7.011
R2779 VNB.n932 VNB.n929 7.011
R2780 VNB.n927 VNB.n925 7.011
R2781 VNB.n991 VNB.n988 7.011
R2782 VNB.n986 VNB.n984 7.011
R2783 VNB.n1066 VNB.n1063 7.011
R2784 VNB.n1061 VNB.n1059 7.011
R2785 VNB.n1118 VNB.n1115 7.011
R2786 VNB.n1113 VNB.n1111 7.011
R2787 VNB.n1170 VNB.n1167 7.011
R2788 VNB.n1165 VNB.n1163 7.011
R2789 VNB.n1238 VNB.n1235 7.011
R2790 VNB.n1233 VNB.n1231 7.011
R2791 VNB.n19 VNB.n16 7.011
R2792 VNB.n14 VNB.n12 7.011
R2793 VNB.n62 VNB.n60 7.011
R2794 VNB.n58 VNB.n56 7.011
R2795 VNB.n121 VNB.n120 7.01
R2796 VNB.n113 VNB.n112 7.01
R2797 VNB.n118 VNB.n117 7.01
R2798 VNB.n180 VNB.n179 7.01
R2799 VNB.n172 VNB.n171 7.01
R2800 VNB.n177 VNB.n176 7.01
R2801 VNB.n232 VNB.n231 7.01
R2802 VNB.n224 VNB.n223 7.01
R2803 VNB.n229 VNB.n228 7.01
R2804 VNB.n307 VNB.n306 7.01
R2805 VNB.n299 VNB.n298 7.01
R2806 VNB.n304 VNB.n303 7.01
R2807 VNB.n359 VNB.n358 7.01
R2808 VNB.n351 VNB.n350 7.01
R2809 VNB.n356 VNB.n355 7.01
R2810 VNB.n418 VNB.n417 7.01
R2811 VNB.n410 VNB.n409 7.01
R2812 VNB.n415 VNB.n414 7.01
R2813 VNB.n486 VNB.n485 7.01
R2814 VNB.n478 VNB.n477 7.01
R2815 VNB.n483 VNB.n482 7.01
R2816 VNB.n554 VNB.n553 7.01
R2817 VNB.n546 VNB.n545 7.01
R2818 VNB.n551 VNB.n550 7.01
R2819 VNB.n606 VNB.n605 7.01
R2820 VNB.n598 VNB.n597 7.01
R2821 VNB.n603 VNB.n602 7.01
R2822 VNB.n681 VNB.n680 7.01
R2823 VNB.n673 VNB.n672 7.01
R2824 VNB.n678 VNB.n677 7.01
R2825 VNB.n740 VNB.n739 7.01
R2826 VNB.n732 VNB.n731 7.01
R2827 VNB.n737 VNB.n736 7.01
R2828 VNB.n799 VNB.n798 7.01
R2829 VNB.n791 VNB.n790 7.01
R2830 VNB.n796 VNB.n795 7.01
R2831 VNB.n867 VNB.n866 7.01
R2832 VNB.n859 VNB.n858 7.01
R2833 VNB.n864 VNB.n863 7.01
R2834 VNB.n935 VNB.n934 7.01
R2835 VNB.n927 VNB.n926 7.01
R2836 VNB.n932 VNB.n931 7.01
R2837 VNB.n994 VNB.n993 7.01
R2838 VNB.n986 VNB.n985 7.01
R2839 VNB.n991 VNB.n990 7.01
R2840 VNB.n1069 VNB.n1068 7.01
R2841 VNB.n1061 VNB.n1060 7.01
R2842 VNB.n1066 VNB.n1065 7.01
R2843 VNB.n1121 VNB.n1120 7.01
R2844 VNB.n1113 VNB.n1112 7.01
R2845 VNB.n1118 VNB.n1117 7.01
R2846 VNB.n1173 VNB.n1172 7.01
R2847 VNB.n1165 VNB.n1164 7.01
R2848 VNB.n1170 VNB.n1169 7.01
R2849 VNB.n1241 VNB.n1240 7.01
R2850 VNB.n1233 VNB.n1232 7.01
R2851 VNB.n1238 VNB.n1237 7.01
R2852 VNB.n22 VNB.n21 7.01
R2853 VNB.n14 VNB.n13 7.01
R2854 VNB.n19 VNB.n18 7.01
R2855 VNB.n65 VNB.n64 7.01
R2856 VNB.n58 VNB.n57 7.01
R2857 VNB.n62 VNB.n61 7.01
R2858 VNB.n1314 VNB.n1313 7.01
R2859 VNB.n1310 VNB.n1309 6.788
R2860 VNB.n1305 VNB.n1304 6.788
R2861 VNB.n79 VNB.n69 6.111
R2862 VNB.n1302 VNB.n1301 6.111
R2863 VNB.n79 VNB.n78 6.1
R2864 VNB.n1301 VNB.n51 6.1
R2865 VNB.n97 VNB.n92 2.511
R2866 VNB.n156 VNB.n151 2.511
R2867 VNB.n208 VNB.n205 2.511
R2868 VNB.n335 VNB.n332 2.511
R2869 VNB.n394 VNB.n389 2.511
R2870 VNB.n582 VNB.n579 2.511
R2871 VNB.n716 VNB.n711 2.511
R2872 VNB.n775 VNB.n770 2.511
R2873 VNB.n970 VNB.n965 2.511
R2874 VNB.n1097 VNB.n1094 2.511
R2875 VNB.n1149 VNB.n1146 2.511
R2876 VNB.n48 VNB.n43 2.511
R2877 VNB.n95 VNB.n93 1.99
R2878 VNB.n154 VNB.n152 1.99
R2879 VNB.n392 VNB.n390 1.99
R2880 VNB.n714 VNB.n712 1.99
R2881 VNB.n773 VNB.n771 1.99
R2882 VNB.n968 VNB.n966 1.99
R2883 VNB.n46 VNB.n44 1.99
R2884 VNB.n283 VNB.n277 1.255
R2885 VNB.n462 VNB.n459 1.255
R2886 VNB.n530 VNB.n527 1.255
R2887 VNB.n657 VNB.n651 1.255
R2888 VNB.n843 VNB.n840 1.255
R2889 VNB.n911 VNB.n908 1.255
R2890 VNB.n1045 VNB.n1039 1.255
R2891 VNB.n1217 VNB.n1214 1.255
R2892 VNB.n1285 VNB.n1282 1.255
R2893 VNB.n1315 VNB.n1306 0.921
R2894 VNB.n1315 VNB.n1310 0.476
R2895 VNB.n1315 VNB.n1305 0.475
R2896 VNB.n128 VNB.n106 0.272
R2897 VNB.n187 VNB.n165 0.272
R2898 VNB.n239 VNB.n217 0.272
R2899 VNB.n314 VNB.n292 0.272
R2900 VNB.n366 VNB.n344 0.272
R2901 VNB.n425 VNB.n403 0.272
R2902 VNB.n493 VNB.n471 0.272
R2903 VNB.n561 VNB.n539 0.272
R2904 VNB.n613 VNB.n591 0.272
R2905 VNB.n688 VNB.n666 0.272
R2906 VNB.n747 VNB.n725 0.272
R2907 VNB.n806 VNB.n784 0.272
R2908 VNB.n874 VNB.n852 0.272
R2909 VNB.n942 VNB.n920 0.272
R2910 VNB.n1001 VNB.n979 0.272
R2911 VNB.n1076 VNB.n1054 0.272
R2912 VNB.n1128 VNB.n1106 0.272
R2913 VNB.n1180 VNB.n1158 0.272
R2914 VNB.n1248 VNB.n1226 0.272
R2915 VNB.n1295 VNB.n1294 0.272
R2916 VNB.n119 VNB.n113 0.246
R2917 VNB.n120 VNB.n119 0.246
R2918 VNB.n119 VNB.n118 0.246
R2919 VNB.n178 VNB.n172 0.246
R2920 VNB.n179 VNB.n178 0.246
R2921 VNB.n178 VNB.n177 0.246
R2922 VNB.n230 VNB.n224 0.246
R2923 VNB.n231 VNB.n230 0.246
R2924 VNB.n230 VNB.n229 0.246
R2925 VNB.n305 VNB.n299 0.246
R2926 VNB.n306 VNB.n305 0.246
R2927 VNB.n305 VNB.n304 0.246
R2928 VNB.n357 VNB.n351 0.246
R2929 VNB.n358 VNB.n357 0.246
R2930 VNB.n357 VNB.n356 0.246
R2931 VNB.n416 VNB.n410 0.246
R2932 VNB.n417 VNB.n416 0.246
R2933 VNB.n416 VNB.n415 0.246
R2934 VNB.n484 VNB.n478 0.246
R2935 VNB.n485 VNB.n484 0.246
R2936 VNB.n484 VNB.n483 0.246
R2937 VNB.n552 VNB.n546 0.246
R2938 VNB.n553 VNB.n552 0.246
R2939 VNB.n552 VNB.n551 0.246
R2940 VNB.n604 VNB.n598 0.246
R2941 VNB.n605 VNB.n604 0.246
R2942 VNB.n604 VNB.n603 0.246
R2943 VNB.n679 VNB.n673 0.246
R2944 VNB.n680 VNB.n679 0.246
R2945 VNB.n679 VNB.n678 0.246
R2946 VNB.n738 VNB.n732 0.246
R2947 VNB.n739 VNB.n738 0.246
R2948 VNB.n738 VNB.n737 0.246
R2949 VNB.n797 VNB.n791 0.246
R2950 VNB.n798 VNB.n797 0.246
R2951 VNB.n797 VNB.n796 0.246
R2952 VNB.n865 VNB.n859 0.246
R2953 VNB.n866 VNB.n865 0.246
R2954 VNB.n865 VNB.n864 0.246
R2955 VNB.n933 VNB.n927 0.246
R2956 VNB.n934 VNB.n933 0.246
R2957 VNB.n933 VNB.n932 0.246
R2958 VNB.n992 VNB.n986 0.246
R2959 VNB.n993 VNB.n992 0.246
R2960 VNB.n992 VNB.n991 0.246
R2961 VNB.n1067 VNB.n1061 0.246
R2962 VNB.n1068 VNB.n1067 0.246
R2963 VNB.n1067 VNB.n1066 0.246
R2964 VNB.n1119 VNB.n1113 0.246
R2965 VNB.n1120 VNB.n1119 0.246
R2966 VNB.n1119 VNB.n1118 0.246
R2967 VNB.n1171 VNB.n1165 0.246
R2968 VNB.n1172 VNB.n1171 0.246
R2969 VNB.n1171 VNB.n1170 0.246
R2970 VNB.n1239 VNB.n1233 0.246
R2971 VNB.n1240 VNB.n1239 0.246
R2972 VNB.n1239 VNB.n1238 0.246
R2973 VNB.n20 VNB.n14 0.246
R2974 VNB.n21 VNB.n20 0.246
R2975 VNB.n20 VNB.n19 0.246
R2976 VNB.n63 VNB.n58 0.246
R2977 VNB.n64 VNB.n63 0.246
R2978 VNB.n63 VNB.n62 0.246
R2979 VNB.n1315 VNB.n1314 0.246
R2980 VNB.n81 VNB.n80 0.136
R2981 VNB.n87 VNB.n81 0.136
R2982 VNB.n98 VNB.n87 0.136
R2983 VNB.n102 VNB.n98 0.136
R2984 VNB.n106 VNB.n102 0.136
R2985 VNB.n132 VNB.n128 0.136
R2986 VNB.n136 VNB.n132 0.136
R2987 VNB.n140 VNB.n136 0.136
R2988 VNB.n146 VNB.n140 0.136
R2989 VNB.n157 VNB.n146 0.136
R2990 VNB.n161 VNB.n157 0.136
R2991 VNB.n165 VNB.n161 0.136
R2992 VNB.n191 VNB.n187 0.136
R2993 VNB.n195 VNB.n191 0.136
R2994 VNB.n199 VNB.n195 0.136
R2995 VNB.n203 VNB.n199 0.136
R2996 VNB.n209 VNB.n203 0.136
R2997 VNB.n213 VNB.n209 0.136
R2998 VNB.n217 VNB.n213 0.136
R2999 VNB.n243 VNB.n239 0.136
R3000 VNB.n247 VNB.n243 0.136
R3001 VNB.n251 VNB.n247 0.136
R3002 VNB.n255 VNB.n251 0.136
R3003 VNB.n259 VNB.n255 0.136
R3004 VNB.n263 VNB.n259 0.136
R3005 VNB.n267 VNB.n263 0.136
R3006 VNB.n272 VNB.n267 0.136
R3007 VNB.n284 VNB.n272 0.136
R3008 VNB.n288 VNB.n284 0.136
R3009 VNB.n292 VNB.n288 0.136
R3010 VNB.n318 VNB.n314 0.136
R3011 VNB.n322 VNB.n318 0.136
R3012 VNB.n326 VNB.n322 0.136
R3013 VNB.n330 VNB.n326 0.136
R3014 VNB.n336 VNB.n330 0.136
R3015 VNB.n340 VNB.n336 0.136
R3016 VNB.n344 VNB.n340 0.136
R3017 VNB.n370 VNB.n366 0.136
R3018 VNB.n374 VNB.n370 0.136
R3019 VNB.n378 VNB.n374 0.136
R3020 VNB.n384 VNB.n378 0.136
R3021 VNB.n395 VNB.n384 0.136
R3022 VNB.n399 VNB.n395 0.136
R3023 VNB.n403 VNB.n399 0.136
R3024 VNB.n429 VNB.n425 0.136
R3025 VNB.n433 VNB.n429 0.136
R3026 VNB.n437 VNB.n433 0.136
R3027 VNB.n441 VNB.n437 0.136
R3028 VNB.n445 VNB.n441 0.136
R3029 VNB.n449 VNB.n445 0.136
R3030 VNB.n453 VNB.n449 0.136
R3031 VNB.n457 VNB.n453 0.136
R3032 VNB.n463 VNB.n457 0.136
R3033 VNB.n467 VNB.n463 0.136
R3034 VNB.n471 VNB.n467 0.136
R3035 VNB.n497 VNB.n493 0.136
R3036 VNB.n501 VNB.n497 0.136
R3037 VNB.n505 VNB.n501 0.136
R3038 VNB.n509 VNB.n505 0.136
R3039 VNB.n513 VNB.n509 0.136
R3040 VNB.n517 VNB.n513 0.136
R3041 VNB.n521 VNB.n517 0.136
R3042 VNB.n525 VNB.n521 0.136
R3043 VNB.n531 VNB.n525 0.136
R3044 VNB.n535 VNB.n531 0.136
R3045 VNB.n539 VNB.n535 0.136
R3046 VNB.n565 VNB.n561 0.136
R3047 VNB.n569 VNB.n565 0.136
R3048 VNB.n573 VNB.n569 0.136
R3049 VNB.n577 VNB.n573 0.136
R3050 VNB.n583 VNB.n577 0.136
R3051 VNB.n587 VNB.n583 0.136
R3052 VNB.n591 VNB.n587 0.136
R3053 VNB.n617 VNB.n613 0.136
R3054 VNB.n621 VNB.n617 0.136
R3055 VNB.n625 VNB.n621 0.136
R3056 VNB.n629 VNB.n625 0.136
R3057 VNB.n633 VNB.n629 0.136
R3058 VNB.n637 VNB.n633 0.136
R3059 VNB.n641 VNB.n637 0.136
R3060 VNB.n646 VNB.n641 0.136
R3061 VNB.n658 VNB.n646 0.136
R3062 VNB.n662 VNB.n658 0.136
R3063 VNB.n666 VNB.n662 0.136
R3064 VNB.n692 VNB.n688 0.136
R3065 VNB.n696 VNB.n692 0.136
R3066 VNB.n700 VNB.n696 0.136
R3067 VNB.n706 VNB.n700 0.136
R3068 VNB.n717 VNB.n706 0.136
R3069 VNB.n721 VNB.n717 0.136
R3070 VNB.n725 VNB.n721 0.136
R3071 VNB.n751 VNB.n747 0.136
R3072 VNB.n755 VNB.n751 0.136
R3073 VNB.n759 VNB.n755 0.136
R3074 VNB.n765 VNB.n759 0.136
R3075 VNB.n776 VNB.n765 0.136
R3076 VNB.n780 VNB.n776 0.136
R3077 VNB.n784 VNB.n780 0.136
R3078 VNB.n810 VNB.n806 0.136
R3079 VNB.n814 VNB.n810 0.136
R3080 VNB.n818 VNB.n814 0.136
R3081 VNB.n822 VNB.n818 0.136
R3082 VNB.n826 VNB.n822 0.136
R3083 VNB.n830 VNB.n826 0.136
R3084 VNB.n834 VNB.n830 0.136
R3085 VNB.n838 VNB.n834 0.136
R3086 VNB.n844 VNB.n838 0.136
R3087 VNB.n848 VNB.n844 0.136
R3088 VNB.n852 VNB.n848 0.136
R3089 VNB.n878 VNB.n874 0.136
R3090 VNB.n882 VNB.n878 0.136
R3091 VNB.n886 VNB.n882 0.136
R3092 VNB.n890 VNB.n886 0.136
R3093 VNB.n894 VNB.n890 0.136
R3094 VNB.n898 VNB.n894 0.136
R3095 VNB.n902 VNB.n898 0.136
R3096 VNB.n906 VNB.n902 0.136
R3097 VNB.n912 VNB.n906 0.136
R3098 VNB.n916 VNB.n912 0.136
R3099 VNB.n920 VNB.n916 0.136
R3100 VNB.n946 VNB.n942 0.136
R3101 VNB.n950 VNB.n946 0.136
R3102 VNB.n954 VNB.n950 0.136
R3103 VNB.n960 VNB.n954 0.136
R3104 VNB.n971 VNB.n960 0.136
R3105 VNB.n975 VNB.n971 0.136
R3106 VNB.n979 VNB.n975 0.136
R3107 VNB.n1005 VNB.n1001 0.136
R3108 VNB.n1009 VNB.n1005 0.136
R3109 VNB.n1013 VNB.n1009 0.136
R3110 VNB.n1017 VNB.n1013 0.136
R3111 VNB.n1021 VNB.n1017 0.136
R3112 VNB.n1025 VNB.n1021 0.136
R3113 VNB.n1029 VNB.n1025 0.136
R3114 VNB.n1034 VNB.n1029 0.136
R3115 VNB.n1046 VNB.n1034 0.136
R3116 VNB.n1050 VNB.n1046 0.136
R3117 VNB.n1054 VNB.n1050 0.136
R3118 VNB.n1080 VNB.n1076 0.136
R3119 VNB.n1084 VNB.n1080 0.136
R3120 VNB.n1088 VNB.n1084 0.136
R3121 VNB.n1092 VNB.n1088 0.136
R3122 VNB.n1098 VNB.n1092 0.136
R3123 VNB.n1102 VNB.n1098 0.136
R3124 VNB.n1106 VNB.n1102 0.136
R3125 VNB.n1132 VNB.n1128 0.136
R3126 VNB.n1136 VNB.n1132 0.136
R3127 VNB.n1140 VNB.n1136 0.136
R3128 VNB.n1144 VNB.n1140 0.136
R3129 VNB.n1150 VNB.n1144 0.136
R3130 VNB.n1154 VNB.n1150 0.136
R3131 VNB.n1158 VNB.n1154 0.136
R3132 VNB.n1184 VNB.n1180 0.136
R3133 VNB.n1188 VNB.n1184 0.136
R3134 VNB.n1192 VNB.n1188 0.136
R3135 VNB.n1196 VNB.n1192 0.136
R3136 VNB.n1200 VNB.n1196 0.136
R3137 VNB.n1204 VNB.n1200 0.136
R3138 VNB.n1208 VNB.n1204 0.136
R3139 VNB.n1212 VNB.n1208 0.136
R3140 VNB.n1218 VNB.n1212 0.136
R3141 VNB.n1222 VNB.n1218 0.136
R3142 VNB.n1226 VNB.n1222 0.136
R3143 VNB.n1252 VNB.n1248 0.136
R3144 VNB.n1256 VNB.n1252 0.136
R3145 VNB.n1260 VNB.n1256 0.136
R3146 VNB.n1264 VNB.n1260 0.136
R3147 VNB.n1268 VNB.n1264 0.136
R3148 VNB.n1272 VNB.n1268 0.136
R3149 VNB.n1276 VNB.n1272 0.136
R3150 VNB.n1280 VNB.n1276 0.136
R3151 VNB.n1286 VNB.n1280 0.136
R3152 VNB.n1290 VNB.n1286 0.136
R3153 VNB.n1294 VNB.n1290 0.136
R3154 VNB.n1296 VNB.n1295 0.136
R3155 VNB.n1297 VNB.n1296 0.136
R3156 VNB.n1298 VNB.n1297 0.136
R3157 VNB.n1299 VNB.n1298 0.136
R3158 VNB.n1300 VNB.n1299 0.136
R3159 a_217_1004.n5 a_217_1004.t7 512.525
R3160 a_217_1004.n3 a_217_1004.t9 512.525
R3161 a_217_1004.n5 a_217_1004.t8 371.139
R3162 a_217_1004.n3 a_217_1004.t6 371.139
R3163 a_217_1004.n6 a_217_1004.n5 226.225
R3164 a_217_1004.n4 a_217_1004.n3 225.866
R3165 a_217_1004.n4 a_217_1004.t5 218.057
R3166 a_217_1004.n6 a_217_1004.t10 217.698
R3167 a_217_1004.n8 a_217_1004.n2 215.652
R3168 a_217_1004.n10 a_217_1004.n8 147.503
R3169 a_217_1004.n7 a_217_1004.n4 79.488
R3170 a_217_1004.n8 a_217_1004.n7 77.314
R3171 a_217_1004.n2 a_217_1004.n1 76.002
R3172 a_217_1004.n7 a_217_1004.n6 76
R3173 a_217_1004.n10 a_217_1004.n9 15.218
R3174 a_217_1004.n0 a_217_1004.t2 14.282
R3175 a_217_1004.n0 a_217_1004.t3 14.282
R3176 a_217_1004.n1 a_217_1004.t1 14.282
R3177 a_217_1004.n1 a_217_1004.t0 14.282
R3178 a_217_1004.n2 a_217_1004.n0 12.85
R3179 a_217_1004.n11 a_217_1004.n10 12.014
R3180 a_1719_75.n4 a_1719_75.n3 19.724
R3181 a_1719_75.t0 a_1719_75.n5 11.595
R3182 a_1719_75.t0 a_1719_75.n4 9.207
R3183 a_1719_75.n2 a_1719_75.n0 8.543
R3184 a_1719_75.t0 a_1719_75.n2 3.034
R3185 a_1719_75.n2 a_1719_75.n1 0.443
R3186 a_14869_1005.n4 a_14869_1005.n3 195.987
R3187 a_14869_1005.n2 a_14869_1005.t5 89.553
R3188 a_14869_1005.n4 a_14869_1005.n0 75.271
R3189 a_14869_1005.n3 a_14869_1005.n2 75.214
R3190 a_14869_1005.n5 a_14869_1005.n4 36.517
R3191 a_14869_1005.n3 a_14869_1005.t6 14.338
R3192 a_14869_1005.n1 a_14869_1005.t4 14.282
R3193 a_14869_1005.n1 a_14869_1005.t7 14.282
R3194 a_14869_1005.n0 a_14869_1005.t1 14.282
R3195 a_14869_1005.n0 a_14869_1005.t0 14.282
R3196 a_14869_1005.t3 a_14869_1005.n5 14.282
R3197 a_14869_1005.n5 a_14869_1005.t2 14.282
R3198 a_14869_1005.n2 a_14869_1005.n1 12.119
R3199 a_1265_943.n6 a_1265_943.t10 454.685
R3200 a_1265_943.n8 a_1265_943.t13 454.685
R3201 a_1265_943.n4 a_1265_943.t6 454.685
R3202 a_1265_943.n6 a_1265_943.t5 428.979
R3203 a_1265_943.n8 a_1265_943.t9 428.979
R3204 a_1265_943.n4 a_1265_943.t8 428.979
R3205 a_1265_943.n7 a_1265_943.t11 248.006
R3206 a_1265_943.n9 a_1265_943.t12 248.006
R3207 a_1265_943.n5 a_1265_943.t7 248.006
R3208 a_1265_943.n14 a_1265_943.n12 220.639
R3209 a_1265_943.n12 a_1265_943.n3 135.994
R3210 a_1265_943.n7 a_1265_943.n6 81.941
R3211 a_1265_943.n9 a_1265_943.n8 81.941
R3212 a_1265_943.n5 a_1265_943.n4 81.941
R3213 a_1265_943.n11 a_1265_943.n5 81.396
R3214 a_1265_943.n10 a_1265_943.n9 79.491
R3215 a_1265_943.n3 a_1265_943.n2 76.002
R3216 a_1265_943.n10 a_1265_943.n7 76
R3217 a_1265_943.n12 a_1265_943.n11 76
R3218 a_1265_943.n14 a_1265_943.n13 30
R3219 a_1265_943.n15 a_1265_943.n0 24.383
R3220 a_1265_943.n15 a_1265_943.n14 23.684
R3221 a_1265_943.n1 a_1265_943.t3 14.282
R3222 a_1265_943.n1 a_1265_943.t2 14.282
R3223 a_1265_943.n2 a_1265_943.t0 14.282
R3224 a_1265_943.n2 a_1265_943.t1 14.282
R3225 a_1265_943.n3 a_1265_943.n1 12.85
R3226 a_1265_943.n11 a_1265_943.n10 2.947
R3227 a_1905_1004.n6 a_1905_1004.t8 480.392
R3228 a_1905_1004.n6 a_1905_1004.t9 403.272
R3229 a_1905_1004.n8 a_1905_1004.n5 233.952
R3230 a_1905_1004.n7 a_1905_1004.t7 213.869
R3231 a_1905_1004.n7 a_1905_1004.n6 161.6
R3232 a_1905_1004.n8 a_1905_1004.n7 153.315
R3233 a_1905_1004.n10 a_1905_1004.n8 143.492
R3234 a_1905_1004.n4 a_1905_1004.n3 79.232
R3235 a_1905_1004.n5 a_1905_1004.n4 63.152
R3236 a_1905_1004.n10 a_1905_1004.n9 30
R3237 a_1905_1004.n11 a_1905_1004.n0 24.383
R3238 a_1905_1004.n11 a_1905_1004.n10 23.684
R3239 a_1905_1004.n5 a_1905_1004.n1 16.08
R3240 a_1905_1004.n4 a_1905_1004.n2 16.08
R3241 a_1905_1004.n1 a_1905_1004.t1 14.282
R3242 a_1905_1004.n1 a_1905_1004.t0 14.282
R3243 a_1905_1004.n2 a_1905_1004.t5 14.282
R3244 a_1905_1004.n2 a_1905_1004.t6 14.282
R3245 a_1905_1004.n3 a_1905_1004.t3 14.282
R3246 a_1905_1004.n3 a_1905_1004.t4 14.282
R3247 a_5101_1004.n6 a_5101_1004.t8 512.525
R3248 a_5101_1004.n4 a_5101_1004.t5 512.525
R3249 a_5101_1004.n6 a_5101_1004.t10 371.139
R3250 a_5101_1004.n4 a_5101_1004.t9 371.139
R3251 a_5101_1004.n7 a_5101_1004.n6 226.225
R3252 a_5101_1004.n5 a_5101_1004.n4 225.866
R3253 a_5101_1004.n5 a_5101_1004.t7 218.057
R3254 a_5101_1004.n7 a_5101_1004.t6 217.698
R3255 a_5101_1004.n9 a_5101_1004.n3 215.652
R3256 a_5101_1004.n11 a_5101_1004.n9 140.981
R3257 a_5101_1004.n8 a_5101_1004.n5 79.488
R3258 a_5101_1004.n9 a_5101_1004.n8 77.314
R3259 a_5101_1004.n3 a_5101_1004.n2 76.002
R3260 a_5101_1004.n8 a_5101_1004.n7 76
R3261 a_5101_1004.n11 a_5101_1004.n10 30
R3262 a_5101_1004.n12 a_5101_1004.n0 24.383
R3263 a_5101_1004.n12 a_5101_1004.n11 23.684
R3264 a_5101_1004.n1 a_5101_1004.t1 14.282
R3265 a_5101_1004.n1 a_5101_1004.t0 14.282
R3266 a_5101_1004.n2 a_5101_1004.t4 14.282
R3267 a_5101_1004.n2 a_5101_1004.t3 14.282
R3268 a_5101_1004.n3 a_5101_1004.n1 12.85
R3269 a_10111_383.n6 a_10111_383.t12 480.392
R3270 a_10111_383.n8 a_10111_383.t11 472.359
R3271 a_10111_383.n6 a_10111_383.t9 403.272
R3272 a_10111_383.n8 a_10111_383.t7 384.527
R3273 a_10111_383.n7 a_10111_383.t10 320.08
R3274 a_10111_383.n9 a_10111_383.t8 277.772
R3275 a_10111_383.n13 a_10111_383.n11 249.364
R3276 a_10111_383.n11 a_10111_383.n5 127.401
R3277 a_10111_383.n10 a_10111_383.n7 83.304
R3278 a_10111_383.n10 a_10111_383.n9 80.032
R3279 a_10111_383.n4 a_10111_383.n3 79.232
R3280 a_10111_383.n11 a_10111_383.n10 76
R3281 a_10111_383.n9 a_10111_383.n8 67.001
R3282 a_10111_383.n5 a_10111_383.n4 63.152
R3283 a_10111_383.n7 a_10111_383.n6 55.388
R3284 a_10111_383.n13 a_10111_383.n12 30
R3285 a_10111_383.n14 a_10111_383.n0 24.383
R3286 a_10111_383.n14 a_10111_383.n13 23.684
R3287 a_10111_383.n5 a_10111_383.n1 16.08
R3288 a_10111_383.n4 a_10111_383.n2 16.08
R3289 a_10111_383.n1 a_10111_383.t5 14.282
R3290 a_10111_383.n1 a_10111_383.t4 14.282
R3291 a_10111_383.n2 a_10111_383.t2 14.282
R3292 a_10111_383.n2 a_10111_383.t3 14.282
R3293 a_10111_383.n3 a_10111_383.t1 14.282
R3294 a_10111_383.n3 a_10111_383.t0 14.282
R3295 a_9985_1004.n5 a_9985_1004.t9 512.525
R3296 a_9985_1004.n3 a_9985_1004.t7 512.525
R3297 a_9985_1004.n5 a_9985_1004.t5 371.139
R3298 a_9985_1004.n3 a_9985_1004.t10 371.139
R3299 a_9985_1004.n6 a_9985_1004.n5 226.225
R3300 a_9985_1004.n4 a_9985_1004.n3 225.866
R3301 a_9985_1004.n4 a_9985_1004.t8 218.057
R3302 a_9985_1004.n6 a_9985_1004.t6 217.698
R3303 a_9985_1004.n8 a_9985_1004.n2 215.652
R3304 a_9985_1004.n10 a_9985_1004.n8 147.503
R3305 a_9985_1004.n7 a_9985_1004.n4 79.488
R3306 a_9985_1004.n8 a_9985_1004.n7 77.314
R3307 a_9985_1004.n2 a_9985_1004.n1 76.002
R3308 a_9985_1004.n7 a_9985_1004.n6 76
R3309 a_9985_1004.n10 a_9985_1004.n9 15.218
R3310 a_9985_1004.n0 a_9985_1004.t2 14.282
R3311 a_9985_1004.n0 a_9985_1004.t3 14.282
R3312 a_9985_1004.n1 a_9985_1004.t1 14.282
R3313 a_9985_1004.n1 a_9985_1004.t0 14.282
R3314 a_9985_1004.n2 a_9985_1004.n0 12.85
R3315 a_9985_1004.n11 a_9985_1004.n10 12.014
R3316 a_12470_73.t0 a_12470_73.n1 34.62
R3317 a_12470_73.t0 a_12470_73.n0 8.137
R3318 a_12470_73.t0 a_12470_73.n2 4.69
R3319 a_10806_182.n10 a_10806_182.n8 82.852
R3320 a_10806_182.n7 a_10806_182.n6 32.833
R3321 a_10806_182.n8 a_10806_182.t1 32.416
R3322 a_10806_182.n10 a_10806_182.n9 27.2
R3323 a_10806_182.n11 a_10806_182.n0 23.498
R3324 a_10806_182.n3 a_10806_182.n2 23.284
R3325 a_10806_182.n11 a_10806_182.n10 22.4
R3326 a_10806_182.n7 a_10806_182.n4 19.017
R3327 a_10806_182.n6 a_10806_182.n5 13.494
R3328 a_10806_182.t1 a_10806_182.n1 7.04
R3329 a_10806_182.t1 a_10806_182.n3 5.727
R3330 a_10806_182.n8 a_10806_182.n7 1.435
R3331 a_15430_73.n2 a_15430_73.n0 34.602
R3332 a_15430_73.n2 a_15430_73.n1 2.138
R3333 a_15430_73.t0 a_15430_73.n2 0.069
R3334 a_11673_1004.n6 a_11673_1004.t7 480.392
R3335 a_11673_1004.n6 a_11673_1004.t8 403.272
R3336 a_11673_1004.n8 a_11673_1004.n5 233.952
R3337 a_11673_1004.n7 a_11673_1004.t9 213.869
R3338 a_11673_1004.n7 a_11673_1004.n6 161.6
R3339 a_11673_1004.n8 a_11673_1004.n7 153.315
R3340 a_11673_1004.n10 a_11673_1004.n8 143.492
R3341 a_11673_1004.n4 a_11673_1004.n3 79.232
R3342 a_11673_1004.n5 a_11673_1004.n4 63.152
R3343 a_11673_1004.n10 a_11673_1004.n9 30
R3344 a_11673_1004.n11 a_11673_1004.n0 24.383
R3345 a_11673_1004.n11 a_11673_1004.n10 23.684
R3346 a_11673_1004.n5 a_11673_1004.n1 16.08
R3347 a_11673_1004.n4 a_11673_1004.n2 16.08
R3348 a_11673_1004.n1 a_11673_1004.t3 14.282
R3349 a_11673_1004.n1 a_11673_1004.t2 14.282
R3350 a_11673_1004.n2 a_11673_1004.t6 14.282
R3351 a_11673_1004.n2 a_11673_1004.t5 14.282
R3352 a_11673_1004.n3 a_11673_1004.t1 14.282
R3353 a_11673_1004.n3 a_11673_1004.t0 14.282
R3354 a_13781_75.n1 a_13781_75.n0 25.576
R3355 a_13781_75.n3 a_13781_75.n2 9.111
R3356 a_13781_75.n7 a_13781_75.n5 7.859
R3357 a_13781_75.t0 a_13781_75.n7 3.034
R3358 a_13781_75.n5 a_13781_75.n3 1.964
R3359 a_13781_75.n5 a_13781_75.n4 1.964
R3360 a_13781_75.t0 a_13781_75.n1 1.871
R3361 a_13781_75.n7 a_13781_75.n6 0.443
R3362 a_14062_182.n12 a_14062_182.n5 96.467
R3363 a_14062_182.t0 a_14062_182.n1 46.91
R3364 a_14062_182.n9 a_14062_182.n7 34.805
R3365 a_14062_182.n9 a_14062_182.n8 32.622
R3366 a_14062_182.t0 a_14062_182.n12 32.417
R3367 a_14062_182.n5 a_14062_182.n4 22.349
R3368 a_14062_182.n11 a_14062_182.n9 19.017
R3369 a_14062_182.n1 a_14062_182.n0 17.006
R3370 a_14062_182.n5 a_14062_182.n3 8.443
R3371 a_14062_182.t0 a_14062_182.n2 8.137
R3372 a_14062_182.n7 a_14062_182.n6 7.5
R3373 a_14062_182.n11 a_14062_182.n10 7.5
R3374 a_14062_182.n12 a_14062_182.n11 1.435
R3375 a_13241_1004.n9 a_13241_1004.t7 512.525
R3376 a_13241_1004.n6 a_13241_1004.t13 512.525
R3377 a_13241_1004.n4 a_13241_1004.t5 477.179
R3378 a_13241_1004.n4 a_13241_1004.t11 406.485
R3379 a_13241_1004.n9 a_13241_1004.t10 371.139
R3380 a_13241_1004.n6 a_13241_1004.t9 371.139
R3381 a_13241_1004.n10 a_13241_1004.t6 350.821
R3382 a_13241_1004.n5 a_13241_1004.t12 346.633
R3383 a_13241_1004.n7 a_13241_1004.t8 340.206
R3384 a_13241_1004.n14 a_13241_1004.n12 273.745
R3385 a_13241_1004.n10 a_13241_1004.n9 93.101
R3386 a_13241_1004.n7 a_13241_1004.n6 89.615
R3387 a_13241_1004.n12 a_13241_1004.n3 82.888
R3388 a_13241_1004.n8 a_13241_1004.n5 78.675
R3389 a_13241_1004.n12 a_13241_1004.n11 77.315
R3390 a_13241_1004.n3 a_13241_1004.n2 76.002
R3391 a_13241_1004.n8 a_13241_1004.n7 76
R3392 a_13241_1004.n11 a_13241_1004.n10 76
R3393 a_13241_1004.n14 a_13241_1004.n13 30
R3394 a_13241_1004.n5 a_13241_1004.n4 29.194
R3395 a_13241_1004.n15 a_13241_1004.n0 24.383
R3396 a_13241_1004.n15 a_13241_1004.n14 23.684
R3397 a_13241_1004.n1 a_13241_1004.t0 14.282
R3398 a_13241_1004.n1 a_13241_1004.t2 14.282
R3399 a_13241_1004.n2 a_13241_1004.t3 14.282
R3400 a_13241_1004.n2 a_13241_1004.t4 14.282
R3401 a_13241_1004.n3 a_13241_1004.n1 12.85
R3402 a_13241_1004.n11 a_13241_1004.n8 3.219
R3403 a_757_75.n1 a_757_75.n0 25.576
R3404 a_757_75.n3 a_757_75.n2 9.111
R3405 a_757_75.n7 a_757_75.n5 7.859
R3406 a_757_75.t0 a_757_75.n7 3.034
R3407 a_757_75.n5 a_757_75.n3 1.964
R3408 a_757_75.n5 a_757_75.n4 1.964
R3409 a_757_75.t0 a_757_75.n1 1.871
R3410 a_757_75.n7 a_757_75.n6 0.443
R3411 a_1038_182.n12 a_1038_182.n10 82.852
R3412 a_1038_182.n13 a_1038_182.n0 49.6
R3413 a_1038_182.t1 a_1038_182.n2 46.91
R3414 a_1038_182.n7 a_1038_182.n5 34.805
R3415 a_1038_182.n7 a_1038_182.n6 32.622
R3416 a_1038_182.n10 a_1038_182.t1 32.416
R3417 a_1038_182.n12 a_1038_182.n11 27.2
R3418 a_1038_182.n13 a_1038_182.n12 22.4
R3419 a_1038_182.n9 a_1038_182.n7 19.017
R3420 a_1038_182.n2 a_1038_182.n1 17.006
R3421 a_1038_182.n5 a_1038_182.n4 7.5
R3422 a_1038_182.n9 a_1038_182.n8 7.5
R3423 a_1038_182.t1 a_1038_182.n3 7.04
R3424 a_1038_182.n10 a_1038_182.n9 1.435
R3425 a_2702_73.t0 a_2702_73.n1 34.62
R3426 a_2702_73.t0 a_2702_73.n0 8.137
R3427 a_2702_73.t0 a_2702_73.n2 4.69
R3428 a_13136_73.t0 a_13136_73.n1 34.62
R3429 a_13136_73.t0 a_13136_73.n0 8.137
R3430 a_13136_73.t0 a_13136_73.n2 4.69
R3431 a_343_383.n6 a_343_383.t12 480.392
R3432 a_343_383.n8 a_343_383.t7 472.359
R3433 a_343_383.n6 a_343_383.t9 403.272
R3434 a_343_383.n8 a_343_383.t10 384.527
R3435 a_343_383.n7 a_343_383.t11 320.08
R3436 a_343_383.n9 a_343_383.t8 277.772
R3437 a_343_383.n13 a_343_383.n11 249.364
R3438 a_343_383.n11 a_343_383.n5 127.401
R3439 a_343_383.n10 a_343_383.n7 83.304
R3440 a_343_383.n10 a_343_383.n9 80.032
R3441 a_343_383.n4 a_343_383.n3 79.232
R3442 a_343_383.n11 a_343_383.n10 76
R3443 a_343_383.n9 a_343_383.n8 67.001
R3444 a_343_383.n5 a_343_383.n4 63.152
R3445 a_343_383.n7 a_343_383.n6 55.388
R3446 a_343_383.n14 a_343_383.n0 55.263
R3447 a_343_383.n13 a_343_383.n12 30
R3448 a_343_383.n14 a_343_383.n13 23.684
R3449 a_343_383.n5 a_343_383.n1 16.08
R3450 a_343_383.n4 a_343_383.n2 16.08
R3451 a_343_383.n1 a_343_383.t3 14.282
R3452 a_343_383.n1 a_343_383.t2 14.282
R3453 a_343_383.n2 a_343_383.t1 14.282
R3454 a_343_383.n2 a_343_383.t0 14.282
R3455 a_343_383.n3 a_343_383.t6 14.282
R3456 a_343_383.n3 a_343_383.t5 14.282
R3457 a_8252_73.n12 a_8252_73.n11 26.811
R3458 a_8252_73.n6 a_8252_73.n5 24.977
R3459 a_8252_73.n2 a_8252_73.n1 24.877
R3460 a_8252_73.t0 a_8252_73.n2 12.677
R3461 a_8252_73.t0 a_8252_73.n3 11.595
R3462 a_8252_73.t1 a_8252_73.n8 8.137
R3463 a_8252_73.t0 a_8252_73.n4 7.273
R3464 a_8252_73.t0 a_8252_73.n0 6.109
R3465 a_8252_73.t1 a_8252_73.n7 4.864
R3466 a_8252_73.t0 a_8252_73.n12 2.074
R3467 a_8252_73.n7 a_8252_73.n6 1.13
R3468 a_8252_73.n12 a_8252_73.t1 0.937
R3469 a_8252_73.t1 a_8252_73.n10 0.804
R3470 a_8252_73.n10 a_8252_73.n9 0.136
R3471 a_112_73.n12 a_112_73.n11 26.811
R3472 a_112_73.n6 a_112_73.n5 24.977
R3473 a_112_73.n2 a_112_73.n1 24.877
R3474 a_112_73.t0 a_112_73.n2 12.677
R3475 a_112_73.t0 a_112_73.n3 11.595
R3476 a_112_73.t1 a_112_73.n8 8.137
R3477 a_112_73.t0 a_112_73.n4 7.273
R3478 a_112_73.t0 a_112_73.n0 6.109
R3479 a_112_73.t1 a_112_73.n7 4.864
R3480 a_112_73.t0 a_112_73.n12 2.074
R3481 a_112_73.n7 a_112_73.n6 1.13
R3482 a_112_73.n12 a_112_73.t1 0.937
R3483 a_112_73.t1 a_112_73.n10 0.804
R3484 a_112_73.n10 a_112_73.n9 0.136
R3485 a_13367_383.n6 a_13367_383.t9 472.359
R3486 a_13367_383.n6 a_13367_383.t7 384.527
R3487 a_13367_383.n7 a_13367_383.t8 277.772
R3488 a_13367_383.n10 a_13367_383.n8 249.704
R3489 a_13367_383.n8 a_13367_383.n7 156.035
R3490 a_13367_383.n8 a_13367_383.n5 127.74
R3491 a_13367_383.n4 a_13367_383.n3 79.232
R3492 a_13367_383.n7 a_13367_383.n6 67.001
R3493 a_13367_383.n5 a_13367_383.n4 63.152
R3494 a_13367_383.n11 a_13367_383.n0 55.263
R3495 a_13367_383.n10 a_13367_383.n9 30
R3496 a_13367_383.n11 a_13367_383.n10 23.684
R3497 a_13367_383.n5 a_13367_383.n1 16.08
R3498 a_13367_383.n4 a_13367_383.n2 16.08
R3499 a_13367_383.n1 a_13367_383.t4 14.282
R3500 a_13367_383.n1 a_13367_383.t3 14.282
R3501 a_13367_383.n2 a_13367_383.t6 14.282
R3502 a_13367_383.n2 a_13367_383.t5 14.282
R3503 a_13367_383.n3 a_13367_383.t1 14.282
R3504 a_13367_383.n3 a_13367_383.t0 14.282
R3505 a_5641_75.n1 a_5641_75.n0 25.576
R3506 a_5641_75.n3 a_5641_75.n2 9.111
R3507 a_5641_75.n7 a_5641_75.n5 7.859
R3508 a_5641_75.t0 a_5641_75.n7 3.034
R3509 a_5641_75.n5 a_5641_75.n3 1.964
R3510 a_5641_75.n5 a_5641_75.n4 1.964
R3511 a_5641_75.t0 a_5641_75.n1 1.871
R3512 a_5641_75.n7 a_5641_75.n6 0.443
R3513 a_4294_182.n9 a_4294_182.n7 82.852
R3514 a_4294_182.n3 a_4294_182.n1 44.628
R3515 a_4294_182.t0 a_4294_182.n9 32.417
R3516 a_4294_182.n7 a_4294_182.n6 27.2
R3517 a_4294_182.n5 a_4294_182.n4 23.498
R3518 a_4294_182.n3 a_4294_182.n2 23.284
R3519 a_4294_182.n7 a_4294_182.n5 22.4
R3520 a_4294_182.t0 a_4294_182.n11 20.241
R3521 a_4294_182.n11 a_4294_182.n10 13.494
R3522 a_4294_182.t0 a_4294_182.n0 8.137
R3523 a_4294_182.t0 a_4294_182.n3 5.727
R3524 a_4294_182.n9 a_4294_182.n8 1.435
R3525 a_11768_182.n9 a_11768_182.n7 82.852
R3526 a_11768_182.n3 a_11768_182.n1 44.628
R3527 a_11768_182.t0 a_11768_182.n9 32.417
R3528 a_11768_182.n7 a_11768_182.n6 27.2
R3529 a_11768_182.n5 a_11768_182.n4 23.498
R3530 a_11768_182.n3 a_11768_182.n2 23.284
R3531 a_11768_182.n7 a_11768_182.n5 22.4
R3532 a_11768_182.t0 a_11768_182.n11 20.241
R3533 a_11768_182.n11 a_11768_182.n10 13.494
R3534 a_11768_182.t0 a_11768_182.n0 8.137
R3535 a_11768_182.t0 a_11768_182.n3 5.727
R3536 a_11768_182.n9 a_11768_182.n8 1.435
R3537 a_2000_182.n8 a_2000_182.n6 96.467
R3538 a_2000_182.n3 a_2000_182.n1 44.628
R3539 a_2000_182.t0 a_2000_182.n8 32.417
R3540 a_2000_182.n3 a_2000_182.n2 23.284
R3541 a_2000_182.n6 a_2000_182.n5 22.349
R3542 a_2000_182.t0 a_2000_182.n10 20.241
R3543 a_2000_182.n10 a_2000_182.n9 13.494
R3544 a_2000_182.n6 a_2000_182.n4 8.443
R3545 a_2000_182.t0 a_2000_182.n0 8.137
R3546 a_2000_182.t0 a_2000_182.n3 5.727
R3547 a_2000_182.n8 a_2000_182.n7 1.435
R3548 a_3368_73.n12 a_3368_73.n11 26.811
R3549 a_3368_73.n6 a_3368_73.n5 24.977
R3550 a_3368_73.n2 a_3368_73.n1 24.877
R3551 a_3368_73.t0 a_3368_73.n2 12.677
R3552 a_3368_73.t0 a_3368_73.n3 11.595
R3553 a_3368_73.t1 a_3368_73.n8 8.137
R3554 a_3368_73.t0 a_3368_73.n4 7.273
R3555 a_3368_73.t0 a_3368_73.n0 6.109
R3556 a_3368_73.t1 a_3368_73.n7 4.864
R3557 a_3368_73.t0 a_3368_73.n12 2.074
R3558 a_3368_73.n7 a_3368_73.n6 1.13
R3559 a_3368_73.n12 a_3368_73.t1 0.937
R3560 a_3368_73.t1 a_3368_73.n10 0.804
R3561 a_3368_73.n10 a_3368_73.n9 0.136
R3562 a_14764_73.n1 a_14764_73.n0 32.249
R3563 a_14764_73.t0 a_14764_73.n5 7.911
R3564 a_14764_73.n4 a_14764_73.n2 4.032
R3565 a_14764_73.n4 a_14764_73.n3 3.644
R3566 a_14764_73.t0 a_14764_73.n1 2.534
R3567 a_14764_73.t0 a_14764_73.n4 1.099
R3568 a_6603_75.n5 a_6603_75.n4 19.724
R3569 a_6603_75.t0 a_6603_75.n3 11.595
R3570 a_6603_75.t0 a_6603_75.n5 9.207
R3571 a_6603_75.n2 a_6603_75.n1 2.455
R3572 a_6603_75.n2 a_6603_75.n0 1.32
R3573 a_6603_75.t0 a_6603_75.n2 0.246
R3574 a_4013_75.n5 a_4013_75.n4 19.724
R3575 a_4013_75.t0 a_4013_75.n3 11.595
R3576 a_4013_75.t0 a_4013_75.n5 9.207
R3577 a_4013_75.n2 a_4013_75.n1 2.455
R3578 a_4013_75.n2 a_4013_75.n0 1.32
R3579 a_4013_75.t0 a_4013_75.n2 0.246
R3580 a_5922_182.n10 a_5922_182.n8 82.852
R3581 a_5922_182.n11 a_5922_182.n0 49.6
R3582 a_5922_182.n7 a_5922_182.n6 32.833
R3583 a_5922_182.n8 a_5922_182.t1 32.416
R3584 a_5922_182.n10 a_5922_182.n9 27.2
R3585 a_5922_182.n3 a_5922_182.n2 23.284
R3586 a_5922_182.n11 a_5922_182.n10 22.4
R3587 a_5922_182.n7 a_5922_182.n4 19.017
R3588 a_5922_182.n6 a_5922_182.n5 13.494
R3589 a_5922_182.t1 a_5922_182.n1 7.04
R3590 a_5922_182.t1 a_5922_182.n3 5.727
R3591 a_5922_182.n8 a_5922_182.n7 1.435
R3592 a_7586_73.n12 a_7586_73.n11 26.811
R3593 a_7586_73.n6 a_7586_73.n5 24.977
R3594 a_7586_73.n2 a_7586_73.n1 24.877
R3595 a_7586_73.t0 a_7586_73.n2 12.677
R3596 a_7586_73.t0 a_7586_73.n3 11.595
R3597 a_7586_73.t1 a_7586_73.n8 8.137
R3598 a_7586_73.t0 a_7586_73.n4 7.273
R3599 a_7586_73.t0 a_7586_73.n0 6.109
R3600 a_7586_73.t1 a_7586_73.n7 4.864
R3601 a_7586_73.t0 a_7586_73.n12 2.074
R3602 a_7586_73.n7 a_7586_73.n6 1.13
R3603 a_7586_73.n12 a_7586_73.t1 0.937
R3604 a_7586_73.t1 a_7586_73.n10 0.804
R3605 a_7586_73.n10 a_7586_73.n9 0.136
R3606 a_10525_75.n1 a_10525_75.n0 25.576
R3607 a_10525_75.n3 a_10525_75.n2 9.111
R3608 a_10525_75.n7 a_10525_75.n6 2.455
R3609 a_10525_75.n5 a_10525_75.n3 1.964
R3610 a_10525_75.n5 a_10525_75.n4 1.964
R3611 a_10525_75.t0 a_10525_75.n1 1.871
R3612 a_10525_75.n7 a_10525_75.n5 0.636
R3613 a_10525_75.t0 a_10525_75.n7 0.246
R3614 a_16096_73.t0 a_16096_73.n1 34.62
R3615 a_16096_73.t0 a_16096_73.n0 8.137
R3616 a_16096_73.t0 a_16096_73.n2 4.69
R3617 a_4996_73.t0 a_4996_73.n1 34.62
R3618 a_4996_73.t0 a_4996_73.n0 8.137
R3619 a_4996_73.t0 a_4996_73.n2 4.69
R3620 a_9178_182.n10 a_9178_182.n8 82.852
R3621 a_9178_182.n7 a_9178_182.n6 32.833
R3622 a_9178_182.n8 a_9178_182.t1 32.416
R3623 a_9178_182.n10 a_9178_182.n9 27.2
R3624 a_9178_182.n11 a_9178_182.n0 23.498
R3625 a_9178_182.n3 a_9178_182.n2 23.284
R3626 a_9178_182.n11 a_9178_182.n10 22.4
R3627 a_9178_182.n7 a_9178_182.n4 19.017
R3628 a_9178_182.n6 a_9178_182.n5 13.494
R3629 a_9178_182.t1 a_9178_182.n1 7.04
R3630 a_9178_182.t1 a_9178_182.n3 5.727
R3631 a_9178_182.n8 a_9178_182.n7 1.435
R3632 a_11487_75.n5 a_11487_75.n4 19.724
R3633 a_11487_75.t0 a_11487_75.n3 11.595
R3634 a_11487_75.t0 a_11487_75.n5 9.207
R3635 a_11487_75.n2 a_11487_75.n1 2.455
R3636 a_11487_75.n2 a_11487_75.n0 1.32
R3637 a_11487_75.t0 a_11487_75.n2 0.246
R3638 a_8897_75.n5 a_8897_75.n4 19.724
R3639 a_8897_75.t0 a_8897_75.n3 11.595
R3640 a_8897_75.t0 a_8897_75.n5 9.207
R3641 a_8897_75.n2 a_8897_75.n1 2.455
R3642 a_8897_75.n2 a_8897_75.n0 1.32
R3643 a_8897_75.t0 a_8897_75.n2 0.246
C6 VPB VNB 62.14fF
C7 a_8897_75.n0 VNB 0.10fF
C8 a_8897_75.n1 VNB 0.04fF
C9 a_8897_75.n2 VNB 0.03fF
C10 a_8897_75.n3 VNB 0.07fF
C11 a_8897_75.n4 VNB 0.08fF
C12 a_8897_75.n5 VNB 0.06fF
C13 a_11487_75.n0 VNB 0.10fF
C14 a_11487_75.n1 VNB 0.04fF
C15 a_11487_75.n2 VNB 0.03fF
C16 a_11487_75.n3 VNB 0.07fF
C17 a_11487_75.n4 VNB 0.08fF
C18 a_11487_75.n5 VNB 0.06fF
C19 a_9178_182.n0 VNB 0.02fF
C20 a_9178_182.n1 VNB 0.09fF
C21 a_9178_182.n2 VNB 0.13fF
C22 a_9178_182.n3 VNB 0.11fF
C23 a_9178_182.t1 VNB 0.30fF
C24 a_9178_182.n4 VNB 0.09fF
C25 a_9178_182.n5 VNB 0.06fF
C26 a_9178_182.n6 VNB 0.01fF
C27 a_9178_182.n7 VNB 0.03fF
C28 a_9178_182.n8 VNB 0.11fF
C29 a_9178_182.n9 VNB 0.02fF
C30 a_9178_182.n10 VNB 0.05fF
C31 a_9178_182.n11 VNB 0.03fF
C32 a_4996_73.n0 VNB 0.05fF
C33 a_4996_73.n1 VNB 0.12fF
C34 a_4996_73.n2 VNB 0.04fF
C35 a_16096_73.n0 VNB 0.06fF
C36 a_16096_73.n1 VNB 0.13fF
C37 a_16096_73.n2 VNB 0.04fF
C38 a_10525_75.n0 VNB 0.09fF
C39 a_10525_75.n1 VNB 0.10fF
C40 a_10525_75.n2 VNB 0.05fF
C41 a_10525_75.n3 VNB 0.03fF
C42 a_10525_75.n4 VNB 0.04fF
C43 a_10525_75.n5 VNB 0.03fF
C44 a_10525_75.n6 VNB 0.04fF
C45 a_7586_73.n0 VNB 0.02fF
C46 a_7586_73.n1 VNB 0.10fF
C47 a_7586_73.n2 VNB 0.06fF
C48 a_7586_73.n3 VNB 0.06fF
C49 a_7586_73.n4 VNB 0.00fF
C50 a_7586_73.n5 VNB 0.04fF
C51 a_7586_73.n6 VNB 0.05fF
C52 a_7586_73.n7 VNB 0.02fF
C53 a_7586_73.n8 VNB 0.05fF
C54 a_7586_73.n9 VNB 0.08fF
C55 a_7586_73.n10 VNB 0.17fF
C56 a_7586_73.t1 VNB 0.23fF
C57 a_7586_73.n11 VNB 0.09fF
C58 a_7586_73.n12 VNB 0.00fF
C59 a_5922_182.n0 VNB 0.02fF
C60 a_5922_182.n1 VNB 0.09fF
C61 a_5922_182.n2 VNB 0.13fF
C62 a_5922_182.n3 VNB 0.11fF
C63 a_5922_182.t1 VNB 0.30fF
C64 a_5922_182.n4 VNB 0.09fF
C65 a_5922_182.n5 VNB 0.06fF
C66 a_5922_182.n6 VNB 0.01fF
C67 a_5922_182.n7 VNB 0.03fF
C68 a_5922_182.n8 VNB 0.11fF
C69 a_5922_182.n9 VNB 0.02fF
C70 a_5922_182.n10 VNB 0.05fF
C71 a_5922_182.n11 VNB 0.02fF
C72 a_4013_75.n0 VNB 0.10fF
C73 a_4013_75.n1 VNB 0.04fF
C74 a_4013_75.n2 VNB 0.03fF
C75 a_4013_75.n3 VNB 0.07fF
C76 a_4013_75.n4 VNB 0.08fF
C77 a_4013_75.n5 VNB 0.06fF
C78 a_6603_75.n0 VNB 0.10fF
C79 a_6603_75.n1 VNB 0.04fF
C80 a_6603_75.n2 VNB 0.03fF
C81 a_6603_75.n3 VNB 0.07fF
C82 a_6603_75.n4 VNB 0.08fF
C83 a_6603_75.n5 VNB 0.06fF
C84 a_14764_73.n0 VNB 0.11fF
C85 a_14764_73.n1 VNB 0.09fF
C86 a_14764_73.n2 VNB 0.08fF
C87 a_14764_73.n3 VNB 0.02fF
C88 a_14764_73.n4 VNB 0.01fF
C89 a_14764_73.n5 VNB 0.06fF
C90 a_3368_73.n0 VNB 0.02fF
C91 a_3368_73.n1 VNB 0.10fF
C92 a_3368_73.n2 VNB 0.06fF
C93 a_3368_73.n3 VNB 0.06fF
C94 a_3368_73.n4 VNB 0.00fF
C95 a_3368_73.n5 VNB 0.04fF
C96 a_3368_73.n6 VNB 0.05fF
C97 a_3368_73.n7 VNB 0.02fF
C98 a_3368_73.n8 VNB 0.05fF
C99 a_3368_73.n9 VNB 0.08fF
C100 a_3368_73.n10 VNB 0.17fF
C101 a_3368_73.t1 VNB 0.23fF
C102 a_3368_73.n11 VNB 0.09fF
C103 a_3368_73.n12 VNB 0.00fF
C104 a_2000_182.n0 VNB 0.07fF
C105 a_2000_182.n1 VNB 0.09fF
C106 a_2000_182.n2 VNB 0.13fF
C107 a_2000_182.n3 VNB 0.11fF
C108 a_2000_182.n4 VNB 0.02fF
C109 a_2000_182.n5 VNB 0.03fF
C110 a_2000_182.n6 VNB 0.06fF
C111 a_2000_182.n7 VNB 0.03fF
C112 a_2000_182.n8 VNB 0.12fF
C113 a_2000_182.n9 VNB 0.06fF
C114 a_2000_182.n10 VNB 0.01fF
C115 a_2000_182.t0 VNB 0.33fF
C116 a_11768_182.n0 VNB 0.07fF
C117 a_11768_182.n1 VNB 0.09fF
C118 a_11768_182.n2 VNB 0.13fF
C119 a_11768_182.n3 VNB 0.11fF
C120 a_11768_182.n4 VNB 0.02fF
C121 a_11768_182.n5 VNB 0.03fF
C122 a_11768_182.n6 VNB 0.02fF
C123 a_11768_182.n7 VNB 0.05fF
C124 a_11768_182.n8 VNB 0.03fF
C125 a_11768_182.n9 VNB 0.11fF
C126 a_11768_182.n10 VNB 0.06fF
C127 a_11768_182.n11 VNB 0.01fF
C128 a_11768_182.t0 VNB 0.33fF
C129 a_4294_182.n0 VNB 0.07fF
C130 a_4294_182.n1 VNB 0.09fF
C131 a_4294_182.n2 VNB 0.13fF
C132 a_4294_182.n3 VNB 0.11fF
C133 a_4294_182.n4 VNB 0.02fF
C134 a_4294_182.n5 VNB 0.03fF
C135 a_4294_182.n6 VNB 0.02fF
C136 a_4294_182.n7 VNB 0.05fF
C137 a_4294_182.n8 VNB 0.03fF
C138 a_4294_182.n9 VNB 0.11fF
C139 a_4294_182.n10 VNB 0.06fF
C140 a_4294_182.n11 VNB 0.01fF
C141 a_4294_182.t0 VNB 0.33fF
C142 a_5641_75.n0 VNB 0.09fF
C143 a_5641_75.n1 VNB 0.10fF
C144 a_5641_75.n2 VNB 0.05fF
C145 a_5641_75.n3 VNB 0.03fF
C146 a_5641_75.n4 VNB 0.04fF
C147 a_5641_75.n5 VNB 0.11fF
C148 a_5641_75.n6 VNB 0.04fF
C149 a_13367_383.n0 VNB 0.05fF
C150 a_13367_383.n1 VNB 0.69fF
C151 a_13367_383.n2 VNB 0.69fF
C152 a_13367_383.n3 VNB 0.81fF
C153 a_13367_383.n4 VNB 0.25fF
C154 a_13367_383.n5 VNB 0.33fF
C155 a_13367_383.n6 VNB 0.37fF
C156 a_13367_383.t8 VNB 0.73fF
C157 a_13367_383.n7 VNB 1.09fF
C158 a_13367_383.n8 VNB 1.18fF
C159 a_13367_383.n9 VNB 0.05fF
C160 a_13367_383.n10 VNB 0.44fF
C161 a_13367_383.n11 VNB 0.06fF
C162 a_112_73.n0 VNB 0.02fF
C163 a_112_73.n1 VNB 0.10fF
C164 a_112_73.n2 VNB 0.06fF
C165 a_112_73.n3 VNB 0.06fF
C166 a_112_73.n4 VNB 0.00fF
C167 a_112_73.n5 VNB 0.04fF
C168 a_112_73.n6 VNB 0.05fF
C169 a_112_73.n7 VNB 0.02fF
C170 a_112_73.n8 VNB 0.05fF
C171 a_112_73.n9 VNB 0.07fF
C172 a_112_73.n10 VNB 0.17fF
C173 a_112_73.t1 VNB 0.22fF
C174 a_112_73.n11 VNB 0.09fF
C175 a_112_73.n12 VNB 0.00fF
C176 a_8252_73.n0 VNB 0.02fF
C177 a_8252_73.n1 VNB 0.10fF
C178 a_8252_73.n2 VNB 0.06fF
C179 a_8252_73.n3 VNB 0.06fF
C180 a_8252_73.n4 VNB 0.00fF
C181 a_8252_73.n5 VNB 0.04fF
C182 a_8252_73.n6 VNB 0.05fF
C183 a_8252_73.n7 VNB 0.02fF
C184 a_8252_73.n8 VNB 0.05fF
C185 a_8252_73.n9 VNB 0.08fF
C186 a_8252_73.n10 VNB 0.17fF
C187 a_8252_73.t1 VNB 0.23fF
C188 a_8252_73.n11 VNB 0.09fF
C189 a_8252_73.n12 VNB 0.00fF
C190 a_343_383.n0 VNB 0.06fF
C191 a_343_383.n1 VNB 0.76fF
C192 a_343_383.n2 VNB 0.76fF
C193 a_343_383.n3 VNB 0.89fF
C194 a_343_383.n4 VNB 0.28fF
C195 a_343_383.n5 VNB 0.36fF
C196 a_343_383.n6 VNB 0.46fF
C197 a_343_383.n7 VNB 0.66fF
C198 a_343_383.n8 VNB 0.41fF
C199 a_343_383.t8 VNB 0.81fF
C200 a_343_383.n9 VNB 0.56fF
C201 a_343_383.n10 VNB 3.54fF
C202 a_343_383.n11 VNB 0.63fF
C203 a_343_383.n12 VNB 0.06fF
C204 a_343_383.n13 VNB 0.49fF
C205 a_343_383.n14 VNB 0.06fF
C206 a_13136_73.n0 VNB 0.05fF
C207 a_13136_73.n1 VNB 0.12fF
C208 a_13136_73.n2 VNB 0.04fF
C209 a_2702_73.n0 VNB 0.05fF
C210 a_2702_73.n1 VNB 0.12fF
C211 a_2702_73.n2 VNB 0.04fF
C212 a_1038_182.n0 VNB 0.02fF
C213 a_1038_182.n1 VNB 0.07fF
C214 a_1038_182.n2 VNB 0.13fF
C215 a_1038_182.n3 VNB 0.09fF
C216 a_1038_182.t1 VNB 0.25fF
C217 a_1038_182.n4 VNB 0.05fF
C218 a_1038_182.n5 VNB 0.06fF
C219 a_1038_182.n6 VNB 0.07fF
C220 a_1038_182.n7 VNB 0.07fF
C221 a_1038_182.n8 VNB 0.03fF
C222 a_1038_182.n9 VNB 0.01fF
C223 a_1038_182.n10 VNB 0.11fF
C224 a_1038_182.n11 VNB 0.02fF
C225 a_1038_182.n12 VNB 0.05fF
C226 a_1038_182.n13 VNB 0.02fF
C227 a_757_75.n0 VNB 0.09fF
C228 a_757_75.n1 VNB 0.10fF
C229 a_757_75.n2 VNB 0.05fF
C230 a_757_75.n3 VNB 0.03fF
C231 a_757_75.n4 VNB 0.04fF
C232 a_757_75.n5 VNB 0.11fF
C233 a_757_75.n6 VNB 0.04fF
C234 a_13241_1004.n0 VNB 0.04fF
C235 a_13241_1004.n1 VNB 0.56fF
C236 a_13241_1004.n2 VNB 0.66fF
C237 a_13241_1004.n3 VNB 0.24fF
C238 a_13241_1004.n4 VNB 0.31fF
C239 a_13241_1004.n5 VNB 0.43fF
C240 a_13241_1004.n6 VNB 0.28fF
C241 a_13241_1004.n7 VNB 0.50fF
C242 a_13241_1004.n8 VNB 1.05fF
C243 a_13241_1004.n9 VNB 0.27fF
C244 a_13241_1004.n10 VNB 0.51fF
C245 a_13241_1004.n11 VNB 0.74fF
C246 a_13241_1004.n12 VNB 0.44fF
C247 a_13241_1004.n13 VNB 0.04fF
C248 a_13241_1004.n14 VNB 0.39fF
C249 a_13241_1004.n15 VNB 0.06fF
C250 a_14062_182.n0 VNB 0.07fF
C251 a_14062_182.n1 VNB 0.13fF
C252 a_14062_182.n2 VNB 0.07fF
C253 a_14062_182.n3 VNB 0.02fF
C254 a_14062_182.n4 VNB 0.03fF
C255 a_14062_182.n5 VNB 0.06fF
C256 a_14062_182.n6 VNB 0.05fF
C257 a_14062_182.n7 VNB 0.06fF
C258 a_14062_182.n8 VNB 0.07fF
C259 a_14062_182.n9 VNB 0.07fF
C260 a_14062_182.n10 VNB 0.03fF
C261 a_14062_182.n11 VNB 0.01fF
C262 a_14062_182.n12 VNB 0.12fF
C263 a_14062_182.t0 VNB 0.28fF
C264 a_13781_75.n0 VNB 0.09fF
C265 a_13781_75.n1 VNB 0.10fF
C266 a_13781_75.n2 VNB 0.05fF
C267 a_13781_75.n3 VNB 0.03fF
C268 a_13781_75.n4 VNB 0.04fF
C269 a_13781_75.n5 VNB 0.11fF
C270 a_13781_75.n6 VNB 0.04fF
C271 a_11673_1004.n0 VNB 0.04fF
C272 a_11673_1004.n1 VNB 0.56fF
C273 a_11673_1004.n2 VNB 0.56fF
C274 a_11673_1004.n3 VNB 0.65fF
C275 a_11673_1004.n4 VNB 0.21fF
C276 a_11673_1004.n5 VNB 0.39fF
C277 a_11673_1004.n6 VNB 0.46fF
C278 a_11673_1004.n7 VNB 0.57fF
C279 a_11673_1004.n8 VNB 0.65fF
C280 a_11673_1004.n9 VNB 0.04fF
C281 a_11673_1004.n10 VNB 0.23fF
C282 a_11673_1004.n11 VNB 0.06fF
C283 a_15430_73.n0 VNB 0.13fF
C284 a_15430_73.n1 VNB 0.13fF
C285 a_15430_73.n2 VNB 0.14fF
C286 a_10806_182.n0 VNB 0.02fF
C287 a_10806_182.n1 VNB 0.09fF
C288 a_10806_182.n2 VNB 0.13fF
C289 a_10806_182.n3 VNB 0.11fF
C290 a_10806_182.t1 VNB 0.30fF
C291 a_10806_182.n4 VNB 0.09fF
C292 a_10806_182.n5 VNB 0.06fF
C293 a_10806_182.n6 VNB 0.01fF
C294 a_10806_182.n7 VNB 0.03fF
C295 a_10806_182.n8 VNB 0.11fF
C296 a_10806_182.n9 VNB 0.02fF
C297 a_10806_182.n10 VNB 0.05fF
C298 a_10806_182.n11 VNB 0.03fF
C299 a_12470_73.n0 VNB 0.05fF
C300 a_12470_73.n1 VNB 0.12fF
C301 a_12470_73.n2 VNB 0.04fF
C302 a_9985_1004.n0 VNB 0.72fF
C303 a_9985_1004.n1 VNB 0.85fF
C304 a_9985_1004.n2 VNB 0.51fF
C305 a_9985_1004.n3 VNB 0.55fF
C306 a_9985_1004.n4 VNB 0.64fF
C307 a_9985_1004.n5 VNB 0.56fF
C308 a_9985_1004.n6 VNB 0.61fF
C309 a_9985_1004.n7 VNB 1.53fF
C310 a_9985_1004.n8 VNB 0.59fF
C311 a_9985_1004.n9 VNB 0.11fF
C312 a_9985_1004.n10 VNB 0.28fF
C313 a_9985_1004.n11 VNB 0.06fF
C314 a_10111_383.n0 VNB 0.06fF
C315 a_10111_383.n1 VNB 0.86fF
C316 a_10111_383.n2 VNB 0.86fF
C317 a_10111_383.n3 VNB 1.01fF
C318 a_10111_383.n4 VNB 0.32fF
C319 a_10111_383.n5 VNB 0.41fF
C320 a_10111_383.n6 VNB 0.52fF
C321 a_10111_383.n7 VNB 0.75fF
C322 a_10111_383.n8 VNB 0.46fF
C323 a_10111_383.t8 VNB 0.92fF
C324 a_10111_383.n9 VNB 0.64fF
C325 a_10111_383.n10 VNB 4.03fF
C326 a_10111_383.n11 VNB 0.72fF
C327 a_10111_383.n12 VNB 0.06fF
C328 a_10111_383.n13 VNB 0.55fF
C329 a_10111_383.n14 VNB 0.09fF
C330 a_5101_1004.n0 VNB 0.05fF
C331 a_5101_1004.n1 VNB 0.71fF
C332 a_5101_1004.n2 VNB 0.85fF
C333 a_5101_1004.n3 VNB 0.51fF
C334 a_5101_1004.n4 VNB 0.55fF
C335 a_5101_1004.n5 VNB 0.64fF
C336 a_5101_1004.n6 VNB 0.55fF
C337 a_5101_1004.n7 VNB 0.61fF
C338 a_5101_1004.n8 VNB 1.53fF
C339 a_5101_1004.n9 VNB 0.57fF
C340 a_5101_1004.n10 VNB 0.05fF
C341 a_5101_1004.n11 VNB 0.29fF
C342 a_5101_1004.n12 VNB 0.07fF
C343 a_1905_1004.n0 VNB 0.04fF
C344 a_1905_1004.n1 VNB 0.53fF
C345 a_1905_1004.n2 VNB 0.53fF
C346 a_1905_1004.n3 VNB 0.63fF
C347 a_1905_1004.n4 VNB 0.20fF
C348 a_1905_1004.n5 VNB 0.38fF
C349 a_1905_1004.n6 VNB 0.45fF
C350 a_1905_1004.n7 VNB 0.55fF
C351 a_1905_1004.n8 VNB 0.62fF
C352 a_1905_1004.n9 VNB 0.03fF
C353 a_1905_1004.n10 VNB 0.22fF
C354 a_1905_1004.n11 VNB 0.05fF
C355 a_1265_943.n0 VNB 0.06fF
C356 a_1265_943.n1 VNB 0.80fF
C357 a_1265_943.n2 VNB 0.95fF
C358 a_1265_943.n3 VNB 0.43fF
C359 a_1265_943.n4 VNB 0.54fF
C360 a_1265_943.t7 VNB 0.82fF
C361 a_1265_943.n5 VNB 0.61fF
C362 a_1265_943.n6 VNB 0.54fF
C363 a_1265_943.t11 VNB 0.82fF
C364 a_1265_943.n7 VNB 0.54fF
C365 a_1265_943.n8 VNB 0.54fF
C366 a_1265_943.t12 VNB 0.82fF
C367 a_1265_943.n9 VNB 0.57fF
C368 a_1265_943.n10 VNB 1.72fF
C369 a_1265_943.n11 VNB 2.32fF
C370 a_1265_943.n12 VNB 0.63fF
C371 a_1265_943.n13 VNB 0.05fF
C372 a_1265_943.n14 VNB 0.47fF
C373 a_1265_943.n15 VNB 0.08fF
C374 a_14869_1005.n0 VNB 0.41fF
C375 a_14869_1005.n1 VNB 0.33fF
C376 a_14869_1005.n2 VNB 0.23fF
C377 a_14869_1005.n3 VNB 0.63fF
C378 a_14869_1005.n4 VNB 0.28fF
C379 a_14869_1005.n5 VNB 0.37fF
C380 a_1719_75.n0 VNB 0.20fF
C381 a_1719_75.n1 VNB 0.04fF
C382 a_1719_75.n2 VNB 0.01fF
C383 a_1719_75.n3 VNB 0.08fF
C384 a_1719_75.n4 VNB 0.06fF
C385 a_1719_75.n5 VNB 0.07fF
C386 a_217_1004.n0 VNB 0.54fF
C387 a_217_1004.n1 VNB 0.64fF
C388 a_217_1004.n2 VNB 0.38fF
C389 a_217_1004.n3 VNB 0.42fF
C390 a_217_1004.n4 VNB 0.48fF
C391 a_217_1004.n5 VNB 0.42fF
C392 a_217_1004.n6 VNB 0.46fF
C393 a_217_1004.n7 VNB 1.15fF
C394 a_217_1004.n8 VNB 0.44fF
C395 a_217_1004.n9 VNB 0.08fF
C396 a_217_1004.n10 VNB 0.21fF
C397 a_217_1004.n11 VNB 0.05fF
C398 a_9880_73.n0 VNB 0.05fF
C399 a_9880_73.n1 VNB 0.02fF
C400 a_9880_73.n2 VNB 0.12fF
C401 a_9880_73.n3 VNB 0.04fF
C402 a_9880_73.n4 VNB 0.17fF
C403 a_8483_383.n0 VNB 0.05fF
C404 a_8483_383.n1 VNB 0.73fF
C405 a_8483_383.n2 VNB 0.73fF
C406 a_8483_383.n3 VNB 0.85fF
C407 a_8483_383.n4 VNB 0.27fF
C408 a_8483_383.n5 VNB 0.35fF
C409 a_8483_383.n6 VNB 0.39fF
C410 a_8483_383.t7 VNB 0.77fF
C411 a_8483_383.n7 VNB 1.15fF
C412 a_8483_383.n8 VNB 1.25fF
C413 a_8483_383.n9 VNB 0.05fF
C414 a_8483_383.n10 VNB 0.47fF
C415 a_8483_383.n11 VNB 0.07fF
C416 a_8357_1004.n0 VNB 1.04fF
C417 a_8357_1004.n1 VNB 1.23fF
C418 a_8357_1004.n2 VNB 0.74fF
C419 a_8357_1004.n3 VNB 0.56fF
C420 a_8357_1004.n4 VNB 0.63fF
C421 a_8357_1004.t12 VNB 1.12fF
C422 a_8357_1004.n5 VNB 1.88fF
C423 a_8357_1004.n6 VNB 1.44fF
C424 a_8357_1004.t8 VNB 0.96fF
C425 a_8357_1004.n7 VNB 1.67fF
C426 a_8357_1004.n8 VNB 0.80fF
C427 a_8357_1004.n9 VNB 0.89fF
C428 a_8357_1004.n10 VNB 9.30fF
C429 a_8357_1004.n11 VNB 0.85fF
C430 a_8357_1004.n12 VNB 0.16fF
C431 a_8357_1004.n13 VNB 0.40fF
C432 a_8357_1004.n14 VNB 0.09fF
C433 a_11033_943.n0 VNB 0.07fF
C434 a_11033_943.n1 VNB 0.93fF
C435 a_11033_943.n2 VNB 1.10fF
C436 a_11033_943.n3 VNB 0.50fF
C437 a_11033_943.n4 VNB 0.62fF
C438 a_11033_943.t12 VNB 0.95fF
C439 a_11033_943.n5 VNB 0.71fF
C440 a_11033_943.n6 VNB 0.62fF
C441 a_11033_943.t8 VNB 0.95fF
C442 a_11033_943.n7 VNB 0.63fF
C443 a_11033_943.n8 VNB 0.62fF
C444 a_11033_943.t5 VNB 0.95fF
C445 a_11033_943.n9 VNB 0.67fF
C446 a_11033_943.n10 VNB 2.00fF
C447 a_11033_943.n11 VNB 2.70fF
C448 a_11033_943.n12 VNB 0.73fF
C449 a_11033_943.n13 VNB 0.06fF
C450 a_11033_943.n14 VNB 0.54fF
C451 a_11033_943.n15 VNB 0.09fF
C452 a_3599_383.n0 VNB 0.05fF
C453 a_3599_383.n1 VNB 0.71fF
C454 a_3599_383.n2 VNB 0.71fF
C455 a_3599_383.n3 VNB 0.83fF
C456 a_3599_383.n4 VNB 0.26fF
C457 a_3599_383.n5 VNB 0.34fF
C458 a_3599_383.n6 VNB 0.38fF
C459 a_3599_383.t8 VNB 0.75fF
C460 a_3599_383.n7 VNB 1.11fF
C461 a_3599_383.n8 VNB 1.20fF
C462 a_3599_383.n9 VNB 0.06fF
C463 a_3599_383.n10 VNB 0.45fF
C464 a_3599_383.n11 VNB 0.06fF
C465 a_15533_1005.n0 VNB 0.28fF
C466 a_15533_1005.n1 VNB 0.35fF
C467 a_15533_1005.n2 VNB 0.25fF
C468 a_15533_1005.n3 VNB 0.56fF
C469 a_15533_1005.n4 VNB 0.20fF
C470 a_15533_1005.n5 VNB 0.29fF
C471 a_15044_181.n0 VNB 0.42fF
C472 a_15044_181.n1 VNB 0.51fF
C473 a_15044_181.n2 VNB 0.48fF
C474 a_15044_181.n3 VNB 0.04fF
C475 a_15044_181.n4 VNB 0.05fF
C476 a_15044_181.n5 VNB 0.03fF
C477 a_15044_181.n6 VNB 0.09fF
C478 a_15044_181.n7 VNB 0.04fF
C479 a_15044_181.n8 VNB 0.05fF
C480 a_15044_181.n9 VNB 0.11fF
C481 a_15044_181.n10 VNB 1.09fF
C482 a_15044_181.n11 VNB 0.43fF
C483 a_15044_181.n12 VNB 0.08fF
C484 a_15044_181.n13 VNB 0.04fF
C485 a_15044_181.n14 VNB 0.04fF
C486 a_3473_1004.n0 VNB 1.31fF
C487 a_3473_1004.n1 VNB 1.55fF
C488 a_3473_1004.n2 VNB 0.79fF
C489 a_3473_1004.n3 VNB 0.89fF
C490 a_3473_1004.n4 VNB 1.15fF
C491 a_3473_1004.n5 VNB 1.42fF
C492 a_3473_1004.t7 VNB 1.09fF
C493 a_3473_1004.n6 VNB 0.93fF
C494 a_3473_1004.n7 VNB 5.04fF
C495 a_3473_1004.n8 VNB 0.86fF
C496 a_3473_1004.n9 VNB 1.15fF
C497 a_3473_1004.n10 VNB 20.24fF
C498 a_3473_1004.n11 VNB 1.07fF
C499 a_3473_1004.n12 VNB 0.21fF
C500 a_3473_1004.n13 VNB 0.67fF
C501 a_3473_1004.n14 VNB 0.11fF
C502 VPB.n0 VNB 0.03fF
C503 VPB.n1 VNB 0.04fF
C504 VPB.n2 VNB 0.02fF
C505 VPB.n3 VNB 0.14fF
C506 VPB.n5 VNB 0.02fF
C507 VPB.n6 VNB 0.02fF
C508 VPB.n7 VNB 0.02fF
C509 VPB.n8 VNB 0.02fF
C510 VPB.n10 VNB 0.02fF
C511 VPB.n11 VNB 0.02fF
C512 VPB.n12 VNB 0.02fF
C513 VPB.n14 VNB 0.10fF
C514 VPB.n15 VNB 0.02fF
C515 VPB.n16 VNB 0.02fF
C516 VPB.n17 VNB 0.02fF
C517 VPB.n18 VNB 0.04fF
C518 VPB.n19 VNB 0.02fF
C519 VPB.n20 VNB 0.25fF
C520 VPB.n21 VNB 0.04fF
C521 VPB.n23 VNB 0.02fF
C522 VPB.n24 VNB 0.02fF
C523 VPB.n25 VNB 0.02fF
C524 VPB.n26 VNB 0.02fF
C525 VPB.n28 VNB 0.02fF
C526 VPB.n29 VNB 0.02fF
C527 VPB.n30 VNB 0.02fF
C528 VPB.n32 VNB 0.28fF
C529 VPB.n34 VNB 0.03fF
C530 VPB.n35 VNB 0.02fF
C531 VPB.n36 VNB 0.03fF
C532 VPB.n37 VNB 0.03fF
C533 VPB.n38 VNB 0.28fF
C534 VPB.n39 VNB 0.01fF
C535 VPB.n40 VNB 0.02fF
C536 VPB.n41 VNB 0.24fF
C537 VPB.n42 VNB 0.02fF
C538 VPB.n43 VNB 0.01fF
C539 VPB.n44 VNB 0.05fF
C540 VPB.n45 VNB 0.14fF
C541 VPB.n46 VNB 0.16fF
C542 VPB.n47 VNB 0.02fF
C543 VPB.n48 VNB 0.02fF
C544 VPB.n49 VNB 0.14fF
C545 VPB.n50 VNB 0.15fF
C546 VPB.n51 VNB 0.02fF
C547 VPB.n52 VNB 0.02fF
C548 VPB.n53 VNB 0.02fF
C549 VPB.n54 VNB 0.14fF
C550 VPB.n55 VNB 0.15fF
C551 VPB.n56 VNB 0.02fF
C552 VPB.n57 VNB 0.02fF
C553 VPB.n58 VNB 0.14fF
C554 VPB.n59 VNB 0.16fF
C555 VPB.n60 VNB 0.02fF
C556 VPB.n61 VNB 0.02fF
C557 VPB.n62 VNB 0.06fF
C558 VPB.n63 VNB 0.24fF
C559 VPB.n64 VNB 0.02fF
C560 VPB.n65 VNB 0.01fF
C561 VPB.n66 VNB 0.02fF
C562 VPB.n67 VNB 0.02fF
C563 VPB.n68 VNB 0.02fF
C564 VPB.n69 VNB 0.14fF
C565 VPB.n70 VNB 0.03fF
C566 VPB.n71 VNB 0.02fF
C567 VPB.n72 VNB 0.05fF
C568 VPB.n73 VNB 0.01fF
C569 VPB.n75 VNB 0.02fF
C570 VPB.n76 VNB 0.02fF
C571 VPB.n77 VNB 0.02fF
C572 VPB.n78 VNB 0.02fF
C573 VPB.n81 VNB 0.02fF
C574 VPB.n83 VNB 0.46fF
C575 VPB.n85 VNB 0.04fF
C576 VPB.n86 VNB 0.04fF
C577 VPB.n87 VNB 0.28fF
C578 VPB.n88 VNB 0.03fF
C579 VPB.n89 VNB 0.04fF
C580 VPB.n90 VNB 0.28fF
C581 VPB.n91 VNB 0.02fF
C582 VPB.n92 VNB 0.02fF
C583 VPB.n93 VNB 0.28fF
C584 VPB.n94 VNB 0.02fF
C585 VPB.n95 VNB 0.02fF
C586 VPB.n96 VNB 0.28fF
C587 VPB.n97 VNB 0.02fF
C588 VPB.n98 VNB 0.02fF
C589 VPB.n99 VNB 0.00fF
C590 VPB.n100 VNB 0.10fF
C591 VPB.n101 VNB 0.02fF
C592 VPB.n102 VNB 0.28fF
C593 VPB.n103 VNB 0.02fF
C594 VPB.n104 VNB 0.02fF
C595 VPB.n105 VNB 0.02fF
C596 VPB.n106 VNB 0.28fF
C597 VPB.n107 VNB 0.02fF
C598 VPB.n108 VNB 0.02fF
C599 VPB.n109 VNB 0.02fF
C600 VPB.n110 VNB 0.28fF
C601 VPB.n111 VNB 0.02fF
C602 VPB.n112 VNB 0.02fF
C603 VPB.n113 VNB 0.02fF
C604 VPB.n114 VNB 0.28fF
C605 VPB.n115 VNB 0.01fF
C606 VPB.n116 VNB 0.02fF
C607 VPB.n117 VNB 0.04fF
C608 VPB.n118 VNB 0.02fF
C609 VPB.n119 VNB 0.02fF
C610 VPB.n120 VNB 0.02fF
C611 VPB.n121 VNB 0.04fF
C612 VPB.n122 VNB 0.02fF
C613 VPB.n123 VNB 0.20fF
C614 VPB.n124 VNB 0.04fF
C615 VPB.n126 VNB 0.02fF
C616 VPB.n127 VNB 0.02fF
C617 VPB.n128 VNB 0.02fF
C618 VPB.n129 VNB 0.02fF
C619 VPB.n131 VNB 0.02fF
C620 VPB.n132 VNB 0.02fF
C621 VPB.n133 VNB 0.02fF
C622 VPB.n135 VNB 0.28fF
C623 VPB.n137 VNB 0.03fF
C624 VPB.n138 VNB 0.02fF
C625 VPB.n139 VNB 0.03fF
C626 VPB.n140 VNB 0.03fF
C627 VPB.n141 VNB 0.28fF
C628 VPB.n142 VNB 0.01fF
C629 VPB.n143 VNB 0.02fF
C630 VPB.n144 VNB 0.04fF
C631 VPB.n145 VNB 0.28fF
C632 VPB.n146 VNB 0.02fF
C633 VPB.n147 VNB 0.02fF
C634 VPB.n148 VNB 0.02fF
C635 VPB.n149 VNB 0.28fF
C636 VPB.n150 VNB 0.02fF
C637 VPB.n151 VNB 0.02fF
C638 VPB.n152 VNB 0.02fF
C639 VPB.n153 VNB 0.28fF
C640 VPB.n154 VNB 0.02fF
C641 VPB.n155 VNB 0.02fF
C642 VPB.n156 VNB 0.02fF
C643 VPB.n157 VNB 0.28fF
C644 VPB.n158 VNB 0.02fF
C645 VPB.n159 VNB 0.02fF
C646 VPB.n160 VNB 0.02fF
C647 VPB.n161 VNB 0.28fF
C648 VPB.n162 VNB 0.02fF
C649 VPB.n163 VNB 0.02fF
C650 VPB.n164 VNB 0.02fF
C651 VPB.n165 VNB 0.28fF
C652 VPB.n166 VNB 0.02fF
C653 VPB.n167 VNB 0.02fF
C654 VPB.n168 VNB 0.02fF
C655 VPB.n169 VNB 0.28fF
C656 VPB.n170 VNB 0.01fF
C657 VPB.n171 VNB 0.02fF
C658 VPB.n172 VNB 0.04fF
C659 VPB.n173 VNB 0.02fF
C660 VPB.n174 VNB 0.02fF
C661 VPB.n175 VNB 0.02fF
C662 VPB.n176 VNB 0.04fF
C663 VPB.n177 VNB 0.02fF
C664 VPB.n178 VNB 0.20fF
C665 VPB.n179 VNB 0.04fF
C666 VPB.n181 VNB 0.02fF
C667 VPB.n182 VNB 0.02fF
C668 VPB.n183 VNB 0.02fF
C669 VPB.n184 VNB 0.02fF
C670 VPB.n186 VNB 0.02fF
C671 VPB.n187 VNB 0.02fF
C672 VPB.n188 VNB 0.02fF
C673 VPB.n190 VNB 0.28fF
C674 VPB.n192 VNB 0.03fF
C675 VPB.n193 VNB 0.02fF
C676 VPB.n194 VNB 0.03fF
C677 VPB.n195 VNB 0.03fF
C678 VPB.n196 VNB 0.28fF
C679 VPB.n197 VNB 0.01fF
C680 VPB.n198 VNB 0.02fF
C681 VPB.n199 VNB 0.04fF
C682 VPB.n200 VNB 0.06fF
C683 VPB.n201 VNB 0.24fF
C684 VPB.n202 VNB 0.02fF
C685 VPB.n203 VNB 0.01fF
C686 VPB.n204 VNB 0.02fF
C687 VPB.n205 VNB 0.14fF
C688 VPB.n206 VNB 0.16fF
C689 VPB.n207 VNB 0.02fF
C690 VPB.n208 VNB 0.02fF
C691 VPB.n209 VNB 0.02fF
C692 VPB.n210 VNB 0.10fF
C693 VPB.n211 VNB 0.02fF
C694 VPB.n212 VNB 0.14fF
C695 VPB.n213 VNB 0.15fF
C696 VPB.n214 VNB 0.02fF
C697 VPB.n215 VNB 0.02fF
C698 VPB.n216 VNB 0.02fF
C699 VPB.n217 VNB 0.14fF
C700 VPB.n218 VNB 0.15fF
C701 VPB.n219 VNB 0.02fF
C702 VPB.n220 VNB 0.02fF
C703 VPB.n221 VNB 0.02fF
C704 VPB.n222 VNB 0.14fF
C705 VPB.n223 VNB 0.16fF
C706 VPB.n224 VNB 0.02fF
C707 VPB.n225 VNB 0.02fF
C708 VPB.n226 VNB 0.02fF
C709 VPB.n227 VNB 0.06fF
C710 VPB.n228 VNB 0.24fF
C711 VPB.n229 VNB 0.02fF
C712 VPB.n230 VNB 0.01fF
C713 VPB.n231 VNB 0.02fF
C714 VPB.n232 VNB 0.28fF
C715 VPB.n233 VNB 0.01fF
C716 VPB.n234 VNB 0.02fF
C717 VPB.n235 VNB 0.04fF
C718 VPB.n236 VNB 0.02fF
C719 VPB.n237 VNB 0.02fF
C720 VPB.n238 VNB 0.02fF
C721 VPB.n239 VNB 0.04fF
C722 VPB.n240 VNB 0.02fF
C723 VPB.n241 VNB 0.24fF
C724 VPB.n242 VNB 0.04fF
C725 VPB.n244 VNB 0.02fF
C726 VPB.n245 VNB 0.02fF
C727 VPB.n246 VNB 0.02fF
C728 VPB.n247 VNB 0.02fF
C729 VPB.n249 VNB 0.02fF
C730 VPB.n250 VNB 0.02fF
C731 VPB.n251 VNB 0.02fF
C732 VPB.n253 VNB 0.28fF
C733 VPB.n255 VNB 0.03fF
C734 VPB.n256 VNB 0.02fF
C735 VPB.n257 VNB 0.03fF
C736 VPB.n258 VNB 0.03fF
C737 VPB.n259 VNB 0.28fF
C738 VPB.n260 VNB 0.01fF
C739 VPB.n261 VNB 0.02fF
C740 VPB.n262 VNB 0.04fF
C741 VPB.n263 VNB 0.28fF
C742 VPB.n264 VNB 0.02fF
C743 VPB.n265 VNB 0.02fF
C744 VPB.n266 VNB 0.02fF
C745 VPB.n267 VNB 0.05fF
C746 VPB.n268 VNB 0.21fF
C747 VPB.n269 VNB 0.02fF
C748 VPB.n270 VNB 0.01fF
C749 VPB.n271 VNB 0.02fF
C750 VPB.n272 VNB 0.14fF
C751 VPB.n273 VNB 0.16fF
C752 VPB.n274 VNB 0.02fF
C753 VPB.n275 VNB 0.02fF
C754 VPB.n276 VNB 0.02fF
C755 VPB.n277 VNB 0.10fF
C756 VPB.n278 VNB 0.02fF
C757 VPB.n279 VNB 0.14fF
C758 VPB.n280 VNB 0.16fF
C759 VPB.n281 VNB 0.02fF
C760 VPB.n282 VNB 0.02fF
C761 VPB.n283 VNB 0.02fF
C762 VPB.n284 VNB 0.14fF
C763 VPB.n285 VNB 0.15fF
C764 VPB.n286 VNB 0.02fF
C765 VPB.n287 VNB 0.02fF
C766 VPB.n288 VNB 0.02fF
C767 VPB.n289 VNB 0.14fF
C768 VPB.n290 VNB 0.15fF
C769 VPB.n291 VNB 0.02fF
C770 VPB.n292 VNB 0.02fF
C771 VPB.n293 VNB 0.02fF
C772 VPB.n294 VNB 0.10fF
C773 VPB.n295 VNB 0.02fF
C774 VPB.n296 VNB 0.14fF
C775 VPB.n297 VNB 0.16fF
C776 VPB.n298 VNB 0.02fF
C777 VPB.n299 VNB 0.02fF
C778 VPB.n300 VNB 0.02fF
C779 VPB.n301 VNB 0.14fF
C780 VPB.n302 VNB 0.16fF
C781 VPB.n303 VNB 0.02fF
C782 VPB.n304 VNB 0.02fF
C783 VPB.n305 VNB 0.02fF
C784 VPB.n306 VNB 0.06fF
C785 VPB.n307 VNB 0.21fF
C786 VPB.n308 VNB 0.02fF
C787 VPB.n309 VNB 0.01fF
C788 VPB.n310 VNB 0.02fF
C789 VPB.n311 VNB 0.28fF
C790 VPB.n312 VNB 0.02fF
C791 VPB.n313 VNB 0.02fF
C792 VPB.n314 VNB 0.02fF
C793 VPB.n315 VNB 0.28fF
C794 VPB.n316 VNB 0.01fF
C795 VPB.n317 VNB 0.02fF
C796 VPB.n318 VNB 0.04fF
C797 VPB.n319 VNB 0.02fF
C798 VPB.n320 VNB 0.02fF
C799 VPB.n321 VNB 0.02fF
C800 VPB.n322 VNB 0.04fF
C801 VPB.n323 VNB 0.02fF
C802 VPB.n324 VNB 0.24fF
C803 VPB.n325 VNB 0.04fF
C804 VPB.n327 VNB 0.02fF
C805 VPB.n328 VNB 0.02fF
C806 VPB.n329 VNB 0.02fF
C807 VPB.n330 VNB 0.02fF
C808 VPB.n332 VNB 0.02fF
C809 VPB.n333 VNB 0.02fF
C810 VPB.n334 VNB 0.02fF
C811 VPB.n336 VNB 0.28fF
C812 VPB.n338 VNB 0.03fF
C813 VPB.n339 VNB 0.02fF
C814 VPB.n340 VNB 0.03fF
C815 VPB.n341 VNB 0.03fF
C816 VPB.n342 VNB 0.28fF
C817 VPB.n343 VNB 0.01fF
C818 VPB.n344 VNB 0.02fF
C819 VPB.n345 VNB 0.04fF
C820 VPB.n346 VNB 0.05fF
C821 VPB.n347 VNB 0.24fF
C822 VPB.n348 VNB 0.02fF
C823 VPB.n349 VNB 0.01fF
C824 VPB.n350 VNB 0.02fF
C825 VPB.n351 VNB 0.14fF
C826 VPB.n352 VNB 0.16fF
C827 VPB.n353 VNB 0.02fF
C828 VPB.n354 VNB 0.02fF
C829 VPB.n355 VNB 0.02fF
C830 VPB.n356 VNB 0.10fF
C831 VPB.n357 VNB 0.02fF
C832 VPB.n358 VNB 0.14fF
C833 VPB.n359 VNB 0.15fF
C834 VPB.n360 VNB 0.02fF
C835 VPB.n361 VNB 0.02fF
C836 VPB.n362 VNB 0.02fF
C837 VPB.n363 VNB 0.14fF
C838 VPB.n364 VNB 0.15fF
C839 VPB.n365 VNB 0.02fF
C840 VPB.n366 VNB 0.02fF
C841 VPB.n367 VNB 0.02fF
C842 VPB.n368 VNB 0.14fF
C843 VPB.n369 VNB 0.16fF
C844 VPB.n370 VNB 0.02fF
C845 VPB.n371 VNB 0.02fF
C846 VPB.n372 VNB 0.02fF
C847 VPB.n373 VNB 0.06fF
C848 VPB.n374 VNB 0.24fF
C849 VPB.n375 VNB 0.02fF
C850 VPB.n376 VNB 0.01fF
C851 VPB.n377 VNB 0.02fF
C852 VPB.n378 VNB 0.28fF
C853 VPB.n379 VNB 0.01fF
C854 VPB.n380 VNB 0.02fF
C855 VPB.n381 VNB 0.04fF
C856 VPB.n382 VNB 0.02fF
C857 VPB.n383 VNB 0.02fF
C858 VPB.n384 VNB 0.02fF
C859 VPB.n385 VNB 0.04fF
C860 VPB.n386 VNB 0.02fF
C861 VPB.n387 VNB 0.20fF
C862 VPB.n388 VNB 0.04fF
C863 VPB.n390 VNB 0.02fF
C864 VPB.n391 VNB 0.02fF
C865 VPB.n392 VNB 0.02fF
C866 VPB.n393 VNB 0.02fF
C867 VPB.n395 VNB 0.02fF
C868 VPB.n396 VNB 0.02fF
C869 VPB.n397 VNB 0.02fF
C870 VPB.n399 VNB 0.28fF
C871 VPB.n401 VNB 0.03fF
C872 VPB.n402 VNB 0.02fF
C873 VPB.n403 VNB 0.03fF
C874 VPB.n404 VNB 0.03fF
C875 VPB.n405 VNB 0.28fF
C876 VPB.n406 VNB 0.01fF
C877 VPB.n407 VNB 0.02fF
C878 VPB.n408 VNB 0.04fF
C879 VPB.n409 VNB 0.05fF
C880 VPB.n410 VNB 0.24fF
C881 VPB.n411 VNB 0.02fF
C882 VPB.n412 VNB 0.01fF
C883 VPB.n413 VNB 0.02fF
C884 VPB.n414 VNB 0.14fF
C885 VPB.n415 VNB 0.16fF
C886 VPB.n416 VNB 0.02fF
C887 VPB.n417 VNB 0.02fF
C888 VPB.n418 VNB 0.02fF
C889 VPB.n419 VNB 0.10fF
C890 VPB.n420 VNB 0.02fF
C891 VPB.n421 VNB 0.14fF
C892 VPB.n422 VNB 0.15fF
C893 VPB.n423 VNB 0.02fF
C894 VPB.n424 VNB 0.02fF
C895 VPB.n425 VNB 0.02fF
C896 VPB.n426 VNB 0.14fF
C897 VPB.n427 VNB 0.15fF
C898 VPB.n428 VNB 0.02fF
C899 VPB.n429 VNB 0.02fF
C900 VPB.n430 VNB 0.02fF
C901 VPB.n431 VNB 0.14fF
C902 VPB.n432 VNB 0.16fF
C903 VPB.n433 VNB 0.02fF
C904 VPB.n434 VNB 0.02fF
C905 VPB.n435 VNB 0.02fF
C906 VPB.n436 VNB 0.06fF
C907 VPB.n437 VNB 0.24fF
C908 VPB.n438 VNB 0.02fF
C909 VPB.n439 VNB 0.01fF
C910 VPB.n440 VNB 0.02fF
C911 VPB.n441 VNB 0.28fF
C912 VPB.n442 VNB 0.01fF
C913 VPB.n443 VNB 0.02fF
C914 VPB.n444 VNB 0.04fF
C915 VPB.n445 VNB 0.02fF
C916 VPB.n446 VNB 0.02fF
C917 VPB.n447 VNB 0.02fF
C918 VPB.n448 VNB 0.04fF
C919 VPB.n449 VNB 0.02fF
C920 VPB.n450 VNB 0.24fF
C921 VPB.n451 VNB 0.04fF
C922 VPB.n453 VNB 0.02fF
C923 VPB.n454 VNB 0.02fF
C924 VPB.n455 VNB 0.02fF
C925 VPB.n456 VNB 0.02fF
C926 VPB.n458 VNB 0.02fF
C927 VPB.n459 VNB 0.02fF
C928 VPB.n460 VNB 0.02fF
C929 VPB.n462 VNB 0.28fF
C930 VPB.n464 VNB 0.03fF
C931 VPB.n465 VNB 0.02fF
C932 VPB.n466 VNB 0.03fF
C933 VPB.n467 VNB 0.03fF
C934 VPB.n468 VNB 0.28fF
C935 VPB.n469 VNB 0.01fF
C936 VPB.n470 VNB 0.02fF
C937 VPB.n471 VNB 0.04fF
C938 VPB.n472 VNB 0.28fF
C939 VPB.n473 VNB 0.02fF
C940 VPB.n474 VNB 0.02fF
C941 VPB.n475 VNB 0.02fF
C942 VPB.n476 VNB 0.05fF
C943 VPB.n477 VNB 0.21fF
C944 VPB.n478 VNB 0.02fF
C945 VPB.n479 VNB 0.01fF
C946 VPB.n480 VNB 0.02fF
C947 VPB.n481 VNB 0.14fF
C948 VPB.n482 VNB 0.16fF
C949 VPB.n483 VNB 0.02fF
C950 VPB.n484 VNB 0.02fF
C951 VPB.n485 VNB 0.02fF
C952 VPB.n486 VNB 0.10fF
C953 VPB.n487 VNB 0.02fF
C954 VPB.n488 VNB 0.14fF
C955 VPB.n489 VNB 0.16fF
C956 VPB.n490 VNB 0.02fF
C957 VPB.n491 VNB 0.02fF
C958 VPB.n492 VNB 0.02fF
C959 VPB.n493 VNB 0.14fF
C960 VPB.n494 VNB 0.15fF
C961 VPB.n495 VNB 0.02fF
C962 VPB.n496 VNB 0.02fF
C963 VPB.n497 VNB 0.02fF
C964 VPB.n498 VNB 0.14fF
C965 VPB.n499 VNB 0.15fF
C966 VPB.n500 VNB 0.02fF
C967 VPB.n501 VNB 0.02fF
C968 VPB.n502 VNB 0.02fF
C969 VPB.n503 VNB 0.10fF
C970 VPB.n504 VNB 0.02fF
C971 VPB.n505 VNB 0.14fF
C972 VPB.n506 VNB 0.16fF
C973 VPB.n507 VNB 0.02fF
C974 VPB.n508 VNB 0.02fF
C975 VPB.n509 VNB 0.02fF
C976 VPB.n510 VNB 0.14fF
C977 VPB.n511 VNB 0.16fF
C978 VPB.n512 VNB 0.02fF
C979 VPB.n513 VNB 0.02fF
C980 VPB.n514 VNB 0.02fF
C981 VPB.n515 VNB 0.06fF
C982 VPB.n516 VNB 0.21fF
C983 VPB.n517 VNB 0.02fF
C984 VPB.n518 VNB 0.01fF
C985 VPB.n519 VNB 0.02fF
C986 VPB.n520 VNB 0.28fF
C987 VPB.n521 VNB 0.02fF
C988 VPB.n522 VNB 0.02fF
C989 VPB.n523 VNB 0.02fF
C990 VPB.n524 VNB 0.28fF
C991 VPB.n525 VNB 0.01fF
C992 VPB.n526 VNB 0.02fF
C993 VPB.n527 VNB 0.04fF
C994 VPB.n528 VNB 0.02fF
C995 VPB.n529 VNB 0.02fF
C996 VPB.n530 VNB 0.02fF
C997 VPB.n531 VNB 0.04fF
C998 VPB.n532 VNB 0.02fF
C999 VPB.n533 VNB 0.29fF
C1000 VPB.n534 VNB 0.04fF
C1001 VPB.n536 VNB 0.02fF
C1002 VPB.n537 VNB 0.02fF
C1003 VPB.n538 VNB 0.02fF
C1004 VPB.n539 VNB 0.02fF
C1005 VPB.n541 VNB 0.02fF
C1006 VPB.n542 VNB 0.02fF
C1007 VPB.n543 VNB 0.02fF
C1008 VPB.n545 VNB 0.28fF
C1009 VPB.n547 VNB 0.03fF
C1010 VPB.n548 VNB 0.02fF
C1011 VPB.n549 VNB 0.03fF
C1012 VPB.n550 VNB 0.03fF
C1013 VPB.n551 VNB 0.28fF
C1014 VPB.n552 VNB 0.01fF
C1015 VPB.n553 VNB 0.02fF
C1016 VPB.n554 VNB 0.04fF
C1017 VPB.n555 VNB 0.28fF
C1018 VPB.n556 VNB 0.02fF
C1019 VPB.n557 VNB 0.02fF
C1020 VPB.n558 VNB 0.02fF
C1021 VPB.n559 VNB 0.05fF
C1022 VPB.n560 VNB 0.21fF
C1023 VPB.n561 VNB 0.02fF
C1024 VPB.n562 VNB 0.01fF
C1025 VPB.n563 VNB 0.02fF
C1026 VPB.n564 VNB 0.14fF
C1027 VPB.n565 VNB 0.16fF
C1028 VPB.n566 VNB 0.02fF
C1029 VPB.n567 VNB 0.02fF
C1030 VPB.n568 VNB 0.02fF
C1031 VPB.n569 VNB 0.10fF
C1032 VPB.n570 VNB 0.02fF
C1033 VPB.n571 VNB 0.14fF
C1034 VPB.n572 VNB 0.16fF
C1035 VPB.n573 VNB 0.02fF
C1036 VPB.n574 VNB 0.02fF
C1037 VPB.n575 VNB 0.02fF
C1038 VPB.n576 VNB 0.14fF
C1039 VPB.n577 VNB 0.15fF
C1040 VPB.n578 VNB 0.02fF
C1041 VPB.n579 VNB 0.02fF
C1042 VPB.n580 VNB 0.02fF
C1043 VPB.n581 VNB 0.14fF
C1044 VPB.n582 VNB 0.15fF
C1045 VPB.n583 VNB 0.02fF
C1046 VPB.n584 VNB 0.02fF
C1047 VPB.n585 VNB 0.02fF
C1048 VPB.n586 VNB 0.10fF
C1049 VPB.n587 VNB 0.02fF
C1050 VPB.n588 VNB 0.14fF
C1051 VPB.n589 VNB 0.16fF
C1052 VPB.n590 VNB 0.02fF
C1053 VPB.n591 VNB 0.02fF
C1054 VPB.n592 VNB 0.02fF
C1055 VPB.n593 VNB 0.14fF
C1056 VPB.n594 VNB 0.16fF
C1057 VPB.n595 VNB 0.02fF
C1058 VPB.n596 VNB 0.02fF
C1059 VPB.n597 VNB 0.02fF
C1060 VPB.n598 VNB 0.06fF
C1061 VPB.n599 VNB 0.21fF
C1062 VPB.n600 VNB 0.02fF
C1063 VPB.n601 VNB 0.01fF
C1064 VPB.n602 VNB 0.02fF
C1065 VPB.n603 VNB 0.28fF
C1066 VPB.n604 VNB 0.02fF
C1067 VPB.n605 VNB 0.02fF
C1068 VPB.n606 VNB 0.02fF
C1069 VPB.n607 VNB 0.28fF
C1070 VPB.n608 VNB 0.01fF
C1071 VPB.n609 VNB 0.02fF
C1072 VPB.n610 VNB 0.04fF
C1073 VPB.n611 VNB 0.02fF
C1074 VPB.n612 VNB 0.02fF
C1075 VPB.n613 VNB 0.02fF
C1076 VPB.n614 VNB 0.04fF
C1077 VPB.n615 VNB 0.02fF
C1078 VPB.n616 VNB 0.24fF
C1079 VPB.n617 VNB 0.04fF
C1080 VPB.n619 VNB 0.02fF
C1081 VPB.n620 VNB 0.02fF
C1082 VPB.n621 VNB 0.02fF
C1083 VPB.n622 VNB 0.02fF
C1084 VPB.n624 VNB 0.02fF
C1085 VPB.n625 VNB 0.02fF
C1086 VPB.n626 VNB 0.02fF
C1087 VPB.n628 VNB 0.28fF
C1088 VPB.n630 VNB 0.03fF
C1089 VPB.n631 VNB 0.02fF
C1090 VPB.n632 VNB 0.03fF
C1091 VPB.n633 VNB 0.03fF
C1092 VPB.n634 VNB 0.28fF
C1093 VPB.n635 VNB 0.01fF
C1094 VPB.n636 VNB 0.02fF
C1095 VPB.n637 VNB 0.04fF
C1096 VPB.n638 VNB 0.05fF
C1097 VPB.n639 VNB 0.24fF
C1098 VPB.n640 VNB 0.02fF
C1099 VPB.n641 VNB 0.01fF
C1100 VPB.n642 VNB 0.02fF
C1101 VPB.n643 VNB 0.14fF
C1102 VPB.n644 VNB 0.16fF
C1103 VPB.n645 VNB 0.02fF
C1104 VPB.n646 VNB 0.02fF
C1105 VPB.n647 VNB 0.02fF
C1106 VPB.n648 VNB 0.10fF
C1107 VPB.n649 VNB 0.02fF
C1108 VPB.n650 VNB 0.14fF
C1109 VPB.n651 VNB 0.15fF
C1110 VPB.n652 VNB 0.02fF
C1111 VPB.n653 VNB 0.02fF
C1112 VPB.n654 VNB 0.02fF
C1113 VPB.n655 VNB 0.14fF
C1114 VPB.n656 VNB 0.15fF
C1115 VPB.n657 VNB 0.02fF
C1116 VPB.n658 VNB 0.02fF
C1117 VPB.n659 VNB 0.02fF
C1118 VPB.n660 VNB 0.14fF
C1119 VPB.n661 VNB 0.16fF
C1120 VPB.n662 VNB 0.02fF
C1121 VPB.n663 VNB 0.02fF
C1122 VPB.n664 VNB 0.02fF
C1123 VPB.n665 VNB 0.06fF
C1124 VPB.n666 VNB 0.24fF
C1125 VPB.n667 VNB 0.02fF
C1126 VPB.n668 VNB 0.01fF
C1127 VPB.n669 VNB 0.02fF
C1128 VPB.n670 VNB 0.28fF
C1129 VPB.n671 VNB 0.01fF
C1130 VPB.n672 VNB 0.02fF
C1131 VPB.n673 VNB 0.04fF
C1132 VPB.n674 VNB 0.02fF
C1133 VPB.n675 VNB 0.02fF
C1134 VPB.n676 VNB 0.02fF
C1135 VPB.n677 VNB 0.04fF
C1136 VPB.n678 VNB 0.02fF
C1137 VPB.n679 VNB 0.24fF
C1138 VPB.n680 VNB 0.04fF
C1139 VPB.n682 VNB 0.02fF
C1140 VPB.n683 VNB 0.02fF
C1141 VPB.n684 VNB 0.02fF
C1142 VPB.n685 VNB 0.02fF
C1143 VPB.n687 VNB 0.02fF
C1144 VPB.n688 VNB 0.02fF
C1145 VPB.n689 VNB 0.02fF
C1146 VPB.n691 VNB 0.28fF
C1147 VPB.n693 VNB 0.03fF
C1148 VPB.n694 VNB 0.02fF
C1149 VPB.n695 VNB 0.03fF
C1150 VPB.n696 VNB 0.03fF
C1151 VPB.n697 VNB 0.28fF
C1152 VPB.n698 VNB 0.01fF
C1153 VPB.n699 VNB 0.02fF
C1154 VPB.n700 VNB 0.04fF
C1155 VPB.n701 VNB 0.28fF
C1156 VPB.n702 VNB 0.02fF
C1157 VPB.n703 VNB 0.02fF
C1158 VPB.n704 VNB 0.02fF
C1159 VPB.n705 VNB 0.05fF
C1160 VPB.n706 VNB 0.21fF
C1161 VPB.n707 VNB 0.02fF
C1162 VPB.n708 VNB 0.01fF
C1163 VPB.n709 VNB 0.02fF
C1164 VPB.n710 VNB 0.14fF
C1165 VPB.n711 VNB 0.16fF
C1166 VPB.n712 VNB 0.02fF
C1167 VPB.n713 VNB 0.02fF
C1168 VPB.n714 VNB 0.02fF
C1169 VPB.n715 VNB 0.10fF
C1170 VPB.n716 VNB 0.02fF
C1171 VPB.n717 VNB 0.14fF
C1172 VPB.n718 VNB 0.16fF
C1173 VPB.n719 VNB 0.02fF
C1174 VPB.n720 VNB 0.02fF
C1175 VPB.n721 VNB 0.02fF
C1176 VPB.n722 VNB 0.14fF
C1177 VPB.n723 VNB 0.15fF
C1178 VPB.n724 VNB 0.02fF
C1179 VPB.n725 VNB 0.02fF
C1180 VPB.n726 VNB 0.02fF
C1181 VPB.n727 VNB 0.14fF
C1182 VPB.n728 VNB 0.15fF
C1183 VPB.n729 VNB 0.02fF
C1184 VPB.n730 VNB 0.02fF
C1185 VPB.n731 VNB 0.02fF
C1186 VPB.n732 VNB 0.10fF
C1187 VPB.n733 VNB 0.02fF
C1188 VPB.n734 VNB 0.14fF
C1189 VPB.n735 VNB 0.16fF
C1190 VPB.n736 VNB 0.02fF
C1191 VPB.n737 VNB 0.02fF
C1192 VPB.n738 VNB 0.02fF
C1193 VPB.n739 VNB 0.14fF
C1194 VPB.n740 VNB 0.16fF
C1195 VPB.n741 VNB 0.02fF
C1196 VPB.n742 VNB 0.02fF
C1197 VPB.n743 VNB 0.02fF
C1198 VPB.n744 VNB 0.06fF
C1199 VPB.n745 VNB 0.21fF
C1200 VPB.n746 VNB 0.02fF
C1201 VPB.n747 VNB 0.01fF
C1202 VPB.n748 VNB 0.02fF
C1203 VPB.n749 VNB 0.28fF
C1204 VPB.n750 VNB 0.02fF
C1205 VPB.n751 VNB 0.02fF
C1206 VPB.n752 VNB 0.02fF
C1207 VPB.n753 VNB 0.28fF
C1208 VPB.n754 VNB 0.01fF
C1209 VPB.n755 VNB 0.02fF
C1210 VPB.n756 VNB 0.04fF
C1211 VPB.n757 VNB 0.02fF
C1212 VPB.n758 VNB 0.02fF
C1213 VPB.n759 VNB 0.02fF
C1214 VPB.n760 VNB 0.04fF
C1215 VPB.n761 VNB 0.02fF
C1216 VPB.n762 VNB 0.24fF
C1217 VPB.n763 VNB 0.04fF
C1218 VPB.n765 VNB 0.02fF
C1219 VPB.n766 VNB 0.02fF
C1220 VPB.n767 VNB 0.02fF
C1221 VPB.n768 VNB 0.02fF
C1222 VPB.n770 VNB 0.02fF
C1223 VPB.n771 VNB 0.02fF
C1224 VPB.n772 VNB 0.02fF
C1225 VPB.n774 VNB 0.28fF
C1226 VPB.n776 VNB 0.03fF
C1227 VPB.n777 VNB 0.02fF
C1228 VPB.n778 VNB 0.03fF
C1229 VPB.n779 VNB 0.03fF
C1230 VPB.n780 VNB 0.28fF
C1231 VPB.n781 VNB 0.01fF
C1232 VPB.n782 VNB 0.02fF
C1233 VPB.n783 VNB 0.04fF
C1234 VPB.n784 VNB 0.05fF
C1235 VPB.n785 VNB 0.24fF
C1236 VPB.n786 VNB 0.02fF
C1237 VPB.n787 VNB 0.01fF
C1238 VPB.n788 VNB 0.02fF
C1239 VPB.n789 VNB 0.14fF
C1240 VPB.n790 VNB 0.16fF
C1241 VPB.n791 VNB 0.02fF
C1242 VPB.n792 VNB 0.02fF
C1243 VPB.n793 VNB 0.02fF
C1244 VPB.n794 VNB 0.10fF
C1245 VPB.n795 VNB 0.02fF
C1246 VPB.n796 VNB 0.14fF
C1247 VPB.n797 VNB 0.15fF
C1248 VPB.n798 VNB 0.02fF
C1249 VPB.n799 VNB 0.02fF
C1250 VPB.n800 VNB 0.02fF
C1251 VPB.n801 VNB 0.14fF
C1252 VPB.n802 VNB 0.15fF
C1253 VPB.n803 VNB 0.02fF
C1254 VPB.n804 VNB 0.02fF
C1255 VPB.n805 VNB 0.02fF
C1256 VPB.n806 VNB 0.14fF
C1257 VPB.n807 VNB 0.16fF
C1258 VPB.n808 VNB 0.02fF
C1259 VPB.n809 VNB 0.02fF
C1260 VPB.n810 VNB 0.02fF
C1261 VPB.n811 VNB 0.06fF
C1262 VPB.n812 VNB 0.24fF
C1263 VPB.n813 VNB 0.02fF
C1264 VPB.n814 VNB 0.01fF
C1265 VPB.n815 VNB 0.02fF
C1266 VPB.n816 VNB 0.28fF
C1267 VPB.n817 VNB 0.01fF
C1268 VPB.n818 VNB 0.02fF
C1269 VPB.n819 VNB 0.04fF
C1270 VPB.n820 VNB 0.02fF
C1271 VPB.n821 VNB 0.02fF
C1272 VPB.n822 VNB 0.02fF
C1273 VPB.n823 VNB 0.04fF
C1274 VPB.n824 VNB 0.02fF
C1275 VPB.n825 VNB 0.20fF
C1276 VPB.n826 VNB 0.04fF
C1277 VPB.n828 VNB 0.02fF
C1278 VPB.n829 VNB 0.02fF
C1279 VPB.n830 VNB 0.02fF
C1280 VPB.n831 VNB 0.02fF
C1281 VPB.n833 VNB 0.02fF
C1282 VPB.n834 VNB 0.02fF
C1283 VPB.n835 VNB 0.02fF
C1284 VPB.n837 VNB 0.28fF
C1285 VPB.n839 VNB 0.03fF
C1286 VPB.n840 VNB 0.02fF
C1287 VPB.n841 VNB 0.03fF
C1288 VPB.n842 VNB 0.03fF
C1289 VPB.n843 VNB 0.28fF
C1290 VPB.n844 VNB 0.01fF
C1291 VPB.n845 VNB 0.02fF
C1292 VPB.n846 VNB 0.04fF
C1293 VPB.n847 VNB 0.05fF
C1294 VPB.n848 VNB 0.24fF
C1295 VPB.n849 VNB 0.02fF
C1296 VPB.n850 VNB 0.01fF
C1297 VPB.n851 VNB 0.02fF
C1298 VPB.n852 VNB 0.14fF
C1299 VPB.n853 VNB 0.16fF
C1300 VPB.n854 VNB 0.02fF
C1301 VPB.n855 VNB 0.02fF
C1302 VPB.n856 VNB 0.02fF
C1303 VPB.n857 VNB 0.10fF
C1304 VPB.n858 VNB 0.02fF
C1305 VPB.n859 VNB 0.14fF
C1306 VPB.n860 VNB 0.15fF
C1307 VPB.n861 VNB 0.02fF
C1308 VPB.n862 VNB 0.02fF
C1309 VPB.n863 VNB 0.02fF
C1310 VPB.n864 VNB 0.14fF
C1311 VPB.n865 VNB 0.15fF
C1312 VPB.n866 VNB 0.02fF
C1313 VPB.n867 VNB 0.02fF
C1314 VPB.n868 VNB 0.02fF
C1315 VPB.n869 VNB 0.14fF
C1316 VPB.n870 VNB 0.16fF
C1317 VPB.n871 VNB 0.02fF
C1318 VPB.n872 VNB 0.02fF
C1319 VPB.n873 VNB 0.02fF
C1320 VPB.n874 VNB 0.06fF
C1321 VPB.n875 VNB 0.24fF
C1322 VPB.n876 VNB 0.02fF
C1323 VPB.n877 VNB 0.01fF
C1324 VPB.n878 VNB 0.02fF
C1325 VPB.n879 VNB 0.28fF
C1326 VPB.n880 VNB 0.01fF
C1327 VPB.n881 VNB 0.02fF
C1328 VPB.n882 VNB 0.04fF
C1329 VPB.n883 VNB 0.02fF
C1330 VPB.n884 VNB 0.02fF
C1331 VPB.n885 VNB 0.02fF
C1332 VPB.n886 VNB 0.04fF
C1333 VPB.n887 VNB 0.02fF
C1334 VPB.n888 VNB 0.24fF
C1335 VPB.n889 VNB 0.04fF
C1336 VPB.n891 VNB 0.02fF
C1337 VPB.n892 VNB 0.02fF
C1338 VPB.n893 VNB 0.02fF
C1339 VPB.n894 VNB 0.02fF
C1340 VPB.n896 VNB 0.02fF
C1341 VPB.n897 VNB 0.02fF
C1342 VPB.n898 VNB 0.02fF
C1343 VPB.n900 VNB 0.28fF
C1344 VPB.n902 VNB 0.03fF
C1345 VPB.n903 VNB 0.02fF
C1346 VPB.n904 VNB 0.03fF
C1347 VPB.n905 VNB 0.03fF
C1348 VPB.n906 VNB 0.28fF
C1349 VPB.n907 VNB 0.01fF
C1350 VPB.n908 VNB 0.02fF
C1351 VPB.n909 VNB 0.04fF
C1352 VPB.n910 VNB 0.28fF
C1353 VPB.n911 VNB 0.02fF
C1354 VPB.n912 VNB 0.02fF
C1355 VPB.n913 VNB 0.02fF
C1356 VPB.n914 VNB 0.05fF
C1357 VPB.n915 VNB 0.21fF
C1358 VPB.n916 VNB 0.02fF
C1359 VPB.n917 VNB 0.01fF
C1360 VPB.n918 VNB 0.02fF
C1361 VPB.n919 VNB 0.14fF
C1362 VPB.n920 VNB 0.16fF
C1363 VPB.n921 VNB 0.02fF
C1364 VPB.n922 VNB 0.02fF
C1365 VPB.n923 VNB 0.02fF
C1366 VPB.n924 VNB 0.10fF
C1367 VPB.n925 VNB 0.02fF
C1368 VPB.n926 VNB 0.14fF
C1369 VPB.n927 VNB 0.16fF
C1370 VPB.n928 VNB 0.02fF
C1371 VPB.n929 VNB 0.02fF
C1372 VPB.n930 VNB 0.02fF
C1373 VPB.n931 VNB 0.14fF
C1374 VPB.n932 VNB 0.15fF
C1375 VPB.n933 VNB 0.02fF
C1376 VPB.n934 VNB 0.02fF
C1377 VPB.n935 VNB 0.02fF
C1378 VPB.n936 VNB 0.14fF
C1379 VPB.n937 VNB 0.15fF
C1380 VPB.n938 VNB 0.02fF
C1381 VPB.n939 VNB 0.02fF
C1382 VPB.n940 VNB 0.02fF
C1383 VPB.n941 VNB 0.10fF
C1384 VPB.n942 VNB 0.02fF
C1385 VPB.n943 VNB 0.14fF
C1386 VPB.n944 VNB 0.16fF
C1387 VPB.n945 VNB 0.02fF
C1388 VPB.n946 VNB 0.02fF
C1389 VPB.n947 VNB 0.02fF
C1390 VPB.n948 VNB 0.14fF
C1391 VPB.n949 VNB 0.16fF
C1392 VPB.n950 VNB 0.02fF
C1393 VPB.n951 VNB 0.02fF
C1394 VPB.n952 VNB 0.02fF
C1395 VPB.n953 VNB 0.06fF
C1396 VPB.n954 VNB 0.21fF
C1397 VPB.n955 VNB 0.02fF
C1398 VPB.n956 VNB 0.01fF
C1399 VPB.n957 VNB 0.02fF
C1400 VPB.n958 VNB 0.28fF
C1401 VPB.n959 VNB 0.02fF
C1402 VPB.n960 VNB 0.02fF
C1403 VPB.n961 VNB 0.02fF
C1404 VPB.n962 VNB 0.28fF
C1405 VPB.n963 VNB 0.01fF
C1406 VPB.n964 VNB 0.02fF
C1407 VPB.n965 VNB 0.04fF
C1408 VPB.n966 VNB 0.02fF
C1409 VPB.n967 VNB 0.02fF
C1410 VPB.n968 VNB 0.02fF
C1411 VPB.n969 VNB 0.04fF
C1412 VPB.n970 VNB 0.02fF
C1413 VPB.n971 VNB 0.29fF
C1414 VPB.n972 VNB 0.04fF
C1415 VPB.n974 VNB 0.02fF
C1416 VPB.n975 VNB 0.02fF
C1417 VPB.n976 VNB 0.02fF
C1418 VPB.n977 VNB 0.02fF
C1419 VPB.n979 VNB 0.02fF
C1420 VPB.n980 VNB 0.02fF
C1421 VPB.n981 VNB 0.02fF
C1422 VPB.n983 VNB 0.28fF
C1423 VPB.n985 VNB 0.03fF
C1424 VPB.n986 VNB 0.02fF
C1425 VPB.n987 VNB 0.03fF
C1426 VPB.n988 VNB 0.03fF
C1427 VPB.n989 VNB 0.28fF
C1428 VPB.n990 VNB 0.01fF
C1429 VPB.n991 VNB 0.02fF
C1430 VPB.n992 VNB 0.04fF
C1431 VPB.n993 VNB 0.28fF
C1432 VPB.n994 VNB 0.02fF
C1433 VPB.n995 VNB 0.02fF
C1434 VPB.n996 VNB 0.02fF
C1435 VPB.n997 VNB 0.05fF
C1436 VPB.n998 VNB 0.21fF
C1437 VPB.n999 VNB 0.02fF
C1438 VPB.n1000 VNB 0.01fF
C1439 VPB.n1001 VNB 0.02fF
C1440 VPB.n1002 VNB 0.14fF
C1441 VPB.n1003 VNB 0.16fF
C1442 VPB.n1004 VNB 0.02fF
C1443 VPB.n1005 VNB 0.02fF
C1444 VPB.n1006 VNB 0.02fF
C1445 VPB.n1007 VNB 0.10fF
C1446 VPB.n1008 VNB 0.02fF
C1447 VPB.n1009 VNB 0.14fF
C1448 VPB.n1010 VNB 0.16fF
C1449 VPB.n1011 VNB 0.02fF
C1450 VPB.n1012 VNB 0.02fF
C1451 VPB.n1013 VNB 0.02fF
C1452 VPB.n1014 VNB 0.14fF
C1453 VPB.n1015 VNB 0.15fF
C1454 VPB.n1016 VNB 0.02fF
C1455 VPB.n1017 VNB 0.02fF
C1456 VPB.n1018 VNB 0.02fF
C1457 VPB.n1019 VNB 0.14fF
C1458 VPB.n1020 VNB 0.15fF
C1459 VPB.n1021 VNB 0.02fF
C1460 VPB.n1022 VNB 0.02fF
C1461 VPB.n1023 VNB 0.02fF
C1462 VPB.n1024 VNB 0.10fF
C1463 VPB.n1025 VNB 0.02fF
C1464 VPB.n1026 VNB 0.14fF
C1465 VPB.n1027 VNB 0.16fF
C1466 VPB.n1028 VNB 0.02fF
C1467 VPB.n1029 VNB 0.02fF
C1468 VPB.n1030 VNB 0.02fF
C1469 VPB.n1031 VNB 0.14fF
C1470 VPB.n1032 VNB 0.16fF
C1471 VPB.n1033 VNB 0.02fF
C1472 VPB.n1034 VNB 0.02fF
C1473 VPB.n1035 VNB 0.02fF
C1474 VPB.n1036 VNB 0.06fF
C1475 VPB.n1037 VNB 0.21fF
C1476 VPB.n1038 VNB 0.02fF
C1477 VPB.n1039 VNB 0.01fF
C1478 VPB.n1040 VNB 0.02fF
C1479 VPB.n1041 VNB 0.28fF
C1480 VPB.n1042 VNB 0.02fF
C1481 VPB.n1043 VNB 0.02fF
C1482 VPB.n1044 VNB 0.02fF
C1483 VPB.n1045 VNB 0.28fF
C1484 VPB.n1046 VNB 0.01fF
C1485 VPB.n1047 VNB 0.02fF
C1486 VPB.n1048 VNB 0.04fF
C1487 VPB.n1049 VNB 0.02fF
C1488 VPB.n1050 VNB 0.02fF
C1489 VPB.n1051 VNB 0.02fF
C1490 VPB.n1052 VNB 0.04fF
C1491 VPB.n1053 VNB 0.02fF
C1492 VPB.n1054 VNB 0.24fF
C1493 VPB.n1055 VNB 0.04fF
C1494 VPB.n1057 VNB 0.02fF
C1495 VPB.n1058 VNB 0.02fF
C1496 VPB.n1059 VNB 0.02fF
C1497 VPB.n1060 VNB 0.02fF
C1498 VPB.n1062 VNB 0.02fF
C1499 VPB.n1063 VNB 0.02fF
C1500 VPB.n1064 VNB 0.02fF
C1501 VPB.n1066 VNB 0.28fF
C1502 VPB.n1068 VNB 0.03fF
C1503 VPB.n1069 VNB 0.02fF
C1504 VPB.n1070 VNB 0.03fF
C1505 VPB.n1071 VNB 0.03fF
C1506 VPB.n1072 VNB 0.28fF
C1507 VPB.n1073 VNB 0.01fF
C1508 VPB.n1074 VNB 0.02fF
C1509 VPB.n1075 VNB 0.04fF
C1510 VPB.n1076 VNB 0.05fF
C1511 VPB.n1077 VNB 0.24fF
C1512 VPB.n1078 VNB 0.02fF
C1513 VPB.n1079 VNB 0.01fF
C1514 VPB.n1080 VNB 0.02fF
C1515 VPB.n1081 VNB 0.14fF
C1516 VPB.n1082 VNB 0.16fF
C1517 VPB.n1083 VNB 0.02fF
C1518 VPB.n1084 VNB 0.02fF
C1519 VPB.n1085 VNB 0.02fF
C1520 VPB.n1086 VNB 0.10fF
C1521 VPB.n1087 VNB 0.02fF
C1522 VPB.n1088 VNB 0.14fF
C1523 VPB.n1089 VNB 0.15fF
C1524 VPB.n1090 VNB 0.02fF
C1525 VPB.n1091 VNB 0.02fF
C1526 VPB.n1092 VNB 0.02fF
C1527 VPB.n1093 VNB 0.14fF
C1528 VPB.n1094 VNB 0.15fF
C1529 VPB.n1095 VNB 0.02fF
C1530 VPB.n1096 VNB 0.02fF
C1531 VPB.n1097 VNB 0.02fF
C1532 VPB.n1098 VNB 0.14fF
C1533 VPB.n1099 VNB 0.16fF
C1534 VPB.n1100 VNB 0.02fF
C1535 VPB.n1101 VNB 0.02fF
C1536 VPB.n1102 VNB 0.02fF
C1537 VPB.n1103 VNB 0.06fF
C1538 VPB.n1104 VNB 0.24fF
C1539 VPB.n1105 VNB 0.02fF
C1540 VPB.n1106 VNB 0.01fF
C1541 VPB.n1107 VNB 0.02fF
C1542 VPB.n1108 VNB 0.28fF
C1543 VPB.n1109 VNB 0.01fF
C1544 VPB.n1110 VNB 0.02fF
C1545 VPB.n1111 VNB 0.04fF
C1546 VPB.n1112 VNB 0.02fF
C1547 VPB.n1113 VNB 0.02fF
C1548 VPB.n1114 VNB 0.02fF
C1549 VPB.n1115 VNB 0.04fF
C1550 VPB.n1116 VNB 0.02fF
C1551 VPB.n1117 VNB 0.24fF
C1552 VPB.n1118 VNB 0.04fF
C1553 VPB.n1120 VNB 0.02fF
C1554 VPB.n1121 VNB 0.02fF
C1555 VPB.n1122 VNB 0.02fF
C1556 VPB.n1123 VNB 0.02fF
C1557 VPB.n1125 VNB 0.02fF
C1558 VPB.n1126 VNB 0.02fF
C1559 VPB.n1127 VNB 0.02fF
C1560 VPB.n1129 VNB 0.28fF
C1561 VPB.n1131 VNB 0.03fF
C1562 VPB.n1132 VNB 0.02fF
C1563 VPB.n1133 VNB 0.03fF
C1564 VPB.n1134 VNB 0.03fF
C1565 VPB.n1135 VNB 0.28fF
C1566 VPB.n1136 VNB 0.01fF
C1567 VPB.n1137 VNB 0.02fF
C1568 VPB.n1138 VNB 0.04fF
C1569 VPB.n1139 VNB 0.28fF
C1570 VPB.n1140 VNB 0.02fF
C1571 VPB.n1141 VNB 0.02fF
C1572 VPB.n1142 VNB 0.02fF
C1573 VPB.n1143 VNB 0.05fF
C1574 VPB.n1144 VNB 0.21fF
C1575 VPB.n1145 VNB 0.02fF
C1576 VPB.n1146 VNB 0.01fF
C1577 VPB.n1147 VNB 0.02fF
C1578 VPB.n1148 VNB 0.14fF
C1579 VPB.n1149 VNB 0.16fF
C1580 VPB.n1150 VNB 0.02fF
C1581 VPB.n1151 VNB 0.02fF
C1582 VPB.n1152 VNB 0.02fF
C1583 VPB.n1153 VNB 0.10fF
C1584 VPB.n1154 VNB 0.02fF
C1585 VPB.n1155 VNB 0.14fF
C1586 VPB.n1156 VNB 0.16fF
C1587 VPB.n1157 VNB 0.02fF
C1588 VPB.n1158 VNB 0.02fF
C1589 VPB.n1159 VNB 0.02fF
C1590 VPB.n1160 VNB 0.14fF
C1591 VPB.n1161 VNB 0.15fF
C1592 VPB.n1162 VNB 0.02fF
C1593 VPB.n1163 VNB 0.02fF
C1594 VPB.n1164 VNB 0.02fF
C1595 VPB.n1165 VNB 0.14fF
C1596 VPB.n1166 VNB 0.15fF
C1597 VPB.n1167 VNB 0.02fF
C1598 VPB.n1168 VNB 0.02fF
C1599 VPB.n1169 VNB 0.02fF
C1600 VPB.n1170 VNB 0.10fF
C1601 VPB.n1171 VNB 0.02fF
C1602 VPB.n1172 VNB 0.14fF
C1603 VPB.n1173 VNB 0.16fF
C1604 VPB.n1174 VNB 0.02fF
C1605 VPB.n1175 VNB 0.02fF
C1606 VPB.n1176 VNB 0.02fF
C1607 VPB.n1177 VNB 0.14fF
C1608 VPB.n1178 VNB 0.16fF
C1609 VPB.n1179 VNB 0.02fF
C1610 VPB.n1180 VNB 0.02fF
C1611 VPB.n1181 VNB 0.02fF
C1612 VPB.n1182 VNB 0.06fF
C1613 VPB.n1183 VNB 0.21fF
C1614 VPB.n1184 VNB 0.02fF
C1615 VPB.n1185 VNB 0.01fF
C1616 VPB.n1186 VNB 0.02fF
C1617 VPB.n1187 VNB 0.28fF
C1618 VPB.n1188 VNB 0.02fF
C1619 VPB.n1189 VNB 0.02fF
C1620 VPB.n1190 VNB 0.02fF
C1621 VPB.n1191 VNB 0.28fF
C1622 VPB.n1192 VNB 0.01fF
C1623 VPB.n1193 VNB 0.02fF
C1624 VPB.n1194 VNB 0.04fF
C1625 VPB.n1195 VNB 0.02fF
C1626 VPB.n1196 VNB 0.02fF
C1627 VPB.n1197 VNB 0.02fF
C1628 VPB.n1198 VNB 0.04fF
C1629 VPB.n1199 VNB 0.02fF
C1630 VPB.n1200 VNB 0.24fF
C1631 VPB.n1201 VNB 0.04fF
C1632 VPB.n1203 VNB 0.02fF
C1633 VPB.n1204 VNB 0.02fF
C1634 VPB.n1205 VNB 0.02fF
C1635 VPB.n1206 VNB 0.02fF
C1636 VPB.n1208 VNB 0.02fF
C1637 VPB.n1209 VNB 0.02fF
C1638 VPB.n1210 VNB 0.02fF
C1639 VPB.n1212 VNB 0.28fF
C1640 VPB.n1214 VNB 0.03fF
C1641 VPB.n1215 VNB 0.02fF
C1642 VPB.n1216 VNB 0.03fF
C1643 VPB.n1217 VNB 0.03fF
C1644 VPB.n1218 VNB 0.28fF
C1645 VPB.n1219 VNB 0.01fF
C1646 VPB.n1220 VNB 0.02fF
C1647 VPB.n1221 VNB 0.04fF
C1648 VPB.n1222 VNB 0.05fF
C1649 VPB.n1223 VNB 0.24fF
C1650 VPB.n1224 VNB 0.02fF
C1651 VPB.n1225 VNB 0.01fF
C1652 VPB.n1226 VNB 0.02fF
C1653 VPB.n1227 VNB 0.14fF
C1654 VPB.n1228 VNB 0.16fF
C1655 VPB.n1229 VNB 0.02fF
C1656 VPB.n1230 VNB 0.02fF
C1657 VPB.n1231 VNB 0.02fF
C1658 VPB.n1232 VNB 0.10fF
C1659 VPB.n1233 VNB 0.02fF
C1660 VPB.n1234 VNB 0.14fF
C1661 VPB.n1235 VNB 0.15fF
C1662 VPB.n1236 VNB 0.02fF
C1663 VPB.n1237 VNB 0.02fF
C1664 VPB.n1238 VNB 0.02fF
C1665 VPB.n1239 VNB 0.14fF
C1666 VPB.n1240 VNB 0.15fF
C1667 VPB.n1241 VNB 0.02fF
C1668 VPB.n1242 VNB 0.02fF
C1669 VPB.n1243 VNB 0.02fF
C1670 VPB.n1244 VNB 0.14fF
C1671 VPB.n1245 VNB 0.16fF
C1672 VPB.n1246 VNB 0.02fF
C1673 VPB.n1247 VNB 0.02fF
C1674 VPB.n1248 VNB 0.02fF
C1675 VPB.n1249 VNB 0.06fF
C1676 VPB.n1250 VNB 0.24fF
C1677 VPB.n1251 VNB 0.02fF
C1678 VPB.n1252 VNB 0.01fF
C1679 VPB.n1253 VNB 0.02fF
C1680 VPB.n1254 VNB 0.28fF
C1681 VPB.n1255 VNB 0.01fF
C1682 VPB.n1256 VNB 0.02fF
C1683 VPB.n1257 VNB 0.04fF
C1684 VPB.n1258 VNB 0.02fF
C1685 VPB.n1259 VNB 0.02fF
C1686 VPB.n1260 VNB 0.02fF
C1687 VPB.n1261 VNB 0.04fF
C1688 VPB.n1262 VNB 0.02fF
C1689 VPB.n1263 VNB 0.20fF
C1690 VPB.n1264 VNB 0.04fF
C1691 VPB.n1266 VNB 0.02fF
C1692 VPB.n1267 VNB 0.02fF
C1693 VPB.n1268 VNB 0.02fF
C1694 VPB.n1269 VNB 0.02fF
C1695 VPB.n1271 VNB 0.02fF
C1696 VPB.n1272 VNB 0.02fF
C1697 VPB.n1273 VNB 0.02fF
C1698 VPB.n1275 VNB 0.28fF
C1699 VPB.n1277 VNB 0.03fF
C1700 VPB.n1278 VNB 0.02fF
C1701 VPB.n1279 VNB 0.03fF
C1702 VPB.n1280 VNB 0.03fF
C1703 VPB.n1281 VNB 0.28fF
C1704 VPB.n1282 VNB 0.01fF
C1705 VPB.n1283 VNB 0.02fF
C1706 VPB.n1284 VNB 0.04fF
C1707 VPB.n1285 VNB 0.05fF
C1708 VPB.n1286 VNB 0.24fF
C1709 VPB.n1287 VNB 0.02fF
C1710 VPB.n1288 VNB 0.01fF
C1711 VPB.n1289 VNB 0.02fF
C1712 VPB.n1290 VNB 0.14fF
C1713 VPB.n1291 VNB 0.16fF
C1714 VPB.n1292 VNB 0.02fF
C1715 VPB.n1293 VNB 0.02fF
C1716 VPB.n1294 VNB 0.02fF
C1717 VPB.n1295 VNB 0.10fF
C1718 VPB.n1296 VNB 0.02fF
C1719 VPB.n1297 VNB 0.14fF
C1720 VPB.n1298 VNB 0.15fF
C1721 VPB.n1299 VNB 0.02fF
C1722 VPB.n1300 VNB 0.02fF
C1723 VPB.n1301 VNB 0.02fF
C1724 VPB.n1302 VNB 0.14fF
C1725 VPB.n1303 VNB 0.15fF
C1726 VPB.n1304 VNB 0.02fF
C1727 VPB.n1305 VNB 0.02fF
C1728 VPB.n1306 VNB 0.02fF
C1729 VPB.n1307 VNB 0.14fF
C1730 VPB.n1308 VNB 0.16fF
C1731 VPB.n1309 VNB 0.02fF
C1732 VPB.n1310 VNB 0.02fF
C1733 VPB.n1311 VNB 0.02fF
C1734 VPB.n1312 VNB 0.06fF
C1735 VPB.n1313 VNB 0.24fF
C1736 VPB.n1314 VNB 0.02fF
C1737 VPB.n1315 VNB 0.01fF
C1738 VPB.n1316 VNB 0.02fF
C1739 VPB.n1317 VNB 0.28fF
C1740 VPB.n1318 VNB 0.01fF
C1741 VPB.n1319 VNB 0.02fF
C1742 VPB.n1320 VNB 0.04fF
C1743 VPB.n1321 VNB 0.02fF
C1744 VPB.n1322 VNB 0.02fF
C1745 VPB.n1323 VNB 0.02fF
C1746 VPB.n1324 VNB 0.04fF
C1747 VPB.n1325 VNB 0.02fF
C1748 VPB.n1326 VNB 0.24fF
C1749 VPB.n1327 VNB 0.04fF
C1750 VPB.n1329 VNB 0.02fF
C1751 VPB.n1330 VNB 0.02fF
C1752 VPB.n1331 VNB 0.02fF
C1753 VPB.n1332 VNB 0.02fF
C1754 VPB.n1334 VNB 0.02fF
C1755 VPB.n1335 VNB 0.02fF
C1756 VPB.n1336 VNB 0.02fF
C1757 VPB.n1338 VNB 0.28fF
C1758 VPB.n1340 VNB 0.03fF
C1759 VPB.n1341 VNB 0.02fF
C1760 VPB.n1342 VNB 0.03fF
C1761 VPB.n1343 VNB 0.03fF
C1762 VPB.n1344 VNB 0.28fF
C1763 VPB.n1345 VNB 0.01fF
C1764 VPB.n1346 VNB 0.02fF
C1765 VPB.n1347 VNB 0.04fF
C1766 VPB.n1348 VNB 0.28fF
C1767 VPB.n1349 VNB 0.02fF
C1768 VPB.n1350 VNB 0.02fF
C1769 VPB.n1351 VNB 0.02fF
C1770 VPB.n1352 VNB 0.05fF
C1771 VPB.n1353 VNB 0.21fF
C1772 VPB.n1354 VNB 0.02fF
C1773 VPB.n1355 VNB 0.01fF
C1774 VPB.n1356 VNB 0.02fF
C1775 VPB.n1357 VNB 0.14fF
C1776 VPB.n1358 VNB 0.16fF
C1777 VPB.n1359 VNB 0.02fF
C1778 VPB.n1360 VNB 0.02fF
C1779 VPB.n1361 VNB 0.02fF
C1780 VPB.n1362 VNB 0.10fF
C1781 VPB.n1363 VNB 0.02fF
C1782 VPB.n1364 VNB 0.14fF
C1783 VPB.n1365 VNB 0.16fF
C1784 VPB.n1366 VNB 0.02fF
C1785 VPB.n1367 VNB 0.02fF
C1786 VPB.n1368 VNB 0.02fF
C1787 VPB.n1369 VNB 0.14fF
C1788 VPB.n1370 VNB 0.15fF
C1789 VPB.n1371 VNB 0.02fF
C1790 VPB.n1372 VNB 0.02fF
C1791 VPB.n1373 VNB 0.02fF
C1792 VPB.n1374 VNB 0.14fF
C1793 VPB.n1375 VNB 0.15fF
C1794 VPB.n1376 VNB 0.02fF
C1795 VPB.n1377 VNB 0.02fF
C1796 VPB.n1378 VNB 0.02fF
C1797 VPB.n1379 VNB 0.10fF
C1798 VPB.n1380 VNB 0.02fF
C1799 VPB.n1381 VNB 0.14fF
C1800 VPB.n1382 VNB 0.16fF
C1801 VPB.n1383 VNB 0.02fF
C1802 VPB.n1384 VNB 0.02fF
C1803 VPB.n1385 VNB 0.02fF
C1804 VPB.n1386 VNB 0.14fF
C1805 VPB.n1387 VNB 0.16fF
C1806 VPB.n1388 VNB 0.02fF
C1807 VPB.n1389 VNB 0.02fF
C1808 VPB.n1390 VNB 0.02fF
C1809 VPB.n1391 VNB 0.06fF
C1810 VPB.n1392 VNB 0.21fF
C1811 VPB.n1393 VNB 0.02fF
C1812 VPB.n1394 VNB 0.01fF
C1813 VPB.n1395 VNB 0.02fF
C1814 VPB.n1396 VNB 0.28fF
C1815 VPB.n1397 VNB 0.02fF
C1816 VPB.n1398 VNB 0.02fF
C1817 VPB.n1399 VNB 0.02fF
C1818 VPB.n1400 VNB 0.28fF
C1819 VPB.n1401 VNB 0.01fF
C1820 VPB.n1402 VNB 0.02fF
C1821 VPB.n1403 VNB 0.04fF
C1822 VPB.n1404 VNB 0.02fF
C1823 VPB.n1405 VNB 0.02fF
C1824 VPB.n1406 VNB 0.02fF
C1825 VPB.n1407 VNB 0.04fF
C1826 VPB.n1408 VNB 0.02fF
C1827 VPB.n1409 VNB 0.29fF
C1828 VPB.n1410 VNB 0.04fF
C1829 VPB.n1412 VNB 0.02fF
C1830 VPB.n1413 VNB 0.02fF
C1831 VPB.n1414 VNB 0.02fF
C1832 VPB.n1415 VNB 0.02fF
C1833 VPB.n1417 VNB 0.02fF
C1834 VPB.n1418 VNB 0.02fF
C1835 VPB.n1419 VNB 0.02fF
C1836 VPB.n1421 VNB 0.28fF
C1837 VPB.n1423 VNB 0.03fF
C1838 VPB.n1424 VNB 0.02fF
C1839 VPB.n1425 VNB 0.03fF
C1840 VPB.n1426 VNB 0.03fF
C1841 VPB.n1427 VNB 0.28fF
C1842 VPB.n1428 VNB 0.01fF
C1843 VPB.n1429 VNB 0.02fF
C1844 VPB.n1430 VNB 0.04fF
C1845 VPB.n1431 VNB 0.28fF
C1846 VPB.n1432 VNB 0.02fF
C1847 VPB.n1433 VNB 0.02fF
C1848 VPB.n1434 VNB 0.02fF
C1849 VPB.n1435 VNB 0.05fF
C1850 VPB.n1436 VNB 0.21fF
C1851 VPB.n1437 VNB 0.02fF
C1852 VPB.n1438 VNB 0.01fF
C1853 VPB.n1439 VNB 0.02fF
C1854 VPB.n1440 VNB 0.14fF
C1855 VPB.n1441 VNB 0.16fF
C1856 VPB.n1442 VNB 0.02fF
C1857 VPB.n1443 VNB 0.02fF
C1858 VPB.n1444 VNB 0.02fF
C1859 VPB.n1445 VNB 0.10fF
C1860 VPB.n1446 VNB 0.02fF
C1861 VPB.n1447 VNB 0.14fF
C1862 VPB.n1448 VNB 0.16fF
C1863 VPB.n1449 VNB 0.02fF
C1864 VPB.n1450 VNB 0.02fF
C1865 VPB.n1451 VNB 0.02fF
C1866 VPB.n1452 VNB 0.14fF
C1867 VPB.n1453 VNB 0.15fF
C1868 VPB.n1454 VNB 0.02fF
C1869 VPB.n1455 VNB 0.02fF
C1870 VPB.n1456 VNB 0.02fF
C1871 VPB.n1457 VNB 0.14fF
C1872 VPB.n1458 VNB 0.15fF
C1873 VPB.n1459 VNB 0.02fF
C1874 VPB.n1460 VNB 0.02fF
C1875 VPB.n1461 VNB 0.02fF
C1876 VPB.n1462 VNB 0.10fF
C1877 VPB.n1463 VNB 0.02fF
C1878 VPB.n1464 VNB 0.14fF
C1879 VPB.n1465 VNB 0.16fF
C1880 VPB.n1466 VNB 0.02fF
C1881 VPB.n1467 VNB 0.02fF
C1882 VPB.n1468 VNB 0.02fF
C1883 VPB.n1469 VNB 0.14fF
C1884 VPB.n1470 VNB 0.16fF
C1885 VPB.n1471 VNB 0.02fF
C1886 VPB.n1472 VNB 0.02fF
C1887 VPB.n1473 VNB 0.02fF
C1888 VPB.n1474 VNB 0.06fF
C1889 VPB.n1475 VNB 0.21fF
C1890 VPB.n1476 VNB 0.02fF
C1891 VPB.n1477 VNB 0.01fF
C1892 VPB.n1478 VNB 0.02fF
C1893 VPB.n1479 VNB 0.28fF
C1894 VPB.n1480 VNB 0.02fF
C1895 VPB.n1481 VNB 0.02fF
C1896 VPB.n1482 VNB 0.02fF
C1897 VPB.n1483 VNB 0.28fF
C1898 VPB.n1484 VNB 0.01fF
C1899 VPB.n1485 VNB 0.02fF
C1900 VPB.n1486 VNB 0.04fF
C1901 VPB.n1487 VNB 0.04fF
C1902 VPB.n1488 VNB 0.02fF
C1903 VPB.n1489 VNB 0.02fF
C1904 VPB.n1490 VNB 0.02fF
C1905 VPB.n1491 VNB 0.02fF
C1906 VPB.n1492 VNB 0.10fF
C1907 VPB.n1493 VNB 0.00fF
C1908 VPB.n1494 VNB 0.04fF
C1909 VPB.n1495 VNB 0.02fF
C1910 VPB.n1496 VNB 0.02fF
C1911 VPB.n1497 VNB 0.02fF
C1912 VPB.n1498 VNB 0.04fF
C1913 VPB.n1499 VNB 0.04fF
C1914 VPB.n1501 VNB 0.43fF
C1915 a_5227_383.n0 VNB 0.07fF
C1916 a_5227_383.n1 VNB 0.90fF
C1917 a_5227_383.n2 VNB 0.90fF
C1918 a_5227_383.n3 VNB 1.05fF
C1919 a_5227_383.n4 VNB 0.33fF
C1920 a_5227_383.n5 VNB 0.43fF
C1921 a_5227_383.n6 VNB 0.54fF
C1922 a_5227_383.n7 VNB 0.78fF
C1923 a_5227_383.n8 VNB 0.48fF
C1924 a_5227_383.t12 VNB 0.95fF
C1925 a_5227_383.n9 VNB 0.67fF
C1926 a_5227_383.n10 VNB 4.19fF
C1927 a_5227_383.n11 VNB 0.74fF
C1928 a_5227_383.n12 VNB 0.06fF
C1929 a_5227_383.n13 VNB 0.58fF
C1930 a_5227_383.n14 VNB 0.09fF
C1931 a_6789_1004.n0 VNB 0.56fF
C1932 a_6789_1004.n1 VNB 0.56fF
C1933 a_6789_1004.n2 VNB 0.65fF
C1934 a_6789_1004.n3 VNB 0.21fF
C1935 a_6789_1004.n4 VNB 0.39fF
C1936 a_6789_1004.n5 VNB 0.46fF
C1937 a_6789_1004.n6 VNB 0.57fF
C1938 a_6789_1004.n7 VNB 0.66fF
C1939 a_6789_1004.n8 VNB 0.09fF
C1940 a_6789_1004.n9 VNB 0.22fF
C1941 a_6789_1004.n10 VNB 0.05fF
C1942 a_6884_182.n0 VNB 0.02fF
C1943 a_6884_182.n1 VNB 0.07fF
C1944 a_6884_182.n2 VNB 0.13fF
C1945 a_6884_182.n3 VNB 0.09fF
C1946 a_6884_182.t1 VNB 0.25fF
C1947 a_6884_182.n4 VNB 0.05fF
C1948 a_6884_182.n5 VNB 0.06fF
C1949 a_6884_182.n6 VNB 0.07fF
C1950 a_6884_182.n7 VNB 0.07fF
C1951 a_6884_182.n8 VNB 0.03fF
C1952 a_6884_182.n9 VNB 0.01fF
C1953 a_6884_182.n10 VNB 0.11fF
C1954 a_6884_182.n11 VNB 0.02fF
C1955 a_6884_182.n12 VNB 0.05fF
C1956 a_6884_182.n13 VNB 0.03fF
C1957 a_6149_943.n0 VNB 0.07fF
C1958 a_6149_943.n1 VNB 0.96fF
C1959 a_6149_943.n2 VNB 1.14fF
C1960 a_6149_943.n3 VNB 0.52fF
C1961 a_6149_943.n4 VNB 0.65fF
C1962 a_6149_943.t10 VNB 0.99fF
C1963 a_6149_943.n5 VNB 0.73fF
C1964 a_6149_943.n6 VNB 0.65fF
C1965 a_6149_943.t5 VNB 0.98fF
C1966 a_6149_943.n7 VNB 0.66fF
C1967 a_6149_943.n8 VNB 0.65fF
C1968 a_6149_943.t13 VNB 0.99fF
C1969 a_6149_943.n9 VNB 0.69fF
C1970 a_6149_943.n10 VNB 2.06fF
C1971 a_6149_943.n11 VNB 2.79fF
C1972 a_6149_943.n12 VNB 0.76fF
C1973 a_6149_943.n13 VNB 0.06fF
C1974 a_6149_943.n14 VNB 0.56fF
C1975 a_6149_943.n15 VNB 0.10fF
.ends
