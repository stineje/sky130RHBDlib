* SPICE3 file created from DFFRNQNX1.ext - technology: sky130A

.subckt DFFRNQNX1 QN D CLK RN VPB VNB
M1000 QN a_4151_943.t7 a_3924_182.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1001 VPB.t29 a_147_159.t7 a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_599_943.t4 a_1304_166# VPB.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t20 a_599_943.t7 a_2141_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPB.t13 CLK a_277_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t24 a_277_1004.t8 QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=1.74p ps=13.74u
M1006 a_599_943.t1 RN VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 QN a_4151_943.t5 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_147_159.t4 CLK VPB.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_4151_943.t1 QN VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VNB QN a_4626_73.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1011 VNB a_147_159.t14 a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t0 a_599_943.t9 a_277_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPB.t27 a_147_159.t8 a_2141_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VNB a_599_943.t8 a_2036_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPB.t17 a_2141_1004.t6 a_147_159.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_147_159.t0 RN VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_4151_943.t3 a_147_159.t9 VPB.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_277_1004.t5 a_147_159.t10 VPB.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VNB a_277_1004.t7 a_3643_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPB.t22 a_277_1004.t10 a_599_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPB.t7 RN a_599_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t16 a_4151_943.t6 QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VNB a_2141_1004.t5 a_2681_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_277_1004.t3 CLK VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2141_1004.t0 a_599_943.t10 VPB.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 QN a_277_1004.t11 VPB.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPB.t11 a_1304_166# a_599_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPB.t6 RN QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_599_943.t5 a_277_1004.t12 VPB.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_277_1004.t6 a_599_943.t11 VPB.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2141_1004.t2 a_147_159.t13 VPB.t26 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 QN RN VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_147_159.t6 a_2141_1004.t7 VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VNB a_277_1004.t9 a_1053_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPB.t14 CLK a_147_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPB.t3 QN a_4151_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPB.t8 RN a_147_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPB.t30 a_147_159.t15 a_4151_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB a_1304_166# 0.05fF
C1 VPB RN 0.17fF
C2 VPB CLK 0.75fF
C3 a_1304_166# RN 0.18fF
C4 VPB QN 1.85fF
C5 a_1304_166# CLK 0.04fF
C6 CLK RN 0.26fF
C7 RN QN 0.12fF
R0 a_147_159.n10 a_147_159.t7 512.525
R1 a_147_159.n8 a_147_159.t8 472.359
R2 a_147_159.n6 a_147_159.t15 472.359
R3 a_147_159.n8 a_147_159.t13 384.527
R4 a_147_159.n6 a_147_159.t9 384.527
R5 a_147_159.n10 a_147_159.t10 371.139
R6 a_147_159.n11 a_147_159.t14 324.268
R7 a_147_159.n9 a_147_159.t12 277.772
R8 a_147_159.n7 a_147_159.t11 277.772
R9 a_147_159.n16 a_147_159.n14 249.704
R10 a_147_159.n14 a_147_159.n5 127.74
R11 a_147_159.n11 a_147_159.n10 119.654
R12 a_147_159.n12 a_147_159.n11 83.572
R13 a_147_159.n13 a_147_159.n7 81.396
R14 a_147_159.n4 a_147_159.n3 79.232
R15 a_147_159.n12 a_147_159.n9 76
R16 a_147_159.n14 a_147_159.n13 76
R17 a_147_159.n9 a_147_159.n8 67.001
R18 a_147_159.n7 a_147_159.n6 67.001
R19 a_147_159.n5 a_147_159.n4 63.152
R20 a_147_159.n16 a_147_159.n15 30
R21 a_147_159.n17 a_147_159.n0 24.383
R22 a_147_159.n17 a_147_159.n16 23.684
R23 a_147_159.n5 a_147_159.n1 16.08
R24 a_147_159.n4 a_147_159.n2 16.08
R25 a_147_159.n1 a_147_159.t1 14.282
R26 a_147_159.n1 a_147_159.t0 14.282
R27 a_147_159.n2 a_147_159.t3 14.282
R28 a_147_159.n2 a_147_159.t4 14.282
R29 a_147_159.n3 a_147_159.t5 14.282
R30 a_147_159.n3 a_147_159.t6 14.282
R31 a_147_159.n13 a_147_159.n12 4.035
R32 a_277_1004.n7 a_277_1004.t10 512.525
R33 a_277_1004.n5 a_277_1004.t8 512.525
R34 a_277_1004.n7 a_277_1004.t12 371.139
R35 a_277_1004.n5 a_277_1004.t11 371.139
R36 a_277_1004.n8 a_277_1004.t9 297.715
R37 a_277_1004.n6 a_277_1004.t7 297.715
R38 a_277_1004.n12 a_277_1004.n10 229.673
R39 a_277_1004.n10 a_277_1004.n4 154.293
R40 a_277_1004.n8 a_277_1004.n7 146.207
R41 a_277_1004.n6 a_277_1004.n5 146.207
R42 a_277_1004.n9 a_277_1004.n6 85.476
R43 a_277_1004.n3 a_277_1004.n2 79.232
R44 a_277_1004.n10 a_277_1004.n9 77.315
R45 a_277_1004.n9 a_277_1004.n8 76
R46 a_277_1004.n4 a_277_1004.n3 63.152
R47 a_277_1004.n4 a_277_1004.n0 16.08
R48 a_277_1004.n3 a_277_1004.n1 16.08
R49 a_277_1004.n12 a_277_1004.n11 15.218
R50 a_277_1004.n0 a_277_1004.t0 14.282
R51 a_277_1004.n0 a_277_1004.t6 14.282
R52 a_277_1004.n1 a_277_1004.t2 14.282
R53 a_277_1004.n1 a_277_1004.t3 14.282
R54 a_277_1004.n2 a_277_1004.t4 14.282
R55 a_277_1004.n2 a_277_1004.t5 14.282
R56 a_277_1004.n13 a_277_1004.n12 12.014
R57 VPB VPB.n473 126.832
R58 VPB.n40 VPB.n38 94.117
R59 VPB.n395 VPB.n393 94.117
R60 VPB.n332 VPB.n330 94.117
R61 VPB.n129 VPB.n127 94.117
R62 VPB.n255 VPB.n253 94.117
R63 VPB.n268 VPB.n267 80.104
R64 VPB.n139 VPB.n138 80.104
R65 VPB.n408 VPB.n407 80.104
R66 VPB.n50 VPB.n49 80.104
R67 VPB.n216 VPB.n215 76
R68 VPB.n221 VPB.n220 76
R69 VPB.n226 VPB.n225 76
R70 VPB.n230 VPB.n229 76
R71 VPB.n257 VPB.n256 76
R72 VPB.n261 VPB.n260 76
R73 VPB.n266 VPB.n265 76
R74 VPB.n271 VPB.n270 76
R75 VPB.n278 VPB.n277 76
R76 VPB.n283 VPB.n282 76
R77 VPB.n288 VPB.n287 76
R78 VPB.n295 VPB.n294 76
R79 VPB.n300 VPB.n299 76
R80 VPB.n305 VPB.n304 76
R81 VPB.n309 VPB.n308 76
R82 VPB.n313 VPB.n312 76
R83 VPB.n328 VPB.n325 76
R84 VPB.n334 VPB.n333 76
R85 VPB.n339 VPB.n338 76
R86 VPB.n344 VPB.n343 76
R87 VPB.n351 VPB.n350 76
R88 VPB.n356 VPB.n355 76
R89 VPB.n361 VPB.n360 76
R90 VPB.n366 VPB.n365 76
R91 VPB.n370 VPB.n369 76
R92 VPB.n397 VPB.n396 76
R93 VPB.n401 VPB.n400 76
R94 VPB.n406 VPB.n405 76
R95 VPB.n411 VPB.n410 76
R96 VPB.n418 VPB.n417 76
R97 VPB.n423 VPB.n422 76
R98 VPB.n428 VPB.n427 76
R99 VPB.n435 VPB.n434 76
R100 VPB.n440 VPB.n439 76
R101 VPB.n445 VPB.n444 76
R102 VPB.n449 VPB.n448 76
R103 VPB.n453 VPB.n452 76
R104 VPB.n466 VPB.n465 76
R105 VPB.n297 VPB.n296 75.654
R106 VPB.n161 VPB.n160 75.654
R107 VPB.n437 VPB.n436 75.654
R108 VPB.n72 VPB.n71 75.654
R109 VPB.n22 VPB.n21 61.764
R110 VPB.n377 VPB.n376 61.764
R111 VPB.n88 VPB.n87 61.764
R112 VPB.n111 VPB.n110 61.764
R113 VPB.n237 VPB.n236 61.764
R114 VPB.n78 VPB.t28 55.106
R115 VPB.n441 VPB.t21 55.106
R116 VPB.n362 VPB.t19 55.106
R117 VPB.n167 VPB.t18 55.106
R118 VPB.n301 VPB.t23 55.106
R119 VPB.n222 VPB.t2 55.106
R120 VPB.n45 VPB.t0 55.106
R121 VPB.n402 VPB.t7 55.106
R122 VPB.n335 VPB.t27 55.106
R123 VPB.n134 VPB.t8 55.106
R124 VPB.n262 VPB.t16 55.106
R125 VPB.n205 VPB.t30 55.106
R126 VPB.n202 VPB.n201 48.952
R127 VPB.n275 VPB.n274 48.952
R128 VPB.n143 VPB.n142 48.952
R129 VPB.n341 VPB.n340 48.952
R130 VPB.n415 VPB.n414 48.952
R131 VPB.n54 VPB.n53 48.952
R132 VPB.n218 VPB.n217 44.502
R133 VPB.n292 VPB.n291 44.502
R134 VPB.n157 VPB.n156 44.502
R135 VPB.n358 VPB.n357 44.502
R136 VPB.n432 VPB.n431 44.502
R137 VPB.n68 VPB.n67 44.502
R138 VPB.n66 VPB.n14 40.824
R139 VPB.n57 VPB.n15 40.824
R140 VPB.n430 VPB.n429 40.824
R141 VPB.n413 VPB.n412 40.824
R142 VPB.n346 VPB.n345 40.824
R143 VPB.n155 VPB.n103 40.824
R144 VPB.n146 VPB.n104 40.824
R145 VPB.n290 VPB.n289 40.824
R146 VPB.n273 VPB.n272 40.824
R147 VPB.n196 VPB.n195 40.824
R148 VPB.n210 VPB.n209 35.118
R149 VPB.n470 VPB.n466 20.452
R150 VPB.n194 VPB.n191 20.452
R151 VPB.n198 VPB.n197 17.801
R152 VPB.n280 VPB.n279 17.801
R153 VPB.n148 VPB.n147 17.801
R154 VPB.n348 VPB.n347 17.801
R155 VPB.n420 VPB.n419 17.801
R156 VPB.n59 VPB.n58 17.801
R157 VPB.n14 VPB.t12 14.282
R158 VPB.n14 VPB.t29 14.282
R159 VPB.n15 VPB.t31 14.282
R160 VPB.n15 VPB.t13 14.282
R161 VPB.n429 VPB.t10 14.282
R162 VPB.n429 VPB.t22 14.282
R163 VPB.n412 VPB.t4 14.282
R164 VPB.n412 VPB.t11 14.282
R165 VPB.n345 VPB.t26 14.282
R166 VPB.n345 VPB.t20 14.282
R167 VPB.n103 VPB.t15 14.282
R168 VPB.n103 VPB.t17 14.282
R169 VPB.n104 VPB.t9 14.282
R170 VPB.n104 VPB.t14 14.282
R171 VPB.n289 VPB.t5 14.282
R172 VPB.n289 VPB.t24 14.282
R173 VPB.n272 VPB.t1 14.282
R174 VPB.n272 VPB.t6 14.282
R175 VPB.n195 VPB.t25 14.282
R176 VPB.n195 VPB.t3 14.282
R177 VPB.n194 VPB.n193 13.653
R178 VPB.n193 VPB.n192 13.653
R179 VPB.n208 VPB.n207 13.653
R180 VPB.n207 VPB.n206 13.653
R181 VPB.n204 VPB.n203 13.653
R182 VPB.n203 VPB.n202 13.653
R183 VPB.n200 VPB.n199 13.653
R184 VPB.n199 VPB.n198 13.653
R185 VPB.n215 VPB.n214 13.653
R186 VPB.n214 VPB.n213 13.653
R187 VPB.n220 VPB.n219 13.653
R188 VPB.n219 VPB.n218 13.653
R189 VPB.n225 VPB.n224 13.653
R190 VPB.n224 VPB.n223 13.653
R191 VPB.n229 VPB.n228 13.653
R192 VPB.n228 VPB.n227 13.653
R193 VPB.n256 VPB.n255 13.653
R194 VPB.n255 VPB.n254 13.653
R195 VPB.n260 VPB.n259 13.653
R196 VPB.n259 VPB.n258 13.653
R197 VPB.n265 VPB.n264 13.653
R198 VPB.n264 VPB.n263 13.653
R199 VPB.n270 VPB.n269 13.653
R200 VPB.n269 VPB.n268 13.653
R201 VPB.n277 VPB.n276 13.653
R202 VPB.n276 VPB.n275 13.653
R203 VPB.n282 VPB.n281 13.653
R204 VPB.n281 VPB.n280 13.653
R205 VPB.n287 VPB.n286 13.653
R206 VPB.n286 VPB.n285 13.653
R207 VPB.n294 VPB.n293 13.653
R208 VPB.n293 VPB.n292 13.653
R209 VPB.n299 VPB.n298 13.653
R210 VPB.n298 VPB.n297 13.653
R211 VPB.n304 VPB.n303 13.653
R212 VPB.n303 VPB.n302 13.653
R213 VPB.n308 VPB.n307 13.653
R214 VPB.n307 VPB.n306 13.653
R215 VPB.n312 VPB.n311 13.653
R216 VPB.n311 VPB.n310 13.653
R217 VPB.n130 VPB.n129 13.653
R218 VPB.n129 VPB.n128 13.653
R219 VPB.n133 VPB.n132 13.653
R220 VPB.n132 VPB.n131 13.653
R221 VPB.n137 VPB.n136 13.653
R222 VPB.n136 VPB.n135 13.653
R223 VPB.n141 VPB.n140 13.653
R224 VPB.n140 VPB.n139 13.653
R225 VPB.n145 VPB.n144 13.653
R226 VPB.n144 VPB.n143 13.653
R227 VPB.n150 VPB.n149 13.653
R228 VPB.n149 VPB.n148 13.653
R229 VPB.n154 VPB.n153 13.653
R230 VPB.n153 VPB.n152 13.653
R231 VPB.n159 VPB.n158 13.653
R232 VPB.n158 VPB.n157 13.653
R233 VPB.n163 VPB.n162 13.653
R234 VPB.n162 VPB.n161 13.653
R235 VPB.n166 VPB.n165 13.653
R236 VPB.n165 VPB.n164 13.653
R237 VPB.n170 VPB.n169 13.653
R238 VPB.n169 VPB.n168 13.653
R239 VPB.n328 VPB.n327 13.653
R240 VPB.n327 VPB.n326 13.653
R241 VPB.n333 VPB.n332 13.653
R242 VPB.n332 VPB.n331 13.653
R243 VPB.n338 VPB.n337 13.653
R244 VPB.n337 VPB.n336 13.653
R245 VPB.n343 VPB.n342 13.653
R246 VPB.n342 VPB.n341 13.653
R247 VPB.n350 VPB.n349 13.653
R248 VPB.n349 VPB.n348 13.653
R249 VPB.n355 VPB.n354 13.653
R250 VPB.n354 VPB.n353 13.653
R251 VPB.n360 VPB.n359 13.653
R252 VPB.n359 VPB.n358 13.653
R253 VPB.n365 VPB.n364 13.653
R254 VPB.n364 VPB.n363 13.653
R255 VPB.n369 VPB.n368 13.653
R256 VPB.n368 VPB.n367 13.653
R257 VPB.n396 VPB.n395 13.653
R258 VPB.n395 VPB.n394 13.653
R259 VPB.n400 VPB.n399 13.653
R260 VPB.n399 VPB.n398 13.653
R261 VPB.n405 VPB.n404 13.653
R262 VPB.n404 VPB.n403 13.653
R263 VPB.n410 VPB.n409 13.653
R264 VPB.n409 VPB.n408 13.653
R265 VPB.n417 VPB.n416 13.653
R266 VPB.n416 VPB.n415 13.653
R267 VPB.n422 VPB.n421 13.653
R268 VPB.n421 VPB.n420 13.653
R269 VPB.n427 VPB.n426 13.653
R270 VPB.n426 VPB.n425 13.653
R271 VPB.n434 VPB.n433 13.653
R272 VPB.n433 VPB.n432 13.653
R273 VPB.n439 VPB.n438 13.653
R274 VPB.n438 VPB.n437 13.653
R275 VPB.n444 VPB.n443 13.653
R276 VPB.n443 VPB.n442 13.653
R277 VPB.n448 VPB.n447 13.653
R278 VPB.n447 VPB.n446 13.653
R279 VPB.n452 VPB.n451 13.653
R280 VPB.n451 VPB.n450 13.653
R281 VPB.n41 VPB.n40 13.653
R282 VPB.n40 VPB.n39 13.653
R283 VPB.n44 VPB.n43 13.653
R284 VPB.n43 VPB.n42 13.653
R285 VPB.n48 VPB.n47 13.653
R286 VPB.n47 VPB.n46 13.653
R287 VPB.n52 VPB.n51 13.653
R288 VPB.n51 VPB.n50 13.653
R289 VPB.n56 VPB.n55 13.653
R290 VPB.n55 VPB.n54 13.653
R291 VPB.n61 VPB.n60 13.653
R292 VPB.n60 VPB.n59 13.653
R293 VPB.n65 VPB.n64 13.653
R294 VPB.n64 VPB.n63 13.653
R295 VPB.n70 VPB.n69 13.653
R296 VPB.n69 VPB.n68 13.653
R297 VPB.n74 VPB.n73 13.653
R298 VPB.n73 VPB.n72 13.653
R299 VPB.n77 VPB.n76 13.653
R300 VPB.n76 VPB.n75 13.653
R301 VPB.n81 VPB.n80 13.653
R302 VPB.n80 VPB.n79 13.653
R303 VPB.n466 VPB.n0 13.653
R304 VPB VPB.n0 13.653
R305 VPB.n213 VPB.n212 13.35
R306 VPB.n285 VPB.n284 13.35
R307 VPB.n152 VPB.n151 13.35
R308 VPB.n353 VPB.n352 13.35
R309 VPB.n425 VPB.n424 13.35
R310 VPB.n63 VPB.n62 13.35
R311 VPB.n470 VPB.n469 13.276
R312 VPB.n469 VPB.n467 13.276
R313 VPB.n36 VPB.n18 13.276
R314 VPB.n18 VPB.n16 13.276
R315 VPB.n391 VPB.n373 13.276
R316 VPB.n373 VPB.n371 13.276
R317 VPB.n102 VPB.n84 13.276
R318 VPB.n84 VPB.n82 13.276
R319 VPB.n125 VPB.n107 13.276
R320 VPB.n107 VPB.n105 13.276
R321 VPB.n251 VPB.n233 13.276
R322 VPB.n233 VPB.n231 13.276
R323 VPB.n204 VPB.n200 13.276
R324 VPB.n256 VPB.n252 13.276
R325 VPB.n130 VPB.n126 13.276
R326 VPB.n133 VPB.n130 13.276
R327 VPB.n141 VPB.n137 13.276
R328 VPB.n145 VPB.n141 13.276
R329 VPB.n154 VPB.n150 13.276
R330 VPB.n163 VPB.n159 13.276
R331 VPB.n166 VPB.n163 13.276
R332 VPB.n328 VPB.n170 13.276
R333 VPB.n329 VPB.n328 13.276
R334 VPB.n333 VPB.n329 13.276
R335 VPB.n396 VPB.n392 13.276
R336 VPB.n41 VPB.n37 13.276
R337 VPB.n44 VPB.n41 13.276
R338 VPB.n52 VPB.n48 13.276
R339 VPB.n56 VPB.n52 13.276
R340 VPB.n65 VPB.n61 13.276
R341 VPB.n74 VPB.n70 13.276
R342 VPB.n77 VPB.n74 13.276
R343 VPB.n466 VPB.n81 13.276
R344 VPB.n191 VPB.n173 13.276
R345 VPB.n173 VPB.n171 13.276
R346 VPB.n178 VPB.n176 12.796
R347 VPB.n178 VPB.n177 12.564
R348 VPB.n170 VPB.n167 12.558
R349 VPB.n81 VPB.n78 12.558
R350 VPB.n134 VPB.n133 12.2
R351 VPB.n45 VPB.n44 12.2
R352 VPB.n187 VPB.n186 12.198
R353 VPB.n184 VPB.n183 12.198
R354 VPB.n184 VPB.n181 12.198
R355 VPB.n205 VPB.n204 11.841
R356 VPB.n150 VPB.n146 9.329
R357 VPB.n61 VPB.n57 9.329
R358 VPB.n155 VPB.n154 8.97
R359 VPB.n66 VPB.n65 8.97
R360 VPB.n191 VPB.n190 7.5
R361 VPB.n176 VPB.n175 7.5
R362 VPB.n183 VPB.n182 7.5
R363 VPB.n181 VPB.n180 7.5
R364 VPB.n173 VPB.n172 7.5
R365 VPB.n188 VPB.n174 7.5
R366 VPB.n233 VPB.n232 7.5
R367 VPB.n246 VPB.n245 7.5
R368 VPB.n240 VPB.n239 7.5
R369 VPB.n242 VPB.n241 7.5
R370 VPB.n235 VPB.n234 7.5
R371 VPB.n251 VPB.n250 7.5
R372 VPB.n107 VPB.n106 7.5
R373 VPB.n120 VPB.n119 7.5
R374 VPB.n114 VPB.n113 7.5
R375 VPB.n116 VPB.n115 7.5
R376 VPB.n109 VPB.n108 7.5
R377 VPB.n125 VPB.n124 7.5
R378 VPB.n84 VPB.n83 7.5
R379 VPB.n97 VPB.n96 7.5
R380 VPB.n91 VPB.n90 7.5
R381 VPB.n93 VPB.n92 7.5
R382 VPB.n86 VPB.n85 7.5
R383 VPB.n102 VPB.n101 7.5
R384 VPB.n373 VPB.n372 7.5
R385 VPB.n386 VPB.n385 7.5
R386 VPB.n380 VPB.n379 7.5
R387 VPB.n382 VPB.n381 7.5
R388 VPB.n375 VPB.n374 7.5
R389 VPB.n391 VPB.n390 7.5
R390 VPB.n18 VPB.n17 7.5
R391 VPB.n31 VPB.n30 7.5
R392 VPB.n25 VPB.n24 7.5
R393 VPB.n27 VPB.n26 7.5
R394 VPB.n20 VPB.n19 7.5
R395 VPB.n36 VPB.n35 7.5
R396 VPB.n469 VPB.n468 7.5
R397 VPB.n12 VPB.n11 7.5
R398 VPB.n6 VPB.n5 7.5
R399 VPB.n8 VPB.n7 7.5
R400 VPB.n2 VPB.n1 7.5
R401 VPB.n471 VPB.n470 7.5
R402 VPB.n37 VPB.n36 7.176
R403 VPB.n392 VPB.n391 7.176
R404 VPB.n329 VPB.n102 7.176
R405 VPB.n126 VPB.n125 7.176
R406 VPB.n252 VPB.n251 7.176
R407 VPB.n247 VPB.n244 6.729
R408 VPB.n243 VPB.n240 6.729
R409 VPB.n238 VPB.n235 6.729
R410 VPB.n121 VPB.n118 6.729
R411 VPB.n117 VPB.n114 6.729
R412 VPB.n112 VPB.n109 6.729
R413 VPB.n98 VPB.n95 6.729
R414 VPB.n94 VPB.n91 6.729
R415 VPB.n89 VPB.n86 6.729
R416 VPB.n387 VPB.n384 6.729
R417 VPB.n383 VPB.n380 6.729
R418 VPB.n378 VPB.n375 6.729
R419 VPB.n32 VPB.n29 6.729
R420 VPB.n28 VPB.n25 6.729
R421 VPB.n23 VPB.n20 6.729
R422 VPB.n13 VPB.n10 6.729
R423 VPB.n9 VPB.n6 6.729
R424 VPB.n4 VPB.n2 6.729
R425 VPB.n238 VPB.n237 6.728
R426 VPB.n243 VPB.n242 6.728
R427 VPB.n247 VPB.n246 6.728
R428 VPB.n250 VPB.n249 6.728
R429 VPB.n112 VPB.n111 6.728
R430 VPB.n117 VPB.n116 6.728
R431 VPB.n121 VPB.n120 6.728
R432 VPB.n124 VPB.n123 6.728
R433 VPB.n89 VPB.n88 6.728
R434 VPB.n94 VPB.n93 6.728
R435 VPB.n98 VPB.n97 6.728
R436 VPB.n101 VPB.n100 6.728
R437 VPB.n378 VPB.n377 6.728
R438 VPB.n383 VPB.n382 6.728
R439 VPB.n387 VPB.n386 6.728
R440 VPB.n390 VPB.n389 6.728
R441 VPB.n23 VPB.n22 6.728
R442 VPB.n28 VPB.n27 6.728
R443 VPB.n32 VPB.n31 6.728
R444 VPB.n35 VPB.n34 6.728
R445 VPB.n4 VPB.n3 6.728
R446 VPB.n9 VPB.n8 6.728
R447 VPB.n13 VPB.n12 6.728
R448 VPB.n472 VPB.n471 6.728
R449 VPB.n200 VPB.n196 6.458
R450 VPB.n350 VPB.n346 6.458
R451 VPB.n190 VPB.n189 6.398
R452 VPB.n209 VPB.n194 6.112
R453 VPB.n209 VPB.n208 6.101
R454 VPB.n294 VPB.n290 4.305
R455 VPB.n159 VPB.n155 4.305
R456 VPB.n434 VPB.n430 4.305
R457 VPB.n70 VPB.n66 4.305
R458 VPB.n277 VPB.n273 3.947
R459 VPB.n146 VPB.n145 3.947
R460 VPB.n417 VPB.n413 3.947
R461 VPB.n57 VPB.n56 3.947
R462 VPB.n225 VPB.n222 1.794
R463 VPB.n365 VPB.n362 1.794
R464 VPB.n208 VPB.n205 1.435
R465 VPB.n338 VPB.n335 1.435
R466 VPB.n188 VPB.n179 1.402
R467 VPB.n188 VPB.n184 1.402
R468 VPB.n188 VPB.n185 1.402
R469 VPB.n188 VPB.n187 1.402
R470 VPB.n265 VPB.n262 1.076
R471 VPB.n137 VPB.n134 1.076
R472 VPB.n405 VPB.n402 1.076
R473 VPB.n48 VPB.n45 1.076
R474 VPB.n189 VPB.n188 0.735
R475 VPB.n188 VPB.n178 0.735
R476 VPB.n304 VPB.n301 0.717
R477 VPB.n167 VPB.n166 0.717
R478 VPB.n444 VPB.n441 0.717
R479 VPB.n78 VPB.n77 0.717
R480 VPB.n248 VPB.n247 0.387
R481 VPB.n248 VPB.n243 0.387
R482 VPB.n248 VPB.n238 0.387
R483 VPB.n249 VPB.n248 0.387
R484 VPB.n122 VPB.n121 0.387
R485 VPB.n122 VPB.n117 0.387
R486 VPB.n122 VPB.n112 0.387
R487 VPB.n123 VPB.n122 0.387
R488 VPB.n99 VPB.n98 0.387
R489 VPB.n99 VPB.n94 0.387
R490 VPB.n99 VPB.n89 0.387
R491 VPB.n100 VPB.n99 0.387
R492 VPB.n388 VPB.n387 0.387
R493 VPB.n388 VPB.n383 0.387
R494 VPB.n388 VPB.n378 0.387
R495 VPB.n389 VPB.n388 0.387
R496 VPB.n33 VPB.n32 0.387
R497 VPB.n33 VPB.n28 0.387
R498 VPB.n33 VPB.n23 0.387
R499 VPB.n34 VPB.n33 0.387
R500 VPB.n473 VPB.n13 0.387
R501 VPB.n473 VPB.n9 0.387
R502 VPB.n473 VPB.n4 0.387
R503 VPB.n473 VPB.n472 0.387
R504 VPB.n257 VPB.n230 0.272
R505 VPB.n314 VPB.n313 0.272
R506 VPB.n397 VPB.n370 0.272
R507 VPB.n454 VPB.n453 0.272
R508 VPB.n465 VPB 0.198
R509 VPB.n211 VPB.n210 0.136
R510 VPB.n216 VPB.n211 0.136
R511 VPB.n221 VPB.n216 0.136
R512 VPB.n226 VPB.n221 0.136
R513 VPB.n230 VPB.n226 0.136
R514 VPB.n261 VPB.n257 0.136
R515 VPB.n266 VPB.n261 0.136
R516 VPB.n271 VPB.n266 0.136
R517 VPB.n278 VPB.n271 0.136
R518 VPB.n283 VPB.n278 0.136
R519 VPB.n288 VPB.n283 0.136
R520 VPB.n295 VPB.n288 0.136
R521 VPB.n300 VPB.n295 0.136
R522 VPB.n305 VPB.n300 0.136
R523 VPB.n309 VPB.n305 0.136
R524 VPB.n313 VPB.n309 0.136
R525 VPB.n315 VPB.n314 0.136
R526 VPB.n316 VPB.n315 0.136
R527 VPB.n317 VPB.n316 0.136
R528 VPB.n318 VPB.n317 0.136
R529 VPB.n319 VPB.n318 0.136
R530 VPB.n320 VPB.n319 0.136
R531 VPB.n321 VPB.n320 0.136
R532 VPB.n322 VPB.n321 0.136
R533 VPB.n323 VPB.n322 0.136
R534 VPB.n324 VPB.n323 0.136
R535 VPB.n325 VPB.n324 0.136
R536 VPB.n325 VPB 0.136
R537 VPB.n334 VPB 0.136
R538 VPB.n339 VPB.n334 0.136
R539 VPB.n344 VPB.n339 0.136
R540 VPB.n351 VPB.n344 0.136
R541 VPB.n356 VPB.n351 0.136
R542 VPB.n361 VPB.n356 0.136
R543 VPB.n366 VPB.n361 0.136
R544 VPB.n370 VPB.n366 0.136
R545 VPB.n401 VPB.n397 0.136
R546 VPB.n406 VPB.n401 0.136
R547 VPB.n411 VPB.n406 0.136
R548 VPB.n418 VPB.n411 0.136
R549 VPB.n423 VPB.n418 0.136
R550 VPB.n428 VPB.n423 0.136
R551 VPB.n435 VPB.n428 0.136
R552 VPB.n440 VPB.n435 0.136
R553 VPB.n445 VPB.n440 0.136
R554 VPB.n449 VPB.n445 0.136
R555 VPB.n453 VPB.n449 0.136
R556 VPB.n455 VPB.n454 0.136
R557 VPB.n456 VPB.n455 0.136
R558 VPB.n457 VPB.n456 0.136
R559 VPB.n458 VPB.n457 0.136
R560 VPB.n459 VPB.n458 0.136
R561 VPB.n460 VPB.n459 0.136
R562 VPB.n461 VPB.n460 0.136
R563 VPB.n462 VPB.n461 0.136
R564 VPB.n463 VPB.n462 0.136
R565 VPB.n464 VPB.n463 0.136
R566 VPB.n465 VPB.n464 0.136
R567 a_599_943.n6 a_599_943.t7 480.392
R568 a_599_943.n8 a_599_943.t11 454.685
R569 a_599_943.n8 a_599_943.t9 428.979
R570 a_599_943.n6 a_599_943.t10 403.272
R571 a_599_943.n7 a_599_943.t8 266.974
R572 a_599_943.n9 a_599_943.t12 221.453
R573 a_599_943.n13 a_599_943.n11 196.598
R574 a_599_943.n11 a_599_943.n5 180.846
R575 a_599_943.n9 a_599_943.n8 108.494
R576 a_599_943.n7 a_599_943.n6 108.494
R577 a_599_943.n10 a_599_943.n9 80.035
R578 a_599_943.n4 a_599_943.n3 79.232
R579 a_599_943.n10 a_599_943.n7 77.315
R580 a_599_943.n11 a_599_943.n10 76
R581 a_599_943.n5 a_599_943.n4 63.152
R582 a_599_943.n13 a_599_943.n12 30
R583 a_599_943.n14 a_599_943.n0 24.383
R584 a_599_943.n14 a_599_943.n13 23.684
R585 a_599_943.n5 a_599_943.n1 16.08
R586 a_599_943.n4 a_599_943.n2 16.08
R587 a_599_943.n1 a_599_943.t0 14.282
R588 a_599_943.n1 a_599_943.t1 14.282
R589 a_599_943.n2 a_599_943.t3 14.282
R590 a_599_943.n2 a_599_943.t4 14.282
R591 a_599_943.n3 a_599_943.t6 14.282
R592 a_599_943.n3 a_599_943.t5 14.282
R593 a_91_75.t0 a_91_75.n0 117.777
R594 a_91_75.n2 a_91_75.n1 55.228
R595 a_91_75.n4 a_91_75.n3 9.111
R596 a_91_75.n8 a_91_75.n6 7.859
R597 a_91_75.t0 a_91_75.n2 4.04
R598 a_91_75.t0 a_91_75.n8 3.034
R599 a_91_75.n6 a_91_75.n4 1.964
R600 a_91_75.n6 a_91_75.n5 1.964
R601 a_91_75.n8 a_91_75.n7 0.443
R602 a_372_182.n10 a_372_182.n8 82.852
R603 a_372_182.n11 a_372_182.n0 49.6
R604 a_372_182.n7 a_372_182.n6 32.833
R605 a_372_182.n8 a_372_182.t1 32.416
R606 a_372_182.n10 a_372_182.n9 27.2
R607 a_372_182.n3 a_372_182.n2 23.284
R608 a_372_182.n11 a_372_182.n10 22.4
R609 a_372_182.n7 a_372_182.n4 19.017
R610 a_372_182.n6 a_372_182.n5 13.494
R611 a_372_182.t1 a_372_182.n1 7.04
R612 a_372_182.t1 a_372_182.n3 5.727
R613 a_372_182.n8 a_372_182.n7 1.435
R614 a_3643_75.t0 a_3643_75.n0 117.777
R615 a_3643_75.n2 a_3643_75.n1 55.228
R616 a_3643_75.n4 a_3643_75.n3 9.111
R617 a_3643_75.n8 a_3643_75.n6 7.859
R618 a_3643_75.t0 a_3643_75.n2 4.04
R619 a_3643_75.t0 a_3643_75.n8 3.034
R620 a_3643_75.n6 a_3643_75.n4 1.964
R621 a_3643_75.n6 a_3643_75.n5 1.964
R622 a_3643_75.n8 a_3643_75.n7 0.443
R623 VNB VNB.n407 300.778
R624 VNB.n191 VNB.n190 199.897
R625 VNB.n84 VNB.n83 199.897
R626 VNB.n67 VNB.n66 199.897
R627 VNB.n317 VNB.n316 199.897
R628 VNB.n15 VNB.n14 199.897
R629 VNB.n93 VNB.n91 154.509
R630 VNB.n200 VNB.n198 154.509
R631 VNB.n326 VNB.n324 154.509
R632 VNB.n267 VNB.n265 154.509
R633 VNB.n24 VNB.n22 154.509
R634 VNB.n358 VNB.n357 147.75
R635 VNB.n157 VNB.n156 121.366
R636 VNB.n283 VNB.n282 121.366
R637 VNB.n370 VNB.n367 121.366
R638 VNB.n236 VNB.n235 85.559
R639 VNB.n122 VNB.n73 85.559
R640 VNB.n53 VNB.n4 85.559
R641 VNB.n394 VNB.n393 76
R642 VNB.n381 VNB.n380 76
R643 VNB.n377 VNB.n376 76
R644 VNB.n373 VNB.n372 76
R645 VNB.n361 VNB.n360 76
R646 VNB.n356 VNB.n355 76
R647 VNB.n352 VNB.n351 76
R648 VNB.n348 VNB.n347 76
R649 VNB.n344 VNB.n343 76
R650 VNB.n340 VNB.n339 76
R651 VNB.n336 VNB.n335 76
R652 VNB.n332 VNB.n331 76
R653 VNB.n328 VNB.n327 76
R654 VNB.n306 VNB.n305 76
R655 VNB.n302 VNB.n301 76
R656 VNB.n298 VNB.n297 76
R657 VNB.n287 VNB.n286 76
R658 VNB.n281 VNB.n280 76
R659 VNB.n277 VNB.n276 76
R660 VNB.n273 VNB.n272 76
R661 VNB.n269 VNB.n268 76
R662 VNB.n263 VNB.n260 76
R663 VNB.n248 VNB.n247 76
R664 VNB.n244 VNB.n243 76
R665 VNB.n240 VNB.n239 76
R666 VNB.n234 VNB.n233 76
R667 VNB.n230 VNB.n229 76
R668 VNB.n226 VNB.n225 76
R669 VNB.n222 VNB.n221 76
R670 VNB.n218 VNB.n217 76
R671 VNB.n214 VNB.n213 76
R672 VNB.n210 VNB.n209 76
R673 VNB.n206 VNB.n205 76
R674 VNB.n202 VNB.n201 76
R675 VNB.n180 VNB.n179 76
R676 VNB.n176 VNB.n175 76
R677 VNB.n172 VNB.n171 76
R678 VNB.n161 VNB.n160 76
R679 VNB.n366 VNB.n365 64.552
R680 VNB.n166 VNB.n165 63.835
R681 VNB.n292 VNB.n291 63.835
R682 VNB.n238 VNB.n237 41.971
R683 VNB.n120 VNB.n119 41.971
R684 VNB.n51 VNB.n50 41.971
R685 VNB.n158 VNB.n157 36.937
R686 VNB.n284 VNB.n283 36.937
R687 VNB.n370 VNB.n369 36.937
R688 VNB.n154 VNB.n153 35.118
R689 VNB.n369 VNB.n368 29.844
R690 VNB.n165 VNB.n164 28.421
R691 VNB.n291 VNB.n290 28.421
R692 VNB.n365 VNB.n364 28.421
R693 VNB.n169 VNB.n168 27.855
R694 VNB.n295 VNB.n294 27.855
R695 VNB.n165 VNB.n163 25.263
R696 VNB.n291 VNB.n289 25.263
R697 VNB.n365 VNB.n363 25.263
R698 VNB.n163 VNB.n162 24.383
R699 VNB.n289 VNB.n288 24.383
R700 VNB.n363 VNB.n362 24.383
R701 VNB.n143 VNB.n140 20.452
R702 VNB.n395 VNB.n394 20.452
R703 VNB.n170 VNB.n169 16.721
R704 VNB.n296 VNB.n295 16.721
R705 VNB.n152 VNB.n151 13.653
R706 VNB.n151 VNB.n150 13.653
R707 VNB.n149 VNB.n148 13.653
R708 VNB.n148 VNB.n147 13.653
R709 VNB.n146 VNB.n145 13.653
R710 VNB.n145 VNB.n144 13.653
R711 VNB.n160 VNB.n159 13.653
R712 VNB.n159 VNB.n158 13.653
R713 VNB.n171 VNB.n170 13.653
R714 VNB.n175 VNB.n174 13.653
R715 VNB.n174 VNB.n173 13.653
R716 VNB.n179 VNB.n178 13.653
R717 VNB.n178 VNB.n177 13.653
R718 VNB.n201 VNB.n200 13.653
R719 VNB.n200 VNB.n199 13.653
R720 VNB.n205 VNB.n204 13.653
R721 VNB.n204 VNB.n203 13.653
R722 VNB.n209 VNB.n208 13.653
R723 VNB.n208 VNB.n207 13.653
R724 VNB.n213 VNB.n212 13.653
R725 VNB.n212 VNB.n211 13.653
R726 VNB.n217 VNB.n216 13.653
R727 VNB.n216 VNB.n215 13.653
R728 VNB.n221 VNB.n220 13.653
R729 VNB.n220 VNB.n219 13.653
R730 VNB.n225 VNB.n224 13.653
R731 VNB.n224 VNB.n223 13.653
R732 VNB.n229 VNB.n228 13.653
R733 VNB.n228 VNB.n227 13.653
R734 VNB.n233 VNB.n232 13.653
R735 VNB.n232 VNB.n231 13.653
R736 VNB.n239 VNB.n238 13.653
R737 VNB.n243 VNB.n242 13.653
R738 VNB.n242 VNB.n241 13.653
R739 VNB.n247 VNB.n246 13.653
R740 VNB.n246 VNB.n245 13.653
R741 VNB.n94 VNB.n93 13.653
R742 VNB.n93 VNB.n92 13.653
R743 VNB.n97 VNB.n96 13.653
R744 VNB.n96 VNB.n95 13.653
R745 VNB.n100 VNB.n99 13.653
R746 VNB.n99 VNB.n98 13.653
R747 VNB.n103 VNB.n102 13.653
R748 VNB.n102 VNB.n101 13.653
R749 VNB.n106 VNB.n105 13.653
R750 VNB.n105 VNB.n104 13.653
R751 VNB.n109 VNB.n108 13.653
R752 VNB.n108 VNB.n107 13.653
R753 VNB.n112 VNB.n111 13.653
R754 VNB.n111 VNB.n110 13.653
R755 VNB.n115 VNB.n114 13.653
R756 VNB.n114 VNB.n113 13.653
R757 VNB.n118 VNB.n117 13.653
R758 VNB.n117 VNB.n116 13.653
R759 VNB.n121 VNB.n120 13.653
R760 VNB.n125 VNB.n124 13.653
R761 VNB.n124 VNB.n123 13.653
R762 VNB.n263 VNB.n262 13.653
R763 VNB.n262 VNB.n261 13.653
R764 VNB.n268 VNB.n267 13.653
R765 VNB.n267 VNB.n266 13.653
R766 VNB.n272 VNB.n271 13.653
R767 VNB.n271 VNB.n270 13.653
R768 VNB.n276 VNB.n275 13.653
R769 VNB.n275 VNB.n274 13.653
R770 VNB.n280 VNB.n279 13.653
R771 VNB.n279 VNB.n278 13.653
R772 VNB.n286 VNB.n285 13.653
R773 VNB.n285 VNB.n284 13.653
R774 VNB.n297 VNB.n296 13.653
R775 VNB.n301 VNB.n300 13.653
R776 VNB.n300 VNB.n299 13.653
R777 VNB.n305 VNB.n304 13.653
R778 VNB.n304 VNB.n303 13.653
R779 VNB.n327 VNB.n326 13.653
R780 VNB.n326 VNB.n325 13.653
R781 VNB.n331 VNB.n330 13.653
R782 VNB.n330 VNB.n329 13.653
R783 VNB.n335 VNB.n334 13.653
R784 VNB.n334 VNB.n333 13.653
R785 VNB.n339 VNB.n338 13.653
R786 VNB.n338 VNB.n337 13.653
R787 VNB.n343 VNB.n342 13.653
R788 VNB.n342 VNB.n341 13.653
R789 VNB.n347 VNB.n346 13.653
R790 VNB.n346 VNB.n345 13.653
R791 VNB.n351 VNB.n350 13.653
R792 VNB.n350 VNB.n349 13.653
R793 VNB.n355 VNB.n354 13.653
R794 VNB.n354 VNB.n353 13.653
R795 VNB.n360 VNB.n359 13.653
R796 VNB.n359 VNB.n358 13.653
R797 VNB.n372 VNB.n371 13.653
R798 VNB.n371 VNB.n370 13.653
R799 VNB.n376 VNB.n375 13.653
R800 VNB.n375 VNB.n374 13.653
R801 VNB.n380 VNB.n379 13.653
R802 VNB.n379 VNB.n378 13.653
R803 VNB.n25 VNB.n24 13.653
R804 VNB.n24 VNB.n23 13.653
R805 VNB.n28 VNB.n27 13.653
R806 VNB.n27 VNB.n26 13.653
R807 VNB.n31 VNB.n30 13.653
R808 VNB.n30 VNB.n29 13.653
R809 VNB.n34 VNB.n33 13.653
R810 VNB.n33 VNB.n32 13.653
R811 VNB.n37 VNB.n36 13.653
R812 VNB.n36 VNB.n35 13.653
R813 VNB.n40 VNB.n39 13.653
R814 VNB.n39 VNB.n38 13.653
R815 VNB.n43 VNB.n42 13.653
R816 VNB.n42 VNB.n41 13.653
R817 VNB.n46 VNB.n45 13.653
R818 VNB.n45 VNB.n44 13.653
R819 VNB.n49 VNB.n48 13.653
R820 VNB.n48 VNB.n47 13.653
R821 VNB.n52 VNB.n51 13.653
R822 VNB.n56 VNB.n55 13.653
R823 VNB.n55 VNB.n54 13.653
R824 VNB.n394 VNB.n0 13.653
R825 VNB VNB.n0 13.653
R826 VNB.n143 VNB.n142 13.653
R827 VNB.n142 VNB.n141 13.653
R828 VNB.n402 VNB.n399 13.577
R829 VNB.n128 VNB.n126 13.276
R830 VNB.n140 VNB.n128 13.276
R831 VNB.n183 VNB.n181 13.276
R832 VNB.n196 VNB.n183 13.276
R833 VNB.n76 VNB.n74 13.276
R834 VNB.n89 VNB.n76 13.276
R835 VNB.n59 VNB.n57 13.276
R836 VNB.n72 VNB.n59 13.276
R837 VNB.n309 VNB.n307 13.276
R838 VNB.n322 VNB.n309 13.276
R839 VNB.n7 VNB.n5 13.276
R840 VNB.n20 VNB.n7 13.276
R841 VNB.n152 VNB.n149 13.276
R842 VNB.n149 VNB.n146 13.276
R843 VNB.n201 VNB.n197 13.276
R844 VNB.n94 VNB.n90 13.276
R845 VNB.n97 VNB.n94 13.276
R846 VNB.n100 VNB.n97 13.276
R847 VNB.n103 VNB.n100 13.276
R848 VNB.n106 VNB.n103 13.276
R849 VNB.n109 VNB.n106 13.276
R850 VNB.n112 VNB.n109 13.276
R851 VNB.n115 VNB.n112 13.276
R852 VNB.n118 VNB.n115 13.276
R853 VNB.n121 VNB.n118 13.276
R854 VNB.n263 VNB.n125 13.276
R855 VNB.n264 VNB.n263 13.276
R856 VNB.n268 VNB.n264 13.276
R857 VNB.n327 VNB.n323 13.276
R858 VNB.n25 VNB.n21 13.276
R859 VNB.n28 VNB.n25 13.276
R860 VNB.n31 VNB.n28 13.276
R861 VNB.n34 VNB.n31 13.276
R862 VNB.n37 VNB.n34 13.276
R863 VNB.n40 VNB.n37 13.276
R864 VNB.n43 VNB.n40 13.276
R865 VNB.n46 VNB.n43 13.276
R866 VNB.n49 VNB.n46 13.276
R867 VNB.n52 VNB.n49 13.276
R868 VNB.n394 VNB.n56 13.276
R869 VNB.n3 VNB.n1 13.276
R870 VNB.n395 VNB.n3 13.276
R871 VNB.n125 VNB.n122 12.02
R872 VNB.n56 VNB.n53 12.02
R873 VNB.n404 VNB.n403 7.5
R874 VNB.n189 VNB.n188 7.5
R875 VNB.n185 VNB.n184 7.5
R876 VNB.n183 VNB.n182 7.5
R877 VNB.n196 VNB.n195 7.5
R878 VNB.n82 VNB.n81 7.5
R879 VNB.n78 VNB.n77 7.5
R880 VNB.n76 VNB.n75 7.5
R881 VNB.n89 VNB.n88 7.5
R882 VNB.n65 VNB.n64 7.5
R883 VNB.n61 VNB.n60 7.5
R884 VNB.n59 VNB.n58 7.5
R885 VNB.n72 VNB.n71 7.5
R886 VNB.n315 VNB.n314 7.5
R887 VNB.n311 VNB.n310 7.5
R888 VNB.n309 VNB.n308 7.5
R889 VNB.n322 VNB.n321 7.5
R890 VNB.n13 VNB.n12 7.5
R891 VNB.n9 VNB.n8 7.5
R892 VNB.n7 VNB.n6 7.5
R893 VNB.n20 VNB.n19 7.5
R894 VNB.n396 VNB.n395 7.5
R895 VNB.n3 VNB.n2 7.5
R896 VNB.n401 VNB.n400 7.5
R897 VNB.n134 VNB.n133 7.5
R898 VNB.n130 VNB.n129 7.5
R899 VNB.n128 VNB.n127 7.5
R900 VNB.n140 VNB.n139 7.5
R901 VNB.n197 VNB.n196 7.176
R902 VNB.n90 VNB.n89 7.176
R903 VNB.n264 VNB.n72 7.176
R904 VNB.n323 VNB.n322 7.176
R905 VNB.n21 VNB.n20 7.176
R906 VNB.n406 VNB.n404 7.011
R907 VNB.n192 VNB.n189 7.011
R908 VNB.n187 VNB.n185 7.011
R909 VNB.n85 VNB.n82 7.011
R910 VNB.n80 VNB.n78 7.011
R911 VNB.n68 VNB.n65 7.011
R912 VNB.n63 VNB.n61 7.011
R913 VNB.n318 VNB.n315 7.011
R914 VNB.n313 VNB.n311 7.011
R915 VNB.n16 VNB.n13 7.011
R916 VNB.n11 VNB.n9 7.011
R917 VNB.n136 VNB.n134 7.011
R918 VNB.n132 VNB.n130 7.011
R919 VNB.n195 VNB.n194 7.01
R920 VNB.n187 VNB.n186 7.01
R921 VNB.n192 VNB.n191 7.01
R922 VNB.n88 VNB.n87 7.01
R923 VNB.n80 VNB.n79 7.01
R924 VNB.n85 VNB.n84 7.01
R925 VNB.n71 VNB.n70 7.01
R926 VNB.n63 VNB.n62 7.01
R927 VNB.n68 VNB.n67 7.01
R928 VNB.n321 VNB.n320 7.01
R929 VNB.n313 VNB.n312 7.01
R930 VNB.n318 VNB.n317 7.01
R931 VNB.n19 VNB.n18 7.01
R932 VNB.n11 VNB.n10 7.01
R933 VNB.n16 VNB.n15 7.01
R934 VNB.n139 VNB.n138 7.01
R935 VNB.n132 VNB.n131 7.01
R936 VNB.n136 VNB.n135 7.01
R937 VNB.n406 VNB.n405 7.01
R938 VNB.n402 VNB.n401 6.788
R939 VNB.n397 VNB.n396 6.788
R940 VNB.n153 VNB.n143 6.111
R941 VNB.n153 VNB.n152 6.1
R942 VNB.n171 VNB.n166 2.511
R943 VNB.n297 VNB.n292 2.511
R944 VNB.n169 VNB.n167 1.99
R945 VNB.n295 VNB.n293 1.99
R946 VNB.n239 VNB.n236 1.255
R947 VNB.n122 VNB.n121 1.255
R948 VNB.n372 VNB.n366 1.255
R949 VNB.n53 VNB.n52 1.255
R950 VNB.n407 VNB.n398 0.921
R951 VNB.n407 VNB.n402 0.476
R952 VNB.n407 VNB.n397 0.475
R953 VNB.n202 VNB.n180 0.272
R954 VNB.n249 VNB.n248 0.272
R955 VNB.n328 VNB.n306 0.272
R956 VNB.n382 VNB.n381 0.272
R957 VNB.n193 VNB.n187 0.246
R958 VNB.n194 VNB.n193 0.246
R959 VNB.n193 VNB.n192 0.246
R960 VNB.n86 VNB.n80 0.246
R961 VNB.n87 VNB.n86 0.246
R962 VNB.n86 VNB.n85 0.246
R963 VNB.n69 VNB.n63 0.246
R964 VNB.n70 VNB.n69 0.246
R965 VNB.n69 VNB.n68 0.246
R966 VNB.n319 VNB.n313 0.246
R967 VNB.n320 VNB.n319 0.246
R968 VNB.n319 VNB.n318 0.246
R969 VNB.n17 VNB.n11 0.246
R970 VNB.n18 VNB.n17 0.246
R971 VNB.n17 VNB.n16 0.246
R972 VNB.n137 VNB.n132 0.246
R973 VNB.n138 VNB.n137 0.246
R974 VNB.n137 VNB.n136 0.246
R975 VNB.n407 VNB.n406 0.246
R976 VNB.n393 VNB 0.198
R977 VNB.n155 VNB.n154 0.136
R978 VNB.n161 VNB.n155 0.136
R979 VNB.n172 VNB.n161 0.136
R980 VNB.n176 VNB.n172 0.136
R981 VNB.n180 VNB.n176 0.136
R982 VNB.n206 VNB.n202 0.136
R983 VNB.n210 VNB.n206 0.136
R984 VNB.n214 VNB.n210 0.136
R985 VNB.n218 VNB.n214 0.136
R986 VNB.n222 VNB.n218 0.136
R987 VNB.n226 VNB.n222 0.136
R988 VNB.n230 VNB.n226 0.136
R989 VNB.n234 VNB.n230 0.136
R990 VNB.n240 VNB.n234 0.136
R991 VNB.n244 VNB.n240 0.136
R992 VNB.n248 VNB.n244 0.136
R993 VNB.n250 VNB.n249 0.136
R994 VNB.n251 VNB.n250 0.136
R995 VNB.n252 VNB.n251 0.136
R996 VNB.n253 VNB.n252 0.136
R997 VNB.n254 VNB.n253 0.136
R998 VNB.n255 VNB.n254 0.136
R999 VNB.n256 VNB.n255 0.136
R1000 VNB.n257 VNB.n256 0.136
R1001 VNB.n258 VNB.n257 0.136
R1002 VNB.n259 VNB.n258 0.136
R1003 VNB.n260 VNB.n259 0.136
R1004 VNB.n260 VNB 0.136
R1005 VNB.n269 VNB 0.136
R1006 VNB.n273 VNB.n269 0.136
R1007 VNB.n277 VNB.n273 0.136
R1008 VNB.n281 VNB.n277 0.136
R1009 VNB.n287 VNB.n281 0.136
R1010 VNB.n298 VNB.n287 0.136
R1011 VNB.n302 VNB.n298 0.136
R1012 VNB.n306 VNB.n302 0.136
R1013 VNB.n332 VNB.n328 0.136
R1014 VNB.n336 VNB.n332 0.136
R1015 VNB.n340 VNB.n336 0.136
R1016 VNB.n344 VNB.n340 0.136
R1017 VNB.n348 VNB.n344 0.136
R1018 VNB.n352 VNB.n348 0.136
R1019 VNB.n356 VNB.n352 0.136
R1020 VNB.n361 VNB.n356 0.136
R1021 VNB.n373 VNB.n361 0.136
R1022 VNB.n377 VNB.n373 0.136
R1023 VNB.n381 VNB.n377 0.136
R1024 VNB.n383 VNB.n382 0.136
R1025 VNB.n384 VNB.n383 0.136
R1026 VNB.n385 VNB.n384 0.136
R1027 VNB.n386 VNB.n385 0.136
R1028 VNB.n387 VNB.n386 0.136
R1029 VNB.n388 VNB.n387 0.136
R1030 VNB.n389 VNB.n388 0.136
R1031 VNB.n390 VNB.n389 0.136
R1032 VNB.n391 VNB.n390 0.136
R1033 VNB.n392 VNB.n391 0.136
R1034 VNB.n393 VNB.n392 0.136
R1035 a_2141_1004.n4 a_2141_1004.t6 512.525
R1036 a_2141_1004.n4 a_2141_1004.t7 371.139
R1037 a_2141_1004.n5 a_2141_1004.t5 271.162
R1038 a_2141_1004.n8 a_2141_1004.n6 194.086
R1039 a_2141_1004.n5 a_2141_1004.n4 172.76
R1040 a_2141_1004.n6 a_2141_1004.n3 162.547
R1041 a_2141_1004.n6 a_2141_1004.n5 153.315
R1042 a_2141_1004.n3 a_2141_1004.n2 76.002
R1043 a_2141_1004.n8 a_2141_1004.n7 30
R1044 a_2141_1004.n9 a_2141_1004.n0 24.383
R1045 a_2141_1004.n9 a_2141_1004.n8 23.684
R1046 a_2141_1004.n1 a_2141_1004.t3 14.282
R1047 a_2141_1004.n1 a_2141_1004.t2 14.282
R1048 a_2141_1004.n2 a_2141_1004.t1 14.282
R1049 a_2141_1004.n2 a_2141_1004.t0 14.282
R1050 a_2141_1004.n3 a_2141_1004.n1 12.85
R1051 a_4626_73.n5 a_4626_73.n4 24.877
R1052 a_4626_73.t0 a_4626_73.n5 12.677
R1053 a_4626_73.t0 a_4626_73.n3 11.595
R1054 a_4626_73.t0 a_4626_73.n6 8.137
R1055 a_4626_73.n2 a_4626_73.n0 4.031
R1056 a_4626_73.n2 a_4626_73.n1 3.644
R1057 a_4626_73.t0 a_4626_73.n2 1.093
R1058 a_4151_943.n3 a_4151_943.t5 454.685
R1059 a_4151_943.n3 a_4151_943.t6 428.979
R1060 a_4151_943.n4 a_4151_943.t7 248.006
R1061 a_4151_943.n7 a_4151_943.n5 227.161
R1062 a_4151_943.n5 a_4151_943.n4 154.947
R1063 a_4151_943.n5 a_4151_943.n2 135.994
R1064 a_4151_943.n4 a_4151_943.n3 81.941
R1065 a_4151_943.n2 a_4151_943.n1 76.002
R1066 a_4151_943.n7 a_4151_943.n6 15.218
R1067 a_4151_943.n0 a_4151_943.t2 14.282
R1068 a_4151_943.n0 a_4151_943.t3 14.282
R1069 a_4151_943.n1 a_4151_943.t0 14.282
R1070 a_4151_943.n1 a_4151_943.t1 14.282
R1071 a_4151_943.n2 a_4151_943.n0 12.85
R1072 a_4151_943.n8 a_4151_943.n7 12.014
R1073 a_1334_182.n9 a_1334_182.n7 82.852
R1074 a_1334_182.n3 a_1334_182.n1 44.628
R1075 a_1334_182.t0 a_1334_182.n9 32.417
R1076 a_1334_182.n7 a_1334_182.n6 27.2
R1077 a_1334_182.n5 a_1334_182.n4 23.498
R1078 a_1334_182.n3 a_1334_182.n2 23.284
R1079 a_1334_182.n7 a_1334_182.n5 22.4
R1080 a_1334_182.t0 a_1334_182.n11 20.241
R1081 a_1334_182.n11 a_1334_182.n10 13.494
R1082 a_1334_182.t0 a_1334_182.n0 8.137
R1083 a_1334_182.t0 a_1334_182.n3 5.727
R1084 a_1334_182.n9 a_1334_182.n8 1.435
R1085 a_2036_73.n12 a_2036_73.n11 26.811
R1086 a_2036_73.n6 a_2036_73.n5 24.977
R1087 a_2036_73.n2 a_2036_73.n1 24.877
R1088 a_2036_73.t0 a_2036_73.n2 12.677
R1089 a_2036_73.t0 a_2036_73.n3 11.595
R1090 a_2036_73.t1 a_2036_73.n8 8.137
R1091 a_2036_73.t0 a_2036_73.n4 7.273
R1092 a_2036_73.t0 a_2036_73.n0 6.109
R1093 a_2036_73.t1 a_2036_73.n7 4.864
R1094 a_2036_73.t0 a_2036_73.n12 2.074
R1095 a_2036_73.n7 a_2036_73.n6 1.13
R1096 a_2036_73.n12 a_2036_73.t1 0.937
R1097 a_2036_73.t1 a_2036_73.n10 0.804
R1098 a_2036_73.n10 a_2036_73.n9 0.136
R1099 a_2681_75.n1 a_2681_75.n0 25.576
R1100 a_2681_75.n3 a_2681_75.n2 9.111
R1101 a_2681_75.n7 a_2681_75.n5 7.859
R1102 a_2681_75.t0 a_2681_75.n7 3.034
R1103 a_2681_75.n5 a_2681_75.n3 1.964
R1104 a_2681_75.n5 a_2681_75.n4 1.964
R1105 a_2681_75.t0 a_2681_75.n1 1.871
R1106 a_2681_75.n7 a_2681_75.n6 0.443
R1107 a_3924_182.n10 a_3924_182.n8 82.852
R1108 a_3924_182.n11 a_3924_182.n0 49.6
R1109 a_3924_182.n7 a_3924_182.n6 32.833
R1110 a_3924_182.n8 a_3924_182.t1 32.416
R1111 a_3924_182.n10 a_3924_182.n9 27.2
R1112 a_3924_182.n3 a_3924_182.n2 23.284
R1113 a_3924_182.n11 a_3924_182.n10 22.4
R1114 a_3924_182.n7 a_3924_182.n4 19.017
R1115 a_3924_182.n6 a_3924_182.n5 13.494
R1116 a_3924_182.t1 a_3924_182.n1 7.04
R1117 a_3924_182.t1 a_3924_182.n3 5.727
R1118 a_3924_182.n8 a_3924_182.n7 1.435
R1119 a_1053_75.n1 a_1053_75.n0 25.576
R1120 a_1053_75.n3 a_1053_75.n2 9.111
R1121 a_1053_75.n7 a_1053_75.n6 2.455
R1122 a_1053_75.n5 a_1053_75.n3 1.964
R1123 a_1053_75.n5 a_1053_75.n4 1.964
R1124 a_1053_75.t0 a_1053_75.n1 1.871
R1125 a_1053_75.n7 a_1053_75.n5 0.636
R1126 a_1053_75.t0 a_1053_75.n7 0.246
R1127 a_2962_182.n8 a_2962_182.n6 96.467
R1128 a_2962_182.n3 a_2962_182.n1 44.628
R1129 a_2962_182.t0 a_2962_182.n8 32.417
R1130 a_2962_182.n3 a_2962_182.n2 23.284
R1131 a_2962_182.n6 a_2962_182.n5 22.349
R1132 a_2962_182.t0 a_2962_182.n10 20.241
R1133 a_2962_182.n10 a_2962_182.n9 13.494
R1134 a_2962_182.n6 a_2962_182.n4 8.443
R1135 a_2962_182.t0 a_2962_182.n0 8.137
R1136 a_2962_182.t0 a_2962_182.n3 5.727
R1137 a_2962_182.n8 a_2962_182.n7 1.435
C8 VPB VNB 20.02fF
C9 a_2962_182.n0 VNB 0.07fF
C10 a_2962_182.n1 VNB 0.09fF
C11 a_2962_182.n2 VNB 0.13fF
C12 a_2962_182.n3 VNB 0.11fF
C13 a_2962_182.n4 VNB 0.02fF
C14 a_2962_182.n5 VNB 0.03fF
C15 a_2962_182.n6 VNB 0.06fF
C16 a_2962_182.n7 VNB 0.03fF
C17 a_2962_182.n8 VNB 0.12fF
C18 a_2962_182.n9 VNB 0.06fF
C19 a_2962_182.n10 VNB 0.01fF
C20 a_2962_182.t0 VNB 0.33fF
C21 a_1053_75.n0 VNB 0.09fF
C22 a_1053_75.n1 VNB 0.10fF
C23 a_1053_75.n2 VNB 0.05fF
C24 a_1053_75.n3 VNB 0.03fF
C25 a_1053_75.n4 VNB 0.04fF
C26 a_1053_75.n5 VNB 0.03fF
C27 a_1053_75.n6 VNB 0.04fF
C28 a_3924_182.n0 VNB 0.02fF
C29 a_3924_182.n1 VNB 0.09fF
C30 a_3924_182.n2 VNB 0.13fF
C31 a_3924_182.n3 VNB 0.11fF
C32 a_3924_182.n4 VNB 0.09fF
C33 a_3924_182.n5 VNB 0.06fF
C34 a_3924_182.n6 VNB 0.01fF
C35 a_3924_182.n7 VNB 0.03fF
C36 a_3924_182.n8 VNB 0.11fF
C37 a_3924_182.n9 VNB 0.02fF
C38 a_3924_182.n10 VNB 0.05fF
C39 a_3924_182.n11 VNB 0.02fF
C40 a_2681_75.n0 VNB 0.09fF
C41 a_2681_75.n1 VNB 0.10fF
C42 a_2681_75.n2 VNB 0.05fF
C43 a_2681_75.n3 VNB 0.03fF
C44 a_2681_75.n4 VNB 0.04fF
C45 a_2681_75.n5 VNB 0.11fF
C46 a_2681_75.n6 VNB 0.04fF
C47 a_2036_73.n0 VNB 0.02fF
C48 a_2036_73.n1 VNB 0.10fF
C49 a_2036_73.n2 VNB 0.06fF
C50 a_2036_73.n3 VNB 0.06fF
C51 a_2036_73.n4 VNB 0.00fF
C52 a_2036_73.n5 VNB 0.04fF
C53 a_2036_73.n6 VNB 0.05fF
C54 a_2036_73.n7 VNB 0.02fF
C55 a_2036_73.n8 VNB 0.05fF
C56 a_2036_73.n9 VNB 0.08fF
C57 a_2036_73.n10 VNB 0.17fF
C58 a_2036_73.t1 VNB 0.23fF
C59 a_2036_73.n11 VNB 0.09fF
C60 a_2036_73.n12 VNB 0.00fF
C61 a_1334_182.n0 VNB 0.07fF
C62 a_1334_182.n1 VNB 0.09fF
C63 a_1334_182.n2 VNB 0.13fF
C64 a_1334_182.n3 VNB 0.11fF
C65 a_1334_182.n4 VNB 0.02fF
C66 a_1334_182.n5 VNB 0.03fF
C67 a_1334_182.n6 VNB 0.02fF
C68 a_1334_182.n7 VNB 0.05fF
C69 a_1334_182.n8 VNB 0.03fF
C70 a_1334_182.n9 VNB 0.11fF
C71 a_1334_182.n10 VNB 0.06fF
C72 a_1334_182.n11 VNB 0.01fF
C73 a_1334_182.t0 VNB 0.33fF
C74 a_4151_943.n0 VNB 0.54fF
C75 a_4151_943.n1 VNB 0.64fF
C76 a_4151_943.n2 VNB 0.29fF
C77 a_4151_943.n3 VNB 0.37fF
C78 a_4151_943.n4 VNB 0.74fF
C79 a_4151_943.n5 VNB 0.81fF
C80 a_4151_943.n6 VNB 0.09fF
C81 a_4151_943.n7 VNB 0.31fF
C82 a_4151_943.n8 VNB 0.05fF
C83 a_4626_73.n0 VNB 0.07fF
C84 a_4626_73.n1 VNB 0.02fF
C85 a_4626_73.n2 VNB 0.01fF
C86 a_4626_73.n3 VNB 0.06fF
C87 a_4626_73.n4 VNB 0.10fF
C88 a_4626_73.n5 VNB 0.06fF
C89 a_4626_73.n6 VNB 0.05fF
C90 a_2141_1004.n0 VNB 0.04fF
C91 a_2141_1004.n1 VNB 0.52fF
C92 a_2141_1004.n2 VNB 0.62fF
C93 a_2141_1004.n3 VNB 0.31fF
C94 a_2141_1004.n4 VNB 0.34fF
C95 a_2141_1004.n5 VNB 0.64fF
C96 a_2141_1004.n6 VNB 0.59fF
C97 a_2141_1004.n7 VNB 0.03fF
C98 a_2141_1004.n8 VNB 0.28fF
C99 a_2141_1004.n9 VNB 0.05fF
C100 a_3643_75.n0 VNB 0.03fF
C101 a_3643_75.n1 VNB 0.10fF
C102 a_3643_75.n2 VNB 0.10fF
C103 a_3643_75.n3 VNB 0.05fF
C104 a_3643_75.n4 VNB 0.03fF
C105 a_3643_75.n5 VNB 0.04fF
C106 a_3643_75.n6 VNB 0.11fF
C107 a_3643_75.n7 VNB 0.04fF
C108 a_372_182.n0 VNB 0.02fF
C109 a_372_182.n1 VNB 0.09fF
C110 a_372_182.n2 VNB 0.13fF
C111 a_372_182.n3 VNB 0.11fF
C112 a_372_182.t1 VNB 0.30fF
C113 a_372_182.n4 VNB 0.09fF
C114 a_372_182.n5 VNB 0.06fF
C115 a_372_182.n6 VNB 0.01fF
C116 a_372_182.n7 VNB 0.03fF
C117 a_372_182.n8 VNB 0.11fF
C118 a_372_182.n9 VNB 0.02fF
C119 a_372_182.n10 VNB 0.05fF
C120 a_372_182.n11 VNB 0.02fF
C121 a_91_75.n0 VNB 0.03fF
C122 a_91_75.n1 VNB 0.10fF
C123 a_91_75.n2 VNB 0.10fF
C124 a_91_75.n3 VNB 0.04fF
C125 a_91_75.n4 VNB 0.03fF
C126 a_91_75.n5 VNB 0.03fF
C127 a_91_75.n6 VNB 0.11fF
C128 a_91_75.n7 VNB 0.04fF
C129 a_599_943.n0 VNB 0.04fF
C130 a_599_943.n1 VNB 0.57fF
C131 a_599_943.n2 VNB 0.57fF
C132 a_599_943.n3 VNB 0.66fF
C133 a_599_943.n4 VNB 0.21fF
C134 a_599_943.n5 VNB 0.34fF
C135 a_599_943.n6 VNB 0.41fF
C136 a_599_943.n7 VNB 0.41fF
C137 a_599_943.n8 VNB 0.41fF
C138 a_599_943.t12 VNB 0.54fF
C139 a_599_943.n9 VNB 0.40fF
C140 a_599_943.n10 VNB 1.31fF
C141 a_599_943.n11 VNB 0.47fF
C142 a_599_943.n12 VNB 0.04fF
C143 a_599_943.n13 VNB 0.30fF
C144 a_599_943.n14 VNB 0.06fF
C145 VPB.n0 VNB 0.03fF
C146 VPB.n1 VNB 0.04fF
C147 VPB.n2 VNB 0.02fF
C148 VPB.n3 VNB 0.18fF
C149 VPB.n5 VNB 0.02fF
C150 VPB.n6 VNB 0.02fF
C151 VPB.n7 VNB 0.02fF
C152 VPB.n8 VNB 0.02fF
C153 VPB.n10 VNB 0.02fF
C154 VPB.n11 VNB 0.02fF
C155 VPB.n12 VNB 0.02fF
C156 VPB.n14 VNB 0.10fF
C157 VPB.n15 VNB 0.10fF
C158 VPB.n16 VNB 0.02fF
C159 VPB.n17 VNB 0.02fF
C160 VPB.n18 VNB 0.02fF
C161 VPB.n19 VNB 0.04fF
C162 VPB.n20 VNB 0.02fF
C163 VPB.n21 VNB 0.29fF
C164 VPB.n22 VNB 0.04fF
C165 VPB.n24 VNB 0.02fF
C166 VPB.n25 VNB 0.02fF
C167 VPB.n26 VNB 0.02fF
C168 VPB.n27 VNB 0.02fF
C169 VPB.n29 VNB 0.02fF
C170 VPB.n30 VNB 0.02fF
C171 VPB.n31 VNB 0.02fF
C172 VPB.n33 VNB 0.27fF
C173 VPB.n35 VNB 0.03fF
C174 VPB.n36 VNB 0.02fF
C175 VPB.n37 VNB 0.03fF
C176 VPB.n38 VNB 0.03fF
C177 VPB.n39 VNB 0.27fF
C178 VPB.n40 VNB 0.01fF
C179 VPB.n41 VNB 0.02fF
C180 VPB.n42 VNB 0.27fF
C181 VPB.n43 VNB 0.02fF
C182 VPB.n44 VNB 0.02fF
C183 VPB.n45 VNB 0.05fF
C184 VPB.n46 VNB 0.20fF
C185 VPB.n47 VNB 0.02fF
C186 VPB.n48 VNB 0.01fF
C187 VPB.n49 VNB 0.14fF
C188 VPB.n50 VNB 0.16fF
C189 VPB.n51 VNB 0.02fF
C190 VPB.n52 VNB 0.02fF
C191 VPB.n53 VNB 0.14fF
C192 VPB.n54 VNB 0.16fF
C193 VPB.n55 VNB 0.02fF
C194 VPB.n56 VNB 0.02fF
C195 VPB.n57 VNB 0.02fF
C196 VPB.n58 VNB 0.14fF
C197 VPB.n59 VNB 0.15fF
C198 VPB.n60 VNB 0.02fF
C199 VPB.n61 VNB 0.02fF
C200 VPB.n62 VNB 0.14fF
C201 VPB.n63 VNB 0.15fF
C202 VPB.n64 VNB 0.02fF
C203 VPB.n65 VNB 0.02fF
C204 VPB.n66 VNB 0.02fF
C205 VPB.n67 VNB 0.14fF
C206 VPB.n68 VNB 0.16fF
C207 VPB.n69 VNB 0.02fF
C208 VPB.n70 VNB 0.02fF
C209 VPB.n71 VNB 0.14fF
C210 VPB.n72 VNB 0.16fF
C211 VPB.n73 VNB 0.02fF
C212 VPB.n74 VNB 0.02fF
C213 VPB.n75 VNB 0.21fF
C214 VPB.n76 VNB 0.02fF
C215 VPB.n77 VNB 0.01fF
C216 VPB.n78 VNB 0.06fF
C217 VPB.n79 VNB 0.27fF
C218 VPB.n80 VNB 0.02fF
C219 VPB.n81 VNB 0.02fF
C220 VPB.n82 VNB 0.02fF
C221 VPB.n83 VNB 0.02fF
C222 VPB.n84 VNB 0.02fF
C223 VPB.n85 VNB 0.04fF
C224 VPB.n86 VNB 0.02fF
C225 VPB.n87 VNB 0.24fF
C226 VPB.n88 VNB 0.04fF
C227 VPB.n90 VNB 0.02fF
C228 VPB.n91 VNB 0.02fF
C229 VPB.n92 VNB 0.02fF
C230 VPB.n93 VNB 0.02fF
C231 VPB.n95 VNB 0.02fF
C232 VPB.n96 VNB 0.02fF
C233 VPB.n97 VNB 0.02fF
C234 VPB.n99 VNB 0.27fF
C235 VPB.n101 VNB 0.03fF
C236 VPB.n102 VNB 0.02fF
C237 VPB.n103 VNB 0.10fF
C238 VPB.n104 VNB 0.10fF
C239 VPB.n105 VNB 0.02fF
C240 VPB.n106 VNB 0.02fF
C241 VPB.n107 VNB 0.02fF
C242 VPB.n108 VNB 0.04fF
C243 VPB.n109 VNB 0.02fF
C244 VPB.n110 VNB 0.28fF
C245 VPB.n111 VNB 0.04fF
C246 VPB.n113 VNB 0.02fF
C247 VPB.n114 VNB 0.02fF
C248 VPB.n115 VNB 0.02fF
C249 VPB.n116 VNB 0.02fF
C250 VPB.n118 VNB 0.02fF
C251 VPB.n119 VNB 0.02fF
C252 VPB.n120 VNB 0.02fF
C253 VPB.n122 VNB 0.27fF
C254 VPB.n124 VNB 0.03fF
C255 VPB.n125 VNB 0.02fF
C256 VPB.n126 VNB 0.03fF
C257 VPB.n127 VNB 0.03fF
C258 VPB.n128 VNB 0.27fF
C259 VPB.n129 VNB 0.01fF
C260 VPB.n130 VNB 0.02fF
C261 VPB.n131 VNB 0.27fF
C262 VPB.n132 VNB 0.02fF
C263 VPB.n133 VNB 0.02fF
C264 VPB.n134 VNB 0.05fF
C265 VPB.n135 VNB 0.20fF
C266 VPB.n136 VNB 0.02fF
C267 VPB.n137 VNB 0.01fF
C268 VPB.n138 VNB 0.14fF
C269 VPB.n139 VNB 0.16fF
C270 VPB.n140 VNB 0.02fF
C271 VPB.n141 VNB 0.02fF
C272 VPB.n142 VNB 0.14fF
C273 VPB.n143 VNB 0.16fF
C274 VPB.n144 VNB 0.02fF
C275 VPB.n145 VNB 0.02fF
C276 VPB.n146 VNB 0.02fF
C277 VPB.n147 VNB 0.14fF
C278 VPB.n148 VNB 0.15fF
C279 VPB.n149 VNB 0.02fF
C280 VPB.n150 VNB 0.02fF
C281 VPB.n151 VNB 0.14fF
C282 VPB.n152 VNB 0.15fF
C283 VPB.n153 VNB 0.02fF
C284 VPB.n154 VNB 0.02fF
C285 VPB.n155 VNB 0.02fF
C286 VPB.n156 VNB 0.14fF
C287 VPB.n157 VNB 0.16fF
C288 VPB.n158 VNB 0.02fF
C289 VPB.n159 VNB 0.02fF
C290 VPB.n160 VNB 0.14fF
C291 VPB.n161 VNB 0.16fF
C292 VPB.n162 VNB 0.02fF
C293 VPB.n163 VNB 0.02fF
C294 VPB.n164 VNB 0.21fF
C295 VPB.n165 VNB 0.02fF
C296 VPB.n166 VNB 0.01fF
C297 VPB.n167 VNB 0.06fF
C298 VPB.n168 VNB 0.27fF
C299 VPB.n169 VNB 0.02fF
C300 VPB.n170 VNB 0.02fF
C301 VPB.n171 VNB 0.02fF
C302 VPB.n172 VNB 0.02fF
C303 VPB.n173 VNB 0.02fF
C304 VPB.n174 VNB 0.14fF
C305 VPB.n175 VNB 0.03fF
C306 VPB.n176 VNB 0.02fF
C307 VPB.n177 VNB 0.05fF
C308 VPB.n178 VNB 0.01fF
C309 VPB.n180 VNB 0.02fF
C310 VPB.n181 VNB 0.02fF
C311 VPB.n182 VNB 0.02fF
C312 VPB.n183 VNB 0.02fF
C313 VPB.n186 VNB 0.02fF
C314 VPB.n188 VNB 0.45fF
C315 VPB.n190 VNB 0.04fF
C316 VPB.n191 VNB 0.04fF
C317 VPB.n192 VNB 0.27fF
C318 VPB.n193 VNB 0.03fF
C319 VPB.n194 VNB 0.03fF
C320 VPB.n195 VNB 0.10fF
C321 VPB.n196 VNB 0.02fF
C322 VPB.n197 VNB 0.14fF
C323 VPB.n198 VNB 0.15fF
C324 VPB.n199 VNB 0.02fF
C325 VPB.n200 VNB 0.02fF
C326 VPB.n201 VNB 0.14fF
C327 VPB.n202 VNB 0.16fF
C328 VPB.n203 VNB 0.02fF
C329 VPB.n204 VNB 0.02fF
C330 VPB.n205 VNB 0.05fF
C331 VPB.n206 VNB 0.23fF
C332 VPB.n207 VNB 0.02fF
C333 VPB.n208 VNB 0.01fF
C334 VPB.n209 VNB 0.00fF
C335 VPB.n210 VNB 0.09fF
C336 VPB.n211 VNB 0.02fF
C337 VPB.n212 VNB 0.14fF
C338 VPB.n213 VNB 0.15fF
C339 VPB.n214 VNB 0.02fF
C340 VPB.n215 VNB 0.02fF
C341 VPB.n216 VNB 0.02fF
C342 VPB.n217 VNB 0.14fF
C343 VPB.n218 VNB 0.16fF
C344 VPB.n219 VNB 0.02fF
C345 VPB.n220 VNB 0.02fF
C346 VPB.n221 VNB 0.02fF
C347 VPB.n222 VNB 0.06fF
C348 VPB.n223 VNB 0.23fF
C349 VPB.n224 VNB 0.02fF
C350 VPB.n225 VNB 0.01fF
C351 VPB.n226 VNB 0.02fF
C352 VPB.n227 VNB 0.27fF
C353 VPB.n228 VNB 0.01fF
C354 VPB.n229 VNB 0.02fF
C355 VPB.n230 VNB 0.04fF
C356 VPB.n231 VNB 0.02fF
C357 VPB.n232 VNB 0.02fF
C358 VPB.n233 VNB 0.02fF
C359 VPB.n234 VNB 0.04fF
C360 VPB.n235 VNB 0.02fF
C361 VPB.n236 VNB 0.24fF
C362 VPB.n237 VNB 0.04fF
C363 VPB.n239 VNB 0.02fF
C364 VPB.n240 VNB 0.02fF
C365 VPB.n241 VNB 0.02fF
C366 VPB.n242 VNB 0.02fF
C367 VPB.n244 VNB 0.02fF
C368 VPB.n245 VNB 0.02fF
C369 VPB.n246 VNB 0.02fF
C370 VPB.n248 VNB 0.27fF
C371 VPB.n250 VNB 0.03fF
C372 VPB.n251 VNB 0.02fF
C373 VPB.n252 VNB 0.03fF
C374 VPB.n253 VNB 0.03fF
C375 VPB.n254 VNB 0.27fF
C376 VPB.n255 VNB 0.01fF
C377 VPB.n256 VNB 0.02fF
C378 VPB.n257 VNB 0.04fF
C379 VPB.n258 VNB 0.27fF
C380 VPB.n259 VNB 0.02fF
C381 VPB.n260 VNB 0.02fF
C382 VPB.n261 VNB 0.02fF
C383 VPB.n262 VNB 0.05fF
C384 VPB.n263 VNB 0.20fF
C385 VPB.n264 VNB 0.02fF
C386 VPB.n265 VNB 0.01fF
C387 VPB.n266 VNB 0.02fF
C388 VPB.n267 VNB 0.14fF
C389 VPB.n268 VNB 0.16fF
C390 VPB.n269 VNB 0.02fF
C391 VPB.n270 VNB 0.02fF
C392 VPB.n271 VNB 0.02fF
C393 VPB.n272 VNB 0.10fF
C394 VPB.n273 VNB 0.02fF
C395 VPB.n274 VNB 0.14fF
C396 VPB.n275 VNB 0.16fF
C397 VPB.n276 VNB 0.02fF
C398 VPB.n277 VNB 0.02fF
C399 VPB.n278 VNB 0.02fF
C400 VPB.n279 VNB 0.14fF
C401 VPB.n280 VNB 0.15fF
C402 VPB.n281 VNB 0.02fF
C403 VPB.n282 VNB 0.02fF
C404 VPB.n283 VNB 0.02fF
C405 VPB.n284 VNB 0.14fF
C406 VPB.n285 VNB 0.15fF
C407 VPB.n286 VNB 0.02fF
C408 VPB.n287 VNB 0.02fF
C409 VPB.n288 VNB 0.02fF
C410 VPB.n289 VNB 0.10fF
C411 VPB.n290 VNB 0.02fF
C412 VPB.n291 VNB 0.14fF
C413 VPB.n292 VNB 0.16fF
C414 VPB.n293 VNB 0.02fF
C415 VPB.n294 VNB 0.02fF
C416 VPB.n295 VNB 0.02fF
C417 VPB.n296 VNB 0.14fF
C418 VPB.n297 VNB 0.16fF
C419 VPB.n298 VNB 0.02fF
C420 VPB.n299 VNB 0.02fF
C421 VPB.n300 VNB 0.02fF
C422 VPB.n301 VNB 0.06fF
C423 VPB.n302 VNB 0.21fF
C424 VPB.n303 VNB 0.02fF
C425 VPB.n304 VNB 0.01fF
C426 VPB.n305 VNB 0.02fF
C427 VPB.n306 VNB 0.27fF
C428 VPB.n307 VNB 0.02fF
C429 VPB.n308 VNB 0.02fF
C430 VPB.n309 VNB 0.02fF
C431 VPB.n310 VNB 0.27fF
C432 VPB.n311 VNB 0.01fF
C433 VPB.n312 VNB 0.02fF
C434 VPB.n313 VNB 0.04fF
C435 VPB.n314 VNB 0.04fF
C436 VPB.n315 VNB 0.02fF
C437 VPB.n316 VNB 0.02fF
C438 VPB.n317 VNB 0.02fF
C439 VPB.n318 VNB 0.02fF
C440 VPB.n319 VNB 0.02fF
C441 VPB.n320 VNB 0.02fF
C442 VPB.n321 VNB 0.02fF
C443 VPB.n322 VNB 0.02fF
C444 VPB.n323 VNB 0.02fF
C445 VPB.n324 VNB 0.02fF
C446 VPB.n325 VNB 0.02fF
C447 VPB.n326 VNB 0.27fF
C448 VPB.n327 VNB 0.01fF
C449 VPB.n328 VNB 0.02fF
C450 VPB.n329 VNB 0.03fF
C451 VPB.n330 VNB 0.03fF
C452 VPB.n331 VNB 0.27fF
C453 VPB.n332 VNB 0.01fF
C454 VPB.n333 VNB 0.02fF
C455 VPB.n334 VNB 0.02fF
C456 VPB.n335 VNB 0.05fF
C457 VPB.n336 VNB 0.23fF
C458 VPB.n337 VNB 0.02fF
C459 VPB.n338 VNB 0.01fF
C460 VPB.n339 VNB 0.02fF
C461 VPB.n340 VNB 0.14fF
C462 VPB.n341 VNB 0.16fF
C463 VPB.n342 VNB 0.02fF
C464 VPB.n343 VNB 0.02fF
C465 VPB.n344 VNB 0.02fF
C466 VPB.n345 VNB 0.10fF
C467 VPB.n346 VNB 0.02fF
C468 VPB.n347 VNB 0.14fF
C469 VPB.n348 VNB 0.15fF
C470 VPB.n349 VNB 0.02fF
C471 VPB.n350 VNB 0.02fF
C472 VPB.n351 VNB 0.02fF
C473 VPB.n352 VNB 0.14fF
C474 VPB.n353 VNB 0.15fF
C475 VPB.n354 VNB 0.02fF
C476 VPB.n355 VNB 0.02fF
C477 VPB.n356 VNB 0.02fF
C478 VPB.n357 VNB 0.14fF
C479 VPB.n358 VNB 0.16fF
C480 VPB.n359 VNB 0.02fF
C481 VPB.n360 VNB 0.02fF
C482 VPB.n361 VNB 0.02fF
C483 VPB.n362 VNB 0.06fF
C484 VPB.n363 VNB 0.23fF
C485 VPB.n364 VNB 0.02fF
C486 VPB.n365 VNB 0.01fF
C487 VPB.n366 VNB 0.02fF
C488 VPB.n367 VNB 0.27fF
C489 VPB.n368 VNB 0.01fF
C490 VPB.n369 VNB 0.02fF
C491 VPB.n370 VNB 0.04fF
C492 VPB.n371 VNB 0.02fF
C493 VPB.n372 VNB 0.02fF
C494 VPB.n373 VNB 0.02fF
C495 VPB.n374 VNB 0.04fF
C496 VPB.n375 VNB 0.02fF
C497 VPB.n376 VNB 0.24fF
C498 VPB.n377 VNB 0.04fF
C499 VPB.n379 VNB 0.02fF
C500 VPB.n380 VNB 0.02fF
C501 VPB.n381 VNB 0.02fF
C502 VPB.n382 VNB 0.02fF
C503 VPB.n384 VNB 0.02fF
C504 VPB.n385 VNB 0.02fF
C505 VPB.n386 VNB 0.02fF
C506 VPB.n388 VNB 0.27fF
C507 VPB.n390 VNB 0.03fF
C508 VPB.n391 VNB 0.02fF
C509 VPB.n392 VNB 0.03fF
C510 VPB.n393 VNB 0.03fF
C511 VPB.n394 VNB 0.27fF
C512 VPB.n395 VNB 0.01fF
C513 VPB.n396 VNB 0.02fF
C514 VPB.n397 VNB 0.04fF
C515 VPB.n398 VNB 0.27fF
C516 VPB.n399 VNB 0.02fF
C517 VPB.n400 VNB 0.02fF
C518 VPB.n401 VNB 0.02fF
C519 VPB.n402 VNB 0.05fF
C520 VPB.n403 VNB 0.20fF
C521 VPB.n404 VNB 0.02fF
C522 VPB.n405 VNB 0.01fF
C523 VPB.n406 VNB 0.02fF
C524 VPB.n407 VNB 0.14fF
C525 VPB.n408 VNB 0.16fF
C526 VPB.n409 VNB 0.02fF
C527 VPB.n410 VNB 0.02fF
C528 VPB.n411 VNB 0.02fF
C529 VPB.n412 VNB 0.10fF
C530 VPB.n413 VNB 0.02fF
C531 VPB.n414 VNB 0.14fF
C532 VPB.n415 VNB 0.16fF
C533 VPB.n416 VNB 0.02fF
C534 VPB.n417 VNB 0.02fF
C535 VPB.n418 VNB 0.02fF
C536 VPB.n419 VNB 0.14fF
C537 VPB.n420 VNB 0.15fF
C538 VPB.n421 VNB 0.02fF
C539 VPB.n422 VNB 0.02fF
C540 VPB.n423 VNB 0.02fF
C541 VPB.n424 VNB 0.14fF
C542 VPB.n425 VNB 0.15fF
C543 VPB.n426 VNB 0.02fF
C544 VPB.n427 VNB 0.02fF
C545 VPB.n428 VNB 0.02fF
C546 VPB.n429 VNB 0.10fF
C547 VPB.n430 VNB 0.02fF
C548 VPB.n431 VNB 0.14fF
C549 VPB.n432 VNB 0.16fF
C550 VPB.n433 VNB 0.02fF
C551 VPB.n434 VNB 0.02fF
C552 VPB.n435 VNB 0.02fF
C553 VPB.n436 VNB 0.14fF
C554 VPB.n437 VNB 0.16fF
C555 VPB.n438 VNB 0.02fF
C556 VPB.n439 VNB 0.02fF
C557 VPB.n440 VNB 0.02fF
C558 VPB.n441 VNB 0.06fF
C559 VPB.n442 VNB 0.21fF
C560 VPB.n443 VNB 0.02fF
C561 VPB.n444 VNB 0.01fF
C562 VPB.n445 VNB 0.02fF
C563 VPB.n446 VNB 0.27fF
C564 VPB.n447 VNB 0.02fF
C565 VPB.n448 VNB 0.02fF
C566 VPB.n449 VNB 0.02fF
C567 VPB.n450 VNB 0.27fF
C568 VPB.n451 VNB 0.01fF
C569 VPB.n452 VNB 0.02fF
C570 VPB.n453 VNB 0.04fF
C571 VPB.n454 VNB 0.04fF
C572 VPB.n455 VNB 0.02fF
C573 VPB.n456 VNB 0.02fF
C574 VPB.n457 VNB 0.02fF
C575 VPB.n458 VNB 0.02fF
C576 VPB.n459 VNB 0.02fF
C577 VPB.n460 VNB 0.02fF
C578 VPB.n461 VNB 0.02fF
C579 VPB.n462 VNB 0.02fF
C580 VPB.n463 VNB 0.02fF
C581 VPB.n464 VNB 0.02fF
C582 VPB.n465 VNB 0.03fF
C583 VPB.n466 VNB 0.03fF
C584 VPB.n467 VNB 0.02fF
C585 VPB.n468 VNB 0.02fF
C586 VPB.n469 VNB 0.02fF
C587 VPB.n470 VNB 0.04fF
C588 VPB.n471 VNB 0.04fF
C589 VPB.n473 VNB 0.42fF
C590 a_277_1004.n0 VNB 0.74fF
C591 a_277_1004.n1 VNB 0.74fF
C592 a_277_1004.n2 VNB 0.87fF
C593 a_277_1004.n3 VNB 0.27fF
C594 a_277_1004.n4 VNB 0.40fF
C595 a_277_1004.n5 VNB 0.44fF
C596 a_277_1004.n6 VNB 0.82fF
C597 a_277_1004.n7 VNB 0.44fF
C598 a_277_1004.n8 VNB 0.65fF
C599 a_277_1004.n9 VNB 3.25fF
C600 a_277_1004.n10 VNB 0.63fF
C601 a_277_1004.n11 VNB 0.11fF
C602 a_277_1004.n12 VNB 0.42fF
C603 a_277_1004.n13 VNB 0.06fF
C604 a_147_159.n0 VNB 0.06fF
C605 a_147_159.n1 VNB 0.74fF
C606 a_147_159.n2 VNB 0.74fF
C607 a_147_159.n3 VNB 0.86fF
C608 a_147_159.n4 VNB 0.27fF
C609 a_147_159.n5 VNB 0.35fF
C610 a_147_159.n6 VNB 0.40fF
C611 a_147_159.t11 VNB 0.79fF
C612 a_147_159.n7 VNB 0.57fF
C613 a_147_159.n8 VNB 0.40fF
C614 a_147_159.t12 VNB 0.78fF
C615 a_147_159.n9 VNB 0.51fF
C616 a_147_159.n10 VNB 0.39fF
C617 a_147_159.n11 VNB 0.76fF
C618 a_147_159.n12 VNB 2.88fF
C619 a_147_159.n13 VNB 2.27fF
C620 a_147_159.n14 VNB 0.61fF
C621 a_147_159.n15 VNB 0.05fF
C622 a_147_159.n16 VNB 0.47fF
C623 a_147_159.n17 VNB 0.07fF
.ends
