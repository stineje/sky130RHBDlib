// File: INVX1.spi.INVX1.pxi
// Created: Tue Oct 15 15:49:25 2024
// 
simulator lang=spectre
x_PM_INVX1\%GND ( GND N_GND_c_3_p N_GND_c_4_p N_GND_c_12_p N_GND_c_1_p \
 N_GND_c_2_p N_GND_M0_noxref_s )  PM_INVX1\%GND
x_PM_INVX1\%VDD ( VDD N_VDD_c_45_p N_VDD_c_32_p N_VDD_c_27_n N_VDD_c_28_n \
 N_VDD_M1_noxref_s N_VDD_M2_noxref_d )  PM_INVX1\%VDD
x_PM_INVX1\%A ( A A A A A A A N_A_c_50_n N_A_M0_noxref_g N_A_M1_noxref_g \
 N_A_M2_noxref_g N_A_c_55_n N_A_c_85_p N_A_c_86_p N_A_c_57_n N_A_c_73_n \
 N_A_c_74_n N_A_c_58_n N_A_c_78_p N_A_c_59_n N_A_c_61_n N_A_c_62_n )  \
 PM_INVX1\%A
x_PM_INVX1\%Y ( Y Y Y Y Y Y Y N_Y_c_97_n N_Y_c_118_n N_Y_c_107_n N_Y_c_109_n \
 N_Y_M0_noxref_d N_Y_M1_noxref_d )  PM_INVX1\%Y
cc_1 ( N_GND_c_1_p N_VDD_c_27_n ) capacitor c=0.00989031f //x=0.63 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_28_n ) capacitor c=0.00989031f //x=1.6 //y=0 \
 //x2=1.48 //y2=7.4
cc_3 ( N_GND_c_3_p N_A_c_50_n ) capacitor c=0.00203213f //x=1.48 //y=0 \
 //x2=0.74 //y2=2.085
cc_4 ( N_GND_c_4_p N_A_c_50_n ) capacitor c=8.01092e-19 //x=1.03 //y=0.535 \
 //x2=0.74 //y2=2.085
cc_5 ( N_GND_c_1_p N_A_c_50_n ) capacitor c=0.0293771f //x=0.63 //y=0 \
 //x2=0.74 //y2=2.085
cc_6 ( N_GND_c_2_p N_A_c_50_n ) capacitor c=0.00118981f //x=1.6 //y=0 \
 //x2=0.74 //y2=2.085
cc_7 ( N_GND_M0_noxref_s N_A_c_50_n ) capacitor c=0.0107239f //x=0.495 \
 //y=0.37 //x2=0.74 //y2=2.085
cc_8 ( N_GND_c_4_p N_A_c_55_n ) capacitor c=0.0120496f //x=1.03 //y=0.535 \
 //x2=0.85 //y2=0.91
cc_9 ( N_GND_M0_noxref_s N_A_c_55_n ) capacitor c=0.0315727f //x=0.495 \
 //y=0.37 //x2=0.85 //y2=0.91
cc_10 ( N_GND_c_1_p N_A_c_57_n ) capacitor c=0.0124051f //x=0.63 //y=0 \
 //x2=0.85 //y2=1.92
cc_11 ( N_GND_M0_noxref_s N_A_c_58_n ) capacitor c=0.00483274f //x=0.495 \
 //y=0.37 //x2=1.225 //y2=0.755
cc_12 ( N_GND_c_12_p N_A_c_59_n ) capacitor c=0.0118602f //x=1.515 //y=0.535 \
 //x2=1.38 //y2=0.91
cc_13 ( N_GND_M0_noxref_s N_A_c_59_n ) capacitor c=0.0143355f //x=0.495 \
 //y=0.37 //x2=1.38 //y2=0.91
cc_14 ( N_GND_M0_noxref_s N_A_c_61_n ) capacitor c=0.0074042f //x=0.495 \
 //y=0.37 //x2=1.38 //y2=1.255
cc_15 ( N_GND_c_4_p N_A_c_62_n ) capacitor c=2.1838e-19 //x=1.03 //y=0.535 \
 //x2=0.74 //y2=2.085
cc_16 ( N_GND_c_1_p N_A_c_62_n ) capacitor c=0.0108179f //x=0.63 //y=0 \
 //x2=0.74 //y2=2.085
cc_17 ( N_GND_M0_noxref_s N_A_c_62_n ) capacitor c=0.00650244f //x=0.495 \
 //y=0.37 //x2=0.74 //y2=2.085
cc_18 ( N_GND_c_1_p Y ) capacitor c=8.10282e-19 //x=0.63 //y=0 //x2=1.48 \
 //y2=2.22
cc_19 ( N_GND_c_3_p N_Y_c_97_n ) capacitor c=0.0021242f //x=1.48 //y=0 \
 //x2=1.395 //y2=2.08
cc_20 ( N_GND_c_2_p N_Y_c_97_n ) capacitor c=0.0301661f //x=1.6 //y=0 \
 //x2=1.395 //y2=2.08
cc_21 ( N_GND_M0_noxref_s N_Y_c_97_n ) capacitor c=0.00999304f //x=0.495 \
 //y=0.37 //x2=1.395 //y2=2.08
cc_22 ( N_GND_c_3_p N_Y_M0_noxref_d ) capacitor c=0.00194883f //x=1.48 //y=0 \
 //x2=0.925 //y2=0.91
cc_23 ( N_GND_c_4_p N_Y_M0_noxref_d ) capacitor c=0.0146043f //x=1.03 \
 //y=0.535 //x2=0.925 //y2=0.91
cc_24 ( N_GND_c_1_p N_Y_M0_noxref_d ) capacitor c=0.0094373f //x=0.63 //y=0 \
 //x2=0.925 //y2=0.91
cc_25 ( N_GND_c_2_p N_Y_M0_noxref_d ) capacitor c=0.00973758f //x=1.6 //y=0 \
 //x2=0.925 //y2=0.91
cc_26 ( N_GND_M0_noxref_s N_Y_M0_noxref_d ) capacitor c=0.076995f //x=0.495 \
 //y=0.37 //x2=0.925 //y2=0.91
cc_27 ( N_VDD_c_27_n N_A_c_50_n ) capacitor c=0.0276175f //x=0.74 //y=7.4 \
 //x2=0.74 //y2=2.085
cc_28 ( N_VDD_c_28_n N_A_c_50_n ) capacitor c=0.00144809f //x=1.48 //y=7.4 \
 //x2=0.74 //y2=2.085
cc_29 ( N_VDD_M1_noxref_s N_A_c_50_n ) capacitor c=0.00938034f //x=0.54 \
 //y=5.02 //x2=0.74 //y2=2.085
cc_30 ( N_VDD_c_32_p N_A_M1_noxref_g ) capacitor c=0.00748034f //x=1.47 \
 //y=7.4 //x2=0.895 //y2=6.02
cc_31 ( N_VDD_c_27_n N_A_M1_noxref_g ) capacitor c=0.0241676f //x=0.74 //y=7.4 \
 //x2=0.895 //y2=6.02
cc_32 ( N_VDD_M1_noxref_s N_A_M1_noxref_g ) capacitor c=0.0528676f //x=0.54 \
 //y=5.02 //x2=0.895 //y2=6.02
cc_33 ( N_VDD_c_32_p N_A_M2_noxref_g ) capacitor c=0.00697478f //x=1.47 \
 //y=7.4 //x2=1.335 //y2=6.02
cc_34 ( N_VDD_M2_noxref_d N_A_M2_noxref_g ) capacitor c=0.0528676f //x=1.41 \
 //y=5.02 //x2=1.335 //y2=6.02
cc_35 ( N_VDD_c_28_n N_A_c_73_n ) capacitor c=0.0287802f //x=1.48 //y=7.4 \
 //x2=1.26 //y2=4.79
cc_36 ( N_VDD_c_27_n N_A_c_74_n ) capacitor c=0.011132f //x=0.74 //y=7.4 \
 //x2=0.97 //y2=4.79
cc_37 ( N_VDD_M1_noxref_s N_A_c_74_n ) capacitor c=0.00665831f //x=0.54 \
 //y=5.02 //x2=0.97 //y2=4.79
cc_38 ( N_VDD_c_27_n Y ) capacitor c=4.80934e-19 //x=0.74 //y=7.4 //x2=1.48 \
 //y2=2.22
cc_39 ( N_VDD_c_28_n Y ) capacitor c=0.0232778f //x=1.48 //y=7.4 //x2=1.48 \
 //y2=2.22
cc_40 ( N_VDD_c_32_p N_Y_c_107_n ) capacitor c=8.92854e-19 //x=1.47 //y=7.4 \
 //x2=1.395 //y2=4.58
cc_41 ( N_VDD_M2_noxref_d N_Y_c_107_n ) capacitor c=0.00644908f //x=1.41 \
 //y=5.02 //x2=1.395 //y2=4.58
cc_42 ( N_VDD_c_27_n N_Y_c_109_n ) capacitor c=0.0179238f //x=0.74 //y=7.4 \
 //x2=1.2 //y2=4.58
cc_43 ( N_VDD_c_45_p N_Y_M1_noxref_d ) capacitor c=0.00722811f //x=1.48 \
 //y=7.4 //x2=0.97 //y2=5.02
cc_44 ( N_VDD_c_32_p N_Y_M1_noxref_d ) capacitor c=0.0139004f //x=1.47 //y=7.4 \
 //x2=0.97 //y2=5.02
cc_45 ( N_VDD_c_28_n N_Y_M1_noxref_d ) capacitor c=0.0219131f //x=1.48 //y=7.4 \
 //x2=0.97 //y2=5.02
cc_46 ( N_VDD_M1_noxref_s N_Y_M1_noxref_d ) capacitor c=0.0843065f //x=0.54 \
 //y=5.02 //x2=0.97 //y2=5.02
cc_47 ( N_VDD_M2_noxref_d N_Y_M1_noxref_d ) capacitor c=0.0832641f //x=1.41 \
 //y=5.02 //x2=0.97 //y2=5.02
cc_48 ( N_A_c_50_n Y ) capacitor c=0.0739084f //x=0.74 //y=2.085 //x2=1.48 \
 //y2=2.22
cc_49 ( N_A_c_62_n Y ) capacitor c=8.49451e-19 //x=0.74 //y=2.085 //x2=1.48 \
 //y2=2.22
cc_50 ( N_A_c_78_p N_Y_c_97_n ) capacitor c=0.0023507f //x=1.225 //y=1.41 \
 //x2=1.395 //y2=2.08
cc_51 ( N_A_c_62_n N_Y_c_118_n ) capacitor c=0.0167852f //x=0.74 //y=2.085 \
 //x2=1.195 //y2=2.08
cc_52 ( N_A_c_73_n N_Y_c_107_n ) capacitor c=0.0107726f //x=1.26 //y=4.79 \
 //x2=1.395 //y2=4.58
cc_53 ( N_A_c_50_n N_Y_c_109_n ) capacitor c=0.0250789f //x=0.74 //y=2.085 \
 //x2=1.2 //y2=4.58
cc_54 ( N_A_c_74_n N_Y_c_109_n ) capacitor c=0.00962086f //x=0.97 //y=4.79 \
 //x2=1.2 //y2=4.58
cc_55 ( N_A_c_50_n N_Y_M0_noxref_d ) capacitor c=0.0175773f //x=0.74 //y=2.085 \
 //x2=0.925 //y2=0.91
cc_56 ( N_A_c_55_n N_Y_M0_noxref_d ) capacitor c=0.00218556f //x=0.85 //y=0.91 \
 //x2=0.925 //y2=0.91
cc_57 ( N_A_c_85_p N_Y_M0_noxref_d ) capacitor c=0.00347355f //x=0.85 \
 //y=1.255 //x2=0.925 //y2=0.91
cc_58 ( N_A_c_86_p N_Y_M0_noxref_d ) capacitor c=0.00742431f //x=0.85 \
 //y=1.565 //x2=0.925 //y2=0.91
cc_59 ( N_A_c_57_n N_Y_M0_noxref_d ) capacitor c=0.00957707f //x=0.85 //y=1.92 \
 //x2=0.925 //y2=0.91
cc_60 ( N_A_c_58_n N_Y_M0_noxref_d ) capacitor c=0.00220879f //x=1.225 \
 //y=0.755 //x2=0.925 //y2=0.91
cc_61 ( N_A_c_78_p N_Y_M0_noxref_d ) capacitor c=0.0138447f //x=1.225 //y=1.41 \
 //x2=0.925 //y2=0.91
cc_62 ( N_A_c_59_n N_Y_M0_noxref_d ) capacitor c=0.00218624f //x=1.38 //y=0.91 \
 //x2=0.925 //y2=0.91
cc_63 ( N_A_c_61_n N_Y_M0_noxref_d ) capacitor c=0.00601286f //x=1.38 \
 //y=1.255 //x2=0.925 //y2=0.91
cc_64 ( N_A_M1_noxref_g N_Y_M1_noxref_d ) capacitor c=0.0219309f //x=0.895 \
 //y=6.02 //x2=0.97 //y2=5.02
cc_65 ( N_A_M2_noxref_g N_Y_M1_noxref_d ) capacitor c=0.021902f //x=1.335 \
 //y=6.02 //x2=0.97 //y2=5.02
cc_66 ( N_A_c_73_n N_Y_M1_noxref_d ) capacitor c=0.0148755f //x=1.26 //y=4.79 \
 //x2=0.97 //y2=5.02
cc_67 ( N_A_c_74_n N_Y_M1_noxref_d ) capacitor c=0.00307344f //x=0.97 //y=4.79 \
 //x2=0.97 //y2=5.02
