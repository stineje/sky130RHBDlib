* SPICE3 file created from FA.ext - technology: sky130A

.subckt FA SUM COUT A B CIN VDD GND
X0 COUT or2x1_pcell_0/m1_547_649# VSUBS VSUBS nshort w=3 l=0.15
X1 VDD or2x1_pcell_0/m1_547_649# COUT VDD pshort w=2 l=0.15
X2 VDD m1_5455_575# or2x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X3 or2x1_pcell_0/m1_547_649# m1_6565_649# or2x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X4 or2x1_pcell_0/m1_547_649# m1_5455_575# VSUBS VSUBS nshort w=3 l=0.15
X5 or2x1_pcell_0/m1_547_649# m1_6565_649# VSUBS VSUBS nshort w=3 l=0.15
X6 GND A xor2X1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X7 GND xor2X1_pcell_0/m1_939_797# xor2X1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X8 VDD A xor2X1_pcell_0/a_761_1330# VDD pshort w=2 l=0.15
X9 m1_2421_427# xor2X1_pcell_0/m1_315_501# xor2X1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X10 m1_2421_427# B xor2X1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X11 m1_2421_427# xor2X1_pcell_0/m1_939_797# xor2X1_pcell_0/a_761_1330# VDD pshort w=2 l=0.15
X12 VDD B xor2X1_pcell_0/a_1427_1330# VDD pshort w=2 l=0.15
X13 m1_2421_427# xor2X1_pcell_0/m1_315_501# xor2X1_pcell_0/a_1427_1330# VDD pshort w=2 l=0.15
X14 xor2X1_pcell_0/m1_315_501# A GND GND nshort w=3 l=0.15
X15 VDD A xor2X1_pcell_0/m1_315_501# VDD pshort w=2 l=0.15
X16 xor2X1_pcell_0/m1_939_797# B xor2X1_pcell_0/li1_M1_contact_2/VSUBS xor2X1_pcell_0/li1_M1_contact_2/VSUBS nshort w=3 l=0.15
X17 VDD B xor2X1_pcell_0/m1_939_797# VDD pshort w=2 l=0.15
X18 m1_5455_575# and2x1_pcell_0/m1_547_649# VSUBS VSUBS nshort w=3 l=0.15
X19 VDD and2x1_pcell_0/m1_547_649# m1_5455_575# VDD pshort w=2 l=0.15
X20 VSUBS CIN and2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# VSUBS nshort w=3 l=0.15
X21 and2x1_pcell_0/m1_547_649# m1_2421_427# and2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# VSUBS nshort w=3 l=0.15
X22 VDD CIN and2x1_pcell_0/m1_547_649# VDD pshort w=2 l=0.15
X23 VDD m1_2421_427# and2x1_pcell_0/m1_547_649# VDD pshort w=2 l=0.15
X24 xor2X1_pcell_1/pmos2_1_3/VSUBS m1_2421_427# xor2X1_pcell_1/nmos_bottom_0/a_0_0# xor2X1_pcell_1/pmos2_1_3/VSUBS nshort w=3 l=0.15
X25 xor2X1_pcell_1/pmos2_1_3/VSUBS xor2X1_pcell_1/m1_939_797# xor2X1_pcell_1/nmos_bottom_1/a_0_0# xor2X1_pcell_1/pmos2_1_3/VSUBS nshort w=3 l=0.15
X26 VDD m1_2421_427# xor2X1_pcell_1/a_761_1330# VDD pshort w=2 l=0.15
X27 SUM xor2X1_pcell_1/m1_315_501# xor2X1_pcell_1/nmos_bottom_1/a_0_0# xor2X1_pcell_1/pmos2_1_3/VSUBS nshort w=3 l=0.15
X28 SUM CIN xor2X1_pcell_1/nmos_bottom_0/a_0_0# xor2X1_pcell_1/pmos2_1_3/VSUBS nshort w=3 l=0.15
X29 SUM xor2X1_pcell_1/m1_939_797# xor2X1_pcell_1/a_761_1330# VDD pshort w=2 l=0.15
X30 VDD CIN xor2X1_pcell_1/a_1427_1330# VDD pshort w=2 l=0.15
X31 SUM xor2X1_pcell_1/m1_315_501# xor2X1_pcell_1/a_1427_1330# VDD pshort w=2 l=0.15
X32 xor2X1_pcell_1/m1_315_501# m1_2421_427# xor2X1_pcell_1/pmos2_1_3/VSUBS xor2X1_pcell_1/pmos2_1_3/VSUBS nshort w=3 l=0.15
X33 VDD m1_2421_427# xor2X1_pcell_1/m1_315_501# VDD pshort w=2 l=0.15
X34 xor2X1_pcell_1/m1_939_797# CIN xor2X1_pcell_1/li1_M1_contact_2/VSUBS xor2X1_pcell_1/li1_M1_contact_2/VSUBS nshort w=3 l=0.15
X35 VDD CIN xor2X1_pcell_1/m1_939_797# VDD pshort w=2 l=0.15
X36 m1_6565_649# and2x1_pcell_1/m1_547_649# VSUBS VSUBS nshort w=3 l=0.15
X37 VDD and2x1_pcell_1/m1_547_649# m1_6565_649# VDD pshort w=2 l=0.15
X38 VSUBS B and2x1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# VSUBS nshort w=3 l=0.15
X39 and2x1_pcell_1/m1_547_649# A and2x1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# VSUBS nshort w=3 l=0.15
X40 VDD B and2x1_pcell_1/m1_547_649# VDD pshort w=2 l=0.15
X41 VDD A and2x1_pcell_1/m1_547_649# VDD pshort w=2 l=0.15
C0 VDD xor2X1_pcell_1/li1_M1_contact_2/VSUBS 15.33fF
.ends
