* SPICE3 file created from XOR2X1.ext - technology: sky130A

.subckt XOR2X1 Y A B VDD GND
M1000 Y a_185_209.t4 a_1222_101.t1 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.14u as=0p ps=0u
M1001 a_575_1051.t1 A.t2 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y.t1 a_185_209.t3 a_1241_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t1 B.t0 a_807_990.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_807_990.t0 B.t1 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_185_209.t1 A.t3 VDD.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B.t3 a_556_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_575_1051.t2 a_807_990.t3 Y.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1241_1051.t3 B.t4 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y.t5 a_807_990.t4 a_575_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1241_1051.t1 a_185_209.t5 Y.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 GND a_807_990.t5 a_1222_101.t0 nshort w=-1.605u l=1.765u
+  ad=2.6398p pd=19.34u as=0p ps=0u
M1012 VDD.t5 A.t4 a_575_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VDD.t6 A.t5 a_185_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 GND A.t1 a_556_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD.t2 B.t5 a_1241_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 B Y 0.62fF
C1 B A 0.04fF
C2 VDD Y 0.53fF
C3 VDD A 0.50fF
C4 Y A 0.08fF
C5 B VDD 0.60fF
R0 A.n2 A.t5 512.525
R1 A.n0 A.t2 480.392
R2 A.n0 A.t4 403.272
R3 A.n2 A.t3 371.139
R4 A.n1 A.t1 336.586
R5 A.n3 A.t0 290.093
R6 A.n3 A.n2 93.541
R7 A.n4 A.n1 77.859
R8 A.n4 A.n3 76
R9 A.n1 A.n0 45.7
R10 A.n4 A 0.046
R11 GND.n27 GND.n25 219.745
R12 GND.n89 GND.n88 219.745
R13 GND.n118 GND.n117 219.745
R14 GND.n27 GND.n26 85.529
R15 GND.n89 GND.n87 85.529
R16 GND.n118 GND.n116 85.529
R17 GND.n45 GND.n44 84.842
R18 GND.n8 GND.n1 76.145
R19 GND.n57 GND.n56 76
R20 GND.n8 GND.n7 76
R21 GND.n14 GND.n13 76
R22 GND.n21 GND.n20 76
R23 GND.n24 GND.n23 76
R24 GND.n31 GND.n30 76
R25 GND.n34 GND.n33 76
R26 GND.n37 GND.n36 76
R27 GND.n40 GND.n39 76
R28 GND.n43 GND.n42 76
R29 GND.n48 GND.n47 76
R30 GND.n51 GND.n50 76
R31 GND.n54 GND.n53 76
R32 GND.n122 GND.n121 76
R33 GND.n115 GND.n114 76
R34 GND.n112 GND.n111 76
R35 GND.n109 GND.n108 76
R36 GND.n106 GND.n105 76
R37 GND.n103 GND.n102 76
R38 GND.n95 GND.n94 76
R39 GND.n92 GND.n91 76
R40 GND.n85 GND.n84 76
R41 GND.n82 GND.n81 76
R42 GND.n74 GND.n73 76
R43 GND.n66 GND.n65 76
R44 GND.n100 GND.n99 63.835
R45 GND.n62 GND.t2 39.412
R46 GND.n78 GND.n77 35.01
R47 GND.n99 GND.n98 28.421
R48 GND.n99 GND.n97 25.263
R49 GND.n97 GND.n96 24.383
R50 GND.n5 GND.n4 19.735
R51 GND.n12 GND.n11 19.735
R52 GND.n19 GND.n18 19.735
R53 GND.n79 GND.n78 19.735
R54 GND.n71 GND.n70 19.735
R55 GND.n64 GND.n63 19.735
R56 GND.n78 GND.n76 19.017
R57 GND.n10 GND.t0 18.552
R58 GND.n62 GND.n61 17.185
R59 GND.n30 GND.n28 14.167
R60 GND.n121 GND.n119 14.167
R61 GND.n91 GND.n90 14.167
R62 GND.n65 GND.n58 13.653
R63 GND.n73 GND.n72 13.653
R64 GND.n81 GND.n80 13.653
R65 GND.n84 GND.n83 13.653
R66 GND.n91 GND.n86 13.653
R67 GND.n94 GND.n93 13.653
R68 GND.n102 GND.n101 13.653
R69 GND.n105 GND.n104 13.653
R70 GND.n108 GND.n107 13.653
R71 GND.n111 GND.n110 13.653
R72 GND.n114 GND.n113 13.653
R73 GND.n121 GND.n120 13.653
R74 GND.n53 GND.n52 13.653
R75 GND.n50 GND.n49 13.653
R76 GND.n47 GND.n46 13.653
R77 GND.n42 GND.n41 13.653
R78 GND.n39 GND.n38 13.653
R79 GND.n36 GND.n35 13.653
R80 GND.n33 GND.n32 13.653
R81 GND.n30 GND.n29 13.653
R82 GND.n23 GND.n22 13.653
R83 GND.n20 GND.n15 13.653
R84 GND.n13 GND.n9 13.653
R85 GND.n7 GND.n6 13.653
R86 GND.n18 GND.n17 13.608
R87 GND.n4 GND.n3 10.853
R88 GND.n3 GND.n2 10.417
R89 GND.n17 GND.n16 7.858
R90 GND.n76 GND.n75 7.5
R91 GND.n69 GND.n68 7.5
R92 GND.n28 GND.n27 7.312
R93 GND.n90 GND.n89 7.312
R94 GND.n119 GND.n118 7.312
R95 GND.n63 GND.n62 6.139
R96 GND.n60 GND.n59 4.551
R97 GND.n20 GND.n19 3.935
R98 GND.n47 GND.n45 3.935
R99 GND.n102 GND.n100 3.935
R100 GND.n81 GND.n79 3.935
R101 GND.n7 GND.n5 3.541
R102 GND.n65 GND.n64 3.541
R103 GND.t2 GND.n60 2.238
R104 GND.n68 GND.n67 1.935
R105 GND.n1 GND.n0 0.596
R106 GND.n56 GND.n55 0.596
R107 GND.n11 GND.n10 0.358
R108 GND.n70 GND.n69 0.358
R109 GND.n31 GND.n24 0.29
R110 GND.n92 GND.n85 0.29
R111 GND.n57 GND 0.207
R112 GND.n13 GND.n12 0.196
R113 GND.n73 GND.n71 0.196
R114 GND.n43 GND.n40 0.181
R115 GND.n109 GND.n106 0.181
R116 GND.n14 GND.n8 0.157
R117 GND.n21 GND.n14 0.157
R118 GND.n82 GND.n74 0.157
R119 GND.n74 GND.n66 0.157
R120 GND.n24 GND.n21 0.145
R121 GND.n34 GND.n31 0.145
R122 GND.n37 GND.n34 0.145
R123 GND.n40 GND.n37 0.145
R124 GND.n48 GND.n43 0.145
R125 GND.n51 GND.n48 0.145
R126 GND.n54 GND.n51 0.145
R127 GND GND.n54 0.145
R128 GND GND.n122 0.145
R129 GND.n122 GND.n115 0.145
R130 GND.n115 GND.n112 0.145
R131 GND.n112 GND.n109 0.145
R132 GND.n106 GND.n103 0.145
R133 GND.n103 GND.n95 0.145
R134 GND.n95 GND.n92 0.145
R135 GND.n85 GND.n82 0.145
R136 GND.n66 GND.n57 0.145
R137 a_185_209.n1 a_185_209.t3 477.179
R138 a_185_209.n1 a_185_209.t5 406.485
R139 a_185_209.n2 a_185_209.t4 269.148
R140 a_185_209.n5 a_185_209.n3 185.537
R141 a_185_209.n3 a_185_209.n0 184.007
R142 a_185_209.n3 a_185_209.n2 156.579
R143 a_185_209.n2 a_185_209.n1 125.359
R144 a_185_209.n5 a_185_209.n4 15.218
R145 a_185_209.n0 a_185_209.t0 14.282
R146 a_185_209.n0 a_185_209.t1 14.282
R147 a_185_209.n6 a_185_209.n5 12.014
R148 a_556_101.t0 a_556_101.n1 34.62
R149 a_556_101.t0 a_556_101.n0 8.137
R150 a_556_101.t0 a_556_101.n2 4.69
R151 VDD.n170 VDD.n168 144.705
R152 VDD.n68 VDD.n66 144.705
R153 VDD.n101 VDD.n99 144.705
R154 VDD.n26 VDD.n25 77.792
R155 VDD.n36 VDD.n35 77.792
R156 VDD.n160 VDD.n159 77.792
R157 VDD.n149 VDD.n148 77.792
R158 VDD.n29 VDD.n23 76.145
R159 VDD.n29 VDD.n28 76
R160 VDD.n33 VDD.n32 76
R161 VDD.n39 VDD.n38 76
R162 VDD.n43 VDD.n42 76
R163 VDD.n70 VDD.n69 76
R164 VDD.n74 VDD.n73 76
R165 VDD.n78 VDD.n77 76
R166 VDD.n82 VDD.n81 76
R167 VDD.n87 VDD.n86 76
R168 VDD.n94 VDD.n93 76
R169 VDD.n98 VDD.n97 76
R170 VDD.n124 VDD.n123 76
R171 VDD.n226 VDD.n225 76
R172 VDD.n222 VDD.n221 76
R173 VDD.n218 VDD.n217 76
R174 VDD.n214 VDD.n213 76
R175 VDD.n210 VDD.n209 76
R176 VDD.n205 VDD.n204 76
R177 VDD.n198 VDD.n197 76
R178 VDD.n194 VDD.n193 76
R179 VDD.n167 VDD.n166 76
R180 VDD.n163 VDD.n162 76
R181 VDD.n157 VDD.n156 76
R182 VDD.n153 VDD.n152 76
R183 VDD.n147 VDD.n146 76
R184 VDD.n200 VDD.n199 65.585
R185 VDD.n89 VDD.n88 65.585
R186 VDD.n151 VDD.t7 55.106
R187 VDD.n158 VDD.t6 55.106
R188 VDD.n34 VDD.t0 55.106
R189 VDD.n24 VDD.t1 55.106
R190 VDD.n106 VDD.n105 36.774
R191 VDD.n48 VDD.n47 36.774
R192 VDD.n186 VDD.n185 36.774
R193 VDD.n91 VDD.n90 32.032
R194 VDD.n202 VDD.n201 32.032
R195 VDD.n146 VDD.n143 21.841
R196 VDD.n23 VDD.n20 21.841
R197 VDD.n199 VDD.t4 14.282
R198 VDD.n199 VDD.t5 14.282
R199 VDD.n88 VDD.t3 14.282
R200 VDD.n88 VDD.t2 14.282
R201 VDD.n143 VDD.n126 14.167
R202 VDD.n126 VDD.n125 14.167
R203 VDD.n121 VDD.n103 14.167
R204 VDD.n103 VDD.n102 14.167
R205 VDD.n64 VDD.n45 14.167
R206 VDD.n45 VDD.n44 14.167
R207 VDD.n191 VDD.n172 14.167
R208 VDD.n172 VDD.n171 14.167
R209 VDD.n20 VDD.n19 14.167
R210 VDD.n19 VDD.n17 14.167
R211 VDD.n69 VDD.n65 14.167
R212 VDD.n123 VDD.n122 14.167
R213 VDD.n193 VDD.n192 14.167
R214 VDD.n23 VDD.n22 13.653
R215 VDD.n22 VDD.n21 13.653
R216 VDD.n28 VDD.n27 13.653
R217 VDD.n27 VDD.n26 13.653
R218 VDD.n32 VDD.n31 13.653
R219 VDD.n31 VDD.n30 13.653
R220 VDD.n38 VDD.n37 13.653
R221 VDD.n37 VDD.n36 13.653
R222 VDD.n42 VDD.n41 13.653
R223 VDD.n41 VDD.n40 13.653
R224 VDD.n69 VDD.n68 13.653
R225 VDD.n68 VDD.n67 13.653
R226 VDD.n73 VDD.n72 13.653
R227 VDD.n72 VDD.n71 13.653
R228 VDD.n77 VDD.n76 13.653
R229 VDD.n76 VDD.n75 13.653
R230 VDD.n81 VDD.n80 13.653
R231 VDD.n80 VDD.n79 13.653
R232 VDD.n86 VDD.n85 13.653
R233 VDD.n85 VDD.n84 13.653
R234 VDD.n93 VDD.n92 13.653
R235 VDD.n92 VDD.n91 13.653
R236 VDD.n97 VDD.n96 13.653
R237 VDD.n96 VDD.n95 13.653
R238 VDD.n123 VDD.n101 13.653
R239 VDD.n101 VDD.n100 13.653
R240 VDD.n225 VDD.n224 13.653
R241 VDD.n224 VDD.n223 13.653
R242 VDD.n221 VDD.n220 13.653
R243 VDD.n220 VDD.n219 13.653
R244 VDD.n217 VDD.n216 13.653
R245 VDD.n216 VDD.n215 13.653
R246 VDD.n213 VDD.n212 13.653
R247 VDD.n212 VDD.n211 13.653
R248 VDD.n209 VDD.n208 13.653
R249 VDD.n208 VDD.n207 13.653
R250 VDD.n204 VDD.n203 13.653
R251 VDD.n203 VDD.n202 13.653
R252 VDD.n197 VDD.n196 13.653
R253 VDD.n196 VDD.n195 13.653
R254 VDD.n193 VDD.n170 13.653
R255 VDD.n170 VDD.n169 13.653
R256 VDD.n166 VDD.n165 13.653
R257 VDD.n165 VDD.n164 13.653
R258 VDD.n162 VDD.n161 13.653
R259 VDD.n161 VDD.n160 13.653
R260 VDD.n156 VDD.n155 13.653
R261 VDD.n155 VDD.n154 13.653
R262 VDD.n152 VDD.n150 13.653
R263 VDD.n150 VDD.n149 13.653
R264 VDD.n146 VDD.n145 13.653
R265 VDD.n145 VDD.n144 13.653
R266 VDD.n4 VDD.n2 12.915
R267 VDD.n4 VDD.n3 12.66
R268 VDD.n13 VDD.n12 12.343
R269 VDD.n10 VDD.n9 12.343
R270 VDD.n10 VDD.n7 12.343
R271 VDD.n122 VDD.n121 7.674
R272 VDD.n65 VDD.n64 7.674
R273 VDD.n192 VDD.n191 7.674
R274 VDD.n59 VDD.n58 7.5
R275 VDD.n53 VDD.n52 7.5
R276 VDD.n55 VDD.n54 7.5
R277 VDD.n50 VDD.n49 7.5
R278 VDD.n64 VDD.n63 7.5
R279 VDD.n116 VDD.n115 7.5
R280 VDD.n110 VDD.n109 7.5
R281 VDD.n112 VDD.n111 7.5
R282 VDD.n118 VDD.n108 7.5
R283 VDD.n118 VDD.n106 7.5
R284 VDD.n121 VDD.n120 7.5
R285 VDD.n176 VDD.n175 7.5
R286 VDD.n179 VDD.n178 7.5
R287 VDD.n181 VDD.n180 7.5
R288 VDD.n184 VDD.n183 7.5
R289 VDD.n191 VDD.n190 7.5
R290 VDD.n138 VDD.n137 7.5
R291 VDD.n132 VDD.n131 7.5
R292 VDD.n134 VDD.n133 7.5
R293 VDD.n140 VDD.n130 7.5
R294 VDD.n140 VDD.n128 7.5
R295 VDD.n143 VDD.n142 7.5
R296 VDD.n20 VDD.n16 7.5
R297 VDD.n2 VDD.n1 7.5
R298 VDD.n9 VDD.n8 7.5
R299 VDD.n7 VDD.n6 7.5
R300 VDD.n19 VDD.n18 7.5
R301 VDD.n14 VDD.n0 7.5
R302 VDD.n51 VDD.n48 6.772
R303 VDD.n62 VDD.n46 6.772
R304 VDD.n60 VDD.n57 6.772
R305 VDD.n56 VDD.n53 6.772
R306 VDD.n119 VDD.n104 6.772
R307 VDD.n117 VDD.n114 6.772
R308 VDD.n113 VDD.n110 6.772
R309 VDD.n141 VDD.n127 6.772
R310 VDD.n139 VDD.n136 6.772
R311 VDD.n135 VDD.n132 6.772
R312 VDD.n51 VDD.n50 6.772
R313 VDD.n56 VDD.n55 6.772
R314 VDD.n60 VDD.n59 6.772
R315 VDD.n63 VDD.n62 6.772
R316 VDD.n113 VDD.n112 6.772
R317 VDD.n117 VDD.n116 6.772
R318 VDD.n120 VDD.n119 6.772
R319 VDD.n135 VDD.n134 6.772
R320 VDD.n139 VDD.n138 6.772
R321 VDD.n142 VDD.n141 6.772
R322 VDD.n190 VDD.n189 6.772
R323 VDD.n177 VDD.n174 6.772
R324 VDD.n182 VDD.n179 6.772
R325 VDD.n187 VDD.n184 6.772
R326 VDD.n187 VDD.n186 6.772
R327 VDD.n182 VDD.n181 6.772
R328 VDD.n177 VDD.n176 6.772
R329 VDD.n189 VDD.n173 6.772
R330 VDD.n16 VDD.n15 6.458
R331 VDD.n108 VDD.n107 6.202
R332 VDD.n130 VDD.n129 6.202
R333 VDD.n93 VDD.n89 5.903
R334 VDD.n204 VDD.n200 5.903
R335 VDD.n84 VDD.n83 4.576
R336 VDD.n207 VDD.n206 4.576
R337 VDD.n28 VDD.n24 1.967
R338 VDD.n38 VDD.n34 1.967
R339 VDD.n162 VDD.n158 1.967
R340 VDD.n152 VDD.n151 1.967
R341 VDD.n14 VDD.n5 1.329
R342 VDD.n14 VDD.n10 1.329
R343 VDD.n14 VDD.n11 1.329
R344 VDD.n14 VDD.n13 1.329
R345 VDD.n15 VDD.n14 0.696
R346 VDD.n14 VDD.n4 0.696
R347 VDD.n61 VDD.n60 0.365
R348 VDD.n61 VDD.n56 0.365
R349 VDD.n61 VDD.n51 0.365
R350 VDD.n62 VDD.n61 0.365
R351 VDD.n118 VDD.n117 0.365
R352 VDD.n118 VDD.n113 0.365
R353 VDD.n119 VDD.n118 0.365
R354 VDD.n140 VDD.n139 0.365
R355 VDD.n140 VDD.n135 0.365
R356 VDD.n141 VDD.n140 0.365
R357 VDD.n188 VDD.n187 0.365
R358 VDD.n188 VDD.n182 0.365
R359 VDD.n188 VDD.n177 0.365
R360 VDD.n189 VDD.n188 0.365
R361 VDD.n70 VDD.n43 0.29
R362 VDD.n194 VDD.n167 0.29
R363 VDD.n147 VDD 0.207
R364 VDD.n87 VDD.n82 0.181
R365 VDD.n214 VDD.n210 0.181
R366 VDD.n33 VDD.n29 0.157
R367 VDD.n39 VDD.n33 0.157
R368 VDD.n163 VDD.n157 0.157
R369 VDD.n157 VDD.n153 0.157
R370 VDD.n43 VDD.n39 0.145
R371 VDD.n74 VDD.n70 0.145
R372 VDD.n78 VDD.n74 0.145
R373 VDD.n82 VDD.n78 0.145
R374 VDD.n94 VDD.n87 0.145
R375 VDD.n98 VDD.n94 0.145
R376 VDD.n124 VDD.n98 0.145
R377 VDD VDD.n124 0.145
R378 VDD VDD.n226 0.145
R379 VDD.n226 VDD.n222 0.145
R380 VDD.n222 VDD.n218 0.145
R381 VDD.n218 VDD.n214 0.145
R382 VDD.n210 VDD.n205 0.145
R383 VDD.n205 VDD.n198 0.145
R384 VDD.n198 VDD.n194 0.145
R385 VDD.n167 VDD.n163 0.145
R386 VDD.n153 VDD.n147 0.145
R387 a_575_1051.n0 a_575_1051.t2 101.66
R388 a_575_1051.n0 a_575_1051.t0 101.66
R389 a_575_1051.n0 a_575_1051.t3 14.294
R390 a_575_1051.t1 a_575_1051.n0 14.282
R391 a_1241_1051.n0 a_1241_1051.t1 101.66
R392 a_1241_1051.n0 a_1241_1051.t2 101.66
R393 a_1241_1051.t0 a_1241_1051.n0 14.294
R394 a_1241_1051.n0 a_1241_1051.t3 14.282
R395 Y.n8 Y.n7 232.332
R396 Y.n5 Y.n4 210.593
R397 Y.n5 Y.n0 165.336
R398 Y.n8 Y.n6 165.336
R399 Y Y.n8 78.357
R400 Y.n9 Y.n5 76
R401 Y.n4 Y.n3 30
R402 Y.n2 Y.n1 24.383
R403 Y.n4 Y.n2 23.684
R404 Y.n0 Y.t0 14.282
R405 Y.n0 Y.t1 14.282
R406 Y.n6 Y.t4 14.282
R407 Y.n6 Y.t5 14.282
R408 Y.n9 Y 0.046
R409 B.n0 B.t1 512.525
R410 B.n3 B.t4 480.392
R411 B.n3 B.t5 403.272
R412 B.n1 B.t3 372.349
R413 B.n0 B.t0 371.139
R414 B.n1 B.t2 157.328
R415 B.n2 B.n1 132.764
R416 B B.n3 124.329
R417 B.n2 B.n0 93.541
R418 B.n4 B.n2 76
R419 B.n4 B 0.046
R420 a_807_990.n0 a_807_990.t4 477.179
R421 a_807_990.n0 a_807_990.t3 406.485
R422 a_807_990.n4 a_807_990.t5 384.505
R423 a_807_990.n5 a_807_990.n0 228.016
R424 a_807_990.n4 a_807_990.n3 167.985
R425 a_807_990.n6 a_807_990.n5 130.9
R426 a_807_990.n5 a_807_990.n4 79.658
R427 a_807_990.n3 a_807_990.n2 22.578
R428 a_807_990.t1 a_807_990.n6 14.282
R429 a_807_990.n6 a_807_990.t0 14.282
R430 a_807_990.n3 a_807_990.n1 8.58
R431 a_1222_101.n12 a_1222_101.n11 26.811
R432 a_1222_101.n6 a_1222_101.n5 24.977
R433 a_1222_101.n2 a_1222_101.n1 24.877
R434 a_1222_101.t0 a_1222_101.n2 12.677
R435 a_1222_101.t0 a_1222_101.n3 11.595
R436 a_1222_101.t1 a_1222_101.n8 8.137
R437 a_1222_101.t0 a_1222_101.n4 7.273
R438 a_1222_101.t0 a_1222_101.n0 6.109
R439 a_1222_101.t1 a_1222_101.n7 4.864
R440 a_1222_101.t0 a_1222_101.n12 2.074
R441 a_1222_101.n7 a_1222_101.n6 1.13
R442 a_1222_101.n12 a_1222_101.t1 0.937
R443 a_1222_101.t1 a_1222_101.n10 0.804
R444 a_1222_101.n10 a_1222_101.n9 0.136
C6 VDD GND 9.14fF
C7 a_1222_101.n0 GND 0.02fF
C8 a_1222_101.n1 GND 0.10fF
C9 a_1222_101.n2 GND 0.06fF
C10 a_1222_101.n3 GND 0.06fF
C11 a_1222_101.n4 GND 0.00fF
C12 a_1222_101.n5 GND 0.04fF
C13 a_1222_101.n6 GND 0.05fF
C14 a_1222_101.n7 GND 0.02fF
C15 a_1222_101.n8 GND 0.05fF
C16 a_1222_101.n9 GND 0.08fF
C17 a_1222_101.n10 GND 0.17fF
C18 a_1222_101.n11 GND 0.09fF
C19 a_1222_101.n12 GND 0.00fF
C20 a_807_990.n0 GND 1.12fF
C21 a_807_990.n1 GND 0.07fF
C22 a_807_990.n2 GND 0.08fF
C23 a_807_990.n3 GND 0.36fF
C24 a_807_990.n4 GND 1.35fF
C25 a_807_990.n5 GND 1.36fF
C26 a_807_990.n6 GND 1.07fF
C27 Y.n0 GND 1.10fF
C28 Y.n1 GND 0.07fF
C29 Y.n2 GND 0.09fF
C30 Y.n3 GND 0.06fF
C31 Y.n4 GND 0.49fF
C32 Y.n5 GND 0.73fF
C33 Y.n6 GND 1.10fF
C34 Y.n7 GND 0.66fF
C35 Y.n8 GND 0.80fF
C36 Y.n9 GND 0.05fF
C37 a_1241_1051.n0 GND 0.52fF
C38 a_575_1051.n0 GND 0.52fF
C39 VDD.n0 GND 0.12fF
C40 VDD.n1 GND 0.02fF
C41 VDD.n2 GND 0.02fF
C42 VDD.n3 GND 0.04fF
C43 VDD.n4 GND 0.01fF
C44 VDD.n6 GND 0.02fF
C45 VDD.n7 GND 0.02fF
C46 VDD.n8 GND 0.02fF
C47 VDD.n9 GND 0.02fF
C48 VDD.n12 GND 0.02fF
C49 VDD.n14 GND 0.45fF
C50 VDD.n16 GND 0.03fF
C51 VDD.n17 GND 0.02fF
C52 VDD.n18 GND 0.02fF
C53 VDD.n19 GND 0.02fF
C54 VDD.n20 GND 0.03fF
C55 VDD.n21 GND 0.27fF
C56 VDD.n22 GND 0.02fF
C57 VDD.n23 GND 0.03fF
C58 VDD.n24 GND 0.06fF
C59 VDD.n25 GND 0.14fF
C60 VDD.n26 GND 0.20fF
C61 VDD.n27 GND 0.01fF
C62 VDD.n28 GND 0.01fF
C63 VDD.n29 GND 0.07fF
C64 VDD.n30 GND 0.16fF
C65 VDD.n31 GND 0.01fF
C66 VDD.n32 GND 0.02fF
C67 VDD.n33 GND 0.02fF
C68 VDD.n34 GND 0.06fF
C69 VDD.n35 GND 0.14fF
C70 VDD.n36 GND 0.20fF
C71 VDD.n37 GND 0.01fF
C72 VDD.n38 GND 0.01fF
C73 VDD.n39 GND 0.02fF
C74 VDD.n40 GND 0.27fF
C75 VDD.n41 GND 0.01fF
C76 VDD.n42 GND 0.02fF
C77 VDD.n43 GND 0.03fF
C78 VDD.n44 GND 0.02fF
C79 VDD.n45 GND 0.02fF
C80 VDD.n46 GND 0.02fF
C81 VDD.n47 GND 0.18fF
C82 VDD.n48 GND 0.04fF
C83 VDD.n49 GND 0.03fF
C84 VDD.n50 GND 0.02fF
C85 VDD.n52 GND 0.02fF
C86 VDD.n53 GND 0.02fF
C87 VDD.n54 GND 0.02fF
C88 VDD.n55 GND 0.02fF
C89 VDD.n57 GND 0.02fF
C90 VDD.n58 GND 0.02fF
C91 VDD.n59 GND 0.02fF
C92 VDD.n61 GND 0.27fF
C93 VDD.n63 GND 0.02fF
C94 VDD.n64 GND 0.02fF
C95 VDD.n65 GND 0.03fF
C96 VDD.n66 GND 0.02fF
C97 VDD.n67 GND 0.27fF
C98 VDD.n68 GND 0.01fF
C99 VDD.n69 GND 0.02fF
C100 VDD.n70 GND 0.03fF
C101 VDD.n71 GND 0.27fF
C102 VDD.n72 GND 0.01fF
C103 VDD.n73 GND 0.02fF
C104 VDD.n74 GND 0.02fF
C105 VDD.n75 GND 0.27fF
C106 VDD.n76 GND 0.01fF
C107 VDD.n77 GND 0.02fF
C108 VDD.n78 GND 0.02fF
C109 VDD.n79 GND 0.30fF
C110 VDD.n80 GND 0.01fF
C111 VDD.n81 GND 0.03fF
C112 VDD.n82 GND 0.03fF
C113 VDD.n83 GND 0.17fF
C114 VDD.n84 GND 0.14fF
C115 VDD.n85 GND 0.01fF
C116 VDD.n86 GND 0.02fF
C117 VDD.n87 GND 0.03fF
C118 VDD.n88 GND 0.10fF
C119 VDD.n89 GND 0.03fF
C120 VDD.n90 GND 0.13fF
C121 VDD.n91 GND 0.16fF
C122 VDD.n92 GND 0.01fF
C123 VDD.n93 GND 0.02fF
C124 VDD.n94 GND 0.02fF
C125 VDD.n95 GND 0.24fF
C126 VDD.n96 GND 0.01fF
C127 VDD.n97 GND 0.02fF
C128 VDD.n98 GND 0.02fF
C129 VDD.n99 GND 0.02fF
C130 VDD.n100 GND 0.27fF
C131 VDD.n101 GND 0.01fF
C132 VDD.n102 GND 0.02fF
C133 VDD.n103 GND 0.02fF
C134 VDD.n104 GND 0.02fF
C135 VDD.n105 GND 0.21fF
C136 VDD.n106 GND 0.04fF
C137 VDD.n107 GND 0.03fF
C138 VDD.n108 GND 0.02fF
C139 VDD.n109 GND 0.02fF
C140 VDD.n110 GND 0.02fF
C141 VDD.n111 GND 0.02fF
C142 VDD.n112 GND 0.02fF
C143 VDD.n114 GND 0.02fF
C144 VDD.n115 GND 0.02fF
C145 VDD.n116 GND 0.02fF
C146 VDD.n118 GND 0.27fF
C147 VDD.n120 GND 0.02fF
C148 VDD.n121 GND 0.02fF
C149 VDD.n122 GND 0.03fF
C150 VDD.n123 GND 0.02fF
C151 VDD.n124 GND 0.02fF
C152 VDD.n125 GND 0.02fF
C153 VDD.n126 GND 0.02fF
C154 VDD.n127 GND 0.02fF
C155 VDD.n128 GND 0.12fF
C156 VDD.n129 GND 0.03fF
C157 VDD.n130 GND 0.02fF
C158 VDD.n131 GND 0.02fF
C159 VDD.n132 GND 0.02fF
C160 VDD.n133 GND 0.02fF
C161 VDD.n134 GND 0.02fF
C162 VDD.n136 GND 0.02fF
C163 VDD.n137 GND 0.02fF
C164 VDD.n138 GND 0.02fF
C165 VDD.n140 GND 0.45fF
C166 VDD.n142 GND 0.03fF
C167 VDD.n143 GND 0.03fF
C168 VDD.n144 GND 0.27fF
C169 VDD.n145 GND 0.02fF
C170 VDD.n146 GND 0.03fF
C171 VDD.n147 GND 0.03fF
C172 VDD.n148 GND 0.14fF
C173 VDD.n149 GND 0.20fF
C174 VDD.n150 GND 0.01fF
C175 VDD.n151 GND 0.06fF
C176 VDD.n152 GND 0.01fF
C177 VDD.n153 GND 0.02fF
C178 VDD.n154 GND 0.16fF
C179 VDD.n155 GND 0.01fF
C180 VDD.n156 GND 0.02fF
C181 VDD.n157 GND 0.02fF
C182 VDD.n158 GND 0.06fF
C183 VDD.n159 GND 0.14fF
C184 VDD.n160 GND 0.20fF
C185 VDD.n161 GND 0.01fF
C186 VDD.n162 GND 0.01fF
C187 VDD.n163 GND 0.02fF
C188 VDD.n164 GND 0.27fF
C189 VDD.n165 GND 0.01fF
C190 VDD.n166 GND 0.02fF
C191 VDD.n167 GND 0.03fF
C192 VDD.n168 GND 0.02fF
C193 VDD.n169 GND 0.27fF
C194 VDD.n170 GND 0.01fF
C195 VDD.n171 GND 0.02fF
C196 VDD.n172 GND 0.02fF
C197 VDD.n173 GND 0.02fF
C198 VDD.n174 GND 0.02fF
C199 VDD.n175 GND 0.02fF
C200 VDD.n176 GND 0.02fF
C201 VDD.n178 GND 0.02fF
C202 VDD.n179 GND 0.02fF
C203 VDD.n180 GND 0.02fF
C204 VDD.n181 GND 0.02fF
C205 VDD.n183 GND 0.03fF
C206 VDD.n184 GND 0.02fF
C207 VDD.n185 GND 0.18fF
C208 VDD.n186 GND 0.04fF
C209 VDD.n188 GND 0.27fF
C210 VDD.n190 GND 0.02fF
C211 VDD.n191 GND 0.02fF
C212 VDD.n192 GND 0.03fF
C213 VDD.n193 GND 0.02fF
C214 VDD.n194 GND 0.03fF
C215 VDD.n195 GND 0.24fF
C216 VDD.n196 GND 0.01fF
C217 VDD.n197 GND 0.02fF
C218 VDD.n198 GND 0.02fF
C219 VDD.n199 GND 0.10fF
C220 VDD.n200 GND 0.03fF
C221 VDD.n201 GND 0.13fF
C222 VDD.n202 GND 0.16fF
C223 VDD.n203 GND 0.01fF
C224 VDD.n204 GND 0.02fF
C225 VDD.n205 GND 0.02fF
C226 VDD.n206 GND 0.17fF
C227 VDD.n207 GND 0.14fF
C228 VDD.n208 GND 0.01fF
C229 VDD.n209 GND 0.02fF
C230 VDD.n210 GND 0.03fF
C231 VDD.n211 GND 0.30fF
C232 VDD.n212 GND 0.01fF
C233 VDD.n213 GND 0.03fF
C234 VDD.n214 GND 0.03fF
C235 VDD.n215 GND 0.27fF
C236 VDD.n216 GND 0.01fF
C237 VDD.n217 GND 0.02fF
C238 VDD.n218 GND 0.02fF
C239 VDD.n219 GND 0.27fF
C240 VDD.n220 GND 0.01fF
C241 VDD.n221 GND 0.02fF
C242 VDD.n222 GND 0.02fF
C243 VDD.n223 GND 0.27fF
C244 VDD.n224 GND 0.01fF
C245 VDD.n225 GND 0.02fF
C246 VDD.n226 GND 0.02fF
C247 a_556_101.n0 GND 0.05fF
C248 a_556_101.n1 GND 0.12fF
C249 a_556_101.n2 GND 0.04fF
C250 a_185_209.n0 GND 0.99fF
C251 a_185_209.n1 GND 0.53fF
C252 a_185_209.n2 GND 1.23fF
C253 a_185_209.n3 GND 1.29fF
C254 a_185_209.n4 GND 0.11fF
C255 a_185_209.n5 GND 0.32fF
C256 a_185_209.n6 GND 0.06fF
.ends
