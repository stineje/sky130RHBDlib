* SPICE3 file created from AO3X1.ext - technology: sky130A

.subckt AO3X1 A B C Y VDD VSS
X0 VDD A a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0.00336 pd=2.736 as=0 ps=0 w=2 l=0.15 M=2
X1 VDD a_217_1050 a_797_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X2 VDD a_864_209 Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.0058 ps=4.58 w=2 l=0.15 M=2
X3 VDD B a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X4 a_797_1051 C a_864_209 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X5 VSS A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0.0032565 pd=2.261 as=0 ps=0 w=3 l=0.15
X6 a_864_209 a_217_1050 VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X7 a_217_1050 B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X8 a_864_209 C VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X9 Y a_864_209 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
C0 a_217_1050 VDD 2.17f
C1 VDD VSS 3.28f
.ends
