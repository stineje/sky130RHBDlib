* SPICE3 file created from TMRDFFSNRNQX1.ext - technology: sky130A

.subckt TMRDFFSNRNQX1 Q D CLK SN RN VDD GND
M1000 VDD.t60 a_10219_989.t7 a_17533_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_15669_1050.t4 a_15991_989.t7 VDD.t65 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 GND a_6049_1050.t8 a_7787_103.t0 nshort w=-1.605u l=1.765u
+  ad=4.9019p pd=41.07u as=0p ps=0u
M1003 VDD.t42 a_11821_1050.t7 a_12143_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_13105_989.t0 CLK.t1 VDD.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 GND a_6371_989.t8 a_9711_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1006 VDD.t94 SN.t0 a_15991_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 GND D.t4 a_5863_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t77 SN.t1 a_10219_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_13745_1050.t3 a_11821_1050.t8 VDD.t43 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VDD.t35 a_12143_989.t7 a_15669_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_6049_1050.t1 a_6371_989.t7 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VDD.t69 a_2201_1050.t7 a_1561_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VDD.t49 a_7333_989.t7 a_7973_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t61 a_10219_989.t8 a_9897_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_4447_989.t3 SN.t2 VDD.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_17708_209.t2 a_4447_989.t8 a_18197_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_17533_1051.t7 a_4447_989.t9 a_18197_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VDD.t19 CLK.t2 a_6371_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_7333_989.t4 RN.t0 VDD.t106 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 GND a_11821_1050.t9 a_12597_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t54 D.t1 a_6049_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 GND a_13745_1050.t7 a_14521_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_7973_1050.t4 SN.t4 VDD.t78 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_18197_1051.t4 a_10219_989.t9 a_17708_209.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 VDD.t38 a_15991_989.t9 a_17533_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 GND a_9897_1050.t7 a_10673_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1027 GND a_7973_1050.t7 a_8749_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1028 VDD.t68 D.t2 a_277_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q a_17708_209.t7 GND.t15 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1030 VDD.t86 D.t3 a_11821_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 GND D.t5 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1032 VDD.t85 RN.t2 a_15669_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_599_989.t3 CLK.t3 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VDD.t105 RN.t3 a_9897_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_11821_1050.t1 a_12143_989.t8 VDD.t36 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 VDD.t10 CLK.t4 a_1561_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VDD.t33 a_13105_989.t9 a_13745_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 GND a_15991_989.t11 a_17428_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1039 VDD.t102 a_277_1050.t7 a_2201_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_7333_989.t1 CLK.t6 VDD.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_10219_989.t0 SN.t5 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VDD.t75 a_7333_989.t8 a_6371_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 VDD.t16 CLK.t7 a_12143_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_13105_989.t3 RN.t4 VDD.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 GND a_11821_1050.t10 a_13559_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1046 GND a_12143_989.t9 a_15483_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1047 VDD.t80 RN.t5 a_277_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_6371_989.t4 a_6049_1050.t9 VDD.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_17533_1051.t4 a_15991_989.t10 VDD.t39 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 VDD.t109 a_7973_1050.t8 a_7333_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 VDD.t93 a_9897_1050.t8 a_10219_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 a_12143_989.t0 CLK.t8 VDD.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_599_989.t6 a_1561_989.t7 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_15991_989.t0 a_15669_1050.t7 VDD.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 VDD.t104 RN.t7 a_1561_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_9897_1050.t2 a_6371_989.t9 VDD.t88 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 GND a_15669_1050.t8 a_16445_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_4125_1050.t3 a_599_989.t8 VDD.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 VDD.t112 SN.t6 a_2201_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 a_4125_1050.t2 a_4447_989.t10 VDD.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 VDD.t72 a_6371_989.t10 a_6049_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_18197_1051.t7 a_15991_989.t12 a_17533_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_1561_989.t0 CLK.t9 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 VDD.t81 a_599_989.t9 a_277_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 a_13745_1050.t4 SN.t7 VDD.t51 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_17533_1051.t5 a_10219_989.t11 VDD.t59 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_12143_989.t2 a_11821_1050.t11 VDD.t98 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 VDD.t47 a_13745_1050.t8 a_13105_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_15991_989.t6 SN.t10 VDD.t97 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 VDD.t100 a_17708_209.t8 Q.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_15669_1050.t6 a_12143_989.t10 VDD.t108 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_4125_1050.t5 RN.t9 VDD.t79 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 GND a_277_1050.t8 a_2015_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1074 VDD.t73 a_1561_989.t8 a_2201_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 VDD.t84 RN.t10 a_6049_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 a_7333_989.t6 a_7973_1050.t9 VDD.t113 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 a_7973_1050.t0 a_7333_989.t9 VDD.t70 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 a_9897_1050.t4 a_10219_989.t12 VDD.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VDD.t34 a_13105_989.t10 a_15991_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_1561_989.t3 a_2201_1050.t8 VDD.t50 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 a_18197_1051.t0 a_4447_989.t13 a_17533_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 VDD.t1 a_4125_1050.t8 a_4447_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_6371_989.t0 CLK.t12 VDD.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 VDD.t20 CLK.t13 a_7333_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_6049_1050.t0 D.t6 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_17708_209.t3 a_10219_989.t13 a_18197_1051.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 a_277_1050.t0 D.t7 VDD.t89 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 VDD.t13 CLK.t14 a_13105_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_15991_989.t1 a_13105_989.t11 VDD.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 a_10219_989.t2 a_7333_989.t10 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 VDD.t99 a_11821_1050.t12 a_13745_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 VDD.t30 a_13105_989.t12 a_12143_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_15669_1050.t0 RN.t13 VDD.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 GND a_2201_1050.t9 a_2977_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1095 VDD.t64 a_277_1050.t9 a_599_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 a_9897_1050.t0 RN.t14 VDD.t48 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 VDD.t7 RN.t15 a_11821_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 VDD.t74 a_1561_989.t11 a_599_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 a_13745_1050.t1 a_13105_989.t13 VDD.t32 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 GND a_277_1050.t10 a_1053_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1101 VDD.t91 SN.t12 a_4447_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_18197_1051.t3 a_4447_989.t14 a_17708_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 VDD.t37 a_15991_989.t13 a_15669_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_6371_989.t2 a_7333_989.t12 VDD.t53 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 VDD.t67 RN.t17 a_7333_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VDD.t82 SN.t13 a_7973_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 a_277_1050.t5 RN.t18 VDD.t40 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 a_11821_1050.t3 RN.t19 VDD.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 VDD.t76 SN.t14 a_13745_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_10219_989.t5 a_9897_1050.t9 VDD.t92 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 GND a_599_989.t11 a_3939_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1112 VDD.t11 CLK.t15 a_599_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 a_1561_989.t5 RN.t20 VDD.t103 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1114 VDD.t107 a_12143_989.t12 a_11821_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 VDD.t111 a_1561_989.t13 a_4447_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 a_2201_1050.t2 SN.t15 VDD.t96 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_12143_989.t5 a_13105_989.t14 VDD.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 VDD.t6 RN.t21 a_4125_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 VDD.t22 RN.t22 a_13105_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 a_599_989.t0 a_277_1050.t11 VDD.t101 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 VDD.t58 a_6049_1050.t10 a_7973_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 a_277_1050.t4 a_599_989.t10 VDD.t87 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 a_11821_1050.t2 D.t8 VDD.t52 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1124 GND a_6049_1050.t7 a_6825_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1125 a_13105_989.t6 a_13745_1050.t9 VDD.t46 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1126 GND a_4125_1050.t7 a_4901_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1127 VDD.t41 a_15669_1050.t9 a_15991_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1128 a_7973_1050.t5 a_6049_1050.t11 VDD.t57 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1129 VDD.t110 a_6371_989.t12 a_9897_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1130 a_2201_1050.t1 a_277_1050.t12 VDD.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1131 VDD.t4 a_7333_989.t15 a_10219_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1132 Q.t1 a_17708_209.t9 VDD.t26 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1133 a_2201_1050.t5 a_1561_989.t14 VDD.t90 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1134 VDD.t44 a_599_989.t12 a_4125_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1135 a_6049_1050.t3 RN.t26 VDD.t63 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1136 GND a_4447_989.t7 a_18760_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1137 GND a_15991_989.t8 a_18094_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1138 VDD.t95 a_4447_989.t15 a_4125_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1139 a_17533_1051.t2 a_15991_989.t14 a_18197_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1140 a_4447_989.t0 a_4125_1050.t9 VDD.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1141 VDD.t55 a_6049_1050.t12 a_6371_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1142 a_4447_989.t4 a_1561_989.t15 VDD.t83 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1143 GND D.t0 a_11635_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD SN 0.30fF
C1 VDD Q 0.76fF
C2 D SN 0.31fF
C3 RN SN 16.07fF
C4 CLK SN 0.63fF
C5 VDD D 5.87fF
C6 VDD RN 0.48fF
C7 VDD CLK 1.65fF
C8 D RN 2.36fF
C9 D CLK 12.06fF
C10 RN CLK 1.11fF
R0 CLK.n18 CLK.t15 459.505
R1 CLK.n15 CLK.t4 459.505
R2 CLK.n12 CLK.t2 459.505
R3 CLK.n7 CLK.t13 459.505
R4 CLK.n4 CLK.t7 459.505
R5 CLK.n0 CLK.t14 459.505
R6 CLK.n18 CLK.t3 384.527
R7 CLK.n15 CLK.t9 384.527
R8 CLK.n12 CLK.t12 384.527
R9 CLK.n7 CLK.t6 384.527
R10 CLK.n4 CLK.t8 384.527
R11 CLK.n0 CLK.t1 384.527
R12 CLK.n16 CLK.t0 322.151
R13 CLK.n8 CLK.t5 322.151
R14 CLK.n1 CLK.t10 322.151
R15 CLK.n20 CLK.t17 321.792
R16 CLK.n10 CLK.t16 320.152
R17 CLK.n2 CLK.t11 320.152
R18 CLK.n19 CLK 152
R19 CLK.n6 CLK.n5 75.989
R20 CLK.n14 CLK.n13 75.989
R21 CLK.n3 CLK.n2 75.568
R22 CLK.n11 CLK.n10 75.568
R23 CLK.n3 CLK.n1 56.374
R24 CLK.n21 CLK.n20 49.379
R25 CLK.n9 CLK.n8 49.342
R26 CLK.n17 CLK.n16 49.342
R27 CLK.n1 CLK.n0 27.599
R28 CLK.n8 CLK.n7 27.599
R29 CLK.n16 CLK.n15 27.599
R30 CLK.n19 CLK.n18 21.475
R31 CLK.n13 CLK.n12 21.475
R32 CLK.n5 CLK.n4 21.475
R33 CLK.n9 CLK.n6 14.076
R34 CLK.n17 CLK.n14 14.076
R35 CLK.n11 CLK.n9 7.032
R36 CLK.n21 CLK.n17 7.032
R37 CLK.n20 CLK.n19 3.3
R38 CLK.n21 CLK 0.046
R39 CLK.n6 CLK.n3 0.023
R40 CLK.n14 CLK.n11 0.023
R41 a_2977_103.t0 a_2977_103.n0 117.777
R42 a_2977_103.n2 a_2977_103.n1 55.228
R43 a_2977_103.n4 a_2977_103.n3 9.111
R44 a_2977_103.n8 a_2977_103.n6 7.859
R45 a_2977_103.t0 a_2977_103.n2 4.04
R46 a_2977_103.t0 a_2977_103.n8 3.034
R47 a_2977_103.n6 a_2977_103.n4 1.964
R48 a_2977_103.n6 a_2977_103.n5 1.964
R49 a_2977_103.n8 a_2977_103.n7 0.443
R50 a_3258_210.n12 a_3258_210.n10 82.852
R51 a_3258_210.n13 a_3258_210.n0 49.6
R52 a_3258_210.t1 a_3258_210.n2 46.91
R53 a_3258_210.n7 a_3258_210.n5 34.805
R54 a_3258_210.n7 a_3258_210.n6 32.622
R55 a_3258_210.n10 a_3258_210.t1 32.416
R56 a_3258_210.n12 a_3258_210.n11 27.2
R57 a_3258_210.n13 a_3258_210.n12 22.4
R58 a_3258_210.n9 a_3258_210.n7 19.017
R59 a_3258_210.n2 a_3258_210.n1 17.006
R60 a_3258_210.n5 a_3258_210.n4 7.5
R61 a_3258_210.n9 a_3258_210.n8 7.5
R62 a_3258_210.t1 a_3258_210.n3 7.04
R63 a_3258_210.n10 a_3258_210.n9 1.435
R64 a_13105_989.n7 a_13105_989.t13 454.685
R65 a_13105_989.n9 a_13105_989.t14 454.685
R66 a_13105_989.n5 a_13105_989.t11 454.685
R67 a_13105_989.n7 a_13105_989.t9 428.979
R68 a_13105_989.n9 a_13105_989.t12 428.979
R69 a_13105_989.n5 a_13105_989.t10 428.979
R70 a_13105_989.n8 a_13105_989.t7 264.512
R71 a_13105_989.n6 a_13105_989.t8 264.512
R72 a_13105_989.n10 a_13105_989.t15 264.173
R73 a_13105_989.n15 a_13105_989.n13 246.179
R74 a_13105_989.n13 a_13105_989.n4 144.246
R75 a_13105_989.n12 a_13105_989.n6 82.484
R76 a_13105_989.n11 a_13105_989.n10 79.495
R77 a_13105_989.n3 a_13105_989.n2 79.232
R78 a_13105_989.n11 a_13105_989.n8 76
R79 a_13105_989.n13 a_13105_989.n12 76
R80 a_13105_989.n8 a_13105_989.n7 71.894
R81 a_13105_989.n6 a_13105_989.n5 71.894
R82 a_13105_989.n10 a_13105_989.n9 71.555
R83 a_13105_989.n4 a_13105_989.n3 63.152
R84 a_13105_989.n4 a_13105_989.n0 16.08
R85 a_13105_989.n3 a_13105_989.n1 16.08
R86 a_13105_989.n15 a_13105_989.n14 15.218
R87 a_13105_989.n0 a_13105_989.t2 14.282
R88 a_13105_989.n0 a_13105_989.t3 14.282
R89 a_13105_989.n1 a_13105_989.t1 14.282
R90 a_13105_989.n1 a_13105_989.t0 14.282
R91 a_13105_989.n2 a_13105_989.t4 14.282
R92 a_13105_989.n2 a_13105_989.t6 14.282
R93 a_13105_989.n16 a_13105_989.n15 12.014
R94 a_13105_989.n12 a_13105_989.n11 4.035
R95 a_13840_210.n12 a_13840_210.n5 96.467
R96 a_13840_210.t0 a_13840_210.n1 46.91
R97 a_13840_210.n9 a_13840_210.n7 34.805
R98 a_13840_210.n9 a_13840_210.n8 32.622
R99 a_13840_210.t0 a_13840_210.n12 32.417
R100 a_13840_210.n5 a_13840_210.n4 22.349
R101 a_13840_210.n11 a_13840_210.n9 19.017
R102 a_13840_210.n1 a_13840_210.n0 17.006
R103 a_13840_210.n5 a_13840_210.n3 8.443
R104 a_13840_210.t0 a_13840_210.n2 8.137
R105 a_13840_210.n7 a_13840_210.n6 7.5
R106 a_13840_210.n11 a_13840_210.n10 7.5
R107 a_13840_210.n12 a_13840_210.n11 1.435
R108 a_13745_1050.n5 a_13745_1050.t8 512.525
R109 a_13745_1050.n5 a_13745_1050.t9 371.139
R110 a_13745_1050.n6 a_13745_1050.t7 234.562
R111 a_13745_1050.n7 a_13745_1050.n4 223.905
R112 a_13745_1050.n6 a_13745_1050.n5 215.819
R113 a_13745_1050.n9 a_13745_1050.n7 166.52
R114 a_13745_1050.n7 a_13745_1050.n6 153.315
R115 a_13745_1050.n3 a_13745_1050.n2 79.232
R116 a_13745_1050.n4 a_13745_1050.n3 63.152
R117 a_13745_1050.n4 a_13745_1050.n0 16.08
R118 a_13745_1050.n3 a_13745_1050.n1 16.08
R119 a_13745_1050.n9 a_13745_1050.n8 15.218
R120 a_13745_1050.n0 a_13745_1050.t2 14.282
R121 a_13745_1050.n0 a_13745_1050.t1 14.282
R122 a_13745_1050.n1 a_13745_1050.t5 14.282
R123 a_13745_1050.n1 a_13745_1050.t4 14.282
R124 a_13745_1050.n2 a_13745_1050.t6 14.282
R125 a_13745_1050.n2 a_13745_1050.t3 14.282
R126 a_13745_1050.n10 a_13745_1050.n9 12.014
R127 a_6049_1050.n7 a_6049_1050.t12 512.525
R128 a_6049_1050.n5 a_6049_1050.t10 512.525
R129 a_6049_1050.n7 a_6049_1050.t9 371.139
R130 a_6049_1050.n5 a_6049_1050.t11 371.139
R131 a_6049_1050.n8 a_6049_1050.t7 234.921
R132 a_6049_1050.n6 a_6049_1050.t8 234.921
R133 a_6049_1050.n10 a_6049_1050.n4 223.546
R134 a_6049_1050.n8 a_6049_1050.n7 215.46
R135 a_6049_1050.n6 a_6049_1050.n5 215.46
R136 a_6049_1050.n12 a_6049_1050.n10 166.879
R137 a_6049_1050.n9 a_6049_1050.n6 79.491
R138 a_6049_1050.n3 a_6049_1050.n2 79.232
R139 a_6049_1050.n10 a_6049_1050.n9 77.315
R140 a_6049_1050.n9 a_6049_1050.n8 76
R141 a_6049_1050.n4 a_6049_1050.n3 63.152
R142 a_6049_1050.n4 a_6049_1050.n0 16.08
R143 a_6049_1050.n3 a_6049_1050.n1 16.08
R144 a_6049_1050.n12 a_6049_1050.n11 15.218
R145 a_6049_1050.n0 a_6049_1050.t4 14.282
R146 a_6049_1050.n0 a_6049_1050.t1 14.282
R147 a_6049_1050.n1 a_6049_1050.t6 14.282
R148 a_6049_1050.n1 a_6049_1050.t3 14.282
R149 a_6049_1050.n2 a_6049_1050.t2 14.282
R150 a_6049_1050.n2 a_6049_1050.t0 14.282
R151 a_6049_1050.n13 a_6049_1050.n12 12.014
R152 a_6825_103.t0 a_6825_103.n0 117.777
R153 a_6825_103.n2 a_6825_103.n1 55.228
R154 a_6825_103.n4 a_6825_103.n3 9.111
R155 a_6825_103.n8 a_6825_103.n6 7.859
R156 a_6825_103.t0 a_6825_103.n2 4.04
R157 a_6825_103.t0 a_6825_103.n8 3.034
R158 a_6825_103.n6 a_6825_103.n4 1.964
R159 a_6825_103.n6 a_6825_103.n5 1.964
R160 a_6825_103.n8 a_6825_103.n7 0.443
R161 GND.n30 GND.n29 219.745
R162 GND.n60 GND.n58 219.745
R163 GND.n90 GND.n88 219.745
R164 GND.n487 GND.n486 219.745
R165 GND.n529 GND.n527 219.745
R166 GND.n571 GND.n569 219.745
R167 GND.n613 GND.n611 219.745
R168 GND.n655 GND.n653 219.745
R169 GND.n697 GND.n695 219.745
R170 GND.n742 GND.n740 219.745
R171 GND.n784 GND.n782 219.745
R172 GND.n829 GND.n827 219.745
R173 GND.n871 GND.n869 219.745
R174 GND.n417 GND.n415 219.745
R175 GND.n375 GND.n373 219.745
R176 GND.n333 GND.n331 219.745
R177 GND.n291 GND.n289 219.745
R178 GND.n249 GND.n247 219.745
R179 GND.n204 GND.n202 219.745
R180 GND.n162 GND.n160 219.745
R181 GND.n120 GND.n119 219.745
R182 GND.n151 GND.n150 85.559
R183 GND.n193 GND.n192 85.559
R184 GND.n280 GND.n279 85.559
R185 GND.n322 GND.n321 85.559
R186 GND.n364 GND.n363 85.559
R187 GND.n406 GND.n405 85.559
R188 GND.n880 GND.n879 85.559
R189 GND.n838 GND.n837 85.559
R190 GND.n751 GND.n750 85.559
R191 GND.n664 GND.n663 85.559
R192 GND.n622 GND.n621 85.559
R193 GND.n580 GND.n579 85.559
R194 GND.n538 GND.n537 85.559
R195 GND.n496 GND.n495 85.559
R196 GND.n454 GND.n453 85.559
R197 GND.n30 GND.n28 85.529
R198 GND.n60 GND.n59 85.529
R199 GND.n90 GND.n89 85.529
R200 GND.n487 GND.n485 85.529
R201 GND.n529 GND.n528 85.529
R202 GND.n571 GND.n570 85.529
R203 GND.n613 GND.n612 85.529
R204 GND.n655 GND.n654 85.529
R205 GND.n697 GND.n696 85.529
R206 GND.n742 GND.n741 85.529
R207 GND.n784 GND.n783 85.529
R208 GND.n829 GND.n828 85.529
R209 GND.n871 GND.n870 85.529
R210 GND.n417 GND.n416 85.529
R211 GND.n375 GND.n374 85.529
R212 GND.n333 GND.n332 85.529
R213 GND.n291 GND.n290 85.529
R214 GND.n249 GND.n248 85.529
R215 GND.n204 GND.n203 85.529
R216 GND.n162 GND.n161 85.529
R217 GND.n120 GND.n118 85.529
R218 GND.n78 GND.n77 84.842
R219 GND.n108 GND.n107 84.842
R220 GND.n48 GND.n47 84.842
R221 GND.n9 GND.n1 76.145
R222 GND.n448 GND.n447 76
R223 GND.n73 GND.n72 76
R224 GND.n76 GND.n75 76
R225 GND.n81 GND.n80 76
R226 GND.n84 GND.n83 76
R227 GND.n87 GND.n86 76
R228 GND.n94 GND.n93 76
R229 GND.n97 GND.n96 76
R230 GND.n100 GND.n99 76
R231 GND.n103 GND.n102 76
R232 GND.n106 GND.n105 76
R233 GND.n111 GND.n110 76
R234 GND.n114 GND.n113 76
R235 GND.n117 GND.n116 76
R236 GND.n124 GND.n123 76
R237 GND.n127 GND.n126 76
R238 GND.n130 GND.n129 76
R239 GND.n133 GND.n132 76
R240 GND.n136 GND.n135 76
R241 GND.n139 GND.n138 76
R242 GND.n142 GND.n141 76
R243 GND.n145 GND.n144 76
R244 GND.n148 GND.n147 76
R245 GND.n153 GND.n152 76
R246 GND.n156 GND.n155 76
R247 GND.n159 GND.n158 76
R248 GND.n166 GND.n165 76
R249 GND.n169 GND.n168 76
R250 GND.n172 GND.n171 76
R251 GND.n175 GND.n174 76
R252 GND.n178 GND.n177 76
R253 GND.n181 GND.n180 76
R254 GND.n184 GND.n183 76
R255 GND.n187 GND.n186 76
R256 GND.n190 GND.n189 76
R257 GND.n195 GND.n194 76
R258 GND.n198 GND.n197 76
R259 GND.n201 GND.n200 76
R260 GND.n208 GND.n207 76
R261 GND.n211 GND.n210 76
R262 GND.n214 GND.n213 76
R263 GND.n217 GND.n216 76
R264 GND.n220 GND.n219 76
R265 GND.n223 GND.n222 76
R266 GND.n226 GND.n225 76
R267 GND.n229 GND.n228 76
R268 GND.n232 GND.n231 76
R269 GND.n240 GND.n239 76
R270 GND.n243 GND.n242 76
R271 GND.n246 GND.n245 76
R272 GND.n253 GND.n252 76
R273 GND.n256 GND.n255 76
R274 GND.n259 GND.n258 76
R275 GND.n262 GND.n261 76
R276 GND.n265 GND.n264 76
R277 GND.n268 GND.n267 76
R278 GND.n271 GND.n270 76
R279 GND.n274 GND.n273 76
R280 GND.n277 GND.n276 76
R281 GND.n282 GND.n281 76
R282 GND.n285 GND.n284 76
R283 GND.n288 GND.n287 76
R284 GND.n295 GND.n294 76
R285 GND.n298 GND.n297 76
R286 GND.n301 GND.n300 76
R287 GND.n304 GND.n303 76
R288 GND.n307 GND.n306 76
R289 GND.n310 GND.n309 76
R290 GND.n313 GND.n312 76
R291 GND.n316 GND.n315 76
R292 GND.n319 GND.n318 76
R293 GND.n324 GND.n323 76
R294 GND.n327 GND.n326 76
R295 GND.n330 GND.n329 76
R296 GND.n337 GND.n336 76
R297 GND.n340 GND.n339 76
R298 GND.n343 GND.n342 76
R299 GND.n346 GND.n345 76
R300 GND.n349 GND.n348 76
R301 GND.n352 GND.n351 76
R302 GND.n355 GND.n354 76
R303 GND.n358 GND.n357 76
R304 GND.n361 GND.n360 76
R305 GND.n366 GND.n365 76
R306 GND.n369 GND.n368 76
R307 GND.n372 GND.n371 76
R308 GND.n379 GND.n378 76
R309 GND.n382 GND.n381 76
R310 GND.n385 GND.n384 76
R311 GND.n388 GND.n387 76
R312 GND.n391 GND.n390 76
R313 GND.n394 GND.n393 76
R314 GND.n397 GND.n396 76
R315 GND.n400 GND.n399 76
R316 GND.n403 GND.n402 76
R317 GND.n408 GND.n407 76
R318 GND.n411 GND.n410 76
R319 GND.n414 GND.n413 76
R320 GND.n421 GND.n420 76
R321 GND.n424 GND.n423 76
R322 GND.n427 GND.n426 76
R323 GND.n430 GND.n429 76
R324 GND.n433 GND.n432 76
R325 GND.n436 GND.n435 76
R326 GND.n439 GND.n438 76
R327 GND.n442 GND.n441 76
R328 GND.n445 GND.n444 76
R329 GND.n882 GND.n881 76
R330 GND.n877 GND.n876 76
R331 GND.n874 GND.n873 76
R332 GND.n867 GND.n866 76
R333 GND.n864 GND.n863 76
R334 GND.n861 GND.n860 76
R335 GND.n858 GND.n857 76
R336 GND.n855 GND.n854 76
R337 GND.n852 GND.n851 76
R338 GND.n849 GND.n848 76
R339 GND.n846 GND.n845 76
R340 GND.n843 GND.n842 76
R341 GND.n840 GND.n839 76
R342 GND.n835 GND.n834 76
R343 GND.n832 GND.n831 76
R344 GND.n825 GND.n824 76
R345 GND.n822 GND.n821 76
R346 GND.n819 GND.n818 76
R347 GND.n816 GND.n815 76
R348 GND.n813 GND.n812 76
R349 GND.n810 GND.n809 76
R350 GND.n807 GND.n806 76
R351 GND.n804 GND.n803 76
R352 GND.n801 GND.n800 76
R353 GND.n798 GND.n797 76
R354 GND.n790 GND.n789 76
R355 GND.n787 GND.n786 76
R356 GND.n780 GND.n779 76
R357 GND.n777 GND.n776 76
R358 GND.n774 GND.n773 76
R359 GND.n771 GND.n770 76
R360 GND.n768 GND.n767 76
R361 GND.n765 GND.n764 76
R362 GND.n762 GND.n761 76
R363 GND.n759 GND.n758 76
R364 GND.n756 GND.n755 76
R365 GND.n753 GND.n752 76
R366 GND.n748 GND.n747 76
R367 GND.n745 GND.n744 76
R368 GND.n738 GND.n737 76
R369 GND.n735 GND.n734 76
R370 GND.n732 GND.n731 76
R371 GND.n729 GND.n728 76
R372 GND.n726 GND.n725 76
R373 GND.n723 GND.n722 76
R374 GND.n720 GND.n719 76
R375 GND.n717 GND.n716 76
R376 GND.n714 GND.n713 76
R377 GND.n711 GND.n710 76
R378 GND.n703 GND.n702 76
R379 GND.n700 GND.n699 76
R380 GND.n693 GND.n692 76
R381 GND.n690 GND.n689 76
R382 GND.n687 GND.n686 76
R383 GND.n684 GND.n683 76
R384 GND.n681 GND.n680 76
R385 GND.n678 GND.n677 76
R386 GND.n675 GND.n674 76
R387 GND.n672 GND.n671 76
R388 GND.n669 GND.n668 76
R389 GND.n666 GND.n665 76
R390 GND.n661 GND.n660 76
R391 GND.n658 GND.n657 76
R392 GND.n651 GND.n650 76
R393 GND.n648 GND.n647 76
R394 GND.n645 GND.n644 76
R395 GND.n642 GND.n641 76
R396 GND.n639 GND.n638 76
R397 GND.n636 GND.n635 76
R398 GND.n633 GND.n632 76
R399 GND.n630 GND.n629 76
R400 GND.n627 GND.n626 76
R401 GND.n624 GND.n623 76
R402 GND.n619 GND.n618 76
R403 GND.n616 GND.n615 76
R404 GND.n609 GND.n608 76
R405 GND.n606 GND.n605 76
R406 GND.n603 GND.n602 76
R407 GND.n600 GND.n599 76
R408 GND.n597 GND.n596 76
R409 GND.n594 GND.n593 76
R410 GND.n591 GND.n590 76
R411 GND.n588 GND.n587 76
R412 GND.n585 GND.n584 76
R413 GND.n582 GND.n581 76
R414 GND.n577 GND.n576 76
R415 GND.n574 GND.n573 76
R416 GND.n567 GND.n566 76
R417 GND.n564 GND.n563 76
R418 GND.n561 GND.n560 76
R419 GND.n558 GND.n557 76
R420 GND.n555 GND.n554 76
R421 GND.n552 GND.n551 76
R422 GND.n549 GND.n548 76
R423 GND.n546 GND.n545 76
R424 GND.n543 GND.n542 76
R425 GND.n540 GND.n539 76
R426 GND.n535 GND.n534 76
R427 GND.n532 GND.n531 76
R428 GND.n525 GND.n524 76
R429 GND.n522 GND.n521 76
R430 GND.n519 GND.n518 76
R431 GND.n516 GND.n515 76
R432 GND.n513 GND.n512 76
R433 GND.n510 GND.n509 76
R434 GND.n507 GND.n506 76
R435 GND.n504 GND.n503 76
R436 GND.n501 GND.n500 76
R437 GND.n498 GND.n497 76
R438 GND.n493 GND.n492 76
R439 GND.n490 GND.n489 76
R440 GND.n483 GND.n482 76
R441 GND.n480 GND.n479 76
R442 GND.n477 GND.n476 76
R443 GND.n474 GND.n473 76
R444 GND.n471 GND.n470 76
R445 GND.n468 GND.n467 76
R446 GND.n465 GND.n464 76
R447 GND.n462 GND.n461 76
R448 GND.n459 GND.n458 76
R449 GND.n456 GND.n455 76
R450 GND.n451 GND.n450 76
R451 GND.n9 GND.n8 76
R452 GND.n17 GND.n16 76
R453 GND.n24 GND.n23 76
R454 GND.n27 GND.n26 76
R455 GND.n34 GND.n33 76
R456 GND.n37 GND.n36 76
R457 GND.n40 GND.n39 76
R458 GND.n43 GND.n42 76
R459 GND.n46 GND.n45 76
R460 GND.n51 GND.n50 76
R461 GND.n54 GND.n53 76
R462 GND.n57 GND.n56 76
R463 GND.n64 GND.n63 76
R464 GND.n67 GND.n66 76
R465 GND.n70 GND.n69 76
R466 GND.n238 GND.n237 64.552
R467 GND.n796 GND.n795 64.552
R468 GND.n709 GND.n708 64.552
R469 GND.n5 GND.n4 35.01
R470 GND.n3 GND.n2 29.127
R471 GND.n237 GND.n236 28.421
R472 GND.n795 GND.n794 28.421
R473 GND.n708 GND.n707 28.421
R474 GND.n237 GND.n235 25.263
R475 GND.n795 GND.n793 25.263
R476 GND.n708 GND.n706 25.263
R477 GND.n235 GND.n234 24.383
R478 GND.n793 GND.n792 24.383
R479 GND.n706 GND.n705 24.383
R480 GND.n12 GND.t15 20.794
R481 GND.n6 GND.n5 19.735
R482 GND.n14 GND.n13 19.735
R483 GND.n21 GND.n20 19.735
R484 GND.n5 GND.n3 19.017
R485 GND.n33 GND.n31 14.167
R486 GND.n63 GND.n61 14.167
R487 GND.n93 GND.n91 14.167
R488 GND.n123 GND.n121 14.167
R489 GND.n165 GND.n163 14.167
R490 GND.n207 GND.n205 14.167
R491 GND.n252 GND.n250 14.167
R492 GND.n294 GND.n292 14.167
R493 GND.n336 GND.n334 14.167
R494 GND.n378 GND.n376 14.167
R495 GND.n420 GND.n418 14.167
R496 GND.n873 GND.n872 14.167
R497 GND.n831 GND.n830 14.167
R498 GND.n786 GND.n785 14.167
R499 GND.n744 GND.n743 14.167
R500 GND.n699 GND.n698 14.167
R501 GND.n657 GND.n656 14.167
R502 GND.n615 GND.n614 14.167
R503 GND.n573 GND.n572 14.167
R504 GND.n531 GND.n530 14.167
R505 GND.n489 GND.n488 14.167
R506 GND.n450 GND.n449 13.653
R507 GND.n455 GND.n452 13.653
R508 GND.n458 GND.n457 13.653
R509 GND.n461 GND.n460 13.653
R510 GND.n464 GND.n463 13.653
R511 GND.n467 GND.n466 13.653
R512 GND.n470 GND.n469 13.653
R513 GND.n473 GND.n472 13.653
R514 GND.n476 GND.n475 13.653
R515 GND.n479 GND.n478 13.653
R516 GND.n482 GND.n481 13.653
R517 GND.n489 GND.n484 13.653
R518 GND.n492 GND.n491 13.653
R519 GND.n497 GND.n494 13.653
R520 GND.n500 GND.n499 13.653
R521 GND.n503 GND.n502 13.653
R522 GND.n506 GND.n505 13.653
R523 GND.n509 GND.n508 13.653
R524 GND.n512 GND.n511 13.653
R525 GND.n515 GND.n514 13.653
R526 GND.n518 GND.n517 13.653
R527 GND.n521 GND.n520 13.653
R528 GND.n524 GND.n523 13.653
R529 GND.n531 GND.n526 13.653
R530 GND.n534 GND.n533 13.653
R531 GND.n539 GND.n536 13.653
R532 GND.n542 GND.n541 13.653
R533 GND.n545 GND.n544 13.653
R534 GND.n548 GND.n547 13.653
R535 GND.n551 GND.n550 13.653
R536 GND.n554 GND.n553 13.653
R537 GND.n557 GND.n556 13.653
R538 GND.n560 GND.n559 13.653
R539 GND.n563 GND.n562 13.653
R540 GND.n566 GND.n565 13.653
R541 GND.n573 GND.n568 13.653
R542 GND.n576 GND.n575 13.653
R543 GND.n581 GND.n578 13.653
R544 GND.n584 GND.n583 13.653
R545 GND.n587 GND.n586 13.653
R546 GND.n590 GND.n589 13.653
R547 GND.n593 GND.n592 13.653
R548 GND.n596 GND.n595 13.653
R549 GND.n599 GND.n598 13.653
R550 GND.n602 GND.n601 13.653
R551 GND.n605 GND.n604 13.653
R552 GND.n608 GND.n607 13.653
R553 GND.n615 GND.n610 13.653
R554 GND.n618 GND.n617 13.653
R555 GND.n623 GND.n620 13.653
R556 GND.n626 GND.n625 13.653
R557 GND.n629 GND.n628 13.653
R558 GND.n632 GND.n631 13.653
R559 GND.n635 GND.n634 13.653
R560 GND.n638 GND.n637 13.653
R561 GND.n641 GND.n640 13.653
R562 GND.n644 GND.n643 13.653
R563 GND.n647 GND.n646 13.653
R564 GND.n650 GND.n649 13.653
R565 GND.n657 GND.n652 13.653
R566 GND.n660 GND.n659 13.653
R567 GND.n665 GND.n662 13.653
R568 GND.n668 GND.n667 13.653
R569 GND.n671 GND.n670 13.653
R570 GND.n674 GND.n673 13.653
R571 GND.n677 GND.n676 13.653
R572 GND.n680 GND.n679 13.653
R573 GND.n683 GND.n682 13.653
R574 GND.n686 GND.n685 13.653
R575 GND.n689 GND.n688 13.653
R576 GND.n692 GND.n691 13.653
R577 GND.n699 GND.n694 13.653
R578 GND.n702 GND.n701 13.653
R579 GND.n710 GND.n704 13.653
R580 GND.n713 GND.n712 13.653
R581 GND.n716 GND.n715 13.653
R582 GND.n719 GND.n718 13.653
R583 GND.n722 GND.n721 13.653
R584 GND.n725 GND.n724 13.653
R585 GND.n728 GND.n727 13.653
R586 GND.n731 GND.n730 13.653
R587 GND.n734 GND.n733 13.653
R588 GND.n737 GND.n736 13.653
R589 GND.n744 GND.n739 13.653
R590 GND.n747 GND.n746 13.653
R591 GND.n752 GND.n749 13.653
R592 GND.n755 GND.n754 13.653
R593 GND.n758 GND.n757 13.653
R594 GND.n761 GND.n760 13.653
R595 GND.n764 GND.n763 13.653
R596 GND.n767 GND.n766 13.653
R597 GND.n770 GND.n769 13.653
R598 GND.n773 GND.n772 13.653
R599 GND.n776 GND.n775 13.653
R600 GND.n779 GND.n778 13.653
R601 GND.n786 GND.n781 13.653
R602 GND.n789 GND.n788 13.653
R603 GND.n797 GND.n791 13.653
R604 GND.n800 GND.n799 13.653
R605 GND.n803 GND.n802 13.653
R606 GND.n806 GND.n805 13.653
R607 GND.n809 GND.n808 13.653
R608 GND.n812 GND.n811 13.653
R609 GND.n815 GND.n814 13.653
R610 GND.n818 GND.n817 13.653
R611 GND.n821 GND.n820 13.653
R612 GND.n824 GND.n823 13.653
R613 GND.n831 GND.n826 13.653
R614 GND.n834 GND.n833 13.653
R615 GND.n839 GND.n836 13.653
R616 GND.n842 GND.n841 13.653
R617 GND.n845 GND.n844 13.653
R618 GND.n848 GND.n847 13.653
R619 GND.n851 GND.n850 13.653
R620 GND.n854 GND.n853 13.653
R621 GND.n857 GND.n856 13.653
R622 GND.n860 GND.n859 13.653
R623 GND.n863 GND.n862 13.653
R624 GND.n866 GND.n865 13.653
R625 GND.n873 GND.n868 13.653
R626 GND.n876 GND.n875 13.653
R627 GND.n881 GND.n878 13.653
R628 GND.n444 GND.n443 13.653
R629 GND.n441 GND.n440 13.653
R630 GND.n438 GND.n437 13.653
R631 GND.n435 GND.n434 13.653
R632 GND.n432 GND.n431 13.653
R633 GND.n429 GND.n428 13.653
R634 GND.n426 GND.n425 13.653
R635 GND.n423 GND.n422 13.653
R636 GND.n420 GND.n419 13.653
R637 GND.n413 GND.n412 13.653
R638 GND.n410 GND.n409 13.653
R639 GND.n407 GND.n404 13.653
R640 GND.n402 GND.n401 13.653
R641 GND.n399 GND.n398 13.653
R642 GND.n396 GND.n395 13.653
R643 GND.n393 GND.n392 13.653
R644 GND.n390 GND.n389 13.653
R645 GND.n387 GND.n386 13.653
R646 GND.n384 GND.n383 13.653
R647 GND.n381 GND.n380 13.653
R648 GND.n378 GND.n377 13.653
R649 GND.n371 GND.n370 13.653
R650 GND.n368 GND.n367 13.653
R651 GND.n365 GND.n362 13.653
R652 GND.n360 GND.n359 13.653
R653 GND.n357 GND.n356 13.653
R654 GND.n354 GND.n353 13.653
R655 GND.n351 GND.n350 13.653
R656 GND.n348 GND.n347 13.653
R657 GND.n345 GND.n344 13.653
R658 GND.n342 GND.n341 13.653
R659 GND.n339 GND.n338 13.653
R660 GND.n336 GND.n335 13.653
R661 GND.n329 GND.n328 13.653
R662 GND.n326 GND.n325 13.653
R663 GND.n323 GND.n320 13.653
R664 GND.n318 GND.n317 13.653
R665 GND.n315 GND.n314 13.653
R666 GND.n312 GND.n311 13.653
R667 GND.n309 GND.n308 13.653
R668 GND.n306 GND.n305 13.653
R669 GND.n303 GND.n302 13.653
R670 GND.n300 GND.n299 13.653
R671 GND.n297 GND.n296 13.653
R672 GND.n294 GND.n293 13.653
R673 GND.n287 GND.n286 13.653
R674 GND.n284 GND.n283 13.653
R675 GND.n281 GND.n278 13.653
R676 GND.n276 GND.n275 13.653
R677 GND.n273 GND.n272 13.653
R678 GND.n270 GND.n269 13.653
R679 GND.n267 GND.n266 13.653
R680 GND.n264 GND.n263 13.653
R681 GND.n261 GND.n260 13.653
R682 GND.n258 GND.n257 13.653
R683 GND.n255 GND.n254 13.653
R684 GND.n252 GND.n251 13.653
R685 GND.n245 GND.n244 13.653
R686 GND.n242 GND.n241 13.653
R687 GND.n239 GND.n233 13.653
R688 GND.n231 GND.n230 13.653
R689 GND.n228 GND.n227 13.653
R690 GND.n225 GND.n224 13.653
R691 GND.n222 GND.n221 13.653
R692 GND.n219 GND.n218 13.653
R693 GND.n216 GND.n215 13.653
R694 GND.n213 GND.n212 13.653
R695 GND.n210 GND.n209 13.653
R696 GND.n207 GND.n206 13.653
R697 GND.n200 GND.n199 13.653
R698 GND.n197 GND.n196 13.653
R699 GND.n194 GND.n191 13.653
R700 GND.n189 GND.n188 13.653
R701 GND.n186 GND.n185 13.653
R702 GND.n183 GND.n182 13.653
R703 GND.n180 GND.n179 13.653
R704 GND.n177 GND.n176 13.653
R705 GND.n174 GND.n173 13.653
R706 GND.n171 GND.n170 13.653
R707 GND.n168 GND.n167 13.653
R708 GND.n165 GND.n164 13.653
R709 GND.n158 GND.n157 13.653
R710 GND.n155 GND.n154 13.653
R711 GND.n152 GND.n149 13.653
R712 GND.n147 GND.n146 13.653
R713 GND.n144 GND.n143 13.653
R714 GND.n141 GND.n140 13.653
R715 GND.n138 GND.n137 13.653
R716 GND.n135 GND.n134 13.653
R717 GND.n132 GND.n131 13.653
R718 GND.n129 GND.n128 13.653
R719 GND.n126 GND.n125 13.653
R720 GND.n123 GND.n122 13.653
R721 GND.n116 GND.n115 13.653
R722 GND.n113 GND.n112 13.653
R723 GND.n110 GND.n109 13.653
R724 GND.n105 GND.n104 13.653
R725 GND.n102 GND.n101 13.653
R726 GND.n99 GND.n98 13.653
R727 GND.n96 GND.n95 13.653
R728 GND.n93 GND.n92 13.653
R729 GND.n86 GND.n85 13.653
R730 GND.n83 GND.n82 13.653
R731 GND.n80 GND.n79 13.653
R732 GND.n75 GND.n74 13.653
R733 GND.n72 GND.n71 13.653
R734 GND.n8 GND.n7 13.653
R735 GND.n16 GND.n15 13.653
R736 GND.n23 GND.n22 13.653
R737 GND.n26 GND.n25 13.653
R738 GND.n33 GND.n32 13.653
R739 GND.n36 GND.n35 13.653
R740 GND.n39 GND.n38 13.653
R741 GND.n42 GND.n41 13.653
R742 GND.n45 GND.n44 13.653
R743 GND.n50 GND.n49 13.653
R744 GND.n53 GND.n52 13.653
R745 GND.n56 GND.n55 13.653
R746 GND.n63 GND.n62 13.653
R747 GND.n66 GND.n65 13.653
R748 GND.n69 GND.n68 13.653
R749 GND.n20 GND.n19 12.837
R750 GND.n19 GND.n18 7.566
R751 GND.n31 GND.n30 7.312
R752 GND.n61 GND.n60 7.312
R753 GND.n91 GND.n90 7.312
R754 GND.n488 GND.n487 7.312
R755 GND.n530 GND.n529 7.312
R756 GND.n572 GND.n571 7.312
R757 GND.n614 GND.n613 7.312
R758 GND.n656 GND.n655 7.312
R759 GND.n698 GND.n697 7.312
R760 GND.n743 GND.n742 7.312
R761 GND.n785 GND.n784 7.312
R762 GND.n830 GND.n829 7.312
R763 GND.n872 GND.n871 7.312
R764 GND.n418 GND.n417 7.312
R765 GND.n376 GND.n375 7.312
R766 GND.n334 GND.n333 7.312
R767 GND.n292 GND.n291 7.312
R768 GND.n250 GND.n249 7.312
R769 GND.n205 GND.n204 7.312
R770 GND.n163 GND.n162 7.312
R771 GND.n121 GND.n120 7.312
R772 GND.n11 GND.n10 4.551
R773 GND.n8 GND.n6 3.935
R774 GND.n50 GND.n48 3.935
R775 GND.n80 GND.n78 3.935
R776 GND.n110 GND.n108 3.935
R777 GND.n23 GND.n21 3.541
R778 GND.t15 GND.n11 2.238
R779 GND.n447 GND.n446 0.596
R780 GND.n1 GND.n0 0.596
R781 GND.n13 GND.n12 0.358
R782 GND.n34 GND.n27 0.29
R783 GND.n64 GND.n57 0.29
R784 GND.n94 GND.n87 0.29
R785 GND.n124 GND.n117 0.29
R786 GND.n166 GND.n159 0.29
R787 GND.n208 GND.n201 0.29
R788 GND.n253 GND.n246 0.29
R789 GND.n295 GND.n288 0.29
R790 GND.n337 GND.n330 0.29
R791 GND.n379 GND.n372 0.29
R792 GND.n421 GND.n414 0.29
R793 GND.n874 GND.n867 0.29
R794 GND.n832 GND.n825 0.29
R795 GND.n787 GND.n780 0.29
R796 GND.n745 GND.n738 0.29
R797 GND.n700 GND.n693 0.29
R798 GND.n658 GND.n651 0.29
R799 GND.n616 GND.n609 0.29
R800 GND.n574 GND.n567 0.29
R801 GND.n532 GND.n525 0.29
R802 GND.n490 GND.n483 0.29
R803 GND.n448 GND 0.207
R804 GND.n142 GND.n139 0.197
R805 GND.n184 GND.n181 0.197
R806 GND.n226 GND.n223 0.197
R807 GND.n271 GND.n268 0.197
R808 GND.n313 GND.n310 0.197
R809 GND.n355 GND.n352 0.197
R810 GND.n397 GND.n394 0.197
R811 GND.n439 GND.n436 0.197
R812 GND.n852 GND.n849 0.197
R813 GND.n810 GND.n807 0.197
R814 GND.n765 GND.n762 0.197
R815 GND.n723 GND.n720 0.197
R816 GND.n678 GND.n675 0.197
R817 GND.n636 GND.n633 0.197
R818 GND.n594 GND.n591 0.197
R819 GND.n552 GND.n549 0.197
R820 GND.n510 GND.n507 0.197
R821 GND.n468 GND.n465 0.197
R822 GND.n16 GND.n14 0.196
R823 GND.n152 GND.n151 0.196
R824 GND.n194 GND.n193 0.196
R825 GND.n239 GND.n238 0.196
R826 GND.n281 GND.n280 0.196
R827 GND.n323 GND.n322 0.196
R828 GND.n365 GND.n364 0.196
R829 GND.n407 GND.n406 0.196
R830 GND.n881 GND.n880 0.196
R831 GND.n839 GND.n838 0.196
R832 GND.n797 GND.n796 0.196
R833 GND.n752 GND.n751 0.196
R834 GND.n710 GND.n709 0.196
R835 GND.n665 GND.n664 0.196
R836 GND.n623 GND.n622 0.196
R837 GND.n581 GND.n580 0.196
R838 GND.n539 GND.n538 0.196
R839 GND.n497 GND.n496 0.196
R840 GND.n455 GND.n454 0.196
R841 GND.n46 GND.n43 0.181
R842 GND.n76 GND.n73 0.181
R843 GND.n106 GND.n103 0.181
R844 GND.n17 GND.n9 0.157
R845 GND.n24 GND.n17 0.157
R846 GND.n27 GND.n24 0.145
R847 GND.n37 GND.n34 0.145
R848 GND.n40 GND.n37 0.145
R849 GND.n43 GND.n40 0.145
R850 GND.n51 GND.n46 0.145
R851 GND.n54 GND.n51 0.145
R852 GND.n57 GND.n54 0.145
R853 GND.n67 GND.n64 0.145
R854 GND.n70 GND.n67 0.145
R855 GND.n73 GND.n70 0.145
R856 GND.n81 GND.n76 0.145
R857 GND.n84 GND.n81 0.145
R858 GND.n87 GND.n84 0.145
R859 GND.n97 GND.n94 0.145
R860 GND.n100 GND.n97 0.145
R861 GND.n103 GND.n100 0.145
R862 GND.n111 GND.n106 0.145
R863 GND.n114 GND.n111 0.145
R864 GND.n117 GND.n114 0.145
R865 GND.n127 GND.n124 0.145
R866 GND.n130 GND.n127 0.145
R867 GND.n133 GND.n130 0.145
R868 GND.n136 GND.n133 0.145
R869 GND.n139 GND.n136 0.145
R870 GND.n145 GND.n142 0.145
R871 GND.n148 GND.n145 0.145
R872 GND.n153 GND.n148 0.145
R873 GND.n156 GND.n153 0.145
R874 GND.n159 GND.n156 0.145
R875 GND.n169 GND.n166 0.145
R876 GND.n172 GND.n169 0.145
R877 GND.n175 GND.n172 0.145
R878 GND.n178 GND.n175 0.145
R879 GND.n181 GND.n178 0.145
R880 GND.n187 GND.n184 0.145
R881 GND.n190 GND.n187 0.145
R882 GND.n195 GND.n190 0.145
R883 GND.n198 GND.n195 0.145
R884 GND.n201 GND.n198 0.145
R885 GND.n211 GND.n208 0.145
R886 GND.n214 GND.n211 0.145
R887 GND.n217 GND.n214 0.145
R888 GND.n220 GND.n217 0.145
R889 GND.n223 GND.n220 0.145
R890 GND.n229 GND.n226 0.145
R891 GND.n232 GND.n229 0.145
R892 GND.n240 GND.n232 0.145
R893 GND.n243 GND.n240 0.145
R894 GND.n246 GND.n243 0.145
R895 GND.n256 GND.n253 0.145
R896 GND.n259 GND.n256 0.145
R897 GND.n262 GND.n259 0.145
R898 GND.n265 GND.n262 0.145
R899 GND.n268 GND.n265 0.145
R900 GND.n274 GND.n271 0.145
R901 GND.n277 GND.n274 0.145
R902 GND.n282 GND.n277 0.145
R903 GND.n285 GND.n282 0.145
R904 GND.n288 GND.n285 0.145
R905 GND.n298 GND.n295 0.145
R906 GND.n301 GND.n298 0.145
R907 GND.n304 GND.n301 0.145
R908 GND.n307 GND.n304 0.145
R909 GND.n310 GND.n307 0.145
R910 GND.n316 GND.n313 0.145
R911 GND.n319 GND.n316 0.145
R912 GND.n324 GND.n319 0.145
R913 GND.n327 GND.n324 0.145
R914 GND.n330 GND.n327 0.145
R915 GND.n340 GND.n337 0.145
R916 GND.n343 GND.n340 0.145
R917 GND.n346 GND.n343 0.145
R918 GND.n349 GND.n346 0.145
R919 GND.n352 GND.n349 0.145
R920 GND.n358 GND.n355 0.145
R921 GND.n361 GND.n358 0.145
R922 GND.n366 GND.n361 0.145
R923 GND.n369 GND.n366 0.145
R924 GND.n372 GND.n369 0.145
R925 GND.n382 GND.n379 0.145
R926 GND.n385 GND.n382 0.145
R927 GND.n388 GND.n385 0.145
R928 GND.n391 GND.n388 0.145
R929 GND.n394 GND.n391 0.145
R930 GND.n400 GND.n397 0.145
R931 GND.n403 GND.n400 0.145
R932 GND.n408 GND.n403 0.145
R933 GND.n411 GND.n408 0.145
R934 GND.n414 GND.n411 0.145
R935 GND.n424 GND.n421 0.145
R936 GND.n427 GND.n424 0.145
R937 GND.n430 GND.n427 0.145
R938 GND.n433 GND.n430 0.145
R939 GND.n436 GND.n433 0.145
R940 GND.n442 GND.n439 0.145
R941 GND.n445 GND.n442 0.145
R942 GND.n882 GND.n877 0.145
R943 GND.n877 GND.n874 0.145
R944 GND.n867 GND.n864 0.145
R945 GND.n864 GND.n861 0.145
R946 GND.n861 GND.n858 0.145
R947 GND.n858 GND.n855 0.145
R948 GND.n855 GND.n852 0.145
R949 GND.n849 GND.n846 0.145
R950 GND.n846 GND.n843 0.145
R951 GND.n843 GND.n840 0.145
R952 GND.n840 GND.n835 0.145
R953 GND.n835 GND.n832 0.145
R954 GND.n825 GND.n822 0.145
R955 GND.n822 GND.n819 0.145
R956 GND.n819 GND.n816 0.145
R957 GND.n816 GND.n813 0.145
R958 GND.n813 GND.n810 0.145
R959 GND.n807 GND.n804 0.145
R960 GND.n804 GND.n801 0.145
R961 GND.n801 GND.n798 0.145
R962 GND.n798 GND.n790 0.145
R963 GND.n790 GND.n787 0.145
R964 GND.n780 GND.n777 0.145
R965 GND.n777 GND.n774 0.145
R966 GND.n774 GND.n771 0.145
R967 GND.n771 GND.n768 0.145
R968 GND.n768 GND.n765 0.145
R969 GND.n762 GND.n759 0.145
R970 GND.n759 GND.n756 0.145
R971 GND.n756 GND.n753 0.145
R972 GND.n753 GND.n748 0.145
R973 GND.n748 GND.n745 0.145
R974 GND.n738 GND.n735 0.145
R975 GND.n735 GND.n732 0.145
R976 GND.n732 GND.n729 0.145
R977 GND.n729 GND.n726 0.145
R978 GND.n726 GND.n723 0.145
R979 GND.n720 GND.n717 0.145
R980 GND.n717 GND.n714 0.145
R981 GND.n714 GND.n711 0.145
R982 GND.n711 GND.n703 0.145
R983 GND.n703 GND.n700 0.145
R984 GND.n693 GND.n690 0.145
R985 GND.n690 GND.n687 0.145
R986 GND.n687 GND.n684 0.145
R987 GND.n684 GND.n681 0.145
R988 GND.n681 GND.n678 0.145
R989 GND.n675 GND.n672 0.145
R990 GND.n672 GND.n669 0.145
R991 GND.n669 GND.n666 0.145
R992 GND.n666 GND.n661 0.145
R993 GND.n661 GND.n658 0.145
R994 GND.n651 GND.n648 0.145
R995 GND.n648 GND.n645 0.145
R996 GND.n645 GND.n642 0.145
R997 GND.n642 GND.n639 0.145
R998 GND.n639 GND.n636 0.145
R999 GND.n633 GND.n630 0.145
R1000 GND.n630 GND.n627 0.145
R1001 GND.n627 GND.n624 0.145
R1002 GND.n624 GND.n619 0.145
R1003 GND.n619 GND.n616 0.145
R1004 GND.n609 GND.n606 0.145
R1005 GND.n606 GND.n603 0.145
R1006 GND.n603 GND.n600 0.145
R1007 GND.n600 GND.n597 0.145
R1008 GND.n597 GND.n594 0.145
R1009 GND.n591 GND.n588 0.145
R1010 GND.n588 GND.n585 0.145
R1011 GND.n585 GND.n582 0.145
R1012 GND.n582 GND.n577 0.145
R1013 GND.n577 GND.n574 0.145
R1014 GND.n567 GND.n564 0.145
R1015 GND.n564 GND.n561 0.145
R1016 GND.n561 GND.n558 0.145
R1017 GND.n558 GND.n555 0.145
R1018 GND.n555 GND.n552 0.145
R1019 GND.n549 GND.n546 0.145
R1020 GND.n546 GND.n543 0.145
R1021 GND.n543 GND.n540 0.145
R1022 GND.n540 GND.n535 0.145
R1023 GND.n535 GND.n532 0.145
R1024 GND.n525 GND.n522 0.145
R1025 GND.n522 GND.n519 0.145
R1026 GND.n519 GND.n516 0.145
R1027 GND.n516 GND.n513 0.145
R1028 GND.n513 GND.n510 0.145
R1029 GND.n507 GND.n504 0.145
R1030 GND.n504 GND.n501 0.145
R1031 GND.n501 GND.n498 0.145
R1032 GND.n498 GND.n493 0.145
R1033 GND.n493 GND.n490 0.145
R1034 GND.n483 GND.n480 0.145
R1035 GND.n480 GND.n477 0.145
R1036 GND.n477 GND.n474 0.145
R1037 GND.n474 GND.n471 0.145
R1038 GND.n471 GND.n468 0.145
R1039 GND.n465 GND.n462 0.145
R1040 GND.n462 GND.n459 0.145
R1041 GND.n459 GND.n456 0.145
R1042 GND.n456 GND.n451 0.145
R1043 GND.n451 GND.n448 0.145
R1044 GND GND.n882 0.086
R1045 GND GND.n445 0.058
R1046 a_10219_989.n5 a_10219_989.t9 475.572
R1047 a_10219_989.n7 a_10219_989.t7 469.145
R1048 a_10219_989.n11 a_10219_989.t12 454.685
R1049 a_10219_989.n11 a_10219_989.t8 428.979
R1050 a_10219_989.n7 a_10219_989.t11 384.527
R1051 a_10219_989.n5 a_10219_989.t13 384.527
R1052 a_10219_989.n8 a_10219_989.t14 294.278
R1053 a_10219_989.n6 a_10219_989.t10 294.278
R1054 a_10219_989.n12 a_10219_989.t15 184.853
R1055 a_10219_989.n15 a_10219_989.n13 166.52
R1056 a_10219_989.n13 a_10219_989.n12 156.035
R1057 a_10219_989.n12 a_10219_989.n11 151.553
R1058 a_10219_989.n10 a_10219_989.n4 144.246
R1059 a_10219_989.n10 a_10219_989.n9 99.225
R1060 a_10219_989.n9 a_10219_989.n6 80.851
R1061 a_10219_989.n13 a_10219_989.n10 79.658
R1062 a_10219_989.n3 a_10219_989.n2 79.232
R1063 a_10219_989.n9 a_10219_989.n8 76
R1064 a_10219_989.n4 a_10219_989.n3 63.152
R1065 a_10219_989.n6 a_10219_989.n5 57.842
R1066 a_10219_989.n8 a_10219_989.n7 56.833
R1067 a_10219_989.n4 a_10219_989.n0 16.08
R1068 a_10219_989.n3 a_10219_989.n1 16.08
R1069 a_10219_989.n15 a_10219_989.n14 15.218
R1070 a_10219_989.n0 a_10219_989.t1 14.282
R1071 a_10219_989.n0 a_10219_989.t2 14.282
R1072 a_10219_989.n1 a_10219_989.t4 14.282
R1073 a_10219_989.n1 a_10219_989.t0 14.282
R1074 a_10219_989.n2 a_10219_989.t6 14.282
R1075 a_10219_989.n2 a_10219_989.t5 14.282
R1076 a_10219_989.n16 a_10219_989.n15 12.014
R1077 a_17533_1051.n3 a_17533_1051.n2 195.987
R1078 a_17533_1051.n4 a_17533_1051.t7 89.553
R1079 a_17533_1051.n2 a_17533_1051.n1 75.271
R1080 a_17533_1051.n4 a_17533_1051.n3 75.214
R1081 a_17533_1051.n2 a_17533_1051.n0 36.519
R1082 a_17533_1051.n3 a_17533_1051.t1 14.338
R1083 a_17533_1051.n0 a_17533_1051.t6 14.282
R1084 a_17533_1051.n0 a_17533_1051.t5 14.282
R1085 a_17533_1051.n1 a_17533_1051.t3 14.282
R1086 a_17533_1051.n1 a_17533_1051.t4 14.282
R1087 a_17533_1051.t0 a_17533_1051.n5 14.282
R1088 a_17533_1051.n5 a_17533_1051.t2 14.282
R1089 a_17533_1051.n5 a_17533_1051.n4 12.122
R1090 VDD.n951 VDD.n949 144.705
R1091 VDD.n1032 VDD.n1030 144.705
R1092 VDD.n1113 VDD.n1111 144.705
R1093 VDD.n1194 VDD.n1192 144.705
R1094 VDD.n1275 VDD.n1273 144.705
R1095 VDD.n1356 VDD.n1354 144.705
R1096 VDD.n1437 VDD.n1435 144.705
R1097 VDD.n1518 VDD.n1516 144.705
R1098 VDD.n1599 VDD.n1597 144.705
R1099 VDD.n804 VDD.n802 144.705
R1100 VDD.n1680 VDD.n1678 144.705
R1101 VDD.n723 VDD.n721 144.705
R1102 VDD.n642 VDD.n640 144.705
R1103 VDD.n561 VDD.n559 144.705
R1104 VDD.n480 VDD.n478 144.705
R1105 VDD.n399 VDD.n397 144.705
R1106 VDD.n318 VDD.n316 144.705
R1107 VDD.n237 VDD.n235 144.705
R1108 VDD.n176 VDD.n174 144.705
R1109 VDD.n122 VDD.n120 144.705
R1110 VDD.n68 VDD.n66 144.705
R1111 VDD.n26 VDD.n25 77.792
R1112 VDD.n35 VDD.n34 77.792
R1113 VDD.n29 VDD.n23 76.145
R1114 VDD.n29 VDD.n28 76
R1115 VDD.n33 VDD.n32 76
R1116 VDD.n39 VDD.n38 76
R1117 VDD.n43 VDD.n42 76
R1118 VDD.n70 VDD.n69 76
R1119 VDD.n74 VDD.n73 76
R1120 VDD.n78 VDD.n77 76
R1121 VDD.n82 VDD.n81 76
R1122 VDD.n86 VDD.n85 76
R1123 VDD.n90 VDD.n89 76
R1124 VDD.n94 VDD.n93 76
R1125 VDD.n98 VDD.n97 76
R1126 VDD.n124 VDD.n123 76
R1127 VDD.n128 VDD.n127 76
R1128 VDD.n132 VDD.n131 76
R1129 VDD.n136 VDD.n135 76
R1130 VDD.n140 VDD.n139 76
R1131 VDD.n144 VDD.n143 76
R1132 VDD.n148 VDD.n147 76
R1133 VDD.n152 VDD.n151 76
R1134 VDD.n178 VDD.n177 76
R1135 VDD.n183 VDD.n182 76
R1136 VDD.n188 VDD.n187 76
R1137 VDD.n194 VDD.n193 76
R1138 VDD.n199 VDD.n198 76
R1139 VDD.n204 VDD.n203 76
R1140 VDD.n209 VDD.n208 76
R1141 VDD.n213 VDD.n212 76
R1142 VDD.n239 VDD.n238 76
R1143 VDD.n243 VDD.n242 76
R1144 VDD.n247 VDD.n246 76
R1145 VDD.n252 VDD.n251 76
R1146 VDD.n259 VDD.n258 76
R1147 VDD.n264 VDD.n263 76
R1148 VDD.n269 VDD.n268 76
R1149 VDD.n276 VDD.n275 76
R1150 VDD.n281 VDD.n280 76
R1151 VDD.n286 VDD.n285 76
R1152 VDD.n290 VDD.n289 76
R1153 VDD.n294 VDD.n293 76
R1154 VDD.n320 VDD.n319 76
R1155 VDD.n324 VDD.n323 76
R1156 VDD.n328 VDD.n327 76
R1157 VDD.n333 VDD.n332 76
R1158 VDD.n340 VDD.n339 76
R1159 VDD.n345 VDD.n344 76
R1160 VDD.n350 VDD.n349 76
R1161 VDD.n357 VDD.n356 76
R1162 VDD.n362 VDD.n361 76
R1163 VDD.n367 VDD.n366 76
R1164 VDD.n371 VDD.n370 76
R1165 VDD.n375 VDD.n374 76
R1166 VDD.n401 VDD.n400 76
R1167 VDD.n405 VDD.n404 76
R1168 VDD.n409 VDD.n408 76
R1169 VDD.n414 VDD.n413 76
R1170 VDD.n421 VDD.n420 76
R1171 VDD.n426 VDD.n425 76
R1172 VDD.n431 VDD.n430 76
R1173 VDD.n438 VDD.n437 76
R1174 VDD.n443 VDD.n442 76
R1175 VDD.n448 VDD.n447 76
R1176 VDD.n452 VDD.n451 76
R1177 VDD.n456 VDD.n455 76
R1178 VDD.n482 VDD.n481 76
R1179 VDD.n486 VDD.n485 76
R1180 VDD.n490 VDD.n489 76
R1181 VDD.n495 VDD.n494 76
R1182 VDD.n502 VDD.n501 76
R1183 VDD.n507 VDD.n506 76
R1184 VDD.n512 VDD.n511 76
R1185 VDD.n519 VDD.n518 76
R1186 VDD.n524 VDD.n523 76
R1187 VDD.n529 VDD.n528 76
R1188 VDD.n533 VDD.n532 76
R1189 VDD.n537 VDD.n536 76
R1190 VDD.n563 VDD.n562 76
R1191 VDD.n567 VDD.n566 76
R1192 VDD.n571 VDD.n570 76
R1193 VDD.n576 VDD.n575 76
R1194 VDD.n583 VDD.n582 76
R1195 VDD.n588 VDD.n587 76
R1196 VDD.n593 VDD.n592 76
R1197 VDD.n600 VDD.n599 76
R1198 VDD.n605 VDD.n604 76
R1199 VDD.n610 VDD.n609 76
R1200 VDD.n614 VDD.n613 76
R1201 VDD.n618 VDD.n617 76
R1202 VDD.n644 VDD.n643 76
R1203 VDD.n648 VDD.n647 76
R1204 VDD.n652 VDD.n651 76
R1205 VDD.n657 VDD.n656 76
R1206 VDD.n664 VDD.n663 76
R1207 VDD.n669 VDD.n668 76
R1208 VDD.n674 VDD.n673 76
R1209 VDD.n681 VDD.n680 76
R1210 VDD.n686 VDD.n685 76
R1211 VDD.n691 VDD.n690 76
R1212 VDD.n695 VDD.n694 76
R1213 VDD.n699 VDD.n698 76
R1214 VDD.n725 VDD.n724 76
R1215 VDD.n729 VDD.n728 76
R1216 VDD.n733 VDD.n732 76
R1217 VDD.n738 VDD.n737 76
R1218 VDD.n745 VDD.n744 76
R1219 VDD.n750 VDD.n749 76
R1220 VDD.n755 VDD.n754 76
R1221 VDD.n762 VDD.n761 76
R1222 VDD.n767 VDD.n766 76
R1223 VDD.n772 VDD.n771 76
R1224 VDD.n776 VDD.n775 76
R1225 VDD.n780 VDD.n779 76
R1226 VDD.n806 VDD.n805 76
R1227 VDD.n810 VDD.n809 76
R1228 VDD.n814 VDD.n813 76
R1229 VDD.n819 VDD.n818 76
R1230 VDD.n826 VDD.n825 76
R1231 VDD.n831 VDD.n830 76
R1232 VDD.n836 VDD.n835 76
R1233 VDD.n843 VDD.n842 76
R1234 VDD.n848 VDD.n847 76
R1235 VDD.n1691 VDD.n1690 76
R1236 VDD.n1686 VDD.n1685 76
R1237 VDD.n1682 VDD.n1681 76
R1238 VDD.n1656 VDD.n1655 76
R1239 VDD.n1652 VDD.n1651 76
R1240 VDD.n1648 VDD.n1647 76
R1241 VDD.n1644 VDD.n1643 76
R1242 VDD.n1639 VDD.n1638 76
R1243 VDD.n1632 VDD.n1631 76
R1244 VDD.n1627 VDD.n1626 76
R1245 VDD.n1622 VDD.n1621 76
R1246 VDD.n1615 VDD.n1614 76
R1247 VDD.n1610 VDD.n1609 76
R1248 VDD.n1605 VDD.n1604 76
R1249 VDD.n1601 VDD.n1600 76
R1250 VDD.n1575 VDD.n1574 76
R1251 VDD.n1571 VDD.n1570 76
R1252 VDD.n1567 VDD.n1566 76
R1253 VDD.n1563 VDD.n1562 76
R1254 VDD.n1558 VDD.n1557 76
R1255 VDD.n1551 VDD.n1550 76
R1256 VDD.n1546 VDD.n1545 76
R1257 VDD.n1541 VDD.n1540 76
R1258 VDD.n1534 VDD.n1533 76
R1259 VDD.n1529 VDD.n1528 76
R1260 VDD.n1524 VDD.n1523 76
R1261 VDD.n1520 VDD.n1519 76
R1262 VDD.n1494 VDD.n1493 76
R1263 VDD.n1490 VDD.n1489 76
R1264 VDD.n1486 VDD.n1485 76
R1265 VDD.n1482 VDD.n1481 76
R1266 VDD.n1477 VDD.n1476 76
R1267 VDD.n1470 VDD.n1469 76
R1268 VDD.n1465 VDD.n1464 76
R1269 VDD.n1460 VDD.n1459 76
R1270 VDD.n1453 VDD.n1452 76
R1271 VDD.n1448 VDD.n1447 76
R1272 VDD.n1443 VDD.n1442 76
R1273 VDD.n1439 VDD.n1438 76
R1274 VDD.n1413 VDD.n1412 76
R1275 VDD.n1409 VDD.n1408 76
R1276 VDD.n1405 VDD.n1404 76
R1277 VDD.n1401 VDD.n1400 76
R1278 VDD.n1396 VDD.n1395 76
R1279 VDD.n1389 VDD.n1388 76
R1280 VDD.n1384 VDD.n1383 76
R1281 VDD.n1379 VDD.n1378 76
R1282 VDD.n1372 VDD.n1371 76
R1283 VDD.n1367 VDD.n1366 76
R1284 VDD.n1362 VDD.n1361 76
R1285 VDD.n1358 VDD.n1357 76
R1286 VDD.n1332 VDD.n1331 76
R1287 VDD.n1328 VDD.n1327 76
R1288 VDD.n1324 VDD.n1323 76
R1289 VDD.n1320 VDD.n1319 76
R1290 VDD.n1315 VDD.n1314 76
R1291 VDD.n1308 VDD.n1307 76
R1292 VDD.n1303 VDD.n1302 76
R1293 VDD.n1298 VDD.n1297 76
R1294 VDD.n1291 VDD.n1290 76
R1295 VDD.n1286 VDD.n1285 76
R1296 VDD.n1281 VDD.n1280 76
R1297 VDD.n1277 VDD.n1276 76
R1298 VDD.n1251 VDD.n1250 76
R1299 VDD.n1247 VDD.n1246 76
R1300 VDD.n1243 VDD.n1242 76
R1301 VDD.n1239 VDD.n1238 76
R1302 VDD.n1234 VDD.n1233 76
R1303 VDD.n1227 VDD.n1226 76
R1304 VDD.n1222 VDD.n1221 76
R1305 VDD.n1217 VDD.n1216 76
R1306 VDD.n1210 VDD.n1209 76
R1307 VDD.n1205 VDD.n1204 76
R1308 VDD.n1200 VDD.n1199 76
R1309 VDD.n1196 VDD.n1195 76
R1310 VDD.n1170 VDD.n1169 76
R1311 VDD.n1166 VDD.n1165 76
R1312 VDD.n1162 VDD.n1161 76
R1313 VDD.n1158 VDD.n1157 76
R1314 VDD.n1153 VDD.n1152 76
R1315 VDD.n1146 VDD.n1145 76
R1316 VDD.n1141 VDD.n1140 76
R1317 VDD.n1136 VDD.n1135 76
R1318 VDD.n1129 VDD.n1128 76
R1319 VDD.n1124 VDD.n1123 76
R1320 VDD.n1119 VDD.n1118 76
R1321 VDD.n1115 VDD.n1114 76
R1322 VDD.n1089 VDD.n1088 76
R1323 VDD.n1085 VDD.n1084 76
R1324 VDD.n1081 VDD.n1080 76
R1325 VDD.n1077 VDD.n1076 76
R1326 VDD.n1072 VDD.n1071 76
R1327 VDD.n1065 VDD.n1064 76
R1328 VDD.n1060 VDD.n1059 76
R1329 VDD.n1055 VDD.n1054 76
R1330 VDD.n1048 VDD.n1047 76
R1331 VDD.n1043 VDD.n1042 76
R1332 VDD.n1038 VDD.n1037 76
R1333 VDD.n1034 VDD.n1033 76
R1334 VDD.n1008 VDD.n1007 76
R1335 VDD.n1004 VDD.n1003 76
R1336 VDD.n1000 VDD.n999 76
R1337 VDD.n996 VDD.n995 76
R1338 VDD.n991 VDD.n990 76
R1339 VDD.n984 VDD.n983 76
R1340 VDD.n979 VDD.n978 76
R1341 VDD.n974 VDD.n973 76
R1342 VDD.n967 VDD.n966 76
R1343 VDD.n962 VDD.n961 76
R1344 VDD.n957 VDD.n956 76
R1345 VDD.n953 VDD.n952 76
R1346 VDD.n926 VDD.n925 76
R1347 VDD.n922 VDD.n921 76
R1348 VDD.n918 VDD.n917 76
R1349 VDD.n914 VDD.n913 76
R1350 VDD.n909 VDD.n908 76
R1351 VDD.n902 VDD.n901 76
R1352 VDD.n897 VDD.n896 76
R1353 VDD.n892 VDD.n891 76
R1354 VDD.n885 VDD.n884 76
R1355 VDD.n880 VDD.n879 76
R1356 VDD.n875 VDD.n874 76
R1357 VDD.n871 VDD.n870 76
R1358 VDD.n249 VDD.n248 64.064
R1359 VDD.n330 VDD.n329 64.064
R1360 VDD.n411 VDD.n410 64.064
R1361 VDD.n492 VDD.n491 64.064
R1362 VDD.n573 VDD.n572 64.064
R1363 VDD.n654 VDD.n653 64.064
R1364 VDD.n735 VDD.n734 64.064
R1365 VDD.n816 VDD.n815 64.064
R1366 VDD.n1641 VDD.n1640 64.064
R1367 VDD.n1560 VDD.n1559 64.064
R1368 VDD.n1479 VDD.n1478 64.064
R1369 VDD.n1398 VDD.n1397 64.064
R1370 VDD.n1317 VDD.n1316 64.064
R1371 VDD.n1236 VDD.n1235 64.064
R1372 VDD.n1155 VDD.n1154 64.064
R1373 VDD.n1074 VDD.n1073 64.064
R1374 VDD.n993 VDD.n992 64.064
R1375 VDD.n911 VDD.n910 64.064
R1376 VDD.n278 VDD.n277 59.488
R1377 VDD.n359 VDD.n358 59.488
R1378 VDD.n440 VDD.n439 59.488
R1379 VDD.n521 VDD.n520 59.488
R1380 VDD.n602 VDD.n601 59.488
R1381 VDD.n683 VDD.n682 59.488
R1382 VDD.n764 VDD.n763 59.488
R1383 VDD.n845 VDD.n844 59.488
R1384 VDD.n1612 VDD.n1611 59.488
R1385 VDD.n1531 VDD.n1530 59.488
R1386 VDD.n1450 VDD.n1449 59.488
R1387 VDD.n1369 VDD.n1368 59.488
R1388 VDD.n1288 VDD.n1287 59.488
R1389 VDD.n1207 VDD.n1206 59.488
R1390 VDD.n1126 VDD.n1125 59.488
R1391 VDD.n1045 VDD.n1044 59.488
R1392 VDD.n964 VDD.n963 59.488
R1393 VDD.n882 VDD.n881 59.488
R1394 VDD.n205 VDD.t39 55.465
R1395 VDD.n179 VDD.t60 55.465
R1396 VDD.n876 VDD.t89 55.106
R1397 VDD.n958 VDD.t101 55.106
R1398 VDD.n1039 VDD.t27 55.106
R1399 VDD.n1120 VDD.t50 55.106
R1400 VDD.n1201 VDD.t28 55.106
R1401 VDD.n1282 VDD.t45 55.106
R1402 VDD.n1363 VDD.t0 55.106
R1403 VDD.n1444 VDD.t56 55.106
R1404 VDD.n1525 VDD.t57 55.106
R1405 VDD.n1606 VDD.t113 55.106
R1406 VDD.n1687 VDD.t88 55.106
R1407 VDD.n768 VDD.t92 55.106
R1408 VDD.n687 VDD.t52 55.106
R1409 VDD.n606 VDD.t98 55.106
R1410 VDD.n525 VDD.t43 55.106
R1411 VDD.n444 VDD.t46 55.106
R1412 VDD.n363 VDD.t108 55.106
R1413 VDD.n282 VDD.t25 55.106
R1414 VDD.n37 VDD.t26 55.106
R1415 VDD.n24 VDD.t100 55.106
R1416 VDD.n917 VDD.t81 55.106
R1417 VDD.n999 VDD.t74 55.106
R1418 VDD.n1080 VDD.t73 55.106
R1419 VDD.n1161 VDD.t104 55.106
R1420 VDD.n1242 VDD.t95 55.106
R1421 VDD.n1323 VDD.t111 55.106
R1422 VDD.n1404 VDD.t72 55.106
R1423 VDD.n1485 VDD.t75 55.106
R1424 VDD.n1566 VDD.t49 55.106
R1425 VDD.n1647 VDD.t67 55.106
R1426 VDD.n813 VDD.t61 55.106
R1427 VDD.n732 VDD.t4 55.106
R1428 VDD.n651 VDD.t107 55.106
R1429 VDD.n570 VDD.t30 55.106
R1430 VDD.n489 VDD.t33 55.106
R1431 VDD.n408 VDD.t22 55.106
R1432 VDD.n327 VDD.t37 55.106
R1433 VDD.n246 VDD.t34 55.106
R1434 VDD.n190 VDD.n189 41.183
R1435 VDD.n887 VDD.n886 40.824
R1436 VDD.n907 VDD.n906 40.824
R1437 VDD.n969 VDD.n968 40.824
R1438 VDD.n989 VDD.n988 40.824
R1439 VDD.n1050 VDD.n1049 40.824
R1440 VDD.n1070 VDD.n1069 40.824
R1441 VDD.n1131 VDD.n1130 40.824
R1442 VDD.n1151 VDD.n1150 40.824
R1443 VDD.n1212 VDD.n1211 40.824
R1444 VDD.n1232 VDD.n1231 40.824
R1445 VDD.n1293 VDD.n1292 40.824
R1446 VDD.n1313 VDD.n1312 40.824
R1447 VDD.n1374 VDD.n1373 40.824
R1448 VDD.n1394 VDD.n1393 40.824
R1449 VDD.n1455 VDD.n1454 40.824
R1450 VDD.n1475 VDD.n1474 40.824
R1451 VDD.n1536 VDD.n1535 40.824
R1452 VDD.n1556 VDD.n1555 40.824
R1453 VDD.n1617 VDD.n1616 40.824
R1454 VDD.n1637 VDD.n1636 40.824
R1455 VDD.n838 VDD.n837 40.824
R1456 VDD.n824 VDD.n823 40.824
R1457 VDD.n757 VDD.n756 40.824
R1458 VDD.n743 VDD.n742 40.824
R1459 VDD.n676 VDD.n675 40.824
R1460 VDD.n662 VDD.n661 40.824
R1461 VDD.n595 VDD.n594 40.824
R1462 VDD.n581 VDD.n580 40.824
R1463 VDD.n514 VDD.n513 40.824
R1464 VDD.n500 VDD.n499 40.824
R1465 VDD.n433 VDD.n432 40.824
R1466 VDD.n419 VDD.n418 40.824
R1467 VDD.n352 VDD.n351 40.824
R1468 VDD.n338 VDD.n337 40.824
R1469 VDD.n271 VDD.n270 40.824
R1470 VDD.n257 VDD.n256 40.824
R1471 VDD.n1013 VDD.n1012 36.774
R1472 VDD.n1094 VDD.n1093 36.774
R1473 VDD.n1175 VDD.n1174 36.774
R1474 VDD.n1256 VDD.n1255 36.774
R1475 VDD.n1337 VDD.n1336 36.774
R1476 VDD.n1418 VDD.n1417 36.774
R1477 VDD.n1499 VDD.n1498 36.774
R1478 VDD.n1580 VDD.n1579 36.774
R1479 VDD.n1661 VDD.n1660 36.774
R1480 VDD.n785 VDD.n784 36.774
R1481 VDD.n704 VDD.n703 36.774
R1482 VDD.n623 VDD.n622 36.774
R1483 VDD.n542 VDD.n541 36.774
R1484 VDD.n461 VDD.n460 36.774
R1485 VDD.n380 VDD.n379 36.774
R1486 VDD.n299 VDD.n298 36.774
R1487 VDD.n218 VDD.n217 36.774
R1488 VDD.n157 VDD.n156 36.774
R1489 VDD.n103 VDD.n102 36.774
R1490 VDD.n48 VDD.n47 36.774
R1491 VDD.n942 VDD.n941 36.774
R1492 VDD.n185 VDD.n184 36.608
R1493 VDD.n201 VDD.n200 32.032
R1494 VDD.n254 VDD.n253 27.456
R1495 VDD.n335 VDD.n334 27.456
R1496 VDD.n416 VDD.n415 27.456
R1497 VDD.n497 VDD.n496 27.456
R1498 VDD.n578 VDD.n577 27.456
R1499 VDD.n659 VDD.n658 27.456
R1500 VDD.n740 VDD.n739 27.456
R1501 VDD.n821 VDD.n820 27.456
R1502 VDD.n1634 VDD.n1633 27.456
R1503 VDD.n1553 VDD.n1552 27.456
R1504 VDD.n1472 VDD.n1471 27.456
R1505 VDD.n1391 VDD.n1390 27.456
R1506 VDD.n1310 VDD.n1309 27.456
R1507 VDD.n1229 VDD.n1228 27.456
R1508 VDD.n1148 VDD.n1147 27.456
R1509 VDD.n1067 VDD.n1066 27.456
R1510 VDD.n986 VDD.n985 27.456
R1511 VDD.n904 VDD.n903 27.456
R1512 VDD.n273 VDD.n272 22.88
R1513 VDD.n354 VDD.n353 22.88
R1514 VDD.n435 VDD.n434 22.88
R1515 VDD.n516 VDD.n515 22.88
R1516 VDD.n597 VDD.n596 22.88
R1517 VDD.n678 VDD.n677 22.88
R1518 VDD.n759 VDD.n758 22.88
R1519 VDD.n840 VDD.n839 22.88
R1520 VDD.n1619 VDD.n1618 22.88
R1521 VDD.n1538 VDD.n1537 22.88
R1522 VDD.n1457 VDD.n1456 22.88
R1523 VDD.n1376 VDD.n1375 22.88
R1524 VDD.n1295 VDD.n1294 22.88
R1525 VDD.n1214 VDD.n1213 22.88
R1526 VDD.n1133 VDD.n1132 22.88
R1527 VDD.n1052 VDD.n1051 22.88
R1528 VDD.n971 VDD.n970 22.88
R1529 VDD.n889 VDD.n888 22.88
R1530 VDD.n870 VDD.n867 21.841
R1531 VDD.n23 VDD.n20 21.841
R1532 VDD.n886 VDD.t40 14.282
R1533 VDD.n886 VDD.t68 14.282
R1534 VDD.n906 VDD.t87 14.282
R1535 VDD.n906 VDD.t80 14.282
R1536 VDD.n968 VDD.t18 14.282
R1537 VDD.n968 VDD.t64 14.282
R1538 VDD.n988 VDD.t5 14.282
R1539 VDD.n988 VDD.t11 14.282
R1540 VDD.n1049 VDD.t96 14.282
R1541 VDD.n1049 VDD.t102 14.282
R1542 VDD.n1069 VDD.t90 14.282
R1543 VDD.n1069 VDD.t112 14.282
R1544 VDD.n1130 VDD.t12 14.282
R1545 VDD.n1130 VDD.t69 14.282
R1546 VDD.n1150 VDD.t103 14.282
R1547 VDD.n1150 VDD.t10 14.282
R1548 VDD.n1211 VDD.t79 14.282
R1549 VDD.n1211 VDD.t44 14.282
R1550 VDD.n1231 VDD.t9 14.282
R1551 VDD.n1231 VDD.t6 14.282
R1552 VDD.n1292 VDD.t71 14.282
R1553 VDD.n1292 VDD.t1 14.282
R1554 VDD.n1312 VDD.t83 14.282
R1555 VDD.n1312 VDD.t91 14.282
R1556 VDD.n1373 VDD.t63 14.282
R1557 VDD.n1373 VDD.t54 14.282
R1558 VDD.n1393 VDD.t2 14.282
R1559 VDD.n1393 VDD.t84 14.282
R1560 VDD.n1454 VDD.t17 14.282
R1561 VDD.n1454 VDD.t55 14.282
R1562 VDD.n1474 VDD.t53 14.282
R1563 VDD.n1474 VDD.t19 14.282
R1564 VDD.n1535 VDD.t78 14.282
R1565 VDD.n1535 VDD.t58 14.282
R1566 VDD.n1555 VDD.t70 14.282
R1567 VDD.n1555 VDD.t82 14.282
R1568 VDD.n1616 VDD.t21 14.282
R1569 VDD.n1616 VDD.t109 14.282
R1570 VDD.n1636 VDD.t106 14.282
R1571 VDD.n1636 VDD.t20 14.282
R1572 VDD.n837 VDD.t48 14.282
R1573 VDD.n837 VDD.t110 14.282
R1574 VDD.n823 VDD.t62 14.282
R1575 VDD.n823 VDD.t105 14.282
R1576 VDD.n756 VDD.t3 14.282
R1577 VDD.n756 VDD.t93 14.282
R1578 VDD.n742 VDD.t8 14.282
R1579 VDD.n742 VDD.t77 14.282
R1580 VDD.n675 VDD.t66 14.282
R1581 VDD.n675 VDD.t86 14.282
R1582 VDD.n661 VDD.t36 14.282
R1583 VDD.n661 VDD.t7 14.282
R1584 VDD.n594 VDD.t15 14.282
R1585 VDD.n594 VDD.t42 14.282
R1586 VDD.n580 VDD.t29 14.282
R1587 VDD.n580 VDD.t16 14.282
R1588 VDD.n513 VDD.t51 14.282
R1589 VDD.n513 VDD.t99 14.282
R1590 VDD.n499 VDD.t32 14.282
R1591 VDD.n499 VDD.t76 14.282
R1592 VDD.n432 VDD.t14 14.282
R1593 VDD.n432 VDD.t47 14.282
R1594 VDD.n418 VDD.t24 14.282
R1595 VDD.n418 VDD.t13 14.282
R1596 VDD.n351 VDD.t23 14.282
R1597 VDD.n351 VDD.t35 14.282
R1598 VDD.n337 VDD.t65 14.282
R1599 VDD.n337 VDD.t85 14.282
R1600 VDD.n270 VDD.t97 14.282
R1601 VDD.n270 VDD.t41 14.282
R1602 VDD.n256 VDD.t31 14.282
R1603 VDD.n256 VDD.t94 14.282
R1604 VDD.n189 VDD.t59 14.282
R1605 VDD.n189 VDD.t38 14.282
R1606 VDD.n867 VDD.n850 14.167
R1607 VDD.n850 VDD.n849 14.167
R1608 VDD.n1028 VDD.n1010 14.167
R1609 VDD.n1010 VDD.n1009 14.167
R1610 VDD.n1109 VDD.n1091 14.167
R1611 VDD.n1091 VDD.n1090 14.167
R1612 VDD.n1190 VDD.n1172 14.167
R1613 VDD.n1172 VDD.n1171 14.167
R1614 VDD.n1271 VDD.n1253 14.167
R1615 VDD.n1253 VDD.n1252 14.167
R1616 VDD.n1352 VDD.n1334 14.167
R1617 VDD.n1334 VDD.n1333 14.167
R1618 VDD.n1433 VDD.n1415 14.167
R1619 VDD.n1415 VDD.n1414 14.167
R1620 VDD.n1514 VDD.n1496 14.167
R1621 VDD.n1496 VDD.n1495 14.167
R1622 VDD.n1595 VDD.n1577 14.167
R1623 VDD.n1577 VDD.n1576 14.167
R1624 VDD.n1676 VDD.n1658 14.167
R1625 VDD.n1658 VDD.n1657 14.167
R1626 VDD.n800 VDD.n782 14.167
R1627 VDD.n782 VDD.n781 14.167
R1628 VDD.n719 VDD.n701 14.167
R1629 VDD.n701 VDD.n700 14.167
R1630 VDD.n638 VDD.n620 14.167
R1631 VDD.n620 VDD.n619 14.167
R1632 VDD.n557 VDD.n539 14.167
R1633 VDD.n539 VDD.n538 14.167
R1634 VDD.n476 VDD.n458 14.167
R1635 VDD.n458 VDD.n457 14.167
R1636 VDD.n395 VDD.n377 14.167
R1637 VDD.n377 VDD.n376 14.167
R1638 VDD.n314 VDD.n296 14.167
R1639 VDD.n296 VDD.n295 14.167
R1640 VDD.n233 VDD.n215 14.167
R1641 VDD.n215 VDD.n214 14.167
R1642 VDD.n172 VDD.n154 14.167
R1643 VDD.n154 VDD.n153 14.167
R1644 VDD.n118 VDD.n100 14.167
R1645 VDD.n100 VDD.n99 14.167
R1646 VDD.n64 VDD.n45 14.167
R1647 VDD.n45 VDD.n44 14.167
R1648 VDD.n947 VDD.n928 14.167
R1649 VDD.n928 VDD.n927 14.167
R1650 VDD.n20 VDD.n19 14.167
R1651 VDD.n19 VDD.n17 14.167
R1652 VDD.n69 VDD.n65 14.167
R1653 VDD.n123 VDD.n119 14.167
R1654 VDD.n177 VDD.n173 14.167
R1655 VDD.n238 VDD.n234 14.167
R1656 VDD.n319 VDD.n315 14.167
R1657 VDD.n400 VDD.n396 14.167
R1658 VDD.n481 VDD.n477 14.167
R1659 VDD.n562 VDD.n558 14.167
R1660 VDD.n643 VDD.n639 14.167
R1661 VDD.n724 VDD.n720 14.167
R1662 VDD.n805 VDD.n801 14.167
R1663 VDD.n1681 VDD.n1677 14.167
R1664 VDD.n1600 VDD.n1596 14.167
R1665 VDD.n1519 VDD.n1515 14.167
R1666 VDD.n1438 VDD.n1434 14.167
R1667 VDD.n1357 VDD.n1353 14.167
R1668 VDD.n1276 VDD.n1272 14.167
R1669 VDD.n1195 VDD.n1191 14.167
R1670 VDD.n1114 VDD.n1110 14.167
R1671 VDD.n1033 VDD.n1029 14.167
R1672 VDD.n952 VDD.n948 14.167
R1673 VDD.n266 VDD.n265 13.728
R1674 VDD.n347 VDD.n346 13.728
R1675 VDD.n428 VDD.n427 13.728
R1676 VDD.n509 VDD.n508 13.728
R1677 VDD.n590 VDD.n589 13.728
R1678 VDD.n671 VDD.n670 13.728
R1679 VDD.n752 VDD.n751 13.728
R1680 VDD.n833 VDD.n832 13.728
R1681 VDD.n1624 VDD.n1623 13.728
R1682 VDD.n1543 VDD.n1542 13.728
R1683 VDD.n1462 VDD.n1461 13.728
R1684 VDD.n1381 VDD.n1380 13.728
R1685 VDD.n1300 VDD.n1299 13.728
R1686 VDD.n1219 VDD.n1218 13.728
R1687 VDD.n1138 VDD.n1137 13.728
R1688 VDD.n1057 VDD.n1056 13.728
R1689 VDD.n976 VDD.n975 13.728
R1690 VDD.n894 VDD.n893 13.728
R1691 VDD.n23 VDD.n22 13.653
R1692 VDD.n22 VDD.n21 13.653
R1693 VDD.n28 VDD.n27 13.653
R1694 VDD.n27 VDD.n26 13.653
R1695 VDD.n32 VDD.n31 13.653
R1696 VDD.n31 VDD.n30 13.653
R1697 VDD.n38 VDD.n36 13.653
R1698 VDD.n36 VDD.n35 13.653
R1699 VDD.n42 VDD.n41 13.653
R1700 VDD.n41 VDD.n40 13.653
R1701 VDD.n69 VDD.n68 13.653
R1702 VDD.n68 VDD.n67 13.653
R1703 VDD.n73 VDD.n72 13.653
R1704 VDD.n72 VDD.n71 13.653
R1705 VDD.n77 VDD.n76 13.653
R1706 VDD.n76 VDD.n75 13.653
R1707 VDD.n81 VDD.n80 13.653
R1708 VDD.n80 VDD.n79 13.653
R1709 VDD.n85 VDD.n84 13.653
R1710 VDD.n84 VDD.n83 13.653
R1711 VDD.n89 VDD.n88 13.653
R1712 VDD.n88 VDD.n87 13.653
R1713 VDD.n93 VDD.n92 13.653
R1714 VDD.n92 VDD.n91 13.653
R1715 VDD.n97 VDD.n96 13.653
R1716 VDD.n96 VDD.n95 13.653
R1717 VDD.n123 VDD.n122 13.653
R1718 VDD.n122 VDD.n121 13.653
R1719 VDD.n127 VDD.n126 13.653
R1720 VDD.n126 VDD.n125 13.653
R1721 VDD.n131 VDD.n130 13.653
R1722 VDD.n130 VDD.n129 13.653
R1723 VDD.n135 VDD.n134 13.653
R1724 VDD.n134 VDD.n133 13.653
R1725 VDD.n139 VDD.n138 13.653
R1726 VDD.n138 VDD.n137 13.653
R1727 VDD.n143 VDD.n142 13.653
R1728 VDD.n142 VDD.n141 13.653
R1729 VDD.n147 VDD.n146 13.653
R1730 VDD.n146 VDD.n145 13.653
R1731 VDD.n151 VDD.n150 13.653
R1732 VDD.n150 VDD.n149 13.653
R1733 VDD.n177 VDD.n176 13.653
R1734 VDD.n176 VDD.n175 13.653
R1735 VDD.n182 VDD.n181 13.653
R1736 VDD.n181 VDD.n180 13.653
R1737 VDD.n187 VDD.n186 13.653
R1738 VDD.n186 VDD.n185 13.653
R1739 VDD.n193 VDD.n192 13.653
R1740 VDD.n192 VDD.n191 13.653
R1741 VDD.n198 VDD.n197 13.653
R1742 VDD.n197 VDD.n196 13.653
R1743 VDD.n203 VDD.n202 13.653
R1744 VDD.n202 VDD.n201 13.653
R1745 VDD.n208 VDD.n207 13.653
R1746 VDD.n207 VDD.n206 13.653
R1747 VDD.n212 VDD.n211 13.653
R1748 VDD.n211 VDD.n210 13.653
R1749 VDD.n238 VDD.n237 13.653
R1750 VDD.n237 VDD.n236 13.653
R1751 VDD.n242 VDD.n241 13.653
R1752 VDD.n241 VDD.n240 13.653
R1753 VDD.n246 VDD.n245 13.653
R1754 VDD.n245 VDD.n244 13.653
R1755 VDD.n251 VDD.n250 13.653
R1756 VDD.n250 VDD.n249 13.653
R1757 VDD.n258 VDD.n255 13.653
R1758 VDD.n255 VDD.n254 13.653
R1759 VDD.n263 VDD.n262 13.653
R1760 VDD.n262 VDD.n261 13.653
R1761 VDD.n268 VDD.n267 13.653
R1762 VDD.n267 VDD.n266 13.653
R1763 VDD.n275 VDD.n274 13.653
R1764 VDD.n274 VDD.n273 13.653
R1765 VDD.n280 VDD.n279 13.653
R1766 VDD.n279 VDD.n278 13.653
R1767 VDD.n285 VDD.n284 13.653
R1768 VDD.n284 VDD.n283 13.653
R1769 VDD.n289 VDD.n288 13.653
R1770 VDD.n288 VDD.n287 13.653
R1771 VDD.n293 VDD.n292 13.653
R1772 VDD.n292 VDD.n291 13.653
R1773 VDD.n319 VDD.n318 13.653
R1774 VDD.n318 VDD.n317 13.653
R1775 VDD.n323 VDD.n322 13.653
R1776 VDD.n322 VDD.n321 13.653
R1777 VDD.n327 VDD.n326 13.653
R1778 VDD.n326 VDD.n325 13.653
R1779 VDD.n332 VDD.n331 13.653
R1780 VDD.n331 VDD.n330 13.653
R1781 VDD.n339 VDD.n336 13.653
R1782 VDD.n336 VDD.n335 13.653
R1783 VDD.n344 VDD.n343 13.653
R1784 VDD.n343 VDD.n342 13.653
R1785 VDD.n349 VDD.n348 13.653
R1786 VDD.n348 VDD.n347 13.653
R1787 VDD.n356 VDD.n355 13.653
R1788 VDD.n355 VDD.n354 13.653
R1789 VDD.n361 VDD.n360 13.653
R1790 VDD.n360 VDD.n359 13.653
R1791 VDD.n366 VDD.n365 13.653
R1792 VDD.n365 VDD.n364 13.653
R1793 VDD.n370 VDD.n369 13.653
R1794 VDD.n369 VDD.n368 13.653
R1795 VDD.n374 VDD.n373 13.653
R1796 VDD.n373 VDD.n372 13.653
R1797 VDD.n400 VDD.n399 13.653
R1798 VDD.n399 VDD.n398 13.653
R1799 VDD.n404 VDD.n403 13.653
R1800 VDD.n403 VDD.n402 13.653
R1801 VDD.n408 VDD.n407 13.653
R1802 VDD.n407 VDD.n406 13.653
R1803 VDD.n413 VDD.n412 13.653
R1804 VDD.n412 VDD.n411 13.653
R1805 VDD.n420 VDD.n417 13.653
R1806 VDD.n417 VDD.n416 13.653
R1807 VDD.n425 VDD.n424 13.653
R1808 VDD.n424 VDD.n423 13.653
R1809 VDD.n430 VDD.n429 13.653
R1810 VDD.n429 VDD.n428 13.653
R1811 VDD.n437 VDD.n436 13.653
R1812 VDD.n436 VDD.n435 13.653
R1813 VDD.n442 VDD.n441 13.653
R1814 VDD.n441 VDD.n440 13.653
R1815 VDD.n447 VDD.n446 13.653
R1816 VDD.n446 VDD.n445 13.653
R1817 VDD.n451 VDD.n450 13.653
R1818 VDD.n450 VDD.n449 13.653
R1819 VDD.n455 VDD.n454 13.653
R1820 VDD.n454 VDD.n453 13.653
R1821 VDD.n481 VDD.n480 13.653
R1822 VDD.n480 VDD.n479 13.653
R1823 VDD.n485 VDD.n484 13.653
R1824 VDD.n484 VDD.n483 13.653
R1825 VDD.n489 VDD.n488 13.653
R1826 VDD.n488 VDD.n487 13.653
R1827 VDD.n494 VDD.n493 13.653
R1828 VDD.n493 VDD.n492 13.653
R1829 VDD.n501 VDD.n498 13.653
R1830 VDD.n498 VDD.n497 13.653
R1831 VDD.n506 VDD.n505 13.653
R1832 VDD.n505 VDD.n504 13.653
R1833 VDD.n511 VDD.n510 13.653
R1834 VDD.n510 VDD.n509 13.653
R1835 VDD.n518 VDD.n517 13.653
R1836 VDD.n517 VDD.n516 13.653
R1837 VDD.n523 VDD.n522 13.653
R1838 VDD.n522 VDD.n521 13.653
R1839 VDD.n528 VDD.n527 13.653
R1840 VDD.n527 VDD.n526 13.653
R1841 VDD.n532 VDD.n531 13.653
R1842 VDD.n531 VDD.n530 13.653
R1843 VDD.n536 VDD.n535 13.653
R1844 VDD.n535 VDD.n534 13.653
R1845 VDD.n562 VDD.n561 13.653
R1846 VDD.n561 VDD.n560 13.653
R1847 VDD.n566 VDD.n565 13.653
R1848 VDD.n565 VDD.n564 13.653
R1849 VDD.n570 VDD.n569 13.653
R1850 VDD.n569 VDD.n568 13.653
R1851 VDD.n575 VDD.n574 13.653
R1852 VDD.n574 VDD.n573 13.653
R1853 VDD.n582 VDD.n579 13.653
R1854 VDD.n579 VDD.n578 13.653
R1855 VDD.n587 VDD.n586 13.653
R1856 VDD.n586 VDD.n585 13.653
R1857 VDD.n592 VDD.n591 13.653
R1858 VDD.n591 VDD.n590 13.653
R1859 VDD.n599 VDD.n598 13.653
R1860 VDD.n598 VDD.n597 13.653
R1861 VDD.n604 VDD.n603 13.653
R1862 VDD.n603 VDD.n602 13.653
R1863 VDD.n609 VDD.n608 13.653
R1864 VDD.n608 VDD.n607 13.653
R1865 VDD.n613 VDD.n612 13.653
R1866 VDD.n612 VDD.n611 13.653
R1867 VDD.n617 VDD.n616 13.653
R1868 VDD.n616 VDD.n615 13.653
R1869 VDD.n643 VDD.n642 13.653
R1870 VDD.n642 VDD.n641 13.653
R1871 VDD.n647 VDD.n646 13.653
R1872 VDD.n646 VDD.n645 13.653
R1873 VDD.n651 VDD.n650 13.653
R1874 VDD.n650 VDD.n649 13.653
R1875 VDD.n656 VDD.n655 13.653
R1876 VDD.n655 VDD.n654 13.653
R1877 VDD.n663 VDD.n660 13.653
R1878 VDD.n660 VDD.n659 13.653
R1879 VDD.n668 VDD.n667 13.653
R1880 VDD.n667 VDD.n666 13.653
R1881 VDD.n673 VDD.n672 13.653
R1882 VDD.n672 VDD.n671 13.653
R1883 VDD.n680 VDD.n679 13.653
R1884 VDD.n679 VDD.n678 13.653
R1885 VDD.n685 VDD.n684 13.653
R1886 VDD.n684 VDD.n683 13.653
R1887 VDD.n690 VDD.n689 13.653
R1888 VDD.n689 VDD.n688 13.653
R1889 VDD.n694 VDD.n693 13.653
R1890 VDD.n693 VDD.n692 13.653
R1891 VDD.n698 VDD.n697 13.653
R1892 VDD.n697 VDD.n696 13.653
R1893 VDD.n724 VDD.n723 13.653
R1894 VDD.n723 VDD.n722 13.653
R1895 VDD.n728 VDD.n727 13.653
R1896 VDD.n727 VDD.n726 13.653
R1897 VDD.n732 VDD.n731 13.653
R1898 VDD.n731 VDD.n730 13.653
R1899 VDD.n737 VDD.n736 13.653
R1900 VDD.n736 VDD.n735 13.653
R1901 VDD.n744 VDD.n741 13.653
R1902 VDD.n741 VDD.n740 13.653
R1903 VDD.n749 VDD.n748 13.653
R1904 VDD.n748 VDD.n747 13.653
R1905 VDD.n754 VDD.n753 13.653
R1906 VDD.n753 VDD.n752 13.653
R1907 VDD.n761 VDD.n760 13.653
R1908 VDD.n760 VDD.n759 13.653
R1909 VDD.n766 VDD.n765 13.653
R1910 VDD.n765 VDD.n764 13.653
R1911 VDD.n771 VDD.n770 13.653
R1912 VDD.n770 VDD.n769 13.653
R1913 VDD.n775 VDD.n774 13.653
R1914 VDD.n774 VDD.n773 13.653
R1915 VDD.n779 VDD.n778 13.653
R1916 VDD.n778 VDD.n777 13.653
R1917 VDD.n805 VDD.n804 13.653
R1918 VDD.n804 VDD.n803 13.653
R1919 VDD.n809 VDD.n808 13.653
R1920 VDD.n808 VDD.n807 13.653
R1921 VDD.n813 VDD.n812 13.653
R1922 VDD.n812 VDD.n811 13.653
R1923 VDD.n818 VDD.n817 13.653
R1924 VDD.n817 VDD.n816 13.653
R1925 VDD.n825 VDD.n822 13.653
R1926 VDD.n822 VDD.n821 13.653
R1927 VDD.n830 VDD.n829 13.653
R1928 VDD.n829 VDD.n828 13.653
R1929 VDD.n835 VDD.n834 13.653
R1930 VDD.n834 VDD.n833 13.653
R1931 VDD.n842 VDD.n841 13.653
R1932 VDD.n841 VDD.n840 13.653
R1933 VDD.n847 VDD.n846 13.653
R1934 VDD.n846 VDD.n845 13.653
R1935 VDD.n1690 VDD.n1689 13.653
R1936 VDD.n1689 VDD.n1688 13.653
R1937 VDD.n1685 VDD.n1684 13.653
R1938 VDD.n1684 VDD.n1683 13.653
R1939 VDD.n1681 VDD.n1680 13.653
R1940 VDD.n1680 VDD.n1679 13.653
R1941 VDD.n1655 VDD.n1654 13.653
R1942 VDD.n1654 VDD.n1653 13.653
R1943 VDD.n1651 VDD.n1650 13.653
R1944 VDD.n1650 VDD.n1649 13.653
R1945 VDD.n1647 VDD.n1646 13.653
R1946 VDD.n1646 VDD.n1645 13.653
R1947 VDD.n1643 VDD.n1642 13.653
R1948 VDD.n1642 VDD.n1641 13.653
R1949 VDD.n1638 VDD.n1635 13.653
R1950 VDD.n1635 VDD.n1634 13.653
R1951 VDD.n1631 VDD.n1630 13.653
R1952 VDD.n1630 VDD.n1629 13.653
R1953 VDD.n1626 VDD.n1625 13.653
R1954 VDD.n1625 VDD.n1624 13.653
R1955 VDD.n1621 VDD.n1620 13.653
R1956 VDD.n1620 VDD.n1619 13.653
R1957 VDD.n1614 VDD.n1613 13.653
R1958 VDD.n1613 VDD.n1612 13.653
R1959 VDD.n1609 VDD.n1608 13.653
R1960 VDD.n1608 VDD.n1607 13.653
R1961 VDD.n1604 VDD.n1603 13.653
R1962 VDD.n1603 VDD.n1602 13.653
R1963 VDD.n1600 VDD.n1599 13.653
R1964 VDD.n1599 VDD.n1598 13.653
R1965 VDD.n1574 VDD.n1573 13.653
R1966 VDD.n1573 VDD.n1572 13.653
R1967 VDD.n1570 VDD.n1569 13.653
R1968 VDD.n1569 VDD.n1568 13.653
R1969 VDD.n1566 VDD.n1565 13.653
R1970 VDD.n1565 VDD.n1564 13.653
R1971 VDD.n1562 VDD.n1561 13.653
R1972 VDD.n1561 VDD.n1560 13.653
R1973 VDD.n1557 VDD.n1554 13.653
R1974 VDD.n1554 VDD.n1553 13.653
R1975 VDD.n1550 VDD.n1549 13.653
R1976 VDD.n1549 VDD.n1548 13.653
R1977 VDD.n1545 VDD.n1544 13.653
R1978 VDD.n1544 VDD.n1543 13.653
R1979 VDD.n1540 VDD.n1539 13.653
R1980 VDD.n1539 VDD.n1538 13.653
R1981 VDD.n1533 VDD.n1532 13.653
R1982 VDD.n1532 VDD.n1531 13.653
R1983 VDD.n1528 VDD.n1527 13.653
R1984 VDD.n1527 VDD.n1526 13.653
R1985 VDD.n1523 VDD.n1522 13.653
R1986 VDD.n1522 VDD.n1521 13.653
R1987 VDD.n1519 VDD.n1518 13.653
R1988 VDD.n1518 VDD.n1517 13.653
R1989 VDD.n1493 VDD.n1492 13.653
R1990 VDD.n1492 VDD.n1491 13.653
R1991 VDD.n1489 VDD.n1488 13.653
R1992 VDD.n1488 VDD.n1487 13.653
R1993 VDD.n1485 VDD.n1484 13.653
R1994 VDD.n1484 VDD.n1483 13.653
R1995 VDD.n1481 VDD.n1480 13.653
R1996 VDD.n1480 VDD.n1479 13.653
R1997 VDD.n1476 VDD.n1473 13.653
R1998 VDD.n1473 VDD.n1472 13.653
R1999 VDD.n1469 VDD.n1468 13.653
R2000 VDD.n1468 VDD.n1467 13.653
R2001 VDD.n1464 VDD.n1463 13.653
R2002 VDD.n1463 VDD.n1462 13.653
R2003 VDD.n1459 VDD.n1458 13.653
R2004 VDD.n1458 VDD.n1457 13.653
R2005 VDD.n1452 VDD.n1451 13.653
R2006 VDD.n1451 VDD.n1450 13.653
R2007 VDD.n1447 VDD.n1446 13.653
R2008 VDD.n1446 VDD.n1445 13.653
R2009 VDD.n1442 VDD.n1441 13.653
R2010 VDD.n1441 VDD.n1440 13.653
R2011 VDD.n1438 VDD.n1437 13.653
R2012 VDD.n1437 VDD.n1436 13.653
R2013 VDD.n1412 VDD.n1411 13.653
R2014 VDD.n1411 VDD.n1410 13.653
R2015 VDD.n1408 VDD.n1407 13.653
R2016 VDD.n1407 VDD.n1406 13.653
R2017 VDD.n1404 VDD.n1403 13.653
R2018 VDD.n1403 VDD.n1402 13.653
R2019 VDD.n1400 VDD.n1399 13.653
R2020 VDD.n1399 VDD.n1398 13.653
R2021 VDD.n1395 VDD.n1392 13.653
R2022 VDD.n1392 VDD.n1391 13.653
R2023 VDD.n1388 VDD.n1387 13.653
R2024 VDD.n1387 VDD.n1386 13.653
R2025 VDD.n1383 VDD.n1382 13.653
R2026 VDD.n1382 VDD.n1381 13.653
R2027 VDD.n1378 VDD.n1377 13.653
R2028 VDD.n1377 VDD.n1376 13.653
R2029 VDD.n1371 VDD.n1370 13.653
R2030 VDD.n1370 VDD.n1369 13.653
R2031 VDD.n1366 VDD.n1365 13.653
R2032 VDD.n1365 VDD.n1364 13.653
R2033 VDD.n1361 VDD.n1360 13.653
R2034 VDD.n1360 VDD.n1359 13.653
R2035 VDD.n1357 VDD.n1356 13.653
R2036 VDD.n1356 VDD.n1355 13.653
R2037 VDD.n1331 VDD.n1330 13.653
R2038 VDD.n1330 VDD.n1329 13.653
R2039 VDD.n1327 VDD.n1326 13.653
R2040 VDD.n1326 VDD.n1325 13.653
R2041 VDD.n1323 VDD.n1322 13.653
R2042 VDD.n1322 VDD.n1321 13.653
R2043 VDD.n1319 VDD.n1318 13.653
R2044 VDD.n1318 VDD.n1317 13.653
R2045 VDD.n1314 VDD.n1311 13.653
R2046 VDD.n1311 VDD.n1310 13.653
R2047 VDD.n1307 VDD.n1306 13.653
R2048 VDD.n1306 VDD.n1305 13.653
R2049 VDD.n1302 VDD.n1301 13.653
R2050 VDD.n1301 VDD.n1300 13.653
R2051 VDD.n1297 VDD.n1296 13.653
R2052 VDD.n1296 VDD.n1295 13.653
R2053 VDD.n1290 VDD.n1289 13.653
R2054 VDD.n1289 VDD.n1288 13.653
R2055 VDD.n1285 VDD.n1284 13.653
R2056 VDD.n1284 VDD.n1283 13.653
R2057 VDD.n1280 VDD.n1279 13.653
R2058 VDD.n1279 VDD.n1278 13.653
R2059 VDD.n1276 VDD.n1275 13.653
R2060 VDD.n1275 VDD.n1274 13.653
R2061 VDD.n1250 VDD.n1249 13.653
R2062 VDD.n1249 VDD.n1248 13.653
R2063 VDD.n1246 VDD.n1245 13.653
R2064 VDD.n1245 VDD.n1244 13.653
R2065 VDD.n1242 VDD.n1241 13.653
R2066 VDD.n1241 VDD.n1240 13.653
R2067 VDD.n1238 VDD.n1237 13.653
R2068 VDD.n1237 VDD.n1236 13.653
R2069 VDD.n1233 VDD.n1230 13.653
R2070 VDD.n1230 VDD.n1229 13.653
R2071 VDD.n1226 VDD.n1225 13.653
R2072 VDD.n1225 VDD.n1224 13.653
R2073 VDD.n1221 VDD.n1220 13.653
R2074 VDD.n1220 VDD.n1219 13.653
R2075 VDD.n1216 VDD.n1215 13.653
R2076 VDD.n1215 VDD.n1214 13.653
R2077 VDD.n1209 VDD.n1208 13.653
R2078 VDD.n1208 VDD.n1207 13.653
R2079 VDD.n1204 VDD.n1203 13.653
R2080 VDD.n1203 VDD.n1202 13.653
R2081 VDD.n1199 VDD.n1198 13.653
R2082 VDD.n1198 VDD.n1197 13.653
R2083 VDD.n1195 VDD.n1194 13.653
R2084 VDD.n1194 VDD.n1193 13.653
R2085 VDD.n1169 VDD.n1168 13.653
R2086 VDD.n1168 VDD.n1167 13.653
R2087 VDD.n1165 VDD.n1164 13.653
R2088 VDD.n1164 VDD.n1163 13.653
R2089 VDD.n1161 VDD.n1160 13.653
R2090 VDD.n1160 VDD.n1159 13.653
R2091 VDD.n1157 VDD.n1156 13.653
R2092 VDD.n1156 VDD.n1155 13.653
R2093 VDD.n1152 VDD.n1149 13.653
R2094 VDD.n1149 VDD.n1148 13.653
R2095 VDD.n1145 VDD.n1144 13.653
R2096 VDD.n1144 VDD.n1143 13.653
R2097 VDD.n1140 VDD.n1139 13.653
R2098 VDD.n1139 VDD.n1138 13.653
R2099 VDD.n1135 VDD.n1134 13.653
R2100 VDD.n1134 VDD.n1133 13.653
R2101 VDD.n1128 VDD.n1127 13.653
R2102 VDD.n1127 VDD.n1126 13.653
R2103 VDD.n1123 VDD.n1122 13.653
R2104 VDD.n1122 VDD.n1121 13.653
R2105 VDD.n1118 VDD.n1117 13.653
R2106 VDD.n1117 VDD.n1116 13.653
R2107 VDD.n1114 VDD.n1113 13.653
R2108 VDD.n1113 VDD.n1112 13.653
R2109 VDD.n1088 VDD.n1087 13.653
R2110 VDD.n1087 VDD.n1086 13.653
R2111 VDD.n1084 VDD.n1083 13.653
R2112 VDD.n1083 VDD.n1082 13.653
R2113 VDD.n1080 VDD.n1079 13.653
R2114 VDD.n1079 VDD.n1078 13.653
R2115 VDD.n1076 VDD.n1075 13.653
R2116 VDD.n1075 VDD.n1074 13.653
R2117 VDD.n1071 VDD.n1068 13.653
R2118 VDD.n1068 VDD.n1067 13.653
R2119 VDD.n1064 VDD.n1063 13.653
R2120 VDD.n1063 VDD.n1062 13.653
R2121 VDD.n1059 VDD.n1058 13.653
R2122 VDD.n1058 VDD.n1057 13.653
R2123 VDD.n1054 VDD.n1053 13.653
R2124 VDD.n1053 VDD.n1052 13.653
R2125 VDD.n1047 VDD.n1046 13.653
R2126 VDD.n1046 VDD.n1045 13.653
R2127 VDD.n1042 VDD.n1041 13.653
R2128 VDD.n1041 VDD.n1040 13.653
R2129 VDD.n1037 VDD.n1036 13.653
R2130 VDD.n1036 VDD.n1035 13.653
R2131 VDD.n1033 VDD.n1032 13.653
R2132 VDD.n1032 VDD.n1031 13.653
R2133 VDD.n1007 VDD.n1006 13.653
R2134 VDD.n1006 VDD.n1005 13.653
R2135 VDD.n1003 VDD.n1002 13.653
R2136 VDD.n1002 VDD.n1001 13.653
R2137 VDD.n999 VDD.n998 13.653
R2138 VDD.n998 VDD.n997 13.653
R2139 VDD.n995 VDD.n994 13.653
R2140 VDD.n994 VDD.n993 13.653
R2141 VDD.n990 VDD.n987 13.653
R2142 VDD.n987 VDD.n986 13.653
R2143 VDD.n983 VDD.n982 13.653
R2144 VDD.n982 VDD.n981 13.653
R2145 VDD.n978 VDD.n977 13.653
R2146 VDD.n977 VDD.n976 13.653
R2147 VDD.n973 VDD.n972 13.653
R2148 VDD.n972 VDD.n971 13.653
R2149 VDD.n966 VDD.n965 13.653
R2150 VDD.n965 VDD.n964 13.653
R2151 VDD.n961 VDD.n960 13.653
R2152 VDD.n960 VDD.n959 13.653
R2153 VDD.n956 VDD.n955 13.653
R2154 VDD.n955 VDD.n954 13.653
R2155 VDD.n952 VDD.n951 13.653
R2156 VDD.n951 VDD.n950 13.653
R2157 VDD.n925 VDD.n924 13.653
R2158 VDD.n924 VDD.n923 13.653
R2159 VDD.n921 VDD.n920 13.653
R2160 VDD.n920 VDD.n919 13.653
R2161 VDD.n917 VDD.n916 13.653
R2162 VDD.n916 VDD.n915 13.653
R2163 VDD.n913 VDD.n912 13.653
R2164 VDD.n912 VDD.n911 13.653
R2165 VDD.n908 VDD.n905 13.653
R2166 VDD.n905 VDD.n904 13.653
R2167 VDD.n901 VDD.n900 13.653
R2168 VDD.n900 VDD.n899 13.653
R2169 VDD.n896 VDD.n895 13.653
R2170 VDD.n895 VDD.n894 13.653
R2171 VDD.n891 VDD.n890 13.653
R2172 VDD.n890 VDD.n889 13.653
R2173 VDD.n884 VDD.n883 13.653
R2174 VDD.n883 VDD.n882 13.653
R2175 VDD.n879 VDD.n878 13.653
R2176 VDD.n878 VDD.n877 13.653
R2177 VDD.n874 VDD.n873 13.653
R2178 VDD.n873 VDD.n872 13.653
R2179 VDD.n870 VDD.n869 13.653
R2180 VDD.n869 VDD.n868 13.653
R2181 VDD.n4 VDD.n2 12.915
R2182 VDD.n4 VDD.n3 12.66
R2183 VDD.n12 VDD.n11 12.343
R2184 VDD.n12 VDD.n9 12.343
R2185 VDD.n7 VDD.n6 12.343
R2186 VDD.n261 VDD.n260 9.152
R2187 VDD.n342 VDD.n341 9.152
R2188 VDD.n423 VDD.n422 9.152
R2189 VDD.n504 VDD.n503 9.152
R2190 VDD.n585 VDD.n584 9.152
R2191 VDD.n666 VDD.n665 9.152
R2192 VDD.n747 VDD.n746 9.152
R2193 VDD.n828 VDD.n827 9.152
R2194 VDD.n1629 VDD.n1628 9.152
R2195 VDD.n1548 VDD.n1547 9.152
R2196 VDD.n1467 VDD.n1466 9.152
R2197 VDD.n1386 VDD.n1385 9.152
R2198 VDD.n1305 VDD.n1304 9.152
R2199 VDD.n1224 VDD.n1223 9.152
R2200 VDD.n1143 VDD.n1142 9.152
R2201 VDD.n1062 VDD.n1061 9.152
R2202 VDD.n981 VDD.n980 9.152
R2203 VDD.n899 VDD.n898 9.152
R2204 VDD.n193 VDD.n190 8.658
R2205 VDD.n1029 VDD.n1028 7.674
R2206 VDD.n1110 VDD.n1109 7.674
R2207 VDD.n1191 VDD.n1190 7.674
R2208 VDD.n1272 VDD.n1271 7.674
R2209 VDD.n1353 VDD.n1352 7.674
R2210 VDD.n1434 VDD.n1433 7.674
R2211 VDD.n1515 VDD.n1514 7.674
R2212 VDD.n1596 VDD.n1595 7.674
R2213 VDD.n1677 VDD.n1676 7.674
R2214 VDD.n801 VDD.n800 7.674
R2215 VDD.n720 VDD.n719 7.674
R2216 VDD.n639 VDD.n638 7.674
R2217 VDD.n558 VDD.n557 7.674
R2218 VDD.n477 VDD.n476 7.674
R2219 VDD.n396 VDD.n395 7.674
R2220 VDD.n315 VDD.n314 7.674
R2221 VDD.n234 VDD.n233 7.674
R2222 VDD.n173 VDD.n172 7.674
R2223 VDD.n119 VDD.n118 7.674
R2224 VDD.n65 VDD.n64 7.674
R2225 VDD.n948 VDD.n947 7.674
R2226 VDD.n59 VDD.n58 7.5
R2227 VDD.n53 VDD.n52 7.5
R2228 VDD.n55 VDD.n54 7.5
R2229 VDD.n50 VDD.n49 7.5
R2230 VDD.n64 VDD.n63 7.5
R2231 VDD.n113 VDD.n112 7.5
R2232 VDD.n107 VDD.n106 7.5
R2233 VDD.n109 VDD.n108 7.5
R2234 VDD.n115 VDD.n105 7.5
R2235 VDD.n115 VDD.n103 7.5
R2236 VDD.n118 VDD.n117 7.5
R2237 VDD.n167 VDD.n166 7.5
R2238 VDD.n161 VDD.n160 7.5
R2239 VDD.n163 VDD.n162 7.5
R2240 VDD.n169 VDD.n159 7.5
R2241 VDD.n169 VDD.n157 7.5
R2242 VDD.n172 VDD.n171 7.5
R2243 VDD.n228 VDD.n227 7.5
R2244 VDD.n222 VDD.n221 7.5
R2245 VDD.n224 VDD.n223 7.5
R2246 VDD.n230 VDD.n220 7.5
R2247 VDD.n230 VDD.n218 7.5
R2248 VDD.n233 VDD.n232 7.5
R2249 VDD.n309 VDD.n308 7.5
R2250 VDD.n303 VDD.n302 7.5
R2251 VDD.n305 VDD.n304 7.5
R2252 VDD.n311 VDD.n301 7.5
R2253 VDD.n311 VDD.n299 7.5
R2254 VDD.n314 VDD.n313 7.5
R2255 VDD.n390 VDD.n389 7.5
R2256 VDD.n384 VDD.n383 7.5
R2257 VDD.n386 VDD.n385 7.5
R2258 VDD.n392 VDD.n382 7.5
R2259 VDD.n392 VDD.n380 7.5
R2260 VDD.n395 VDD.n394 7.5
R2261 VDD.n471 VDD.n470 7.5
R2262 VDD.n465 VDD.n464 7.5
R2263 VDD.n467 VDD.n466 7.5
R2264 VDD.n473 VDD.n463 7.5
R2265 VDD.n473 VDD.n461 7.5
R2266 VDD.n476 VDD.n475 7.5
R2267 VDD.n552 VDD.n551 7.5
R2268 VDD.n546 VDD.n545 7.5
R2269 VDD.n548 VDD.n547 7.5
R2270 VDD.n554 VDD.n544 7.5
R2271 VDD.n554 VDD.n542 7.5
R2272 VDD.n557 VDD.n556 7.5
R2273 VDD.n633 VDD.n632 7.5
R2274 VDD.n627 VDD.n626 7.5
R2275 VDD.n629 VDD.n628 7.5
R2276 VDD.n635 VDD.n625 7.5
R2277 VDD.n635 VDD.n623 7.5
R2278 VDD.n638 VDD.n637 7.5
R2279 VDD.n714 VDD.n713 7.5
R2280 VDD.n708 VDD.n707 7.5
R2281 VDD.n710 VDD.n709 7.5
R2282 VDD.n716 VDD.n706 7.5
R2283 VDD.n716 VDD.n704 7.5
R2284 VDD.n719 VDD.n718 7.5
R2285 VDD.n795 VDD.n794 7.5
R2286 VDD.n789 VDD.n788 7.5
R2287 VDD.n791 VDD.n790 7.5
R2288 VDD.n797 VDD.n787 7.5
R2289 VDD.n797 VDD.n785 7.5
R2290 VDD.n800 VDD.n799 7.5
R2291 VDD.n1671 VDD.n1670 7.5
R2292 VDD.n1665 VDD.n1664 7.5
R2293 VDD.n1667 VDD.n1666 7.5
R2294 VDD.n1673 VDD.n1663 7.5
R2295 VDD.n1673 VDD.n1661 7.5
R2296 VDD.n1676 VDD.n1675 7.5
R2297 VDD.n1590 VDD.n1589 7.5
R2298 VDD.n1584 VDD.n1583 7.5
R2299 VDD.n1586 VDD.n1585 7.5
R2300 VDD.n1592 VDD.n1582 7.5
R2301 VDD.n1592 VDD.n1580 7.5
R2302 VDD.n1595 VDD.n1594 7.5
R2303 VDD.n1509 VDD.n1508 7.5
R2304 VDD.n1503 VDD.n1502 7.5
R2305 VDD.n1505 VDD.n1504 7.5
R2306 VDD.n1511 VDD.n1501 7.5
R2307 VDD.n1511 VDD.n1499 7.5
R2308 VDD.n1514 VDD.n1513 7.5
R2309 VDD.n1428 VDD.n1427 7.5
R2310 VDD.n1422 VDD.n1421 7.5
R2311 VDD.n1424 VDD.n1423 7.5
R2312 VDD.n1430 VDD.n1420 7.5
R2313 VDD.n1430 VDD.n1418 7.5
R2314 VDD.n1433 VDD.n1432 7.5
R2315 VDD.n1347 VDD.n1346 7.5
R2316 VDD.n1341 VDD.n1340 7.5
R2317 VDD.n1343 VDD.n1342 7.5
R2318 VDD.n1349 VDD.n1339 7.5
R2319 VDD.n1349 VDD.n1337 7.5
R2320 VDD.n1352 VDD.n1351 7.5
R2321 VDD.n1266 VDD.n1265 7.5
R2322 VDD.n1260 VDD.n1259 7.5
R2323 VDD.n1262 VDD.n1261 7.5
R2324 VDD.n1268 VDD.n1258 7.5
R2325 VDD.n1268 VDD.n1256 7.5
R2326 VDD.n1271 VDD.n1270 7.5
R2327 VDD.n1185 VDD.n1184 7.5
R2328 VDD.n1179 VDD.n1178 7.5
R2329 VDD.n1181 VDD.n1180 7.5
R2330 VDD.n1187 VDD.n1177 7.5
R2331 VDD.n1187 VDD.n1175 7.5
R2332 VDD.n1190 VDD.n1189 7.5
R2333 VDD.n1104 VDD.n1103 7.5
R2334 VDD.n1098 VDD.n1097 7.5
R2335 VDD.n1100 VDD.n1099 7.5
R2336 VDD.n1106 VDD.n1096 7.5
R2337 VDD.n1106 VDD.n1094 7.5
R2338 VDD.n1109 VDD.n1108 7.5
R2339 VDD.n1023 VDD.n1022 7.5
R2340 VDD.n1017 VDD.n1016 7.5
R2341 VDD.n1019 VDD.n1018 7.5
R2342 VDD.n1025 VDD.n1015 7.5
R2343 VDD.n1025 VDD.n1013 7.5
R2344 VDD.n1028 VDD.n1027 7.5
R2345 VDD.n932 VDD.n931 7.5
R2346 VDD.n935 VDD.n934 7.5
R2347 VDD.n937 VDD.n936 7.5
R2348 VDD.n940 VDD.n939 7.5
R2349 VDD.n947 VDD.n946 7.5
R2350 VDD.n862 VDD.n861 7.5
R2351 VDD.n856 VDD.n855 7.5
R2352 VDD.n858 VDD.n857 7.5
R2353 VDD.n864 VDD.n854 7.5
R2354 VDD.n864 VDD.n852 7.5
R2355 VDD.n867 VDD.n866 7.5
R2356 VDD.n20 VDD.n16 7.5
R2357 VDD.n2 VDD.n1 7.5
R2358 VDD.n6 VDD.n5 7.5
R2359 VDD.n11 VDD.n10 7.5
R2360 VDD.n19 VDD.n18 7.5
R2361 VDD.n14 VDD.n0 7.5
R2362 VDD.n51 VDD.n48 6.772
R2363 VDD.n62 VDD.n46 6.772
R2364 VDD.n60 VDD.n57 6.772
R2365 VDD.n56 VDD.n53 6.772
R2366 VDD.n116 VDD.n101 6.772
R2367 VDD.n114 VDD.n111 6.772
R2368 VDD.n110 VDD.n107 6.772
R2369 VDD.n170 VDD.n155 6.772
R2370 VDD.n168 VDD.n165 6.772
R2371 VDD.n164 VDD.n161 6.772
R2372 VDD.n231 VDD.n216 6.772
R2373 VDD.n229 VDD.n226 6.772
R2374 VDD.n225 VDD.n222 6.772
R2375 VDD.n312 VDD.n297 6.772
R2376 VDD.n310 VDD.n307 6.772
R2377 VDD.n306 VDD.n303 6.772
R2378 VDD.n393 VDD.n378 6.772
R2379 VDD.n391 VDD.n388 6.772
R2380 VDD.n387 VDD.n384 6.772
R2381 VDD.n474 VDD.n459 6.772
R2382 VDD.n472 VDD.n469 6.772
R2383 VDD.n468 VDD.n465 6.772
R2384 VDD.n555 VDD.n540 6.772
R2385 VDD.n553 VDD.n550 6.772
R2386 VDD.n549 VDD.n546 6.772
R2387 VDD.n636 VDD.n621 6.772
R2388 VDD.n634 VDD.n631 6.772
R2389 VDD.n630 VDD.n627 6.772
R2390 VDD.n717 VDD.n702 6.772
R2391 VDD.n715 VDD.n712 6.772
R2392 VDD.n711 VDD.n708 6.772
R2393 VDD.n798 VDD.n783 6.772
R2394 VDD.n796 VDD.n793 6.772
R2395 VDD.n792 VDD.n789 6.772
R2396 VDD.n1674 VDD.n1659 6.772
R2397 VDD.n1672 VDD.n1669 6.772
R2398 VDD.n1668 VDD.n1665 6.772
R2399 VDD.n1593 VDD.n1578 6.772
R2400 VDD.n1591 VDD.n1588 6.772
R2401 VDD.n1587 VDD.n1584 6.772
R2402 VDD.n1512 VDD.n1497 6.772
R2403 VDD.n1510 VDD.n1507 6.772
R2404 VDD.n1506 VDD.n1503 6.772
R2405 VDD.n1431 VDD.n1416 6.772
R2406 VDD.n1429 VDD.n1426 6.772
R2407 VDD.n1425 VDD.n1422 6.772
R2408 VDD.n1350 VDD.n1335 6.772
R2409 VDD.n1348 VDD.n1345 6.772
R2410 VDD.n1344 VDD.n1341 6.772
R2411 VDD.n1269 VDD.n1254 6.772
R2412 VDD.n1267 VDD.n1264 6.772
R2413 VDD.n1263 VDD.n1260 6.772
R2414 VDD.n1188 VDD.n1173 6.772
R2415 VDD.n1186 VDD.n1183 6.772
R2416 VDD.n1182 VDD.n1179 6.772
R2417 VDD.n1107 VDD.n1092 6.772
R2418 VDD.n1105 VDD.n1102 6.772
R2419 VDD.n1101 VDD.n1098 6.772
R2420 VDD.n1026 VDD.n1011 6.772
R2421 VDD.n1024 VDD.n1021 6.772
R2422 VDD.n1020 VDD.n1017 6.772
R2423 VDD.n865 VDD.n851 6.772
R2424 VDD.n863 VDD.n860 6.772
R2425 VDD.n859 VDD.n856 6.772
R2426 VDD.n51 VDD.n50 6.772
R2427 VDD.n56 VDD.n55 6.772
R2428 VDD.n60 VDD.n59 6.772
R2429 VDD.n63 VDD.n62 6.772
R2430 VDD.n110 VDD.n109 6.772
R2431 VDD.n114 VDD.n113 6.772
R2432 VDD.n117 VDD.n116 6.772
R2433 VDD.n164 VDD.n163 6.772
R2434 VDD.n168 VDD.n167 6.772
R2435 VDD.n171 VDD.n170 6.772
R2436 VDD.n225 VDD.n224 6.772
R2437 VDD.n229 VDD.n228 6.772
R2438 VDD.n232 VDD.n231 6.772
R2439 VDD.n306 VDD.n305 6.772
R2440 VDD.n310 VDD.n309 6.772
R2441 VDD.n313 VDD.n312 6.772
R2442 VDD.n387 VDD.n386 6.772
R2443 VDD.n391 VDD.n390 6.772
R2444 VDD.n394 VDD.n393 6.772
R2445 VDD.n468 VDD.n467 6.772
R2446 VDD.n472 VDD.n471 6.772
R2447 VDD.n475 VDD.n474 6.772
R2448 VDD.n549 VDD.n548 6.772
R2449 VDD.n553 VDD.n552 6.772
R2450 VDD.n556 VDD.n555 6.772
R2451 VDD.n630 VDD.n629 6.772
R2452 VDD.n634 VDD.n633 6.772
R2453 VDD.n637 VDD.n636 6.772
R2454 VDD.n711 VDD.n710 6.772
R2455 VDD.n715 VDD.n714 6.772
R2456 VDD.n718 VDD.n717 6.772
R2457 VDD.n792 VDD.n791 6.772
R2458 VDD.n796 VDD.n795 6.772
R2459 VDD.n799 VDD.n798 6.772
R2460 VDD.n1668 VDD.n1667 6.772
R2461 VDD.n1672 VDD.n1671 6.772
R2462 VDD.n1675 VDD.n1674 6.772
R2463 VDD.n1587 VDD.n1586 6.772
R2464 VDD.n1591 VDD.n1590 6.772
R2465 VDD.n1594 VDD.n1593 6.772
R2466 VDD.n1506 VDD.n1505 6.772
R2467 VDD.n1510 VDD.n1509 6.772
R2468 VDD.n1513 VDD.n1512 6.772
R2469 VDD.n1425 VDD.n1424 6.772
R2470 VDD.n1429 VDD.n1428 6.772
R2471 VDD.n1432 VDD.n1431 6.772
R2472 VDD.n1344 VDD.n1343 6.772
R2473 VDD.n1348 VDD.n1347 6.772
R2474 VDD.n1351 VDD.n1350 6.772
R2475 VDD.n1263 VDD.n1262 6.772
R2476 VDD.n1267 VDD.n1266 6.772
R2477 VDD.n1270 VDD.n1269 6.772
R2478 VDD.n1182 VDD.n1181 6.772
R2479 VDD.n1186 VDD.n1185 6.772
R2480 VDD.n1189 VDD.n1188 6.772
R2481 VDD.n1101 VDD.n1100 6.772
R2482 VDD.n1105 VDD.n1104 6.772
R2483 VDD.n1108 VDD.n1107 6.772
R2484 VDD.n1020 VDD.n1019 6.772
R2485 VDD.n1024 VDD.n1023 6.772
R2486 VDD.n1027 VDD.n1026 6.772
R2487 VDD.n859 VDD.n858 6.772
R2488 VDD.n863 VDD.n862 6.772
R2489 VDD.n866 VDD.n865 6.772
R2490 VDD.n946 VDD.n945 6.772
R2491 VDD.n933 VDD.n930 6.772
R2492 VDD.n938 VDD.n935 6.772
R2493 VDD.n943 VDD.n940 6.772
R2494 VDD.n943 VDD.n942 6.772
R2495 VDD.n938 VDD.n937 6.772
R2496 VDD.n933 VDD.n932 6.772
R2497 VDD.n945 VDD.n929 6.772
R2498 VDD.n275 VDD.n271 6.69
R2499 VDD.n356 VDD.n352 6.69
R2500 VDD.n437 VDD.n433 6.69
R2501 VDD.n518 VDD.n514 6.69
R2502 VDD.n599 VDD.n595 6.69
R2503 VDD.n680 VDD.n676 6.69
R2504 VDD.n761 VDD.n757 6.69
R2505 VDD.n842 VDD.n838 6.69
R2506 VDD.n1621 VDD.n1617 6.69
R2507 VDD.n1540 VDD.n1536 6.69
R2508 VDD.n1459 VDD.n1455 6.69
R2509 VDD.n1378 VDD.n1374 6.69
R2510 VDD.n1297 VDD.n1293 6.69
R2511 VDD.n1216 VDD.n1212 6.69
R2512 VDD.n1135 VDD.n1131 6.69
R2513 VDD.n1054 VDD.n1050 6.69
R2514 VDD.n973 VDD.n969 6.69
R2515 VDD.n891 VDD.n887 6.69
R2516 VDD.n16 VDD.n15 6.458
R2517 VDD.n258 VDD.n257 6.296
R2518 VDD.n339 VDD.n338 6.296
R2519 VDD.n420 VDD.n419 6.296
R2520 VDD.n501 VDD.n500 6.296
R2521 VDD.n582 VDD.n581 6.296
R2522 VDD.n663 VDD.n662 6.296
R2523 VDD.n744 VDD.n743 6.296
R2524 VDD.n825 VDD.n824 6.296
R2525 VDD.n1638 VDD.n1637 6.296
R2526 VDD.n1557 VDD.n1556 6.296
R2527 VDD.n1476 VDD.n1475 6.296
R2528 VDD.n1395 VDD.n1394 6.296
R2529 VDD.n1314 VDD.n1313 6.296
R2530 VDD.n1233 VDD.n1232 6.296
R2531 VDD.n1152 VDD.n1151 6.296
R2532 VDD.n1071 VDD.n1070 6.296
R2533 VDD.n990 VDD.n989 6.296
R2534 VDD.n908 VDD.n907 6.296
R2535 VDD.n105 VDD.n104 6.202
R2536 VDD.n159 VDD.n158 6.202
R2537 VDD.n220 VDD.n219 6.202
R2538 VDD.n301 VDD.n300 6.202
R2539 VDD.n382 VDD.n381 6.202
R2540 VDD.n463 VDD.n462 6.202
R2541 VDD.n544 VDD.n543 6.202
R2542 VDD.n625 VDD.n624 6.202
R2543 VDD.n706 VDD.n705 6.202
R2544 VDD.n787 VDD.n786 6.202
R2545 VDD.n1663 VDD.n1662 6.202
R2546 VDD.n1582 VDD.n1581 6.202
R2547 VDD.n1501 VDD.n1500 6.202
R2548 VDD.n1420 VDD.n1419 6.202
R2549 VDD.n1339 VDD.n1338 6.202
R2550 VDD.n1258 VDD.n1257 6.202
R2551 VDD.n1177 VDD.n1176 6.202
R2552 VDD.n1096 VDD.n1095 6.202
R2553 VDD.n1015 VDD.n1014 6.202
R2554 VDD.n854 VDD.n853 6.202
R2555 VDD.n196 VDD.n195 4.576
R2556 VDD.n208 VDD.n205 2.754
R2557 VDD.n182 VDD.n179 2.361
R2558 VDD.n28 VDD.n24 1.967
R2559 VDD.n38 VDD.n37 1.967
R2560 VDD.n14 VDD.n7 1.329
R2561 VDD.n14 VDD.n8 1.329
R2562 VDD.n14 VDD.n12 1.329
R2563 VDD.n14 VDD.n13 1.329
R2564 VDD.n15 VDD.n14 0.696
R2565 VDD.n14 VDD.n4 0.696
R2566 VDD.n285 VDD.n282 0.393
R2567 VDD.n366 VDD.n363 0.393
R2568 VDD.n447 VDD.n444 0.393
R2569 VDD.n528 VDD.n525 0.393
R2570 VDD.n609 VDD.n606 0.393
R2571 VDD.n690 VDD.n687 0.393
R2572 VDD.n771 VDD.n768 0.393
R2573 VDD.n1690 VDD.n1687 0.393
R2574 VDD.n1609 VDD.n1606 0.393
R2575 VDD.n1528 VDD.n1525 0.393
R2576 VDD.n1447 VDD.n1444 0.393
R2577 VDD.n1366 VDD.n1363 0.393
R2578 VDD.n1285 VDD.n1282 0.393
R2579 VDD.n1204 VDD.n1201 0.393
R2580 VDD.n1123 VDD.n1120 0.393
R2581 VDD.n1042 VDD.n1039 0.393
R2582 VDD.n961 VDD.n958 0.393
R2583 VDD.n879 VDD.n876 0.393
R2584 VDD.n61 VDD.n60 0.365
R2585 VDD.n61 VDD.n56 0.365
R2586 VDD.n61 VDD.n51 0.365
R2587 VDD.n62 VDD.n61 0.365
R2588 VDD.n115 VDD.n114 0.365
R2589 VDD.n115 VDD.n110 0.365
R2590 VDD.n116 VDD.n115 0.365
R2591 VDD.n169 VDD.n168 0.365
R2592 VDD.n169 VDD.n164 0.365
R2593 VDD.n170 VDD.n169 0.365
R2594 VDD.n230 VDD.n229 0.365
R2595 VDD.n230 VDD.n225 0.365
R2596 VDD.n231 VDD.n230 0.365
R2597 VDD.n311 VDD.n310 0.365
R2598 VDD.n311 VDD.n306 0.365
R2599 VDD.n312 VDD.n311 0.365
R2600 VDD.n392 VDD.n391 0.365
R2601 VDD.n392 VDD.n387 0.365
R2602 VDD.n393 VDD.n392 0.365
R2603 VDD.n473 VDD.n472 0.365
R2604 VDD.n473 VDD.n468 0.365
R2605 VDD.n474 VDD.n473 0.365
R2606 VDD.n554 VDD.n553 0.365
R2607 VDD.n554 VDD.n549 0.365
R2608 VDD.n555 VDD.n554 0.365
R2609 VDD.n635 VDD.n634 0.365
R2610 VDD.n635 VDD.n630 0.365
R2611 VDD.n636 VDD.n635 0.365
R2612 VDD.n716 VDD.n715 0.365
R2613 VDD.n716 VDD.n711 0.365
R2614 VDD.n717 VDD.n716 0.365
R2615 VDD.n797 VDD.n796 0.365
R2616 VDD.n797 VDD.n792 0.365
R2617 VDD.n798 VDD.n797 0.365
R2618 VDD.n1673 VDD.n1672 0.365
R2619 VDD.n1673 VDD.n1668 0.365
R2620 VDD.n1674 VDD.n1673 0.365
R2621 VDD.n1592 VDD.n1591 0.365
R2622 VDD.n1592 VDD.n1587 0.365
R2623 VDD.n1593 VDD.n1592 0.365
R2624 VDD.n1511 VDD.n1510 0.365
R2625 VDD.n1511 VDD.n1506 0.365
R2626 VDD.n1512 VDD.n1511 0.365
R2627 VDD.n1430 VDD.n1429 0.365
R2628 VDD.n1430 VDD.n1425 0.365
R2629 VDD.n1431 VDD.n1430 0.365
R2630 VDD.n1349 VDD.n1348 0.365
R2631 VDD.n1349 VDD.n1344 0.365
R2632 VDD.n1350 VDD.n1349 0.365
R2633 VDD.n1268 VDD.n1267 0.365
R2634 VDD.n1268 VDD.n1263 0.365
R2635 VDD.n1269 VDD.n1268 0.365
R2636 VDD.n1187 VDD.n1186 0.365
R2637 VDD.n1187 VDD.n1182 0.365
R2638 VDD.n1188 VDD.n1187 0.365
R2639 VDD.n1106 VDD.n1105 0.365
R2640 VDD.n1106 VDD.n1101 0.365
R2641 VDD.n1107 VDD.n1106 0.365
R2642 VDD.n1025 VDD.n1024 0.365
R2643 VDD.n1025 VDD.n1020 0.365
R2644 VDD.n1026 VDD.n1025 0.365
R2645 VDD.n864 VDD.n863 0.365
R2646 VDD.n864 VDD.n859 0.365
R2647 VDD.n865 VDD.n864 0.365
R2648 VDD.n944 VDD.n943 0.365
R2649 VDD.n944 VDD.n938 0.365
R2650 VDD.n944 VDD.n933 0.365
R2651 VDD.n945 VDD.n944 0.365
R2652 VDD.n70 VDD.n43 0.29
R2653 VDD.n124 VDD.n98 0.29
R2654 VDD.n178 VDD.n152 0.29
R2655 VDD.n239 VDD.n213 0.29
R2656 VDD.n320 VDD.n294 0.29
R2657 VDD.n401 VDD.n375 0.29
R2658 VDD.n482 VDD.n456 0.29
R2659 VDD.n563 VDD.n537 0.29
R2660 VDD.n644 VDD.n618 0.29
R2661 VDD.n725 VDD.n699 0.29
R2662 VDD.n806 VDD.n780 0.29
R2663 VDD.n1682 VDD.n1656 0.29
R2664 VDD.n1601 VDD.n1575 0.29
R2665 VDD.n1520 VDD.n1494 0.29
R2666 VDD.n1439 VDD.n1413 0.29
R2667 VDD.n1358 VDD.n1332 0.29
R2668 VDD.n1277 VDD.n1251 0.29
R2669 VDD.n1196 VDD.n1170 0.29
R2670 VDD.n1115 VDD.n1089 0.29
R2671 VDD.n1034 VDD.n1008 0.29
R2672 VDD.n953 VDD.n926 0.29
R2673 VDD.n871 VDD 0.207
R2674 VDD.n269 VDD.n264 0.197
R2675 VDD.n350 VDD.n345 0.197
R2676 VDD.n431 VDD.n426 0.197
R2677 VDD.n512 VDD.n507 0.197
R2678 VDD.n593 VDD.n588 0.197
R2679 VDD.n674 VDD.n669 0.197
R2680 VDD.n755 VDD.n750 0.197
R2681 VDD.n836 VDD.n831 0.197
R2682 VDD.n1632 VDD.n1627 0.197
R2683 VDD.n1551 VDD.n1546 0.197
R2684 VDD.n1470 VDD.n1465 0.197
R2685 VDD.n1389 VDD.n1384 0.197
R2686 VDD.n1308 VDD.n1303 0.197
R2687 VDD.n1227 VDD.n1222 0.197
R2688 VDD.n1146 VDD.n1141 0.197
R2689 VDD.n1065 VDD.n1060 0.197
R2690 VDD.n984 VDD.n979 0.197
R2691 VDD.n902 VDD.n897 0.197
R2692 VDD.n86 VDD.n82 0.181
R2693 VDD.n140 VDD.n136 0.181
R2694 VDD.n199 VDD.n194 0.181
R2695 VDD.n33 VDD.n29 0.157
R2696 VDD.n39 VDD.n33 0.157
R2697 VDD.n43 VDD.n39 0.145
R2698 VDD.n74 VDD.n70 0.145
R2699 VDD.n78 VDD.n74 0.145
R2700 VDD.n82 VDD.n78 0.145
R2701 VDD.n90 VDD.n86 0.145
R2702 VDD.n94 VDD.n90 0.145
R2703 VDD.n98 VDD.n94 0.145
R2704 VDD.n128 VDD.n124 0.145
R2705 VDD.n132 VDD.n128 0.145
R2706 VDD.n136 VDD.n132 0.145
R2707 VDD.n144 VDD.n140 0.145
R2708 VDD.n148 VDD.n144 0.145
R2709 VDD.n152 VDD.n148 0.145
R2710 VDD.n183 VDD.n178 0.145
R2711 VDD.n188 VDD.n183 0.145
R2712 VDD.n194 VDD.n188 0.145
R2713 VDD.n204 VDD.n199 0.145
R2714 VDD.n209 VDD.n204 0.145
R2715 VDD.n213 VDD.n209 0.145
R2716 VDD.n243 VDD.n239 0.145
R2717 VDD.n247 VDD.n243 0.145
R2718 VDD.n252 VDD.n247 0.145
R2719 VDD.n259 VDD.n252 0.145
R2720 VDD.n264 VDD.n259 0.145
R2721 VDD.n276 VDD.n269 0.145
R2722 VDD.n281 VDD.n276 0.145
R2723 VDD.n286 VDD.n281 0.145
R2724 VDD.n290 VDD.n286 0.145
R2725 VDD.n294 VDD.n290 0.145
R2726 VDD.n324 VDD.n320 0.145
R2727 VDD.n328 VDD.n324 0.145
R2728 VDD.n333 VDD.n328 0.145
R2729 VDD.n340 VDD.n333 0.145
R2730 VDD.n345 VDD.n340 0.145
R2731 VDD.n357 VDD.n350 0.145
R2732 VDD.n362 VDD.n357 0.145
R2733 VDD.n367 VDD.n362 0.145
R2734 VDD.n371 VDD.n367 0.145
R2735 VDD.n375 VDD.n371 0.145
R2736 VDD.n405 VDD.n401 0.145
R2737 VDD.n409 VDD.n405 0.145
R2738 VDD.n414 VDD.n409 0.145
R2739 VDD.n421 VDD.n414 0.145
R2740 VDD.n426 VDD.n421 0.145
R2741 VDD.n438 VDD.n431 0.145
R2742 VDD.n443 VDD.n438 0.145
R2743 VDD.n448 VDD.n443 0.145
R2744 VDD.n452 VDD.n448 0.145
R2745 VDD.n456 VDD.n452 0.145
R2746 VDD.n486 VDD.n482 0.145
R2747 VDD.n490 VDD.n486 0.145
R2748 VDD.n495 VDD.n490 0.145
R2749 VDD.n502 VDD.n495 0.145
R2750 VDD.n507 VDD.n502 0.145
R2751 VDD.n519 VDD.n512 0.145
R2752 VDD.n524 VDD.n519 0.145
R2753 VDD.n529 VDD.n524 0.145
R2754 VDD.n533 VDD.n529 0.145
R2755 VDD.n537 VDD.n533 0.145
R2756 VDD.n567 VDD.n563 0.145
R2757 VDD.n571 VDD.n567 0.145
R2758 VDD.n576 VDD.n571 0.145
R2759 VDD.n583 VDD.n576 0.145
R2760 VDD.n588 VDD.n583 0.145
R2761 VDD.n600 VDD.n593 0.145
R2762 VDD.n605 VDD.n600 0.145
R2763 VDD.n610 VDD.n605 0.145
R2764 VDD.n614 VDD.n610 0.145
R2765 VDD.n618 VDD.n614 0.145
R2766 VDD.n648 VDD.n644 0.145
R2767 VDD.n652 VDD.n648 0.145
R2768 VDD.n657 VDD.n652 0.145
R2769 VDD.n664 VDD.n657 0.145
R2770 VDD.n669 VDD.n664 0.145
R2771 VDD.n681 VDD.n674 0.145
R2772 VDD.n686 VDD.n681 0.145
R2773 VDD.n691 VDD.n686 0.145
R2774 VDD.n695 VDD.n691 0.145
R2775 VDD.n699 VDD.n695 0.145
R2776 VDD.n729 VDD.n725 0.145
R2777 VDD.n733 VDD.n729 0.145
R2778 VDD.n738 VDD.n733 0.145
R2779 VDD.n745 VDD.n738 0.145
R2780 VDD.n750 VDD.n745 0.145
R2781 VDD.n762 VDD.n755 0.145
R2782 VDD.n767 VDD.n762 0.145
R2783 VDD.n772 VDD.n767 0.145
R2784 VDD.n776 VDD.n772 0.145
R2785 VDD.n780 VDD.n776 0.145
R2786 VDD.n810 VDD.n806 0.145
R2787 VDD.n814 VDD.n810 0.145
R2788 VDD.n819 VDD.n814 0.145
R2789 VDD.n826 VDD.n819 0.145
R2790 VDD.n831 VDD.n826 0.145
R2791 VDD.n843 VDD.n836 0.145
R2792 VDD.n848 VDD.n843 0.145
R2793 VDD.n1691 VDD.n1686 0.145
R2794 VDD.n1686 VDD.n1682 0.145
R2795 VDD.n1656 VDD.n1652 0.145
R2796 VDD.n1652 VDD.n1648 0.145
R2797 VDD.n1648 VDD.n1644 0.145
R2798 VDD.n1644 VDD.n1639 0.145
R2799 VDD.n1639 VDD.n1632 0.145
R2800 VDD.n1627 VDD.n1622 0.145
R2801 VDD.n1622 VDD.n1615 0.145
R2802 VDD.n1615 VDD.n1610 0.145
R2803 VDD.n1610 VDD.n1605 0.145
R2804 VDD.n1605 VDD.n1601 0.145
R2805 VDD.n1575 VDD.n1571 0.145
R2806 VDD.n1571 VDD.n1567 0.145
R2807 VDD.n1567 VDD.n1563 0.145
R2808 VDD.n1563 VDD.n1558 0.145
R2809 VDD.n1558 VDD.n1551 0.145
R2810 VDD.n1546 VDD.n1541 0.145
R2811 VDD.n1541 VDD.n1534 0.145
R2812 VDD.n1534 VDD.n1529 0.145
R2813 VDD.n1529 VDD.n1524 0.145
R2814 VDD.n1524 VDD.n1520 0.145
R2815 VDD.n1494 VDD.n1490 0.145
R2816 VDD.n1490 VDD.n1486 0.145
R2817 VDD.n1486 VDD.n1482 0.145
R2818 VDD.n1482 VDD.n1477 0.145
R2819 VDD.n1477 VDD.n1470 0.145
R2820 VDD.n1465 VDD.n1460 0.145
R2821 VDD.n1460 VDD.n1453 0.145
R2822 VDD.n1453 VDD.n1448 0.145
R2823 VDD.n1448 VDD.n1443 0.145
R2824 VDD.n1443 VDD.n1439 0.145
R2825 VDD.n1413 VDD.n1409 0.145
R2826 VDD.n1409 VDD.n1405 0.145
R2827 VDD.n1405 VDD.n1401 0.145
R2828 VDD.n1401 VDD.n1396 0.145
R2829 VDD.n1396 VDD.n1389 0.145
R2830 VDD.n1384 VDD.n1379 0.145
R2831 VDD.n1379 VDD.n1372 0.145
R2832 VDD.n1372 VDD.n1367 0.145
R2833 VDD.n1367 VDD.n1362 0.145
R2834 VDD.n1362 VDD.n1358 0.145
R2835 VDD.n1332 VDD.n1328 0.145
R2836 VDD.n1328 VDD.n1324 0.145
R2837 VDD.n1324 VDD.n1320 0.145
R2838 VDD.n1320 VDD.n1315 0.145
R2839 VDD.n1315 VDD.n1308 0.145
R2840 VDD.n1303 VDD.n1298 0.145
R2841 VDD.n1298 VDD.n1291 0.145
R2842 VDD.n1291 VDD.n1286 0.145
R2843 VDD.n1286 VDD.n1281 0.145
R2844 VDD.n1281 VDD.n1277 0.145
R2845 VDD.n1251 VDD.n1247 0.145
R2846 VDD.n1247 VDD.n1243 0.145
R2847 VDD.n1243 VDD.n1239 0.145
R2848 VDD.n1239 VDD.n1234 0.145
R2849 VDD.n1234 VDD.n1227 0.145
R2850 VDD.n1222 VDD.n1217 0.145
R2851 VDD.n1217 VDD.n1210 0.145
R2852 VDD.n1210 VDD.n1205 0.145
R2853 VDD.n1205 VDD.n1200 0.145
R2854 VDD.n1200 VDD.n1196 0.145
R2855 VDD.n1170 VDD.n1166 0.145
R2856 VDD.n1166 VDD.n1162 0.145
R2857 VDD.n1162 VDD.n1158 0.145
R2858 VDD.n1158 VDD.n1153 0.145
R2859 VDD.n1153 VDD.n1146 0.145
R2860 VDD.n1141 VDD.n1136 0.145
R2861 VDD.n1136 VDD.n1129 0.145
R2862 VDD.n1129 VDD.n1124 0.145
R2863 VDD.n1124 VDD.n1119 0.145
R2864 VDD.n1119 VDD.n1115 0.145
R2865 VDD.n1089 VDD.n1085 0.145
R2866 VDD.n1085 VDD.n1081 0.145
R2867 VDD.n1081 VDD.n1077 0.145
R2868 VDD.n1077 VDD.n1072 0.145
R2869 VDD.n1072 VDD.n1065 0.145
R2870 VDD.n1060 VDD.n1055 0.145
R2871 VDD.n1055 VDD.n1048 0.145
R2872 VDD.n1048 VDD.n1043 0.145
R2873 VDD.n1043 VDD.n1038 0.145
R2874 VDD.n1038 VDD.n1034 0.145
R2875 VDD.n1008 VDD.n1004 0.145
R2876 VDD.n1004 VDD.n1000 0.145
R2877 VDD.n1000 VDD.n996 0.145
R2878 VDD.n996 VDD.n991 0.145
R2879 VDD.n991 VDD.n984 0.145
R2880 VDD.n979 VDD.n974 0.145
R2881 VDD.n974 VDD.n967 0.145
R2882 VDD.n967 VDD.n962 0.145
R2883 VDD.n962 VDD.n957 0.145
R2884 VDD.n957 VDD.n953 0.145
R2885 VDD.n926 VDD.n922 0.145
R2886 VDD.n922 VDD.n918 0.145
R2887 VDD.n918 VDD.n914 0.145
R2888 VDD.n914 VDD.n909 0.145
R2889 VDD.n909 VDD.n902 0.145
R2890 VDD.n897 VDD.n892 0.145
R2891 VDD.n892 VDD.n885 0.145
R2892 VDD.n885 VDD.n880 0.145
R2893 VDD.n880 VDD.n875 0.145
R2894 VDD.n875 VDD.n871 0.145
R2895 VDD VDD.n1691 0.086
R2896 VDD VDD.n848 0.058
R2897 a_15991_989.n2 a_15991_989.t9 512.525
R2898 a_15991_989.n0 a_15991_989.t14 477.179
R2899 a_15991_989.n5 a_15991_989.t7 454.685
R2900 a_15991_989.n5 a_15991_989.t13 428.979
R2901 a_15991_989.n0 a_15991_989.t12 406.485
R2902 a_15991_989.n2 a_15991_989.t10 371.139
R2903 a_15991_989.n1 a_15991_989.t8 363.924
R2904 a_15991_989.n4 a_15991_989.t11 303.606
R2905 a_15991_989.n6 a_15991_989.t15 184.853
R2906 a_15991_989.n11 a_15991_989.n10 159.998
R2907 a_15991_989.n11 a_15991_989.n6 156.035
R2908 a_15991_989.n12 a_15991_989.n4 153.043
R2909 a_15991_989.n6 a_15991_989.n5 151.553
R2910 a_15991_989.n16 a_15991_989.n12 144.246
R2911 a_15991_989.n3 a_15991_989.n1 101.359
R2912 a_15991_989.n12 a_15991_989.n11 79.658
R2913 a_15991_989.n15 a_15991_989.n14 79.232
R2914 a_15991_989.n3 a_15991_989.n2 71.88
R2915 a_15991_989.n16 a_15991_989.n15 63.152
R2916 a_15991_989.n4 a_15991_989.n3 53.891
R2917 a_15991_989.n10 a_15991_989.n9 30
R2918 a_15991_989.n8 a_15991_989.n7 24.383
R2919 a_15991_989.n10 a_15991_989.n8 23.684
R2920 a_15991_989.n15 a_15991_989.n13 16.08
R2921 a_15991_989.n17 a_15991_989.n16 16.078
R2922 a_15991_989.n1 a_15991_989.n0 15.776
R2923 a_15991_989.n13 a_15991_989.t5 14.282
R2924 a_15991_989.n13 a_15991_989.t6 14.282
R2925 a_15991_989.n14 a_15991_989.t4 14.282
R2926 a_15991_989.n14 a_15991_989.t0 14.282
R2927 a_15991_989.t2 a_15991_989.n17 14.282
R2928 a_15991_989.n17 a_15991_989.t1 14.282
R2929 a_15669_1050.n0 a_15669_1050.t9 512.525
R2930 a_15669_1050.n0 a_15669_1050.t7 371.139
R2931 a_15669_1050.n1 a_15669_1050.t8 287.668
R2932 a_15669_1050.n6 a_15669_1050.n5 213.104
R2933 a_15669_1050.n10 a_15669_1050.n6 170.799
R2934 a_15669_1050.n1 a_15669_1050.n0 162.713
R2935 a_15669_1050.n6 a_15669_1050.n1 153.315
R2936 a_15669_1050.n9 a_15669_1050.n8 79.232
R2937 a_15669_1050.n10 a_15669_1050.n9 63.152
R2938 a_15669_1050.n5 a_15669_1050.n4 30
R2939 a_15669_1050.n3 a_15669_1050.n2 24.383
R2940 a_15669_1050.n5 a_15669_1050.n3 23.684
R2941 a_15669_1050.n9 a_15669_1050.n7 16.08
R2942 a_15669_1050.n11 a_15669_1050.n10 16.078
R2943 a_15669_1050.n7 a_15669_1050.t5 14.282
R2944 a_15669_1050.n7 a_15669_1050.t0 14.282
R2945 a_15669_1050.n8 a_15669_1050.t1 14.282
R2946 a_15669_1050.n8 a_15669_1050.t6 14.282
R2947 a_15669_1050.n11 a_15669_1050.t3 14.282
R2948 a_15669_1050.t4 a_15669_1050.n11 14.282
R2949 a_11821_1050.n7 a_11821_1050.t7 512.525
R2950 a_11821_1050.n5 a_11821_1050.t12 512.525
R2951 a_11821_1050.n7 a_11821_1050.t11 371.139
R2952 a_11821_1050.n5 a_11821_1050.t8 371.139
R2953 a_11821_1050.n8 a_11821_1050.t9 234.921
R2954 a_11821_1050.n6 a_11821_1050.t10 234.921
R2955 a_11821_1050.n10 a_11821_1050.n4 223.546
R2956 a_11821_1050.n8 a_11821_1050.n7 215.46
R2957 a_11821_1050.n6 a_11821_1050.n5 215.46
R2958 a_11821_1050.n12 a_11821_1050.n10 166.879
R2959 a_11821_1050.n9 a_11821_1050.n6 79.491
R2960 a_11821_1050.n3 a_11821_1050.n2 79.232
R2961 a_11821_1050.n10 a_11821_1050.n9 77.315
R2962 a_11821_1050.n9 a_11821_1050.n8 76
R2963 a_11821_1050.n4 a_11821_1050.n3 63.152
R2964 a_11821_1050.n4 a_11821_1050.n0 16.08
R2965 a_11821_1050.n3 a_11821_1050.n1 16.08
R2966 a_11821_1050.n12 a_11821_1050.n11 15.218
R2967 a_11821_1050.n0 a_11821_1050.t6 14.282
R2968 a_11821_1050.n0 a_11821_1050.t1 14.282
R2969 a_11821_1050.n1 a_11821_1050.t0 14.282
R2970 a_11821_1050.n1 a_11821_1050.t3 14.282
R2971 a_11821_1050.n2 a_11821_1050.t4 14.282
R2972 a_11821_1050.n2 a_11821_1050.t2 14.282
R2973 a_11821_1050.n13 a_11821_1050.n12 12.014
R2974 a_12143_989.n1 a_12143_989.t7 512.525
R2975 a_12143_989.n3 a_12143_989.t8 454.685
R2976 a_12143_989.n3 a_12143_989.t12 428.979
R2977 a_12143_989.n1 a_12143_989.t10 371.139
R2978 a_12143_989.n2 a_12143_989.t9 287.668
R2979 a_12143_989.n4 a_12143_989.t11 237.959
R2980 a_12143_989.n10 a_12143_989.n9 213.104
R2981 a_12143_989.n11 a_12143_989.n10 170.799
R2982 a_12143_989.n2 a_12143_989.n1 162.713
R2983 a_12143_989.n4 a_12143_989.n3 98.447
R2984 a_12143_989.n5 a_12143_989.n2 84.388
R2985 a_12143_989.n5 a_12143_989.n4 80.035
R2986 a_12143_989.n13 a_12143_989.n12 79.232
R2987 a_12143_989.n10 a_12143_989.n5 76
R2988 a_12143_989.n13 a_12143_989.n11 63.152
R2989 a_12143_989.n9 a_12143_989.n8 30
R2990 a_12143_989.n7 a_12143_989.n6 24.383
R2991 a_12143_989.n9 a_12143_989.n7 23.684
R2992 a_12143_989.n11 a_12143_989.n0 16.08
R2993 a_12143_989.n14 a_12143_989.n13 16.078
R2994 a_12143_989.n0 a_12143_989.t6 14.282
R2995 a_12143_989.n0 a_12143_989.t5 14.282
R2996 a_12143_989.n12 a_12143_989.t3 14.282
R2997 a_12143_989.n12 a_12143_989.t2 14.282
R2998 a_12143_989.t1 a_12143_989.n14 14.282
R2999 a_12143_989.n14 a_12143_989.t0 14.282
R3000 a_4125_1050.n5 a_4125_1050.t8 512.525
R3001 a_4125_1050.n5 a_4125_1050.t9 371.139
R3002 a_4125_1050.n6 a_4125_1050.t7 287.668
R3003 a_4125_1050.n9 a_4125_1050.n7 219.626
R3004 a_4125_1050.n7 a_4125_1050.n4 170.799
R3005 a_4125_1050.n6 a_4125_1050.n5 162.713
R3006 a_4125_1050.n7 a_4125_1050.n6 153.315
R3007 a_4125_1050.n3 a_4125_1050.n2 79.232
R3008 a_4125_1050.n4 a_4125_1050.n3 63.152
R3009 a_4125_1050.n4 a_4125_1050.n0 16.08
R3010 a_4125_1050.n3 a_4125_1050.n1 16.08
R3011 a_4125_1050.n9 a_4125_1050.n8 15.218
R3012 a_4125_1050.n0 a_4125_1050.t6 14.282
R3013 a_4125_1050.n0 a_4125_1050.t2 14.282
R3014 a_4125_1050.n1 a_4125_1050.t1 14.282
R3015 a_4125_1050.n1 a_4125_1050.t5 14.282
R3016 a_4125_1050.n2 a_4125_1050.t4 14.282
R3017 a_4125_1050.n2 a_4125_1050.t3 14.282
R3018 a_4125_1050.n10 a_4125_1050.n9 12.014
R3019 a_4901_103.n5 a_4901_103.n4 19.724
R3020 a_4901_103.t0 a_4901_103.n3 11.595
R3021 a_4901_103.t0 a_4901_103.n5 9.207
R3022 a_4901_103.n2 a_4901_103.n1 2.455
R3023 a_4901_103.n2 a_4901_103.n0 1.32
R3024 a_4901_103.t0 a_4901_103.n2 0.246
R3025 SN.n14 SN.t6 479.223
R3026 SN.n11 SN.t12 479.223
R3027 SN.n8 SN.t13 479.223
R3028 SN.n5 SN.t1 479.223
R3029 SN.n2 SN.t14 479.223
R3030 SN.n0 SN.t0 479.223
R3031 SN.n14 SN.t15 375.52
R3032 SN.n11 SN.t2 375.52
R3033 SN.n8 SN.t4 375.52
R3034 SN.n5 SN.t5 375.52
R3035 SN.n2 SN.t7 375.52
R3036 SN.n0 SN.t10 375.52
R3037 SN.n12 SN.n11 201.982
R3038 SN.n6 SN.n5 201.982
R3039 SN.n1 SN.n0 201.982
R3040 SN.n3 SN.n2 199.731
R3041 SN.n9 SN.n8 199.731
R3042 SN.n15 SN.n14 199.731
R3043 SN.n12 SN.t17 141.649
R3044 SN.n6 SN.t8 141.649
R3045 SN.n1 SN.t9 141.649
R3046 SN.n15 SN.t16 128.128
R3047 SN.n9 SN.t3 128.128
R3048 SN.n3 SN.t11 128.128
R3049 SN.n4 SN.n1 86.561
R3050 SN.n7 SN.n6 76
R3051 SN.n13 SN.n12 76
R3052 SN.n4 SN.n3 49.346
R3053 SN.n10 SN.n9 49.346
R3054 SN.n16 SN.n15 49.346
R3055 SN.n7 SN.n4 10.564
R3056 SN.n13 SN.n10 10.564
R3057 SN.n10 SN.n7 10.561
R3058 SN.n16 SN.n13 10.561
R3059 SN.n16 SN 0.046
R3060 a_6371_989.n1 a_6371_989.t12 512.525
R3061 a_6371_989.n3 a_6371_989.t7 454.685
R3062 a_6371_989.n3 a_6371_989.t10 428.979
R3063 a_6371_989.n1 a_6371_989.t9 371.139
R3064 a_6371_989.n2 a_6371_989.t8 287.668
R3065 a_6371_989.n4 a_6371_989.t11 237.959
R3066 a_6371_989.n7 a_6371_989.n6 234.843
R3067 a_6371_989.n8 a_6371_989.n7 170.799
R3068 a_6371_989.n2 a_6371_989.n1 162.713
R3069 a_6371_989.n4 a_6371_989.n3 98.447
R3070 a_6371_989.n5 a_6371_989.n2 84.388
R3071 a_6371_989.n5 a_6371_989.n4 80.035
R3072 a_6371_989.n10 a_6371_989.n9 79.232
R3073 a_6371_989.n7 a_6371_989.n5 76
R3074 a_6371_989.n10 a_6371_989.n8 63.152
R3075 a_6371_989.n8 a_6371_989.n0 16.08
R3076 a_6371_989.n11 a_6371_989.n10 16.078
R3077 a_6371_989.n0 a_6371_989.t5 14.282
R3078 a_6371_989.n0 a_6371_989.t2 14.282
R3079 a_6371_989.n9 a_6371_989.t3 14.282
R3080 a_6371_989.n9 a_6371_989.t4 14.282
R3081 a_6371_989.t1 a_6371_989.n11 14.282
R3082 a_6371_989.n11 a_6371_989.t0 14.282
R3083 a_4447_989.n3 a_4447_989.t14 512.525
R3084 a_4447_989.n2 a_4447_989.t13 512.525
R3085 a_4447_989.n7 a_4447_989.t10 454.685
R3086 a_4447_989.n7 a_4447_989.t15 428.979
R3087 a_4447_989.n3 a_4447_989.t8 371.139
R3088 a_4447_989.n2 a_4447_989.t9 371.139
R3089 a_4447_989.n4 a_4447_989.n3 265.439
R3090 a_4447_989.n13 a_4447_989.n12 202.074
R3091 a_4447_989.n8 a_4447_989.t12 200.159
R3092 a_4447_989.n14 a_4447_989.n13 197.352
R3093 a_4447_989.n6 a_4447_989.n2 185.78
R3094 a_4447_989.n4 a_4447_989.t7 176.995
R3095 a_4447_989.n5 a_4447_989.t11 170.569
R3096 a_4447_989.n5 a_4447_989.n4 153.043
R3097 a_4447_989.n8 a_4447_989.n7 125
R3098 a_4447_989.n9 a_4447_989.n6 123.293
R3099 a_4447_989.n9 a_4447_989.n8 80.035
R3100 a_4447_989.n6 a_4447_989.n5 79.658
R3101 a_4447_989.n16 a_4447_989.n15 79.231
R3102 a_4447_989.n13 a_4447_989.n9 76
R3103 a_4447_989.n15 a_4447_989.n14 63.152
R3104 a_4447_989.n12 a_4447_989.n11 22.578
R3105 a_4447_989.n14 a_4447_989.n1 16.08
R3106 a_4447_989.n15 a_4447_989.n0 16.08
R3107 a_4447_989.n1 a_4447_989.t6 14.282
R3108 a_4447_989.n1 a_4447_989.t4 14.282
R3109 a_4447_989.n0 a_4447_989.t2 14.282
R3110 a_4447_989.n0 a_4447_989.t3 14.282
R3111 a_4447_989.t1 a_4447_989.n16 14.282
R3112 a_4447_989.n16 a_4447_989.t0 14.282
R3113 a_4447_989.n12 a_4447_989.n10 8.58
R3114 a_18760_101.t0 a_18760_101.n1 34.62
R3115 a_18760_101.t0 a_18760_101.n0 8.137
R3116 a_18760_101.t0 a_18760_101.n2 4.69
R3117 a_18094_101.t0 a_18094_101.n0 34.606
R3118 a_18094_101.t0 a_18094_101.n1 2.115
R3119 a_2201_1050.n1 a_2201_1050.t7 512.525
R3120 a_2201_1050.n1 a_2201_1050.t8 371.139
R3121 a_2201_1050.n2 a_2201_1050.t9 234.562
R3122 a_2201_1050.n5 a_2201_1050.n4 223.905
R3123 a_2201_1050.n2 a_2201_1050.n1 215.819
R3124 a_2201_1050.n4 a_2201_1050.n3 181.737
R3125 a_2201_1050.n4 a_2201_1050.n2 153.315
R3126 a_2201_1050.n7 a_2201_1050.n6 79.232
R3127 a_2201_1050.n7 a_2201_1050.n5 63.152
R3128 a_2201_1050.n5 a_2201_1050.n0 16.08
R3129 a_2201_1050.n8 a_2201_1050.n7 16.078
R3130 a_2201_1050.n0 a_2201_1050.t4 14.282
R3131 a_2201_1050.n0 a_2201_1050.t5 14.282
R3132 a_2201_1050.n6 a_2201_1050.t6 14.282
R3133 a_2201_1050.n6 a_2201_1050.t1 14.282
R3134 a_2201_1050.t3 a_2201_1050.n8 14.282
R3135 a_2201_1050.n8 a_2201_1050.t2 14.282
R3136 a_1561_989.n3 a_1561_989.t14 454.685
R3137 a_1561_989.n5 a_1561_989.t7 454.685
R3138 a_1561_989.n1 a_1561_989.t15 454.685
R3139 a_1561_989.n3 a_1561_989.t8 428.979
R3140 a_1561_989.n5 a_1561_989.t11 428.979
R3141 a_1561_989.n1 a_1561_989.t13 428.979
R3142 a_1561_989.n4 a_1561_989.t9 264.512
R3143 a_1561_989.n2 a_1561_989.t12 264.512
R3144 a_1561_989.n6 a_1561_989.t10 264.173
R3145 a_1561_989.n10 a_1561_989.n9 261.396
R3146 a_1561_989.n11 a_1561_989.n10 144.246
R3147 a_1561_989.n8 a_1561_989.n2 82.484
R3148 a_1561_989.n7 a_1561_989.n6 79.495
R3149 a_1561_989.n13 a_1561_989.n12 79.232
R3150 a_1561_989.n7 a_1561_989.n4 76
R3151 a_1561_989.n10 a_1561_989.n8 76
R3152 a_1561_989.n4 a_1561_989.n3 71.894
R3153 a_1561_989.n2 a_1561_989.n1 71.894
R3154 a_1561_989.n6 a_1561_989.n5 71.555
R3155 a_1561_989.n13 a_1561_989.n11 63.152
R3156 a_1561_989.n11 a_1561_989.n0 16.08
R3157 a_1561_989.n14 a_1561_989.n13 16.078
R3158 a_1561_989.n0 a_1561_989.t6 14.282
R3159 a_1561_989.n0 a_1561_989.t5 14.282
R3160 a_1561_989.n12 a_1561_989.t4 14.282
R3161 a_1561_989.n12 a_1561_989.t3 14.282
R3162 a_1561_989.t1 a_1561_989.n14 14.282
R3163 a_1561_989.n14 a_1561_989.t0 14.282
R3164 a_1561_989.n8 a_1561_989.n7 4.035
R3165 a_7333_989.n3 a_7333_989.t9 454.685
R3166 a_7333_989.n5 a_7333_989.t12 454.685
R3167 a_7333_989.n1 a_7333_989.t10 454.685
R3168 a_7333_989.n3 a_7333_989.t7 428.979
R3169 a_7333_989.n5 a_7333_989.t8 428.979
R3170 a_7333_989.n1 a_7333_989.t15 428.979
R3171 a_7333_989.n4 a_7333_989.t13 264.512
R3172 a_7333_989.n2 a_7333_989.t14 264.512
R3173 a_7333_989.n6 a_7333_989.t11 264.173
R3174 a_7333_989.n10 a_7333_989.n9 261.396
R3175 a_7333_989.n11 a_7333_989.n10 144.246
R3176 a_7333_989.n8 a_7333_989.n2 82.484
R3177 a_7333_989.n7 a_7333_989.n6 79.495
R3178 a_7333_989.n13 a_7333_989.n12 79.232
R3179 a_7333_989.n7 a_7333_989.n4 76
R3180 a_7333_989.n10 a_7333_989.n8 76
R3181 a_7333_989.n4 a_7333_989.n3 71.894
R3182 a_7333_989.n2 a_7333_989.n1 71.894
R3183 a_7333_989.n6 a_7333_989.n5 71.555
R3184 a_7333_989.n13 a_7333_989.n11 63.152
R3185 a_7333_989.n11 a_7333_989.n0 16.08
R3186 a_7333_989.n14 a_7333_989.n13 16.078
R3187 a_7333_989.n0 a_7333_989.t2 14.282
R3188 a_7333_989.n0 a_7333_989.t4 14.282
R3189 a_7333_989.n12 a_7333_989.t5 14.282
R3190 a_7333_989.n12 a_7333_989.t6 14.282
R3191 a_7333_989.n14 a_7333_989.t0 14.282
R3192 a_7333_989.t1 a_7333_989.n14 14.282
R3193 a_7333_989.n8 a_7333_989.n7 4.035
R3194 a_7973_1050.n0 a_7973_1050.t8 512.525
R3195 a_7973_1050.n0 a_7973_1050.t9 371.139
R3196 a_7973_1050.n1 a_7973_1050.t7 234.562
R3197 a_7973_1050.n10 a_7973_1050.n6 223.905
R3198 a_7973_1050.n1 a_7973_1050.n0 215.819
R3199 a_7973_1050.n6 a_7973_1050.n5 159.998
R3200 a_7973_1050.n6 a_7973_1050.n1 153.315
R3201 a_7973_1050.n9 a_7973_1050.n8 79.232
R3202 a_7973_1050.n10 a_7973_1050.n9 63.152
R3203 a_7973_1050.n5 a_7973_1050.n4 30
R3204 a_7973_1050.n3 a_7973_1050.n2 24.383
R3205 a_7973_1050.n5 a_7973_1050.n3 23.684
R3206 a_7973_1050.n9 a_7973_1050.n7 16.08
R3207 a_7973_1050.n11 a_7973_1050.n10 16.078
R3208 a_7973_1050.n7 a_7973_1050.t3 14.282
R3209 a_7973_1050.n7 a_7973_1050.t4 14.282
R3210 a_7973_1050.n8 a_7973_1050.t6 14.282
R3211 a_7973_1050.n8 a_7973_1050.t5 14.282
R3212 a_7973_1050.t1 a_7973_1050.n11 14.282
R3213 a_7973_1050.n11 a_7973_1050.t0 14.282
R3214 a_9897_1050.n2 a_9897_1050.t8 512.525
R3215 a_9897_1050.n2 a_9897_1050.t9 371.139
R3216 a_9897_1050.n3 a_9897_1050.t7 287.668
R3217 a_9897_1050.n8 a_9897_1050.n7 213.104
R3218 a_9897_1050.n9 a_9897_1050.n8 170.799
R3219 a_9897_1050.n3 a_9897_1050.n2 162.713
R3220 a_9897_1050.n8 a_9897_1050.n3 153.315
R3221 a_9897_1050.n11 a_9897_1050.n10 79.231
R3222 a_9897_1050.n10 a_9897_1050.n9 63.152
R3223 a_9897_1050.n7 a_9897_1050.n6 30
R3224 a_9897_1050.n5 a_9897_1050.n4 24.383
R3225 a_9897_1050.n7 a_9897_1050.n5 23.684
R3226 a_9897_1050.n9 a_9897_1050.n1 16.08
R3227 a_9897_1050.n10 a_9897_1050.n0 16.08
R3228 a_9897_1050.n1 a_9897_1050.t5 14.282
R3229 a_9897_1050.n1 a_9897_1050.t4 14.282
R3230 a_9897_1050.n0 a_9897_1050.t6 14.282
R3231 a_9897_1050.n0 a_9897_1050.t0 14.282
R3232 a_9897_1050.n11 a_9897_1050.t1 14.282
R3233 a_9897_1050.t2 a_9897_1050.n11 14.282
R3234 a_18197_1051.n4 a_18197_1051.n3 196.002
R3235 a_18197_1051.n2 a_18197_1051.t4 89.553
R3236 a_18197_1051.n4 a_18197_1051.n0 75.271
R3237 a_18197_1051.n3 a_18197_1051.n2 75.214
R3238 a_18197_1051.n5 a_18197_1051.n4 36.519
R3239 a_18197_1051.n3 a_18197_1051.t2 14.338
R3240 a_18197_1051.n1 a_18197_1051.t5 14.282
R3241 a_18197_1051.n1 a_18197_1051.t3 14.282
R3242 a_18197_1051.n0 a_18197_1051.t6 14.282
R3243 a_18197_1051.n0 a_18197_1051.t7 14.282
R3244 a_18197_1051.t1 a_18197_1051.n5 14.282
R3245 a_18197_1051.n5 a_18197_1051.t0 14.282
R3246 a_18197_1051.n2 a_18197_1051.n1 12.119
R3247 a_17708_209.n1 a_17708_209.t8 512.525
R3248 a_17708_209.n1 a_17708_209.t9 371.139
R3249 a_17708_209.n2 a_17708_209.t7 263.54
R3250 a_17708_209.n13 a_17708_209.n12 216.728
R3251 a_17708_209.n13 a_17708_209.n2 153.043
R3252 a_17708_209.n14 a_17708_209.n13 126.664
R3253 a_17708_209.n2 a_17708_209.n1 120.094
R3254 a_17708_209.n10 a_17708_209.n5 111.94
R3255 a_17708_209.n10 a_17708_209.n9 98.501
R3256 a_17708_209.n12 a_17708_209.n10 78.403
R3257 a_17708_209.n15 a_17708_209.n14 75.27
R3258 a_17708_209.n12 a_17708_209.n11 42.274
R3259 a_17708_209.n9 a_17708_209.n8 30
R3260 a_17708_209.n7 a_17708_209.n6 24.383
R3261 a_17708_209.n9 a_17708_209.n7 23.684
R3262 a_17708_209.n5 a_17708_209.n4 22.578
R3263 a_17708_209.n0 a_17708_209.t4 14.282
R3264 a_17708_209.n0 a_17708_209.t3 14.282
R3265 a_17708_209.n15 a_17708_209.t1 14.282
R3266 a_17708_209.t2 a_17708_209.n15 14.282
R3267 a_17708_209.n14 a_17708_209.n0 12.119
R3268 a_17708_209.n5 a_17708_209.n3 8.58
R3269 RN.n23 RN.t5 479.223
R3270 RN.n17 RN.t21 479.223
R3271 RN.n14 RN.t10 479.223
R3272 RN.n8 RN.t3 479.223
R3273 RN.n5 RN.t15 479.223
R3274 RN.n0 RN.t2 479.223
R3275 RN.n20 RN.t20 454.685
R3276 RN.n11 RN.t0 454.685
R3277 RN.n2 RN.t4 454.685
R3278 RN.n20 RN.t7 428.979
R3279 RN.n11 RN.t17 428.979
R3280 RN.n2 RN.t22 428.979
R3281 RN.n23 RN.t18 375.52
R3282 RN.n17 RN.t9 375.52
R3283 RN.n14 RN.t26 375.52
R3284 RN.n8 RN.t14 375.52
R3285 RN.n5 RN.t19 375.52
R3286 RN.n0 RN.t13 375.52
R3287 RN.n21 RN.n20 178.106
R3288 RN.n12 RN.n11 178.106
R3289 RN.n3 RN.n2 178.106
R3290 RN.n24 RN.n23 175.429
R3291 RN.n18 RN.n17 175.429
R3292 RN.n15 RN.n14 175.429
R3293 RN.n9 RN.n8 175.429
R3294 RN.n6 RN.n5 175.429
R3295 RN.n1 RN.n0 175.429
R3296 RN.n24 RN.t11 162.048
R3297 RN.n18 RN.t23 162.048
R3298 RN.n15 RN.t1 162.048
R3299 RN.n9 RN.t8 162.048
R3300 RN.n6 RN.t6 162.048
R3301 RN.n1 RN.t12 162.048
R3302 RN.n21 RN.t16 158.3
R3303 RN.n12 RN.t25 158.3
R3304 RN.n3 RN.t24 158.3
R3305 RN.n4 RN.n1 78.675
R3306 RN.n4 RN.n3 76
R3307 RN.n7 RN.n6 76
R3308 RN.n10 RN.n9 76
R3309 RN.n13 RN.n12 76
R3310 RN.n16 RN.n15 76
R3311 RN.n19 RN.n18 76
R3312 RN.n22 RN.n21 76
R3313 RN.n25 RN.n24 76
R3314 RN.n7 RN.n4 11.381
R3315 RN.n16 RN.n13 11.381
R3316 RN.n25 RN.n22 11.381
R3317 RN.n10 RN.n7 7.028
R3318 RN.n19 RN.n16 7.028
R3319 RN.n13 RN.n10 2.675
R3320 RN.n22 RN.n19 2.675
R3321 RN.n25 RN 0.046
R3322 a_5863_103.n4 a_5863_103.n3 19.724
R3323 a_5863_103.t0 a_5863_103.n5 11.595
R3324 a_5863_103.t0 a_5863_103.n4 9.207
R3325 a_5863_103.n2 a_5863_103.n0 8.543
R3326 a_5863_103.t0 a_5863_103.n2 3.034
R3327 a_5863_103.n2 a_5863_103.n1 0.443
R3328 a_6144_210.n8 a_6144_210.n6 96.467
R3329 a_6144_210.n3 a_6144_210.n1 44.628
R3330 a_6144_210.t0 a_6144_210.n8 32.417
R3331 a_6144_210.n3 a_6144_210.n2 23.284
R3332 a_6144_210.n6 a_6144_210.n5 22.349
R3333 a_6144_210.t0 a_6144_210.n10 20.241
R3334 a_6144_210.n10 a_6144_210.n9 13.494
R3335 a_6144_210.n6 a_6144_210.n4 8.443
R3336 a_6144_210.t0 a_6144_210.n0 8.137
R3337 a_6144_210.t0 a_6144_210.n3 5.727
R3338 a_6144_210.n8 a_6144_210.n7 1.435
R3339 D.n5 D.t2 512.525
R3340 D.n2 D.t1 512.525
R3341 D.n0 D.t3 512.525
R3342 D.n5 D.t7 371.139
R3343 D.n2 D.t6 371.139
R3344 D.n0 D.t8 371.139
R3345 D.n6 D.t5 340.774
R3346 D.n3 D.t4 340.774
R3347 D.n1 D.t0 340.774
R3348 D.n6 D.n5 109.607
R3349 D.n3 D.n2 109.607
R3350 D.n1 D.n0 109.607
R3351 D.n4 D.n1 97.175
R3352 D.n4 D.n3 76
R3353 D.n7 D.n6 76
R3354 D.n7 D.n4 21.175
R3355 D.n7 D 0.046
R3356 a_11635_103.n4 a_11635_103.n3 19.724
R3357 a_11635_103.t0 a_11635_103.n5 11.595
R3358 a_11635_103.t0 a_11635_103.n4 9.207
R3359 a_11635_103.n2 a_11635_103.n0 8.543
R3360 a_11635_103.t0 a_11635_103.n2 3.034
R3361 a_11635_103.n2 a_11635_103.n1 0.443
R3362 a_16726_210.n9 a_16726_210.n7 82.852
R3363 a_16726_210.n3 a_16726_210.n1 44.628
R3364 a_16726_210.t0 a_16726_210.n9 32.417
R3365 a_16726_210.n7 a_16726_210.n6 27.2
R3366 a_16726_210.n5 a_16726_210.n4 23.498
R3367 a_16726_210.n3 a_16726_210.n2 23.284
R3368 a_16726_210.n7 a_16726_210.n5 22.4
R3369 a_16726_210.t0 a_16726_210.n11 20.241
R3370 a_16726_210.n11 a_16726_210.n10 13.494
R3371 a_16726_210.t0 a_16726_210.n0 8.137
R3372 a_16726_210.t0 a_16726_210.n3 5.727
R3373 a_16726_210.n9 a_16726_210.n8 1.435
R3374 a_7787_103.n1 a_7787_103.n0 25.576
R3375 a_7787_103.n3 a_7787_103.n2 9.111
R3376 a_7787_103.n7 a_7787_103.n5 7.859
R3377 a_7787_103.t0 a_7787_103.n7 3.034
R3378 a_7787_103.n5 a_7787_103.n3 1.964
R3379 a_7787_103.n5 a_7787_103.n4 1.964
R3380 a_7787_103.t0 a_7787_103.n1 1.871
R3381 a_7787_103.n7 a_7787_103.n6 0.443
R3382 a_8068_210.n8 a_8068_210.n6 96.467
R3383 a_8068_210.n3 a_8068_210.n1 44.628
R3384 a_8068_210.t0 a_8068_210.n8 32.417
R3385 a_8068_210.n3 a_8068_210.n2 23.284
R3386 a_8068_210.n6 a_8068_210.n5 22.349
R3387 a_8068_210.t0 a_8068_210.n10 20.241
R3388 a_8068_210.n10 a_8068_210.n9 13.494
R3389 a_8068_210.n6 a_8068_210.n4 8.443
R3390 a_8068_210.t0 a_8068_210.n0 8.137
R3391 a_8068_210.t0 a_8068_210.n3 5.727
R3392 a_8068_210.n8 a_8068_210.n7 1.435
R3393 a_277_1050.n4 a_277_1050.t9 512.525
R3394 a_277_1050.n2 a_277_1050.t7 512.525
R3395 a_277_1050.n4 a_277_1050.t11 371.139
R3396 a_277_1050.n2 a_277_1050.t12 371.139
R3397 a_277_1050.n5 a_277_1050.t10 234.921
R3398 a_277_1050.n3 a_277_1050.t8 234.921
R3399 a_277_1050.n9 a_277_1050.n8 223.546
R3400 a_277_1050.n5 a_277_1050.n4 215.46
R3401 a_277_1050.n3 a_277_1050.n2 215.46
R3402 a_277_1050.n8 a_277_1050.n7 182.096
R3403 a_277_1050.n6 a_277_1050.n3 79.491
R3404 a_277_1050.n11 a_277_1050.n10 79.231
R3405 a_277_1050.n8 a_277_1050.n6 77.315
R3406 a_277_1050.n6 a_277_1050.n5 76
R3407 a_277_1050.n10 a_277_1050.n9 63.152
R3408 a_277_1050.n9 a_277_1050.n1 16.08
R3409 a_277_1050.n10 a_277_1050.n0 16.08
R3410 a_277_1050.n1 a_277_1050.t3 14.282
R3411 a_277_1050.n1 a_277_1050.t4 14.282
R3412 a_277_1050.n0 a_277_1050.t6 14.282
R3413 a_277_1050.n0 a_277_1050.t5 14.282
R3414 a_277_1050.t1 a_277_1050.n11 14.282
R3415 a_277_1050.n11 a_277_1050.t0 14.282
R3416 a_9711_103.n4 a_9711_103.n3 19.724
R3417 a_9711_103.t0 a_9711_103.n5 11.595
R3418 a_9711_103.t0 a_9711_103.n4 9.207
R3419 a_9711_103.n2 a_9711_103.n0 8.543
R3420 a_9711_103.t0 a_9711_103.n2 3.034
R3421 a_9711_103.n2 a_9711_103.n1 0.443
R3422 a_599_989.n2 a_599_989.t12 512.525
R3423 a_599_989.n4 a_599_989.t10 454.685
R3424 a_599_989.n4 a_599_989.t9 428.979
R3425 a_599_989.n2 a_599_989.t8 371.139
R3426 a_599_989.n3 a_599_989.t11 287.668
R3427 a_599_989.n5 a_599_989.t7 237.959
R3428 a_599_989.n11 a_599_989.n10 213.104
R3429 a_599_989.n12 a_599_989.n11 170.799
R3430 a_599_989.n3 a_599_989.n2 162.713
R3431 a_599_989.n5 a_599_989.n4 98.447
R3432 a_599_989.n6 a_599_989.n3 84.388
R3433 a_599_989.n6 a_599_989.n5 80.035
R3434 a_599_989.n14 a_599_989.n13 79.231
R3435 a_599_989.n11 a_599_989.n6 76
R3436 a_599_989.n13 a_599_989.n12 63.152
R3437 a_599_989.n10 a_599_989.n9 30
R3438 a_599_989.n8 a_599_989.n7 24.383
R3439 a_599_989.n10 a_599_989.n8 23.684
R3440 a_599_989.n12 a_599_989.n1 16.08
R3441 a_599_989.n13 a_599_989.n0 16.08
R3442 a_599_989.n1 a_599_989.t5 14.282
R3443 a_599_989.n1 a_599_989.t6 14.282
R3444 a_599_989.n0 a_599_989.t2 14.282
R3445 a_599_989.n0 a_599_989.t3 14.282
R3446 a_599_989.t1 a_599_989.n14 14.282
R3447 a_599_989.n14 a_599_989.t0 14.282
R3448 a_372_210.n9 a_372_210.n7 82.852
R3449 a_372_210.n3 a_372_210.n1 44.628
R3450 a_372_210.t0 a_372_210.n9 32.417
R3451 a_372_210.n7 a_372_210.n6 27.2
R3452 a_372_210.n5 a_372_210.n4 23.498
R3453 a_372_210.n3 a_372_210.n2 23.284
R3454 a_372_210.n7 a_372_210.n5 22.4
R3455 a_372_210.t0 a_372_210.n11 20.241
R3456 a_372_210.n11 a_372_210.n10 13.494
R3457 a_372_210.t0 a_372_210.n0 8.137
R3458 a_372_210.t0 a_372_210.n3 5.727
R3459 a_372_210.n9 a_372_210.n8 1.435
R3460 a_8749_103.n1 a_8749_103.n0 25.576
R3461 a_8749_103.n3 a_8749_103.n2 9.111
R3462 a_8749_103.n7 a_8749_103.n5 7.859
R3463 a_8749_103.t0 a_8749_103.n7 3.034
R3464 a_8749_103.n5 a_8749_103.n3 1.964
R3465 a_8749_103.n5 a_8749_103.n4 1.964
R3466 a_8749_103.t0 a_8749_103.n1 1.871
R3467 a_8749_103.n7 a_8749_103.n6 0.443
R3468 a_9030_210.n10 a_9030_210.n8 82.852
R3469 a_9030_210.n11 a_9030_210.n0 49.6
R3470 a_9030_210.n7 a_9030_210.n6 32.833
R3471 a_9030_210.n8 a_9030_210.t1 32.416
R3472 a_9030_210.n10 a_9030_210.n9 27.2
R3473 a_9030_210.n3 a_9030_210.n2 23.284
R3474 a_9030_210.n11 a_9030_210.n10 22.4
R3475 a_9030_210.n7 a_9030_210.n4 19.017
R3476 a_9030_210.n6 a_9030_210.n5 13.494
R3477 a_9030_210.t1 a_9030_210.n1 7.04
R3478 a_9030_210.t1 a_9030_210.n3 5.727
R3479 a_9030_210.n8 a_9030_210.n7 1.435
R3480 a_12597_103.n1 a_12597_103.n0 25.576
R3481 a_12597_103.n3 a_12597_103.n2 9.111
R3482 a_12597_103.n7 a_12597_103.n5 7.859
R3483 a_12597_103.t0 a_12597_103.n7 3.034
R3484 a_12597_103.n5 a_12597_103.n3 1.964
R3485 a_12597_103.n5 a_12597_103.n4 1.964
R3486 a_12597_103.t0 a_12597_103.n1 1.871
R3487 a_12597_103.n7 a_12597_103.n6 0.443
R3488 a_14521_103.n1 a_14521_103.n0 25.576
R3489 a_14521_103.n3 a_14521_103.n2 9.111
R3490 a_14521_103.n7 a_14521_103.n5 7.859
R3491 a_14521_103.t0 a_14521_103.n7 3.034
R3492 a_14521_103.n5 a_14521_103.n3 1.964
R3493 a_14521_103.n5 a_14521_103.n4 1.964
R3494 a_14521_103.t0 a_14521_103.n1 1.871
R3495 a_14521_103.n7 a_14521_103.n6 0.443
R3496 a_10673_103.n1 a_10673_103.n0 25.576
R3497 a_10673_103.n3 a_10673_103.n2 9.111
R3498 a_10673_103.n7 a_10673_103.n5 7.859
R3499 a_10673_103.t0 a_10673_103.n7 3.034
R3500 a_10673_103.n5 a_10673_103.n3 1.964
R3501 a_10673_103.n5 a_10673_103.n4 1.964
R3502 a_10673_103.t0 a_10673_103.n1 1.871
R3503 a_10673_103.n7 a_10673_103.n6 0.443
R3504 Q.n2 Q.n1 253.86
R3505 Q.n2 Q.n0 130.901
R3506 Q.n3 Q.n2 76
R3507 Q.n0 Q.t2 14.282
R3508 Q.n0 Q.t1 14.282
R3509 Q.n3 Q 0.046
R3510 a_91_103.n5 a_91_103.n4 19.724
R3511 a_91_103.t0 a_91_103.n3 11.595
R3512 a_91_103.t0 a_91_103.n5 9.207
R3513 a_91_103.n2 a_91_103.n1 2.455
R3514 a_91_103.n2 a_91_103.n0 1.32
R3515 a_91_103.t0 a_91_103.n2 0.246
R3516 a_11916_210.n8 a_11916_210.n6 96.467
R3517 a_11916_210.n3 a_11916_210.n1 44.628
R3518 a_11916_210.t0 a_11916_210.n8 32.417
R3519 a_11916_210.n3 a_11916_210.n2 23.284
R3520 a_11916_210.n6 a_11916_210.n5 22.349
R3521 a_11916_210.t0 a_11916_210.n10 20.241
R3522 a_11916_210.n10 a_11916_210.n9 13.494
R3523 a_11916_210.n6 a_11916_210.n4 8.443
R3524 a_11916_210.t0 a_11916_210.n0 8.137
R3525 a_11916_210.t0 a_11916_210.n3 5.727
R3526 a_11916_210.n8 a_11916_210.n7 1.435
R3527 a_9992_210.n8 a_9992_210.n6 96.467
R3528 a_9992_210.n3 a_9992_210.n1 44.628
R3529 a_9992_210.t0 a_9992_210.n8 32.417
R3530 a_9992_210.n3 a_9992_210.n2 23.284
R3531 a_9992_210.n6 a_9992_210.n5 22.349
R3532 a_9992_210.t0 a_9992_210.n10 20.241
R3533 a_9992_210.n10 a_9992_210.n9 13.494
R3534 a_9992_210.n6 a_9992_210.n4 8.443
R3535 a_9992_210.t0 a_9992_210.n0 8.137
R3536 a_9992_210.t0 a_9992_210.n3 5.727
R3537 a_9992_210.n8 a_9992_210.n7 1.435
R3538 a_17428_101.n1 a_17428_101.n0 32.249
R3539 a_17428_101.t0 a_17428_101.n5 7.911
R3540 a_17428_101.n4 a_17428_101.n2 4.032
R3541 a_17428_101.n4 a_17428_101.n3 3.644
R3542 a_17428_101.t0 a_17428_101.n1 2.534
R3543 a_17428_101.t0 a_17428_101.n4 1.099
R3544 a_13559_103.n5 a_13559_103.n4 19.724
R3545 a_13559_103.t0 a_13559_103.n3 11.595
R3546 a_13559_103.t0 a_13559_103.n5 9.207
R3547 a_13559_103.n2 a_13559_103.n1 2.455
R3548 a_13559_103.n2 a_13559_103.n0 1.32
R3549 a_13559_103.t0 a_13559_103.n2 0.246
R3550 a_15483_103.n4 a_15483_103.n3 19.724
R3551 a_15483_103.t0 a_15483_103.n5 11.595
R3552 a_15483_103.t0 a_15483_103.n4 9.207
R3553 a_15483_103.n2 a_15483_103.n0 8.543
R3554 a_15483_103.t0 a_15483_103.n2 3.034
R3555 a_15483_103.n2 a_15483_103.n1 0.443
R3556 a_14802_210.n10 a_14802_210.n8 82.852
R3557 a_14802_210.n11 a_14802_210.n0 49.6
R3558 a_14802_210.n7 a_14802_210.n6 32.833
R3559 a_14802_210.n8 a_14802_210.t1 32.416
R3560 a_14802_210.n10 a_14802_210.n9 27.2
R3561 a_14802_210.n3 a_14802_210.n2 23.284
R3562 a_14802_210.n11 a_14802_210.n10 22.4
R3563 a_14802_210.n7 a_14802_210.n4 19.017
R3564 a_14802_210.n6 a_14802_210.n5 13.494
R3565 a_14802_210.t1 a_14802_210.n1 7.04
R3566 a_14802_210.t1 a_14802_210.n3 5.727
R3567 a_14802_210.n8 a_14802_210.n7 1.435
R3568 a_10954_210.n8 a_10954_210.n6 96.467
R3569 a_10954_210.n3 a_10954_210.n1 44.628
R3570 a_10954_210.t0 a_10954_210.n8 32.417
R3571 a_10954_210.n3 a_10954_210.n2 23.284
R3572 a_10954_210.n6 a_10954_210.n5 22.349
R3573 a_10954_210.t0 a_10954_210.n10 20.241
R3574 a_10954_210.n10 a_10954_210.n9 13.494
R3575 a_10954_210.n6 a_10954_210.n4 8.443
R3576 a_10954_210.t0 a_10954_210.n0 8.137
R3577 a_10954_210.t0 a_10954_210.n3 5.727
R3578 a_10954_210.n8 a_10954_210.n7 1.435
R3579 a_16445_103.n1 a_16445_103.n0 25.576
R3580 a_16445_103.n3 a_16445_103.n2 9.111
R3581 a_16445_103.n7 a_16445_103.n6 2.455
R3582 a_16445_103.n5 a_16445_103.n3 1.964
R3583 a_16445_103.n5 a_16445_103.n4 1.964
R3584 a_16445_103.t0 a_16445_103.n1 1.871
R3585 a_16445_103.n7 a_16445_103.n5 0.636
R3586 a_16445_103.t0 a_16445_103.n7 0.246
R3587 a_12878_210.n10 a_12878_210.n8 82.852
R3588 a_12878_210.n11 a_12878_210.n0 49.6
R3589 a_12878_210.n7 a_12878_210.n6 32.833
R3590 a_12878_210.n8 a_12878_210.t1 32.416
R3591 a_12878_210.n10 a_12878_210.n9 27.2
R3592 a_12878_210.n3 a_12878_210.n2 23.284
R3593 a_12878_210.n11 a_12878_210.n10 22.4
R3594 a_12878_210.n7 a_12878_210.n4 19.017
R3595 a_12878_210.n6 a_12878_210.n5 13.494
R3596 a_12878_210.t1 a_12878_210.n1 7.04
R3597 a_12878_210.t1 a_12878_210.n3 5.727
R3598 a_12878_210.n8 a_12878_210.n7 1.435
R3599 a_2296_210.n10 a_2296_210.n8 82.852
R3600 a_2296_210.n7 a_2296_210.n6 32.833
R3601 a_2296_210.n8 a_2296_210.t1 32.416
R3602 a_2296_210.n10 a_2296_210.n9 27.2
R3603 a_2296_210.n11 a_2296_210.n0 23.498
R3604 a_2296_210.n3 a_2296_210.n2 23.284
R3605 a_2296_210.n11 a_2296_210.n10 22.4
R3606 a_2296_210.n7 a_2296_210.n4 19.017
R3607 a_2296_210.n6 a_2296_210.n5 13.494
R3608 a_2296_210.t1 a_2296_210.n1 7.04
R3609 a_2296_210.t1 a_2296_210.n3 5.727
R3610 a_2296_210.n8 a_2296_210.n7 1.435
R3611 a_4220_210.n9 a_4220_210.n7 82.852
R3612 a_4220_210.n3 a_4220_210.n1 44.628
R3613 a_4220_210.t0 a_4220_210.n9 32.417
R3614 a_4220_210.n7 a_4220_210.n6 27.2
R3615 a_4220_210.n5 a_4220_210.n4 23.498
R3616 a_4220_210.n3 a_4220_210.n2 23.284
R3617 a_4220_210.n7 a_4220_210.n5 22.4
R3618 a_4220_210.t0 a_4220_210.n11 20.241
R3619 a_4220_210.n11 a_4220_210.n10 13.494
R3620 a_4220_210.t0 a_4220_210.n0 8.137
R3621 a_4220_210.t0 a_4220_210.n3 5.727
R3622 a_4220_210.n9 a_4220_210.n8 1.435
R3623 a_15764_210.n8 a_15764_210.n6 96.467
R3624 a_15764_210.n3 a_15764_210.n1 44.628
R3625 a_15764_210.t0 a_15764_210.n8 32.417
R3626 a_15764_210.n3 a_15764_210.n2 23.284
R3627 a_15764_210.n6 a_15764_210.n5 22.349
R3628 a_15764_210.t0 a_15764_210.n10 20.241
R3629 a_15764_210.n10 a_15764_210.n9 13.494
R3630 a_15764_210.n6 a_15764_210.n4 8.443
R3631 a_15764_210.t0 a_15764_210.n0 8.137
R3632 a_15764_210.t0 a_15764_210.n3 5.727
R3633 a_15764_210.n8 a_15764_210.n7 1.435
R3634 a_2015_103.n5 a_2015_103.n4 19.724
R3635 a_2015_103.t0 a_2015_103.n3 11.595
R3636 a_2015_103.t0 a_2015_103.n5 9.207
R3637 a_2015_103.n2 a_2015_103.n1 2.455
R3638 a_2015_103.n2 a_2015_103.n0 1.32
R3639 a_2015_103.t0 a_2015_103.n2 0.246
R3640 a_1334_210.n10 a_1334_210.n8 82.852
R3641 a_1334_210.n7 a_1334_210.n6 32.833
R3642 a_1334_210.n8 a_1334_210.t1 32.416
R3643 a_1334_210.n10 a_1334_210.n9 27.2
R3644 a_1334_210.n11 a_1334_210.n0 23.498
R3645 a_1334_210.n3 a_1334_210.n2 23.284
R3646 a_1334_210.n11 a_1334_210.n10 22.4
R3647 a_1334_210.n7 a_1334_210.n4 19.017
R3648 a_1334_210.n6 a_1334_210.n5 13.494
R3649 a_1334_210.t1 a_1334_210.n1 7.04
R3650 a_1334_210.t1 a_1334_210.n3 5.727
R3651 a_1334_210.n8 a_1334_210.n7 1.435
R3652 a_7106_210.n10 a_7106_210.n8 82.852
R3653 a_7106_210.n11 a_7106_210.n0 49.6
R3654 a_7106_210.n7 a_7106_210.n6 32.833
R3655 a_7106_210.n8 a_7106_210.t1 32.416
R3656 a_7106_210.n10 a_7106_210.n9 27.2
R3657 a_7106_210.n3 a_7106_210.n2 23.284
R3658 a_7106_210.n11 a_7106_210.n10 22.4
R3659 a_7106_210.n7 a_7106_210.n4 19.017
R3660 a_7106_210.n6 a_7106_210.n5 13.494
R3661 a_7106_210.t1 a_7106_210.n1 7.04
R3662 a_7106_210.t1 a_7106_210.n3 5.727
R3663 a_7106_210.n8 a_7106_210.n7 1.435
R3664 a_5182_210.n10 a_5182_210.n8 82.852
R3665 a_5182_210.n11 a_5182_210.n0 49.6
R3666 a_5182_210.n7 a_5182_210.n6 32.833
R3667 a_5182_210.n8 a_5182_210.t1 32.416
R3668 a_5182_210.n10 a_5182_210.n9 27.2
R3669 a_5182_210.n3 a_5182_210.n2 23.284
R3670 a_5182_210.n11 a_5182_210.n10 22.4
R3671 a_5182_210.n7 a_5182_210.n4 19.017
R3672 a_5182_210.n6 a_5182_210.n5 13.494
R3673 a_5182_210.t1 a_5182_210.n1 7.04
R3674 a_5182_210.t1 a_5182_210.n3 5.727
R3675 a_5182_210.n8 a_5182_210.n7 1.435
R3676 a_1053_103.n5 a_1053_103.n4 19.724
R3677 a_1053_103.t0 a_1053_103.n3 11.595
R3678 a_1053_103.t0 a_1053_103.n5 9.207
R3679 a_1053_103.n2 a_1053_103.n1 2.455
R3680 a_1053_103.n2 a_1053_103.n0 1.32
R3681 a_1053_103.t0 a_1053_103.n2 0.246
R3682 a_3939_103.n5 a_3939_103.n4 19.724
R3683 a_3939_103.t0 a_3939_103.n3 11.595
R3684 a_3939_103.t0 a_3939_103.n5 9.207
R3685 a_3939_103.n2 a_3939_103.n1 2.455
R3686 a_3939_103.n2 a_3939_103.n0 1.32
R3687 a_3939_103.t0 a_3939_103.n2 0.246
C11 SN GND 9.66fF
C12 RN GND 11.16fF
C13 VDD GND 70.77fF
C14 a_3939_103.n0 GND 0.10fF
C15 a_3939_103.n1 GND 0.04fF
C16 a_3939_103.n2 GND 0.03fF
C17 a_3939_103.n3 GND 0.07fF
C18 a_3939_103.n4 GND 0.08fF
C19 a_3939_103.n5 GND 0.06fF
C20 a_1053_103.n0 GND 0.10fF
C21 a_1053_103.n1 GND 0.04fF
C22 a_1053_103.n2 GND 0.03fF
C23 a_1053_103.n3 GND 0.07fF
C24 a_1053_103.n4 GND 0.08fF
C25 a_1053_103.n5 GND 0.06fF
C26 a_5182_210.n0 GND 0.02fF
C27 a_5182_210.n1 GND 0.09fF
C28 a_5182_210.n2 GND 0.13fF
C29 a_5182_210.n3 GND 0.11fF
C30 a_5182_210.t1 GND 0.30fF
C31 a_5182_210.n4 GND 0.09fF
C32 a_5182_210.n5 GND 0.06fF
C33 a_5182_210.n6 GND 0.01fF
C34 a_5182_210.n7 GND 0.03fF
C35 a_5182_210.n8 GND 0.11fF
C36 a_5182_210.n9 GND 0.02fF
C37 a_5182_210.n10 GND 0.05fF
C38 a_5182_210.n11 GND 0.02fF
C39 a_7106_210.n0 GND 0.02fF
C40 a_7106_210.n1 GND 0.09fF
C41 a_7106_210.n2 GND 0.13fF
C42 a_7106_210.n3 GND 0.11fF
C43 a_7106_210.t1 GND 0.30fF
C44 a_7106_210.n4 GND 0.09fF
C45 a_7106_210.n5 GND 0.06fF
C46 a_7106_210.n6 GND 0.01fF
C47 a_7106_210.n7 GND 0.03fF
C48 a_7106_210.n8 GND 0.11fF
C49 a_7106_210.n9 GND 0.02fF
C50 a_7106_210.n10 GND 0.05fF
C51 a_7106_210.n11 GND 0.02fF
C52 a_1334_210.n0 GND 0.02fF
C53 a_1334_210.n1 GND 0.09fF
C54 a_1334_210.n2 GND 0.13fF
C55 a_1334_210.n3 GND 0.11fF
C56 a_1334_210.t1 GND 0.30fF
C57 a_1334_210.n4 GND 0.09fF
C58 a_1334_210.n5 GND 0.06fF
C59 a_1334_210.n6 GND 0.01fF
C60 a_1334_210.n7 GND 0.03fF
C61 a_1334_210.n8 GND 0.11fF
C62 a_1334_210.n9 GND 0.02fF
C63 a_1334_210.n10 GND 0.05fF
C64 a_1334_210.n11 GND 0.03fF
C65 a_2015_103.n0 GND 0.10fF
C66 a_2015_103.n1 GND 0.04fF
C67 a_2015_103.n2 GND 0.03fF
C68 a_2015_103.n3 GND 0.07fF
C69 a_2015_103.n4 GND 0.08fF
C70 a_2015_103.n5 GND 0.06fF
C71 a_15764_210.n0 GND 0.07fF
C72 a_15764_210.n1 GND 0.09fF
C73 a_15764_210.n2 GND 0.13fF
C74 a_15764_210.n3 GND 0.11fF
C75 a_15764_210.n4 GND 0.02fF
C76 a_15764_210.n5 GND 0.03fF
C77 a_15764_210.n6 GND 0.06fF
C78 a_15764_210.n7 GND 0.03fF
C79 a_15764_210.n8 GND 0.12fF
C80 a_15764_210.n9 GND 0.06fF
C81 a_15764_210.n10 GND 0.01fF
C82 a_15764_210.t0 GND 0.33fF
C83 a_4220_210.n0 GND 0.07fF
C84 a_4220_210.n1 GND 0.09fF
C85 a_4220_210.n2 GND 0.13fF
C86 a_4220_210.n3 GND 0.11fF
C87 a_4220_210.n4 GND 0.02fF
C88 a_4220_210.n5 GND 0.03fF
C89 a_4220_210.n6 GND 0.02fF
C90 a_4220_210.n7 GND 0.05fF
C91 a_4220_210.n8 GND 0.03fF
C92 a_4220_210.n9 GND 0.11fF
C93 a_4220_210.n10 GND 0.06fF
C94 a_4220_210.n11 GND 0.01fF
C95 a_4220_210.t0 GND 0.33fF
C96 a_2296_210.n0 GND 0.02fF
C97 a_2296_210.n1 GND 0.09fF
C98 a_2296_210.n2 GND 0.13fF
C99 a_2296_210.n3 GND 0.11fF
C100 a_2296_210.t1 GND 0.30fF
C101 a_2296_210.n4 GND 0.09fF
C102 a_2296_210.n5 GND 0.06fF
C103 a_2296_210.n6 GND 0.01fF
C104 a_2296_210.n7 GND 0.03fF
C105 a_2296_210.n8 GND 0.11fF
C106 a_2296_210.n9 GND 0.02fF
C107 a_2296_210.n10 GND 0.05fF
C108 a_2296_210.n11 GND 0.03fF
C109 a_12878_210.n0 GND 0.02fF
C110 a_12878_210.n1 GND 0.09fF
C111 a_12878_210.n2 GND 0.13fF
C112 a_12878_210.n3 GND 0.11fF
C113 a_12878_210.t1 GND 0.30fF
C114 a_12878_210.n4 GND 0.09fF
C115 a_12878_210.n5 GND 0.06fF
C116 a_12878_210.n6 GND 0.01fF
C117 a_12878_210.n7 GND 0.03fF
C118 a_12878_210.n8 GND 0.11fF
C119 a_12878_210.n9 GND 0.02fF
C120 a_12878_210.n10 GND 0.05fF
C121 a_12878_210.n11 GND 0.02fF
C122 a_16445_103.n0 GND 0.09fF
C123 a_16445_103.n1 GND 0.10fF
C124 a_16445_103.n2 GND 0.05fF
C125 a_16445_103.n3 GND 0.03fF
C126 a_16445_103.n4 GND 0.04fF
C127 a_16445_103.n5 GND 0.03fF
C128 a_16445_103.n6 GND 0.04fF
C129 a_10954_210.n0 GND 0.07fF
C130 a_10954_210.n1 GND 0.09fF
C131 a_10954_210.n2 GND 0.13fF
C132 a_10954_210.n3 GND 0.11fF
C133 a_10954_210.n4 GND 0.02fF
C134 a_10954_210.n5 GND 0.03fF
C135 a_10954_210.n6 GND 0.06fF
C136 a_10954_210.n7 GND 0.03fF
C137 a_10954_210.n8 GND 0.12fF
C138 a_10954_210.n9 GND 0.06fF
C139 a_10954_210.n10 GND 0.01fF
C140 a_10954_210.t0 GND 0.33fF
C141 a_14802_210.n0 GND 0.02fF
C142 a_14802_210.n1 GND 0.09fF
C143 a_14802_210.n2 GND 0.13fF
C144 a_14802_210.n3 GND 0.11fF
C145 a_14802_210.t1 GND 0.30fF
C146 a_14802_210.n4 GND 0.09fF
C147 a_14802_210.n5 GND 0.06fF
C148 a_14802_210.n6 GND 0.01fF
C149 a_14802_210.n7 GND 0.03fF
C150 a_14802_210.n8 GND 0.11fF
C151 a_14802_210.n9 GND 0.02fF
C152 a_14802_210.n10 GND 0.05fF
C153 a_14802_210.n11 GND 0.02fF
C154 a_15483_103.n0 GND 0.20fF
C155 a_15483_103.n1 GND 0.04fF
C156 a_15483_103.n2 GND 0.01fF
C157 a_15483_103.n3 GND 0.08fF
C158 a_15483_103.n4 GND 0.06fF
C159 a_15483_103.n5 GND 0.07fF
C160 a_13559_103.n0 GND 0.10fF
C161 a_13559_103.n1 GND 0.04fF
C162 a_13559_103.n2 GND 0.03fF
C163 a_13559_103.n3 GND 0.07fF
C164 a_13559_103.n4 GND 0.08fF
C165 a_13559_103.n5 GND 0.06fF
C166 a_17428_101.n0 GND 0.11fF
C167 a_17428_101.n1 GND 0.09fF
C168 a_17428_101.n2 GND 0.08fF
C169 a_17428_101.n3 GND 0.02fF
C170 a_17428_101.n4 GND 0.01fF
C171 a_17428_101.n5 GND 0.06fF
C172 a_9992_210.n0 GND 0.07fF
C173 a_9992_210.n1 GND 0.09fF
C174 a_9992_210.n2 GND 0.13fF
C175 a_9992_210.n3 GND 0.11fF
C176 a_9992_210.n4 GND 0.02fF
C177 a_9992_210.n5 GND 0.03fF
C178 a_9992_210.n6 GND 0.06fF
C179 a_9992_210.n7 GND 0.03fF
C180 a_9992_210.n8 GND 0.12fF
C181 a_9992_210.n9 GND 0.06fF
C182 a_9992_210.n10 GND 0.01fF
C183 a_9992_210.t0 GND 0.33fF
C184 a_11916_210.n0 GND 0.07fF
C185 a_11916_210.n1 GND 0.09fF
C186 a_11916_210.n2 GND 0.13fF
C187 a_11916_210.n3 GND 0.11fF
C188 a_11916_210.n4 GND 0.02fF
C189 a_11916_210.n5 GND 0.03fF
C190 a_11916_210.n6 GND 0.06fF
C191 a_11916_210.n7 GND 0.03fF
C192 a_11916_210.n8 GND 0.12fF
C193 a_11916_210.n9 GND 0.06fF
C194 a_11916_210.n10 GND 0.01fF
C195 a_11916_210.t0 GND 0.33fF
C196 a_91_103.n0 GND 0.10fF
C197 a_91_103.n1 GND 0.04fF
C198 a_91_103.n2 GND 0.03fF
C199 a_91_103.n3 GND 0.06fF
C200 a_91_103.n4 GND 0.08fF
C201 a_91_103.n5 GND 0.06fF
C202 Q.n0 GND 0.75fF
C203 Q.n1 GND 0.45fF
C204 Q.n2 GND 0.51fF
C205 Q.n3 GND 0.01fF
C206 a_10673_103.n0 GND 0.09fF
C207 a_10673_103.n1 GND 0.10fF
C208 a_10673_103.n2 GND 0.05fF
C209 a_10673_103.n3 GND 0.03fF
C210 a_10673_103.n4 GND 0.04fF
C211 a_10673_103.n5 GND 0.11fF
C212 a_10673_103.n6 GND 0.04fF
C213 a_14521_103.n0 GND 0.09fF
C214 a_14521_103.n1 GND 0.10fF
C215 a_14521_103.n2 GND 0.05fF
C216 a_14521_103.n3 GND 0.03fF
C217 a_14521_103.n4 GND 0.04fF
C218 a_14521_103.n5 GND 0.11fF
C219 a_14521_103.n6 GND 0.04fF
C220 a_12597_103.n0 GND 0.09fF
C221 a_12597_103.n1 GND 0.10fF
C222 a_12597_103.n2 GND 0.05fF
C223 a_12597_103.n3 GND 0.03fF
C224 a_12597_103.n4 GND 0.04fF
C225 a_12597_103.n5 GND 0.11fF
C226 a_12597_103.n6 GND 0.04fF
C227 a_9030_210.n0 GND 0.02fF
C228 a_9030_210.n1 GND 0.09fF
C229 a_9030_210.n2 GND 0.13fF
C230 a_9030_210.n3 GND 0.11fF
C231 a_9030_210.t1 GND 0.30fF
C232 a_9030_210.n4 GND 0.09fF
C233 a_9030_210.n5 GND 0.06fF
C234 a_9030_210.n6 GND 0.01fF
C235 a_9030_210.n7 GND 0.03fF
C236 a_9030_210.n8 GND 0.11fF
C237 a_9030_210.n9 GND 0.02fF
C238 a_9030_210.n10 GND 0.05fF
C239 a_9030_210.n11 GND 0.02fF
C240 a_8749_103.n0 GND 0.09fF
C241 a_8749_103.n1 GND 0.10fF
C242 a_8749_103.n2 GND 0.05fF
C243 a_8749_103.n3 GND 0.03fF
C244 a_8749_103.n4 GND 0.04fF
C245 a_8749_103.n5 GND 0.11fF
C246 a_8749_103.n6 GND 0.04fF
C247 a_372_210.n0 GND 0.07fF
C248 a_372_210.n1 GND 0.09fF
C249 a_372_210.n2 GND 0.13fF
C250 a_372_210.n3 GND 0.11fF
C251 a_372_210.n4 GND 0.02fF
C252 a_372_210.n5 GND 0.03fF
C253 a_372_210.n6 GND 0.02fF
C254 a_372_210.n7 GND 0.05fF
C255 a_372_210.n8 GND 0.03fF
C256 a_372_210.n9 GND 0.11fF
C257 a_372_210.n10 GND 0.06fF
C258 a_372_210.n11 GND 0.01fF
C259 a_372_210.t0 GND 0.33fF
C260 a_599_989.n0 GND 0.74fF
C261 a_599_989.n1 GND 0.74fF
C262 a_599_989.n2 GND 0.46fF
C263 a_599_989.n3 GND 0.79fF
C264 a_599_989.n4 GND 0.52fF
C265 a_599_989.t7 GND 0.74fF
C266 a_599_989.n5 GND 0.54fF
C267 a_599_989.n6 GND 3.76fF
C268 a_599_989.n7 GND 0.06fF
C269 a_599_989.n8 GND 0.07fF
C270 a_599_989.n9 GND 0.05fF
C271 a_599_989.n10 GND 0.42fF
C272 a_599_989.n11 GND 0.62fF
C273 a_599_989.n12 GND 0.42fF
C274 a_599_989.n13 GND 0.27fF
C275 a_599_989.n14 GND 0.87fF
C276 a_9711_103.n0 GND 0.20fF
C277 a_9711_103.n1 GND 0.04fF
C278 a_9711_103.n2 GND 0.01fF
C279 a_9711_103.n3 GND 0.08fF
C280 a_9711_103.n4 GND 0.06fF
C281 a_9711_103.n5 GND 0.07fF
C282 a_277_1050.n0 GND 0.54fF
C283 a_277_1050.n1 GND 0.54fF
C284 a_277_1050.n2 GND 0.40fF
C285 a_277_1050.n3 GND 0.49fF
C286 a_277_1050.n4 GND 0.40fF
C287 a_277_1050.n5 GND 0.47fF
C288 a_277_1050.n6 GND 1.14fF
C289 a_277_1050.n7 GND 0.34fF
C290 a_277_1050.n8 GND 0.49fF
C291 a_277_1050.n9 GND 0.37fF
C292 a_277_1050.n10 GND 0.20fF
C293 a_277_1050.n11 GND 0.64fF
C294 a_8068_210.n0 GND 0.07fF
C295 a_8068_210.n1 GND 0.09fF
C296 a_8068_210.n2 GND 0.13fF
C297 a_8068_210.n3 GND 0.11fF
C298 a_8068_210.n4 GND 0.02fF
C299 a_8068_210.n5 GND 0.03fF
C300 a_8068_210.n6 GND 0.06fF
C301 a_8068_210.n7 GND 0.03fF
C302 a_8068_210.n8 GND 0.12fF
C303 a_8068_210.n9 GND 0.06fF
C304 a_8068_210.n10 GND 0.01fF
C305 a_8068_210.t0 GND 0.33fF
C306 a_7787_103.n0 GND 0.09fF
C307 a_7787_103.n1 GND 0.10fF
C308 a_7787_103.n2 GND 0.05fF
C309 a_7787_103.n3 GND 0.03fF
C310 a_7787_103.n4 GND 0.04fF
C311 a_7787_103.n5 GND 0.11fF
C312 a_7787_103.n6 GND 0.04fF
C313 a_16726_210.n0 GND 0.07fF
C314 a_16726_210.n1 GND 0.09fF
C315 a_16726_210.n2 GND 0.13fF
C316 a_16726_210.n3 GND 0.11fF
C317 a_16726_210.n4 GND 0.02fF
C318 a_16726_210.n5 GND 0.03fF
C319 a_16726_210.n6 GND 0.02fF
C320 a_16726_210.n7 GND 0.05fF
C321 a_16726_210.n8 GND 0.03fF
C322 a_16726_210.n9 GND 0.11fF
C323 a_16726_210.n10 GND 0.06fF
C324 a_16726_210.n11 GND 0.01fF
C325 a_16726_210.t0 GND 0.33fF
C326 a_11635_103.n0 GND 0.20fF
C327 a_11635_103.n1 GND 0.04fF
C328 a_11635_103.n2 GND 0.01fF
C329 a_11635_103.n3 GND 0.08fF
C330 a_11635_103.n4 GND 0.06fF
C331 a_11635_103.n5 GND 0.07fF
C332 a_6144_210.n0 GND 0.07fF
C333 a_6144_210.n1 GND 0.09fF
C334 a_6144_210.n2 GND 0.13fF
C335 a_6144_210.n3 GND 0.11fF
C336 a_6144_210.n4 GND 0.02fF
C337 a_6144_210.n5 GND 0.03fF
C338 a_6144_210.n6 GND 0.06fF
C339 a_6144_210.n7 GND 0.03fF
C340 a_6144_210.n8 GND 0.12fF
C341 a_6144_210.n9 GND 0.06fF
C342 a_6144_210.n10 GND 0.01fF
C343 a_6144_210.t0 GND 0.33fF
C344 a_5863_103.n0 GND 0.20fF
C345 a_5863_103.n1 GND 0.04fF
C346 a_5863_103.n2 GND 0.01fF
C347 a_5863_103.n3 GND 0.08fF
C348 a_5863_103.n4 GND 0.06fF
C349 a_5863_103.n5 GND 0.07fF
C350 RN.n0 GND 0.92fF
C351 RN.t12 GND 0.84fF
C352 RN.n1 GND 0.71fF
C353 RN.n2 GND 0.90fF
C354 RN.t24 GND 0.86fF
C355 RN.n3 GND 0.69fF
C356 RN.n4 GND 3.65fF
C357 RN.n5 GND 0.92fF
C358 RN.t6 GND 0.84fF
C359 RN.n6 GND 0.69fF
C360 RN.n7 GND 3.96fF
C361 RN.n8 GND 0.92fF
C362 RN.t8 GND 0.84fF
C363 RN.n9 GND 0.69fF
C364 RN.n10 GND 2.11fF
C365 RN.n11 GND 0.90fF
C366 RN.t25 GND 0.86fF
C367 RN.n12 GND 0.69fF
C368 RN.n13 GND 3.04fF
C369 RN.n14 GND 0.92fF
C370 RN.t1 GND 0.84fF
C371 RN.n15 GND 0.69fF
C372 RN.n16 GND 3.96fF
C373 RN.n17 GND 0.92fF
C374 RN.t23 GND 0.84fF
C375 RN.n18 GND 0.69fF
C376 RN.n19 GND 2.11fF
C377 RN.n20 GND 0.90fF
C378 RN.t16 GND 0.86fF
C379 RN.n21 GND 0.69fF
C380 RN.n22 GND 3.04fF
C381 RN.n23 GND 0.92fF
C382 RN.t11 GND 0.84fF
C383 RN.n24 GND 0.69fF
C384 RN.n25 GND 2.46fF
C385 a_17708_209.n0 GND 0.37fF
C386 a_17708_209.n1 GND 0.26fF
C387 a_17708_209.n2 GND 0.48fF
C388 a_17708_209.n3 GND 0.04fF
C389 a_17708_209.n4 GND 0.04fF
C390 a_17708_209.n5 GND 0.10fF
C391 a_17708_209.n6 GND 0.03fF
C392 a_17708_209.n7 GND 0.04fF
C393 a_17708_209.n8 GND 0.03fF
C394 a_17708_209.n9 GND 0.09fF
C395 a_17708_209.n10 GND 0.97fF
C396 a_17708_209.n11 GND 0.12fF
C397 a_17708_209.n12 GND 0.29fF
C398 a_17708_209.n13 GND 0.45fF
C399 a_17708_209.n14 GND 0.23fF
C400 a_17708_209.n15 GND 0.45fF
C401 a_18197_1051.n0 GND 0.36fF
C402 a_18197_1051.n1 GND 0.29fF
C403 a_18197_1051.n2 GND 0.20fF
C404 a_18197_1051.n3 GND 0.57fF
C405 a_18197_1051.n4 GND 0.25fF
C406 a_18197_1051.n5 GND 0.28fF
C407 a_9897_1050.n0 GND 0.57fF
C408 a_9897_1050.n1 GND 0.57fF
C409 a_9897_1050.n2 GND 0.36fF
C410 a_9897_1050.n3 GND 0.69fF
C411 a_9897_1050.n4 GND 0.04fF
C412 a_9897_1050.n5 GND 0.06fF
C413 a_9897_1050.n6 GND 0.04fF
C414 a_9897_1050.n7 GND 0.32fF
C415 a_9897_1050.n8 GND 0.66fF
C416 a_9897_1050.n9 GND 0.32fF
C417 a_9897_1050.n10 GND 0.21fF
C418 a_9897_1050.n11 GND 0.67fF
C419 a_7973_1050.n0 GND 0.42fF
C420 a_7973_1050.n1 GND 0.67fF
C421 a_7973_1050.n2 GND 0.04fF
C422 a_7973_1050.n3 GND 0.06fF
C423 a_7973_1050.n4 GND 0.04fF
C424 a_7973_1050.n5 GND 0.25fF
C425 a_7973_1050.n6 GND 0.66fF
C426 a_7973_1050.n7 GND 0.56fF
C427 a_7973_1050.n8 GND 0.66fF
C428 a_7973_1050.n9 GND 0.21fF
C429 a_7973_1050.n10 GND 0.39fF
C430 a_7973_1050.n11 GND 0.56fF
C431 a_7333_989.n0 GND 0.95fF
C432 a_7333_989.n1 GND 0.61fF
C433 a_7333_989.t14 GND 1.00fF
C434 a_7333_989.n2 GND 0.76fF
C435 a_7333_989.n3 GND 0.61fF
C436 a_7333_989.t13 GND 1.00fF
C437 a_7333_989.n4 GND 0.66fF
C438 a_7333_989.n5 GND 0.61fF
C439 a_7333_989.t11 GND 1.00fF
C440 a_7333_989.n6 GND 0.69fF
C441 a_7333_989.n7 GND 2.24fF
C442 a_7333_989.n8 GND 3.34fF
C443 a_7333_989.n9 GND 0.77fF
C444 a_7333_989.n10 GND 0.85fF
C445 a_7333_989.n11 GND 0.49fF
C446 a_7333_989.n12 GND 1.12fF
C447 a_7333_989.n13 GND 0.35fF
C448 a_7333_989.n14 GND 0.95fF
C449 a_1561_989.n0 GND 0.88fF
C450 a_1561_989.n1 GND 0.56fF
C451 a_1561_989.t12 GND 0.92fF
C452 a_1561_989.n2 GND 0.70fF
C453 a_1561_989.n3 GND 0.56fF
C454 a_1561_989.t9 GND 0.92fF
C455 a_1561_989.n4 GND 0.61fF
C456 a_1561_989.n5 GND 0.56fF
C457 a_1561_989.t10 GND 0.92fF
C458 a_1561_989.n6 GND 0.64fF
C459 a_1561_989.n7 GND 2.06fF
C460 a_1561_989.n8 GND 3.08fF
C461 a_1561_989.n9 GND 0.70fF
C462 a_1561_989.n10 GND 0.79fF
C463 a_1561_989.n11 GND 0.45fF
C464 a_1561_989.n12 GND 1.03fF
C465 a_1561_989.n13 GND 0.32fF
C466 a_1561_989.n14 GND 0.88fF
C467 a_2201_1050.n0 GND 0.51fF
C468 a_2201_1050.n1 GND 0.38fF
C469 a_2201_1050.n2 GND 0.61fF
C470 a_2201_1050.n3 GND 0.32fF
C471 a_2201_1050.n4 GND 0.63fF
C472 a_2201_1050.n5 GND 0.35fF
C473 a_2201_1050.n6 GND 0.60fF
C474 a_2201_1050.n7 GND 0.19fF
C475 a_2201_1050.n8 GND 0.51fF
C476 a_18094_101.n0 GND 0.13fF
C477 a_18094_101.n1 GND 0.15fF
C478 a_18760_101.n0 GND 0.06fF
C479 a_18760_101.n1 GND 0.14fF
C480 a_18760_101.n2 GND 0.04fF
C481 a_4447_989.n0 GND 1.21fF
C482 a_4447_989.n1 GND 1.21fF
C483 a_4447_989.n2 GND 0.86fF
C484 a_4447_989.n3 GND 1.06fF
C485 a_4447_989.n4 GND 1.31fF
C486 a_4447_989.t11 GND 0.99fF
C487 a_4447_989.n5 GND 0.82fF
C488 a_4447_989.n6 GND 5.26fF
C489 a_4447_989.n7 GND 0.92fF
C490 a_4447_989.t12 GND 1.15fF
C491 a_4447_989.n8 GND 0.86fF
C492 a_4447_989.n9 GND 21.24fF
C493 a_4447_989.n10 GND 0.10fF
C494 a_4447_989.n11 GND 0.12fF
C495 a_4447_989.n12 GND 0.63fF
C496 a_4447_989.n13 GND 1.07fF
C497 a_4447_989.n14 GND 0.76fF
C498 a_4447_989.n15 GND 0.45fF
C499 a_4447_989.n16 GND 1.42fF
C500 a_6371_989.n0 GND 0.98fF
C501 a_6371_989.n1 GND 0.62fF
C502 a_6371_989.n2 GND 1.05fF
C503 a_6371_989.n3 GND 0.69fF
C504 a_6371_989.t11 GND 0.98fF
C505 a_6371_989.n4 GND 0.72fF
C506 a_6371_989.n5 GND 4.99fF
C507 a_6371_989.n6 GND 0.73fF
C508 a_6371_989.n7 GND 0.88fF
C509 a_6371_989.n8 GND 0.56fF
C510 a_6371_989.n9 GND 1.15fF
C511 a_6371_989.n10 GND 0.36fF
C512 a_6371_989.n11 GND 0.98fF
C513 SN.n0 GND 0.97fF
C514 SN.t9 GND 0.79fF
C515 SN.n1 GND 0.94fF
C516 SN.n2 GND 0.96fF
C517 SN.t11 GND 0.78fF
C518 SN.n3 GND 0.68fF
C519 SN.n4 GND 6.47fF
C520 SN.n5 GND 0.97fF
C521 SN.t8 GND 0.79fF
C522 SN.n6 GND 0.66fF
C523 SN.n7 GND 4.47fF
C524 SN.n8 GND 0.96fF
C525 SN.t3 GND 0.78fF
C526 SN.n9 GND 0.68fF
C527 SN.n10 GND 4.47fF
C528 SN.n11 GND 0.97fF
C529 SN.t17 GND 0.79fF
C530 SN.n12 GND 0.66fF
C531 SN.n13 GND 4.47fF
C532 SN.t16 GND 0.78fF
C533 SN.n14 GND 0.96fF
C534 SN.n15 GND 0.68fF
C535 SN.n16 GND 2.26fF
C536 a_4901_103.n0 GND 0.10fF
C537 a_4901_103.n1 GND 0.04fF
C538 a_4901_103.n2 GND 0.03fF
C539 a_4901_103.n3 GND 0.07fF
C540 a_4901_103.n4 GND 0.08fF
C541 a_4901_103.n5 GND 0.06fF
C542 a_4125_1050.n0 GND 0.55fF
C543 a_4125_1050.n1 GND 0.55fF
C544 a_4125_1050.n2 GND 0.64fF
C545 a_4125_1050.n3 GND 0.20fF
C546 a_4125_1050.n4 GND 0.31fF
C547 a_4125_1050.n5 GND 0.34fF
C548 a_4125_1050.n6 GND 0.67fF
C549 a_4125_1050.n7 GND 0.65fF
C550 a_4125_1050.n8 GND 0.08fF
C551 a_4125_1050.n9 GND 0.30fF
C552 a_4125_1050.n10 GND 0.05fF
C553 a_12143_989.n0 GND 0.97fF
C554 a_12143_989.n1 GND 0.61fF
C555 a_12143_989.n2 GND 1.04fF
C556 a_12143_989.n3 GND 0.68fF
C557 a_12143_989.t11 GND 0.97fF
C558 a_12143_989.n4 GND 0.71fF
C559 a_12143_989.n5 GND 4.93fF
C560 a_12143_989.n6 GND 0.07fF
C561 a_12143_989.n7 GND 0.10fF
C562 a_12143_989.n8 GND 0.06fF
C563 a_12143_989.n9 GND 0.55fF
C564 a_12143_989.n10 GND 0.81fF
C565 a_12143_989.n11 GND 0.55fF
C566 a_12143_989.n12 GND 1.14fF
C567 a_12143_989.n13 GND 0.36fF
C568 a_12143_989.n14 GND 0.97fF
C569 a_11821_1050.n0 GND 0.71fF
C570 a_11821_1050.n1 GND 0.71fF
C571 a_11821_1050.n2 GND 0.83fF
C572 a_11821_1050.n3 GND 0.26fF
C573 a_11821_1050.n4 GND 0.48fF
C574 a_11821_1050.n5 GND 0.52fF
C575 a_11821_1050.n6 GND 0.64fF
C576 a_11821_1050.n7 GND 0.52fF
C577 a_11821_1050.n8 GND 0.61fF
C578 a_11821_1050.n9 GND 1.49fF
C579 a_11821_1050.n10 GND 0.61fF
C580 a_11821_1050.n11 GND 0.11fF
C581 a_11821_1050.n12 GND 0.30fF
C582 a_11821_1050.n13 GND 0.06fF
C583 a_15669_1050.n0 GND 0.34fF
C584 a_15669_1050.n1 GND 0.65fF
C585 a_15669_1050.n2 GND 0.04fF
C586 a_15669_1050.n3 GND 0.05fF
C587 a_15669_1050.n4 GND 0.03fF
C588 a_15669_1050.n5 GND 0.30fF
C589 a_15669_1050.n6 GND 0.63fF
C590 a_15669_1050.n7 GND 0.53fF
C591 a_15669_1050.n8 GND 0.63fF
C592 a_15669_1050.n9 GND 0.20fF
C593 a_15669_1050.n10 GND 0.31fF
C594 a_15669_1050.n11 GND 0.53fF
C595 a_15991_989.n0 GND 0.29fF
C596 a_15991_989.n1 GND 0.78fF
C597 a_15991_989.n2 GND 0.26fF
C598 a_15991_989.n3 GND 0.53fF
C599 a_15991_989.n4 GND 0.55fF
C600 a_15991_989.n5 GND 0.46fF
C601 a_15991_989.t15 GND 0.51fF
C602 a_15991_989.n6 GND 0.89fF
C603 a_15991_989.n7 GND 0.04fF
C604 a_15991_989.n8 GND 0.06fF
C605 a_15991_989.n9 GND 0.04fF
C606 a_15991_989.n10 GND 0.25fF
C607 a_15991_989.n11 GND 0.81fF
C608 a_15991_989.n12 GND 0.43fF
C609 a_15991_989.n13 GND 0.57fF
C610 a_15991_989.n14 GND 0.67fF
C611 a_15991_989.n15 GND 0.21fF
C612 a_15991_989.n16 GND 0.29fF
C613 a_15991_989.n17 GND 0.57fF
C614 VDD.n0 GND 0.12fF
C615 VDD.n1 GND 0.03fF
C616 VDD.n2 GND 0.02fF
C617 VDD.n3 GND 0.05fF
C618 VDD.n4 GND 0.01fF
C619 VDD.n5 GND 0.02fF
C620 VDD.n6 GND 0.02fF
C621 VDD.n9 GND 0.02fF
C622 VDD.n10 GND 0.02fF
C623 VDD.n11 GND 0.02fF
C624 VDD.n14 GND 0.46fF
C625 VDD.n16 GND 0.03fF
C626 VDD.n17 GND 0.02fF
C627 VDD.n18 GND 0.02fF
C628 VDD.n19 GND 0.02fF
C629 VDD.n20 GND 0.04fF
C630 VDD.n21 GND 0.28fF
C631 VDD.n22 GND 0.02fF
C632 VDD.n23 GND 0.03fF
C633 VDD.n24 GND 0.06fF
C634 VDD.n25 GND 0.15fF
C635 VDD.n26 GND 0.20fF
C636 VDD.n27 GND 0.01fF
C637 VDD.n28 GND 0.01fF
C638 VDD.n29 GND 0.07fF
C639 VDD.n30 GND 0.17fF
C640 VDD.n31 GND 0.01fF
C641 VDD.n32 GND 0.02fF
C642 VDD.n33 GND 0.02fF
C643 VDD.n34 GND 0.15fF
C644 VDD.n35 GND 0.20fF
C645 VDD.n36 GND 0.01fF
C646 VDD.n37 GND 0.06fF
C647 VDD.n38 GND 0.01fF
C648 VDD.n39 GND 0.02fF
C649 VDD.n40 GND 0.28fF
C650 VDD.n41 GND 0.01fF
C651 VDD.n42 GND 0.02fF
C652 VDD.n43 GND 0.03fF
C653 VDD.n44 GND 0.02fF
C654 VDD.n45 GND 0.02fF
C655 VDD.n46 GND 0.02fF
C656 VDD.n47 GND 0.18fF
C657 VDD.n48 GND 0.04fF
C658 VDD.n49 GND 0.04fF
C659 VDD.n50 GND 0.02fF
C660 VDD.n52 GND 0.02fF
C661 VDD.n53 GND 0.02fF
C662 VDD.n54 GND 0.02fF
C663 VDD.n55 GND 0.02fF
C664 VDD.n57 GND 0.02fF
C665 VDD.n58 GND 0.02fF
C666 VDD.n59 GND 0.02fF
C667 VDD.n61 GND 0.28fF
C668 VDD.n63 GND 0.02fF
C669 VDD.n64 GND 0.02fF
C670 VDD.n65 GND 0.03fF
C671 VDD.n66 GND 0.02fF
C672 VDD.n67 GND 0.28fF
C673 VDD.n68 GND 0.01fF
C674 VDD.n69 GND 0.02fF
C675 VDD.n70 GND 0.03fF
C676 VDD.n71 GND 0.28fF
C677 VDD.n72 GND 0.01fF
C678 VDD.n73 GND 0.02fF
C679 VDD.n74 GND 0.02fF
C680 VDD.n75 GND 0.28fF
C681 VDD.n76 GND 0.01fF
C682 VDD.n77 GND 0.02fF
C683 VDD.n78 GND 0.02fF
C684 VDD.n79 GND 0.31fF
C685 VDD.n80 GND 0.01fF
C686 VDD.n81 GND 0.03fF
C687 VDD.n82 GND 0.03fF
C688 VDD.n83 GND 0.31fF
C689 VDD.n84 GND 0.01fF
C690 VDD.n85 GND 0.03fF
C691 VDD.n86 GND 0.03fF
C692 VDD.n87 GND 0.28fF
C693 VDD.n88 GND 0.01fF
C694 VDD.n89 GND 0.02fF
C695 VDD.n90 GND 0.02fF
C696 VDD.n91 GND 0.28fF
C697 VDD.n92 GND 0.01fF
C698 VDD.n93 GND 0.02fF
C699 VDD.n94 GND 0.02fF
C700 VDD.n95 GND 0.28fF
C701 VDD.n96 GND 0.01fF
C702 VDD.n97 GND 0.02fF
C703 VDD.n98 GND 0.03fF
C704 VDD.n99 GND 0.02fF
C705 VDD.n100 GND 0.02fF
C706 VDD.n101 GND 0.02fF
C707 VDD.n102 GND 0.22fF
C708 VDD.n103 GND 0.04fF
C709 VDD.n104 GND 0.03fF
C710 VDD.n105 GND 0.02fF
C711 VDD.n106 GND 0.02fF
C712 VDD.n107 GND 0.02fF
C713 VDD.n108 GND 0.03fF
C714 VDD.n109 GND 0.02fF
C715 VDD.n111 GND 0.02fF
C716 VDD.n112 GND 0.02fF
C717 VDD.n113 GND 0.02fF
C718 VDD.n115 GND 0.28fF
C719 VDD.n117 GND 0.02fF
C720 VDD.n118 GND 0.02fF
C721 VDD.n119 GND 0.03fF
C722 VDD.n120 GND 0.02fF
C723 VDD.n121 GND 0.28fF
C724 VDD.n122 GND 0.01fF
C725 VDD.n123 GND 0.02fF
C726 VDD.n124 GND 0.03fF
C727 VDD.n125 GND 0.28fF
C728 VDD.n126 GND 0.01fF
C729 VDD.n127 GND 0.02fF
C730 VDD.n128 GND 0.02fF
C731 VDD.n129 GND 0.28fF
C732 VDD.n130 GND 0.01fF
C733 VDD.n131 GND 0.02fF
C734 VDD.n132 GND 0.02fF
C735 VDD.n133 GND 0.31fF
C736 VDD.n134 GND 0.01fF
C737 VDD.n135 GND 0.03fF
C738 VDD.n136 GND 0.03fF
C739 VDD.n137 GND 0.31fF
C740 VDD.n138 GND 0.01fF
C741 VDD.n139 GND 0.03fF
C742 VDD.n140 GND 0.03fF
C743 VDD.n141 GND 0.28fF
C744 VDD.n142 GND 0.01fF
C745 VDD.n143 GND 0.02fF
C746 VDD.n144 GND 0.02fF
C747 VDD.n145 GND 0.28fF
C748 VDD.n146 GND 0.01fF
C749 VDD.n147 GND 0.02fF
C750 VDD.n148 GND 0.02fF
C751 VDD.n149 GND 0.28fF
C752 VDD.n150 GND 0.01fF
C753 VDD.n151 GND 0.02fF
C754 VDD.n152 GND 0.03fF
C755 VDD.n153 GND 0.02fF
C756 VDD.n154 GND 0.02fF
C757 VDD.n155 GND 0.02fF
C758 VDD.n156 GND 0.22fF
C759 VDD.n157 GND 0.04fF
C760 VDD.n158 GND 0.03fF
C761 VDD.n159 GND 0.02fF
C762 VDD.n160 GND 0.02fF
C763 VDD.n161 GND 0.02fF
C764 VDD.n162 GND 0.03fF
C765 VDD.n163 GND 0.02fF
C766 VDD.n165 GND 0.02fF
C767 VDD.n166 GND 0.02fF
C768 VDD.n167 GND 0.02fF
C769 VDD.n169 GND 0.28fF
C770 VDD.n171 GND 0.02fF
C771 VDD.n172 GND 0.02fF
C772 VDD.n173 GND 0.03fF
C773 VDD.n174 GND 0.02fF
C774 VDD.n175 GND 0.28fF
C775 VDD.n176 GND 0.01fF
C776 VDD.n177 GND 0.02fF
C777 VDD.n178 GND 0.03fF
C778 VDD.n179 GND 0.06fF
C779 VDD.n180 GND 0.24fF
C780 VDD.n181 GND 0.01fF
C781 VDD.n182 GND 0.01fF
C782 VDD.n183 GND 0.02fF
C783 VDD.n184 GND 0.14fF
C784 VDD.n185 GND 0.17fF
C785 VDD.n186 GND 0.01fF
C786 VDD.n187 GND 0.02fF
C787 VDD.n188 GND 0.02fF
C788 VDD.n189 GND 0.11fF
C789 VDD.n190 GND 0.03fF
C790 VDD.n191 GND 0.31fF
C791 VDD.n192 GND 0.01fF
C792 VDD.n193 GND 0.02fF
C793 VDD.n194 GND 0.03fF
C794 VDD.n195 GND 0.17fF
C795 VDD.n196 GND 0.14fF
C796 VDD.n197 GND 0.01fF
C797 VDD.n198 GND 0.02fF
C798 VDD.n199 GND 0.03fF
C799 VDD.n200 GND 0.14fF
C800 VDD.n201 GND 0.16fF
C801 VDD.n202 GND 0.01fF
C802 VDD.n203 GND 0.02fF
C803 VDD.n204 GND 0.02fF
C804 VDD.n205 GND 0.06fF
C805 VDD.n206 GND 0.25fF
C806 VDD.n207 GND 0.01fF
C807 VDD.n208 GND 0.01fF
C808 VDD.n209 GND 0.02fF
C809 VDD.n210 GND 0.28fF
C810 VDD.n211 GND 0.01fF
C811 VDD.n212 GND 0.02fF
C812 VDD.n213 GND 0.03fF
C813 VDD.n214 GND 0.02fF
C814 VDD.n215 GND 0.02fF
C815 VDD.n216 GND 0.02fF
C816 VDD.n217 GND 0.26fF
C817 VDD.n218 GND 0.04fF
C818 VDD.n219 GND 0.03fF
C819 VDD.n220 GND 0.02fF
C820 VDD.n221 GND 0.02fF
C821 VDD.n222 GND 0.02fF
C822 VDD.n223 GND 0.03fF
C823 VDD.n224 GND 0.02fF
C824 VDD.n226 GND 0.02fF
C825 VDD.n227 GND 0.02fF
C826 VDD.n228 GND 0.02fF
C827 VDD.n230 GND 0.28fF
C828 VDD.n232 GND 0.02fF
C829 VDD.n233 GND 0.02fF
C830 VDD.n234 GND 0.03fF
C831 VDD.n235 GND 0.02fF
C832 VDD.n236 GND 0.28fF
C833 VDD.n237 GND 0.01fF
C834 VDD.n238 GND 0.02fF
C835 VDD.n239 GND 0.03fF
C836 VDD.n240 GND 0.28fF
C837 VDD.n241 GND 0.01fF
C838 VDD.n242 GND 0.02fF
C839 VDD.n243 GND 0.02fF
C840 VDD.n244 GND 0.22fF
C841 VDD.n245 GND 0.01fF
C842 VDD.n246 GND 0.07fF
C843 VDD.n247 GND 0.02fF
C844 VDD.n248 GND 0.14fF
C845 VDD.n249 GND 0.17fF
C846 VDD.n250 GND 0.01fF
C847 VDD.n251 GND 0.02fF
C848 VDD.n252 GND 0.02fF
C849 VDD.n253 GND 0.14fF
C850 VDD.n254 GND 0.16fF
C851 VDD.n255 GND 0.01fF
C852 VDD.n256 GND 0.11fF
C853 VDD.n257 GND 0.02fF
C854 VDD.n258 GND 0.02fF
C855 VDD.n259 GND 0.02fF
C856 VDD.n260 GND 0.18fF
C857 VDD.n261 GND 0.15fF
C858 VDD.n262 GND 0.01fF
C859 VDD.n263 GND 0.02fF
C860 VDD.n264 GND 0.03fF
C861 VDD.n265 GND 0.18fF
C862 VDD.n266 GND 0.15fF
C863 VDD.n267 GND 0.01fF
C864 VDD.n268 GND 0.02fF
C865 VDD.n269 GND 0.03fF
C866 VDD.n270 GND 0.11fF
C867 VDD.n271 GND 0.02fF
C868 VDD.n272 GND 0.14fF
C869 VDD.n273 GND 0.16fF
C870 VDD.n274 GND 0.01fF
C871 VDD.n275 GND 0.02fF
C872 VDD.n276 GND 0.02fF
C873 VDD.n277 GND 0.14fF
C874 VDD.n278 GND 0.17fF
C875 VDD.n279 GND 0.01fF
C876 VDD.n280 GND 0.02fF
C877 VDD.n281 GND 0.02fF
C878 VDD.n282 GND 0.06fF
C879 VDD.n283 GND 0.23fF
C880 VDD.n284 GND 0.01fF
C881 VDD.n285 GND 0.01fF
C882 VDD.n286 GND 0.02fF
C883 VDD.n287 GND 0.28fF
C884 VDD.n288 GND 0.01fF
C885 VDD.n289 GND 0.02fF
C886 VDD.n290 GND 0.02fF
C887 VDD.n291 GND 0.28fF
C888 VDD.n292 GND 0.01fF
C889 VDD.n293 GND 0.02fF
C890 VDD.n294 GND 0.03fF
C891 VDD.n295 GND 0.02fF
C892 VDD.n296 GND 0.02fF
C893 VDD.n297 GND 0.02fF
C894 VDD.n298 GND 0.31fF
C895 VDD.n299 GND 0.04fF
C896 VDD.n300 GND 0.03fF
C897 VDD.n301 GND 0.02fF
C898 VDD.n302 GND 0.02fF
C899 VDD.n303 GND 0.02fF
C900 VDD.n304 GND 0.03fF
C901 VDD.n305 GND 0.02fF
C902 VDD.n307 GND 0.02fF
C903 VDD.n308 GND 0.02fF
C904 VDD.n309 GND 0.02fF
C905 VDD.n311 GND 0.28fF
C906 VDD.n313 GND 0.02fF
C907 VDD.n314 GND 0.02fF
C908 VDD.n315 GND 0.03fF
C909 VDD.n316 GND 0.02fF
C910 VDD.n317 GND 0.28fF
C911 VDD.n318 GND 0.01fF
C912 VDD.n319 GND 0.02fF
C913 VDD.n320 GND 0.03fF
C914 VDD.n321 GND 0.28fF
C915 VDD.n322 GND 0.01fF
C916 VDD.n323 GND 0.02fF
C917 VDD.n324 GND 0.02fF
C918 VDD.n325 GND 0.22fF
C919 VDD.n326 GND 0.01fF
C920 VDD.n327 GND 0.07fF
C921 VDD.n328 GND 0.02fF
C922 VDD.n329 GND 0.14fF
C923 VDD.n330 GND 0.17fF
C924 VDD.n331 GND 0.01fF
C925 VDD.n332 GND 0.02fF
C926 VDD.n333 GND 0.02fF
C927 VDD.n334 GND 0.14fF
C928 VDD.n335 GND 0.16fF
C929 VDD.n336 GND 0.01fF
C930 VDD.n337 GND 0.11fF
C931 VDD.n338 GND 0.02fF
C932 VDD.n339 GND 0.02fF
C933 VDD.n340 GND 0.02fF
C934 VDD.n341 GND 0.18fF
C935 VDD.n342 GND 0.15fF
C936 VDD.n343 GND 0.01fF
C937 VDD.n344 GND 0.02fF
C938 VDD.n345 GND 0.03fF
C939 VDD.n346 GND 0.18fF
C940 VDD.n347 GND 0.15fF
C941 VDD.n348 GND 0.01fF
C942 VDD.n349 GND 0.02fF
C943 VDD.n350 GND 0.03fF
C944 VDD.n351 GND 0.11fF
C945 VDD.n352 GND 0.02fF
C946 VDD.n353 GND 0.14fF
C947 VDD.n354 GND 0.16fF
C948 VDD.n355 GND 0.01fF
C949 VDD.n356 GND 0.02fF
C950 VDD.n357 GND 0.02fF
C951 VDD.n358 GND 0.14fF
C952 VDD.n359 GND 0.17fF
C953 VDD.n360 GND 0.01fF
C954 VDD.n361 GND 0.02fF
C955 VDD.n362 GND 0.02fF
C956 VDD.n363 GND 0.06fF
C957 VDD.n364 GND 0.23fF
C958 VDD.n365 GND 0.01fF
C959 VDD.n366 GND 0.01fF
C960 VDD.n367 GND 0.02fF
C961 VDD.n368 GND 0.28fF
C962 VDD.n369 GND 0.01fF
C963 VDD.n370 GND 0.02fF
C964 VDD.n371 GND 0.02fF
C965 VDD.n372 GND 0.28fF
C966 VDD.n373 GND 0.01fF
C967 VDD.n374 GND 0.02fF
C968 VDD.n375 GND 0.03fF
C969 VDD.n376 GND 0.02fF
C970 VDD.n377 GND 0.02fF
C971 VDD.n378 GND 0.02fF
C972 VDD.n379 GND 0.31fF
C973 VDD.n380 GND 0.04fF
C974 VDD.n381 GND 0.03fF
C975 VDD.n382 GND 0.02fF
C976 VDD.n383 GND 0.02fF
C977 VDD.n384 GND 0.02fF
C978 VDD.n385 GND 0.03fF
C979 VDD.n386 GND 0.02fF
C980 VDD.n388 GND 0.02fF
C981 VDD.n389 GND 0.02fF
C982 VDD.n390 GND 0.02fF
C983 VDD.n392 GND 0.28fF
C984 VDD.n394 GND 0.02fF
C985 VDD.n395 GND 0.02fF
C986 VDD.n396 GND 0.03fF
C987 VDD.n397 GND 0.02fF
C988 VDD.n398 GND 0.28fF
C989 VDD.n399 GND 0.01fF
C990 VDD.n400 GND 0.02fF
C991 VDD.n401 GND 0.03fF
C992 VDD.n402 GND 0.28fF
C993 VDD.n403 GND 0.01fF
C994 VDD.n404 GND 0.02fF
C995 VDD.n405 GND 0.02fF
C996 VDD.n406 GND 0.22fF
C997 VDD.n407 GND 0.01fF
C998 VDD.n408 GND 0.07fF
C999 VDD.n409 GND 0.02fF
C1000 VDD.n410 GND 0.14fF
C1001 VDD.n411 GND 0.17fF
C1002 VDD.n412 GND 0.01fF
C1003 VDD.n413 GND 0.02fF
C1004 VDD.n414 GND 0.02fF
C1005 VDD.n415 GND 0.14fF
C1006 VDD.n416 GND 0.16fF
C1007 VDD.n417 GND 0.01fF
C1008 VDD.n418 GND 0.11fF
C1009 VDD.n419 GND 0.02fF
C1010 VDD.n420 GND 0.02fF
C1011 VDD.n421 GND 0.02fF
C1012 VDD.n422 GND 0.18fF
C1013 VDD.n423 GND 0.15fF
C1014 VDD.n424 GND 0.01fF
C1015 VDD.n425 GND 0.02fF
C1016 VDD.n426 GND 0.03fF
C1017 VDD.n427 GND 0.18fF
C1018 VDD.n428 GND 0.15fF
C1019 VDD.n429 GND 0.01fF
C1020 VDD.n430 GND 0.02fF
C1021 VDD.n431 GND 0.03fF
C1022 VDD.n432 GND 0.11fF
C1023 VDD.n433 GND 0.02fF
C1024 VDD.n434 GND 0.14fF
C1025 VDD.n435 GND 0.16fF
C1026 VDD.n436 GND 0.01fF
C1027 VDD.n437 GND 0.02fF
C1028 VDD.n438 GND 0.02fF
C1029 VDD.n439 GND 0.14fF
C1030 VDD.n440 GND 0.17fF
C1031 VDD.n441 GND 0.01fF
C1032 VDD.n442 GND 0.02fF
C1033 VDD.n443 GND 0.02fF
C1034 VDD.n444 GND 0.06fF
C1035 VDD.n445 GND 0.23fF
C1036 VDD.n446 GND 0.01fF
C1037 VDD.n447 GND 0.01fF
C1038 VDD.n448 GND 0.02fF
C1039 VDD.n449 GND 0.28fF
C1040 VDD.n450 GND 0.01fF
C1041 VDD.n451 GND 0.02fF
C1042 VDD.n452 GND 0.02fF
C1043 VDD.n453 GND 0.28fF
C1044 VDD.n454 GND 0.01fF
C1045 VDD.n455 GND 0.02fF
C1046 VDD.n456 GND 0.03fF
C1047 VDD.n457 GND 0.02fF
C1048 VDD.n458 GND 0.02fF
C1049 VDD.n459 GND 0.02fF
C1050 VDD.n460 GND 0.31fF
C1051 VDD.n461 GND 0.04fF
C1052 VDD.n462 GND 0.03fF
C1053 VDD.n463 GND 0.02fF
C1054 VDD.n464 GND 0.02fF
C1055 VDD.n465 GND 0.02fF
C1056 VDD.n466 GND 0.03fF
C1057 VDD.n467 GND 0.02fF
C1058 VDD.n469 GND 0.02fF
C1059 VDD.n470 GND 0.02fF
C1060 VDD.n471 GND 0.02fF
C1061 VDD.n473 GND 0.28fF
C1062 VDD.n475 GND 0.02fF
C1063 VDD.n476 GND 0.02fF
C1064 VDD.n477 GND 0.03fF
C1065 VDD.n478 GND 0.02fF
C1066 VDD.n479 GND 0.28fF
C1067 VDD.n480 GND 0.01fF
C1068 VDD.n481 GND 0.02fF
C1069 VDD.n482 GND 0.03fF
C1070 VDD.n483 GND 0.28fF
C1071 VDD.n484 GND 0.01fF
C1072 VDD.n485 GND 0.02fF
C1073 VDD.n486 GND 0.02fF
C1074 VDD.n487 GND 0.22fF
C1075 VDD.n488 GND 0.01fF
C1076 VDD.n489 GND 0.07fF
C1077 VDD.n490 GND 0.02fF
C1078 VDD.n491 GND 0.14fF
C1079 VDD.n492 GND 0.17fF
C1080 VDD.n493 GND 0.01fF
C1081 VDD.n494 GND 0.02fF
C1082 VDD.n495 GND 0.02fF
C1083 VDD.n496 GND 0.14fF
C1084 VDD.n497 GND 0.16fF
C1085 VDD.n498 GND 0.01fF
C1086 VDD.n499 GND 0.11fF
C1087 VDD.n500 GND 0.02fF
C1088 VDD.n501 GND 0.02fF
C1089 VDD.n502 GND 0.02fF
C1090 VDD.n503 GND 0.18fF
C1091 VDD.n504 GND 0.15fF
C1092 VDD.n505 GND 0.01fF
C1093 VDD.n506 GND 0.02fF
C1094 VDD.n507 GND 0.03fF
C1095 VDD.n508 GND 0.18fF
C1096 VDD.n509 GND 0.15fF
C1097 VDD.n510 GND 0.01fF
C1098 VDD.n511 GND 0.02fF
C1099 VDD.n512 GND 0.03fF
C1100 VDD.n513 GND 0.11fF
C1101 VDD.n514 GND 0.02fF
C1102 VDD.n515 GND 0.14fF
C1103 VDD.n516 GND 0.16fF
C1104 VDD.n517 GND 0.01fF
C1105 VDD.n518 GND 0.02fF
C1106 VDD.n519 GND 0.02fF
C1107 VDD.n520 GND 0.14fF
C1108 VDD.n521 GND 0.17fF
C1109 VDD.n522 GND 0.01fF
C1110 VDD.n523 GND 0.02fF
C1111 VDD.n524 GND 0.02fF
C1112 VDD.n525 GND 0.06fF
C1113 VDD.n526 GND 0.23fF
C1114 VDD.n527 GND 0.01fF
C1115 VDD.n528 GND 0.01fF
C1116 VDD.n529 GND 0.02fF
C1117 VDD.n530 GND 0.28fF
C1118 VDD.n531 GND 0.01fF
C1119 VDD.n532 GND 0.02fF
C1120 VDD.n533 GND 0.02fF
C1121 VDD.n534 GND 0.28fF
C1122 VDD.n535 GND 0.01fF
C1123 VDD.n536 GND 0.02fF
C1124 VDD.n537 GND 0.03fF
C1125 VDD.n538 GND 0.02fF
C1126 VDD.n539 GND 0.02fF
C1127 VDD.n540 GND 0.02fF
C1128 VDD.n541 GND 0.31fF
C1129 VDD.n542 GND 0.04fF
C1130 VDD.n543 GND 0.03fF
C1131 VDD.n544 GND 0.02fF
C1132 VDD.n545 GND 0.02fF
C1133 VDD.n546 GND 0.02fF
C1134 VDD.n547 GND 0.03fF
C1135 VDD.n548 GND 0.02fF
C1136 VDD.n550 GND 0.02fF
C1137 VDD.n551 GND 0.02fF
C1138 VDD.n552 GND 0.02fF
C1139 VDD.n554 GND 0.28fF
C1140 VDD.n556 GND 0.02fF
C1141 VDD.n557 GND 0.02fF
C1142 VDD.n558 GND 0.03fF
C1143 VDD.n559 GND 0.02fF
C1144 VDD.n560 GND 0.28fF
C1145 VDD.n561 GND 0.01fF
C1146 VDD.n562 GND 0.02fF
C1147 VDD.n563 GND 0.03fF
C1148 VDD.n564 GND 0.28fF
C1149 VDD.n565 GND 0.01fF
C1150 VDD.n566 GND 0.02fF
C1151 VDD.n567 GND 0.02fF
C1152 VDD.n568 GND 0.22fF
C1153 VDD.n569 GND 0.01fF
C1154 VDD.n570 GND 0.07fF
C1155 VDD.n571 GND 0.02fF
C1156 VDD.n572 GND 0.14fF
C1157 VDD.n573 GND 0.17fF
C1158 VDD.n574 GND 0.01fF
C1159 VDD.n575 GND 0.02fF
C1160 VDD.n576 GND 0.02fF
C1161 VDD.n577 GND 0.14fF
C1162 VDD.n578 GND 0.16fF
C1163 VDD.n579 GND 0.01fF
C1164 VDD.n580 GND 0.11fF
C1165 VDD.n581 GND 0.02fF
C1166 VDD.n582 GND 0.02fF
C1167 VDD.n583 GND 0.02fF
C1168 VDD.n584 GND 0.18fF
C1169 VDD.n585 GND 0.15fF
C1170 VDD.n586 GND 0.01fF
C1171 VDD.n587 GND 0.02fF
C1172 VDD.n588 GND 0.03fF
C1173 VDD.n589 GND 0.18fF
C1174 VDD.n590 GND 0.15fF
C1175 VDD.n591 GND 0.01fF
C1176 VDD.n592 GND 0.02fF
C1177 VDD.n593 GND 0.03fF
C1178 VDD.n594 GND 0.11fF
C1179 VDD.n595 GND 0.02fF
C1180 VDD.n596 GND 0.14fF
C1181 VDD.n597 GND 0.16fF
C1182 VDD.n598 GND 0.01fF
C1183 VDD.n599 GND 0.02fF
C1184 VDD.n600 GND 0.02fF
C1185 VDD.n601 GND 0.14fF
C1186 VDD.n602 GND 0.17fF
C1187 VDD.n603 GND 0.01fF
C1188 VDD.n604 GND 0.02fF
C1189 VDD.n605 GND 0.02fF
C1190 VDD.n606 GND 0.06fF
C1191 VDD.n607 GND 0.23fF
C1192 VDD.n608 GND 0.01fF
C1193 VDD.n609 GND 0.01fF
C1194 VDD.n610 GND 0.02fF
C1195 VDD.n611 GND 0.28fF
C1196 VDD.n612 GND 0.01fF
C1197 VDD.n613 GND 0.02fF
C1198 VDD.n614 GND 0.02fF
C1199 VDD.n615 GND 0.28fF
C1200 VDD.n616 GND 0.01fF
C1201 VDD.n617 GND 0.02fF
C1202 VDD.n618 GND 0.03fF
C1203 VDD.n619 GND 0.02fF
C1204 VDD.n620 GND 0.02fF
C1205 VDD.n621 GND 0.02fF
C1206 VDD.n622 GND 0.31fF
C1207 VDD.n623 GND 0.04fF
C1208 VDD.n624 GND 0.03fF
C1209 VDD.n625 GND 0.02fF
C1210 VDD.n626 GND 0.02fF
C1211 VDD.n627 GND 0.02fF
C1212 VDD.n628 GND 0.03fF
C1213 VDD.n629 GND 0.02fF
C1214 VDD.n631 GND 0.02fF
C1215 VDD.n632 GND 0.02fF
C1216 VDD.n633 GND 0.02fF
C1217 VDD.n635 GND 0.28fF
C1218 VDD.n637 GND 0.02fF
C1219 VDD.n638 GND 0.02fF
C1220 VDD.n639 GND 0.03fF
C1221 VDD.n640 GND 0.02fF
C1222 VDD.n641 GND 0.28fF
C1223 VDD.n642 GND 0.01fF
C1224 VDD.n643 GND 0.02fF
C1225 VDD.n644 GND 0.03fF
C1226 VDD.n645 GND 0.28fF
C1227 VDD.n646 GND 0.01fF
C1228 VDD.n647 GND 0.02fF
C1229 VDD.n648 GND 0.02fF
C1230 VDD.n649 GND 0.22fF
C1231 VDD.n650 GND 0.01fF
C1232 VDD.n651 GND 0.07fF
C1233 VDD.n652 GND 0.02fF
C1234 VDD.n653 GND 0.14fF
C1235 VDD.n654 GND 0.17fF
C1236 VDD.n655 GND 0.01fF
C1237 VDD.n656 GND 0.02fF
C1238 VDD.n657 GND 0.02fF
C1239 VDD.n658 GND 0.14fF
C1240 VDD.n659 GND 0.16fF
C1241 VDD.n660 GND 0.01fF
C1242 VDD.n661 GND 0.11fF
C1243 VDD.n662 GND 0.02fF
C1244 VDD.n663 GND 0.02fF
C1245 VDD.n664 GND 0.02fF
C1246 VDD.n665 GND 0.18fF
C1247 VDD.n666 GND 0.15fF
C1248 VDD.n667 GND 0.01fF
C1249 VDD.n668 GND 0.02fF
C1250 VDD.n669 GND 0.03fF
C1251 VDD.n670 GND 0.18fF
C1252 VDD.n671 GND 0.15fF
C1253 VDD.n672 GND 0.01fF
C1254 VDD.n673 GND 0.02fF
C1255 VDD.n674 GND 0.03fF
C1256 VDD.n675 GND 0.11fF
C1257 VDD.n676 GND 0.02fF
C1258 VDD.n677 GND 0.14fF
C1259 VDD.n678 GND 0.16fF
C1260 VDD.n679 GND 0.01fF
C1261 VDD.n680 GND 0.02fF
C1262 VDD.n681 GND 0.02fF
C1263 VDD.n682 GND 0.14fF
C1264 VDD.n683 GND 0.17fF
C1265 VDD.n684 GND 0.01fF
C1266 VDD.n685 GND 0.02fF
C1267 VDD.n686 GND 0.02fF
C1268 VDD.n687 GND 0.06fF
C1269 VDD.n688 GND 0.23fF
C1270 VDD.n689 GND 0.01fF
C1271 VDD.n690 GND 0.01fF
C1272 VDD.n691 GND 0.02fF
C1273 VDD.n692 GND 0.28fF
C1274 VDD.n693 GND 0.01fF
C1275 VDD.n694 GND 0.02fF
C1276 VDD.n695 GND 0.02fF
C1277 VDD.n696 GND 0.28fF
C1278 VDD.n697 GND 0.01fF
C1279 VDD.n698 GND 0.02fF
C1280 VDD.n699 GND 0.03fF
C1281 VDD.n700 GND 0.02fF
C1282 VDD.n701 GND 0.02fF
C1283 VDD.n702 GND 0.02fF
C1284 VDD.n703 GND 0.31fF
C1285 VDD.n704 GND 0.04fF
C1286 VDD.n705 GND 0.03fF
C1287 VDD.n706 GND 0.02fF
C1288 VDD.n707 GND 0.02fF
C1289 VDD.n708 GND 0.02fF
C1290 VDD.n709 GND 0.03fF
C1291 VDD.n710 GND 0.02fF
C1292 VDD.n712 GND 0.02fF
C1293 VDD.n713 GND 0.02fF
C1294 VDD.n714 GND 0.02fF
C1295 VDD.n716 GND 0.28fF
C1296 VDD.n718 GND 0.02fF
C1297 VDD.n719 GND 0.02fF
C1298 VDD.n720 GND 0.03fF
C1299 VDD.n721 GND 0.02fF
C1300 VDD.n722 GND 0.28fF
C1301 VDD.n723 GND 0.01fF
C1302 VDD.n724 GND 0.02fF
C1303 VDD.n725 GND 0.03fF
C1304 VDD.n726 GND 0.28fF
C1305 VDD.n727 GND 0.01fF
C1306 VDD.n728 GND 0.02fF
C1307 VDD.n729 GND 0.02fF
C1308 VDD.n730 GND 0.22fF
C1309 VDD.n731 GND 0.01fF
C1310 VDD.n732 GND 0.07fF
C1311 VDD.n733 GND 0.02fF
C1312 VDD.n734 GND 0.14fF
C1313 VDD.n735 GND 0.17fF
C1314 VDD.n736 GND 0.01fF
C1315 VDD.n737 GND 0.02fF
C1316 VDD.n738 GND 0.02fF
C1317 VDD.n739 GND 0.14fF
C1318 VDD.n740 GND 0.16fF
C1319 VDD.n741 GND 0.01fF
C1320 VDD.n742 GND 0.11fF
C1321 VDD.n743 GND 0.02fF
C1322 VDD.n744 GND 0.02fF
C1323 VDD.n745 GND 0.02fF
C1324 VDD.n746 GND 0.18fF
C1325 VDD.n747 GND 0.15fF
C1326 VDD.n748 GND 0.01fF
C1327 VDD.n749 GND 0.02fF
C1328 VDD.n750 GND 0.03fF
C1329 VDD.n751 GND 0.18fF
C1330 VDD.n752 GND 0.15fF
C1331 VDD.n753 GND 0.01fF
C1332 VDD.n754 GND 0.02fF
C1333 VDD.n755 GND 0.03fF
C1334 VDD.n756 GND 0.11fF
C1335 VDD.n757 GND 0.02fF
C1336 VDD.n758 GND 0.14fF
C1337 VDD.n759 GND 0.16fF
C1338 VDD.n760 GND 0.01fF
C1339 VDD.n761 GND 0.02fF
C1340 VDD.n762 GND 0.02fF
C1341 VDD.n763 GND 0.14fF
C1342 VDD.n764 GND 0.17fF
C1343 VDD.n765 GND 0.01fF
C1344 VDD.n766 GND 0.02fF
C1345 VDD.n767 GND 0.02fF
C1346 VDD.n768 GND 0.06fF
C1347 VDD.n769 GND 0.23fF
C1348 VDD.n770 GND 0.01fF
C1349 VDD.n771 GND 0.01fF
C1350 VDD.n772 GND 0.02fF
C1351 VDD.n773 GND 0.28fF
C1352 VDD.n774 GND 0.01fF
C1353 VDD.n775 GND 0.02fF
C1354 VDD.n776 GND 0.02fF
C1355 VDD.n777 GND 0.28fF
C1356 VDD.n778 GND 0.01fF
C1357 VDD.n779 GND 0.02fF
C1358 VDD.n780 GND 0.03fF
C1359 VDD.n781 GND 0.02fF
C1360 VDD.n782 GND 0.02fF
C1361 VDD.n783 GND 0.02fF
C1362 VDD.n784 GND 0.31fF
C1363 VDD.n785 GND 0.04fF
C1364 VDD.n786 GND 0.03fF
C1365 VDD.n787 GND 0.02fF
C1366 VDD.n788 GND 0.02fF
C1367 VDD.n789 GND 0.02fF
C1368 VDD.n790 GND 0.03fF
C1369 VDD.n791 GND 0.02fF
C1370 VDD.n793 GND 0.02fF
C1371 VDD.n794 GND 0.02fF
C1372 VDD.n795 GND 0.02fF
C1373 VDD.n797 GND 0.28fF
C1374 VDD.n799 GND 0.02fF
C1375 VDD.n800 GND 0.02fF
C1376 VDD.n801 GND 0.03fF
C1377 VDD.n802 GND 0.02fF
C1378 VDD.n803 GND 0.28fF
C1379 VDD.n804 GND 0.01fF
C1380 VDD.n805 GND 0.02fF
C1381 VDD.n806 GND 0.03fF
C1382 VDD.n807 GND 0.28fF
C1383 VDD.n808 GND 0.01fF
C1384 VDD.n809 GND 0.02fF
C1385 VDD.n810 GND 0.02fF
C1386 VDD.n811 GND 0.22fF
C1387 VDD.n812 GND 0.01fF
C1388 VDD.n813 GND 0.07fF
C1389 VDD.n814 GND 0.02fF
C1390 VDD.n815 GND 0.14fF
C1391 VDD.n816 GND 0.17fF
C1392 VDD.n817 GND 0.01fF
C1393 VDD.n818 GND 0.02fF
C1394 VDD.n819 GND 0.02fF
C1395 VDD.n820 GND 0.14fF
C1396 VDD.n821 GND 0.16fF
C1397 VDD.n822 GND 0.01fF
C1398 VDD.n823 GND 0.11fF
C1399 VDD.n824 GND 0.02fF
C1400 VDD.n825 GND 0.02fF
C1401 VDD.n826 GND 0.02fF
C1402 VDD.n827 GND 0.18fF
C1403 VDD.n828 GND 0.15fF
C1404 VDD.n829 GND 0.01fF
C1405 VDD.n830 GND 0.02fF
C1406 VDD.n831 GND 0.03fF
C1407 VDD.n832 GND 0.18fF
C1408 VDD.n833 GND 0.15fF
C1409 VDD.n834 GND 0.01fF
C1410 VDD.n835 GND 0.02fF
C1411 VDD.n836 GND 0.03fF
C1412 VDD.n837 GND 0.11fF
C1413 VDD.n838 GND 0.02fF
C1414 VDD.n839 GND 0.14fF
C1415 VDD.n840 GND 0.16fF
C1416 VDD.n841 GND 0.01fF
C1417 VDD.n842 GND 0.02fF
C1418 VDD.n843 GND 0.02fF
C1419 VDD.n844 GND 0.14fF
C1420 VDD.n845 GND 0.17fF
C1421 VDD.n846 GND 0.01fF
C1422 VDD.n847 GND 0.02fF
C1423 VDD.n848 GND 0.02fF
C1424 VDD.n849 GND 0.02fF
C1425 VDD.n850 GND 0.02fF
C1426 VDD.n851 GND 0.02fF
C1427 VDD.n852 GND 0.20fF
C1428 VDD.n853 GND 0.03fF
C1429 VDD.n854 GND 0.02fF
C1430 VDD.n855 GND 0.02fF
C1431 VDD.n856 GND 0.02fF
C1432 VDD.n857 GND 0.03fF
C1433 VDD.n858 GND 0.02fF
C1434 VDD.n860 GND 0.02fF
C1435 VDD.n861 GND 0.02fF
C1436 VDD.n862 GND 0.02fF
C1437 VDD.n864 GND 0.46fF
C1438 VDD.n866 GND 0.03fF
C1439 VDD.n867 GND 0.04fF
C1440 VDD.n868 GND 0.28fF
C1441 VDD.n869 GND 0.02fF
C1442 VDD.n870 GND 0.03fF
C1443 VDD.n871 GND 0.03fF
C1444 VDD.n872 GND 0.28fF
C1445 VDD.n873 GND 0.01fF
C1446 VDD.n874 GND 0.02fF
C1447 VDD.n875 GND 0.02fF
C1448 VDD.n876 GND 0.06fF
C1449 VDD.n877 GND 0.23fF
C1450 VDD.n878 GND 0.01fF
C1451 VDD.n879 GND 0.01fF
C1452 VDD.n880 GND 0.02fF
C1453 VDD.n881 GND 0.14fF
C1454 VDD.n882 GND 0.17fF
C1455 VDD.n883 GND 0.01fF
C1456 VDD.n884 GND 0.02fF
C1457 VDD.n885 GND 0.02fF
C1458 VDD.n886 GND 0.11fF
C1459 VDD.n887 GND 0.02fF
C1460 VDD.n888 GND 0.14fF
C1461 VDD.n889 GND 0.16fF
C1462 VDD.n890 GND 0.01fF
C1463 VDD.n891 GND 0.02fF
C1464 VDD.n892 GND 0.02fF
C1465 VDD.n893 GND 0.18fF
C1466 VDD.n894 GND 0.15fF
C1467 VDD.n895 GND 0.01fF
C1468 VDD.n896 GND 0.02fF
C1469 VDD.n897 GND 0.03fF
C1470 VDD.n898 GND 0.18fF
C1471 VDD.n899 GND 0.15fF
C1472 VDD.n900 GND 0.01fF
C1473 VDD.n901 GND 0.02fF
C1474 VDD.n902 GND 0.03fF
C1475 VDD.n903 GND 0.14fF
C1476 VDD.n904 GND 0.16fF
C1477 VDD.n905 GND 0.01fF
C1478 VDD.n906 GND 0.11fF
C1479 VDD.n907 GND 0.02fF
C1480 VDD.n908 GND 0.02fF
C1481 VDD.n909 GND 0.02fF
C1482 VDD.n910 GND 0.14fF
C1483 VDD.n911 GND 0.17fF
C1484 VDD.n912 GND 0.01fF
C1485 VDD.n913 GND 0.02fF
C1486 VDD.n914 GND 0.02fF
C1487 VDD.n915 GND 0.22fF
C1488 VDD.n916 GND 0.01fF
C1489 VDD.n917 GND 0.07fF
C1490 VDD.n918 GND 0.02fF
C1491 VDD.n919 GND 0.28fF
C1492 VDD.n920 GND 0.01fF
C1493 VDD.n921 GND 0.02fF
C1494 VDD.n922 GND 0.02fF
C1495 VDD.n923 GND 0.28fF
C1496 VDD.n924 GND 0.01fF
C1497 VDD.n925 GND 0.02fF
C1498 VDD.n926 GND 0.03fF
C1499 VDD.n927 GND 0.02fF
C1500 VDD.n928 GND 0.02fF
C1501 VDD.n929 GND 0.02fF
C1502 VDD.n930 GND 0.02fF
C1503 VDD.n931 GND 0.02fF
C1504 VDD.n932 GND 0.02fF
C1505 VDD.n934 GND 0.02fF
C1506 VDD.n935 GND 0.02fF
C1507 VDD.n936 GND 0.02fF
C1508 VDD.n937 GND 0.02fF
C1509 VDD.n939 GND 0.04fF
C1510 VDD.n940 GND 0.02fF
C1511 VDD.n941 GND 0.31fF
C1512 VDD.n942 GND 0.04fF
C1513 VDD.n944 GND 0.28fF
C1514 VDD.n946 GND 0.02fF
C1515 VDD.n947 GND 0.02fF
C1516 VDD.n948 GND 0.03fF
C1517 VDD.n949 GND 0.02fF
C1518 VDD.n950 GND 0.28fF
C1519 VDD.n951 GND 0.01fF
C1520 VDD.n952 GND 0.02fF
C1521 VDD.n953 GND 0.03fF
C1522 VDD.n954 GND 0.28fF
C1523 VDD.n955 GND 0.01fF
C1524 VDD.n956 GND 0.02fF
C1525 VDD.n957 GND 0.02fF
C1526 VDD.n958 GND 0.06fF
C1527 VDD.n959 GND 0.23fF
C1528 VDD.n960 GND 0.01fF
C1529 VDD.n961 GND 0.01fF
C1530 VDD.n962 GND 0.02fF
C1531 VDD.n963 GND 0.14fF
C1532 VDD.n964 GND 0.17fF
C1533 VDD.n965 GND 0.01fF
C1534 VDD.n966 GND 0.02fF
C1535 VDD.n967 GND 0.02fF
C1536 VDD.n968 GND 0.11fF
C1537 VDD.n969 GND 0.02fF
C1538 VDD.n970 GND 0.14fF
C1539 VDD.n971 GND 0.16fF
C1540 VDD.n972 GND 0.01fF
C1541 VDD.n973 GND 0.02fF
C1542 VDD.n974 GND 0.02fF
C1543 VDD.n975 GND 0.18fF
C1544 VDD.n976 GND 0.15fF
C1545 VDD.n977 GND 0.01fF
C1546 VDD.n978 GND 0.02fF
C1547 VDD.n979 GND 0.03fF
C1548 VDD.n980 GND 0.18fF
C1549 VDD.n981 GND 0.15fF
C1550 VDD.n982 GND 0.01fF
C1551 VDD.n983 GND 0.02fF
C1552 VDD.n984 GND 0.03fF
C1553 VDD.n985 GND 0.14fF
C1554 VDD.n986 GND 0.16fF
C1555 VDD.n987 GND 0.01fF
C1556 VDD.n988 GND 0.11fF
C1557 VDD.n989 GND 0.02fF
C1558 VDD.n990 GND 0.02fF
C1559 VDD.n991 GND 0.02fF
C1560 VDD.n992 GND 0.14fF
C1561 VDD.n993 GND 0.17fF
C1562 VDD.n994 GND 0.01fF
C1563 VDD.n995 GND 0.02fF
C1564 VDD.n996 GND 0.02fF
C1565 VDD.n997 GND 0.22fF
C1566 VDD.n998 GND 0.01fF
C1567 VDD.n999 GND 0.07fF
C1568 VDD.n1000 GND 0.02fF
C1569 VDD.n1001 GND 0.28fF
C1570 VDD.n1002 GND 0.01fF
C1571 VDD.n1003 GND 0.02fF
C1572 VDD.n1004 GND 0.02fF
C1573 VDD.n1005 GND 0.28fF
C1574 VDD.n1006 GND 0.01fF
C1575 VDD.n1007 GND 0.02fF
C1576 VDD.n1008 GND 0.03fF
C1577 VDD.n1009 GND 0.02fF
C1578 VDD.n1010 GND 0.02fF
C1579 VDD.n1011 GND 0.02fF
C1580 VDD.n1012 GND 0.31fF
C1581 VDD.n1013 GND 0.04fF
C1582 VDD.n1014 GND 0.03fF
C1583 VDD.n1015 GND 0.02fF
C1584 VDD.n1016 GND 0.02fF
C1585 VDD.n1017 GND 0.02fF
C1586 VDD.n1018 GND 0.03fF
C1587 VDD.n1019 GND 0.02fF
C1588 VDD.n1021 GND 0.02fF
C1589 VDD.n1022 GND 0.02fF
C1590 VDD.n1023 GND 0.02fF
C1591 VDD.n1025 GND 0.28fF
C1592 VDD.n1027 GND 0.02fF
C1593 VDD.n1028 GND 0.02fF
C1594 VDD.n1029 GND 0.03fF
C1595 VDD.n1030 GND 0.02fF
C1596 VDD.n1031 GND 0.28fF
C1597 VDD.n1032 GND 0.01fF
C1598 VDD.n1033 GND 0.02fF
C1599 VDD.n1034 GND 0.03fF
C1600 VDD.n1035 GND 0.28fF
C1601 VDD.n1036 GND 0.01fF
C1602 VDD.n1037 GND 0.02fF
C1603 VDD.n1038 GND 0.02fF
C1604 VDD.n1039 GND 0.06fF
C1605 VDD.n1040 GND 0.23fF
C1606 VDD.n1041 GND 0.01fF
C1607 VDD.n1042 GND 0.01fF
C1608 VDD.n1043 GND 0.02fF
C1609 VDD.n1044 GND 0.14fF
C1610 VDD.n1045 GND 0.17fF
C1611 VDD.n1046 GND 0.01fF
C1612 VDD.n1047 GND 0.02fF
C1613 VDD.n1048 GND 0.02fF
C1614 VDD.n1049 GND 0.11fF
C1615 VDD.n1050 GND 0.02fF
C1616 VDD.n1051 GND 0.14fF
C1617 VDD.n1052 GND 0.16fF
C1618 VDD.n1053 GND 0.01fF
C1619 VDD.n1054 GND 0.02fF
C1620 VDD.n1055 GND 0.02fF
C1621 VDD.n1056 GND 0.18fF
C1622 VDD.n1057 GND 0.15fF
C1623 VDD.n1058 GND 0.01fF
C1624 VDD.n1059 GND 0.02fF
C1625 VDD.n1060 GND 0.03fF
C1626 VDD.n1061 GND 0.18fF
C1627 VDD.n1062 GND 0.15fF
C1628 VDD.n1063 GND 0.01fF
C1629 VDD.n1064 GND 0.02fF
C1630 VDD.n1065 GND 0.03fF
C1631 VDD.n1066 GND 0.14fF
C1632 VDD.n1067 GND 0.16fF
C1633 VDD.n1068 GND 0.01fF
C1634 VDD.n1069 GND 0.11fF
C1635 VDD.n1070 GND 0.02fF
C1636 VDD.n1071 GND 0.02fF
C1637 VDD.n1072 GND 0.02fF
C1638 VDD.n1073 GND 0.14fF
C1639 VDD.n1074 GND 0.17fF
C1640 VDD.n1075 GND 0.01fF
C1641 VDD.n1076 GND 0.02fF
C1642 VDD.n1077 GND 0.02fF
C1643 VDD.n1078 GND 0.22fF
C1644 VDD.n1079 GND 0.01fF
C1645 VDD.n1080 GND 0.07fF
C1646 VDD.n1081 GND 0.02fF
C1647 VDD.n1082 GND 0.28fF
C1648 VDD.n1083 GND 0.01fF
C1649 VDD.n1084 GND 0.02fF
C1650 VDD.n1085 GND 0.02fF
C1651 VDD.n1086 GND 0.28fF
C1652 VDD.n1087 GND 0.01fF
C1653 VDD.n1088 GND 0.02fF
C1654 VDD.n1089 GND 0.03fF
C1655 VDD.n1090 GND 0.02fF
C1656 VDD.n1091 GND 0.02fF
C1657 VDD.n1092 GND 0.02fF
C1658 VDD.n1093 GND 0.31fF
C1659 VDD.n1094 GND 0.04fF
C1660 VDD.n1095 GND 0.03fF
C1661 VDD.n1096 GND 0.02fF
C1662 VDD.n1097 GND 0.02fF
C1663 VDD.n1098 GND 0.02fF
C1664 VDD.n1099 GND 0.03fF
C1665 VDD.n1100 GND 0.02fF
C1666 VDD.n1102 GND 0.02fF
C1667 VDD.n1103 GND 0.02fF
C1668 VDD.n1104 GND 0.02fF
C1669 VDD.n1106 GND 0.28fF
C1670 VDD.n1108 GND 0.02fF
C1671 VDD.n1109 GND 0.02fF
C1672 VDD.n1110 GND 0.03fF
C1673 VDD.n1111 GND 0.02fF
C1674 VDD.n1112 GND 0.28fF
C1675 VDD.n1113 GND 0.01fF
C1676 VDD.n1114 GND 0.02fF
C1677 VDD.n1115 GND 0.03fF
C1678 VDD.n1116 GND 0.28fF
C1679 VDD.n1117 GND 0.01fF
C1680 VDD.n1118 GND 0.02fF
C1681 VDD.n1119 GND 0.02fF
C1682 VDD.n1120 GND 0.06fF
C1683 VDD.n1121 GND 0.23fF
C1684 VDD.n1122 GND 0.01fF
C1685 VDD.n1123 GND 0.01fF
C1686 VDD.n1124 GND 0.02fF
C1687 VDD.n1125 GND 0.14fF
C1688 VDD.n1126 GND 0.17fF
C1689 VDD.n1127 GND 0.01fF
C1690 VDD.n1128 GND 0.02fF
C1691 VDD.n1129 GND 0.02fF
C1692 VDD.n1130 GND 0.11fF
C1693 VDD.n1131 GND 0.02fF
C1694 VDD.n1132 GND 0.14fF
C1695 VDD.n1133 GND 0.16fF
C1696 VDD.n1134 GND 0.01fF
C1697 VDD.n1135 GND 0.02fF
C1698 VDD.n1136 GND 0.02fF
C1699 VDD.n1137 GND 0.18fF
C1700 VDD.n1138 GND 0.15fF
C1701 VDD.n1139 GND 0.01fF
C1702 VDD.n1140 GND 0.02fF
C1703 VDD.n1141 GND 0.03fF
C1704 VDD.n1142 GND 0.18fF
C1705 VDD.n1143 GND 0.15fF
C1706 VDD.n1144 GND 0.01fF
C1707 VDD.n1145 GND 0.02fF
C1708 VDD.n1146 GND 0.03fF
C1709 VDD.n1147 GND 0.14fF
C1710 VDD.n1148 GND 0.16fF
C1711 VDD.n1149 GND 0.01fF
C1712 VDD.n1150 GND 0.11fF
C1713 VDD.n1151 GND 0.02fF
C1714 VDD.n1152 GND 0.02fF
C1715 VDD.n1153 GND 0.02fF
C1716 VDD.n1154 GND 0.14fF
C1717 VDD.n1155 GND 0.17fF
C1718 VDD.n1156 GND 0.01fF
C1719 VDD.n1157 GND 0.02fF
C1720 VDD.n1158 GND 0.02fF
C1721 VDD.n1159 GND 0.22fF
C1722 VDD.n1160 GND 0.01fF
C1723 VDD.n1161 GND 0.07fF
C1724 VDD.n1162 GND 0.02fF
C1725 VDD.n1163 GND 0.28fF
C1726 VDD.n1164 GND 0.01fF
C1727 VDD.n1165 GND 0.02fF
C1728 VDD.n1166 GND 0.02fF
C1729 VDD.n1167 GND 0.28fF
C1730 VDD.n1168 GND 0.01fF
C1731 VDD.n1169 GND 0.02fF
C1732 VDD.n1170 GND 0.03fF
C1733 VDD.n1171 GND 0.02fF
C1734 VDD.n1172 GND 0.02fF
C1735 VDD.n1173 GND 0.02fF
C1736 VDD.n1174 GND 0.31fF
C1737 VDD.n1175 GND 0.04fF
C1738 VDD.n1176 GND 0.03fF
C1739 VDD.n1177 GND 0.02fF
C1740 VDD.n1178 GND 0.02fF
C1741 VDD.n1179 GND 0.02fF
C1742 VDD.n1180 GND 0.03fF
C1743 VDD.n1181 GND 0.02fF
C1744 VDD.n1183 GND 0.02fF
C1745 VDD.n1184 GND 0.02fF
C1746 VDD.n1185 GND 0.02fF
C1747 VDD.n1187 GND 0.28fF
C1748 VDD.n1189 GND 0.02fF
C1749 VDD.n1190 GND 0.02fF
C1750 VDD.n1191 GND 0.03fF
C1751 VDD.n1192 GND 0.02fF
C1752 VDD.n1193 GND 0.28fF
C1753 VDD.n1194 GND 0.01fF
C1754 VDD.n1195 GND 0.02fF
C1755 VDD.n1196 GND 0.03fF
C1756 VDD.n1197 GND 0.28fF
C1757 VDD.n1198 GND 0.01fF
C1758 VDD.n1199 GND 0.02fF
C1759 VDD.n1200 GND 0.02fF
C1760 VDD.n1201 GND 0.06fF
C1761 VDD.n1202 GND 0.23fF
C1762 VDD.n1203 GND 0.01fF
C1763 VDD.n1204 GND 0.01fF
C1764 VDD.n1205 GND 0.02fF
C1765 VDD.n1206 GND 0.14fF
C1766 VDD.n1207 GND 0.17fF
C1767 VDD.n1208 GND 0.01fF
C1768 VDD.n1209 GND 0.02fF
C1769 VDD.n1210 GND 0.02fF
C1770 VDD.n1211 GND 0.11fF
C1771 VDD.n1212 GND 0.02fF
C1772 VDD.n1213 GND 0.14fF
C1773 VDD.n1214 GND 0.16fF
C1774 VDD.n1215 GND 0.01fF
C1775 VDD.n1216 GND 0.02fF
C1776 VDD.n1217 GND 0.02fF
C1777 VDD.n1218 GND 0.18fF
C1778 VDD.n1219 GND 0.15fF
C1779 VDD.n1220 GND 0.01fF
C1780 VDD.n1221 GND 0.02fF
C1781 VDD.n1222 GND 0.03fF
C1782 VDD.n1223 GND 0.18fF
C1783 VDD.n1224 GND 0.15fF
C1784 VDD.n1225 GND 0.01fF
C1785 VDD.n1226 GND 0.02fF
C1786 VDD.n1227 GND 0.03fF
C1787 VDD.n1228 GND 0.14fF
C1788 VDD.n1229 GND 0.16fF
C1789 VDD.n1230 GND 0.01fF
C1790 VDD.n1231 GND 0.11fF
C1791 VDD.n1232 GND 0.02fF
C1792 VDD.n1233 GND 0.02fF
C1793 VDD.n1234 GND 0.02fF
C1794 VDD.n1235 GND 0.14fF
C1795 VDD.n1236 GND 0.17fF
C1796 VDD.n1237 GND 0.01fF
C1797 VDD.n1238 GND 0.02fF
C1798 VDD.n1239 GND 0.02fF
C1799 VDD.n1240 GND 0.22fF
C1800 VDD.n1241 GND 0.01fF
C1801 VDD.n1242 GND 0.07fF
C1802 VDD.n1243 GND 0.02fF
C1803 VDD.n1244 GND 0.28fF
C1804 VDD.n1245 GND 0.01fF
C1805 VDD.n1246 GND 0.02fF
C1806 VDD.n1247 GND 0.02fF
C1807 VDD.n1248 GND 0.28fF
C1808 VDD.n1249 GND 0.01fF
C1809 VDD.n1250 GND 0.02fF
C1810 VDD.n1251 GND 0.03fF
C1811 VDD.n1252 GND 0.02fF
C1812 VDD.n1253 GND 0.02fF
C1813 VDD.n1254 GND 0.02fF
C1814 VDD.n1255 GND 0.31fF
C1815 VDD.n1256 GND 0.04fF
C1816 VDD.n1257 GND 0.03fF
C1817 VDD.n1258 GND 0.02fF
C1818 VDD.n1259 GND 0.02fF
C1819 VDD.n1260 GND 0.02fF
C1820 VDD.n1261 GND 0.03fF
C1821 VDD.n1262 GND 0.02fF
C1822 VDD.n1264 GND 0.02fF
C1823 VDD.n1265 GND 0.02fF
C1824 VDD.n1266 GND 0.02fF
C1825 VDD.n1268 GND 0.28fF
C1826 VDD.n1270 GND 0.02fF
C1827 VDD.n1271 GND 0.02fF
C1828 VDD.n1272 GND 0.03fF
C1829 VDD.n1273 GND 0.02fF
C1830 VDD.n1274 GND 0.28fF
C1831 VDD.n1275 GND 0.01fF
C1832 VDD.n1276 GND 0.02fF
C1833 VDD.n1277 GND 0.03fF
C1834 VDD.n1278 GND 0.28fF
C1835 VDD.n1279 GND 0.01fF
C1836 VDD.n1280 GND 0.02fF
C1837 VDD.n1281 GND 0.02fF
C1838 VDD.n1282 GND 0.06fF
C1839 VDD.n1283 GND 0.23fF
C1840 VDD.n1284 GND 0.01fF
C1841 VDD.n1285 GND 0.01fF
C1842 VDD.n1286 GND 0.02fF
C1843 VDD.n1287 GND 0.14fF
C1844 VDD.n1288 GND 0.17fF
C1845 VDD.n1289 GND 0.01fF
C1846 VDD.n1290 GND 0.02fF
C1847 VDD.n1291 GND 0.02fF
C1848 VDD.n1292 GND 0.11fF
C1849 VDD.n1293 GND 0.02fF
C1850 VDD.n1294 GND 0.14fF
C1851 VDD.n1295 GND 0.16fF
C1852 VDD.n1296 GND 0.01fF
C1853 VDD.n1297 GND 0.02fF
C1854 VDD.n1298 GND 0.02fF
C1855 VDD.n1299 GND 0.18fF
C1856 VDD.n1300 GND 0.15fF
C1857 VDD.n1301 GND 0.01fF
C1858 VDD.n1302 GND 0.02fF
C1859 VDD.n1303 GND 0.03fF
C1860 VDD.n1304 GND 0.18fF
C1861 VDD.n1305 GND 0.15fF
C1862 VDD.n1306 GND 0.01fF
C1863 VDD.n1307 GND 0.02fF
C1864 VDD.n1308 GND 0.03fF
C1865 VDD.n1309 GND 0.14fF
C1866 VDD.n1310 GND 0.16fF
C1867 VDD.n1311 GND 0.01fF
C1868 VDD.n1312 GND 0.11fF
C1869 VDD.n1313 GND 0.02fF
C1870 VDD.n1314 GND 0.02fF
C1871 VDD.n1315 GND 0.02fF
C1872 VDD.n1316 GND 0.14fF
C1873 VDD.n1317 GND 0.17fF
C1874 VDD.n1318 GND 0.01fF
C1875 VDD.n1319 GND 0.02fF
C1876 VDD.n1320 GND 0.02fF
C1877 VDD.n1321 GND 0.22fF
C1878 VDD.n1322 GND 0.01fF
C1879 VDD.n1323 GND 0.07fF
C1880 VDD.n1324 GND 0.02fF
C1881 VDD.n1325 GND 0.28fF
C1882 VDD.n1326 GND 0.01fF
C1883 VDD.n1327 GND 0.02fF
C1884 VDD.n1328 GND 0.02fF
C1885 VDD.n1329 GND 0.28fF
C1886 VDD.n1330 GND 0.01fF
C1887 VDD.n1331 GND 0.02fF
C1888 VDD.n1332 GND 0.03fF
C1889 VDD.n1333 GND 0.02fF
C1890 VDD.n1334 GND 0.02fF
C1891 VDD.n1335 GND 0.02fF
C1892 VDD.n1336 GND 0.31fF
C1893 VDD.n1337 GND 0.04fF
C1894 VDD.n1338 GND 0.03fF
C1895 VDD.n1339 GND 0.02fF
C1896 VDD.n1340 GND 0.02fF
C1897 VDD.n1341 GND 0.02fF
C1898 VDD.n1342 GND 0.03fF
C1899 VDD.n1343 GND 0.02fF
C1900 VDD.n1345 GND 0.02fF
C1901 VDD.n1346 GND 0.02fF
C1902 VDD.n1347 GND 0.02fF
C1903 VDD.n1349 GND 0.28fF
C1904 VDD.n1351 GND 0.02fF
C1905 VDD.n1352 GND 0.02fF
C1906 VDD.n1353 GND 0.03fF
C1907 VDD.n1354 GND 0.02fF
C1908 VDD.n1355 GND 0.28fF
C1909 VDD.n1356 GND 0.01fF
C1910 VDD.n1357 GND 0.02fF
C1911 VDD.n1358 GND 0.03fF
C1912 VDD.n1359 GND 0.28fF
C1913 VDD.n1360 GND 0.01fF
C1914 VDD.n1361 GND 0.02fF
C1915 VDD.n1362 GND 0.02fF
C1916 VDD.n1363 GND 0.06fF
C1917 VDD.n1364 GND 0.23fF
C1918 VDD.n1365 GND 0.01fF
C1919 VDD.n1366 GND 0.01fF
C1920 VDD.n1367 GND 0.02fF
C1921 VDD.n1368 GND 0.14fF
C1922 VDD.n1369 GND 0.17fF
C1923 VDD.n1370 GND 0.01fF
C1924 VDD.n1371 GND 0.02fF
C1925 VDD.n1372 GND 0.02fF
C1926 VDD.n1373 GND 0.11fF
C1927 VDD.n1374 GND 0.02fF
C1928 VDD.n1375 GND 0.14fF
C1929 VDD.n1376 GND 0.16fF
C1930 VDD.n1377 GND 0.01fF
C1931 VDD.n1378 GND 0.02fF
C1932 VDD.n1379 GND 0.02fF
C1933 VDD.n1380 GND 0.18fF
C1934 VDD.n1381 GND 0.15fF
C1935 VDD.n1382 GND 0.01fF
C1936 VDD.n1383 GND 0.02fF
C1937 VDD.n1384 GND 0.03fF
C1938 VDD.n1385 GND 0.18fF
C1939 VDD.n1386 GND 0.15fF
C1940 VDD.n1387 GND 0.01fF
C1941 VDD.n1388 GND 0.02fF
C1942 VDD.n1389 GND 0.03fF
C1943 VDD.n1390 GND 0.14fF
C1944 VDD.n1391 GND 0.16fF
C1945 VDD.n1392 GND 0.01fF
C1946 VDD.n1393 GND 0.11fF
C1947 VDD.n1394 GND 0.02fF
C1948 VDD.n1395 GND 0.02fF
C1949 VDD.n1396 GND 0.02fF
C1950 VDD.n1397 GND 0.14fF
C1951 VDD.n1398 GND 0.17fF
C1952 VDD.n1399 GND 0.01fF
C1953 VDD.n1400 GND 0.02fF
C1954 VDD.n1401 GND 0.02fF
C1955 VDD.n1402 GND 0.22fF
C1956 VDD.n1403 GND 0.01fF
C1957 VDD.n1404 GND 0.07fF
C1958 VDD.n1405 GND 0.02fF
C1959 VDD.n1406 GND 0.28fF
C1960 VDD.n1407 GND 0.01fF
C1961 VDD.n1408 GND 0.02fF
C1962 VDD.n1409 GND 0.02fF
C1963 VDD.n1410 GND 0.28fF
C1964 VDD.n1411 GND 0.01fF
C1965 VDD.n1412 GND 0.02fF
C1966 VDD.n1413 GND 0.03fF
C1967 VDD.n1414 GND 0.02fF
C1968 VDD.n1415 GND 0.02fF
C1969 VDD.n1416 GND 0.02fF
C1970 VDD.n1417 GND 0.31fF
C1971 VDD.n1418 GND 0.04fF
C1972 VDD.n1419 GND 0.03fF
C1973 VDD.n1420 GND 0.02fF
C1974 VDD.n1421 GND 0.02fF
C1975 VDD.n1422 GND 0.02fF
C1976 VDD.n1423 GND 0.03fF
C1977 VDD.n1424 GND 0.02fF
C1978 VDD.n1426 GND 0.02fF
C1979 VDD.n1427 GND 0.02fF
C1980 VDD.n1428 GND 0.02fF
C1981 VDD.n1430 GND 0.28fF
C1982 VDD.n1432 GND 0.02fF
C1983 VDD.n1433 GND 0.02fF
C1984 VDD.n1434 GND 0.03fF
C1985 VDD.n1435 GND 0.02fF
C1986 VDD.n1436 GND 0.28fF
C1987 VDD.n1437 GND 0.01fF
C1988 VDD.n1438 GND 0.02fF
C1989 VDD.n1439 GND 0.03fF
C1990 VDD.n1440 GND 0.28fF
C1991 VDD.n1441 GND 0.01fF
C1992 VDD.n1442 GND 0.02fF
C1993 VDD.n1443 GND 0.02fF
C1994 VDD.n1444 GND 0.06fF
C1995 VDD.n1445 GND 0.23fF
C1996 VDD.n1446 GND 0.01fF
C1997 VDD.n1447 GND 0.01fF
C1998 VDD.n1448 GND 0.02fF
C1999 VDD.n1449 GND 0.14fF
C2000 VDD.n1450 GND 0.17fF
C2001 VDD.n1451 GND 0.01fF
C2002 VDD.n1452 GND 0.02fF
C2003 VDD.n1453 GND 0.02fF
C2004 VDD.n1454 GND 0.11fF
C2005 VDD.n1455 GND 0.02fF
C2006 VDD.n1456 GND 0.14fF
C2007 VDD.n1457 GND 0.16fF
C2008 VDD.n1458 GND 0.01fF
C2009 VDD.n1459 GND 0.02fF
C2010 VDD.n1460 GND 0.02fF
C2011 VDD.n1461 GND 0.18fF
C2012 VDD.n1462 GND 0.15fF
C2013 VDD.n1463 GND 0.01fF
C2014 VDD.n1464 GND 0.02fF
C2015 VDD.n1465 GND 0.03fF
C2016 VDD.n1466 GND 0.18fF
C2017 VDD.n1467 GND 0.15fF
C2018 VDD.n1468 GND 0.01fF
C2019 VDD.n1469 GND 0.02fF
C2020 VDD.n1470 GND 0.03fF
C2021 VDD.n1471 GND 0.14fF
C2022 VDD.n1472 GND 0.16fF
C2023 VDD.n1473 GND 0.01fF
C2024 VDD.n1474 GND 0.11fF
C2025 VDD.n1475 GND 0.02fF
C2026 VDD.n1476 GND 0.02fF
C2027 VDD.n1477 GND 0.02fF
C2028 VDD.n1478 GND 0.14fF
C2029 VDD.n1479 GND 0.17fF
C2030 VDD.n1480 GND 0.01fF
C2031 VDD.n1481 GND 0.02fF
C2032 VDD.n1482 GND 0.02fF
C2033 VDD.n1483 GND 0.22fF
C2034 VDD.n1484 GND 0.01fF
C2035 VDD.n1485 GND 0.07fF
C2036 VDD.n1486 GND 0.02fF
C2037 VDD.n1487 GND 0.28fF
C2038 VDD.n1488 GND 0.01fF
C2039 VDD.n1489 GND 0.02fF
C2040 VDD.n1490 GND 0.02fF
C2041 VDD.n1491 GND 0.28fF
C2042 VDD.n1492 GND 0.01fF
C2043 VDD.n1493 GND 0.02fF
C2044 VDD.n1494 GND 0.03fF
C2045 VDD.n1495 GND 0.02fF
C2046 VDD.n1496 GND 0.02fF
C2047 VDD.n1497 GND 0.02fF
C2048 VDD.n1498 GND 0.31fF
C2049 VDD.n1499 GND 0.04fF
C2050 VDD.n1500 GND 0.03fF
C2051 VDD.n1501 GND 0.02fF
C2052 VDD.n1502 GND 0.02fF
C2053 VDD.n1503 GND 0.02fF
C2054 VDD.n1504 GND 0.03fF
C2055 VDD.n1505 GND 0.02fF
C2056 VDD.n1507 GND 0.02fF
C2057 VDD.n1508 GND 0.02fF
C2058 VDD.n1509 GND 0.02fF
C2059 VDD.n1511 GND 0.28fF
C2060 VDD.n1513 GND 0.02fF
C2061 VDD.n1514 GND 0.02fF
C2062 VDD.n1515 GND 0.03fF
C2063 VDD.n1516 GND 0.02fF
C2064 VDD.n1517 GND 0.28fF
C2065 VDD.n1518 GND 0.01fF
C2066 VDD.n1519 GND 0.02fF
C2067 VDD.n1520 GND 0.03fF
C2068 VDD.n1521 GND 0.28fF
C2069 VDD.n1522 GND 0.01fF
C2070 VDD.n1523 GND 0.02fF
C2071 VDD.n1524 GND 0.02fF
C2072 VDD.n1525 GND 0.06fF
C2073 VDD.n1526 GND 0.23fF
C2074 VDD.n1527 GND 0.01fF
C2075 VDD.n1528 GND 0.01fF
C2076 VDD.n1529 GND 0.02fF
C2077 VDD.n1530 GND 0.14fF
C2078 VDD.n1531 GND 0.17fF
C2079 VDD.n1532 GND 0.01fF
C2080 VDD.n1533 GND 0.02fF
C2081 VDD.n1534 GND 0.02fF
C2082 VDD.n1535 GND 0.11fF
C2083 VDD.n1536 GND 0.02fF
C2084 VDD.n1537 GND 0.14fF
C2085 VDD.n1538 GND 0.16fF
C2086 VDD.n1539 GND 0.01fF
C2087 VDD.n1540 GND 0.02fF
C2088 VDD.n1541 GND 0.02fF
C2089 VDD.n1542 GND 0.18fF
C2090 VDD.n1543 GND 0.15fF
C2091 VDD.n1544 GND 0.01fF
C2092 VDD.n1545 GND 0.02fF
C2093 VDD.n1546 GND 0.03fF
C2094 VDD.n1547 GND 0.18fF
C2095 VDD.n1548 GND 0.15fF
C2096 VDD.n1549 GND 0.01fF
C2097 VDD.n1550 GND 0.02fF
C2098 VDD.n1551 GND 0.03fF
C2099 VDD.n1552 GND 0.14fF
C2100 VDD.n1553 GND 0.16fF
C2101 VDD.n1554 GND 0.01fF
C2102 VDD.n1555 GND 0.11fF
C2103 VDD.n1556 GND 0.02fF
C2104 VDD.n1557 GND 0.02fF
C2105 VDD.n1558 GND 0.02fF
C2106 VDD.n1559 GND 0.14fF
C2107 VDD.n1560 GND 0.17fF
C2108 VDD.n1561 GND 0.01fF
C2109 VDD.n1562 GND 0.02fF
C2110 VDD.n1563 GND 0.02fF
C2111 VDD.n1564 GND 0.22fF
C2112 VDD.n1565 GND 0.01fF
C2113 VDD.n1566 GND 0.07fF
C2114 VDD.n1567 GND 0.02fF
C2115 VDD.n1568 GND 0.28fF
C2116 VDD.n1569 GND 0.01fF
C2117 VDD.n1570 GND 0.02fF
C2118 VDD.n1571 GND 0.02fF
C2119 VDD.n1572 GND 0.28fF
C2120 VDD.n1573 GND 0.01fF
C2121 VDD.n1574 GND 0.02fF
C2122 VDD.n1575 GND 0.03fF
C2123 VDD.n1576 GND 0.02fF
C2124 VDD.n1577 GND 0.02fF
C2125 VDD.n1578 GND 0.02fF
C2126 VDD.n1579 GND 0.31fF
C2127 VDD.n1580 GND 0.04fF
C2128 VDD.n1581 GND 0.03fF
C2129 VDD.n1582 GND 0.02fF
C2130 VDD.n1583 GND 0.02fF
C2131 VDD.n1584 GND 0.02fF
C2132 VDD.n1585 GND 0.03fF
C2133 VDD.n1586 GND 0.02fF
C2134 VDD.n1588 GND 0.02fF
C2135 VDD.n1589 GND 0.02fF
C2136 VDD.n1590 GND 0.02fF
C2137 VDD.n1592 GND 0.28fF
C2138 VDD.n1594 GND 0.02fF
C2139 VDD.n1595 GND 0.02fF
C2140 VDD.n1596 GND 0.03fF
C2141 VDD.n1597 GND 0.02fF
C2142 VDD.n1598 GND 0.28fF
C2143 VDD.n1599 GND 0.01fF
C2144 VDD.n1600 GND 0.02fF
C2145 VDD.n1601 GND 0.03fF
C2146 VDD.n1602 GND 0.28fF
C2147 VDD.n1603 GND 0.01fF
C2148 VDD.n1604 GND 0.02fF
C2149 VDD.n1605 GND 0.02fF
C2150 VDD.n1606 GND 0.06fF
C2151 VDD.n1607 GND 0.23fF
C2152 VDD.n1608 GND 0.01fF
C2153 VDD.n1609 GND 0.01fF
C2154 VDD.n1610 GND 0.02fF
C2155 VDD.n1611 GND 0.14fF
C2156 VDD.n1612 GND 0.17fF
C2157 VDD.n1613 GND 0.01fF
C2158 VDD.n1614 GND 0.02fF
C2159 VDD.n1615 GND 0.02fF
C2160 VDD.n1616 GND 0.11fF
C2161 VDD.n1617 GND 0.02fF
C2162 VDD.n1618 GND 0.14fF
C2163 VDD.n1619 GND 0.16fF
C2164 VDD.n1620 GND 0.01fF
C2165 VDD.n1621 GND 0.02fF
C2166 VDD.n1622 GND 0.02fF
C2167 VDD.n1623 GND 0.18fF
C2168 VDD.n1624 GND 0.15fF
C2169 VDD.n1625 GND 0.01fF
C2170 VDD.n1626 GND 0.02fF
C2171 VDD.n1627 GND 0.03fF
C2172 VDD.n1628 GND 0.18fF
C2173 VDD.n1629 GND 0.15fF
C2174 VDD.n1630 GND 0.01fF
C2175 VDD.n1631 GND 0.02fF
C2176 VDD.n1632 GND 0.03fF
C2177 VDD.n1633 GND 0.14fF
C2178 VDD.n1634 GND 0.16fF
C2179 VDD.n1635 GND 0.01fF
C2180 VDD.n1636 GND 0.11fF
C2181 VDD.n1637 GND 0.02fF
C2182 VDD.n1638 GND 0.02fF
C2183 VDD.n1639 GND 0.02fF
C2184 VDD.n1640 GND 0.14fF
C2185 VDD.n1641 GND 0.17fF
C2186 VDD.n1642 GND 0.01fF
C2187 VDD.n1643 GND 0.02fF
C2188 VDD.n1644 GND 0.02fF
C2189 VDD.n1645 GND 0.22fF
C2190 VDD.n1646 GND 0.01fF
C2191 VDD.n1647 GND 0.07fF
C2192 VDD.n1648 GND 0.02fF
C2193 VDD.n1649 GND 0.28fF
C2194 VDD.n1650 GND 0.01fF
C2195 VDD.n1651 GND 0.02fF
C2196 VDD.n1652 GND 0.02fF
C2197 VDD.n1653 GND 0.28fF
C2198 VDD.n1654 GND 0.01fF
C2199 VDD.n1655 GND 0.02fF
C2200 VDD.n1656 GND 0.03fF
C2201 VDD.n1657 GND 0.02fF
C2202 VDD.n1658 GND 0.02fF
C2203 VDD.n1659 GND 0.02fF
C2204 VDD.n1660 GND 0.31fF
C2205 VDD.n1661 GND 0.04fF
C2206 VDD.n1662 GND 0.03fF
C2207 VDD.n1663 GND 0.02fF
C2208 VDD.n1664 GND 0.02fF
C2209 VDD.n1665 GND 0.02fF
C2210 VDD.n1666 GND 0.03fF
C2211 VDD.n1667 GND 0.02fF
C2212 VDD.n1669 GND 0.02fF
C2213 VDD.n1670 GND 0.02fF
C2214 VDD.n1671 GND 0.02fF
C2215 VDD.n1673 GND 0.28fF
C2216 VDD.n1675 GND 0.02fF
C2217 VDD.n1676 GND 0.02fF
C2218 VDD.n1677 GND 0.03fF
C2219 VDD.n1678 GND 0.02fF
C2220 VDD.n1679 GND 0.28fF
C2221 VDD.n1680 GND 0.01fF
C2222 VDD.n1681 GND 0.02fF
C2223 VDD.n1682 GND 0.03fF
C2224 VDD.n1683 GND 0.28fF
C2225 VDD.n1684 GND 0.01fF
C2226 VDD.n1685 GND 0.02fF
C2227 VDD.n1686 GND 0.02fF
C2228 VDD.n1687 GND 0.06fF
C2229 VDD.n1688 GND 0.23fF
C2230 VDD.n1689 GND 0.01fF
C2231 VDD.n1690 GND 0.01fF
C2232 VDD.n1691 GND 0.02fF
C2233 a_17533_1051.n0 GND 0.37fF
C2234 a_17533_1051.n1 GND 0.41fF
C2235 a_17533_1051.n2 GND 0.28fF
C2236 a_17533_1051.n3 GND 0.63fF
C2237 a_17533_1051.n4 GND 0.23fF
C2238 a_17533_1051.n5 GND 0.33fF
C2239 a_10219_989.n0 GND 0.99fF
C2240 a_10219_989.n1 GND 0.99fF
C2241 a_10219_989.n2 GND 1.16fF
C2242 a_10219_989.n3 GND 0.37fF
C2243 a_10219_989.n4 GND 0.51fF
C2244 a_10219_989.n5 GND 0.57fF
C2245 a_10219_989.t10 GND 1.08fF
C2246 a_10219_989.n6 GND 0.81fF
C2247 a_10219_989.n7 GND 0.51fF
C2248 a_10219_989.t14 GND 1.09fF
C2249 a_10219_989.n8 GND 0.70fF
C2250 a_10219_989.n9 GND 10.47fF
C2251 a_10219_989.n10 GND 1.61fF
C2252 a_10219_989.n11 GND 0.80fF
C2253 a_10219_989.t15 GND 0.88fF
C2254 a_10219_989.n12 GND 1.55fF
C2255 a_10219_989.n13 GND 1.42fF
C2256 a_10219_989.n14 GND 0.15fF
C2257 a_10219_989.n15 GND 0.42fF
C2258 a_10219_989.n16 GND 0.08fF
C2259 a_6825_103.n0 GND 0.03fF
C2260 a_6825_103.n1 GND 0.10fF
C2261 a_6825_103.n2 GND 0.10fF
C2262 a_6825_103.n3 GND 0.05fF
C2263 a_6825_103.n4 GND 0.03fF
C2264 a_6825_103.n5 GND 0.04fF
C2265 a_6825_103.n6 GND 0.11fF
C2266 a_6825_103.n7 GND 0.04fF
C2267 a_6049_1050.n0 GND 0.71fF
C2268 a_6049_1050.n1 GND 0.71fF
C2269 a_6049_1050.n2 GND 0.83fF
C2270 a_6049_1050.n3 GND 0.26fF
C2271 a_6049_1050.n4 GND 0.48fF
C2272 a_6049_1050.n5 GND 0.52fF
C2273 a_6049_1050.n6 GND 0.64fF
C2274 a_6049_1050.n7 GND 0.52fF
C2275 a_6049_1050.n8 GND 0.61fF
C2276 a_6049_1050.n9 GND 1.49fF
C2277 a_6049_1050.n10 GND 0.61fF
C2278 a_6049_1050.n11 GND 0.11fF
C2279 a_6049_1050.n12 GND 0.30fF
C2280 a_6049_1050.n13 GND 0.06fF
C2281 a_13745_1050.n0 GND 0.56fF
C2282 a_13745_1050.n1 GND 0.56fF
C2283 a_13745_1050.n2 GND 0.66fF
C2284 a_13745_1050.n3 GND 0.21fF
C2285 a_13745_1050.n4 GND 0.39fF
C2286 a_13745_1050.n5 GND 0.42fF
C2287 a_13745_1050.n6 GND 0.67fF
C2288 a_13745_1050.n7 GND 0.67fF
C2289 a_13745_1050.n8 GND 0.09fF
C2290 a_13745_1050.n9 GND 0.24fF
C2291 a_13745_1050.n10 GND 0.05fF
C2292 a_13840_210.n0 GND 0.07fF
C2293 a_13840_210.n1 GND 0.13fF
C2294 a_13840_210.n2 GND 0.07fF
C2295 a_13840_210.n3 GND 0.02fF
C2296 a_13840_210.n4 GND 0.03fF
C2297 a_13840_210.n5 GND 0.06fF
C2298 a_13840_210.n6 GND 0.05fF
C2299 a_13840_210.n7 GND 0.06fF
C2300 a_13840_210.n8 GND 0.07fF
C2301 a_13840_210.n9 GND 0.07fF
C2302 a_13840_210.n10 GND 0.03fF
C2303 a_13840_210.n11 GND 0.01fF
C2304 a_13840_210.n12 GND 0.12fF
C2305 a_13840_210.t0 GND 0.28fF
C2306 a_13105_989.n0 GND 0.90fF
C2307 a_13105_989.n1 GND 0.90fF
C2308 a_13105_989.n2 GND 1.05fF
C2309 a_13105_989.n3 GND 0.33fF
C2310 a_13105_989.n4 GND 0.46fF
C2311 a_13105_989.n5 GND 0.58fF
C2312 a_13105_989.t8 GND 0.94fF
C2313 a_13105_989.n6 GND 0.72fF
C2314 a_13105_989.n7 GND 0.58fF
C2315 a_13105_989.t7 GND 0.94fF
C2316 a_13105_989.n8 GND 0.62fF
C2317 a_13105_989.n9 GND 0.57fF
C2318 a_13105_989.t15 GND 0.94fF
C2319 a_13105_989.n10 GND 0.65fF
C2320 a_13105_989.n11 GND 2.11fF
C2321 a_13105_989.n12 GND 3.15fF
C2322 a_13105_989.n13 GND 0.77fF
C2323 a_13105_989.n14 GND 0.14fF
C2324 a_13105_989.n15 GND 0.54fF
C2325 a_13105_989.n16 GND 0.08fF
C2326 a_3258_210.n0 GND 0.02fF
C2327 a_3258_210.n1 GND 0.07fF
C2328 a_3258_210.n2 GND 0.13fF
C2329 a_3258_210.n3 GND 0.09fF
C2330 a_3258_210.t1 GND 0.25fF
C2331 a_3258_210.n4 GND 0.05fF
C2332 a_3258_210.n5 GND 0.06fF
C2333 a_3258_210.n6 GND 0.07fF
C2334 a_3258_210.n7 GND 0.07fF
C2335 a_3258_210.n8 GND 0.03fF
C2336 a_3258_210.n9 GND 0.01fF
C2337 a_3258_210.n10 GND 0.11fF
C2338 a_3258_210.n11 GND 0.02fF
C2339 a_3258_210.n12 GND 0.05fF
C2340 a_3258_210.n13 GND 0.02fF
C2341 a_2977_103.n0 GND 0.03fF
C2342 a_2977_103.n1 GND 0.10fF
C2343 a_2977_103.n2 GND 0.10fF
C2344 a_2977_103.n3 GND 0.05fF
C2345 a_2977_103.n4 GND 0.03fF
C2346 a_2977_103.n5 GND 0.04fF
C2347 a_2977_103.n6 GND 0.11fF
C2348 a_2977_103.n7 GND 0.04fF
.ends
