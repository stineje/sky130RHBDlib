// File: DFFX1.spi.pex
// Created: Tue Oct 15 15:48:13 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_DFFX1\%GND ( 1 39 43 46 51 61 69 77 83 89 97 105 113 121 132 136 138 \
 141 143 145 148 149 150 151 152 153 )
c263 ( 153 0 ) capacitor c=0.0208017f //x=19.12 //y=0.865
c264 ( 152 0 ) capacitor c=0.0208124f //x=15.79 //y=0.865
c265 ( 151 0 ) capacitor c=0.0208017f //x=12.46 //y=0.865
c266 ( 150 0 ) capacitor c=0.0208017f //x=9.13 //y=0.865
c267 ( 149 0 ) capacitor c=0.0208019f //x=5.8 //y=0.865
c268 ( 148 0 ) capacitor c=0.022675f //x=0.885 //y=0.875
c269 ( 147 0 ) capacitor c=0.00440095f //x=19.24 //y=0
c270 ( 145 0 ) capacitor c=0.107063f //x=18.13 //y=0
c271 ( 144 0 ) capacitor c=0.00440095f //x=15.98 //y=0
c272 ( 143 0 ) capacitor c=0.107594f //x=14.8 //y=0
c273 ( 142 0 ) capacitor c=0.00440095f //x=12.65 //y=0
c274 ( 141 0 ) capacitor c=0.107063f //x=11.47 //y=0
c275 ( 140 0 ) capacitor c=0.00440095f //x=9.25 //y=0
c276 ( 138 0 ) capacitor c=0.107063f //x=8.14 //y=0
c277 ( 137 0 ) capacitor c=0.00440095f //x=5.99 //y=0
c278 ( 136 0 ) capacitor c=0.109996f //x=4.81 //y=0
c279 ( 135 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c280 ( 132 0 ) capacitor c=0.25934f //x=21.09 //y=0
c281 ( 121 0 ) capacitor c=0.0389288f //x=19.225 //y=0
c282 ( 113 0 ) capacitor c=0.0720403f //x=17.96 //y=0
c283 ( 105 0 ) capacitor c=0.0426751f //x=15.895 //y=0
c284 ( 97 0 ) capacitor c=0.0751168f //x=14.63 //y=0
c285 ( 89 0 ) capacitor c=0.0389288f //x=12.565 //y=0
c286 ( 83 0 ) capacitor c=0.0720403f //x=11.3 //y=0
c287 ( 77 0 ) capacitor c=0.0389288f //x=9.235 //y=0
c288 ( 69 0 ) capacitor c=0.0720423f //x=7.97 //y=0
c289 ( 61 0 ) capacitor c=0.0389288f //x=5.905 //y=0
c290 ( 51 0 ) capacitor c=0.131745f //x=4.64 //y=0
c291 ( 46 0 ) capacitor c=0.178285f //x=0.74 //y=0
c292 ( 43 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c293 ( 39 0 ) capacitor c=0.711045f //x=21.09 //y=0
r294 (  130 132 ) resistor r=26.5322 //w=0.357 //l=0.74 //layer=li \
 //thickness=0.1 //x=20.35 //y=0 //x2=21.09 //y2=0
r295 (  128 147 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.395 //y=0 //x2=19.31 //y2=0
r296 (  128 130 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=19.395 //y=0 //x2=20.35 //y2=0
r297 (  123 147 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.31 //y=0.17 //x2=19.31 //y2=0
r298 (  123 153 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=19.31 //y=0.17 //x2=19.31 //y2=0.955
r299 (  122 145 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.3 //y=0 //x2=18.13 //y2=0
r300 (  121 147 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.225 //y=0 //x2=19.31 //y2=0
r301 (  121 122 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=19.225 //y=0 //x2=18.3 //y2=0
r302 (  116 118 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=16.65 //y=0 //x2=17.76 //y2=0
r303 (  114 144 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.065 //y=0 //x2=15.98 //y2=0
r304 (  114 116 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=16.065 //y=0 //x2=16.65 //y2=0
r305 (  113 145 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.96 //y=0 //x2=18.13 //y2=0
r306 (  113 118 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=17.96 //y=0 //x2=17.76 //y2=0
r307 (  109 144 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.98 //y=0.17 //x2=15.98 //y2=0
r308 (  109 152 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=15.98 //y=0.17 //x2=15.98 //y2=0.955
r309 (  106 143 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.97 //y=0 //x2=14.8 //y2=0
r310 (  106 108 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.97 //y=0 //x2=15.54 //y2=0
r311 (  105 144 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.895 //y=0 //x2=15.98 //y2=0
r312 (  105 108 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=15.895 //y=0 //x2=15.54 //y2=0
r313 (  100 102 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=12.95 //y=0 //x2=14.06 //y2=0
r314 (  98 142 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.735 //y=0 //x2=12.65 //y2=0
r315 (  98 100 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=12.735 //y=0 //x2=12.95 //y2=0
r316 (  97 143 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.63 //y=0 //x2=14.8 //y2=0
r317 (  97 102 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.63 //y=0 //x2=14.06 //y2=0
r318 (  93 142 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.65 //y=0.17 //x2=12.65 //y2=0
r319 (  93 151 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=12.65 //y=0.17 //x2=12.65 //y2=0.955
r320 (  90 141 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.64 //y=0 //x2=11.47 //y2=0
r321 (  90 92 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=11.64 //y=0 //x2=11.84 //y2=0
r322 (  89 142 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.565 //y=0 //x2=12.65 //y2=0
r323 (  89 92 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=12.565 //y=0 //x2=11.84 //y2=0
r324 (  84 140 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.405 //y=0 //x2=9.32 //y2=0
r325 (  84 86 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=9.405 //y=0 //x2=10.36 //y2=0
r326 (  83 141 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.3 //y=0 //x2=11.47 //y2=0
r327 (  83 86 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=11.3 //y=0 //x2=10.36 //y2=0
r328 (  79 140 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.32 //y=0.17 //x2=9.32 //y2=0
r329 (  79 150 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=9.32 //y=0.17 //x2=9.32 //y2=0.955
r330 (  78 138 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=0 //x2=8.14 //y2=0
r331 (  77 140 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.235 //y=0 //x2=9.32 //y2=0
r332 (  77 78 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=9.235 //y=0 //x2=8.31 //y2=0
r333 (  72 74 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r334 (  70 137 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.075 //y=0 //x2=5.99 //y2=0
r335 (  70 72 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=6.075 //y=0 //x2=6.66 //y2=0
r336 (  69 138 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=8.14 //y2=0
r337 (  69 74 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=7.77 //y2=0
r338 (  65 137 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.99 //y=0.17 //x2=5.99 //y2=0
r339 (  65 149 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=5.99 //y=0.17 //x2=5.99 //y2=0.955
r340 (  62 136 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=4.81 //y2=0
r341 (  62 64 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=5.55 //y2=0
r342 (  61 137 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.905 //y=0 //x2=5.99 //y2=0
r343 (  61 64 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=5.905 //y=0 //x2=5.55 //y2=0
r344 (  56 58 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r345 (  54 56 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r346 (  52 135 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r347 (  52 54 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r348 (  51 136 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.81 //y2=0
r349 (  51 58 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r350 (  47 135 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r351 (  47 148 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r352 (  43 135 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r353 (  43 46 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r354 (  39 132 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r355 (  37 130 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=0 //x2=20.35 //y2=0
r356 (  37 39 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=0 //x2=21.09 //y2=0
r357 (  35 147 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.24 //y=0 //x2=19.24 //y2=0
r358 (  35 37 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.24 //y=0 //x2=20.35 //y2=0
r359 (  33 118 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=0 //x2=17.76 //y2=0
r360 (  33 35 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=0 //x2=19.24 //y2=0
r361 (  31 116 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=0 //x2=16.65 //y2=0
r362 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=0 //x2=17.76 //y2=0
r363 (  29 108 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.54 //y=0 //x2=15.54 //y2=0
r364 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.54 //y=0 //x2=16.65 //y2=0
r365 (  27 102 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=0 //x2=14.06 //y2=0
r366 (  27 29 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=0 //x2=15.54 //y2=0
r367 (  25 100 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.95 //y=0 //x2=12.95 //y2=0
r368 (  25 27 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.95 //y=0 //x2=14.06 //y2=0
r369 (  23 92 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.84 //y=0 //x2=11.84 //y2=0
r370 (  23 25 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.84 //y=0 //x2=12.95 //y2=0
r371 (  20 86 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r372 (  18 140 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=0 //x2=9.25 //y2=0
r373 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=0 //x2=10.36 //y2=0
r374 (  16 74 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r375 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=9.25 //y2=0
r376 (  14 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r377 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r378 (  12 64 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r379 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r380 (  10 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r381 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r382 (  8 56 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r383 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r384 (  6 54 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r385 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r386 (  3 46 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r387 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r388 (  1 23 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=0 //x2=11.84 //y2=0
r389 (  1 20 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=0 //x2=10.36 //y2=0
ends PM_DFFX1\%GND

subckt PM_DFFX1\%VDD ( 1 52 59 66 76 86 96 102 112 122 132 136 146 156 166 170 \
 180 190 200 204 214 224 234 238 248 258 276 281 286 291 296 300 301 302 303 \
 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 )
c291 ( 319 0 ) capacitor c=0.038101f //x=20.535 //y=5.02
c292 ( 318 0 ) capacitor c=0.0239699f //x=19.655 //y=5.02
c293 ( 317 0 ) capacitor c=0.0492585f //x=18.785 //y=5.02
c294 ( 316 0 ) capacitor c=0.0380439f //x=17.205 //y=5.02
c295 ( 315 0 ) capacitor c=0.0239704f //x=16.325 //y=5.02
c296 ( 314 0 ) capacitor c=0.0492585f //x=15.455 //y=5.02
c297 ( 313 0 ) capacitor c=0.0380384f //x=13.875 //y=5.02
c298 ( 312 0 ) capacitor c=0.0238899f //x=12.995 //y=5.02
c299 ( 311 0 ) capacitor c=0.048923f //x=12.125 //y=5.02
c300 ( 310 0 ) capacitor c=0.0379613f //x=10.545 //y=5.02
c301 ( 309 0 ) capacitor c=0.0238906f //x=9.665 //y=5.02
c302 ( 308 0 ) capacitor c=0.048923f //x=8.795 //y=5.02
c303 ( 307 0 ) capacitor c=0.0379613f //x=7.215 //y=5.02
c304 ( 306 0 ) capacitor c=0.0238906f //x=6.335 //y=5.02
c305 ( 305 0 ) capacitor c=0.0491017f //x=5.465 //y=5.02
c306 ( 304 0 ) capacitor c=0.0450944f //x=3.585 //y=5.02
c307 ( 303 0 ) capacitor c=0.0240346f //x=2.705 //y=5.02
c308 ( 302 0 ) capacitor c=0.0241226f //x=1.825 //y=5.02
c309 ( 301 0 ) capacitor c=0.0530167f //x=0.955 //y=5.02
c310 ( 300 0 ) capacitor c=0.243962f //x=20.72 //y=7.4
c311 ( 298 0 ) capacitor c=0.00591168f //x=19.8 //y=7.4
c312 ( 297 0 ) capacitor c=0.00617226f //x=18.92 //y=7.4
c313 ( 296 0 ) capacitor c=0.116587f //x=18.13 //y=7.4
c314 ( 295 0 ) capacitor c=0.00591168f //x=17.39 //y=7.4
c315 ( 293 0 ) capacitor c=0.00591168f //x=16.47 //y=7.4
c316 ( 292 0 ) capacitor c=0.00617226f //x=15.59 //y=7.4
c317 ( 291 0 ) capacitor c=0.116067f //x=14.8 //y=7.4
c318 ( 290 0 ) capacitor c=0.00591168f //x=14.06 //y=7.4
c319 ( 288 0 ) capacitor c=0.00591168f //x=13.14 //y=7.4
c320 ( 287 0 ) capacitor c=0.00617226f //x=12.26 //y=7.4
c321 ( 286 0 ) capacitor c=0.114265f //x=11.47 //y=7.4
c322 ( 285 0 ) capacitor c=0.00591168f //x=10.73 //y=7.4
c323 ( 283 0 ) capacitor c=0.00591168f //x=9.81 //y=7.4
c324 ( 282 0 ) capacitor c=0.00617226f //x=8.93 //y=7.4
c325 ( 281 0 ) capacitor c=0.114394f //x=8.14 //y=7.4
c326 ( 280 0 ) capacitor c=0.00591168f //x=7.4 //y=7.4
c327 ( 278 0 ) capacitor c=0.00591168f //x=6.48 //y=7.4
c328 ( 277 0 ) capacitor c=0.00617226f //x=5.6 //y=7.4
c329 ( 276 0 ) capacitor c=0.134457f //x=4.81 //y=7.4
c330 ( 275 0 ) capacitor c=0.00617226f //x=3.73 //y=7.4
c331 ( 274 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c332 ( 273 0 ) capacitor c=0.00643014f //x=1.97 //y=7.4
c333 ( 272 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c334 ( 258 0 ) capacitor c=0.0286919f //x=20.595 //y=7.4
c335 ( 248 0 ) capacitor c=0.0291225f //x=19.715 //y=7.4
c336 ( 238 0 ) capacitor c=0.0246165f //x=18.835 //y=7.4
c337 ( 234 0 ) capacitor c=0.0244015f //x=17.96 //y=7.4
c338 ( 224 0 ) capacitor c=0.0291231f //x=17.265 //y=7.4
c339 ( 214 0 ) capacitor c=0.0291225f //x=16.385 //y=7.4
c340 ( 204 0 ) capacitor c=0.0246165f //x=15.505 //y=7.4
c341 ( 200 0 ) capacitor c=0.0244737f //x=14.63 //y=7.4
c342 ( 190 0 ) capacitor c=0.029119f //x=13.935 //y=7.4
c343 ( 180 0 ) capacitor c=0.0290962f //x=13.055 //y=7.4
c344 ( 170 0 ) capacitor c=0.0246165f //x=12.175 //y=7.4
c345 ( 166 0 ) capacitor c=0.0244015f //x=11.3 //y=7.4
c346 ( 156 0 ) capacitor c=0.0290951f //x=10.605 //y=7.4
c347 ( 146 0 ) capacitor c=0.0290962f //x=9.725 //y=7.4
c348 ( 136 0 ) capacitor c=0.0246165f //x=8.845 //y=7.4
c349 ( 132 0 ) capacitor c=0.0244015f //x=7.97 //y=7.4
c350 ( 122 0 ) capacitor c=0.0290951f //x=7.275 //y=7.4
c351 ( 112 0 ) capacitor c=0.0290962f //x=6.395 //y=7.4
c352 ( 102 0 ) capacitor c=0.0246165f //x=5.515 //y=7.4
c353 ( 96 0 ) capacitor c=0.0399852f //x=4.64 //y=7.4
c354 ( 86 0 ) capacitor c=0.0296265f //x=3.645 //y=7.4
c355 ( 76 0 ) capacitor c=0.0290098f //x=2.765 //y=7.4
c356 ( 66 0 ) capacitor c=0.0290308f //x=1.885 //y=7.4
c357 ( 59 0 ) capacitor c=0.234214f //x=0.37 //y=7.4
c358 ( 56 0 ) capacitor c=0.045728f //x=1.005 //y=7.4
c359 ( 52 0 ) capacitor c=0.745722f //x=20.72 //y=7.4
r360 (  262 300 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.68 //y=7.23 //x2=20.68 //y2=7.4
r361 (  262 319 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.68 //y=7.23 //x2=20.68 //y2=6.745
r362 (  259 298 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.885 //y=7.4 //x2=19.8 //y2=7.4
r363 (  259 261 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=19.885 //y=7.4 //x2=19.98 //y2=7.4
r364 (  258 300 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.595 //y=7.4 //x2=20.68 //y2=7.4
r365 (  258 261 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=20.595 //y=7.4 //x2=19.98 //y2=7.4
r366 (  252 298 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.8 //y=7.23 //x2=19.8 //y2=7.4
r367 (  252 318 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=19.8 //y=7.23 //x2=19.8 //y2=6.745
r368 (  249 297 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.005 //y=7.4 //x2=18.92 //y2=7.4
r369 (  249 251 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=19.005 //y=7.4 //x2=19.24 //y2=7.4
r370 (  248 298 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.715 //y=7.4 //x2=19.8 //y2=7.4
r371 (  248 251 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=19.715 //y=7.4 //x2=19.24 //y2=7.4
r372 (  242 297 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.92 //y=7.23 //x2=18.92 //y2=7.4
r373 (  242 317 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=18.92 //y=7.23 //x2=18.92 //y2=6.405
r374 (  239 296 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.3 //y=7.4 //x2=18.13 //y2=7.4
r375 (  239 241 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=18.3 //y=7.4 //x2=18.5 //y2=7.4
r376 (  238 297 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.835 //y=7.4 //x2=18.92 //y2=7.4
r377 (  238 241 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=18.835 //y=7.4 //x2=18.5 //y2=7.4
r378 (  235 295 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.435 //y=7.4 //x2=17.35 //y2=7.4
r379 (  234 296 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.96 //y=7.4 //x2=18.13 //y2=7.4
r380 (  234 235 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=17.96 //y=7.4 //x2=17.435 //y2=7.4
r381 (  228 295 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.35 //y=7.23 //x2=17.35 //y2=7.4
r382 (  228 316 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.35 //y=7.23 //x2=17.35 //y2=6.745
r383 (  225 293 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.555 //y=7.4 //x2=16.47 //y2=7.4
r384 (  225 227 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=16.555 //y=7.4 //x2=16.65 //y2=7.4
r385 (  224 295 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.265 //y=7.4 //x2=17.35 //y2=7.4
r386 (  224 227 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=17.265 //y=7.4 //x2=16.65 //y2=7.4
r387 (  218 293 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.47 //y=7.23 //x2=16.47 //y2=7.4
r388 (  218 315 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.47 //y=7.23 //x2=16.47 //y2=6.745
r389 (  215 292 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.675 //y=7.4 //x2=15.59 //y2=7.4
r390 (  215 217 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=15.675 //y=7.4 //x2=15.91 //y2=7.4
r391 (  214 293 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.385 //y=7.4 //x2=16.47 //y2=7.4
r392 (  214 217 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=16.385 //y=7.4 //x2=15.91 //y2=7.4
r393 (  208 292 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.59 //y=7.23 //x2=15.59 //y2=7.4
r394 (  208 314 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=15.59 //y=7.23 //x2=15.59 //y2=6.405
r395 (  205 291 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.97 //y=7.4 //x2=14.8 //y2=7.4
r396 (  205 207 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=14.97 //y=7.4 //x2=15.17 //y2=7.4
r397 (  204 292 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.505 //y=7.4 //x2=15.59 //y2=7.4
r398 (  204 207 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=15.505 //y=7.4 //x2=15.17 //y2=7.4
r399 (  201 290 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.105 //y=7.4 //x2=14.02 //y2=7.4
r400 (  200 291 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.63 //y=7.4 //x2=14.8 //y2=7.4
r401 (  200 201 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=14.63 //y=7.4 //x2=14.105 //y2=7.4
r402 (  194 290 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.02 //y=7.23 //x2=14.02 //y2=7.4
r403 (  194 313 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.02 //y=7.23 //x2=14.02 //y2=6.745
r404 (  191 288 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.225 //y=7.4 //x2=13.14 //y2=7.4
r405 (  191 193 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=13.225 //y=7.4 //x2=13.32 //y2=7.4
r406 (  190 290 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.935 //y=7.4 //x2=14.02 //y2=7.4
r407 (  190 193 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.935 //y=7.4 //x2=13.32 //y2=7.4
r408 (  184 288 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.14 //y=7.23 //x2=13.14 //y2=7.4
r409 (  184 312 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=13.14 //y=7.23 //x2=13.14 //y2=6.745
r410 (  181 287 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.345 //y=7.4 //x2=12.26 //y2=7.4
r411 (  181 183 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=12.345 //y=7.4 //x2=12.58 //y2=7.4
r412 (  180 288 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.055 //y=7.4 //x2=13.14 //y2=7.4
r413 (  180 183 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=13.055 //y=7.4 //x2=12.58 //y2=7.4
r414 (  174 287 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.26 //y=7.23 //x2=12.26 //y2=7.4
r415 (  174 311 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=12.26 //y=7.23 //x2=12.26 //y2=6.405
r416 (  171 286 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.64 //y=7.4 //x2=11.47 //y2=7.4
r417 (  171 173 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=11.64 //y=7.4 //x2=11.84 //y2=7.4
r418 (  170 287 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.175 //y=7.4 //x2=12.26 //y2=7.4
r419 (  170 173 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=12.175 //y=7.4 //x2=11.84 //y2=7.4
r420 (  167 285 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.775 //y=7.4 //x2=10.69 //y2=7.4
r421 (  166 286 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.3 //y=7.4 //x2=11.47 //y2=7.4
r422 (  166 167 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=11.3 //y=7.4 //x2=10.775 //y2=7.4
r423 (  160 285 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.69 //y=7.23 //x2=10.69 //y2=7.4
r424 (  160 310 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.69 //y=7.23 //x2=10.69 //y2=6.745
r425 (  157 283 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.895 //y=7.4 //x2=9.81 //y2=7.4
r426 (  157 159 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=9.895 //y=7.4 //x2=9.99 //y2=7.4
r427 (  156 285 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.605 //y=7.4 //x2=10.69 //y2=7.4
r428 (  156 159 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.605 //y=7.4 //x2=9.99 //y2=7.4
r429 (  150 283 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.81 //y=7.23 //x2=9.81 //y2=7.4
r430 (  150 309 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.81 //y=7.23 //x2=9.81 //y2=6.745
r431 (  147 282 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.015 //y=7.4 //x2=8.93 //y2=7.4
r432 (  147 149 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=9.015 //y=7.4 //x2=9.25 //y2=7.4
r433 (  146 283 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.725 //y=7.4 //x2=9.81 //y2=7.4
r434 (  146 149 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=9.725 //y=7.4 //x2=9.25 //y2=7.4
r435 (  140 282 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.93 //y=7.23 //x2=8.93 //y2=7.4
r436 (  140 308 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=8.93 //y=7.23 //x2=8.93 //y2=6.405
r437 (  137 281 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=7.4 //x2=8.14 //y2=7.4
r438 (  137 139 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=8.31 //y=7.4 //x2=8.51 //y2=7.4
r439 (  136 282 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.845 //y=7.4 //x2=8.93 //y2=7.4
r440 (  136 139 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=8.845 //y=7.4 //x2=8.51 //y2=7.4
r441 (  133 280 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.445 //y=7.4 //x2=7.36 //y2=7.4
r442 (  132 281 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=8.14 //y2=7.4
r443 (  132 133 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=7.445 //y2=7.4
r444 (  126 280 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.36 //y=7.23 //x2=7.36 //y2=7.4
r445 (  126 307 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.36 //y=7.23 //x2=7.36 //y2=6.745
r446 (  123 278 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.565 //y=7.4 //x2=6.48 //y2=7.4
r447 (  123 125 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=6.565 //y=7.4 //x2=6.66 //y2=7.4
r448 (  122 280 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.275 //y=7.4 //x2=7.36 //y2=7.4
r449 (  122 125 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=7.275 //y=7.4 //x2=6.66 //y2=7.4
r450 (  116 278 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.48 //y=7.23 //x2=6.48 //y2=7.4
r451 (  116 306 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.48 //y=7.23 //x2=6.48 //y2=6.745
r452 (  113 277 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.685 //y=7.4 //x2=5.6 //y2=7.4
r453 (  113 115 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=5.685 //y=7.4 //x2=5.92 //y2=7.4
r454 (  112 278 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.395 //y=7.4 //x2=6.48 //y2=7.4
r455 (  112 115 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=6.395 //y=7.4 //x2=5.92 //y2=7.4
r456 (  106 277 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.6 //y=7.23 //x2=5.6 //y2=7.4
r457 (  106 305 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.6 //y=7.23 //x2=5.6 //y2=6.405
r458 (  103 276 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r459 (  103 105 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=5.18 //y2=7.4
r460 (  102 277 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.515 //y=7.4 //x2=5.6 //y2=7.4
r461 (  102 105 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=5.515 //y=7.4 //x2=5.18 //y2=7.4
r462 (  97 275 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r463 (  97 99 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r464 (  96 276 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r465 (  96 99 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r466 (  90 275 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r467 (  90 304 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r468 (  87 274 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r469 (  87 89 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=3.33 //y2=7.4
r470 (  86 275 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r471 (  86 89 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.33 //y2=7.4
r472 (  80 274 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r473 (  80 303 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r474 (  77 273 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r475 (  77 79 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=2.22 //y2=7.4
r476 (  76 274 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r477 (  76 79 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.22 //y2=7.4
r478 (  70 273 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r479 (  70 302 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r480 (  67 272 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r481 (  67 69 ) resistor r=10.9356 //w=0.357 //l=0.305 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.48 //y2=7.4
r482 (  66 273 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r483 (  66 69 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.48 //y2=7.4
r484 (  60 272 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r485 (  60 301 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r486 (  56 272 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r487 (  56 59 ) resistor r=22.7675 //w=0.357 //l=0.635 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.37 //y2=7.4
r488 (  52 300 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=20.72 //y=7.4 //x2=20.72 //y2=7.4
r489 (  50 261 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=19.98 //y=7.4 //x2=19.98 //y2=7.4
r490 (  50 52 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=7.397 //x2=20.72 //y2=7.397
r491 (  48 251 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=19.24 //y=7.4 //x2=19.24 //y2=7.4
r492 (  48 50 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=19.24 //y=7.397 //x2=19.98 //y2=7.397
r493 (  46 241 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=18.5 //y=7.4 //x2=18.5 //y2=7.4
r494 (  46 48 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=7.397 //x2=19.24 //y2=7.397
r495 (  44 295 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r496 (  44 46 ) resistor r=0.453431 //w=0.306 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.397 //x2=18.5 //y2=7.397
r497 (  42 227 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=16.65 //y=7.4 //x2=16.65 //y2=7.4
r498 (  42 44 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=7.397 //x2=17.39 //y2=7.397
r499 (  40 217 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=15.91 //y=7.4 //x2=15.91 //y2=7.4
r500 (  40 42 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=15.91 //y=7.397 //x2=16.65 //y2=7.397
r501 (  38 207 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r502 (  38 40 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.397 //x2=15.91 //y2=7.397
r503 (  36 290 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=14.06 //y=7.4 //x2=14.06 //y2=7.4
r504 (  36 38 ) resistor r=0.453431 //w=0.306 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=7.397 //x2=15.17 //y2=7.397
r505 (  34 193 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=13.32 //y=7.4 //x2=13.32 //y2=7.4
r506 (  34 36 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=13.32 //y=7.397 //x2=14.06 //y2=7.397
r507 (  32 183 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r508 (  32 34 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.397 //x2=13.32 //y2=7.397
r509 (  30 173 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=11.84 //y=7.4 //x2=11.84 //y2=7.4
r510 (  30 32 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=11.84 //y=7.397 //x2=12.58 //y2=7.397
r511 (  26 159 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=9.99 //y=7.4 //x2=9.99 //y2=7.4
r512 (  24 149 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=9.25 //y=7.4 //x2=9.25 //y2=7.4
r513 (  24 26 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=7.397 //x2=9.99 //y2=7.397
r514 (  22 139 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=8.51 //y=7.4 //x2=8.51 //y2=7.4
r515 (  22 24 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=8.51 //y=7.397 //x2=9.25 //y2=7.397
r516 (  20 280 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=7.4 //y=7.4 //x2=7.4 //y2=7.4
r517 (  20 22 ) resistor r=0.453431 //w=0.306 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.4 //y=7.397 //x2=8.51 //y2=7.397
r518 (  18 125 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r519 (  18 20 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.397 //x2=7.4 //y2=7.397
r520 (  16 115 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=5.92 //y=7.4 //x2=5.92 //y2=7.4
r521 (  16 18 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=7.397 //x2=6.66 //y2=7.397
r522 (  14 105 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=5.18 //y=7.4 //x2=5.18 //y2=7.4
r523 (  14 16 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=5.18 //y=7.397 //x2=5.92 //y2=7.397
r524 (  12 99 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r525 (  12 14 ) resistor r=0.453431 //w=0.306 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.397 //x2=5.18 //y2=7.397
r526 (  10 89 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=7.4 //x2=3.33 //y2=7.4
r527 (  10 12 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=7.397 //x2=4.07 //y2=7.397
r528 (  8 79 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=2.22 //y=7.4 //x2=2.22 //y2=7.4
r529 (  8 10 ) resistor r=0.453431 //w=0.306 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.22 //y=7.397 //x2=3.33 //y2=7.397
r530 (  6 69 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.48 //y=7.4 //x2=1.48 //y2=7.4
r531 (  6 8 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=1.48 //y=7.397 //x2=2.22 //y2=7.397
r532 (  3 59 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=0.37 //y=7.4 //x2=0.37 //y2=7.4
r533 (  3 6 ) resistor r=0.453431 //w=0.306 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.37 //y=7.397 //x2=1.48 //y2=7.397
r534 (  1 285 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=10.73 //y=7.4 //x2=10.73 //y2=7.4
r535 (  1 30 ) resistor r=0.453431 //w=0.306 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=7.397 //x2=11.84 //y2=7.397
r536 (  1 26 ) resistor r=0.302288 //w=0.306 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=7.397 //x2=9.99 //y2=7.397
ends PM_DFFX1\%VDD

subckt PM_DFFX1\%noxref_3 ( 1 2 3 4 12 25 26 37 39 40 44 46 53 54 55 56 57 58 \
 59 63 64 65 70 72 75 76 77 78 79 80 84 86 89 90 95 96 101 110 113 115 116 )
c232 ( 116 0 ) capacitor c=0.0220291f //x=6.775 //y=5.02
c233 ( 115 0 ) capacitor c=0.0217503f //x=5.895 //y=5.02
c234 ( 113 0 ) capacitor c=0.00866655f //x=6.77 //y=0.905
c235 ( 110 0 ) capacitor c=0.0588816f //x=9.25 //y=4.7
c236 ( 101 0 ) capacitor c=0.058931f //x=3.33 //y=4.7
c237 ( 96 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c238 ( 95 0 ) capacitor c=0.0464411f //x=3.33 //y=2.08
c239 ( 90 0 ) capacitor c=0.0318948f //x=9.585 //y=1.21
c240 ( 89 0 ) capacitor c=0.0187384f //x=9.585 //y=0.865
c241 ( 86 0 ) capacitor c=0.0141798f //x=9.43 //y=1.365
c242 ( 84 0 ) capacitor c=0.0149844f //x=9.43 //y=0.71
c243 ( 80 0 ) capacitor c=0.0853292f //x=9.055 //y=1.915
c244 ( 79 0 ) capacitor c=0.0229722f //x=9.055 //y=1.52
c245 ( 78 0 ) capacitor c=0.0234352f //x=9.055 //y=1.21
c246 ( 77 0 ) capacitor c=0.0199343f //x=9.055 //y=0.865
c247 ( 76 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c248 ( 75 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c249 ( 72 0 ) capacitor c=0.0158629f //x=3.695 //y=1.415
c250 ( 70 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c251 ( 65 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c252 ( 64 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c253 ( 63 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c254 ( 59 0 ) capacitor c=0.110275f //x=9.59 //y=6.02
c255 ( 58 0 ) capacitor c=0.154305f //x=9.15 //y=6.02
c256 ( 57 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c257 ( 56 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c258 ( 53 0 ) capacitor c=0.00211606f //x=6.92 //y=5.2
c259 ( 46 0 ) capacitor c=0.0917424f //x=9.25 //y=2.08
c260 ( 44 0 ) capacitor c=0.108359f //x=7.4 //y=3.33
c261 ( 40 0 ) capacitor c=0.00498573f //x=7.045 //y=1.655
c262 ( 39 0 ) capacitor c=0.0136303f //x=7.315 //y=1.655
c263 ( 37 0 ) capacitor c=0.0137516f //x=7.315 //y=5.2
c264 ( 26 0 ) capacitor c=0.00251635f //x=6.125 //y=5.2
c265 ( 25 0 ) capacitor c=0.0142417f //x=6.835 //y=5.2
c266 ( 12 0 ) capacitor c=0.0883349f //x=3.33 //y=2.08
c267 ( 4 0 ) capacitor c=0.0042919f //x=7.515 //y=3.33
c268 ( 3 0 ) capacitor c=0.0617718f //x=9.135 //y=3.33
c269 ( 2 0 ) capacitor c=0.0149802f //x=3.445 //y=3.33
c270 ( 1 0 ) capacitor c=0.108369f //x=7.285 //y=3.33
r271 (  108 110 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=9.15 //y=4.7 //x2=9.25 //y2=4.7
r272 (  95 96 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r273 (  91 110 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=9.59 //y=4.865 //x2=9.25 //y2=4.7
r274 (  90 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.585 //y=1.21 //x2=9.545 //y2=1.365
r275 (  89 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.585 //y=0.865 //x2=9.545 //y2=0.71
r276 (  89 90 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.585 //y=0.865 //x2=9.585 //y2=1.21
r277 (  87 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.21 //y=1.365 //x2=9.095 //y2=1.365
r278 (  86 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.43 //y=1.365 //x2=9.545 //y2=1.365
r279 (  85 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.21 //y=0.71 //x2=9.095 //y2=0.71
r280 (  84 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.43 //y=0.71 //x2=9.545 //y2=0.71
r281 (  84 85 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=9.43 //y=0.71 //x2=9.21 //y2=0.71
r282 (  81 108 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=9.15 //y=4.865 //x2=9.15 //y2=4.7
r283 (  80 105 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.915 //x2=9.25 //y2=2.08
r284 (  79 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.52 //x2=9.095 //y2=1.365
r285 (  79 80 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.52 //x2=9.055 //y2=1.915
r286 (  78 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.21 //x2=9.095 //y2=1.365
r287 (  77 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.055 //y=0.865 //x2=9.095 //y2=0.71
r288 (  77 78 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.055 //y=0.865 //x2=9.055 //y2=1.21
r289 (  76 103 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r290 (  75 102 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r291 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r292 (  73 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r293 (  72 103 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r294 (  71 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r295 (  70 102 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r296 (  70 71 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r297 (  67 101 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r298 (  65 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r299 (  65 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r300 (  64 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r301 (  63 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r302 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r303 (  60 101 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r304 (  59 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.59 //y=6.02 //x2=9.59 //y2=4.865
r305 (  58 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.15 //y=6.02 //x2=9.15 //y2=4.865
r306 (  57 67 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r307 (  56 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r308 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.32 //y=1.365 //x2=9.43 //y2=1.365
r309 (  55 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.32 //y=1.365 //x2=9.21 //y2=1.365
r310 (  54 72 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r311 (  54 73 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r312 (  51 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=4.7 //x2=9.25 //y2=4.7
r313 (  49 51 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=9.25 //y=3.33 //x2=9.25 //y2=4.7
r314 (  46 105 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=2.08 //x2=9.25 //y2=2.08
r315 (  46 49 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.08 //x2=9.25 //y2=3.33
r316 (  42 44 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=7.4 //y=5.115 //x2=7.4 //y2=3.33
r317 (  41 44 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=7.4 //y=1.74 //x2=7.4 //y2=3.33
r318 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.655 //x2=7.4 //y2=1.74
r319 (  39 40 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.655 //x2=7.045 //y2=1.655
r320 (  38 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.005 //y=5.2 //x2=6.92 //y2=5.2
r321 (  37 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.2 //x2=7.4 //y2=5.115
r322 (  37 38 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.2 //x2=7.005 //y2=5.2
r323 (  33 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.96 //y=1.57 //x2=7.045 //y2=1.655
r324 (  33 113 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=6.96 //y=1.57 //x2=6.96 //y2=1
r325 (  27 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.92 //y=5.285 //x2=6.92 //y2=5.2
r326 (  27 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.92 //y=5.285 //x2=6.92 //y2=5.725
r327 (  25 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.835 //y=5.2 //x2=6.92 //y2=5.2
r328 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.835 //y=5.2 //x2=6.125 //y2=5.2
r329 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.04 //y=5.285 //x2=6.125 //y2=5.2
r330 (  19 115 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.04 //y=5.285 //x2=6.04 //y2=5.725
r331 (  17 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r332 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.33 //x2=3.33 //y2=4.7
r333 (  12 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r334 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.33
r335 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.25 //y=3.33 //x2=9.25 //y2=3.33
r336 (  8 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=7.4 \
 //y=3.33 //x2=7.4 //y2=3.33
r337 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.33 //x2=3.33 //y2=3.33
r338 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.515 //y=3.33 //x2=7.4 //y2=3.33
r339 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.135 //y=3.33 //x2=9.25 //y2=3.33
r340 (  3 4 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=9.135 //y=3.33 //x2=7.515 //y2=3.33
r341 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.445 //y=3.33 //x2=3.33 //y2=3.33
r342 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=3.33 //x2=7.4 //y2=3.33
r343 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=3.33 //x2=3.445 //y2=3.33
ends PM_DFFX1\%noxref_3

subckt PM_DFFX1\%noxref_4 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 \
 52 54 57 58 68 71 73 74 )
c150 ( 74 0 ) capacitor c=0.0220291f //x=10.105 //y=5.02
c151 ( 73 0 ) capacitor c=0.0217503f //x=9.225 //y=5.02
c152 ( 71 0 ) capacitor c=0.00866655f //x=10.1 //y=0.905
c153 ( 68 0 ) capacitor c=0.0588816f //x=12.58 //y=4.7
c154 ( 58 0 ) capacitor c=0.0318948f //x=12.915 //y=1.21
c155 ( 57 0 ) capacitor c=0.0187384f //x=12.915 //y=0.865
c156 ( 54 0 ) capacitor c=0.0141798f //x=12.76 //y=1.365
c157 ( 52 0 ) capacitor c=0.0149844f //x=12.76 //y=0.71
c158 ( 48 0 ) capacitor c=0.0853292f //x=12.385 //y=1.915
c159 ( 47 0 ) capacitor c=0.0229722f //x=12.385 //y=1.52
c160 ( 46 0 ) capacitor c=0.0234352f //x=12.385 //y=1.21
c161 ( 45 0 ) capacitor c=0.0199343f //x=12.385 //y=0.865
c162 ( 44 0 ) capacitor c=0.110275f //x=12.92 //y=6.02
c163 ( 43 0 ) capacitor c=0.154305f //x=12.48 //y=6.02
c164 ( 41 0 ) capacitor c=0.00211606f //x=10.25 //y=5.2
c165 ( 34 0 ) capacitor c=0.0911845f //x=12.58 //y=2.08
c166 ( 32 0 ) capacitor c=0.108686f //x=10.73 //y=3.33
c167 ( 28 0 ) capacitor c=0.00525782f //x=10.375 //y=1.655
c168 ( 27 0 ) capacitor c=0.0139525f //x=10.645 //y=1.655
c169 ( 25 0 ) capacitor c=0.0137516f //x=10.645 //y=5.2
c170 ( 14 0 ) capacitor c=0.00251459f //x=9.455 //y=5.2
c171 ( 13 0 ) capacitor c=0.0143643f //x=10.165 //y=5.2
c172 ( 2 0 ) capacitor c=0.00861293f //x=10.845 //y=3.33
c173 ( 1 0 ) capacitor c=0.067133f //x=12.465 //y=3.33
r174 (  66 68 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=12.48 //y=4.7 //x2=12.58 //y2=4.7
r175 (  59 68 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=12.92 //y=4.865 //x2=12.58 //y2=4.7
r176 (  58 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.915 //y=1.21 //x2=12.875 //y2=1.365
r177 (  57 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.915 //y=0.865 //x2=12.875 //y2=0.71
r178 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.915 //y=0.865 //x2=12.915 //y2=1.21
r179 (  55 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.54 //y=1.365 //x2=12.425 //y2=1.365
r180 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.76 //y=1.365 //x2=12.875 //y2=1.365
r181 (  53 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.54 //y=0.71 //x2=12.425 //y2=0.71
r182 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.76 //y=0.71 //x2=12.875 //y2=0.71
r183 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=12.76 //y=0.71 //x2=12.54 //y2=0.71
r184 (  49 66 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=12.48 //y=4.865 //x2=12.48 //y2=4.7
r185 (  48 63 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.915 //x2=12.58 //y2=2.08
r186 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.52 //x2=12.425 //y2=1.365
r187 (  47 48 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.52 //x2=12.385 //y2=1.915
r188 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.21 //x2=12.425 //y2=1.365
r189 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.385 //y=0.865 //x2=12.425 //y2=0.71
r190 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.385 //y=0.865 //x2=12.385 //y2=1.21
r191 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.92 //y=6.02 //x2=12.92 //y2=4.865
r192 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.48 //y=6.02 //x2=12.48 //y2=4.865
r193 (  42 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.65 //y=1.365 //x2=12.76 //y2=1.365
r194 (  42 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.65 //y=1.365 //x2=12.54 //y2=1.365
r195 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.58 //y=4.7 //x2=12.58 //y2=4.7
r196 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=12.58 //y=3.33 //x2=12.58 //y2=4.7
r197 (  34 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.58 //y=2.08 //x2=12.58 //y2=2.08
r198 (  34 37 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=12.58 //y=2.08 //x2=12.58 //y2=3.33
r199 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=10.73 //y=5.115 //x2=10.73 //y2=3.33
r200 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=10.73 //y=1.74 //x2=10.73 //y2=3.33
r201 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.645 //y=1.655 //x2=10.73 //y2=1.74
r202 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=10.645 //y=1.655 //x2=10.375 //y2=1.655
r203 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.335 //y=5.2 //x2=10.25 //y2=5.2
r204 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.645 //y=5.2 //x2=10.73 //y2=5.115
r205 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=10.645 //y=5.2 //x2=10.335 //y2=5.2
r206 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.29 //y=1.57 //x2=10.375 //y2=1.655
r207 (  21 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=10.29 //y=1.57 //x2=10.29 //y2=1
r208 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.25 //y=5.285 //x2=10.25 //y2=5.2
r209 (  15 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=10.25 //y=5.285 //x2=10.25 //y2=5.725
r210 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.165 //y=5.2 //x2=10.25 //y2=5.2
r211 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.165 //y=5.2 //x2=9.455 //y2=5.2
r212 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.37 //y=5.285 //x2=9.455 //y2=5.2
r213 (  7 73 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=9.37 //y=5.285 //x2=9.37 //y2=5.725
r214 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.58 //y=3.33 //x2=12.58 //y2=3.33
r215 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=3.33 //x2=10.73 //y2=3.33
r216 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.845 //y=3.33 //x2=10.73 //y2=3.33
r217 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.465 //y=3.33 //x2=12.58 //y2=3.33
r218 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=12.465 //y=3.33 //x2=10.845 //y2=3.33
ends PM_DFFX1\%noxref_4

subckt PM_DFFX1\%CLK ( 1 2 7 8 9 10 11 12 13 14 15 16 17 19 31 33 43 44 45 46 \
 47 48 49 50 51 53 59 60 61 62 63 68 69 70 75 77 79 85 86 90 99 100 103 )
c205 ( 103 0 ) capacitor c=0.0331838f //x=13.35 //y=4.7
c206 ( 100 0 ) capacitor c=0.0279499f //x=13.32 //y=1.915
c207 ( 99 0 ) capacitor c=0.0437302f //x=13.32 //y=2.08
c208 ( 90 0 ) capacitor c=0.0334842f //x=2.22 //y=4.7
c209 ( 86 0 ) capacitor c=0.0429696f //x=13.885 //y=1.25
c210 ( 85 0 ) capacitor c=0.0192208f //x=13.885 //y=0.905
c211 ( 79 0 ) capacitor c=0.0158629f //x=13.73 //y=1.405
c212 ( 77 0 ) capacitor c=0.0157803f //x=13.73 //y=0.75
c213 ( 75 0 ) capacitor c=0.0299681f //x=13.725 //y=4.79
c214 ( 70 0 ) capacitor c=0.0205163f //x=13.355 //y=1.56
c215 ( 69 0 ) capacitor c=0.0168481f //x=13.355 //y=1.25
c216 ( 68 0 ) capacitor c=0.0174783f //x=13.355 //y=0.905
c217 ( 63 0 ) capacitor c=0.0245352f //x=2.555 //y=4.79
c218 ( 62 0 ) capacitor c=0.0850619f //x=2.31 //y=1.915
c219 ( 61 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c220 ( 60 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c221 ( 59 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c222 ( 53 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c223 ( 51 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c224 ( 50 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c225 ( 49 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c226 ( 48 0 ) capacitor c=0.15358f //x=13.8 //y=6.02
c227 ( 47 0 ) capacitor c=0.110281f //x=13.36 //y=6.02
c228 ( 46 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c229 ( 45 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c230 ( 33 0 ) capacitor c=0.0746615f //x=13.32 //y=2.08
c231 ( 31 0 ) capacitor c=0.00369614f //x=13.32 //y=4.535
c232 ( 19 0 ) capacitor c=0.100158f //x=2.22 //y=2.08
c233 ( 2 0 ) capacitor c=0.0154455f //x=2.335 //y=4.44
c234 ( 1 0 ) capacitor c=0.25713f //x=13.205 //y=4.44
r235 (  105 106 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=13.35 //y=4.79 //x2=13.35 //y2=4.865
r236 (  103 105 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=13.35 //y=4.7 //x2=13.35 //y2=4.79
r237 (  99 100 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=13.32 //y=2.08 //x2=13.32 //y2=1.915
r238 (  92 93 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r239 (  90 92 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r240 (  86 110 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.885 //y=1.25 //x2=13.845 //y2=1.405
r241 (  85 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.885 //y=0.905 //x2=13.845 //y2=0.75
r242 (  85 86 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.885 //y=0.905 //x2=13.885 //y2=1.25
r243 (  80 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.51 //y=1.405 //x2=13.395 //y2=1.405
r244 (  79 110 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.73 //y=1.405 //x2=13.845 //y2=1.405
r245 (  78 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.51 //y=0.75 //x2=13.395 //y2=0.75
r246 (  77 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.73 //y=0.75 //x2=13.845 //y2=0.75
r247 (  77 78 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=13.73 //y=0.75 //x2=13.51 //y2=0.75
r248 (  76 105 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=13.485 //y=4.79 //x2=13.35 //y2=4.79
r249 (  75 82 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=13.725 //y=4.79 //x2=13.8 //y2=4.865
r250 (  75 76 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=13.725 //y=4.79 //x2=13.485 //y2=4.79
r251 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.355 //y=1.56 //x2=13.395 //y2=1.405
r252 (  70 100 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=13.355 //y=1.56 //x2=13.355 //y2=1.915
r253 (  69 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.355 //y=1.25 //x2=13.395 //y2=1.405
r254 (  68 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.355 //y=0.905 //x2=13.395 //y2=0.75
r255 (  68 69 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.355 //y=0.905 //x2=13.355 //y2=1.25
r256 (  64 92 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r257 (  63 65 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r258 (  63 64 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r259 (  62 97 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r260 (  61 95 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r261 (  61 62 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r262 (  60 95 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r263 (  59 94 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r264 (  59 60 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r265 (  54 88 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r266 (  53 95 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r267 (  52 87 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r268 (  51 94 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r269 (  51 52 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r270 (  50 88 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r271 (  49 87 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r272 (  49 50 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r273 (  48 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.8 //y=6.02 //x2=13.8 //y2=4.865
r274 (  47 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.36 //y=6.02 //x2=13.36 //y2=4.865
r275 (  46 65 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r276 (  45 93 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r277 (  44 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.62 //y=1.405 //x2=13.73 //y2=1.405
r278 (  44 80 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.62 //y=1.405 //x2=13.51 //y2=1.405
r279 (  43 53 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r280 (  43 54 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r281 (  42 103 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=13.35 //y=4.7 //x2=13.35 //y2=4.7
r282 (  33 99 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=13.32 //y=2.08 //x2=13.32 //y2=2.08
r283 (  31 42 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=13.32 //y=4.535 //x2=13.335 //y2=4.7
r284 (  29 90 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r285 (  19 97 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r286 (  17 31 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=13.32 //y=4.44 //x2=13.32 //y2=4.535
r287 (  16 17 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=13.32 //y=3.33 //x2=13.32 //y2=4.44
r288 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=13.32 //y=2.96 //x2=13.32 //y2=3.33
r289 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=13.32 //y=2.59 //x2=13.32 //y2=2.96
r290 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=13.32 //y=2.22 //x2=13.32 //y2=2.59
r291 (  13 33 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=13.32 //y=2.22 //x2=13.32 //y2=2.08
r292 (  12 29 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=2.22 //y=4.44 //x2=2.22 //y2=4.7
r293 (  11 12 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.7 //x2=2.22 //y2=4.44
r294 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.33 //x2=2.22 //y2=3.7
r295 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.96 //x2=2.22 //y2=3.33
r296 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.22 //y=2.59 //x2=2.22 //y2=2.96
r297 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.22 //y=2.22 //x2=2.22 //y2=2.59
r298 (  7 19 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.22 //x2=2.22 //y2=2.08
r299 (  6 17 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=13.32 //y=4.44 //x2=13.32 //y2=4.44
r300 (  4 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.22 //y=4.44 //x2=2.22 //y2=4.44
r301 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.335 //y=4.44 //x2=2.22 //y2=4.44
r302 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.205 //y=4.44 //x2=13.32 //y2=4.44
r303 (  1 2 ) resistor r=10.3721 //w=0.131 //l=10.87 //layer=m1 \
 //thickness=0.36 //x=13.205 //y=4.44 //x2=2.335 //y2=4.44
ends PM_DFFX1\%CLK

subckt PM_DFFX1\%noxref_6 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 63 64 65 \
 66 67 68 69 70 71 72 76 78 81 82 86 87 88 89 93 95 98 99 109 118 121 123 124 \
 125 )
c253 ( 125 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c254 ( 124 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c255 ( 123 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c256 ( 121 0 ) capacitor c=0.00872971f //x=3.395 //y=0.915
c257 ( 118 0 ) capacitor c=0.0593152f //x=15.91 //y=4.7
c258 ( 109 0 ) capacitor c=0.0588816f //x=5.92 //y=4.7
c259 ( 99 0 ) capacitor c=0.0318948f //x=16.245 //y=1.21
c260 ( 98 0 ) capacitor c=0.0187384f //x=16.245 //y=0.865
c261 ( 95 0 ) capacitor c=0.0141798f //x=16.09 //y=1.365
c262 ( 93 0 ) capacitor c=0.0149844f //x=16.09 //y=0.71
c263 ( 89 0 ) capacitor c=0.0860049f //x=15.715 //y=1.915
c264 ( 88 0 ) capacitor c=0.0229722f //x=15.715 //y=1.52
c265 ( 87 0 ) capacitor c=0.0234352f //x=15.715 //y=1.21
c266 ( 86 0 ) capacitor c=0.0199343f //x=15.715 //y=0.865
c267 ( 82 0 ) capacitor c=0.0318948f //x=6.255 //y=1.21
c268 ( 81 0 ) capacitor c=0.0187384f //x=6.255 //y=0.865
c269 ( 78 0 ) capacitor c=0.0141798f //x=6.1 //y=1.365
c270 ( 76 0 ) capacitor c=0.0149844f //x=6.1 //y=0.71
c271 ( 72 0 ) capacitor c=0.0860049f //x=5.725 //y=1.915
c272 ( 71 0 ) capacitor c=0.0229722f //x=5.725 //y=1.52
c273 ( 70 0 ) capacitor c=0.0234352f //x=5.725 //y=1.21
c274 ( 69 0 ) capacitor c=0.0199343f //x=5.725 //y=0.865
c275 ( 68 0 ) capacitor c=0.110275f //x=16.25 //y=6.02
c276 ( 67 0 ) capacitor c=0.154305f //x=15.81 //y=6.02
c277 ( 66 0 ) capacitor c=0.110275f //x=6.26 //y=6.02
c278 ( 65 0 ) capacitor c=0.154305f //x=5.82 //y=6.02
c279 ( 62 0 ) capacitor c=0.00106608f //x=3.29 //y=5.155
c280 ( 61 0 ) capacitor c=0.00207162f //x=2.41 //y=5.155
c281 ( 54 0 ) capacitor c=0.096094f //x=15.91 //y=2.08
c282 ( 46 0 ) capacitor c=0.0913801f //x=5.92 //y=2.08
c283 ( 44 0 ) capacitor c=0.109654f //x=4.07 //y=3.7
c284 ( 40 0 ) capacitor c=0.00493499f //x=3.67 //y=1.665
c285 ( 39 0 ) capacitor c=0.0154052f //x=3.985 //y=1.665
c286 ( 33 0 ) capacitor c=0.0284982f //x=3.985 //y=5.155
c287 ( 25 0 ) capacitor c=0.0176448f //x=3.205 //y=5.155
c288 ( 18 0 ) capacitor c=0.00351598f //x=1.615 //y=5.155
c289 ( 17 0 ) capacitor c=0.015419f //x=2.325 //y=5.155
c290 ( 4 0 ) capacitor c=0.00424317f //x=6.035 //y=3.7
c291 ( 3 0 ) capacitor c=0.215066f //x=15.795 //y=3.7
c292 ( 2 0 ) capacitor c=0.0125346f //x=4.185 //y=3.7
c293 ( 1 0 ) capacitor c=0.0285004f //x=5.805 //y=3.7
r294 (  116 118 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=15.81 //y=4.7 //x2=15.91 //y2=4.7
r295 (  107 109 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=5.82 //y=4.7 //x2=5.92 //y2=4.7
r296 (  100 118 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=16.25 //y=4.865 //x2=15.91 //y2=4.7
r297 (  99 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.245 //y=1.21 //x2=16.205 //y2=1.365
r298 (  98 119 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.245 //y=0.865 //x2=16.205 //y2=0.71
r299 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.245 //y=0.865 //x2=16.245 //y2=1.21
r300 (  96 115 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.87 //y=1.365 //x2=15.755 //y2=1.365
r301 (  95 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.09 //y=1.365 //x2=16.205 //y2=1.365
r302 (  94 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.87 //y=0.71 //x2=15.755 //y2=0.71
r303 (  93 119 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.09 //y=0.71 //x2=16.205 //y2=0.71
r304 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=16.09 //y=0.71 //x2=15.87 //y2=0.71
r305 (  90 116 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=15.81 //y=4.865 //x2=15.81 //y2=4.7
r306 (  89 113 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.915 //x2=15.91 //y2=2.08
r307 (  88 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.52 //x2=15.755 //y2=1.365
r308 (  88 89 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.52 //x2=15.715 //y2=1.915
r309 (  87 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.21 //x2=15.755 //y2=1.365
r310 (  86 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.715 //y=0.865 //x2=15.755 //y2=0.71
r311 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.715 //y=0.865 //x2=15.715 //y2=1.21
r312 (  83 109 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=6.26 //y=4.865 //x2=5.92 //y2=4.7
r313 (  82 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.255 //y=1.21 //x2=6.215 //y2=1.365
r314 (  81 110 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.255 //y=0.865 //x2=6.215 //y2=0.71
r315 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.255 //y=0.865 //x2=6.255 //y2=1.21
r316 (  79 106 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.88 //y=1.365 //x2=5.765 //y2=1.365
r317 (  78 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.1 //y=1.365 //x2=6.215 //y2=1.365
r318 (  77 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.88 //y=0.71 //x2=5.765 //y2=0.71
r319 (  76 110 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.1 //y=0.71 //x2=6.215 //y2=0.71
r320 (  76 77 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.1 //y=0.71 //x2=5.88 //y2=0.71
r321 (  73 107 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=5.82 //y=4.865 //x2=5.82 //y2=4.7
r322 (  72 104 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.915 //x2=5.92 //y2=2.08
r323 (  71 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.52 //x2=5.765 //y2=1.365
r324 (  71 72 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.52 //x2=5.725 //y2=1.915
r325 (  70 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.21 //x2=5.765 //y2=1.365
r326 (  69 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.725 //y=0.865 //x2=5.765 //y2=0.71
r327 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.725 //y=0.865 //x2=5.725 //y2=1.21
r328 (  68 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.25 //y=6.02 //x2=16.25 //y2=4.865
r329 (  67 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.81 //y=6.02 //x2=15.81 //y2=4.865
r330 (  66 83 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.26 //y=6.02 //x2=6.26 //y2=4.865
r331 (  65 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.82 //y=6.02 //x2=5.82 //y2=4.865
r332 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.98 //y=1.365 //x2=16.09 //y2=1.365
r333 (  64 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.98 //y=1.365 //x2=15.87 //y2=1.365
r334 (  63 78 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.99 //y=1.365 //x2=6.1 //y2=1.365
r335 (  63 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.99 //y=1.365 //x2=5.88 //y2=1.365
r336 (  59 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.91 //y=4.7 //x2=15.91 //y2=4.7
r337 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=15.91 //y=3.7 //x2=15.91 //y2=4.7
r338 (  54 113 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.91 //y=2.08 //x2=15.91 //y2=2.08
r339 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=15.91 //y=2.08 //x2=15.91 //y2=3.7
r340 (  51 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.7 //x2=5.92 //y2=4.7
r341 (  49 51 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=4.7
r342 (  46 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r343 (  46 49 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=3.7
r344 (  42 44 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=3.7
r345 (  41 44 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=3.7
r346 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r347 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r348 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r349 (  35 121 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r350 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r351 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r352 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r353 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r354 (  27 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r355 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r356 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r357 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r358 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r359 (  19 124 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r360 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r361 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r362 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r363 (  11 123 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r364 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.91 //y=3.7 //x2=15.91 //y2=3.7
r365 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=3.7
r366 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.7 //x2=4.07 //y2=3.7
r367 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=3.7 //x2=5.92 //y2=3.7
r368 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=3.7 //x2=15.91 //y2=3.7
r369 (  3 4 ) resistor r=9.31298 //w=0.131 //l=9.76 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=3.7 //x2=6.035 //y2=3.7
r370 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=3.7 //x2=4.07 //y2=3.7
r371 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.805 //y=3.7 //x2=5.92 //y2=3.7
r372 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.805 //y=3.7 //x2=4.185 //y2=3.7
ends PM_DFFX1\%noxref_6

subckt PM_DFFX1\%QN ( 1 2 7 8 9 10 11 12 13 14 15 16 17 24 25 36 38 39 50 61 \
 62 63 64 65 66 67 68 72 74 77 78 88 91 93 94 )
c147 ( 94 0 ) capacitor c=0.0220291f //x=16.765 //y=5.02
c148 ( 93 0 ) capacitor c=0.0217503f //x=15.885 //y=5.02
c149 ( 91 0 ) capacitor c=0.00866655f //x=16.76 //y=0.905
c150 ( 88 0 ) capacitor c=0.0593152f //x=19.24 //y=4.7
c151 ( 78 0 ) capacitor c=0.0318948f //x=19.575 //y=1.21
c152 ( 77 0 ) capacitor c=0.0187384f //x=19.575 //y=0.865
c153 ( 74 0 ) capacitor c=0.0141798f //x=19.42 //y=1.365
c154 ( 72 0 ) capacitor c=0.0149844f //x=19.42 //y=0.71
c155 ( 68 0 ) capacitor c=0.0853292f //x=19.045 //y=1.915
c156 ( 67 0 ) capacitor c=0.0229722f //x=19.045 //y=1.52
c157 ( 66 0 ) capacitor c=0.0234352f //x=19.045 //y=1.21
c158 ( 65 0 ) capacitor c=0.0199343f //x=19.045 //y=0.865
c159 ( 64 0 ) capacitor c=0.110275f //x=19.58 //y=6.02
c160 ( 63 0 ) capacitor c=0.154305f //x=19.14 //y=6.02
c161 ( 61 0 ) capacitor c=0.0023043f //x=16.91 //y=5.2
c162 ( 50 0 ) capacitor c=0.0933903f //x=19.24 //y=2.08
c163 ( 39 0 ) capacitor c=0.00525782f //x=17.035 //y=1.655
c164 ( 38 0 ) capacitor c=0.0139525f //x=17.305 //y=1.655
c165 ( 36 0 ) capacitor c=0.0140456f //x=17.305 //y=5.2
c166 ( 25 0 ) capacitor c=0.00265417f //x=16.115 //y=5.2
c167 ( 24 0 ) capacitor c=0.0149565f //x=16.825 //y=5.2
c168 ( 7 0 ) capacitor c=0.110168f //x=17.39 //y=2.22
c169 ( 2 0 ) capacitor c=0.0139448f //x=17.505 //y=3.33
c170 ( 1 0 ) capacitor c=0.0671025f //x=19.125 //y=3.33
r171 (  86 88 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=19.14 //y=4.7 //x2=19.24 //y2=4.7
r172 (  79 88 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=19.58 //y=4.865 //x2=19.24 //y2=4.7
r173 (  78 90 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.575 //y=1.21 //x2=19.535 //y2=1.365
r174 (  77 89 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.575 //y=0.865 //x2=19.535 //y2=0.71
r175 (  77 78 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.575 //y=0.865 //x2=19.575 //y2=1.21
r176 (  75 85 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.2 //y=1.365 //x2=19.085 //y2=1.365
r177 (  74 90 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.42 //y=1.365 //x2=19.535 //y2=1.365
r178 (  73 84 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.2 //y=0.71 //x2=19.085 //y2=0.71
r179 (  72 89 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.42 //y=0.71 //x2=19.535 //y2=0.71
r180 (  72 73 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=19.42 //y=0.71 //x2=19.2 //y2=0.71
r181 (  69 86 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=19.14 //y=4.865 //x2=19.14 //y2=4.7
r182 (  68 83 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.915 //x2=19.24 //y2=2.08
r183 (  67 85 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.52 //x2=19.085 //y2=1.365
r184 (  67 68 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.52 //x2=19.045 //y2=1.915
r185 (  66 85 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.21 //x2=19.085 //y2=1.365
r186 (  65 84 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.045 //y=0.865 //x2=19.085 //y2=0.71
r187 (  65 66 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.045 //y=0.865 //x2=19.045 //y2=1.21
r188 (  64 79 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.58 //y=6.02 //x2=19.58 //y2=4.865
r189 (  63 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.14 //y=6.02 //x2=19.14 //y2=4.865
r190 (  62 74 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=19.31 //y=1.365 //x2=19.42 //y2=1.365
r191 (  62 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=19.31 //y=1.365 //x2=19.2 //y2=1.365
r192 (  59 88 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.24 //y=4.7 //x2=19.24 //y2=4.7
r193 (  50 83 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.24 //y=2.08 //x2=19.24 //y2=2.08
r194 (  38 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.305 //y=1.655 //x2=17.39 //y2=1.74
r195 (  38 39 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=17.305 //y=1.655 //x2=17.035 //y2=1.655
r196 (  37 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.995 //y=5.2 //x2=16.91 //y2=5.2
r197 (  36 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.305 //y=5.2 //x2=17.39 //y2=5.115
r198 (  36 37 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=17.305 //y=5.2 //x2=16.995 //y2=5.2
r199 (  32 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.95 //y=1.57 //x2=17.035 //y2=1.655
r200 (  32 91 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.95 //y=1.57 //x2=16.95 //y2=1
r201 (  26 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.91 //y=5.285 //x2=16.91 //y2=5.2
r202 (  26 94 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=16.91 //y=5.285 //x2=16.91 //y2=5.725
r203 (  24 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.825 //y=5.2 //x2=16.91 //y2=5.2
r204 (  24 25 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.825 //y=5.2 //x2=16.115 //y2=5.2
r205 (  18 25 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.03 //y=5.285 //x2=16.115 //y2=5.2
r206 (  18 93 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=16.03 //y=5.285 //x2=16.03 //y2=5.725
r207 (  17 59 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=19.24 //y=4.44 //x2=19.24 //y2=4.7
r208 (  16 17 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=19.24 //y=3.33 //x2=19.24 //y2=4.44
r209 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.24 //y=2.96 //x2=19.24 //y2=3.33
r210 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.24 //y=2.59 //x2=19.24 //y2=2.96
r211 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.24 //y=2.22 //x2=19.24 //y2=2.59
r212 (  13 50 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=19.24 //y=2.22 //x2=19.24 //y2=2.08
r213 (  12 41 ) resistor r=20.877 //w=0.187 //l=0.305 //layer=li \
 //thickness=0.1 //x=17.39 //y=4.81 //x2=17.39 //y2=5.115
r214 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=17.39 //y=4.44 //x2=17.39 //y2=4.81
r215 (  10 11 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.39 //y=3.33 //x2=17.39 //y2=4.44
r216 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=17.39 //y=2.96 //x2=17.39 //y2=3.33
r217 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=17.39 //y=2.59 //x2=17.39 //y2=2.96
r218 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=17.39 //y=2.22 //x2=17.39 //y2=2.59
r219 (  7 40 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li \
 //thickness=0.1 //x=17.39 //y=2.22 //x2=17.39 //y2=1.74
r220 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.24 //y=3.33 //x2=19.24 //y2=3.33
r221 (  4 10 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.39 //y=3.33 //x2=17.39 //y2=3.33
r222 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.505 //y=3.33 //x2=17.39 //y2=3.33
r223 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.125 //y=3.33 //x2=19.24 //y2=3.33
r224 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=19.125 //y=3.33 //x2=17.505 //y2=3.33
ends PM_DFFX1\%QN

subckt PM_DFFX1\%noxref_8 ( 1 2 3 4 5 6 16 23 25 35 36 47 49 50 54 55 57 63 66 \
 67 68 69 70 71 72 73 74 75 76 77 78 79 81 87 88 89 90 94 95 96 101 103 105 \
 111 112 113 114 115 120 122 124 130 131 141 142 145 154 155 158 166 168 169 )
c358 ( 169 0 ) capacitor c=0.0220291f //x=13.435 //y=5.02
c359 ( 168 0 ) capacitor c=0.0217503f //x=12.555 //y=5.02
c360 ( 166 0 ) capacitor c=0.00866655f //x=13.43 //y=0.905
c361 ( 158 0 ) capacitor c=0.0331844f //x=20.01 //y=4.7
c362 ( 155 0 ) capacitor c=0.0279499f //x=19.98 //y=1.915
c363 ( 154 0 ) capacitor c=0.0437302f //x=19.98 //y=2.08
c364 ( 145 0 ) capacitor c=0.0331095f //x=10.02 //y=4.7
c365 ( 142 0 ) capacitor c=0.0279499f //x=9.99 //y=1.915
c366 ( 141 0 ) capacitor c=0.0437302f //x=9.99 //y=2.08
c367 ( 131 0 ) capacitor c=0.0429696f //x=20.545 //y=1.25
c368 ( 130 0 ) capacitor c=0.0192208f //x=20.545 //y=0.905
c369 ( 124 0 ) capacitor c=0.0158629f //x=20.39 //y=1.405
c370 ( 122 0 ) capacitor c=0.0157803f //x=20.39 //y=0.75
c371 ( 120 0 ) capacitor c=0.0306375f //x=20.385 //y=4.79
c372 ( 115 0 ) capacitor c=0.0205163f //x=20.015 //y=1.56
c373 ( 114 0 ) capacitor c=0.0168481f //x=20.015 //y=1.25
c374 ( 113 0 ) capacitor c=0.0174783f //x=20.015 //y=0.905
c375 ( 112 0 ) capacitor c=0.0429696f //x=10.555 //y=1.25
c376 ( 111 0 ) capacitor c=0.0192208f //x=10.555 //y=0.905
c377 ( 105 0 ) capacitor c=0.0158629f //x=10.4 //y=1.405
c378 ( 103 0 ) capacitor c=0.0157803f //x=10.4 //y=0.75
c379 ( 101 0 ) capacitor c=0.0295235f //x=10.395 //y=4.79
c380 ( 96 0 ) capacitor c=0.0205163f //x=10.025 //y=1.56
c381 ( 95 0 ) capacitor c=0.0168481f //x=10.025 //y=1.25
c382 ( 94 0 ) capacitor c=0.0174783f //x=10.025 //y=0.905
c383 ( 90 0 ) capacitor c=0.0559896f //x=1.385 //y=4.79
c384 ( 89 0 ) capacitor c=0.0298189f //x=1.675 //y=4.79
c385 ( 88 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c386 ( 87 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c387 ( 81 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c388 ( 79 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c389 ( 78 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c390 ( 77 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c391 ( 76 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c392 ( 75 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c393 ( 74 0 ) capacitor c=0.15358f //x=20.46 //y=6.02
c394 ( 73 0 ) capacitor c=0.110281f //x=20.02 //y=6.02
c395 ( 72 0 ) capacitor c=0.15358f //x=10.47 //y=6.02
c396 ( 71 0 ) capacitor c=0.110281f //x=10.03 //y=6.02
c397 ( 70 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c398 ( 69 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c399 ( 63 0 ) capacitor c=0.0023043f //x=13.58 //y=5.2
c400 ( 57 0 ) capacitor c=0.0765697f //x=19.98 //y=2.08
c401 ( 55 0 ) capacitor c=0.00453889f //x=19.98 //y=4.535
c402 ( 54 0 ) capacitor c=0.111691f //x=14.06 //y=4.07
c403 ( 50 0 ) capacitor c=0.00525782f //x=13.705 //y=1.655
c404 ( 49 0 ) capacitor c=0.0140405f //x=13.975 //y=1.655
c405 ( 47 0 ) capacitor c=0.0140413f //x=13.975 //y=5.2
c406 ( 36 0 ) capacitor c=0.00251459f //x=12.785 //y=5.2
c407 ( 35 0 ) capacitor c=0.0143105f //x=13.495 //y=5.2
c408 ( 25 0 ) capacitor c=0.0739568f //x=9.99 //y=2.08
c409 ( 23 0 ) capacitor c=0.00453889f //x=9.99 //y=4.535
c410 ( 16 0 ) capacitor c=0.124161f //x=1.11 //y=2.08
c411 ( 6 0 ) capacitor c=0.00579061f //x=14.175 //y=4.07
c412 ( 5 0 ) capacitor c=0.172193f //x=19.865 //y=4.07
c413 ( 4 0 ) capacitor c=0.00412846f //x=10.105 //y=4.07
c414 ( 3 0 ) capacitor c=0.0575172f //x=13.945 //y=4.07
c415 ( 2 0 ) capacitor c=0.0160818f //x=1.225 //y=4.07
c416 ( 1 0 ) capacitor c=0.163284f //x=9.875 //y=4.07
r417 (  160 161 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=20.01 //y=4.79 //x2=20.01 //y2=4.865
r418 (  158 160 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=20.01 //y=4.7 //x2=20.01 //y2=4.79
r419 (  154 155 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=19.98 //y=2.08 //x2=19.98 //y2=1.915
r420 (  147 148 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=10.02 //y=4.79 //x2=10.02 //y2=4.865
r421 (  145 147 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=10.02 //y=4.7 //x2=10.02 //y2=4.79
r422 (  141 142 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=9.99 //y=2.08 //x2=9.99 //y2=1.915
r423 (  131 165 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.545 //y=1.25 //x2=20.505 //y2=1.405
r424 (  130 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.545 //y=0.905 //x2=20.505 //y2=0.75
r425 (  130 131 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.545 //y=0.905 //x2=20.545 //y2=1.25
r426 (  125 163 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.17 //y=1.405 //x2=20.055 //y2=1.405
r427 (  124 165 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.39 //y=1.405 //x2=20.505 //y2=1.405
r428 (  123 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.17 //y=0.75 //x2=20.055 //y2=0.75
r429 (  122 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.39 //y=0.75 //x2=20.505 //y2=0.75
r430 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.39 //y=0.75 //x2=20.17 //y2=0.75
r431 (  121 160 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=20.145 //y=4.79 //x2=20.01 //y2=4.79
r432 (  120 127 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.385 //y=4.79 //x2=20.46 //y2=4.865
r433 (  120 121 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=20.385 //y=4.79 //x2=20.145 //y2=4.79
r434 (  115 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.015 //y=1.56 //x2=20.055 //y2=1.405
r435 (  115 155 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=20.015 //y=1.56 //x2=20.015 //y2=1.915
r436 (  114 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.015 //y=1.25 //x2=20.055 //y2=1.405
r437 (  113 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.015 //y=0.905 //x2=20.055 //y2=0.75
r438 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.015 //y=0.905 //x2=20.015 //y2=1.25
r439 (  112 152 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.555 //y=1.25 //x2=10.515 //y2=1.405
r440 (  111 151 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.555 //y=0.905 //x2=10.515 //y2=0.75
r441 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.555 //y=0.905 //x2=10.555 //y2=1.25
r442 (  106 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.18 //y=1.405 //x2=10.065 //y2=1.405
r443 (  105 152 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.4 //y=1.405 //x2=10.515 //y2=1.405
r444 (  104 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.18 //y=0.75 //x2=10.065 //y2=0.75
r445 (  103 151 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.4 //y=0.75 //x2=10.515 //y2=0.75
r446 (  103 104 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.4 //y=0.75 //x2=10.18 //y2=0.75
r447 (  102 147 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=10.155 //y=4.79 //x2=10.02 //y2=4.79
r448 (  101 108 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.395 //y=4.79 //x2=10.47 //y2=4.865
r449 (  101 102 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=10.395 //y=4.79 //x2=10.155 //y2=4.79
r450 (  96 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.025 //y=1.56 //x2=10.065 //y2=1.405
r451 (  96 142 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=10.025 //y=1.56 //x2=10.025 //y2=1.915
r452 (  95 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.025 //y=1.25 //x2=10.065 //y2=1.405
r453 (  94 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.025 //y=0.905 //x2=10.065 //y2=0.75
r454 (  94 95 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.025 //y=0.905 //x2=10.025 //y2=1.25
r455 (  89 91 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r456 (  89 90 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r457 (  88 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r458 (  87 138 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r459 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r460 (  84 90 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r461 (  84 137 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r462 (  82 133 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r463 (  81 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r464 (  80 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r465 (  79 138 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r466 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r467 (  78 135 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r468 (  77 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r469 (  77 78 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r470 (  76 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r471 (  75 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r472 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r473 (  74 127 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.46 //y=6.02 //x2=20.46 //y2=4.865
r474 (  73 161 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.02 //y=6.02 //x2=20.02 //y2=4.865
r475 (  72 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.47 //y=6.02 //x2=10.47 //y2=4.865
r476 (  71 148 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.03 //y=6.02 //x2=10.03 //y2=4.865
r477 (  70 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r478 (  69 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r479 (  68 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.28 //y=1.405 //x2=20.39 //y2=1.405
r480 (  68 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.28 //y=1.405 //x2=20.17 //y2=1.405
r481 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.29 //y=1.405 //x2=10.4 //y2=1.405
r482 (  67 106 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.29 //y=1.405 //x2=10.18 //y2=1.405
r483 (  66 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r484 (  66 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r485 (  65 158 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.01 //y=4.7 //x2=20.01 //y2=4.7
r486 (  62 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.02 //y=4.7 //x2=10.02 //y2=4.7
r487 (  57 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.98 //y=2.08 //x2=19.98 //y2=2.08
r488 (  57 60 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.08 //x2=19.98 //y2=4.07
r489 (  55 65 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=19.98 //y=4.535 //x2=19.995 //y2=4.7
r490 (  55 60 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=19.98 //y=4.535 //x2=19.98 //y2=4.07
r491 (  52 54 ) resistor r=71.5294 //w=0.187 //l=1.045 //layer=li \
 //thickness=0.1 //x=14.06 //y=5.115 //x2=14.06 //y2=4.07
r492 (  51 54 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=14.06 //y=1.74 //x2=14.06 //y2=4.07
r493 (  49 51 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.975 //y=1.655 //x2=14.06 //y2=1.74
r494 (  49 50 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=13.975 //y=1.655 //x2=13.705 //y2=1.655
r495 (  48 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.665 //y=5.2 //x2=13.58 //y2=5.2
r496 (  47 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.975 //y=5.2 //x2=14.06 //y2=5.115
r497 (  47 48 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=13.975 //y=5.2 //x2=13.665 //y2=5.2
r498 (  43 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.62 //y=1.57 //x2=13.705 //y2=1.655
r499 (  43 166 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=13.62 //y=1.57 //x2=13.62 //y2=1
r500 (  37 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.58 //y=5.285 //x2=13.58 //y2=5.2
r501 (  37 169 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=13.58 //y=5.285 //x2=13.58 //y2=5.725
r502 (  35 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.495 //y=5.2 //x2=13.58 //y2=5.2
r503 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=13.495 //y=5.2 //x2=12.785 //y2=5.2
r504 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.7 //y=5.285 //x2=12.785 //y2=5.2
r505 (  29 168 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=12.7 //y=5.285 //x2=12.7 //y2=5.725
r506 (  25 141 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.99 //y=2.08 //x2=9.99 //y2=2.08
r507 (  25 28 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=9.99 //y=2.08 //x2=9.99 //y2=4.07
r508 (  23 62 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=9.99 //y=4.535 //x2=10.005 //y2=4.7
r509 (  23 28 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=9.99 //y=4.535 //x2=9.99 //y2=4.07
r510 (  21 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r511 (  19 21 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.7
r512 (  16 135 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r513 (  16 19 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.08 //x2=1.11 //y2=4.07
r514 (  14 60 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.98 //y=4.07 //x2=19.98 //y2=4.07
r515 (  12 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=4.07 //x2=14.06 //y2=4.07
r516 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.99 //y=4.07 //x2=9.99 //y2=4.07
r517 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.07
r518 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.175 //y=4.07 //x2=14.06 //y2=4.07
r519 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=4.07 //x2=19.98 //y2=4.07
r520 (  5 6 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=4.07 //x2=14.175 //y2=4.07
r521 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.105 //y=4.07 //x2=9.99 //y2=4.07
r522 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=4.07 //x2=14.06 //y2=4.07
r523 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=4.07 //x2=10.105 //y2=4.07
r524 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=4.07 //x2=1.11 //y2=4.07
r525 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.875 //y=4.07 //x2=9.99 //y2=4.07
r526 (  1 2 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=9.875 //y=4.07 //x2=1.225 //y2=4.07
ends PM_DFFX1\%noxref_8

subckt PM_DFFX1\%Q ( 1 2 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 23 38 39 50 \
 52 53 67 68 69 70 71 72 73 78 80 82 88 89 91 92 95 103 105 106 )
c158 ( 106 0 ) capacitor c=0.0220291f //x=20.095 //y=5.02
c159 ( 105 0 ) capacitor c=0.0217503f //x=19.215 //y=5.02
c160 ( 103 0 ) capacitor c=0.0084702f //x=20.09 //y=0.905
c161 ( 95 0 ) capacitor c=0.0331552f //x=16.68 //y=4.7
c162 ( 92 0 ) capacitor c=0.0279499f //x=16.65 //y=1.915
c163 ( 91 0 ) capacitor c=0.0437302f //x=16.65 //y=2.08
c164 ( 89 0 ) capacitor c=0.0429696f //x=17.215 //y=1.25
c165 ( 88 0 ) capacitor c=0.0192208f //x=17.215 //y=0.905
c166 ( 82 0 ) capacitor c=0.0158629f //x=17.06 //y=1.405
c167 ( 80 0 ) capacitor c=0.0157803f //x=17.06 //y=0.75
c168 ( 78 0 ) capacitor c=0.0299681f //x=17.055 //y=4.79
c169 ( 73 0 ) capacitor c=0.0205163f //x=16.685 //y=1.56
c170 ( 72 0 ) capacitor c=0.0168481f //x=16.685 //y=1.25
c171 ( 71 0 ) capacitor c=0.0174783f //x=16.685 //y=0.905
c172 ( 70 0 ) capacitor c=0.15358f //x=17.13 //y=6.02
c173 ( 69 0 ) capacitor c=0.110281f //x=16.69 //y=6.02
c174 ( 67 0 ) capacitor c=0.0024826f //x=20.24 //y=5.2
c175 ( 53 0 ) capacitor c=0.00525782f //x=20.365 //y=1.655
c176 ( 52 0 ) capacitor c=0.0140375f //x=20.635 //y=1.655
c177 ( 50 0 ) capacitor c=0.0142748f //x=20.635 //y=5.2
c178 ( 39 0 ) capacitor c=0.00265417f //x=19.445 //y=5.2
c179 ( 38 0 ) capacitor c=0.0150828f //x=20.155 //y=5.2
c180 ( 23 0 ) capacitor c=0.0767118f //x=16.65 //y=2.08
c181 ( 21 0 ) capacitor c=0.00453889f //x=16.65 //y=4.535
c182 ( 13 0 ) capacitor c=0.128349f //x=20.72 //y=2.22
c183 ( 2 0 ) capacitor c=0.00699696f //x=16.765 //y=3.7
c184 ( 1 0 ) capacitor c=0.101946f //x=20.605 //y=3.7
r185 (  97 98 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=16.68 //y=4.79 //x2=16.68 //y2=4.865
r186 (  95 97 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=16.68 //y=4.7 //x2=16.68 //y2=4.79
r187 (  91 92 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=16.65 //y=2.08 //x2=16.65 //y2=1.915
r188 (  89 102 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.215 //y=1.25 //x2=17.175 //y2=1.405
r189 (  88 101 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.215 //y=0.905 //x2=17.175 //y2=0.75
r190 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.215 //y=0.905 //x2=17.215 //y2=1.25
r191 (  83 100 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.84 //y=1.405 //x2=16.725 //y2=1.405
r192 (  82 102 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.06 //y=1.405 //x2=17.175 //y2=1.405
r193 (  81 99 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.84 //y=0.75 //x2=16.725 //y2=0.75
r194 (  80 101 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.06 //y=0.75 //x2=17.175 //y2=0.75
r195 (  80 81 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.06 //y=0.75 //x2=16.84 //y2=0.75
r196 (  79 97 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=16.815 //y=4.79 //x2=16.68 //y2=4.79
r197 (  78 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=17.055 //y=4.79 //x2=17.13 //y2=4.865
r198 (  78 79 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=17.055 //y=4.79 //x2=16.815 //y2=4.79
r199 (  73 100 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.685 //y=1.56 //x2=16.725 //y2=1.405
r200 (  73 92 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=16.685 //y=1.56 //x2=16.685 //y2=1.915
r201 (  72 100 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.685 //y=1.25 //x2=16.725 //y2=1.405
r202 (  71 99 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.685 //y=0.905 //x2=16.725 //y2=0.75
r203 (  71 72 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.685 //y=0.905 //x2=16.685 //y2=1.25
r204 (  70 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.13 //y=6.02 //x2=17.13 //y2=4.865
r205 (  69 98 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.69 //y=6.02 //x2=16.69 //y2=4.865
r206 (  68 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.95 //y=1.405 //x2=17.06 //y2=1.405
r207 (  68 83 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.95 //y=1.405 //x2=16.84 //y2=1.405
r208 (  66 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.68 //y=4.7 //x2=16.68 //y2=4.7
r209 (  52 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.635 //y=1.655 //x2=20.72 //y2=1.74
r210 (  52 53 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=20.635 //y=1.655 //x2=20.365 //y2=1.655
r211 (  51 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.325 //y=5.2 //x2=20.24 //y2=5.2
r212 (  50 55 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.635 //y=5.2 //x2=20.72 //y2=5.115
r213 (  50 51 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=20.635 //y=5.2 //x2=20.325 //y2=5.2
r214 (  46 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.28 //y=1.57 //x2=20.365 //y2=1.655
r215 (  46 103 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=20.28 //y=1.57 //x2=20.28 //y2=1
r216 (  40 67 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.24 //y=5.285 //x2=20.24 //y2=5.2
r217 (  40 106 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=20.24 //y=5.285 //x2=20.24 //y2=5.725
r218 (  38 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.155 //y=5.2 //x2=20.24 //y2=5.2
r219 (  38 39 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=20.155 //y=5.2 //x2=19.445 //y2=5.2
r220 (  32 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.36 //y=5.285 //x2=19.445 //y2=5.2
r221 (  32 105 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=19.36 //y=5.285 //x2=19.36 //y2=5.725
r222 (  23 91 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=2.08 //x2=16.65 //y2=2.08
r223 (  21 66 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.535 //x2=16.665 //y2=4.7
r224 (  20 55 ) resistor r=20.877 //w=0.187 //l=0.305 //layer=li \
 //thickness=0.1 //x=20.72 //y=4.81 //x2=20.72 //y2=5.115
r225 (  19 20 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=20.72 //y=4.44 //x2=20.72 //y2=4.81
r226 (  18 19 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=20.72 //y=4.07 //x2=20.72 //y2=4.44
r227 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=20.72 //y=3.7 //x2=20.72 //y2=4.07
r228 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=20.72 //y=3.33 //x2=20.72 //y2=3.7
r229 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.96 //x2=20.72 //y2=3.33
r230 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.59 //x2=20.72 //y2=2.96
r231 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.22 //x2=20.72 //y2=2.59
r232 (  13 54 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.22 //x2=20.72 //y2=1.74
r233 (  12 21 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.44 //x2=16.65 //y2=4.535
r234 (  11 12 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=16.65 //y=3.7 //x2=16.65 //y2=4.44
r235 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=16.65 //y=3.33 //x2=16.65 //y2=3.7
r236 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.96 //x2=16.65 //y2=3.33
r237 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=16.65 //y=2.59 //x2=16.65 //y2=2.96
r238 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=16.65 //y=2.22 //x2=16.65 //y2=2.59
r239 (  7 23 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.22 //x2=16.65 //y2=2.08
r240 (  6 17 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.72 //y=3.7 //x2=20.72 //y2=3.7
r241 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=16.65 //y=3.7 //x2=16.65 //y2=3.7
r242 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.765 //y=3.7 //x2=16.65 //y2=3.7
r243 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=3.7 //x2=20.72 //y2=3.7
r244 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=3.7 //x2=16.765 //y2=3.7
ends PM_DFFX1\%Q

subckt PM_DFFX1\%noxref_10 ( 1 5 9 13 17 35 )
c47 ( 35 0 ) capacitor c=0.0703709f //x=0.455 //y=0.375
c48 ( 17 0 ) capacitor c=0.0221229f //x=2.445 //y=1.59
c49 ( 13 0 ) capacitor c=0.0156939f //x=2.445 //y=0.54
c50 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c51 ( 5 0 ) capacitor c=0.0206412f //x=1.475 //y=1.59
c52 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r53 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r54 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r55 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r56 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r57 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r58 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r59 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r60 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r61 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r62 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r63 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r64 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r65 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r66 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r67 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r68 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r69 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r70 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_DFFX1\%noxref_10

subckt PM_DFFX1\%noxref_11 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.043074f //x=2.965 //y=0.375
c54 ( 28 0 ) capacitor c=0.00465142f //x=1.86 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c57 ( 11 0 ) capacitor c=0.0149771f //x=3.985 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c59 ( 1 0 ) capacitor c=0.0253322f //x=3.015 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_DFFX1\%noxref_11

subckt PM_DFFX1\%D ( 1 2 3 4 6 13 14 15 16 17 18 23 25 27 33 34 36 37 40 )
c73 ( 40 0 ) capacitor c=0.0331095f //x=6.69 //y=4.7
c74 ( 37 0 ) capacitor c=0.0279499f //x=6.66 //y=1.915
c75 ( 36 0 ) capacitor c=0.0437302f //x=6.66 //y=2.08
c76 ( 34 0 ) capacitor c=0.0429696f //x=7.225 //y=1.25
c77 ( 33 0 ) capacitor c=0.0192208f //x=7.225 //y=0.905
c78 ( 27 0 ) capacitor c=0.0158629f //x=7.07 //y=1.405
c79 ( 25 0 ) capacitor c=0.0157803f //x=7.07 //y=0.75
c80 ( 23 0 ) capacitor c=0.0295235f //x=7.065 //y=4.79
c81 ( 18 0 ) capacitor c=0.0205163f //x=6.695 //y=1.56
c82 ( 17 0 ) capacitor c=0.0168481f //x=6.695 //y=1.25
c83 ( 16 0 ) capacitor c=0.0174783f //x=6.695 //y=0.905
c84 ( 15 0 ) capacitor c=0.15358f //x=7.14 //y=6.02
c85 ( 14 0 ) capacitor c=0.110281f //x=6.7 //y=6.02
c86 ( 6 0 ) capacitor c=0.0737925f //x=6.66 //y=2.08
c87 ( 4 0 ) capacitor c=0.00453889f //x=6.66 //y=4.535
r88 (  42 43 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=6.69 //y=4.79 //x2=6.69 //y2=4.865
r89 (  40 42 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=6.69 //y=4.7 //x2=6.69 //y2=4.79
r90 (  36 37 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.66 //y=2.08 //x2=6.66 //y2=1.915
r91 (  34 47 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.225 //y=1.25 //x2=7.185 //y2=1.405
r92 (  33 46 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.225 //y=0.905 //x2=7.185 //y2=0.75
r93 (  33 34 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.225 //y=0.905 //x2=7.225 //y2=1.25
r94 (  28 45 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.85 //y=1.405 //x2=6.735 //y2=1.405
r95 (  27 47 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.07 //y=1.405 //x2=7.185 //y2=1.405
r96 (  26 44 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.85 //y=0.75 //x2=6.735 //y2=0.75
r97 (  25 46 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.07 //y=0.75 //x2=7.185 //y2=0.75
r98 (  25 26 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.07 //y=0.75 //x2=6.85 //y2=0.75
r99 (  24 42 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=6.825 //y=4.79 //x2=6.69 //y2=4.79
r100 (  23 30 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.065 //y=4.79 //x2=7.14 //y2=4.865
r101 (  23 24 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=7.065 //y=4.79 //x2=6.825 //y2=4.79
r102 (  18 45 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.695 //y=1.56 //x2=6.735 //y2=1.405
r103 (  18 37 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=6.695 //y=1.56 //x2=6.695 //y2=1.915
r104 (  17 45 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.695 //y=1.25 //x2=6.735 //y2=1.405
r105 (  16 44 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.695 //y=0.905 //x2=6.735 //y2=0.75
r106 (  16 17 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.695 //y=0.905 //x2=6.695 //y2=1.25
r107 (  15 30 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.14 //y=6.02 //x2=7.14 //y2=4.865
r108 (  14 43 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.7 //y=6.02 //x2=6.7 //y2=4.865
r109 (  13 27 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.96 //y=1.405 //x2=7.07 //y2=1.405
r110 (  13 28 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.96 //y=1.405 //x2=6.85 //y2=1.405
r111 (  12 40 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.69 //y=4.7 //x2=6.69 //y2=4.7
r112 (  6 36 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.08 //x2=6.66 //y2=2.08
r113 (  4 12 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=6.66 //y=4.535 //x2=6.675 //y2=4.7
r114 (  3 4 ) resistor r=107.807 //w=0.187 //l=1.575 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.96 //x2=6.66 //y2=4.535
r115 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=6.66 //y=2.59 //x2=6.66 //y2=2.96
r116 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=6.66 //y=2.22 //x2=6.66 //y2=2.59
r117 (  1 6 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li //thickness=0.1 \
 //x=6.66 //y=2.22 //x2=6.66 //y2=2.08
ends PM_DFFX1\%D

subckt PM_DFFX1\%noxref_13 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0638069f //x=5.37 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=7.445 //y=0.615
c54 ( 13 0 ) capacitor c=0.0148848f //x=7.36 //y=0.53
c55 ( 10 0 ) capacitor c=0.00664066f //x=6.475 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=6.475 //y=0.615
c57 ( 5 0 ) capacitor c=0.0196287f //x=6.39 //y=1.58
c58 ( 1 0 ) capacitor c=0.00828748f //x=5.505 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.445 //y=0.615 //x2=7.445 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=7.445 //y=0.615 //x2=7.445 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.56 //y=0.53 //x2=6.475 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.56 //y=0.53 //x2=6.96 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.36 //y=0.53 //x2=7.445 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.36 //y=0.53 //x2=6.96 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.475 //y=1.495 //x2=6.475 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.475 //y=1.495 //x2=6.475 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.475 //y=0.615 //x2=6.475 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.475 //y=0.615 //x2=6.475 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.59 //y=1.58 //x2=5.505 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.59 //y=1.58 //x2=5.99 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.39 //y=1.58 //x2=6.475 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.39 //y=1.58 //x2=5.99 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.505 //y=1.495 //x2=5.505 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.505 //y=1.495 //x2=5.505 //y2=0.88
ends PM_DFFX1\%noxref_13

subckt PM_DFFX1\%noxref_14 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.0638071f //x=8.7 //y=0.365
c54 ( 17 0 ) capacitor c=0.00722223f //x=10.775 //y=0.615
c55 ( 13 0 ) capacitor c=0.0149613f //x=10.69 //y=0.53
c56 ( 10 0 ) capacitor c=0.00687696f //x=9.805 //y=1.495
c57 ( 9 0 ) capacitor c=0.006761f //x=9.805 //y=0.615
c58 ( 5 0 ) capacitor c=0.0201208f //x=9.72 //y=1.58
c59 ( 1 0 ) capacitor c=0.00828748f //x=8.835 //y=1.495
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=10.775 //y=0.615 //x2=10.775 //y2=0.49
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=10.775 //y=0.615 //x2=10.775 //y2=0.88
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.89 //y=0.53 //x2=9.805 //y2=0.49
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.89 //y=0.53 //x2=10.29 //y2=0.53
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.69 //y=0.53 //x2=10.775 //y2=0.49
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.69 //y=0.53 //x2=10.29 //y2=0.53
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.805 //y=1.495 //x2=9.805 //y2=1.62
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.805 //y=1.495 //x2=9.805 //y2=0.88
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.805 //y=0.615 //x2=9.805 //y2=0.49
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=9.805 //y=0.615 //x2=9.805 //y2=0.88
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.92 //y=1.58 //x2=8.835 //y2=1.62
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.92 //y=1.58 //x2=9.32 //y2=1.58
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.72 //y=1.58 //x2=9.805 //y2=1.62
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.72 //y=1.58 //x2=9.32 //y2=1.58
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.835 //y=1.495 //x2=8.835 //y2=1.62
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.835 //y=1.495 //x2=8.835 //y2=0.88
ends PM_DFFX1\%noxref_14

subckt PM_DFFX1\%noxref_15 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.0637486f //x=12.03 //y=0.365
c54 ( 17 0 ) capacitor c=0.00722223f //x=14.105 //y=0.615
c55 ( 13 0 ) capacitor c=0.0149666f //x=14.02 //y=0.53
c56 ( 10 0 ) capacitor c=0.00687696f //x=13.135 //y=1.495
c57 ( 9 0 ) capacitor c=0.006761f //x=13.135 //y=0.615
c58 ( 5 0 ) capacitor c=0.0201208f //x=13.05 //y=1.58
c59 ( 1 0 ) capacitor c=0.00828748f //x=12.165 //y=1.495
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.105 //y=0.615 //x2=14.105 //y2=0.49
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=14.105 //y=0.615 //x2=14.105 //y2=0.88
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.22 //y=0.53 //x2=13.135 //y2=0.49
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.22 //y=0.53 //x2=13.62 //y2=0.53
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.02 //y=0.53 //x2=14.105 //y2=0.49
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.02 //y=0.53 //x2=13.62 //y2=0.53
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=13.135 //y=1.495 //x2=13.135 //y2=1.62
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.135 //y=1.495 //x2=13.135 //y2=0.88
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=13.135 //y=0.615 //x2=13.135 //y2=0.49
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=13.135 //y=0.615 //x2=13.135 //y2=0.88
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.25 //y=1.58 //x2=12.165 //y2=1.62
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.25 //y=1.58 //x2=12.65 //y2=1.58
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.05 //y=1.58 //x2=13.135 //y2=1.62
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.05 //y=1.58 //x2=12.65 //y2=1.58
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=12.165 //y=1.495 //x2=12.165 //y2=1.62
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=12.165 //y=1.495 //x2=12.165 //y2=0.88
ends PM_DFFX1\%noxref_15

subckt PM_DFFX1\%noxref_16 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0638071f //x=15.36 //y=0.365
c55 ( 17 0 ) capacitor c=0.00722223f //x=17.435 //y=0.615
c56 ( 13 0 ) capacitor c=0.0150745f //x=17.35 //y=0.53
c57 ( 10 0 ) capacitor c=0.00705906f //x=16.465 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=16.465 //y=0.615
c59 ( 5 0 ) capacitor c=0.0207245f //x=16.38 //y=1.58
c60 ( 1 0 ) capacitor c=0.00856252f //x=15.495 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=17.435 //y=0.615 //x2=17.435 //y2=0.49
r62 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=17.435 //y=0.615 //x2=17.435 //y2=0.88
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.55 //y=0.53 //x2=16.465 //y2=0.49
r64 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.55 //y=0.53 //x2=16.95 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.35 //y=0.53 //x2=17.435 //y2=0.49
r66 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.35 //y=0.53 //x2=16.95 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=16.465 //y=1.495 //x2=16.465 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=16.465 //y=1.495 //x2=16.465 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=16.465 //y=0.615 //x2=16.465 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=16.465 //y=0.615 //x2=16.465 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.58 //y=1.58 //x2=15.495 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.58 //y=1.58 //x2=15.98 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.38 //y=1.58 //x2=16.465 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.38 //y=1.58 //x2=15.98 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.495 //y=1.495 //x2=15.495 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.495 //y=1.495 //x2=15.495 //y2=0.88
ends PM_DFFX1\%noxref_16

subckt PM_DFFX1\%noxref_17 ( 1 5 9 10 13 17 29 )
c50 ( 29 0 ) capacitor c=0.0637434f //x=18.69 //y=0.365
c51 ( 17 0 ) capacitor c=0.00722223f //x=20.765 //y=0.615
c52 ( 13 0 ) capacitor c=0.0149664f //x=20.68 //y=0.53
c53 ( 10 0 ) capacitor c=0.00687696f //x=19.795 //y=1.495
c54 ( 9 0 ) capacitor c=0.006761f //x=19.795 //y=0.615
c55 ( 5 0 ) capacitor c=0.0201208f //x=19.71 //y=1.58
c56 ( 1 0 ) capacitor c=0.00828748f //x=18.825 //y=1.495
r57 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=20.765 //y=0.615 //x2=20.765 //y2=0.49
r58 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.765 //y=0.615 //x2=20.765 //y2=0.88
r59 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.88 //y=0.53 //x2=19.795 //y2=0.49
r60 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.88 //y=0.53 //x2=20.28 //y2=0.53
r61 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.68 //y=0.53 //x2=20.765 //y2=0.49
r62 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.68 //y=0.53 //x2=20.28 //y2=0.53
r63 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=19.795 //y=1.495 //x2=19.795 //y2=1.62
r64 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=19.795 //y=1.495 //x2=19.795 //y2=0.88
r65 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=19.795 //y=0.615 //x2=19.795 //y2=0.49
r66 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=19.795 //y=0.615 //x2=19.795 //y2=0.88
r67 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.91 //y=1.58 //x2=18.825 //y2=1.62
r68 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.91 //y=1.58 //x2=19.31 //y2=1.58
r69 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.71 //y=1.58 //x2=19.795 //y2=1.62
r70 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.71 //y=1.58 //x2=19.31 //y2=1.58
r71 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=18.825 //y=1.495 //x2=18.825 //y2=1.62
r72 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=18.825 //y=1.495 //x2=18.825 //y2=0.88
ends PM_DFFX1\%noxref_17

