magic
tech sky130A
magscale 1 2
timestamp 1652450674
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 2277 945 2311 979
rect 131 871 165 905
rect 649 871 683 905
rect 797 871 831 905
rect 1463 871 1497 905
rect 2277 871 2311 905
rect 131 797 165 831
rect 649 797 683 831
rect 797 797 831 831
rect 1463 797 1497 831
rect 2277 797 2311 831
rect 131 723 165 757
rect 649 723 683 757
rect 797 723 831 757
rect 1463 723 1497 757
rect 2277 723 2311 757
rect 131 649 165 683
rect 1463 649 1497 683
rect 2277 649 2311 683
rect 131 575 165 609
rect 649 575 683 609
rect 797 575 831 609
rect 2277 575 2311 609
rect 131 501 165 535
rect 649 501 683 535
rect 797 501 831 535
rect 1463 501 1497 535
rect 2277 501 2311 535
rect 131 427 165 461
rect 649 427 683 461
rect 797 427 831 461
rect 1463 427 1497 461
rect 2277 427 2311 461
<< metal1 >>
rect -34 1446 2476 1514
rect -34 -34 2476 34
use mux2x1_pcell  mux2x1_pcell_0 pcells
timestamp 1652450488
transform 1 0 0 0 1 0
box -87 -34 2529 1550
<< labels >>
rlabel locali 2277 649 2311 683 1 Y
port 1 nsew signal output
rlabel locali 2277 723 2311 757 1 Y
port 1 nsew signal output
rlabel locali 2277 797 2311 831 1 Y
port 1 nsew signal output
rlabel locali 2277 871 2311 905 1 Y
port 1 nsew signal output
rlabel locali 2277 945 2311 979 1 Y
port 1 nsew signal output
rlabel locali 2277 575 2311 609 1 Y
port 1 nsew signal output
rlabel locali 2277 501 2311 535 1 Y
port 1 nsew signal output
rlabel locali 2277 427 2311 461 1 Y
port 1 nsew signal output
rlabel locali 797 723 831 757 1 A0
port 2 nsew signal input
rlabel locali 797 797 831 831 1 A0
port 2 nsew signal input
rlabel locali 797 871 831 905 1 A0
port 2 nsew signal input
rlabel locali 797 575 831 609 1 A0
port 2 nsew signal input
rlabel locali 797 501 831 535 1 A0
port 2 nsew signal input
rlabel locali 797 427 831 461 1 A0
port 2 nsew signal input
rlabel locali 1463 723 1497 757 1 A1
port 3 nsew signal input
rlabel locali 1463 649 1497 683 1 A1
port 3 nsew signal input
rlabel locali 1463 501 1497 535 1 A1
port 3 nsew signal input
rlabel locali 1463 427 1497 461 1 A1
port 3 nsew signal input
rlabel locali 1463 871 1497 905 1 A1
port 3 nsew signal input
rlabel locali 1463 797 1497 831 1 A1
port 3 nsew signal input
rlabel locali 131 575 165 609 1 S
port 4 nsew signal input
rlabel locali 131 649 165 683 1 S
port 4 nsew signal input
rlabel locali 131 723 165 757 1 S
port 4 nsew signal input
rlabel locali 131 797 165 831 1 S
port 4 nsew signal input
rlabel locali 131 871 165 905 1 S
port 4 nsew signal input
rlabel locali 131 501 165 535 1 S
port 4 nsew signal input
rlabel locali 131 427 165 461 1 S
port 4 nsew signal input
rlabel locali 649 871 683 905 1 S
port 4 nsew signal input
rlabel locali 649 797 683 831 1 S
port 4 nsew signal input
rlabel locali 649 723 683 757 1 S
port 4 nsew signal input
rlabel locali 649 575 683 609 1 S
port 4 nsew signal input
rlabel locali 649 501 683 535 1 S
port 4 nsew signal input
rlabel locali 649 427 683 461 1 S
port 4 nsew signal input
rlabel metal1 -34 1446 2476 1514 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 -34 -34 2476 34 1 GND
port 6 nsew ground bidirectional abutment


<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 2442 1480
string LEFsymmetry X Y R90
<< end >>
