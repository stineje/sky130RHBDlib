* SPICE3 file created from DLATCHN.ext - technology: sky130A

.subckt DLATCHN Q D GATE_N VDD GND
M1000 a_3461_1051.t3 Q.t4 VDD.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_n259_209.t1 GATE_N.t0 VDD.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t19 a_n259_209.t3 a_661_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t11 a_1295_209.t3 a_2795_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD.t4 a_1771_1050.t5 a_2405_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_185_209.t1 D.t1 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1295_209.t1 a_661_1050.t5 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t3 D.t2 a_1771_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_661_1050.t0 a_n259_209.t4 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1771_1050.t0 D.t3 VDD.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 Q.t1 a_3007_411.t4 a_2795_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_3461_1051.t1 a_2405_209.t3 a_3007_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 GND a_n259_209.t7 a_1666_101.t0 nshort w=-1.605u l=1.765u
+  ad=8.7946p pd=61.42u as=0p ps=0u
M1013 a_661_1050.t4 a_185_209.t4 VDD.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1771_1050.t4 a_n259_209.t6 VDD.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_2795_1051.t1 a_1295_209.t4 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VDD.t12 Q.t6 a_3461_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VDD.t1 GATE_N.t1 a_n259_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_2405_209.t0 a_1771_1050.t6 VDD.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 Q a_1295_209.t5 GND.t0 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.15u as=0p ps=0u
M1020 Q a_3007_411.t5 GND.t4 nshort w=-1.83u l=2.06u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t15 a_185_209.t5 a_661_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t6 a_n259_209.t8 a_1771_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VDD.t0 D.t4 a_185_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VDD.t14 a_661_1050.t7 a_1295_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_3007_411.t0 a_2405_209.t5 a_3461_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 GND a_185_209.t3 a_556_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_2795_1051.t3 a_3007_411.t6 Q.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 D GATE_N 0.01fF
C1 Q VDD 0.33fF
C2 VDD GATE_N 0.12fF
C3 D VDD 0.19fF
R0 Q.n0 Q.t4 486.819
R1 Q.n0 Q.t6 384.527
R2 Q.n1 Q.t5 250.501
R3 Q.n11 Q.n2 191.889
R4 Q.n11 Q.n10 135.634
R5 Q.n1 Q.n0 133.1
R6 Q.n10 Q.n9 118.016
R7 Q.n5 Q.n3 80.526
R8 Q.n12 Q.n1 77.315
R9 Q.n12 Q.n11 76
R10 Q.n10 Q.n5 48.405
R11 Q.n9 Q.n8 30
R12 Q.n5 Q.n4 30
R13 Q.n7 Q.n6 24.383
R14 Q.n9 Q.n7 23.684
R15 Q.n2 Q.t3 14.282
R16 Q.n2 Q.t1 14.282
R17 Q.n12 Q 0.046
R18 VDD.n253 VDD.n251 144.705
R19 VDD.n321 VDD.n319 144.705
R20 VDD.n382 VDD.n380 144.705
R21 VDD.n184 VDD.n182 144.705
R22 VDD.n407 VDD.n405 144.705
R23 VDD.n138 VDD.n136 144.705
R24 VDD.n80 VDD.n78 144.705
R25 VDD.n143 VDD.n142 77.792
R26 VDD.n153 VDD.n152 77.792
R27 VDD.n397 VDD.n396 77.792
R28 VDD.n386 VDD.n385 77.792
R29 VDD.n290 VDD.n289 77.792
R30 VDD.n280 VDD.n279 77.792
R31 VDD.n243 VDD.n242 77.792
R32 VDD.n232 VDD.n231 77.792
R33 VDD.n40 VDD.n39 76
R34 VDD.n47 VDD.n46 76
R35 VDD.n51 VDD.n50 76
R36 VDD.n55 VDD.n54 76
R37 VDD.n82 VDD.n81 76
R38 VDD.n86 VDD.n85 76
R39 VDD.n90 VDD.n89 76
R40 VDD.n94 VDD.n93 76
R41 VDD.n99 VDD.n98 76
R42 VDD.n106 VDD.n105 76
R43 VDD.n110 VDD.n109 76
R44 VDD.n114 VDD.n113 76
R45 VDD.n140 VDD.n139 76
R46 VDD.n146 VDD.n145 76
R47 VDD.n150 VDD.n149 76
R48 VDD.n156 VDD.n155 76
R49 VDD.n160 VDD.n159 76
R50 VDD.n186 VDD.n185 76
R51 VDD.n191 VDD.n190 76
R52 VDD.n196 VDD.n195 76
R53 VDD.n202 VDD.n201 76
R54 VDD.n207 VDD.n206 76
R55 VDD.n440 VDD.n439 76
R56 VDD.n435 VDD.n434 76
R57 VDD.n430 VDD.n429 76
R58 VDD.n404 VDD.n403 76
R59 VDD.n400 VDD.n399 76
R60 VDD.n394 VDD.n393 76
R61 VDD.n390 VDD.n389 76
R62 VDD.n384 VDD.n383 76
R63 VDD.n358 VDD.n357 76
R64 VDD.n354 VDD.n353 76
R65 VDD.n349 VDD.n348 76
R66 VDD.n344 VDD.n343 76
R67 VDD.n338 VDD.n337 76
R68 VDD.n333 VDD.n332 76
R69 VDD.n328 VDD.n327 76
R70 VDD.n323 VDD.n322 76
R71 VDD.n297 VDD.n296 76
R72 VDD.n293 VDD.n292 76
R73 VDD.n287 VDD.n286 76
R74 VDD.n283 VDD.n282 76
R75 VDD.n277 VDD.n276 76
R76 VDD.n250 VDD.n249 76
R77 VDD.n246 VDD.n245 76
R78 VDD.n240 VDD.n239 76
R79 VDD.n236 VDD.n235 76
R80 VDD.n230 VDD.n229 76
R81 VDD.n234 VDD.t16 55.106
R82 VDD.n241 VDD.t1 55.106
R83 VDD.n278 VDD.t5 55.106
R84 VDD.n288 VDD.t0 55.106
R85 VDD.n324 VDD.t17 55.106
R86 VDD.n388 VDD.t8 55.106
R87 VDD.n395 VDD.t14 55.106
R88 VDD.n431 VDD.t7 55.106
R89 VDD.n151 VDD.t10 55.106
R90 VDD.n141 VDD.t4 55.106
R91 VDD.n350 VDD.t19 55.106
R92 VDD.n189 VDD.t3 55.106
R93 VDD.n101 VDD.n100 41.183
R94 VDD.n42 VDD.n41 41.183
R95 VDD.n340 VDD.n339 40.824
R96 VDD.n200 VDD.n199 40.824
R97 VDD.n302 VDD.n301 36.774
R98 VDD.n363 VDD.n362 36.774
R99 VDD.n412 VDD.n411 36.774
R100 VDD.n165 VDD.n164 36.774
R101 VDD.n119 VDD.n118 36.774
R102 VDD.n60 VDD.n59 36.774
R103 VDD.n269 VDD.n268 36.774
R104 VDD.n193 VDD.n192 36.608
R105 VDD.n346 VDD.n345 36.608
R106 VDD.n34 VDD.n33 34.942
R107 VDD.n44 VDD.n43 32.032
R108 VDD.n103 VDD.n102 32.032
R109 VDD.n437 VDD.n436 32.032
R110 VDD.n330 VDD.n329 32.032
R111 VDD.n229 VDD.n226 21.841
R112 VDD.n23 VDD.n20 21.841
R113 VDD.n339 VDD.t18 14.282
R114 VDD.n339 VDD.t15 14.282
R115 VDD.n199 VDD.t9 14.282
R116 VDD.n199 VDD.t6 14.282
R117 VDD.n100 VDD.t2 14.282
R118 VDD.n100 VDD.t11 14.282
R119 VDD.n41 VDD.t13 14.282
R120 VDD.n41 VDD.t12 14.282
R121 VDD.n226 VDD.n209 14.167
R122 VDD.n209 VDD.n208 14.167
R123 VDD.n317 VDD.n299 14.167
R124 VDD.n299 VDD.n298 14.167
R125 VDD.n378 VDD.n360 14.167
R126 VDD.n360 VDD.n359 14.167
R127 VDD.n427 VDD.n409 14.167
R128 VDD.n409 VDD.n408 14.167
R129 VDD.n180 VDD.n162 14.167
R130 VDD.n162 VDD.n161 14.167
R131 VDD.n134 VDD.n116 14.167
R132 VDD.n116 VDD.n115 14.167
R133 VDD.n76 VDD.n57 14.167
R134 VDD.n57 VDD.n56 14.167
R135 VDD.n274 VDD.n255 14.167
R136 VDD.n255 VDD.n254 14.167
R137 VDD.n20 VDD.n19 14.167
R138 VDD.n19 VDD.n17 14.167
R139 VDD.n32 VDD.n29 14.167
R140 VDD.n29 VDD.n28 14.167
R141 VDD.n81 VDD.n77 14.167
R142 VDD.n139 VDD.n135 14.167
R143 VDD.n185 VDD.n181 14.167
R144 VDD.n429 VDD.n428 14.167
R145 VDD.n383 VDD.n379 14.167
R146 VDD.n322 VDD.n318 14.167
R147 VDD.n276 VDD.n275 14.167
R148 VDD.n23 VDD.n22 13.653
R149 VDD.n22 VDD.n21 13.653
R150 VDD.n32 VDD.n31 13.653
R151 VDD.n31 VDD.n30 13.653
R152 VDD.n29 VDD.n25 13.653
R153 VDD.n25 VDD.n24 13.653
R154 VDD.n28 VDD.n27 13.653
R155 VDD.n27 VDD.n26 13.653
R156 VDD.n39 VDD.n38 13.653
R157 VDD.n38 VDD.n37 13.653
R158 VDD.n46 VDD.n45 13.653
R159 VDD.n45 VDD.n44 13.653
R160 VDD.n50 VDD.n49 13.653
R161 VDD.n49 VDD.n48 13.653
R162 VDD.n54 VDD.n53 13.653
R163 VDD.n53 VDD.n52 13.653
R164 VDD.n81 VDD.n80 13.653
R165 VDD.n80 VDD.n79 13.653
R166 VDD.n85 VDD.n84 13.653
R167 VDD.n84 VDD.n83 13.653
R168 VDD.n89 VDD.n88 13.653
R169 VDD.n88 VDD.n87 13.653
R170 VDD.n93 VDD.n92 13.653
R171 VDD.n92 VDD.n91 13.653
R172 VDD.n98 VDD.n97 13.653
R173 VDD.n97 VDD.n96 13.653
R174 VDD.n105 VDD.n104 13.653
R175 VDD.n104 VDD.n103 13.653
R176 VDD.n109 VDD.n108 13.653
R177 VDD.n108 VDD.n107 13.653
R178 VDD.n113 VDD.n112 13.653
R179 VDD.n112 VDD.n111 13.653
R180 VDD.n139 VDD.n138 13.653
R181 VDD.n138 VDD.n137 13.653
R182 VDD.n145 VDD.n144 13.653
R183 VDD.n144 VDD.n143 13.653
R184 VDD.n149 VDD.n148 13.653
R185 VDD.n148 VDD.n147 13.653
R186 VDD.n155 VDD.n154 13.653
R187 VDD.n154 VDD.n153 13.653
R188 VDD.n159 VDD.n158 13.653
R189 VDD.n158 VDD.n157 13.653
R190 VDD.n185 VDD.n184 13.653
R191 VDD.n184 VDD.n183 13.653
R192 VDD.n190 VDD.n188 13.653
R193 VDD.n188 VDD.n187 13.653
R194 VDD.n195 VDD.n194 13.653
R195 VDD.n194 VDD.n193 13.653
R196 VDD.n201 VDD.n198 13.653
R197 VDD.n198 VDD.n197 13.653
R198 VDD.n206 VDD.n205 13.653
R199 VDD.n205 VDD.n204 13.653
R200 VDD.n439 VDD.n438 13.653
R201 VDD.n438 VDD.n437 13.653
R202 VDD.n434 VDD.n433 13.653
R203 VDD.n433 VDD.n432 13.653
R204 VDD.n429 VDD.n407 13.653
R205 VDD.n407 VDD.n406 13.653
R206 VDD.n403 VDD.n402 13.653
R207 VDD.n402 VDD.n401 13.653
R208 VDD.n399 VDD.n398 13.653
R209 VDD.n398 VDD.n397 13.653
R210 VDD.n393 VDD.n392 13.653
R211 VDD.n392 VDD.n391 13.653
R212 VDD.n389 VDD.n387 13.653
R213 VDD.n387 VDD.n386 13.653
R214 VDD.n383 VDD.n382 13.653
R215 VDD.n382 VDD.n381 13.653
R216 VDD.n357 VDD.n356 13.653
R217 VDD.n356 VDD.n355 13.653
R218 VDD.n353 VDD.n352 13.653
R219 VDD.n352 VDD.n351 13.653
R220 VDD.n348 VDD.n347 13.653
R221 VDD.n347 VDD.n346 13.653
R222 VDD.n343 VDD.n342 13.653
R223 VDD.n342 VDD.n341 13.653
R224 VDD.n337 VDD.n336 13.653
R225 VDD.n336 VDD.n335 13.653
R226 VDD.n332 VDD.n331 13.653
R227 VDD.n331 VDD.n330 13.653
R228 VDD.n327 VDD.n326 13.653
R229 VDD.n326 VDD.n325 13.653
R230 VDD.n322 VDD.n321 13.653
R231 VDD.n321 VDD.n320 13.653
R232 VDD.n296 VDD.n295 13.653
R233 VDD.n295 VDD.n294 13.653
R234 VDD.n292 VDD.n291 13.653
R235 VDD.n291 VDD.n290 13.653
R236 VDD.n286 VDD.n285 13.653
R237 VDD.n285 VDD.n284 13.653
R238 VDD.n282 VDD.n281 13.653
R239 VDD.n281 VDD.n280 13.653
R240 VDD.n276 VDD.n253 13.653
R241 VDD.n253 VDD.n252 13.653
R242 VDD.n249 VDD.n248 13.653
R243 VDD.n248 VDD.n247 13.653
R244 VDD.n245 VDD.n244 13.653
R245 VDD.n244 VDD.n243 13.653
R246 VDD.n239 VDD.n238 13.653
R247 VDD.n238 VDD.n237 13.653
R248 VDD.n235 VDD.n233 13.653
R249 VDD.n233 VDD.n232 13.653
R250 VDD.n229 VDD.n228 13.653
R251 VDD.n228 VDD.n227 13.653
R252 VDD.n4 VDD.n2 12.915
R253 VDD.n4 VDD.n3 12.66
R254 VDD.n13 VDD.n12 12.343
R255 VDD.n11 VDD.n10 12.343
R256 VDD.n8 VDD.n7 12.343
R257 VDD.n201 VDD.n200 8.658
R258 VDD.n343 VDD.n340 8.658
R259 VDD.n318 VDD.n317 7.674
R260 VDD.n379 VDD.n378 7.674
R261 VDD.n428 VDD.n427 7.674
R262 VDD.n181 VDD.n180 7.674
R263 VDD.n135 VDD.n134 7.674
R264 VDD.n77 VDD.n76 7.674
R265 VDD.n275 VDD.n274 7.674
R266 VDD.n71 VDD.n70 7.5
R267 VDD.n65 VDD.n64 7.5
R268 VDD.n67 VDD.n66 7.5
R269 VDD.n62 VDD.n61 7.5
R270 VDD.n76 VDD.n75 7.5
R271 VDD.n129 VDD.n128 7.5
R272 VDD.n123 VDD.n122 7.5
R273 VDD.n125 VDD.n124 7.5
R274 VDD.n131 VDD.n121 7.5
R275 VDD.n131 VDD.n119 7.5
R276 VDD.n134 VDD.n133 7.5
R277 VDD.n175 VDD.n174 7.5
R278 VDD.n169 VDD.n168 7.5
R279 VDD.n171 VDD.n170 7.5
R280 VDD.n177 VDD.n167 7.5
R281 VDD.n177 VDD.n165 7.5
R282 VDD.n180 VDD.n179 7.5
R283 VDD.n422 VDD.n421 7.5
R284 VDD.n416 VDD.n415 7.5
R285 VDD.n418 VDD.n417 7.5
R286 VDD.n424 VDD.n414 7.5
R287 VDD.n424 VDD.n412 7.5
R288 VDD.n427 VDD.n426 7.5
R289 VDD.n373 VDD.n372 7.5
R290 VDD.n367 VDD.n366 7.5
R291 VDD.n369 VDD.n368 7.5
R292 VDD.n375 VDD.n365 7.5
R293 VDD.n375 VDD.n363 7.5
R294 VDD.n378 VDD.n377 7.5
R295 VDD.n312 VDD.n311 7.5
R296 VDD.n306 VDD.n305 7.5
R297 VDD.n308 VDD.n307 7.5
R298 VDD.n314 VDD.n304 7.5
R299 VDD.n314 VDD.n302 7.5
R300 VDD.n317 VDD.n316 7.5
R301 VDD.n259 VDD.n258 7.5
R302 VDD.n262 VDD.n261 7.5
R303 VDD.n264 VDD.n263 7.5
R304 VDD.n267 VDD.n266 7.5
R305 VDD.n274 VDD.n273 7.5
R306 VDD.n221 VDD.n220 7.5
R307 VDD.n215 VDD.n214 7.5
R308 VDD.n217 VDD.n216 7.5
R309 VDD.n223 VDD.n213 7.5
R310 VDD.n223 VDD.n211 7.5
R311 VDD.n226 VDD.n225 7.5
R312 VDD.n20 VDD.n16 7.5
R313 VDD.n2 VDD.n1 7.5
R314 VDD.n7 VDD.n6 7.5
R315 VDD.n10 VDD.n9 7.5
R316 VDD.n19 VDD.n18 7.5
R317 VDD.n14 VDD.n0 7.5
R318 VDD.n63 VDD.n60 6.772
R319 VDD.n74 VDD.n58 6.772
R320 VDD.n72 VDD.n69 6.772
R321 VDD.n68 VDD.n65 6.772
R322 VDD.n132 VDD.n117 6.772
R323 VDD.n130 VDD.n127 6.772
R324 VDD.n126 VDD.n123 6.772
R325 VDD.n178 VDD.n163 6.772
R326 VDD.n176 VDD.n173 6.772
R327 VDD.n172 VDD.n169 6.772
R328 VDD.n425 VDD.n410 6.772
R329 VDD.n423 VDD.n420 6.772
R330 VDD.n419 VDD.n416 6.772
R331 VDD.n376 VDD.n361 6.772
R332 VDD.n374 VDD.n371 6.772
R333 VDD.n370 VDD.n367 6.772
R334 VDD.n315 VDD.n300 6.772
R335 VDD.n313 VDD.n310 6.772
R336 VDD.n309 VDD.n306 6.772
R337 VDD.n224 VDD.n210 6.772
R338 VDD.n222 VDD.n219 6.772
R339 VDD.n218 VDD.n215 6.772
R340 VDD.n63 VDD.n62 6.772
R341 VDD.n68 VDD.n67 6.772
R342 VDD.n72 VDD.n71 6.772
R343 VDD.n75 VDD.n74 6.772
R344 VDD.n126 VDD.n125 6.772
R345 VDD.n130 VDD.n129 6.772
R346 VDD.n133 VDD.n132 6.772
R347 VDD.n172 VDD.n171 6.772
R348 VDD.n176 VDD.n175 6.772
R349 VDD.n179 VDD.n178 6.772
R350 VDD.n419 VDD.n418 6.772
R351 VDD.n423 VDD.n422 6.772
R352 VDD.n426 VDD.n425 6.772
R353 VDD.n370 VDD.n369 6.772
R354 VDD.n374 VDD.n373 6.772
R355 VDD.n377 VDD.n376 6.772
R356 VDD.n309 VDD.n308 6.772
R357 VDD.n313 VDD.n312 6.772
R358 VDD.n316 VDD.n315 6.772
R359 VDD.n218 VDD.n217 6.772
R360 VDD.n222 VDD.n221 6.772
R361 VDD.n225 VDD.n224 6.772
R362 VDD.n273 VDD.n272 6.772
R363 VDD.n260 VDD.n257 6.772
R364 VDD.n265 VDD.n262 6.772
R365 VDD.n270 VDD.n267 6.772
R366 VDD.n270 VDD.n269 6.772
R367 VDD.n265 VDD.n264 6.772
R368 VDD.n260 VDD.n259 6.772
R369 VDD.n272 VDD.n256 6.772
R370 VDD.n33 VDD.n23 6.487
R371 VDD.n33 VDD.n32 6.475
R372 VDD.n16 VDD.n15 6.458
R373 VDD.n121 VDD.n120 6.202
R374 VDD.n167 VDD.n166 6.202
R375 VDD.n414 VDD.n413 6.202
R376 VDD.n365 VDD.n364 6.202
R377 VDD.n304 VDD.n303 6.202
R378 VDD.n213 VDD.n212 6.202
R379 VDD.n46 VDD.n42 5.903
R380 VDD.n105 VDD.n101 5.903
R381 VDD.n37 VDD.n36 4.576
R382 VDD.n96 VDD.n95 4.576
R383 VDD.n204 VDD.n203 4.576
R384 VDD.n335 VDD.n334 4.576
R385 VDD.n434 VDD.n431 2.754
R386 VDD.n327 VDD.n324 2.754
R387 VDD.n190 VDD.n189 2.361
R388 VDD.n353 VDD.n350 2.361
R389 VDD.n145 VDD.n141 1.967
R390 VDD.n155 VDD.n151 1.967
R391 VDD.n399 VDD.n395 1.967
R392 VDD.n389 VDD.n388 1.967
R393 VDD.n292 VDD.n288 1.967
R394 VDD.n282 VDD.n278 1.967
R395 VDD.n245 VDD.n241 1.967
R396 VDD.n235 VDD.n234 1.967
R397 VDD.n14 VDD.n5 1.329
R398 VDD.n14 VDD.n8 1.329
R399 VDD.n14 VDD.n11 1.329
R400 VDD.n14 VDD.n13 1.329
R401 VDD.n15 VDD.n14 0.696
R402 VDD.n14 VDD.n4 0.696
R403 VDD.n73 VDD.n72 0.365
R404 VDD.n73 VDD.n68 0.365
R405 VDD.n73 VDD.n63 0.365
R406 VDD.n74 VDD.n73 0.365
R407 VDD.n131 VDD.n130 0.365
R408 VDD.n131 VDD.n126 0.365
R409 VDD.n132 VDD.n131 0.365
R410 VDD.n177 VDD.n176 0.365
R411 VDD.n177 VDD.n172 0.365
R412 VDD.n178 VDD.n177 0.365
R413 VDD.n424 VDD.n423 0.365
R414 VDD.n424 VDD.n419 0.365
R415 VDD.n425 VDD.n424 0.365
R416 VDD.n375 VDD.n374 0.365
R417 VDD.n375 VDD.n370 0.365
R418 VDD.n376 VDD.n375 0.365
R419 VDD.n314 VDD.n313 0.365
R420 VDD.n314 VDD.n309 0.365
R421 VDD.n315 VDD.n314 0.365
R422 VDD.n223 VDD.n222 0.365
R423 VDD.n223 VDD.n218 0.365
R424 VDD.n224 VDD.n223 0.365
R425 VDD.n271 VDD.n270 0.365
R426 VDD.n271 VDD.n265 0.365
R427 VDD.n271 VDD.n260 0.365
R428 VDD.n272 VDD.n271 0.365
R429 VDD.n82 VDD.n55 0.29
R430 VDD.n140 VDD.n114 0.29
R431 VDD.n186 VDD.n160 0.29
R432 VDD.n430 VDD.n404 0.29
R433 VDD.n384 VDD.n358 0.29
R434 VDD.n323 VDD.n297 0.29
R435 VDD.n277 VDD.n250 0.29
R436 VDD.n230 VDD 0.207
R437 VDD.n40 VDD.n35 0.181
R438 VDD.n99 VDD.n94 0.181
R439 VDD.n207 VDD.n202 0.181
R440 VDD.n344 VDD.n338 0.181
R441 VDD.n150 VDD.n146 0.157
R442 VDD.n156 VDD.n150 0.157
R443 VDD.n400 VDD.n394 0.157
R444 VDD.n394 VDD.n390 0.157
R445 VDD.n293 VDD.n287 0.157
R446 VDD.n287 VDD.n283 0.157
R447 VDD.n246 VDD.n240 0.157
R448 VDD.n240 VDD.n236 0.157
R449 VDD.n35 VDD.n34 0.145
R450 VDD.n47 VDD.n40 0.145
R451 VDD.n51 VDD.n47 0.145
R452 VDD.n55 VDD.n51 0.145
R453 VDD.n86 VDD.n82 0.145
R454 VDD.n90 VDD.n86 0.145
R455 VDD.n94 VDD.n90 0.145
R456 VDD.n106 VDD.n99 0.145
R457 VDD.n110 VDD.n106 0.145
R458 VDD.n114 VDD.n110 0.145
R459 VDD.n146 VDD.n140 0.145
R460 VDD.n160 VDD.n156 0.145
R461 VDD.n191 VDD.n186 0.145
R462 VDD.n196 VDD.n191 0.145
R463 VDD.n202 VDD.n196 0.145
R464 VDD.n440 VDD.n435 0.145
R465 VDD.n435 VDD.n430 0.145
R466 VDD.n404 VDD.n400 0.145
R467 VDD.n390 VDD.n384 0.145
R468 VDD.n358 VDD.n354 0.145
R469 VDD.n354 VDD.n349 0.145
R470 VDD.n349 VDD.n344 0.145
R471 VDD.n338 VDD.n333 0.145
R472 VDD.n333 VDD.n328 0.145
R473 VDD.n328 VDD.n323 0.145
R474 VDD.n297 VDD.n293 0.145
R475 VDD.n283 VDD.n277 0.145
R476 VDD.n250 VDD.n246 0.145
R477 VDD.n236 VDD.n230 0.145
R478 VDD VDD.n207 0.133
R479 VDD VDD.n440 0.012
R480 a_3461_1051.t2 a_3461_1051.n0 101.66
R481 a_3461_1051.n0 a_3461_1051.t1 101.659
R482 a_3461_1051.n0 a_3461_1051.t0 14.294
R483 a_3461_1051.n0 a_3461_1051.t3 14.282
R484 D.n2 D.t4 512.525
R485 D.n0 D.t2 472.359
R486 D.n0 D.t3 384.527
R487 D.n2 D.t1 371.139
R488 D.n1 D.t5 267.725
R489 D.n3 D.t0 263.54
R490 D.n3 D.n2 120.094
R491 D.n1 D.n0 83.507
R492 D.n4 D.n1 82.484
R493 D.n4 D.n3 76
R494 D.n4 D 0.046
R495 GND.n43 GND.n41 219.745
R496 GND.n169 GND.n168 219.745
R497 GND.n204 GND.n202 219.745
R498 GND.n234 GND.n232 219.745
R499 GND.n267 GND.n265 219.745
R500 GND.n120 GND.n118 219.745
R501 GND.n87 GND.n86 219.745
R502 GND.n43 GND.n42 85.529
R503 GND.n169 GND.n167 85.529
R504 GND.n204 GND.n203 85.529
R505 GND.n234 GND.n233 85.529
R506 GND.n267 GND.n266 85.529
R507 GND.n120 GND.n119 85.529
R508 GND.n87 GND.n85 85.529
R509 GND.n275 GND.n274 84.842
R510 GND.n212 GND.n211 84.842
R511 GND.n8 GND.n1 76.145
R512 GND.n139 GND.n138 76
R513 GND.n8 GND.n7 76
R514 GND.n14 GND.n13 76
R515 GND.n17 GND.n16 76
R516 GND.n24 GND.n23 76
R517 GND.n30 GND.n29 76
R518 GND.n37 GND.n36 76
R519 GND.n40 GND.n39 76
R520 GND.n47 GND.n46 76
R521 GND.n54 GND.n53 76
R522 GND.n60 GND.n59 76
R523 GND.n63 GND.n62 76
R524 GND.n69 GND.n68 76
R525 GND.n74 GND.n73 76
R526 GND.n81 GND.n80 76
R527 GND.n84 GND.n83 76
R528 GND.n91 GND.n90 76
R529 GND.n99 GND.n98 76
R530 GND.n107 GND.n106 76
R531 GND.n114 GND.n113 76
R532 GND.n117 GND.n116 76
R533 GND.n124 GND.n123 76
R534 GND.n127 GND.n126 76
R535 GND.n130 GND.n129 76
R536 GND.n133 GND.n132 76
R537 GND.n136 GND.n135 76
R538 GND.n278 GND.n277 76
R539 GND.n273 GND.n272 76
R540 GND.n270 GND.n269 76
R541 GND.n263 GND.n262 76
R542 GND.n260 GND.n259 76
R543 GND.n252 GND.n251 76
R544 GND.n244 GND.n243 76
R545 GND.n237 GND.n236 76
R546 GND.n230 GND.n229 76
R547 GND.n227 GND.n226 76
R548 GND.n224 GND.n223 76
R549 GND.n221 GND.n220 76
R550 GND.n218 GND.n217 76
R551 GND.n215 GND.n214 76
R552 GND.n210 GND.n209 76
R553 GND.n207 GND.n206 76
R554 GND.n200 GND.n199 76
R555 GND.n197 GND.n196 76
R556 GND.n189 GND.n188 76
R557 GND.n181 GND.n180 76
R558 GND.n172 GND.n171 76
R559 GND.n165 GND.n164 76
R560 GND.n162 GND.n161 76
R561 GND.n154 GND.n153 76
R562 GND.n146 GND.n145 76
R563 GND.n33 GND.t8 39.412
R564 GND.n177 GND.t2 39.412
R565 GND.n95 GND.n94 35.01
R566 GND.n256 GND.n255 35.01
R567 GND.n193 GND.n192 35.01
R568 GND.n158 GND.n157 35.01
R569 GND.n93 GND.n92 29.127
R570 GND.n254 GND.n253 29.127
R571 GND.n156 GND.n155 29.127
R572 GND.n102 GND.t7 20.794
R573 GND.n247 GND.t1 20.794
R574 GND.n149 GND.t9 20.794
R575 GND.n27 GND.n26 19.735
R576 GND.n21 GND.n20 19.735
R577 GND.n12 GND.n11 19.735
R578 GND.n5 GND.n4 19.735
R579 GND.n35 GND.n34 19.735
R580 GND.n71 GND.n70 19.735
R581 GND.n66 GND.n65 19.735
R582 GND.n58 GND.n57 19.735
R583 GND.n51 GND.n50 19.735
R584 GND.n79 GND.n78 19.735
R585 GND.n96 GND.n95 19.735
R586 GND.n104 GND.n103 19.735
R587 GND.n112 GND.n111 19.735
R588 GND.n257 GND.n256 19.735
R589 GND.n249 GND.n248 19.735
R590 GND.n242 GND.n241 19.735
R591 GND.n194 GND.n193 19.735
R592 GND.n186 GND.n185 19.735
R593 GND.n179 GND.n178 19.735
R594 GND.n159 GND.n158 19.735
R595 GND.n151 GND.n150 19.735
R596 GND.n144 GND.n143 19.735
R597 GND.n11 GND.t6 19.724
R598 GND.n57 GND.t4 19.724
R599 GND.n70 GND.t0 19.724
R600 GND.n95 GND.n93 19.017
R601 GND.n256 GND.n254 19.017
R602 GND.n193 GND.n191 19.017
R603 GND.n158 GND.n156 19.017
R604 GND.n33 GND.n32 17.185
R605 GND.n177 GND.n176 17.185
R606 GND.n46 GND.n44 14.167
R607 GND.n90 GND.n88 14.167
R608 GND.n123 GND.n121 14.167
R609 GND.n269 GND.n268 14.167
R610 GND.n236 GND.n235 14.167
R611 GND.n206 GND.n205 14.167
R612 GND.n171 GND.n170 14.167
R613 GND.n19 GND.n18 13.654
R614 GND.n145 GND.n140 13.653
R615 GND.n153 GND.n152 13.653
R616 GND.n161 GND.n160 13.653
R617 GND.n164 GND.n163 13.653
R618 GND.n171 GND.n166 13.653
R619 GND.n180 GND.n173 13.653
R620 GND.n188 GND.n187 13.653
R621 GND.n196 GND.n195 13.653
R622 GND.n199 GND.n198 13.653
R623 GND.n206 GND.n201 13.653
R624 GND.n209 GND.n208 13.653
R625 GND.n214 GND.n213 13.653
R626 GND.n217 GND.n216 13.653
R627 GND.n220 GND.n219 13.653
R628 GND.n223 GND.n222 13.653
R629 GND.n226 GND.n225 13.653
R630 GND.n229 GND.n228 13.653
R631 GND.n236 GND.n231 13.653
R632 GND.n243 GND.n238 13.653
R633 GND.n251 GND.n250 13.653
R634 GND.n259 GND.n258 13.653
R635 GND.n262 GND.n261 13.653
R636 GND.n269 GND.n264 13.653
R637 GND.n272 GND.n271 13.653
R638 GND.n277 GND.n276 13.653
R639 GND.n135 GND.n134 13.653
R640 GND.n132 GND.n131 13.653
R641 GND.n129 GND.n128 13.653
R642 GND.n126 GND.n125 13.653
R643 GND.n123 GND.n122 13.653
R644 GND.n116 GND.n115 13.653
R645 GND.n113 GND.n108 13.653
R646 GND.n106 GND.n105 13.653
R647 GND.n98 GND.n97 13.653
R648 GND.n90 GND.n89 13.653
R649 GND.n83 GND.n82 13.653
R650 GND.n80 GND.n75 13.653
R651 GND.n73 GND.n72 13.653
R652 GND.n68 GND.n67 13.653
R653 GND.n62 GND.n61 13.653
R654 GND.n59 GND.n55 13.653
R655 GND.n53 GND.n52 13.653
R656 GND.n46 GND.n45 13.653
R657 GND.n39 GND.n38 13.653
R658 GND.n36 GND.n31 13.653
R659 GND.n29 GND.n28 13.653
R660 GND.n23 GND.n22 13.653
R661 GND.n16 GND.n15 13.653
R662 GND.n13 GND.n9 13.653
R663 GND.n7 GND.n6 13.653
R664 GND.n78 GND.n77 12.837
R665 GND.n111 GND.n110 12.837
R666 GND.n241 GND.n240 12.837
R667 GND.n143 GND.n142 12.837
R668 GND.n4 GND.n3 11.605
R669 GND.n50 GND.n49 11.605
R670 GND.n3 GND.n2 9.809
R671 GND.n49 GND.n48 9.809
R672 GND.n23 GND.n21 8.854
R673 GND.n68 GND.n66 8.854
R674 GND.n77 GND.n76 7.566
R675 GND.n110 GND.n109 7.566
R676 GND.n240 GND.n239 7.566
R677 GND.n142 GND.n141 7.566
R678 GND.n26 GND.n25 7.5
R679 GND.n191 GND.n190 7.5
R680 GND.n184 GND.n183 7.5
R681 GND.n44 GND.n43 7.312
R682 GND.n170 GND.n169 7.312
R683 GND.n205 GND.n204 7.312
R684 GND.n235 GND.n234 7.312
R685 GND.n268 GND.n267 7.312
R686 GND.n121 GND.n120 7.312
R687 GND.n88 GND.n87 7.312
R688 GND.t6 GND.n10 7.04
R689 GND.t4 GND.n56 7.04
R690 GND.n34 GND.n33 6.139
R691 GND.n178 GND.n177 6.139
R692 GND.n20 GND.n19 5.774
R693 GND.n65 GND.n64 5.774
R694 GND.n101 GND.n100 4.551
R695 GND.n246 GND.n245 4.551
R696 GND.n175 GND.n174 4.551
R697 GND.n148 GND.n147 4.551
R698 GND.n13 GND.n12 3.935
R699 GND.n29 GND.n27 3.935
R700 GND.n59 GND.n58 3.935
R701 GND.n73 GND.n71 3.935
R702 GND.n98 GND.n96 3.935
R703 GND.n277 GND.n275 3.935
R704 GND.n259 GND.n257 3.935
R705 GND.n214 GND.n212 3.935
R706 GND.n196 GND.n194 3.935
R707 GND.n161 GND.n159 3.935
R708 GND.n113 GND.n112 3.541
R709 GND.n243 GND.n242 3.541
R710 GND.n180 GND.n179 3.541
R711 GND.n145 GND.n144 3.541
R712 GND.t7 GND.n101 2.238
R713 GND.t1 GND.n246 2.238
R714 GND.t2 GND.n175 2.238
R715 GND.t9 GND.n148 2.238
R716 GND.n183 GND.n182 1.935
R717 GND.n7 GND.n5 0.983
R718 GND.n36 GND.n35 0.983
R719 GND.n53 GND.n51 0.983
R720 GND.n80 GND.n79 0.983
R721 GND.n1 GND.n0 0.596
R722 GND.n138 GND.n137 0.596
R723 GND.n103 GND.n102 0.358
R724 GND.n248 GND.n247 0.358
R725 GND.n185 GND.n184 0.358
R726 GND.n150 GND.n149 0.358
R727 GND.n47 GND.n40 0.29
R728 GND.n91 GND.n84 0.29
R729 GND.n124 GND.n117 0.29
R730 GND.n270 GND.n263 0.29
R731 GND.n237 GND.n230 0.29
R732 GND.n207 GND.n200 0.29
R733 GND.n172 GND.n165 0.29
R734 GND.n139 GND 0.207
R735 GND.n106 GND.n104 0.196
R736 GND.n251 GND.n249 0.196
R737 GND.n188 GND.n186 0.196
R738 GND.n153 GND.n151 0.196
R739 GND.n24 GND.n17 0.181
R740 GND.n69 GND.n63 0.181
R741 GND.n136 GND.n133 0.181
R742 GND.n221 GND.n218 0.181
R743 GND.n107 GND.n99 0.157
R744 GND.n114 GND.n107 0.157
R745 GND.n260 GND.n252 0.157
R746 GND.n252 GND.n244 0.157
R747 GND.n197 GND.n189 0.157
R748 GND.n189 GND.n181 0.157
R749 GND.n162 GND.n154 0.157
R750 GND.n154 GND.n146 0.157
R751 GND.n14 GND.n8 0.145
R752 GND.n17 GND.n14 0.145
R753 GND.n30 GND.n24 0.145
R754 GND.n37 GND.n30 0.145
R755 GND.n40 GND.n37 0.145
R756 GND.n54 GND.n47 0.145
R757 GND.n60 GND.n54 0.145
R758 GND.n63 GND.n60 0.145
R759 GND.n74 GND.n69 0.145
R760 GND.n81 GND.n74 0.145
R761 GND.n84 GND.n81 0.145
R762 GND.n99 GND.n91 0.145
R763 GND.n117 GND.n114 0.145
R764 GND.n127 GND.n124 0.145
R765 GND.n130 GND.n127 0.145
R766 GND.n133 GND.n130 0.145
R767 GND.n278 GND.n273 0.145
R768 GND.n273 GND.n270 0.145
R769 GND.n263 GND.n260 0.145
R770 GND.n244 GND.n237 0.145
R771 GND.n230 GND.n227 0.145
R772 GND.n227 GND.n224 0.145
R773 GND.n224 GND.n221 0.145
R774 GND.n218 GND.n215 0.145
R775 GND.n215 GND.n210 0.145
R776 GND.n210 GND.n207 0.145
R777 GND.n200 GND.n197 0.145
R778 GND.n181 GND.n172 0.145
R779 GND.n165 GND.n162 0.145
R780 GND.n146 GND.n139 0.145
R781 GND GND.n136 0.133
R782 GND GND.n278 0.012
R783 a_185_209.n0 a_185_209.t5 480.392
R784 a_185_209.n0 a_185_209.t4 403.272
R785 a_185_209.n1 a_185_209.t3 283.48
R786 a_185_209.n3 a_185_209.n2 227.307
R787 a_185_209.n4 a_185_209.n3 157.453
R788 a_185_209.n3 a_185_209.n1 153.315
R789 a_185_209.n1 a_185_209.n0 98.447
R790 a_185_209.n4 a_185_209.t0 14.282
R791 a_185_209.t1 a_185_209.n4 14.282
R792 a_556_101.t0 a_556_101.n1 34.62
R793 a_556_101.t0 a_556_101.n0 8.137
R794 a_556_101.t0 a_556_101.n2 4.69
R795 GATE_N.n0 GATE_N.t1 512.525
R796 GATE_N.n0 GATE_N.t0 371.139
R797 GATE_N.n1 GATE_N.n0 199.753
R798 GATE_N.n1 GATE_N.t2 183.881
R799 GATE_N.n2 GATE_N.n1 76
R800 GATE_N.n2 GATE_N 0.046
R801 a_n259_209.n0 a_n259_209.t8 480.392
R802 a_n259_209.n2 a_n259_209.t3 472.359
R803 a_n259_209.n0 a_n259_209.t6 403.272
R804 a_n259_209.n2 a_n259_209.t4 384.527
R805 a_n259_209.n1 a_n259_209.t7 230.374
R806 a_n259_209.n7 a_n259_209.n6 210.559
R807 a_n259_209.n3 a_n259_209.t5 188.066
R808 a_n259_209.n6 a_n259_209.n5 174.201
R809 a_n259_209.n3 a_n259_209.n2 163.166
R810 a_n259_209.n1 a_n259_209.n0 151.553
R811 a_n259_209.n4 a_n259_209.n1 79.491
R812 a_n259_209.n6 a_n259_209.n4 79.491
R813 a_n259_209.n4 a_n259_209.n3 76
R814 a_n259_209.n7 a_n259_209.t0 14.282
R815 a_n259_209.t1 a_n259_209.n7 14.282
R816 a_661_1050.n0 a_661_1050.t7 512.525
R817 a_661_1050.n0 a_661_1050.t5 371.139
R818 a_661_1050.n1 a_661_1050.t6 210.434
R819 a_661_1050.n3 a_661_1050.n2 205.778
R820 a_661_1050.n5 a_661_1050.n3 179.052
R821 a_661_1050.n1 a_661_1050.n0 173.2
R822 a_661_1050.n3 a_661_1050.n1 153.043
R823 a_661_1050.n5 a_661_1050.n4 76.002
R824 a_661_1050.n4 a_661_1050.t3 14.282
R825 a_661_1050.n4 a_661_1050.t4 14.282
R826 a_661_1050.t1 a_661_1050.n6 14.282
R827 a_661_1050.n6 a_661_1050.t0 14.282
R828 a_661_1050.n6 a_661_1050.n5 12.848
R829 a_1295_209.n0 a_1295_209.t4 486.819
R830 a_1295_209.n0 a_1295_209.t3 384.527
R831 a_1295_209.n1 a_1295_209.t5 277.054
R832 a_1295_209.n3 a_1295_209.n2 227.307
R833 a_1295_209.n4 a_1295_209.n3 157.453
R834 a_1295_209.n3 a_1295_209.n1 157.396
R835 a_1295_209.n1 a_1295_209.n0 106.547
R836 a_1295_209.n4 a_1295_209.t0 14.282
R837 a_1295_209.t1 a_1295_209.n4 14.282
R838 a_2795_1051.t2 a_2795_1051.n0 101.66
R839 a_2795_1051.n0 a_2795_1051.t3 101.659
R840 a_2795_1051.n0 a_2795_1051.t0 14.294
R841 a_2795_1051.n0 a_2795_1051.t1 14.282
R842 a_1771_1050.n0 a_1771_1050.t5 512.525
R843 a_1771_1050.n0 a_1771_1050.t6 371.139
R844 a_1771_1050.n1 a_1771_1050.t7 210.434
R845 a_1771_1050.n6 a_1771_1050.n5 184.039
R846 a_1771_1050.n8 a_1771_1050.n6 179.052
R847 a_1771_1050.n1 a_1771_1050.n0 173.2
R848 a_1771_1050.n6 a_1771_1050.n1 153.043
R849 a_1771_1050.n8 a_1771_1050.n7 76.002
R850 a_1771_1050.n5 a_1771_1050.n4 30
R851 a_1771_1050.n3 a_1771_1050.n2 24.383
R852 a_1771_1050.n5 a_1771_1050.n3 23.684
R853 a_1771_1050.n7 a_1771_1050.t3 14.282
R854 a_1771_1050.n7 a_1771_1050.t4 14.282
R855 a_1771_1050.t1 a_1771_1050.n9 14.282
R856 a_1771_1050.n9 a_1771_1050.t0 14.282
R857 a_1771_1050.n9 a_1771_1050.n8 12.848
R858 a_2405_209.n0 a_2405_209.t3 470.752
R859 a_2405_209.n0 a_2405_209.t5 384.527
R860 a_2405_209.n1 a_2405_209.t4 267.725
R861 a_2405_209.n3 a_2405_209.n2 253.86
R862 a_2405_209.n3 a_2405_209.n1 156.307
R863 a_2405_209.n4 a_2405_209.n3 130.9
R864 a_2405_209.n1 a_2405_209.n0 83.62
R865 a_2405_209.t1 a_2405_209.n4 14.282
R866 a_2405_209.n4 a_2405_209.t0 14.282
R867 a_3007_411.n0 a_3007_411.t6 470.752
R868 a_3007_411.n0 a_3007_411.t4 384.527
R869 a_3007_411.n1 a_3007_411.t5 241.172
R870 a_3007_411.n8 a_3007_411.n7 165.335
R871 a_3007_411.n7 a_3007_411.n6 162.187
R872 a_3007_411.n7 a_3007_411.n1 154.947
R873 a_3007_411.n6 a_3007_411.n5 133.539
R874 a_3007_411.n1 a_3007_411.n0 110.173
R875 a_3007_411.n6 a_3007_411.n2 70.262
R876 a_3007_411.n5 a_3007_411.n4 22.578
R877 a_3007_411.t1 a_3007_411.n8 14.282
R878 a_3007_411.n8 a_3007_411.t0 14.282
R879 a_3007_411.n5 a_3007_411.n3 8.58
R880 a_1666_101.t0 a_1666_101.n1 34.62
R881 a_1666_101.t0 a_1666_101.n0 8.137
R882 a_1666_101.t0 a_1666_101.n2 4.69
C4 VDD GND 17.44fF
C5 a_1666_101.n0 GND 0.05fF
C6 a_1666_101.n1 GND 0.12fF
C7 a_1666_101.n2 GND 0.04fF
C8 a_3007_411.n0 GND 0.38fF
C9 a_3007_411.n1 GND 0.84fF
C10 a_3007_411.n2 GND 0.21fF
C11 a_3007_411.n3 GND 0.05fF
C12 a_3007_411.n4 GND 0.06fF
C13 a_3007_411.n5 GND 0.21fF
C14 a_3007_411.n6 GND 0.52fF
C15 a_3007_411.n7 GND 0.84fF
C16 a_3007_411.n8 GND 0.76fF
C17 a_2405_209.n0 GND 0.37fF
C18 a_2405_209.t4 GND 0.67fF
C19 a_2405_209.n1 GND 1.07fF
C20 a_2405_209.n2 GND 0.50fF
C21 a_2405_209.n3 GND 1.18fF
C22 a_2405_209.n4 GND 0.83fF
C23 a_1771_1050.n0 GND 0.33fF
C24 a_1771_1050.t7 GND 0.45fF
C25 a_1771_1050.n1 GND 0.51fF
C26 a_1771_1050.n2 GND 0.04fF
C27 a_1771_1050.n3 GND 0.05fF
C28 a_1771_1050.n4 GND 0.03fF
C29 a_1771_1050.n5 GND 0.24fF
C30 a_1771_1050.n6 GND 0.51fF
C31 a_1771_1050.n7 GND 0.55fF
C32 a_1771_1050.n8 GND 0.30fF
C33 a_1771_1050.n9 GND 0.47fF
C34 a_2795_1051.n0 GND 0.55fF
C35 a_1295_209.n0 GND 0.44fF
C36 a_1295_209.n1 GND 1.26fF
C37 a_1295_209.n2 GND 0.47fF
C38 a_1295_209.n3 GND 1.34fF
C39 a_1295_209.n4 GND 0.88fF
C40 a_661_1050.n0 GND 0.35fF
C41 a_661_1050.t6 GND 0.47fF
C42 a_661_1050.n1 GND 0.53fF
C43 a_661_1050.n2 GND 0.34fF
C44 a_661_1050.n3 GND 0.56fF
C45 a_661_1050.n4 GND 0.58fF
C46 a_661_1050.n5 GND 0.31fF
C47 a_661_1050.n6 GND 0.49fF
C48 a_n259_209.n0 GND 0.42fF
C49 a_n259_209.n1 GND 0.38fF
C50 a_n259_209.n2 GND 0.38fF
C51 a_n259_209.t5 GND 0.46fF
C52 a_n259_209.n3 GND 0.36fF
C53 a_n259_209.n4 GND 1.53fF
C54 a_n259_209.n5 GND 0.31fF
C55 a_n259_209.n6 GND 0.47fF
C56 a_n259_209.n7 GND 0.75fF
C57 a_556_101.n0 GND 0.05fF
C58 a_556_101.n1 GND 0.12fF
C59 a_556_101.n2 GND 0.04fF
C60 a_185_209.n0 GND 0.39fF
C61 a_185_209.n1 GND 0.59fF
C62 a_185_209.n2 GND 0.40fF
C63 a_185_209.n3 GND 0.67fF
C64 a_185_209.n4 GND 0.75fF
C65 a_3461_1051.n0 GND 0.52fF
C66 VDD.n0 GND 0.14fF
C67 VDD.n1 GND 0.02fF
C68 VDD.n2 GND 0.02fF
C69 VDD.n3 GND 0.04fF
C70 VDD.n4 GND 0.01fF
C71 VDD.n6 GND 0.02fF
C72 VDD.n7 GND 0.02fF
C73 VDD.n9 GND 0.02fF
C74 VDD.n10 GND 0.02fF
C75 VDD.n12 GND 0.02fF
C76 VDD.n14 GND 0.43fF
C77 VDD.n16 GND 0.03fF
C78 VDD.n17 GND 0.02fF
C79 VDD.n18 GND 0.02fF
C80 VDD.n19 GND 0.02fF
C81 VDD.n20 GND 0.03fF
C82 VDD.n21 GND 0.26fF
C83 VDD.n22 GND 0.02fF
C84 VDD.n23 GND 0.03fF
C85 VDD.n24 GND 0.26fF
C86 VDD.n25 GND 0.01fF
C87 VDD.n26 GND 0.28fF
C88 VDD.n27 GND 0.01fF
C89 VDD.n28 GND 0.02fF
C90 VDD.n29 GND 0.02fF
C91 VDD.n30 GND 0.26fF
C92 VDD.n31 GND 0.01fF
C93 VDD.n32 GND 0.02fF
C94 VDD.n33 GND 0.00fF
C95 VDD.n34 GND 0.08fF
C96 VDD.n35 GND 0.02fF
C97 VDD.n36 GND 0.16fF
C98 VDD.n37 GND 0.13fF
C99 VDD.n38 GND 0.01fF
C100 VDD.n39 GND 0.02fF
C101 VDD.n40 GND 0.02fF
C102 VDD.n41 GND 0.10fF
C103 VDD.n42 GND 0.02fF
C104 VDD.n43 GND 0.13fF
C105 VDD.n44 GND 0.15fF
C106 VDD.n45 GND 0.01fF
C107 VDD.n46 GND 0.02fF
C108 VDD.n47 GND 0.02fF
C109 VDD.n48 GND 0.23fF
C110 VDD.n49 GND 0.01fF
C111 VDD.n50 GND 0.02fF
C112 VDD.n51 GND 0.02fF
C113 VDD.n52 GND 0.26fF
C114 VDD.n53 GND 0.01fF
C115 VDD.n54 GND 0.02fF
C116 VDD.n55 GND 0.03fF
C117 VDD.n56 GND 0.02fF
C118 VDD.n57 GND 0.02fF
C119 VDD.n58 GND 0.02fF
C120 VDD.n59 GND 0.20fF
C121 VDD.n60 GND 0.04fF
C122 VDD.n61 GND 0.03fF
C123 VDD.n62 GND 0.02fF
C124 VDD.n64 GND 0.02fF
C125 VDD.n65 GND 0.02fF
C126 VDD.n66 GND 0.02fF
C127 VDD.n67 GND 0.02fF
C128 VDD.n69 GND 0.02fF
C129 VDD.n70 GND 0.02fF
C130 VDD.n71 GND 0.02fF
C131 VDD.n73 GND 0.26fF
C132 VDD.n75 GND 0.02fF
C133 VDD.n76 GND 0.02fF
C134 VDD.n77 GND 0.03fF
C135 VDD.n78 GND 0.02fF
C136 VDD.n79 GND 0.26fF
C137 VDD.n80 GND 0.01fF
C138 VDD.n81 GND 0.02fF
C139 VDD.n82 GND 0.03fF
C140 VDD.n83 GND 0.26fF
C141 VDD.n84 GND 0.01fF
C142 VDD.n85 GND 0.02fF
C143 VDD.n86 GND 0.02fF
C144 VDD.n87 GND 0.26fF
C145 VDD.n88 GND 0.01fF
C146 VDD.n89 GND 0.02fF
C147 VDD.n90 GND 0.02fF
C148 VDD.n91 GND 0.28fF
C149 VDD.n92 GND 0.01fF
C150 VDD.n93 GND 0.02fF
C151 VDD.n94 GND 0.02fF
C152 VDD.n95 GND 0.16fF
C153 VDD.n96 GND 0.13fF
C154 VDD.n97 GND 0.01fF
C155 VDD.n98 GND 0.02fF
C156 VDD.n99 GND 0.02fF
C157 VDD.n100 GND 0.10fF
C158 VDD.n101 GND 0.02fF
C159 VDD.n102 GND 0.13fF
C160 VDD.n103 GND 0.15fF
C161 VDD.n104 GND 0.01fF
C162 VDD.n105 GND 0.02fF
C163 VDD.n106 GND 0.02fF
C164 VDD.n107 GND 0.23fF
C165 VDD.n108 GND 0.01fF
C166 VDD.n109 GND 0.02fF
C167 VDD.n110 GND 0.02fF
C168 VDD.n111 GND 0.26fF
C169 VDD.n112 GND 0.01fF
C170 VDD.n113 GND 0.02fF
C171 VDD.n114 GND 0.03fF
C172 VDD.n115 GND 0.02fF
C173 VDD.n116 GND 0.02fF
C174 VDD.n117 GND 0.02fF
C175 VDD.n118 GND 0.17fF
C176 VDD.n119 GND 0.04fF
C177 VDD.n120 GND 0.03fF
C178 VDD.n121 GND 0.02fF
C179 VDD.n122 GND 0.02fF
C180 VDD.n123 GND 0.02fF
C181 VDD.n124 GND 0.02fF
C182 VDD.n125 GND 0.02fF
C183 VDD.n127 GND 0.02fF
C184 VDD.n128 GND 0.02fF
C185 VDD.n129 GND 0.02fF
C186 VDD.n131 GND 0.26fF
C187 VDD.n133 GND 0.02fF
C188 VDD.n134 GND 0.02fF
C189 VDD.n135 GND 0.03fF
C190 VDD.n136 GND 0.02fF
C191 VDD.n137 GND 0.26fF
C192 VDD.n138 GND 0.01fF
C193 VDD.n139 GND 0.02fF
C194 VDD.n140 GND 0.03fF
C195 VDD.n141 GND 0.05fF
C196 VDD.n142 GND 0.14fF
C197 VDD.n143 GND 0.19fF
C198 VDD.n144 GND 0.01fF
C199 VDD.n145 GND 0.01fF
C200 VDD.n146 GND 0.02fF
C201 VDD.n147 GND 0.16fF
C202 VDD.n148 GND 0.01fF
C203 VDD.n149 GND 0.02fF
C204 VDD.n150 GND 0.02fF
C205 VDD.n151 GND 0.06fF
C206 VDD.n152 GND 0.14fF
C207 VDD.n153 GND 0.19fF
C208 VDD.n154 GND 0.01fF
C209 VDD.n155 GND 0.01fF
C210 VDD.n156 GND 0.02fF
C211 VDD.n157 GND 0.26fF
C212 VDD.n158 GND 0.01fF
C213 VDD.n159 GND 0.02fF
C214 VDD.n160 GND 0.03fF
C215 VDD.n161 GND 0.02fF
C216 VDD.n162 GND 0.02fF
C217 VDD.n163 GND 0.02fF
C218 VDD.n164 GND 0.17fF
C219 VDD.n165 GND 0.04fF
C220 VDD.n166 GND 0.03fF
C221 VDD.n167 GND 0.02fF
C222 VDD.n168 GND 0.02fF
C223 VDD.n169 GND 0.02fF
C224 VDD.n170 GND 0.02fF
C225 VDD.n171 GND 0.02fF
C226 VDD.n173 GND 0.02fF
C227 VDD.n174 GND 0.02fF
C228 VDD.n175 GND 0.02fF
C229 VDD.n177 GND 0.26fF
C230 VDD.n179 GND 0.02fF
C231 VDD.n180 GND 0.02fF
C232 VDD.n181 GND 0.03fF
C233 VDD.n182 GND 0.02fF
C234 VDD.n183 GND 0.26fF
C235 VDD.n184 GND 0.01fF
C236 VDD.n185 GND 0.02fF
C237 VDD.n186 GND 0.03fF
C238 VDD.n187 GND 0.23fF
C239 VDD.n188 GND 0.01fF
C240 VDD.n189 GND 0.05fF
C241 VDD.n190 GND 0.01fF
C242 VDD.n191 GND 0.02fF
C243 VDD.n192 GND 0.13fF
C244 VDD.n193 GND 0.16fF
C245 VDD.n194 GND 0.01fF
C246 VDD.n195 GND 0.02fF
C247 VDD.n196 GND 0.02fF
C248 VDD.n197 GND 0.28fF
C249 VDD.n198 GND 0.01fF
C250 VDD.n199 GND 0.10fF
C251 VDD.n200 GND 0.02fF
C252 VDD.n201 GND 0.02fF
C253 VDD.n202 GND 0.02fF
C254 VDD.n203 GND 0.16fF
C255 VDD.n204 GND 0.13fF
C256 VDD.n205 GND 0.01fF
C257 VDD.n206 GND 0.02fF
C258 VDD.n207 GND 0.02fF
C259 VDD.n208 GND 0.02fF
C260 VDD.n209 GND 0.02fF
C261 VDD.n210 GND 0.02fF
C262 VDD.n211 GND 0.11fF
C263 VDD.n212 GND 0.03fF
C264 VDD.n213 GND 0.02fF
C265 VDD.n214 GND 0.02fF
C266 VDD.n215 GND 0.02fF
C267 VDD.n216 GND 0.02fF
C268 VDD.n217 GND 0.02fF
C269 VDD.n219 GND 0.02fF
C270 VDD.n220 GND 0.02fF
C271 VDD.n221 GND 0.02fF
C272 VDD.n223 GND 0.43fF
C273 VDD.n225 GND 0.03fF
C274 VDD.n226 GND 0.03fF
C275 VDD.n227 GND 0.26fF
C276 VDD.n228 GND 0.02fF
C277 VDD.n229 GND 0.03fF
C278 VDD.n230 GND 0.03fF
C279 VDD.n231 GND 0.14fF
C280 VDD.n232 GND 0.19fF
C281 VDD.n233 GND 0.01fF
C282 VDD.n234 GND 0.06fF
C283 VDD.n235 GND 0.01fF
C284 VDD.n236 GND 0.02fF
C285 VDD.n237 GND 0.16fF
C286 VDD.n238 GND 0.01fF
C287 VDD.n239 GND 0.02fF
C288 VDD.n240 GND 0.02fF
C289 VDD.n241 GND 0.05fF
C290 VDD.n242 GND 0.14fF
C291 VDD.n243 GND 0.19fF
C292 VDD.n244 GND 0.01fF
C293 VDD.n245 GND 0.01fF
C294 VDD.n246 GND 0.02fF
C295 VDD.n247 GND 0.26fF
C296 VDD.n248 GND 0.01fF
C297 VDD.n249 GND 0.02fF
C298 VDD.n250 GND 0.03fF
C299 VDD.n251 GND 0.02fF
C300 VDD.n252 GND 0.26fF
C301 VDD.n253 GND 0.01fF
C302 VDD.n254 GND 0.02fF
C303 VDD.n255 GND 0.02fF
C304 VDD.n256 GND 0.02fF
C305 VDD.n257 GND 0.02fF
C306 VDD.n258 GND 0.02fF
C307 VDD.n259 GND 0.02fF
C308 VDD.n261 GND 0.02fF
C309 VDD.n262 GND 0.02fF
C310 VDD.n263 GND 0.02fF
C311 VDD.n264 GND 0.02fF
C312 VDD.n266 GND 0.03fF
C313 VDD.n267 GND 0.02fF
C314 VDD.n268 GND 0.14fF
C315 VDD.n269 GND 0.04fF
C316 VDD.n271 GND 0.26fF
C317 VDD.n273 GND 0.02fF
C318 VDD.n274 GND 0.02fF
C319 VDD.n275 GND 0.03fF
C320 VDD.n276 GND 0.02fF
C321 VDD.n277 GND 0.03fF
C322 VDD.n278 GND 0.06fF
C323 VDD.n279 GND 0.14fF
C324 VDD.n280 GND 0.19fF
C325 VDD.n281 GND 0.01fF
C326 VDD.n282 GND 0.01fF
C327 VDD.n283 GND 0.02fF
C328 VDD.n284 GND 0.16fF
C329 VDD.n285 GND 0.01fF
C330 VDD.n286 GND 0.02fF
C331 VDD.n287 GND 0.02fF
C332 VDD.n288 GND 0.05fF
C333 VDD.n289 GND 0.14fF
C334 VDD.n290 GND 0.19fF
C335 VDD.n291 GND 0.01fF
C336 VDD.n292 GND 0.01fF
C337 VDD.n293 GND 0.02fF
C338 VDD.n294 GND 0.26fF
C339 VDD.n295 GND 0.01fF
C340 VDD.n296 GND 0.02fF
C341 VDD.n297 GND 0.03fF
C342 VDD.n298 GND 0.02fF
C343 VDD.n299 GND 0.02fF
C344 VDD.n300 GND 0.02fF
C345 VDD.n301 GND 0.17fF
C346 VDD.n302 GND 0.04fF
C347 VDD.n303 GND 0.03fF
C348 VDD.n304 GND 0.02fF
C349 VDD.n305 GND 0.02fF
C350 VDD.n306 GND 0.02fF
C351 VDD.n307 GND 0.02fF
C352 VDD.n308 GND 0.02fF
C353 VDD.n310 GND 0.02fF
C354 VDD.n311 GND 0.02fF
C355 VDD.n312 GND 0.02fF
C356 VDD.n314 GND 0.26fF
C357 VDD.n316 GND 0.02fF
C358 VDD.n317 GND 0.02fF
C359 VDD.n318 GND 0.03fF
C360 VDD.n319 GND 0.02fF
C361 VDD.n320 GND 0.26fF
C362 VDD.n321 GND 0.01fF
C363 VDD.n322 GND 0.02fF
C364 VDD.n323 GND 0.03fF
C365 VDD.n324 GND 0.06fF
C366 VDD.n325 GND 0.23fF
C367 VDD.n326 GND 0.01fF
C368 VDD.n327 GND 0.01fF
C369 VDD.n328 GND 0.02fF
C370 VDD.n329 GND 0.13fF
C371 VDD.n330 GND 0.15fF
C372 VDD.n331 GND 0.01fF
C373 VDD.n332 GND 0.02fF
C374 VDD.n333 GND 0.02fF
C375 VDD.n334 GND 0.16fF
C376 VDD.n335 GND 0.13fF
C377 VDD.n336 GND 0.01fF
C378 VDD.n337 GND 0.02fF
C379 VDD.n338 GND 0.02fF
C380 VDD.n339 GND 0.10fF
C381 VDD.n340 GND 0.02fF
C382 VDD.n341 GND 0.28fF
C383 VDD.n342 GND 0.01fF
C384 VDD.n343 GND 0.02fF
C385 VDD.n344 GND 0.02fF
C386 VDD.n345 GND 0.13fF
C387 VDD.n346 GND 0.16fF
C388 VDD.n347 GND 0.01fF
C389 VDD.n348 GND 0.02fF
C390 VDD.n349 GND 0.02fF
C391 VDD.n350 GND 0.05fF
C392 VDD.n351 GND 0.23fF
C393 VDD.n352 GND 0.01fF
C394 VDD.n353 GND 0.01fF
C395 VDD.n354 GND 0.02fF
C396 VDD.n355 GND 0.26fF
C397 VDD.n356 GND 0.01fF
C398 VDD.n357 GND 0.02fF
C399 VDD.n358 GND 0.03fF
C400 VDD.n359 GND 0.02fF
C401 VDD.n360 GND 0.02fF
C402 VDD.n361 GND 0.02fF
C403 VDD.n362 GND 0.17fF
C404 VDD.n363 GND 0.04fF
C405 VDD.n364 GND 0.03fF
C406 VDD.n365 GND 0.02fF
C407 VDD.n366 GND 0.02fF
C408 VDD.n367 GND 0.02fF
C409 VDD.n368 GND 0.02fF
C410 VDD.n369 GND 0.02fF
C411 VDD.n371 GND 0.02fF
C412 VDD.n372 GND 0.02fF
C413 VDD.n373 GND 0.02fF
C414 VDD.n375 GND 0.26fF
C415 VDD.n377 GND 0.02fF
C416 VDD.n378 GND 0.02fF
C417 VDD.n379 GND 0.03fF
C418 VDD.n380 GND 0.02fF
C419 VDD.n381 GND 0.26fF
C420 VDD.n382 GND 0.01fF
C421 VDD.n383 GND 0.02fF
C422 VDD.n384 GND 0.03fF
C423 VDD.n385 GND 0.14fF
C424 VDD.n386 GND 0.19fF
C425 VDD.n387 GND 0.01fF
C426 VDD.n388 GND 0.06fF
C427 VDD.n389 GND 0.01fF
C428 VDD.n390 GND 0.02fF
C429 VDD.n391 GND 0.16fF
C430 VDD.n392 GND 0.01fF
C431 VDD.n393 GND 0.02fF
C432 VDD.n394 GND 0.02fF
C433 VDD.n395 GND 0.05fF
C434 VDD.n396 GND 0.14fF
C435 VDD.n397 GND 0.19fF
C436 VDD.n398 GND 0.01fF
C437 VDD.n399 GND 0.01fF
C438 VDD.n400 GND 0.02fF
C439 VDD.n401 GND 0.26fF
C440 VDD.n402 GND 0.01fF
C441 VDD.n403 GND 0.02fF
C442 VDD.n404 GND 0.03fF
C443 VDD.n405 GND 0.02fF
C444 VDD.n406 GND 0.26fF
C445 VDD.n407 GND 0.01fF
C446 VDD.n408 GND 0.02fF
C447 VDD.n409 GND 0.02fF
C448 VDD.n410 GND 0.02fF
C449 VDD.n411 GND 0.17fF
C450 VDD.n412 GND 0.04fF
C451 VDD.n413 GND 0.03fF
C452 VDD.n414 GND 0.02fF
C453 VDD.n415 GND 0.02fF
C454 VDD.n416 GND 0.02fF
C455 VDD.n417 GND 0.02fF
C456 VDD.n418 GND 0.02fF
C457 VDD.n420 GND 0.02fF
C458 VDD.n421 GND 0.02fF
C459 VDD.n422 GND 0.02fF
C460 VDD.n424 GND 0.26fF
C461 VDD.n426 GND 0.02fF
C462 VDD.n427 GND 0.02fF
C463 VDD.n428 GND 0.03fF
C464 VDD.n429 GND 0.02fF
C465 VDD.n430 GND 0.03fF
C466 VDD.n431 GND 0.06fF
C467 VDD.n432 GND 0.23fF
C468 VDD.n433 GND 0.01fF
C469 VDD.n434 GND 0.01fF
C470 VDD.n435 GND 0.02fF
C471 VDD.n436 GND 0.13fF
C472 VDD.n437 GND 0.15fF
C473 VDD.n438 GND 0.01fF
C474 VDD.n439 GND 0.02fF
C475 VDD.n440 GND 0.01fF
C476 Q.n0 GND 0.40fF
C477 Q.t5 GND 0.52fF
C478 Q.n1 GND 0.41fF
C479 Q.n2 GND 0.72fF
C480 Q.n3 GND 0.06fF
C481 Q.n4 GND 0.04fF
C482 Q.n5 GND 0.13fF
C483 Q.n6 GND 0.04fF
C484 Q.n7 GND 0.06fF
C485 Q.n8 GND 0.04fF
C486 Q.n9 GND 0.19fF
C487 Q.n10 GND 0.37fF
C488 Q.n11 GND 0.39fF
C489 Q.n12 GND 0.35fF
.ends
