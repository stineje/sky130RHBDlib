* SPICE3 file created from OR2X1.ext - technology: sky130A

.subckt OR2X1 Y A B VDD GND
X0 Y or2x1_pcell_0/m1_547_649# GND GND nshort w=3 l=0.15
X1 VDD or2x1_pcell_0/m1_547_649# Y VDD pshort w=2 l=0.15
X2 VDD A or2x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X3 or2x1_pcell_0/m1_547_649# B or2x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X4 or2x1_pcell_0/m1_547_649# A GND GND nshort w=3 l=0.15
X5 or2x1_pcell_0/m1_547_649# B GND GND nshort w=3 l=0.15
C0 VDD GND 3.21fF
.ends
