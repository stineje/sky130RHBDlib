* SPICE3 file created from DFFSNQNX1.ext - technology: sky130A

.subckt DFFSNQNX1 QN D CLK SN VDD VSS
X0 VDD D a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0.001182 pd=9.582 as=0 ps=0 w=2 l=0.15 M=2
X1 VDD a_1265_989 a_1905_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X2 a_3599_411 a_1265_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X3 a_1265_989 CLK a_2702_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X4 a_1905_1050 a_217_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X5 a_4294_210 SN a_4013_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X6 VDD a_343_411 a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X7 VDD a_217_1050 a_343_411 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X8 QN a_3599_411 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.00116 pd=9.16 as=0 ps=0 w=2 l=0.15 M=2
X9 a_1905_1050 a_1265_989 a_2000_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X10 VDD CLK a_343_411 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X11 QN a_343_411 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X12 VDD a_1905_1050 a_1265_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X13 a_343_411 a_1265_989 a_1038_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X14 VDD QN a_3599_411 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X15 VSS a_217_1050 a_757_103 VSS sky130_fd_pr__nfet_01v8 ad=0.0010746 pd=9.42 as=0 ps=0 w=3 l=0.15
X16 VDD a_1265_989 a_343_411 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X17 VSS D a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X18 VSS a_343_411 a_3368_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X19 VDD SN a_3599_411 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X20 a_1905_1050 SN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X21 VSS a_217_1050 a_1719_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X22 a_1038_210 CLK a_757_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X23 VSS a_1905_1050 a_2702_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X24 a_217_1050 a_343_411 a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X25 VDD CLK a_1265_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X26 a_2000_210 SN a_1719_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X27 a_3599_411 a_1265_989 a_4294_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X28 QN a_3599_411 a_3368_101 VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
X29 VSS QN a_4013_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 a_217_1050 VDD 2.52f
C1 a_343_411 CLK 2.41f
C2 a_343_411 VDD 6.03f
C3 a_1265_989 a_343_411 3.02f
C4 QN VDD 2.20f
C5 a_3599_411 VDD 2.82f
C6 a_1265_989 VDD 2.79f
C7 a_1905_1050 VDD 2.82f
C8 VDD VSS 7.98f
.ends
