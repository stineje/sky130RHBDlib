// File: pmos2.spi.PMOS2.pxi
// Created: Tue Oct 15 16:00:16 2024
// 
simulator lang=spectre
x_PM_PMOS2\%noxref_4 ( N_noxref_4_M0_noxref_g N_noxref_4_M1_noxref_g \
 N_noxref_4_c_18_n )  PM_PMOS2\%noxref_4
cc_1 ( noxref_1 noxref_2 ) capacitor c=0.0735271f //x=0.44 //y=-2 //x2=0.87 \
 //y2=-2
cc_2 ( noxref_1 noxref_3 ) capacitor c=0.0149132f //x=0.44 //y=-2 //x2=1.31 \
 //y2=-2
cc_3 ( noxref_1 N_noxref_4_M0_noxref_g ) capacitor c=0.0394719f //x=0.44 \
 //y=-2 //x2=0.795 //y2=-1
cc_4 ( noxref_2 noxref_3 ) capacitor c=0.0735271f //x=0.87 //y=-2 //x2=1.31 \
 //y2=-2
cc_5 ( noxref_2 N_noxref_4_M0_noxref_g ) capacitor c=0.0134243f //x=0.87 \
 //y=-2 //x2=0.795 //y2=-1
cc_6 ( noxref_2 N_noxref_4_M1_noxref_g ) capacitor c=0.0134243f //x=0.87 \
 //y=-2 //x2=1.235 //y2=-1
cc_7 ( noxref_2 N_noxref_4_c_18_n ) capacitor c=0.00261532f //x=0.87 //y=-2 \
 //x2=1.16 //y2=-2.23
cc_8 ( noxref_3 N_noxref_4_M1_noxref_g ) capacitor c=0.0394719f //x=1.31 \
 //y=-2 //x2=1.235 //y2=-1
