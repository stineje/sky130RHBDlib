* SPICE3 file created from VOTERN3X1.ext - technology: sky130A

.subckt VOTERN3X1 YN A B C VPB VNB
M1000 a_217_1005.t1 A VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VNB B a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=0.5373p pd=4.71u as=0p ps=0u
M1002 VNB a_1027_944# a_1444_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_217_1005.t7 a_1027_944# a_881_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_392_181.t5 a_1027_944# a_881_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_392_181.t1 A a_881_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t2 B a_217_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_881_1005.t4 a_1027_944# a_217_1005.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t0 A a_217_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_881_1005.t3 B a_217_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_881_1005.t6 a_1027_944# a_392_181.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_217_1005.t2 B VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_217_1005.t5 B a_881_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VNB B a_778_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_881_1005.t0 A a_392_181.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u






R0 VPB VPB.n109 122.382
R1 VPB.n75 VPB.n73 94.117
R2 VPB.n173 VPB.n171 94.117
R3 VPB.n39 VPB.n38 76
R4 VPB.n43 VPB.n42 76
R5 VPB.n47 VPB.n46 76
R6 VPB.n51 VPB.n50 76
R7 VPB.n77 VPB.n76 76
R8 VPB.n81 VPB.n80 76
R9 VPB.n85 VPB.n84 76
R10 VPB.n89 VPB.n88 76
R11 VPB.n187 VPB.n186 76
R12 VPB.n183 VPB.n182 76
R13 VPB.n179 VPB.n178 76
R14 VPB.n175 VPB.n174 76
R15 VPB.n149 VPB.n148 76
R16 VPB.n145 VPB.n144 76
R17 VPB.n140 VPB.n139 76
R18 VPB.n135 VPB.n134 76
R19 VPB.n128 VPB.n127 76
R20 VPB.n123 VPB.n122 76
R21 VPB.n118 VPB.n117 76
R22 VPB.n113 VPB.n112 76
R23 VPB.n154 VPB.n153 61.764
R24 VPB.n56 VPB.n55 61.764
R25 VPB.n114 VPB.t3 55.465
R26 VPB.n141 VPB.t0 55.465
R27 VPB.n137 VPB.n136 48.952
R28 VPB.n120 VPB.n119 44.502
R29 VPB.n130 VPB.n129 41.183
R30 VPB.n34 VPB.n33 35.118
R31 VPB.n112 VPB.n93 20.452
R32 VPB.n23 VPB.n20 20.452
R33 VPB.n132 VPB.n131 17.801
R34 VPB.n129 VPB.t1 14.282
R35 VPB.n129 VPB.t2 14.282
R36 VPB.n23 VPB.n22 13.653
R37 VPB.n22 VPB.n21 13.653
R38 VPB.n32 VPB.n31 13.653
R39 VPB.n31 VPB.n30 13.653
R40 VPB.n29 VPB.n25 13.653
R41 VPB.n25 VPB.n24 13.653
R42 VPB.n28 VPB.n27 13.653
R43 VPB.n27 VPB.n26 13.653
R44 VPB.n38 VPB.n37 13.653
R45 VPB.n37 VPB.n36 13.653
R46 VPB.n42 VPB.n41 13.653
R47 VPB.n41 VPB.n40 13.653
R48 VPB.n46 VPB.n45 13.653
R49 VPB.n45 VPB.n44 13.653
R50 VPB.n50 VPB.n49 13.653
R51 VPB.n49 VPB.n48 13.653
R52 VPB.n76 VPB.n75 13.653
R53 VPB.n75 VPB.n74 13.653
R54 VPB.n80 VPB.n79 13.653
R55 VPB.n79 VPB.n78 13.653
R56 VPB.n84 VPB.n83 13.653
R57 VPB.n83 VPB.n82 13.653
R58 VPB.n88 VPB.n87 13.653
R59 VPB.n87 VPB.n86 13.653
R60 VPB.n186 VPB.n185 13.653
R61 VPB.n185 VPB.n184 13.653
R62 VPB.n182 VPB.n181 13.653
R63 VPB.n181 VPB.n180 13.653
R64 VPB.n178 VPB.n177 13.653
R65 VPB.n177 VPB.n176 13.653
R66 VPB.n174 VPB.n173 13.653
R67 VPB.n173 VPB.n172 13.653
R68 VPB.n148 VPB.n147 13.653
R69 VPB.n147 VPB.n146 13.653
R70 VPB.n144 VPB.n143 13.653
R71 VPB.n143 VPB.n142 13.653
R72 VPB.n139 VPB.n138 13.653
R73 VPB.n138 VPB.n137 13.653
R74 VPB.n134 VPB.n133 13.653
R75 VPB.n133 VPB.n132 13.653
R76 VPB.n127 VPB.n126 13.653
R77 VPB.n126 VPB.n125 13.653
R78 VPB.n122 VPB.n121 13.653
R79 VPB.n121 VPB.n120 13.653
R80 VPB.n117 VPB.n116 13.653
R81 VPB.n116 VPB.n115 13.653
R82 VPB.n112 VPB.n111 13.653
R83 VPB.n111 VPB.n110 13.653
R84 VPB.n125 VPB.n124 13.35
R85 VPB.n71 VPB.n54 13.276
R86 VPB.n54 VPB.n52 13.276
R87 VPB.n169 VPB.n152 13.276
R88 VPB.n152 VPB.n150 13.276
R89 VPB.n93 VPB.n92 13.276
R90 VPB.n92 VPB.n90 13.276
R91 VPB.n20 VPB.n19 13.276
R92 VPB.n19 VPB.n17 13.276
R93 VPB.n32 VPB.n29 13.276
R94 VPB.n29 VPB.n28 13.276
R95 VPB.n76 VPB.n72 13.276
R96 VPB.n174 VPB.n170 13.276
R97 VPB.n4 VPB.n2 12.796
R98 VPB.n4 VPB.n3 12.564
R99 VPB.n13 VPB.n12 12.198
R100 VPB.n11 VPB.n10 12.198
R101 VPB.n7 VPB.n6 12.198
R102 VPB.n92 VPB.n91 7.5
R103 VPB.n98 VPB.n97 7.5
R104 VPB.n101 VPB.n100 7.5
R105 VPB.n103 VPB.n102 7.5
R106 VPB.n106 VPB.n105 7.5
R107 VPB.n94 VPB.n93 7.5
R108 VPB.n152 VPB.n151 7.5
R109 VPB.n164 VPB.n163 7.5
R110 VPB.n158 VPB.n157 7.5
R111 VPB.n160 VPB.n159 7.5
R112 VPB.n166 VPB.n156 7.5
R113 VPB.n166 VPB.n154 7.5
R114 VPB.n169 VPB.n168 7.5
R115 VPB.n54 VPB.n53 7.5
R116 VPB.n66 VPB.n65 7.5
R117 VPB.n60 VPB.n59 7.5
R118 VPB.n62 VPB.n61 7.5
R119 VPB.n68 VPB.n58 7.5
R120 VPB.n68 VPB.n56 7.5
R121 VPB.n71 VPB.n70 7.5
R122 VPB.n20 VPB.n16 7.5
R123 VPB.n2 VPB.n1 7.5
R124 VPB.n6 VPB.n5 7.5
R125 VPB.n10 VPB.n9 7.5
R126 VPB.n19 VPB.n18 7.5
R127 VPB.n14 VPB.n0 7.5
R128 VPB.n72 VPB.n71 7.176
R129 VPB.n170 VPB.n169 7.176
R130 VPB.n165 VPB.n162 6.729
R131 VPB.n161 VPB.n158 6.729
R132 VPB.n67 VPB.n64 6.729
R133 VPB.n63 VPB.n60 6.729
R134 VPB.n161 VPB.n160 6.728
R135 VPB.n165 VPB.n164 6.728
R136 VPB.n168 VPB.n167 6.728
R137 VPB.n63 VPB.n62 6.728
R138 VPB.n67 VPB.n66 6.728
R139 VPB.n70 VPB.n69 6.728
R140 VPB.n95 VPB.n94 6.728
R141 VPB.n99 VPB.n96 6.728
R142 VPB.n104 VPB.n101 6.728
R143 VPB.n108 VPB.n106 6.728
R144 VPB.n108 VPB.n107 6.728
R145 VPB.n104 VPB.n103 6.728
R146 VPB.n99 VPB.n98 6.728
R147 VPB.n134 VPB.n130 6.458
R148 VPB.n16 VPB.n15 6.398
R149 VPB.n156 VPB.n155 6.166
R150 VPB.n58 VPB.n57 6.166
R151 VPB.n33 VPB.n23 6.112
R152 VPB.n33 VPB.n32 6.101
R153 VPB.n110 VPB 4.45
R154 VPB.n117 VPB.n114 1.794
R155 VPB.n144 VPB.n141 1.435
R156 VPB.n14 VPB.n7 1.402
R157 VPB.n14 VPB.n8 1.402
R158 VPB.n14 VPB.n11 1.402
R159 VPB.n14 VPB.n13 1.402
R160 VPB.n15 VPB.n14 0.735
R161 VPB.n14 VPB.n4 0.735
R162 VPB.n166 VPB.n165 0.387
R163 VPB.n166 VPB.n161 0.387
R164 VPB.n167 VPB.n166 0.387
R165 VPB.n68 VPB.n67 0.387
R166 VPB.n68 VPB.n63 0.387
R167 VPB.n69 VPB.n68 0.387
R168 VPB.n109 VPB.n108 0.387
R169 VPB.n109 VPB.n104 0.387
R170 VPB.n109 VPB.n99 0.387
R171 VPB.n109 VPB.n95 0.387
R172 VPB.n77 VPB.n51 0.272
R173 VPB.n175 VPB.n149 0.272
R174 VPB.n113 VPB 0.198
R175 VPB.n35 VPB.n34 0.136
R176 VPB.n39 VPB.n35 0.136
R177 VPB.n43 VPB.n39 0.136
R178 VPB.n47 VPB.n43 0.136
R179 VPB.n51 VPB.n47 0.136
R180 VPB.n81 VPB.n77 0.136
R181 VPB.n85 VPB.n81 0.136
R182 VPB.n89 VPB.n85 0.136
R183 VPB.n187 VPB.n183 0.136
R184 VPB.n183 VPB.n179 0.136
R185 VPB.n179 VPB.n175 0.136
R186 VPB.n149 VPB.n145 0.136
R187 VPB.n145 VPB.n140 0.136
R188 VPB.n140 VPB.n135 0.136
R189 VPB.n135 VPB.n128 0.136
R190 VPB.n128 VPB.n123 0.136
R191 VPB.n123 VPB.n118 0.136
R192 VPB.n118 VPB.n113 0.136
R193 VPB VPB.n89 0.068
R194 VPB VPB.n187 0.068
R195 a_217_1005.n4 a_217_1005.n3 195.987
R196 a_217_1005.n2 a_217_1005.t7 89.553
R197 a_217_1005.n4 a_217_1005.n0 75.271
R198 a_217_1005.n3 a_217_1005.n2 75.214
R199 a_217_1005.n5 a_217_1005.n4 36.517
R200 a_217_1005.n3 a_217_1005.t4 14.338
R201 a_217_1005.n1 a_217_1005.t6 14.282
R202 a_217_1005.n1 a_217_1005.t5 14.282
R203 a_217_1005.n0 a_217_1005.t3 14.282
R204 a_217_1005.n0 a_217_1005.t2 14.282
R205 a_217_1005.n5 a_217_1005.t0 14.282
R206 a_217_1005.t1 a_217_1005.n5 14.282
R207 a_217_1005.n2 a_217_1005.n1 12.119
R208 a_881_1005.n4 a_881_1005.n3 196.002
R209 a_881_1005.n2 a_881_1005.t0 89.553
R210 a_881_1005.n5 a_881_1005.n4 75.27
R211 a_881_1005.n3 a_881_1005.n2 75.214
R212 a_881_1005.n4 a_881_1005.n0 36.52
R213 a_881_1005.n3 a_881_1005.t7 14.338
R214 a_881_1005.n0 a_881_1005.t5 14.282
R215 a_881_1005.n0 a_881_1005.t4 14.282
R216 a_881_1005.n1 a_881_1005.t1 14.282
R217 a_881_1005.n1 a_881_1005.t6 14.282
R218 a_881_1005.n5 a_881_1005.t2 14.282
R219 a_881_1005.t3 a_881_1005.n5 14.282
R220 a_881_1005.n2 a_881_1005.n1 12.119
R221 a_392_181.n13 a_392_181.n3 336.934
R222 a_392_181.n12 a_392_181.n11 98.501
R223 a_392_181.n12 a_392_181.n7 96.417
R224 a_392_181.n13 a_392_181.n12 78.403
R225 a_392_181.n3 a_392_181.n2 75.271
R226 a_392_181.n16 a_392_181.n0 55.263
R227 a_392_181.n7 a_392_181.n6 30
R228 a_392_181.n11 a_392_181.n10 30
R229 a_392_181.n15 a_392_181.n14 30
R230 a_392_181.n16 a_392_181.n15 25.263
R231 a_392_181.n5 a_392_181.n4 24.383
R232 a_392_181.n9 a_392_181.n8 24.383
R233 a_392_181.n7 a_392_181.n5 23.684
R234 a_392_181.n11 a_392_181.n9 23.684
R235 a_392_181.n15 a_392_181.n13 20.417
R236 a_392_181.n1 a_392_181.t0 14.282
R237 a_392_181.n1 a_392_181.t1 14.282
R238 a_392_181.n2 a_392_181.t4 14.282
R239 a_392_181.n2 a_392_181.t5 14.282
R240 a_392_181.n3 a_392_181.n1 12.119
R241 a_1444_73.t0 a_1444_73.n1 93.333
R242 a_1444_73.n4 a_1444_73.n2 55.07
R243 a_1444_73.t0 a_1444_73.n0 8.137
R244 a_1444_73.n4 a_1444_73.n3 4.619
R245 a_1444_73.t0 a_1444_73.n4 0.071
R246 a_112_73.t0 a_112_73.n0 93.333
R247 a_112_73.n2 a_112_73.n1 51.404
R248 a_112_73.t0 a_112_73.n6 7.911
R249 a_112_73.t0 a_112_73.n2 4.039
R250 a_112_73.n5 a_112_73.n3 4.032
R251 a_112_73.n5 a_112_73.n4 3.644
R252 a_112_73.t0 a_112_73.n5 1.099
R253 a_778_73.t0 a_778_73.n0 93.333
R254 a_778_73.n3 a_778_73.n1 55.048
R255 a_778_73.n3 a_778_73.n2 2.097
R256 a_778_73.t0 a_778_73.n3 0.11
R257 VNB VNB.n166 300.778
R258 VNB.n66 VNB.n65 199.897
R259 VNB.n15 VNB.n14 199.897
R260 VNB.n92 VNB.n90 154.509
R261 VNB.n35 VNB.n33 154.509
R262 VNB.n79 VNB.n72 84.842
R263 VNB.n22 VNB.n21 84.842
R264 VNB.n49 VNB.n4 84.842
R265 VNB.n153 VNB.n152 76
R266 VNB.n141 VNB.n140 76
R267 VNB.n137 VNB.n134 76
R268 VNB.n81 VNB.n80 36.678
R269 VNB.n24 VNB.n23 36.678
R270 VNB.n51 VNB.n50 36.678
R271 VNB.n125 VNB.n124 35.118
R272 VNB.n117 VNB.n114 20.452
R273 VNB.n154 VNB.n153 20.452
R274 VNB.n123 VNB.n122 13.653
R275 VNB.n122 VNB.n121 13.653
R276 VNB.n120 VNB.n119 13.653
R277 VNB.n119 VNB.n118 13.653
R278 VNB.n75 VNB.n74 13.653
R279 VNB.n74 VNB.n73 13.653
R280 VNB.n78 VNB.n77 13.653
R281 VNB.n77 VNB.n76 13.653
R282 VNB.n82 VNB.n81 13.653
R283 VNB.n85 VNB.n84 13.653
R284 VNB.n84 VNB.n83 13.653
R285 VNB.n88 VNB.n87 13.653
R286 VNB.n87 VNB.n86 13.653
R287 VNB.n93 VNB.n92 13.653
R288 VNB.n92 VNB.n91 13.653
R289 VNB.n96 VNB.n95 13.653
R290 VNB.n95 VNB.n94 13.653
R291 VNB.n99 VNB.n98 13.653
R292 VNB.n98 VNB.n97 13.653
R293 VNB.n137 VNB.n136 13.653
R294 VNB.n136 VNB.n135 13.653
R295 VNB.n140 VNB.n139 13.653
R296 VNB.n139 VNB.n138 13.653
R297 VNB.n25 VNB.n24 13.653
R298 VNB.n28 VNB.n27 13.653
R299 VNB.n27 VNB.n26 13.653
R300 VNB.n31 VNB.n30 13.653
R301 VNB.n30 VNB.n29 13.653
R302 VNB.n36 VNB.n35 13.653
R303 VNB.n35 VNB.n34 13.653
R304 VNB.n39 VNB.n38 13.653
R305 VNB.n38 VNB.n37 13.653
R306 VNB.n42 VNB.n41 13.653
R307 VNB.n41 VNB.n40 13.653
R308 VNB.n45 VNB.n44 13.653
R309 VNB.n44 VNB.n43 13.653
R310 VNB.n48 VNB.n47 13.653
R311 VNB.n47 VNB.n46 13.653
R312 VNB.n52 VNB.n51 13.653
R313 VNB.n55 VNB.n54 13.653
R314 VNB.n54 VNB.n53 13.653
R315 VNB.n153 VNB.n0 13.653
R316 VNB VNB.n0 13.653
R317 VNB.n117 VNB.n116 13.653
R318 VNB.n116 VNB.n115 13.653
R319 VNB.n161 VNB.n158 13.577
R320 VNB.n102 VNB.n100 13.276
R321 VNB.n114 VNB.n102 13.276
R322 VNB.n58 VNB.n56 13.276
R323 VNB.n71 VNB.n58 13.276
R324 VNB.n7 VNB.n5 13.276
R325 VNB.n20 VNB.n7 13.276
R326 VNB.n123 VNB.n120 13.276
R327 VNB.n78 VNB.n75 13.276
R328 VNB.n85 VNB.n82 13.276
R329 VNB.n88 VNB.n85 13.276
R330 VNB.n89 VNB.n88 13.276
R331 VNB.n93 VNB.n89 13.276
R332 VNB.n96 VNB.n93 13.276
R333 VNB.n99 VNB.n96 13.276
R334 VNB.n137 VNB.n99 13.276
R335 VNB.n140 VNB.n137 13.276
R336 VNB.n28 VNB.n25 13.276
R337 VNB.n31 VNB.n28 13.276
R338 VNB.n32 VNB.n31 13.276
R339 VNB.n36 VNB.n32 13.276
R340 VNB.n39 VNB.n36 13.276
R341 VNB.n42 VNB.n39 13.276
R342 VNB.n45 VNB.n42 13.276
R343 VNB.n48 VNB.n45 13.276
R344 VNB.n55 VNB.n52 13.276
R345 VNB.n153 VNB.n55 13.276
R346 VNB.n3 VNB.n1 13.276
R347 VNB.n154 VNB.n3 13.276
R348 VNB.n79 VNB.n78 10.764
R349 VNB.n49 VNB.n48 10.764
R350 VNB.n163 VNB.n162 7.5
R351 VNB.n64 VNB.n63 7.5
R352 VNB.n60 VNB.n59 7.5
R353 VNB.n58 VNB.n57 7.5
R354 VNB.n71 VNB.n70 7.5
R355 VNB.n13 VNB.n12 7.5
R356 VNB.n9 VNB.n8 7.5
R357 VNB.n7 VNB.n6 7.5
R358 VNB.n20 VNB.n19 7.5
R359 VNB.n155 VNB.n154 7.5
R360 VNB.n3 VNB.n2 7.5
R361 VNB.n160 VNB.n159 7.5
R362 VNB.n108 VNB.n107 7.5
R363 VNB.n104 VNB.n103 7.5
R364 VNB.n102 VNB.n101 7.5
R365 VNB.n114 VNB.n113 7.5
R366 VNB.n89 VNB.n71 7.176
R367 VNB.n32 VNB.n20 7.176
R368 VNB.n165 VNB.n163 7.011
R369 VNB.n67 VNB.n64 7.011
R370 VNB.n62 VNB.n60 7.011
R371 VNB.n16 VNB.n13 7.011
R372 VNB.n11 VNB.n9 7.011
R373 VNB.n110 VNB.n108 7.011
R374 VNB.n106 VNB.n104 7.011
R375 VNB.n70 VNB.n69 7.01
R376 VNB.n62 VNB.n61 7.01
R377 VNB.n67 VNB.n66 7.01
R378 VNB.n19 VNB.n18 7.01
R379 VNB.n11 VNB.n10 7.01
R380 VNB.n16 VNB.n15 7.01
R381 VNB.n113 VNB.n112 7.01
R382 VNB.n106 VNB.n105 7.01
R383 VNB.n110 VNB.n109 7.01
R384 VNB.n165 VNB.n164 7.01
R385 VNB.n161 VNB.n160 6.788
R386 VNB.n156 VNB.n155 6.788
R387 VNB.n124 VNB.n117 6.111
R388 VNB.n124 VNB.n123 6.1
R389 VNB.n82 VNB.n79 2.511
R390 VNB.n25 VNB.n22 2.511
R391 VNB.n52 VNB.n49 2.511
R392 VNB.n166 VNB.n157 0.921
R393 VNB.n166 VNB.n161 0.476
R394 VNB.n166 VNB.n156 0.475
R395 VNB.n131 VNB.n130 0.272
R396 VNB.n145 VNB.n144 0.272
R397 VNB.n68 VNB.n62 0.246
R398 VNB.n69 VNB.n68 0.246
R399 VNB.n68 VNB.n67 0.246
R400 VNB.n17 VNB.n11 0.246
R401 VNB.n18 VNB.n17 0.246
R402 VNB.n17 VNB.n16 0.246
R403 VNB.n111 VNB.n106 0.246
R404 VNB.n112 VNB.n111 0.246
R405 VNB.n111 VNB.n110 0.246
R406 VNB.n166 VNB.n165 0.246
R407 VNB.n152 VNB 0.198
R408 VNB.n126 VNB.n125 0.136
R409 VNB.n127 VNB.n126 0.136
R410 VNB.n128 VNB.n127 0.136
R411 VNB.n129 VNB.n128 0.136
R412 VNB.n130 VNB.n129 0.136
R413 VNB.n132 VNB.n131 0.136
R414 VNB.n133 VNB.n132 0.136
R415 VNB.n134 VNB.n133 0.136
R416 VNB.n142 VNB.n141 0.136
R417 VNB.n143 VNB.n142 0.136
R418 VNB.n144 VNB.n143 0.136
R419 VNB.n146 VNB.n145 0.136
R420 VNB.n147 VNB.n146 0.136
R421 VNB.n148 VNB.n147 0.136
R422 VNB.n149 VNB.n148 0.136
R423 VNB.n150 VNB.n149 0.136
R424 VNB.n151 VNB.n150 0.136
R425 VNB.n152 VNB.n151 0.136
R426 VNB.n134 VNB 0.068
R427 VNB.n141 VNB 0.068



























































































































































































































.ends
