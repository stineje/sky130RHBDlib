magic
tech sky130A
magscale 1 2
timestamp 1652323009
<< nwell >>
rect 87 786 579 1550
<< pwell >>
rect 34 542 632 544
rect -31 -30 697 542
rect 34 -34 632 -30
<< pdiffc >>
rect 141 1059 175 1093
rect 229 1059 263 1093
rect 405 1059 439 1093
<< psubdiff >>
rect 34 542 632 544
rect 31 482 635 542
rect 31 480 34 482
rect 632 480 635 482
rect 31 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 635 17
rect 31 -30 635 -17
rect 34 -34 632 -30
<< nsubdiff >>
rect 34 1497 632 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 632 1497
rect 34 822 632 884
<< psubdiffcont >>
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
<< poly >>
rect 168 375 198 413
rect 362 382 392 383
<< locali >>
rect 34 1497 632 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 632 1497
rect 34 1446 632 1463
rect 141 1093 175 1111
rect 141 1027 175 1059
rect 229 1093 263 1111
rect 229 1057 263 1059
rect 405 1093 439 1111
rect 405 1057 439 1059
rect 229 1023 535 1057
rect 353 908 361 942
rect 205 433 239 908
rect 353 441 387 908
rect 353 433 357 441
rect 501 348 535 1023
rect 413 314 535 348
rect 413 233 447 314
rect 219 34 253 167
rect 34 32 632 34
rect 31 17 635 32
rect 31 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 635 17
rect 31 -30 635 -17
rect 34 -34 632 -30
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
<< metal1 >>
rect 34 1497 632 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 632 1497
rect 34 1446 632 1463
rect 34 32 632 34
rect 31 17 635 32
rect 31 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 635 17
rect 31 -30 635 -17
rect 34 -34 632 -30
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 223 -1 0 417
box -32 -28 34 26
use nmos_bottom  nmos_bottom_0
timestamp 1651256857
transform -1 0 360 0 1 73
box 0 0 248 302
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 223 -1 0 941
box -32 -28 34 26
use pmos2  pmos2_0
timestamp 1648061063
transform 1 0 43 0 1 1404
box 52 -461 352 42
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 -1 369 1 0 415
box -32 -28 34 26
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1651256895
transform -1 0 554 0 1 73
box 0 0 248 309
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 377 -1 0 941
box -32 -28 34 26
use pmos2  pmos2_1
timestamp 1648061063
transform 1 0 219 0 1 1404
box 52 -461 352 42
use diff_ring_side  diff_ring_side_0
timestamp 1652319726
transform 1 0 666 0 1 0
box -87 -34 87 1550
use diff_ring_side  diff_ring_side_1
timestamp 1652319726
transform 1 0 0 0 1 0
box -87 -34 87 1550
<< end >>
