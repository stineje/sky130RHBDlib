// File: invx1_pcell.spi.INVX1_PCELL.pxi
// Created: Tue Oct 15 15:57:06 2024
// 
simulator lang=spectre
x_PM_INVX1_PCELL\%noxref_2 ( N_noxref_2_c_32_p N_noxref_2_c_19_p \
 N_noxref_2_c_14_n N_noxref_2_c_15_n N_noxref_2_M1_noxref_s \
 N_noxref_2_M2_noxref_d )  PM_INVX1_PCELL\%noxref_2
x_PM_INVX1_PCELL\%noxref_3 ( N_noxref_3_c_37_n N_noxref_3_M0_noxref_g \
 N_noxref_3_M1_noxref_g N_noxref_3_M2_noxref_g N_noxref_3_c_38_n \
 N_noxref_3_c_64_p N_noxref_3_c_65_p N_noxref_3_c_39_n N_noxref_3_c_52_n \
 N_noxref_3_c_53_n N_noxref_3_c_40_n N_noxref_3_c_55_p N_noxref_3_c_41_n \
 N_noxref_3_c_42_n N_noxref_3_c_43_n )  PM_INVX1_PCELL\%noxref_3
x_PM_INVX1_PCELL\%noxref_4 ( N_noxref_4_c_75_n N_noxref_4_c_89_n \
 N_noxref_4_c_78_n N_noxref_4_c_80_n N_noxref_4_c_76_n N_noxref_4_M0_noxref_d \
 N_noxref_4_M1_noxref_d )  PM_INVX1_PCELL\%noxref_4
cc_1 ( noxref_1 N_noxref_2_c_14_n ) capacitor c=0.00989031f //x=0.495 //y=0.37 \
 //x2=0.74 //y2=7.4
cc_2 ( noxref_1 N_noxref_2_c_15_n ) capacitor c=0.00989031f //x=0.495 //y=0.37 \
 //x2=1.48 //y2=7.4
cc_3 ( noxref_1 N_noxref_3_c_37_n ) capacitor c=0.0441241f //x=0.495 //y=0.37 \
 //x2=0.74 //y2=2.085
cc_4 ( noxref_1 N_noxref_3_c_38_n ) capacitor c=0.0436223f //x=0.495 //y=0.37 \
 //x2=0.85 //y2=0.91
cc_5 ( noxref_1 N_noxref_3_c_39_n ) capacitor c=0.0124051f //x=0.495 //y=0.37 \
 //x2=0.85 //y2=1.92
cc_6 ( noxref_1 N_noxref_3_c_40_n ) capacitor c=0.00483274f //x=0.495 //y=0.37 \
 //x2=1.225 //y2=0.755
cc_7 ( noxref_1 N_noxref_3_c_41_n ) capacitor c=0.0261956f //x=0.495 //y=0.37 \
 //x2=1.38 //y2=0.91
cc_8 ( noxref_1 N_noxref_3_c_42_n ) capacitor c=0.0074042f //x=0.495 //y=0.37 \
 //x2=1.38 //y2=1.255
cc_9 ( noxref_1 N_noxref_3_c_43_n ) capacitor c=0.0175388f //x=0.495 //y=0.37 \
 //x2=0.74 //y2=2.085
cc_10 ( noxref_1 N_noxref_4_c_75_n ) capacitor c=0.0422833f //x=0.495 //y=0.37 \
 //x2=1.395 //y2=2.08
cc_11 ( noxref_1 N_noxref_4_c_76_n ) capacitor c=8.10282e-19 //x=0.495 \
 //y=0.37 //x2=1.48 //y2=4.495
cc_12 ( noxref_1 N_noxref_4_M0_noxref_d ) capacitor c=0.112723f //x=0.495 \
 //y=0.37 //x2=0.925 //y2=0.91
cc_13 ( N_noxref_2_c_14_n N_noxref_3_c_37_n ) capacitor c=0.0276175f //x=0.74 \
 //y=7.4 //x2=0.74 //y2=2.085
cc_14 ( N_noxref_2_c_15_n N_noxref_3_c_37_n ) capacitor c=0.00144809f //x=1.48 \
 //y=7.4 //x2=0.74 //y2=2.085
cc_15 ( N_noxref_2_M1_noxref_s N_noxref_3_c_37_n ) capacitor c=0.00938034f \
 //x=0.54 //y=5.02 //x2=0.74 //y2=2.085
cc_16 ( N_noxref_2_c_19_p N_noxref_3_M1_noxref_g ) capacitor c=0.00748034f \
 //x=1.47 //y=7.4 //x2=0.895 //y2=6.02
cc_17 ( N_noxref_2_c_14_n N_noxref_3_M1_noxref_g ) capacitor c=0.0241676f \
 //x=0.74 //y=7.4 //x2=0.895 //y2=6.02
cc_18 ( N_noxref_2_M1_noxref_s N_noxref_3_M1_noxref_g ) capacitor c=0.0528676f \
 //x=0.54 //y=5.02 //x2=0.895 //y2=6.02
cc_19 ( N_noxref_2_c_19_p N_noxref_3_M2_noxref_g ) capacitor c=0.00697478f \
 //x=1.47 //y=7.4 //x2=1.335 //y2=6.02
cc_20 ( N_noxref_2_M2_noxref_d N_noxref_3_M2_noxref_g ) capacitor c=0.0528676f \
 //x=1.41 //y=5.02 //x2=1.335 //y2=6.02
cc_21 ( N_noxref_2_c_15_n N_noxref_3_c_52_n ) capacitor c=0.0287802f //x=1.48 \
 //y=7.4 //x2=1.26 //y2=4.79
cc_22 ( N_noxref_2_c_14_n N_noxref_3_c_53_n ) capacitor c=0.011132f //x=0.74 \
 //y=7.4 //x2=0.97 //y2=4.79
cc_23 ( N_noxref_2_M1_noxref_s N_noxref_3_c_53_n ) capacitor c=0.00665831f \
 //x=0.54 //y=5.02 //x2=0.97 //y2=4.79
cc_24 ( N_noxref_2_c_19_p N_noxref_4_c_78_n ) capacitor c=8.92854e-19 //x=1.47 \
 //y=7.4 //x2=1.395 //y2=4.58
cc_25 ( N_noxref_2_M2_noxref_d N_noxref_4_c_78_n ) capacitor c=0.00644908f \
 //x=1.41 //y=5.02 //x2=1.395 //y2=4.58
cc_26 ( N_noxref_2_c_14_n N_noxref_4_c_80_n ) capacitor c=0.0179238f //x=0.74 \
 //y=7.4 //x2=1.2 //y2=4.58
cc_27 ( N_noxref_2_c_14_n N_noxref_4_c_76_n ) capacitor c=4.80934e-19 //x=0.74 \
 //y=7.4 //x2=1.48 //y2=4.495
cc_28 ( N_noxref_2_c_15_n N_noxref_4_c_76_n ) capacitor c=0.0232778f //x=1.48 \
 //y=7.4 //x2=1.48 //y2=4.495
cc_29 ( N_noxref_2_c_32_p N_noxref_4_M1_noxref_d ) capacitor c=0.00722811f \
 //x=1.48 //y=7.4 //x2=0.97 //y2=5.02
cc_30 ( N_noxref_2_c_19_p N_noxref_4_M1_noxref_d ) capacitor c=0.0139004f \
 //x=1.47 //y=7.4 //x2=0.97 //y2=5.02
cc_31 ( N_noxref_2_c_15_n N_noxref_4_M1_noxref_d ) capacitor c=0.0219131f \
 //x=1.48 //y=7.4 //x2=0.97 //y2=5.02
cc_32 ( N_noxref_2_M1_noxref_s N_noxref_4_M1_noxref_d ) capacitor c=0.0843065f \
 //x=0.54 //y=5.02 //x2=0.97 //y2=5.02
cc_33 ( N_noxref_2_M2_noxref_d N_noxref_4_M1_noxref_d ) capacitor c=0.0832641f \
 //x=1.41 //y=5.02 //x2=0.97 //y2=5.02
cc_34 ( N_noxref_3_c_55_p N_noxref_4_c_75_n ) capacitor c=0.0023507f //x=1.225 \
 //y=1.41 //x2=1.395 //y2=2.08
cc_35 ( N_noxref_3_c_43_n N_noxref_4_c_89_n ) capacitor c=0.0167852f //x=0.74 \
 //y=2.085 //x2=1.195 //y2=2.08
cc_36 ( N_noxref_3_c_52_n N_noxref_4_c_78_n ) capacitor c=0.0107726f //x=1.26 \
 //y=4.79 //x2=1.395 //y2=4.58
cc_37 ( N_noxref_3_c_37_n N_noxref_4_c_80_n ) capacitor c=0.0250789f //x=0.74 \
 //y=2.085 //x2=1.2 //y2=4.58
cc_38 ( N_noxref_3_c_53_n N_noxref_4_c_80_n ) capacitor c=0.00962086f //x=0.97 \
 //y=4.79 //x2=1.2 //y2=4.58
cc_39 ( N_noxref_3_c_37_n N_noxref_4_c_76_n ) capacitor c=0.0739084f //x=0.74 \
 //y=2.085 //x2=1.48 //y2=4.495
cc_40 ( N_noxref_3_c_43_n N_noxref_4_c_76_n ) capacitor c=8.49451e-19 //x=0.74 \
 //y=2.085 //x2=1.48 //y2=4.495
cc_41 ( N_noxref_3_c_37_n N_noxref_4_M0_noxref_d ) capacitor c=0.0175773f \
 //x=0.74 //y=2.085 //x2=0.925 //y2=0.91
cc_42 ( N_noxref_3_c_38_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218556f \
 //x=0.85 //y=0.91 //x2=0.925 //y2=0.91
cc_43 ( N_noxref_3_c_64_p N_noxref_4_M0_noxref_d ) capacitor c=0.00347355f \
 //x=0.85 //y=1.255 //x2=0.925 //y2=0.91
cc_44 ( N_noxref_3_c_65_p N_noxref_4_M0_noxref_d ) capacitor c=0.00742431f \
 //x=0.85 //y=1.565 //x2=0.925 //y2=0.91
cc_45 ( N_noxref_3_c_39_n N_noxref_4_M0_noxref_d ) capacitor c=0.00957707f \
 //x=0.85 //y=1.92 //x2=0.925 //y2=0.91
cc_46 ( N_noxref_3_c_40_n N_noxref_4_M0_noxref_d ) capacitor c=0.00220879f \
 //x=1.225 //y=0.755 //x2=0.925 //y2=0.91
cc_47 ( N_noxref_3_c_55_p N_noxref_4_M0_noxref_d ) capacitor c=0.0138447f \
 //x=1.225 //y=1.41 //x2=0.925 //y2=0.91
cc_48 ( N_noxref_3_c_41_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218624f \
 //x=1.38 //y=0.91 //x2=0.925 //y2=0.91
cc_49 ( N_noxref_3_c_42_n N_noxref_4_M0_noxref_d ) capacitor c=0.00601286f \
 //x=1.38 //y=1.255 //x2=0.925 //y2=0.91
cc_50 ( N_noxref_3_M1_noxref_g N_noxref_4_M1_noxref_d ) capacitor c=0.0219309f \
 //x=0.895 //y=6.02 //x2=0.97 //y2=5.02
cc_51 ( N_noxref_3_M2_noxref_g N_noxref_4_M1_noxref_d ) capacitor c=0.021902f \
 //x=1.335 //y=6.02 //x2=0.97 //y2=5.02
cc_52 ( N_noxref_3_c_52_n N_noxref_4_M1_noxref_d ) capacitor c=0.0148755f \
 //x=1.26 //y=4.79 //x2=0.97 //y2=5.02
cc_53 ( N_noxref_3_c_53_n N_noxref_4_M1_noxref_d ) capacitor c=0.00307344f \
 //x=0.97 //y=4.79 //x2=0.97 //y2=5.02
