magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 638 203
rect 29 -17 63 21
<< scnmos >>
rect 80 47 110 177
rect 152 47 182 177
rect 267 47 297 177
rect 353 47 383 177
rect 439 47 469 177
rect 525 47 555 177
<< scpmoshvt >>
rect 80 297 110 497
rect 166 297 196 497
rect 267 297 297 497
rect 353 297 383 497
rect 439 297 469 497
rect 525 297 555 497
<< ndiff >>
rect 27 161 80 177
rect 27 127 35 161
rect 69 127 80 161
rect 27 93 80 127
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 47 152 177
rect 182 89 267 177
rect 182 55 207 89
rect 241 55 267 89
rect 182 47 267 55
rect 297 153 353 177
rect 297 119 308 153
rect 342 119 353 153
rect 297 47 353 119
rect 383 89 439 177
rect 383 55 394 89
rect 428 55 439 89
rect 383 47 439 55
rect 469 169 525 177
rect 469 135 480 169
rect 514 135 525 169
rect 469 101 525 135
rect 469 67 480 101
rect 514 67 525 101
rect 469 47 525 67
rect 555 89 612 177
rect 555 55 566 89
rect 600 55 612 89
rect 555 47 612 55
<< pdiff >>
rect 27 485 80 497
rect 27 451 35 485
rect 69 451 80 485
rect 27 417 80 451
rect 27 383 35 417
rect 69 383 80 417
rect 27 297 80 383
rect 110 477 166 497
rect 110 443 121 477
rect 155 443 166 477
rect 110 409 166 443
rect 110 375 121 409
rect 155 375 166 409
rect 110 297 166 375
rect 196 489 267 497
rect 196 455 214 489
rect 248 455 267 489
rect 196 421 267 455
rect 196 387 214 421
rect 248 387 267 421
rect 196 297 267 387
rect 297 477 353 497
rect 297 443 308 477
rect 342 443 353 477
rect 297 409 353 443
rect 297 375 308 409
rect 342 375 353 409
rect 297 297 353 375
rect 383 489 439 497
rect 383 455 394 489
rect 428 455 439 489
rect 383 421 439 455
rect 383 387 394 421
rect 428 387 439 421
rect 383 297 439 387
rect 469 477 525 497
rect 469 443 480 477
rect 514 443 525 477
rect 469 409 525 443
rect 469 375 480 409
rect 514 375 525 409
rect 469 341 525 375
rect 469 307 480 341
rect 514 307 525 341
rect 469 297 525 307
rect 555 489 612 497
rect 555 455 566 489
rect 600 455 612 489
rect 555 421 612 455
rect 555 387 566 421
rect 600 387 612 421
rect 555 297 612 387
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 207 55 241 89
rect 308 119 342 153
rect 394 55 428 89
rect 480 135 514 169
rect 480 67 514 101
rect 566 55 600 89
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 121 443 155 477
rect 121 375 155 409
rect 214 455 248 489
rect 214 387 248 421
rect 308 443 342 477
rect 308 375 342 409
rect 394 455 428 489
rect 394 387 428 421
rect 480 443 514 477
rect 480 375 514 409
rect 480 307 514 341
rect 566 455 600 489
rect 566 387 600 421
<< poly >>
rect 80 497 110 523
rect 166 497 196 523
rect 267 497 297 523
rect 353 497 383 523
rect 439 497 469 523
rect 525 497 555 523
rect 80 265 110 297
rect 166 265 196 297
rect 267 265 297 297
rect 353 265 383 297
rect 439 265 469 297
rect 525 265 555 297
rect 43 249 110 265
rect 43 215 53 249
rect 87 215 110 249
rect 43 199 110 215
rect 80 177 110 199
rect 152 249 206 265
rect 152 215 162 249
rect 196 215 206 249
rect 152 199 206 215
rect 267 249 555 265
rect 267 215 283 249
rect 317 215 351 249
rect 385 215 419 249
rect 453 215 487 249
rect 521 215 555 249
rect 267 199 555 215
rect 152 177 182 199
rect 267 177 297 199
rect 353 177 383 199
rect 439 177 469 199
rect 525 177 555 199
rect 80 21 110 47
rect 152 21 182 47
rect 267 21 297 47
rect 353 21 383 47
rect 439 21 469 47
rect 525 21 555 47
<< polycont >>
rect 53 215 87 249
rect 162 215 196 249
rect 283 215 317 249
rect 351 215 385 249
rect 419 215 453 249
rect 487 215 521 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 19 376 85 383
rect 121 477 157 493
rect 155 443 157 477
rect 121 409 157 443
rect 155 375 157 409
rect 198 489 264 527
rect 198 455 214 489
rect 248 455 264 489
rect 198 421 264 455
rect 198 387 214 421
rect 248 387 264 421
rect 306 477 344 493
rect 306 443 308 477
rect 342 443 344 477
rect 306 409 344 443
rect 121 350 157 375
rect 306 375 308 409
rect 342 375 344 409
rect 378 489 444 527
rect 378 455 394 489
rect 428 455 444 489
rect 378 421 444 455
rect 378 387 394 421
rect 428 387 444 421
rect 478 477 516 493
rect 478 443 480 477
rect 514 443 516 477
rect 478 409 516 443
rect 306 352 344 375
rect 478 375 480 409
rect 514 375 516 409
rect 550 489 616 527
rect 550 455 566 489
rect 600 455 616 489
rect 550 421 616 455
rect 550 387 566 421
rect 600 387 616 421
rect 478 353 516 375
rect 478 352 627 353
rect 25 249 87 323
rect 121 316 272 350
rect 230 271 272 316
rect 306 341 627 352
rect 306 307 480 341
rect 514 307 627 341
rect 25 215 53 249
rect 25 199 87 215
rect 121 249 196 265
rect 121 215 162 249
rect 121 199 196 215
rect 230 249 537 271
rect 230 215 283 249
rect 317 215 351 249
rect 385 215 419 249
rect 453 215 487 249
rect 521 215 537 249
rect 230 204 537 215
rect 230 161 272 204
rect 571 169 627 307
rect 19 127 35 161
rect 69 127 272 161
rect 19 123 272 127
rect 306 153 480 169
rect 19 93 85 123
rect 306 119 308 153
rect 342 135 480 153
rect 514 135 627 169
rect 342 123 627 135
rect 342 119 344 123
rect 306 103 344 119
rect 19 59 35 93
rect 69 59 85 93
rect 478 101 516 123
rect 19 51 85 59
rect 191 55 207 89
rect 241 55 257 89
rect 191 17 257 55
rect 378 55 394 89
rect 428 55 444 89
rect 378 17 444 55
rect 478 67 480 101
rect 514 67 516 101
rect 478 51 516 67
rect 550 55 566 89
rect 600 55 616 89
rect 550 17 616 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 581 153 615 187 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 121 221 155 255 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 and2_4
rlabel metal1 s 0 -48 644 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 644 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 3823880
string GDS_START 3818194
string path 0.000 0.000 16.100 0.000 
<< end >>
