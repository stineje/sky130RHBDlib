* SPICE3 file created from AOAI4X1.ext - technology: sky130A

.subckt AOAI4X1 YN A B C D VDD GND
M1000 a_864_209.t2 C.t0 a_797_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 GND A.t1 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=2.2948p pd=16.08u as=0p ps=0u
M1002 GND a_864_209.t4 a_1444_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t3 a_217_1050.t5 a_797_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 YN.t1 D.t0 VDD.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD.t4 A.t0 a_217_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 YN D.t1 a_1444_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1007 VDD.t6 B.t0 a_217_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t8 a_864_209.t5 YN.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_217_1050.t2 A.t2 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_797_1051.t2 C.t1 a_864_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_797_1051.t1 a_217_1050.t7 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VDD.t1 D.t2 YN.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_217_1050.t0 B.t2 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 YN.t3 a_864_209.t6 VDD.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 A VDD 0.08fF
C1 D YN 0.26fF
C2 VDD YN 1.33fF
C3 A B 0.27fF
C4 VDD C 0.07fF
C5 VDD D 0.07fF
C6 VDD B 0.07fF
R0 C.n0 C.t1 470.752
R1 C.n0 C.t0 384.527
R2 C.n1 C.t2 241.172
R3 C.n1 C.n0 110.173
R4 C.n2 C.n1 76
R5 C.n2 C 0.046
R6 a_797_1051.t0 a_797_1051.n0 101.66
R7 a_797_1051.n0 a_797_1051.t2 101.659
R8 a_797_1051.n0 a_797_1051.t3 14.294
R9 a_797_1051.n0 a_797_1051.t1 14.282
R10 a_864_209.n0 a_864_209.t5 480.392
R11 a_864_209.n0 a_864_209.t6 403.272
R12 a_864_209.n10 a_864_209.n9 244.994
R13 a_864_209.n1 a_864_209.t4 203.821
R14 a_864_209.n1 a_864_209.n0 178.106
R15 a_864_209.n9 a_864_209.n1 153.315
R16 a_864_209.n8 a_864_209.n7 133.539
R17 a_864_209.n9 a_864_209.n8 82.528
R18 a_864_209.n4 a_864_209.n2 80.526
R19 a_864_209.n8 a_864_209.n4 48.405
R20 a_864_209.n4 a_864_209.n3 30
R21 a_864_209.n7 a_864_209.n6 22.578
R22 a_864_209.n10 a_864_209.t1 14.282
R23 a_864_209.t2 a_864_209.n10 14.282
R24 a_864_209.n7 a_864_209.n5 8.58
R25 a_217_1050.n4 a_217_1050.t7 486.819
R26 a_217_1050.n4 a_217_1050.t5 384.527
R27 a_217_1050.n6 a_217_1050.n3 232.158
R28 a_217_1050.n5 a_217_1050.t6 197.395
R29 a_217_1050.n5 a_217_1050.n4 186.206
R30 a_217_1050.n6 a_217_1050.n5 153.315
R31 a_217_1050.n8 a_217_1050.n6 130.933
R32 a_217_1050.n3 a_217_1050.n2 76.002
R33 a_217_1050.n8 a_217_1050.n7 30
R34 a_217_1050.n9 a_217_1050.n0 24.383
R35 a_217_1050.n9 a_217_1050.n8 23.684
R36 a_217_1050.n1 a_217_1050.t3 14.282
R37 a_217_1050.n1 a_217_1050.t0 14.282
R38 a_217_1050.n2 a_217_1050.t1 14.282
R39 a_217_1050.n2 a_217_1050.t2 14.282
R40 a_217_1050.n3 a_217_1050.n1 12.85
R41 VDD.n83 VDD.n81 144.705
R42 VDD.n180 VDD.n178 144.705
R43 VDD.n44 VDD.n43 76
R44 VDD.n49 VDD.n48 76
R45 VDD.n54 VDD.n53 76
R46 VDD.n58 VDD.n57 76
R47 VDD.n85 VDD.n84 76
R48 VDD.n89 VDD.n88 76
R49 VDD.n93 VDD.n92 76
R50 VDD.n97 VDD.n96 76
R51 VDD.n198 VDD.n197 76
R52 VDD.n193 VDD.n192 76
R53 VDD.n186 VDD.n185 76
R54 VDD.n182 VDD.n181 76
R55 VDD.n155 VDD.n154 76
R56 VDD.n151 VDD.n150 76
R57 VDD.n146 VDD.n145 76
R58 VDD.n141 VDD.n140 76
R59 VDD.n135 VDD.n134 76
R60 VDD.n130 VDD.n129 76
R61 VDD.n125 VDD.n124 76
R62 VDD.n120 VDD.n119 76
R63 VDD.n121 VDD.t5 55.106
R64 VDD.n50 VDD.t9 55.106
R65 VDD.n147 VDD.t6 55.106
R66 VDD.n33 VDD.t1 55.106
R67 VDD.n188 VDD.n187 41.183
R68 VDD.n137 VDD.n136 40.824
R69 VDD.n28 VDD.n27 40.824
R70 VDD.n63 VDD.n62 36.774
R71 VDD.n171 VDD.n170 36.774
R72 VDD.n25 VDD.n24 36.608
R73 VDD.n143 VDD.n142 36.608
R74 VDD.n38 VDD.n37 34.942
R75 VDD.n46 VDD.n45 32.032
R76 VDD.n190 VDD.n189 32.032
R77 VDD.n127 VDD.n126 32.032
R78 VDD.n119 VDD.n116 21.841
R79 VDD.n23 VDD.n20 21.841
R80 VDD.n136 VDD.t0 14.282
R81 VDD.n136 VDD.t4 14.282
R82 VDD.n187 VDD.t2 14.282
R83 VDD.n187 VDD.t3 14.282
R84 VDD.n27 VDD.t7 14.282
R85 VDD.n27 VDD.t8 14.282
R86 VDD.n116 VDD.n99 14.167
R87 VDD.n99 VDD.n98 14.167
R88 VDD.n79 VDD.n60 14.167
R89 VDD.n60 VDD.n59 14.167
R90 VDD.n176 VDD.n157 14.167
R91 VDD.n157 VDD.n156 14.167
R92 VDD.n20 VDD.n19 14.167
R93 VDD.n19 VDD.n17 14.167
R94 VDD.n32 VDD.n31 14.167
R95 VDD.n84 VDD.n80 14.167
R96 VDD.n181 VDD.n177 14.167
R97 VDD.n23 VDD.n22 13.653
R98 VDD.n22 VDD.n21 13.653
R99 VDD.n36 VDD.n35 13.653
R100 VDD.n35 VDD.n34 13.653
R101 VDD.n32 VDD.n26 13.653
R102 VDD.n26 VDD.n25 13.653
R103 VDD.n31 VDD.n30 13.653
R104 VDD.n30 VDD.n29 13.653
R105 VDD.n43 VDD.n42 13.653
R106 VDD.n42 VDD.n41 13.653
R107 VDD.n48 VDD.n47 13.653
R108 VDD.n47 VDD.n46 13.653
R109 VDD.n53 VDD.n52 13.653
R110 VDD.n52 VDD.n51 13.653
R111 VDD.n57 VDD.n56 13.653
R112 VDD.n56 VDD.n55 13.653
R113 VDD.n84 VDD.n83 13.653
R114 VDD.n83 VDD.n82 13.653
R115 VDD.n88 VDD.n87 13.653
R116 VDD.n87 VDD.n86 13.653
R117 VDD.n92 VDD.n91 13.653
R118 VDD.n91 VDD.n90 13.653
R119 VDD.n96 VDD.n95 13.653
R120 VDD.n95 VDD.n94 13.653
R121 VDD.n197 VDD.n196 13.653
R122 VDD.n196 VDD.n195 13.653
R123 VDD.n192 VDD.n191 13.653
R124 VDD.n191 VDD.n190 13.653
R125 VDD.n185 VDD.n184 13.653
R126 VDD.n184 VDD.n183 13.653
R127 VDD.n181 VDD.n180 13.653
R128 VDD.n180 VDD.n179 13.653
R129 VDD.n154 VDD.n153 13.653
R130 VDD.n153 VDD.n152 13.653
R131 VDD.n150 VDD.n149 13.653
R132 VDD.n149 VDD.n148 13.653
R133 VDD.n145 VDD.n144 13.653
R134 VDD.n144 VDD.n143 13.653
R135 VDD.n140 VDD.n139 13.653
R136 VDD.n139 VDD.n138 13.653
R137 VDD.n134 VDD.n133 13.653
R138 VDD.n133 VDD.n132 13.653
R139 VDD.n129 VDD.n128 13.653
R140 VDD.n128 VDD.n127 13.653
R141 VDD.n124 VDD.n123 13.653
R142 VDD.n123 VDD.n122 13.653
R143 VDD.n119 VDD.n118 13.653
R144 VDD.n118 VDD.n117 13.653
R145 VDD.n4 VDD.n2 12.915
R146 VDD.n4 VDD.n3 12.66
R147 VDD.n13 VDD.n12 12.343
R148 VDD.n11 VDD.n10 12.343
R149 VDD.n7 VDD.n6 12.343
R150 VDD.n33 VDD.n32 11.806
R151 VDD.n31 VDD.n28 8.658
R152 VDD.n140 VDD.n137 8.658
R153 VDD.n80 VDD.n79 7.674
R154 VDD.n177 VDD.n176 7.674
R155 VDD.n74 VDD.n73 7.5
R156 VDD.n68 VDD.n67 7.5
R157 VDD.n70 VDD.n69 7.5
R158 VDD.n65 VDD.n64 7.5
R159 VDD.n79 VDD.n78 7.5
R160 VDD.n161 VDD.n160 7.5
R161 VDD.n164 VDD.n163 7.5
R162 VDD.n166 VDD.n165 7.5
R163 VDD.n169 VDD.n168 7.5
R164 VDD.n176 VDD.n175 7.5
R165 VDD.n111 VDD.n110 7.5
R166 VDD.n105 VDD.n104 7.5
R167 VDD.n107 VDD.n106 7.5
R168 VDD.n113 VDD.n103 7.5
R169 VDD.n113 VDD.n101 7.5
R170 VDD.n116 VDD.n115 7.5
R171 VDD.n20 VDD.n16 7.5
R172 VDD.n2 VDD.n1 7.5
R173 VDD.n6 VDD.n5 7.5
R174 VDD.n10 VDD.n9 7.5
R175 VDD.n19 VDD.n18 7.5
R176 VDD.n14 VDD.n0 7.5
R177 VDD.n66 VDD.n63 6.772
R178 VDD.n77 VDD.n61 6.772
R179 VDD.n75 VDD.n72 6.772
R180 VDD.n71 VDD.n68 6.772
R181 VDD.n114 VDD.n100 6.772
R182 VDD.n112 VDD.n109 6.772
R183 VDD.n108 VDD.n105 6.772
R184 VDD.n66 VDD.n65 6.772
R185 VDD.n71 VDD.n70 6.772
R186 VDD.n75 VDD.n74 6.772
R187 VDD.n78 VDD.n77 6.772
R188 VDD.n108 VDD.n107 6.772
R189 VDD.n112 VDD.n111 6.772
R190 VDD.n115 VDD.n114 6.772
R191 VDD.n175 VDD.n174 6.772
R192 VDD.n162 VDD.n159 6.772
R193 VDD.n167 VDD.n164 6.772
R194 VDD.n172 VDD.n169 6.772
R195 VDD.n172 VDD.n171 6.772
R196 VDD.n167 VDD.n166 6.772
R197 VDD.n162 VDD.n161 6.772
R198 VDD.n174 VDD.n158 6.772
R199 VDD.n37 VDD.n23 6.487
R200 VDD.n37 VDD.n36 6.475
R201 VDD.n16 VDD.n15 6.458
R202 VDD.n103 VDD.n102 6.202
R203 VDD.n192 VDD.n188 5.903
R204 VDD.n41 VDD.n40 4.576
R205 VDD.n195 VDD.n194 4.576
R206 VDD.n132 VDD.n131 4.576
R207 VDD.n53 VDD.n50 2.754
R208 VDD.n124 VDD.n121 2.754
R209 VDD.n36 VDD.n33 2.361
R210 VDD.n150 VDD.n147 2.361
R211 VDD.n14 VDD.n7 1.329
R212 VDD.n14 VDD.n8 1.329
R213 VDD.n14 VDD.n11 1.329
R214 VDD.n14 VDD.n13 1.329
R215 VDD.n15 VDD.n14 0.696
R216 VDD.n14 VDD.n4 0.696
R217 VDD.n76 VDD.n75 0.365
R218 VDD.n76 VDD.n71 0.365
R219 VDD.n76 VDD.n66 0.365
R220 VDD.n77 VDD.n76 0.365
R221 VDD.n113 VDD.n112 0.365
R222 VDD.n113 VDD.n108 0.365
R223 VDD.n114 VDD.n113 0.365
R224 VDD.n173 VDD.n172 0.365
R225 VDD.n173 VDD.n167 0.365
R226 VDD.n173 VDD.n162 0.365
R227 VDD.n174 VDD.n173 0.365
R228 VDD.n85 VDD.n58 0.29
R229 VDD.n182 VDD.n155 0.29
R230 VDD.n120 VDD 0.207
R231 VDD.n44 VDD.n39 0.181
R232 VDD.n141 VDD.n135 0.181
R233 VDD.n39 VDD.n38 0.145
R234 VDD.n49 VDD.n44 0.145
R235 VDD.n54 VDD.n49 0.145
R236 VDD.n58 VDD.n54 0.145
R237 VDD.n89 VDD.n85 0.145
R238 VDD.n93 VDD.n89 0.145
R239 VDD.n97 VDD.n93 0.145
R240 VDD.n198 VDD.n193 0.145
R241 VDD.n193 VDD.n186 0.145
R242 VDD.n186 VDD.n182 0.145
R243 VDD.n155 VDD.n151 0.145
R244 VDD.n151 VDD.n146 0.145
R245 VDD.n146 VDD.n141 0.145
R246 VDD.n135 VDD.n130 0.145
R247 VDD.n130 VDD.n125 0.145
R248 VDD.n125 VDD.n120 0.145
R249 VDD VDD.n97 0.09
R250 VDD VDD.n198 0.09
R251 D.n0 D.t2 472.359
R252 D.n0 D.t0 384.527
R253 D.n1 D.t1 267.725
R254 D.n1 D.n0 83.507
R255 D.n2 D.n1 76
R256 D.n2 D 0.046
R257 YN.n7 YN.n2 205.605
R258 YN.n7 YN.n6 157.486
R259 YN.n2 YN.n1 76.002
R260 YN.n8 YN.n7 76
R261 YN.n6 YN.n5 30
R262 YN.n4 YN.n3 24.383
R263 YN.n6 YN.n4 23.684
R264 YN.n0 YN.t0 14.282
R265 YN.n0 YN.t1 14.282
R266 YN.n1 YN.t4 14.282
R267 YN.n1 YN.t3 14.282
R268 YN.n2 YN.n0 12.85
R269 YN.n8 YN 0.046
R270 A.n0 A.t0 480.392
R271 A.n0 A.t2 403.272
R272 A.n1 A.t1 230.374
R273 A.n1 A.n0 151.553
R274 A.n2 A.n1 76
R275 A.n2 A 0.046
R276 GND.n29 GND.n27 219.745
R277 GND.n85 GND.n84 219.745
R278 GND.n29 GND.n28 85.529
R279 GND.n85 GND.n83 85.529
R280 GND.n55 GND.n54 76
R281 GND.n12 GND.n11 76
R282 GND.n20 GND.n19 76
R283 GND.n23 GND.n22 76
R284 GND.n26 GND.n25 76
R285 GND.n33 GND.n32 76
R286 GND.n40 GND.n39 76
R287 GND.n46 GND.n45 76
R288 GND.n52 GND.n51 76
R289 GND.n103 GND.n102 76
R290 GND.n100 GND.n99 76
R291 GND.n95 GND.n94 76
R292 GND.n88 GND.n87 76
R293 GND.n81 GND.n80 76
R294 GND.n78 GND.n77 76
R295 GND.n75 GND.n74 76
R296 GND.n72 GND.n71 76
R297 GND.n69 GND.n68 76
R298 GND.n66 GND.n65 76
R299 GND.n58 GND.n57 76
R300 GND.n17 GND.n16 63.835
R301 GND.n63 GND.n62 63.835
R302 GND.n8 GND.n7 34.942
R303 GND.n16 GND.n15 28.421
R304 GND.n62 GND.n61 28.421
R305 GND.n16 GND.n14 25.263
R306 GND.n62 GND.n60 25.263
R307 GND.n14 GND.n13 24.383
R308 GND.n60 GND.n59 24.383
R309 GND.n97 GND.n96 19.735
R310 GND.n50 GND.n49 19.735
R311 GND.n44 GND.n43 19.735
R312 GND.n37 GND.n36 19.735
R313 GND.n93 GND.n92 19.735
R314 GND.n43 GND.t3 19.724
R315 GND.n96 GND.t0 19.724
R316 GND.n6 GND.n5 14.167
R317 GND.n5 GND.n4 14.167
R318 GND.n32 GND.n30 14.167
R319 GND.n87 GND.n86 14.167
R320 GND.n57 GND.n56 13.653
R321 GND.n65 GND.n64 13.653
R322 GND.n68 GND.n67 13.653
R323 GND.n71 GND.n70 13.653
R324 GND.n74 GND.n73 13.653
R325 GND.n77 GND.n76 13.653
R326 GND.n80 GND.n79 13.653
R327 GND.n87 GND.n82 13.653
R328 GND.n94 GND.n89 13.653
R329 GND.n99 GND.n98 13.653
R330 GND.n102 GND.n101 13.653
R331 GND.n51 GND.n47 13.653
R332 GND.n45 GND.n41 13.653
R333 GND.n39 GND.n38 13.653
R334 GND.n32 GND.n31 13.653
R335 GND.n25 GND.n24 13.653
R336 GND.n22 GND.n21 13.653
R337 GND.n19 GND.n18 13.653
R338 GND.n11 GND.n10 13.653
R339 GND.n4 GND.n3 13.653
R340 GND.n5 GND.n2 13.653
R341 GND.n6 GND.n1 13.653
R342 GND.n92 GND.n91 12.837
R343 GND.n36 GND.n35 11.605
R344 GND.n35 GND.n34 9.809
R345 GND.n51 GND.n50 8.854
R346 GND.n91 GND.n90 7.566
R347 GND.n30 GND.n29 7.312
R348 GND.n86 GND.n85 7.312
R349 GND.n7 GND.n0 7.083
R350 GND.t3 GND.n42 7.04
R351 GND.n7 GND.n6 6.474
R352 GND.n49 GND.n48 5.774
R353 GND.n19 GND.n17 3.935
R354 GND.n45 GND.n44 3.935
R355 GND.n99 GND.n97 3.935
R356 GND.n65 GND.n63 3.935
R357 GND.n39 GND.n37 0.983
R358 GND.n94 GND.n93 0.983
R359 GND.n54 GND.n53 0.596
R360 GND.n33 GND.n26 0.29
R361 GND.n88 GND.n81 0.29
R362 GND.n55 GND 0.207
R363 GND.n12 GND.n9 0.181
R364 GND.n72 GND.n69 0.181
R365 GND.n9 GND.n8 0.145
R366 GND.n20 GND.n12 0.145
R367 GND.n23 GND.n20 0.145
R368 GND.n26 GND.n23 0.145
R369 GND.n40 GND.n33 0.145
R370 GND.n46 GND.n40 0.145
R371 GND.n52 GND.n46 0.145
R372 GND.n103 GND.n100 0.145
R373 GND.n100 GND.n95 0.145
R374 GND.n95 GND.n88 0.145
R375 GND.n81 GND.n78 0.145
R376 GND.n78 GND.n75 0.145
R377 GND.n75 GND.n72 0.145
R378 GND.n69 GND.n66 0.145
R379 GND.n66 GND.n58 0.145
R380 GND.n58 GND.n55 0.145
R381 GND GND.n52 0.09
R382 GND GND.n103 0.09
R383 a_112_101.n12 a_112_101.n11 26.811
R384 a_112_101.n6 a_112_101.n5 24.977
R385 a_112_101.n2 a_112_101.n1 24.877
R386 a_112_101.t0 a_112_101.n2 12.677
R387 a_112_101.t0 a_112_101.n3 11.595
R388 a_112_101.t1 a_112_101.n8 8.137
R389 a_112_101.t0 a_112_101.n4 7.273
R390 a_112_101.t0 a_112_101.n0 6.109
R391 a_112_101.t1 a_112_101.n7 4.864
R392 a_112_101.t0 a_112_101.n12 2.074
R393 a_112_101.n7 a_112_101.n6 1.13
R394 a_112_101.n12 a_112_101.t1 0.937
R395 a_112_101.t1 a_112_101.n10 0.804
R396 a_112_101.n10 a_112_101.n9 0.136
R397 a_1444_101.t0 a_1444_101.n1 34.62
R398 a_1444_101.t0 a_1444_101.n0 8.137
R399 a_1444_101.t0 a_1444_101.n2 4.69
R400 B.n0 B.t0 472.359
R401 B.n0 B.t2 384.527
R402 B.n1 B.t1 214.619
R403 B.n1 B.n0 136.613
R404 B.n2 B.n1 76
R405 B.n2 B 0.046
C7 VDD GND 8.14fF
C8 a_1444_101.n0 GND 0.05fF
C9 a_1444_101.n1 GND 0.12fF
C10 a_1444_101.n2 GND 0.04fF
C11 a_112_101.n0 GND 0.02fF
C12 a_112_101.n1 GND 0.10fF
C13 a_112_101.n2 GND 0.06fF
C14 a_112_101.n3 GND 0.06fF
C15 a_112_101.n4 GND 0.00fF
C16 a_112_101.n5 GND 0.04fF
C17 a_112_101.n6 GND 0.05fF
C18 a_112_101.n7 GND 0.02fF
C19 a_112_101.n8 GND 0.05fF
C20 a_112_101.n9 GND 0.07fF
C21 a_112_101.n10 GND 0.17fF
C22 a_112_101.t1 GND 0.22fF
C23 a_112_101.n11 GND 0.09fF
C24 a_112_101.n12 GND 0.00fF
C25 YN.n0 GND 0.48fF
C26 YN.n1 GND 0.56fF
C27 YN.n2 GND 0.33fF
C28 YN.n3 GND 0.04fF
C29 YN.n4 GND 0.05fF
C30 YN.n5 GND 0.03fF
C31 YN.n6 GND 0.21fF
C32 YN.n7 GND 0.38fF
C33 YN.n8 GND 0.01fF
C34 VDD.n0 GND 0.14fF
C35 VDD.n1 GND 0.02fF
C36 VDD.n2 GND 0.02fF
C37 VDD.n3 GND 0.04fF
C38 VDD.n4 GND 0.01fF
C39 VDD.n5 GND 0.02fF
C40 VDD.n6 GND 0.02fF
C41 VDD.n9 GND 0.02fF
C42 VDD.n10 GND 0.02fF
C43 VDD.n12 GND 0.02fF
C44 VDD.n14 GND 0.43fF
C45 VDD.n16 GND 0.03fF
C46 VDD.n17 GND 0.02fF
C47 VDD.n18 GND 0.02fF
C48 VDD.n19 GND 0.02fF
C49 VDD.n20 GND 0.03fF
C50 VDD.n21 GND 0.26fF
C51 VDD.n22 GND 0.02fF
C52 VDD.n23 GND 0.03fF
C53 VDD.n24 GND 0.13fF
C54 VDD.n25 GND 0.16fF
C55 VDD.n26 GND 0.01fF
C56 VDD.n27 GND 0.10fF
C57 VDD.n28 GND 0.02fF
C58 VDD.n29 GND 0.28fF
C59 VDD.n30 GND 0.01fF
C60 VDD.n31 GND 0.02fF
C61 VDD.n32 GND 0.02fF
C62 VDD.n33 GND 0.05fF
C63 VDD.n34 GND 0.23fF
C64 VDD.n35 GND 0.01fF
C65 VDD.n36 GND 0.01fF
C66 VDD.n37 GND 0.00fF
C67 VDD.n38 GND 0.08fF
C68 VDD.n39 GND 0.02fF
C69 VDD.n40 GND 0.16fF
C70 VDD.n41 GND 0.13fF
C71 VDD.n42 GND 0.01fF
C72 VDD.n43 GND 0.02fF
C73 VDD.n44 GND 0.02fF
C74 VDD.n45 GND 0.13fF
C75 VDD.n46 GND 0.15fF
C76 VDD.n47 GND 0.01fF
C77 VDD.n48 GND 0.02fF
C78 VDD.n49 GND 0.02fF
C79 VDD.n50 GND 0.06fF
C80 VDD.n51 GND 0.23fF
C81 VDD.n52 GND 0.01fF
C82 VDD.n53 GND 0.01fF
C83 VDD.n54 GND 0.02fF
C84 VDD.n55 GND 0.26fF
C85 VDD.n56 GND 0.01fF
C86 VDD.n57 GND 0.02fF
C87 VDD.n58 GND 0.03fF
C88 VDD.n59 GND 0.02fF
C89 VDD.n60 GND 0.02fF
C90 VDD.n61 GND 0.02fF
C91 VDD.n62 GND 0.20fF
C92 VDD.n63 GND 0.04fF
C93 VDD.n64 GND 0.03fF
C94 VDD.n65 GND 0.02fF
C95 VDD.n67 GND 0.02fF
C96 VDD.n68 GND 0.02fF
C97 VDD.n69 GND 0.02fF
C98 VDD.n70 GND 0.02fF
C99 VDD.n72 GND 0.02fF
C100 VDD.n73 GND 0.02fF
C101 VDD.n74 GND 0.02fF
C102 VDD.n76 GND 0.26fF
C103 VDD.n78 GND 0.02fF
C104 VDD.n79 GND 0.02fF
C105 VDD.n80 GND 0.03fF
C106 VDD.n81 GND 0.02fF
C107 VDD.n82 GND 0.26fF
C108 VDD.n83 GND 0.01fF
C109 VDD.n84 GND 0.02fF
C110 VDD.n85 GND 0.03fF
C111 VDD.n86 GND 0.26fF
C112 VDD.n87 GND 0.01fF
C113 VDD.n88 GND 0.02fF
C114 VDD.n89 GND 0.02fF
C115 VDD.n90 GND 0.26fF
C116 VDD.n91 GND 0.01fF
C117 VDD.n92 GND 0.02fF
C118 VDD.n93 GND 0.02fF
C119 VDD.n94 GND 0.28fF
C120 VDD.n95 GND 0.01fF
C121 VDD.n96 GND 0.02fF
C122 VDD.n97 GND 0.02fF
C123 VDD.n98 GND 0.02fF
C124 VDD.n99 GND 0.02fF
C125 VDD.n100 GND 0.02fF
C126 VDD.n101 GND 0.14fF
C127 VDD.n102 GND 0.03fF
C128 VDD.n103 GND 0.02fF
C129 VDD.n104 GND 0.02fF
C130 VDD.n105 GND 0.02fF
C131 VDD.n106 GND 0.02fF
C132 VDD.n107 GND 0.02fF
C133 VDD.n109 GND 0.02fF
C134 VDD.n110 GND 0.02fF
C135 VDD.n111 GND 0.02fF
C136 VDD.n113 GND 0.43fF
C137 VDD.n115 GND 0.03fF
C138 VDD.n116 GND 0.03fF
C139 VDD.n117 GND 0.26fF
C140 VDD.n118 GND 0.02fF
C141 VDD.n119 GND 0.03fF
C142 VDD.n120 GND 0.03fF
C143 VDD.n121 GND 0.06fF
C144 VDD.n122 GND 0.23fF
C145 VDD.n123 GND 0.01fF
C146 VDD.n124 GND 0.01fF
C147 VDD.n125 GND 0.02fF
C148 VDD.n126 GND 0.13fF
C149 VDD.n127 GND 0.15fF
C150 VDD.n128 GND 0.01fF
C151 VDD.n129 GND 0.02fF
C152 VDD.n130 GND 0.02fF
C153 VDD.n131 GND 0.16fF
C154 VDD.n132 GND 0.13fF
C155 VDD.n133 GND 0.01fF
C156 VDD.n134 GND 0.02fF
C157 VDD.n135 GND 0.02fF
C158 VDD.n136 GND 0.10fF
C159 VDD.n137 GND 0.02fF
C160 VDD.n138 GND 0.28fF
C161 VDD.n139 GND 0.01fF
C162 VDD.n140 GND 0.02fF
C163 VDD.n141 GND 0.02fF
C164 VDD.n142 GND 0.13fF
C165 VDD.n143 GND 0.16fF
C166 VDD.n144 GND 0.01fF
C167 VDD.n145 GND 0.02fF
C168 VDD.n146 GND 0.02fF
C169 VDD.n147 GND 0.05fF
C170 VDD.n148 GND 0.23fF
C171 VDD.n149 GND 0.01fF
C172 VDD.n150 GND 0.01fF
C173 VDD.n151 GND 0.02fF
C174 VDD.n152 GND 0.26fF
C175 VDD.n153 GND 0.01fF
C176 VDD.n154 GND 0.02fF
C177 VDD.n155 GND 0.03fF
C178 VDD.n156 GND 0.02fF
C179 VDD.n157 GND 0.02fF
C180 VDD.n158 GND 0.02fF
C181 VDD.n159 GND 0.02fF
C182 VDD.n160 GND 0.02fF
C183 VDD.n161 GND 0.02fF
C184 VDD.n163 GND 0.02fF
C185 VDD.n164 GND 0.02fF
C186 VDD.n165 GND 0.02fF
C187 VDD.n166 GND 0.02fF
C188 VDD.n168 GND 0.03fF
C189 VDD.n169 GND 0.02fF
C190 VDD.n170 GND 0.20fF
C191 VDD.n171 GND 0.04fF
C192 VDD.n173 GND 0.26fF
C193 VDD.n175 GND 0.02fF
C194 VDD.n176 GND 0.02fF
C195 VDD.n177 GND 0.03fF
C196 VDD.n178 GND 0.02fF
C197 VDD.n179 GND 0.26fF
C198 VDD.n180 GND 0.01fF
C199 VDD.n181 GND 0.02fF
C200 VDD.n182 GND 0.03fF
C201 VDD.n183 GND 0.23fF
C202 VDD.n184 GND 0.01fF
C203 VDD.n185 GND 0.02fF
C204 VDD.n186 GND 0.02fF
C205 VDD.n187 GND 0.10fF
C206 VDD.n188 GND 0.02fF
C207 VDD.n189 GND 0.13fF
C208 VDD.n190 GND 0.15fF
C209 VDD.n191 GND 0.01fF
C210 VDD.n192 GND 0.02fF
C211 VDD.n193 GND 0.02fF
C212 VDD.n194 GND 0.16fF
C213 VDD.n195 GND 0.13fF
C214 VDD.n196 GND 0.01fF
C215 VDD.n197 GND 0.02fF
C216 VDD.n198 GND 0.02fF
C217 a_217_1050.n0 GND 0.03fF
C218 a_217_1050.n1 GND 0.42fF
C219 a_217_1050.n2 GND 0.50fF
C220 a_217_1050.n3 GND 0.32fF
C221 a_217_1050.n4 GND 0.36fF
C222 a_217_1050.t6 GND 0.37fF
C223 a_217_1050.n5 GND 0.45fF
C224 a_217_1050.n6 GND 0.48fF
C225 a_217_1050.n7 GND 0.03fF
C226 a_217_1050.n8 GND 0.16fF
C227 a_217_1050.n9 GND 0.04fF
C228 a_864_209.n0 GND 0.39fF
C229 a_864_209.n1 GND 0.46fF
C230 a_864_209.n2 GND 0.05fF
C231 a_864_209.n3 GND 0.03fF
C232 a_864_209.n4 GND 0.10fF
C233 a_864_209.n5 GND 0.04fF
C234 a_864_209.n6 GND 0.04fF
C235 a_864_209.n7 GND 0.16fF
C236 a_864_209.n8 GND 0.27fF
C237 a_864_209.n9 GND 0.47fF
C238 a_864_209.n10 GND 0.63fF
C239 a_797_1051.n0 GND 0.54fF
.ends
