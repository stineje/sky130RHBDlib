// File: TMRDFFSNRNQX1.spi.pex
// Created: Tue Oct 15 15:53:14 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_TMRDFFSNRNQX1\%GND ( 1 167 171 174 179 189 197 207 215 225 233 243 \
 251 261 269 279 287 297 305 315 323 333 341 351 359 369 377 387 395 405 413 \
 423 431 441 449 459 467 477 485 495 503 511 517 523 531 542 547 551 564 566 \
 568 570 572 574 576 578 580 582 584 586 588 590 592 594 596 598 600 603 605 \
 612 619 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 \
 637 638 639 640 )
c1096 ( 640 0 ) capacitor c=0.0584744f //x=97.065 //y=0.37
c1097 ( 639 0 ) capacitor c=0.0215012f //x=94.23 //y=0.865
c1098 ( 638 0 ) capacitor c=0.0215012f //x=90.9 //y=0.865
c1099 ( 637 0 ) capacitor c=0.0207058f //x=87.57 //y=0.865
c1100 ( 636 0 ) capacitor c=0.0225954f //x=82.655 //y=0.875
c1101 ( 635 0 ) capacitor c=0.0225954f //x=77.845 //y=0.875
c1102 ( 634 0 ) capacitor c=0.0225954f //x=73.035 //y=0.875
c1103 ( 633 0 ) capacitor c=0.0225954f //x=68.225 //y=0.875
c1104 ( 632 0 ) capacitor c=0.0225954f //x=63.415 //y=0.875
c1105 ( 631 0 ) capacitor c=0.0225954f //x=58.605 //y=0.875
c1106 ( 630 0 ) capacitor c=0.0225954f //x=53.795 //y=0.875
c1107 ( 629 0 ) capacitor c=0.0225954f //x=48.985 //y=0.875
c1108 ( 628 0 ) capacitor c=0.0225954f //x=44.175 //y=0.875
c1109 ( 627 0 ) capacitor c=0.0225954f //x=39.365 //y=0.875
c1110 ( 626 0 ) capacitor c=0.0225954f //x=34.555 //y=0.875
c1111 ( 625 0 ) capacitor c=0.0225954f //x=29.745 //y=0.875
c1112 ( 624 0 ) capacitor c=0.0225954f //x=24.935 //y=0.875
c1113 ( 623 0 ) capacitor c=0.0225954f //x=20.125 //y=0.875
c1114 ( 622 0 ) capacitor c=0.0225954f //x=15.315 //y=0.875
c1115 ( 621 0 ) capacitor c=0.0225954f //x=10.505 //y=0.875
c1116 ( 620 0 ) capacitor c=0.0225954f //x=5.695 //y=0.875
c1117 ( 619 0 ) capacitor c=0.022675f //x=0.885 //y=0.875
c1118 ( 612 0 ) capacitor c=0.234368f //x=98.17 //y=0
c1119 ( 605 0 ) capacitor c=0.101943f //x=96.57 //y=0
c1120 ( 604 0 ) capacitor c=0.00440095f //x=94.42 //y=0
c1121 ( 603 0 ) capacitor c=0.101195f //x=93.24 //y=0
c1122 ( 602 0 ) capacitor c=0.00440095f //x=91.02 //y=0
c1123 ( 600 0 ) capacitor c=0.116097f //x=89.91 //y=0
c1124 ( 599 0 ) capacitor c=0.00440095f //x=87.76 //y=0
c1125 ( 598 0 ) capacitor c=0.107313f //x=86.58 //y=0
c1126 ( 597 0 ) capacitor c=0.00440144f //x=82.845 //y=0
c1127 ( 596 0 ) capacitor c=0.106956f //x=81.77 //y=0
c1128 ( 595 0 ) capacitor c=0.00440144f //x=78.035 //y=0
c1129 ( 594 0 ) capacitor c=0.106903f //x=76.96 //y=0
c1130 ( 593 0 ) capacitor c=0.00440144f //x=73.225 //y=0
c1131 ( 592 0 ) capacitor c=0.107052f //x=72.15 //y=0
c1132 ( 591 0 ) capacitor c=0.00440144f //x=68.415 //y=0
c1133 ( 590 0 ) capacitor c=0.107294f //x=67.34 //y=0
c1134 ( 589 0 ) capacitor c=0.00440144f //x=63.605 //y=0
c1135 ( 588 0 ) capacitor c=0.10703f //x=62.53 //y=0
c1136 ( 587 0 ) capacitor c=0.00440144f //x=58.795 //y=0
c1137 ( 586 0 ) capacitor c=0.107024f //x=57.72 //y=0
c1138 ( 585 0 ) capacitor c=0.00440144f //x=53.985 //y=0
c1139 ( 584 0 ) capacitor c=0.10703f //x=52.91 //y=0
c1140 ( 583 0 ) capacitor c=0.00440144f //x=49.175 //y=0
c1141 ( 582 0 ) capacitor c=0.106903f //x=48.1 //y=0
c1142 ( 581 0 ) capacitor c=0.00440144f //x=44.365 //y=0
c1143 ( 580 0 ) capacitor c=0.107052f //x=43.29 //y=0
c1144 ( 579 0 ) capacitor c=0.00440144f //x=39.555 //y=0
c1145 ( 578 0 ) capacitor c=0.107294f //x=38.48 //y=0
c1146 ( 577 0 ) capacitor c=0.00440144f //x=34.745 //y=0
c1147 ( 576 0 ) capacitor c=0.10703f //x=33.67 //y=0
c1148 ( 575 0 ) capacitor c=0.00440144f //x=29.935 //y=0
c1149 ( 574 0 ) capacitor c=0.107024f //x=28.86 //y=0
c1150 ( 573 0 ) capacitor c=0.00440144f //x=25.125 //y=0
c1151 ( 572 0 ) capacitor c=0.10703f //x=24.05 //y=0
c1152 ( 571 0 ) capacitor c=0.00440144f //x=20.315 //y=0
c1153 ( 570 0 ) capacitor c=0.106903f //x=19.24 //y=0
c1154 ( 569 0 ) capacitor c=0.00440144f //x=15.505 //y=0
c1155 ( 568 0 ) capacitor c=0.107052f //x=14.43 //y=0
c1156 ( 567 0 ) capacitor c=0.00440144f //x=10.695 //y=0
c1157 ( 566 0 ) capacitor c=0.107294f //x=9.62 //y=0
c1158 ( 565 0 ) capacitor c=0.00440144f //x=5.885 //y=0
c1159 ( 564 0 ) capacitor c=0.10703f //x=4.81 //y=0
c1160 ( 563 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c1161 ( 554 0 ) capacitor c=0.00583665f //x=98.17 //y=0.45
c1162 ( 551 0 ) capacitor c=0.00542558f //x=98.085 //y=0.535
c1163 ( 550 0 ) capacitor c=0.00479856f //x=97.685 //y=0.45
c1164 ( 547 0 ) capacitor c=0.00707849f //x=97.6 //y=0.535
c1165 ( 542 0 ) capacitor c=0.00588377f //x=97.2 //y=0.45
c1166 ( 539 0 ) capacitor c=0.0190475f //x=97.115 //y=0
c1167 ( 531 0 ) capacitor c=0.0749789f //x=96.4 //y=0
c1168 ( 523 0 ) capacitor c=0.0389876f //x=94.335 //y=0
c1169 ( 517 0 ) capacitor c=0.0716428f //x=93.07 //y=0
c1170 ( 511 0 ) capacitor c=0.0388276f //x=91.005 //y=0
c1171 ( 503 0 ) capacitor c=0.0717274f //x=89.74 //y=0
c1172 ( 495 0 ) capacitor c=0.039094f //x=87.675 //y=0
c1173 ( 485 0 ) capacitor c=0.133361f //x=86.41 //y=0
c1174 ( 477 0 ) capacitor c=0.0339325f //x=82.76 //y=0
c1175 ( 467 0 ) capacitor c=0.133559f //x=81.6 //y=0
c1176 ( 459 0 ) capacitor c=0.0339325f //x=77.95 //y=0
c1177 ( 449 0 ) capacitor c=0.133561f //x=76.79 //y=0
c1178 ( 441 0 ) capacitor c=0.0339325f //x=73.14 //y=0
c1179 ( 431 0 ) capacitor c=0.133362f //x=71.98 //y=0
c1180 ( 423 0 ) capacitor c=0.0339325f //x=68.33 //y=0
c1181 ( 413 0 ) capacitor c=0.133362f //x=67.17 //y=0
c1182 ( 405 0 ) capacitor c=0.0339325f //x=63.52 //y=0
c1183 ( 395 0 ) capacitor c=0.133362f //x=62.36 //y=0
c1184 ( 387 0 ) capacitor c=0.0339325f //x=58.71 //y=0
c1185 ( 377 0 ) capacitor c=0.133362f //x=57.55 //y=0
c1186 ( 369 0 ) capacitor c=0.0339325f //x=53.9 //y=0
c1187 ( 359 0 ) capacitor c=0.133362f //x=52.74 //y=0
c1188 ( 351 0 ) capacitor c=0.0339325f //x=49.09 //y=0
c1189 ( 341 0 ) capacitor c=0.133561f //x=47.93 //y=0
c1190 ( 333 0 ) capacitor c=0.0339325f //x=44.28 //y=0
c1191 ( 323 0 ) capacitor c=0.133362f //x=43.12 //y=0
c1192 ( 315 0 ) capacitor c=0.0339325f //x=39.47 //y=0
c1193 ( 305 0 ) capacitor c=0.133362f //x=38.31 //y=0
c1194 ( 297 0 ) capacitor c=0.0339325f //x=34.66 //y=0
c1195 ( 287 0 ) capacitor c=0.133362f //x=33.5 //y=0
c1196 ( 279 0 ) capacitor c=0.0339325f //x=29.85 //y=0
c1197 ( 269 0 ) capacitor c=0.133362f //x=28.69 //y=0
c1198 ( 261 0 ) capacitor c=0.0339325f //x=25.04 //y=0
c1199 ( 251 0 ) capacitor c=0.133362f //x=23.88 //y=0
c1200 ( 243 0 ) capacitor c=0.0339325f //x=20.23 //y=0
c1201 ( 233 0 ) capacitor c=0.133561f //x=19.07 //y=0
c1202 ( 225 0 ) capacitor c=0.0339325f //x=15.42 //y=0
c1203 ( 215 0 ) capacitor c=0.133362f //x=14.26 //y=0
c1204 ( 207 0 ) capacitor c=0.0339325f //x=10.61 //y=0
c1205 ( 197 0 ) capacitor c=0.133362f //x=9.45 //y=0
c1206 ( 189 0 ) capacitor c=0.0339325f //x=5.8 //y=0
c1207 ( 179 0 ) capacitor c=0.133402f //x=4.64 //y=0
c1208 ( 174 0 ) capacitor c=0.178058f //x=0.74 //y=0
c1209 ( 171 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c1210 ( 167 0 ) capacitor c=2.93672f //x=98.05 //y=0
r1211 (  611 612 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=98.05 //y=0 //x2=98.17 //y2=0
r1212 (  609 611 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=97.685 //y=0 //x2=98.05 //y2=0
r1213 (  608 609 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=97.31 //y=0 //x2=97.685 //y2=0
r1214 (  606 608 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=97.2 //y=0 //x2=97.31 //y2=0
r1215 (  555 640 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=98.17 //y=0.62 //x2=98.17 //y2=0.535
r1216 (  555 640 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=98.17 //y=0.62 //x2=98.17 //y2=1.225
r1217 (  554 640 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=98.17 //y=0.45 //x2=98.17 //y2=0.535
r1218 (  553 612 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=98.17 //y=0.17 //x2=98.17 //y2=0
r1219 (  553 554 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=98.17 //y=0.17 //x2=98.17 //y2=0.45
r1220 (  552 640 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=97.77 //y=0.535 //x2=97.685 //y2=0.535
r1221 (  551 640 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=98.085 //y=0.535 //x2=98.17 //y2=0.535
r1222 (  551 552 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=98.085 //y=0.535 //x2=97.77 //y2=0.535
r1223 (  550 640 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=97.685 //y=0.45 //x2=97.685 //y2=0.535
r1224 (  549 609 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=97.685 //y=0.17 //x2=97.685 //y2=0
r1225 (  549 550 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=97.685 //y=0.17 //x2=97.685 //y2=0.45
r1226 (  548 640 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=97.285 //y=0.535 //x2=97.2 //y2=0.535
r1227 (  547 640 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=97.6 //y=0.535 //x2=97.685 //y2=0.535
r1228 (  547 548 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=97.6 //y=0.535 //x2=97.285 //y2=0.535
r1229 (  543 640 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=97.2 //y=0.62 //x2=97.2 //y2=0.535
r1230 (  543 640 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=97.2 //y=0.62 //x2=97.2 //y2=1.225
r1231 (  542 640 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=97.2 //y=0.45 //x2=97.2 //y2=0.535
r1232 (  541 606 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=97.2 //y=0.17 //x2=97.2 //y2=0
r1233 (  541 542 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=97.2 //y=0.17 //x2=97.2 //y2=0.45
r1234 (  540 605 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=96.74 //y=0 //x2=96.57 //y2=0
r1235 (  539 606 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=97.115 //y=0 //x2=97.2 //y2=0
r1236 (  539 540 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=97.115 //y=0 //x2=96.74 //y2=0
r1237 (  534 536 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=94.72 //y=0 //x2=95.83 //y2=0
r1238 (  532 604 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.505 //y=0 //x2=94.42 //y2=0
r1239 (  532 534 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=94.505 //y=0 //x2=94.72 //y2=0
r1240 (  531 605 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=96.4 //y=0 //x2=96.57 //y2=0
r1241 (  531 536 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=96.4 //y=0 //x2=95.83 //y2=0
r1242 (  527 604 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=94.42 //y=0.17 //x2=94.42 //y2=0
r1243 (  527 639 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=94.42 //y=0.17 //x2=94.42 //y2=0.955
r1244 (  524 603 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=93.41 //y=0 //x2=93.24 //y2=0
r1245 (  524 526 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=93.41 //y=0 //x2=93.61 //y2=0
r1246 (  523 604 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.335 //y=0 //x2=94.42 //y2=0
r1247 (  523 526 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=94.335 //y=0 //x2=93.61 //y2=0
r1248 (  518 602 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.175 //y=0 //x2=91.09 //y2=0
r1249 (  518 520 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=91.175 //y=0 //x2=92.13 //y2=0
r1250 (  517 603 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=93.07 //y=0 //x2=93.24 //y2=0
r1251 (  517 520 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=93.07 //y=0 //x2=92.13 //y2=0
r1252 (  513 602 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=91.09 //y=0.17 //x2=91.09 //y2=0
r1253 (  513 638 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=91.09 //y=0.17 //x2=91.09 //y2=0.955
r1254 (  512 600 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=90.08 //y=0 //x2=89.91 //y2=0
r1255 (  511 602 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.005 //y=0 //x2=91.09 //y2=0
r1256 (  511 512 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=91.005 //y=0 //x2=90.08 //y2=0
r1257 (  506 508 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=88.43 //y=0 //x2=89.54 //y2=0
r1258 (  504 599 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=87.845 //y=0 //x2=87.76 //y2=0
r1259 (  504 506 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=87.845 //y=0 //x2=88.43 //y2=0
r1260 (  503 600 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=89.74 //y=0 //x2=89.91 //y2=0
r1261 (  503 508 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=89.74 //y=0 //x2=89.54 //y2=0
r1262 (  499 599 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=87.76 //y=0.17 //x2=87.76 //y2=0
r1263 (  499 637 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=87.76 //y=0.17 //x2=87.76 //y2=0.955
r1264 (  496 598 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=86.75 //y=0 //x2=86.58 //y2=0
r1265 (  496 498 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=86.75 //y=0 //x2=87.32 //y2=0
r1266 (  495 599 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=87.675 //y=0 //x2=87.76 //y2=0
r1267 (  495 498 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=87.675 //y=0 //x2=87.32 //y2=0
r1268 (  490 492 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=84.73 //y=0 //x2=85.84 //y2=0
r1269 (  488 490 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=83.62 //y=0 //x2=84.73 //y2=0
r1270 (  486 597 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.93 //y=0 //x2=82.845 //y2=0
r1271 (  486 488 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=82.93 //y=0 //x2=83.62 //y2=0
r1272 (  485 598 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=86.41 //y=0 //x2=86.58 //y2=0
r1273 (  485 492 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=86.41 //y=0 //x2=85.84 //y2=0
r1274 (  481 597 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=82.845 //y=0.17 //x2=82.845 //y2=0
r1275 (  481 636 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=82.845 //y=0.17 //x2=82.845 //y2=0.965
r1276 (  478 596 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.94 //y=0 //x2=81.77 //y2=0
r1277 (  478 480 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=81.94 //y=0 //x2=82.51 //y2=0
r1278 (  477 597 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.76 //y=0 //x2=82.845 //y2=0
r1279 (  477 480 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=82.76 //y=0 //x2=82.51 //y2=0
r1280 (  472 474 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=79.92 //y=0 //x2=81.03 //y2=0
r1281 (  470 472 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=78.81 //y=0 //x2=79.92 //y2=0
r1282 (  468 595 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.12 //y=0 //x2=78.035 //y2=0
r1283 (  468 470 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=78.12 //y=0 //x2=78.81 //y2=0
r1284 (  467 596 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.6 //y=0 //x2=81.77 //y2=0
r1285 (  467 474 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=81.6 //y=0 //x2=81.03 //y2=0
r1286 (  463 595 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=78.035 //y=0.17 //x2=78.035 //y2=0
r1287 (  463 635 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=78.035 //y=0.17 //x2=78.035 //y2=0.965
r1288 (  460 594 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.13 //y=0 //x2=76.96 //y2=0
r1289 (  460 462 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=77.13 //y=0 //x2=77.7 //y2=0
r1290 (  459 595 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.95 //y=0 //x2=78.035 //y2=0
r1291 (  459 462 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=77.95 //y=0 //x2=77.7 //y2=0
r1292 (  454 456 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=75.11 //y=0 //x2=76.22 //y2=0
r1293 (  452 454 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=74 //y=0 //x2=75.11 //y2=0
r1294 (  450 593 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.31 //y=0 //x2=73.225 //y2=0
r1295 (  450 452 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=73.31 //y=0 //x2=74 //y2=0
r1296 (  449 594 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.79 //y=0 //x2=76.96 //y2=0
r1297 (  449 456 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=76.79 //y=0 //x2=76.22 //y2=0
r1298 (  445 593 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.225 //y=0.17 //x2=73.225 //y2=0
r1299 (  445 634 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=73.225 //y=0.17 //x2=73.225 //y2=0.965
r1300 (  442 592 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=72.32 //y=0 //x2=72.15 //y2=0
r1301 (  442 444 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=72.32 //y=0 //x2=72.89 //y2=0
r1302 (  441 593 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.14 //y=0 //x2=73.225 //y2=0
r1303 (  441 444 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=73.14 //y=0 //x2=72.89 //y2=0
r1304 (  436 438 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=70.3 //y=0 //x2=71.41 //y2=0
r1305 (  434 436 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=69.19 //y=0 //x2=70.3 //y2=0
r1306 (  432 591 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.5 //y=0 //x2=68.415 //y2=0
r1307 (  432 434 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=68.5 //y=0 //x2=69.19 //y2=0
r1308 (  431 592 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.98 //y=0 //x2=72.15 //y2=0
r1309 (  431 438 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=71.98 //y=0 //x2=71.41 //y2=0
r1310 (  427 591 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.415 //y=0.17 //x2=68.415 //y2=0
r1311 (  427 633 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=68.415 //y=0.17 //x2=68.415 //y2=0.965
r1312 (  424 590 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.51 //y=0 //x2=67.34 //y2=0
r1313 (  424 426 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.51 //y=0 //x2=68.08 //y2=0
r1314 (  423 591 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.33 //y=0 //x2=68.415 //y2=0
r1315 (  423 426 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=68.33 //y=0 //x2=68.08 //y2=0
r1316 (  418 420 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=65.49 //y=0 //x2=66.6 //y2=0
r1317 (  416 418 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=64.38 //y=0 //x2=65.49 //y2=0
r1318 (  414 589 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.69 //y=0 //x2=63.605 //y2=0
r1319 (  414 416 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=63.69 //y=0 //x2=64.38 //y2=0
r1320 (  413 590 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.17 //y=0 //x2=67.34 //y2=0
r1321 (  413 420 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.17 //y=0 //x2=66.6 //y2=0
r1322 (  409 589 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=63.605 //y=0.17 //x2=63.605 //y2=0
r1323 (  409 632 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=63.605 //y=0.17 //x2=63.605 //y2=0.965
r1324 (  406 588 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.7 //y=0 //x2=62.53 //y2=0
r1325 (  406 408 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=62.7 //y=0 //x2=63.27 //y2=0
r1326 (  405 589 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.52 //y=0 //x2=63.605 //y2=0
r1327 (  405 408 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=63.52 //y=0 //x2=63.27 //y2=0
r1328 (  400 402 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=60.68 //y=0 //x2=61.79 //y2=0
r1329 (  398 400 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=59.57 //y=0 //x2=60.68 //y2=0
r1330 (  396 587 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.88 //y=0 //x2=58.795 //y2=0
r1331 (  396 398 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=58.88 //y=0 //x2=59.57 //y2=0
r1332 (  395 588 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.36 //y=0 //x2=62.53 //y2=0
r1333 (  395 402 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=62.36 //y=0 //x2=61.79 //y2=0
r1334 (  391 587 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.795 //y=0.17 //x2=58.795 //y2=0
r1335 (  391 631 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=58.795 //y=0.17 //x2=58.795 //y2=0.965
r1336 (  388 586 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.89 //y=0 //x2=57.72 //y2=0
r1337 (  388 390 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=57.89 //y=0 //x2=58.46 //y2=0
r1338 (  387 587 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.71 //y=0 //x2=58.795 //y2=0
r1339 (  387 390 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=58.71 //y=0 //x2=58.46 //y2=0
r1340 (  382 384 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=55.87 //y=0 //x2=56.98 //y2=0
r1341 (  380 382 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=54.76 //y=0 //x2=55.87 //y2=0
r1342 (  378 585 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.07 //y=0 //x2=53.985 //y2=0
r1343 (  378 380 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=54.07 //y=0 //x2=54.76 //y2=0
r1344 (  377 586 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.55 //y=0 //x2=57.72 //y2=0
r1345 (  377 384 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=57.55 //y=0 //x2=56.98 //y2=0
r1346 (  373 585 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.985 //y=0.17 //x2=53.985 //y2=0
r1347 (  373 630 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=53.985 //y=0.17 //x2=53.985 //y2=0.965
r1348 (  370 584 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.08 //y=0 //x2=52.91 //y2=0
r1349 (  370 372 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=53.08 //y=0 //x2=53.65 //y2=0
r1350 (  369 585 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.9 //y=0 //x2=53.985 //y2=0
r1351 (  369 372 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=53.9 //y=0 //x2=53.65 //y2=0
r1352 (  364 366 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=51.06 //y=0 //x2=52.17 //y2=0
r1353 (  362 364 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=49.95 //y=0 //x2=51.06 //y2=0
r1354 (  360 583 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.26 //y=0 //x2=49.175 //y2=0
r1355 (  360 362 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=49.26 //y=0 //x2=49.95 //y2=0
r1356 (  359 584 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.74 //y=0 //x2=52.91 //y2=0
r1357 (  359 366 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=52.74 //y=0 //x2=52.17 //y2=0
r1358 (  355 583 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.175 //y=0.17 //x2=49.175 //y2=0
r1359 (  355 629 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=49.175 //y=0.17 //x2=49.175 //y2=0.965
r1360 (  352 582 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.27 //y=0 //x2=48.1 //y2=0
r1361 (  352 354 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.27 //y=0 //x2=48.84 //y2=0
r1362 (  351 583 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.09 //y=0 //x2=49.175 //y2=0
r1363 (  351 354 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=49.09 //y=0 //x2=48.84 //y2=0
r1364 (  346 348 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=46.25 //y=0 //x2=47.36 //y2=0
r1365 (  344 346 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=45.14 //y=0 //x2=46.25 //y2=0
r1366 (  342 581 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.45 //y=0 //x2=44.365 //y2=0
r1367 (  342 344 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=44.45 //y=0 //x2=45.14 //y2=0
r1368 (  341 582 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.93 //y=0 //x2=48.1 //y2=0
r1369 (  341 348 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=47.93 //y=0 //x2=47.36 //y2=0
r1370 (  337 581 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.365 //y=0.17 //x2=44.365 //y2=0
r1371 (  337 628 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=44.365 //y=0.17 //x2=44.365 //y2=0.965
r1372 (  334 580 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.46 //y=0 //x2=43.29 //y2=0
r1373 (  334 336 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.46 //y=0 //x2=44.03 //y2=0
r1374 (  333 581 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.28 //y=0 //x2=44.365 //y2=0
r1375 (  333 336 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=44.28 //y=0 //x2=44.03 //y2=0
r1376 (  328 330 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=41.44 //y=0 //x2=42.55 //y2=0
r1377 (  326 328 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=40.33 //y=0 //x2=41.44 //y2=0
r1378 (  324 579 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.64 //y=0 //x2=39.555 //y2=0
r1379 (  324 326 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=39.64 //y=0 //x2=40.33 //y2=0
r1380 (  323 580 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.12 //y=0 //x2=43.29 //y2=0
r1381 (  323 330 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.12 //y=0 //x2=42.55 //y2=0
r1382 (  319 579 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.555 //y=0.17 //x2=39.555 //y2=0
r1383 (  319 627 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=39.555 //y=0.17 //x2=39.555 //y2=0.965
r1384 (  316 578 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.65 //y=0 //x2=38.48 //y2=0
r1385 (  316 318 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.65 //y=0 //x2=39.22 //y2=0
r1386 (  315 579 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.47 //y=0 //x2=39.555 //y2=0
r1387 (  315 318 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=39.47 //y=0 //x2=39.22 //y2=0
r1388 (  310 312 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=36.63 //y=0 //x2=37.74 //y2=0
r1389 (  308 310 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=35.52 //y=0 //x2=36.63 //y2=0
r1390 (  306 577 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.83 //y=0 //x2=34.745 //y2=0
r1391 (  306 308 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=34.83 //y=0 //x2=35.52 //y2=0
r1392 (  305 578 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.31 //y=0 //x2=38.48 //y2=0
r1393 (  305 312 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.31 //y=0 //x2=37.74 //y2=0
r1394 (  301 577 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.745 //y=0.17 //x2=34.745 //y2=0
r1395 (  301 626 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=34.745 //y=0.17 //x2=34.745 //y2=0.965
r1396 (  298 576 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.84 //y=0 //x2=33.67 //y2=0
r1397 (  298 300 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=33.84 //y=0 //x2=34.41 //y2=0
r1398 (  297 577 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.66 //y=0 //x2=34.745 //y2=0
r1399 (  297 300 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=34.66 //y=0 //x2=34.41 //y2=0
r1400 (  292 294 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=31.82 //y=0 //x2=32.93 //y2=0
r1401 (  290 292 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=30.71 //y=0 //x2=31.82 //y2=0
r1402 (  288 575 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.02 //y=0 //x2=29.935 //y2=0
r1403 (  288 290 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=30.02 //y=0 //x2=30.71 //y2=0
r1404 (  287 576 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.5 //y=0 //x2=33.67 //y2=0
r1405 (  287 294 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=33.5 //y=0 //x2=32.93 //y2=0
r1406 (  283 575 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.935 //y=0.17 //x2=29.935 //y2=0
r1407 (  283 625 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=29.935 //y=0.17 //x2=29.935 //y2=0.965
r1408 (  280 574 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.03 //y=0 //x2=28.86 //y2=0
r1409 (  280 282 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=29.03 //y=0 //x2=29.6 //y2=0
r1410 (  279 575 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.85 //y=0 //x2=29.935 //y2=0
r1411 (  279 282 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=29.85 //y=0 //x2=29.6 //y2=0
r1412 (  274 276 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=27.01 //y=0 //x2=28.12 //y2=0
r1413 (  272 274 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=25.9 //y=0 //x2=27.01 //y2=0
r1414 (  270 573 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.21 //y=0 //x2=25.125 //y2=0
r1415 (  270 272 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=25.21 //y=0 //x2=25.9 //y2=0
r1416 (  269 574 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.69 //y=0 //x2=28.86 //y2=0
r1417 (  269 276 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=28.69 //y=0 //x2=28.12 //y2=0
r1418 (  265 573 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.125 //y=0.17 //x2=25.125 //y2=0
r1419 (  265 624 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=25.125 //y=0.17 //x2=25.125 //y2=0.965
r1420 (  262 572 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.22 //y=0 //x2=24.05 //y2=0
r1421 (  262 264 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.22 //y=0 //x2=24.79 //y2=0
r1422 (  261 573 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.04 //y=0 //x2=25.125 //y2=0
r1423 (  261 264 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=25.04 //y=0 //x2=24.79 //y2=0
r1424 (  256 258 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=22.2 //y=0 //x2=23.31 //y2=0
r1425 (  254 256 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.09 //y=0 //x2=22.2 //y2=0
r1426 (  252 571 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.4 //y=0 //x2=20.315 //y2=0
r1427 (  252 254 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=20.4 //y=0 //x2=21.09 //y2=0
r1428 (  251 572 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.88 //y=0 //x2=24.05 //y2=0
r1429 (  251 258 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.88 //y=0 //x2=23.31 //y2=0
r1430 (  247 571 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.315 //y=0.17 //x2=20.315 //y2=0
r1431 (  247 623 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=20.315 //y=0.17 //x2=20.315 //y2=0.965
r1432 (  244 570 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.41 //y=0 //x2=19.24 //y2=0
r1433 (  244 246 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.41 //y=0 //x2=19.98 //y2=0
r1434 (  243 571 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.23 //y=0 //x2=20.315 //y2=0
r1435 (  243 246 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=20.23 //y=0 //x2=19.98 //y2=0
r1436 (  238 240 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.39 //y=0 //x2=18.5 //y2=0
r1437 (  236 238 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=16.28 //y=0 //x2=17.39 //y2=0
r1438 (  234 569 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.59 //y=0 //x2=15.505 //y2=0
r1439 (  234 236 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=15.59 //y=0 //x2=16.28 //y2=0
r1440 (  233 570 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.07 //y=0 //x2=19.24 //y2=0
r1441 (  233 240 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.07 //y=0 //x2=18.5 //y2=0
r1442 (  229 569 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.505 //y=0.17 //x2=15.505 //y2=0
r1443 (  229 622 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=15.505 //y=0.17 //x2=15.505 //y2=0.965
r1444 (  226 568 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=14.43 //y2=0
r1445 (  226 228 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=15.17 //y2=0
r1446 (  225 569 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.42 //y=0 //x2=15.505 //y2=0
r1447 (  225 228 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=15.42 //y=0 //x2=15.17 //y2=0
r1448 (  220 222 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=12.58 //y=0 //x2=13.69 //y2=0
r1449 (  218 220 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r1450 (  216 567 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.78 //y=0 //x2=10.695 //y2=0
r1451 (  216 218 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=10.78 //y=0 //x2=11.47 //y2=0
r1452 (  215 568 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=14.43 //y2=0
r1453 (  215 222 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=13.69 //y2=0
r1454 (  211 567 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.695 //y=0.17 //x2=10.695 //y2=0
r1455 (  211 621 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=10.695 //y=0.17 //x2=10.695 //y2=0.965
r1456 (  208 566 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=9.62 //y2=0
r1457 (  208 210 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=10.36 //y2=0
r1458 (  207 567 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.61 //y=0 //x2=10.695 //y2=0
r1459 (  207 210 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=10.61 //y=0 //x2=10.36 //y2=0
r1460 (  202 204 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.77 //y=0 //x2=8.88 //y2=0
r1461 (  200 202 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r1462 (  198 565 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=5.885 //y2=0
r1463 (  198 200 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=6.66 //y2=0
r1464 (  197 566 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=9.62 //y2=0
r1465 (  197 204 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=8.88 //y2=0
r1466 (  193 565 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0
r1467 (  193 620 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0.965
r1468 (  190 564 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=4.81 //y2=0
r1469 (  190 192 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=5.55 //y2=0
r1470 (  189 565 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.885 //y2=0
r1471 (  189 192 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.55 //y2=0
r1472 (  184 186 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r1473 (  182 184 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r1474 (  180 563 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r1475 (  180 182 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r1476 (  179 564 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.81 //y2=0
r1477 (  179 186 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r1478 (  175 563 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r1479 (  175 619 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r1480 (  171 563 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r1481 (  171 174 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r1482 (  167 611 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=98.05 //y=0 //x2=98.05 //y2=0
r1483 (  165 608 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=97.31 //y=0 //x2=97.31 //y2=0
r1484 (  165 167 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=97.31 //y=0 //x2=98.05 //y2=0
r1485 (  163 536 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=95.83 //y=0 //x2=95.83 //y2=0
r1486 (  163 165 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=95.83 //y=0 //x2=97.31 //y2=0
r1487 (  161 534 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=94.72 //y=0 //x2=94.72 //y2=0
r1488 (  161 163 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=94.72 //y=0 //x2=95.83 //y2=0
r1489 (  159 526 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=93.61 //y=0 //x2=93.61 //y2=0
r1490 (  159 161 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=93.61 //y=0 //x2=94.72 //y2=0
r1491 (  157 520 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=92.13 //y=0 //x2=92.13 //y2=0
r1492 (  157 159 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=92.13 //y=0 //x2=93.61 //y2=0
r1493 (  155 602 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=91.02 //y=0 //x2=91.02 //y2=0
r1494 (  155 157 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=91.02 //y=0 //x2=92.13 //y2=0
r1495 (  153 508 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=89.54 //y=0 //x2=89.54 //y2=0
r1496 (  153 155 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=89.54 //y=0 //x2=91.02 //y2=0
r1497 (  151 506 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=88.43 //y=0 //x2=88.43 //y2=0
r1498 (  151 153 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=88.43 //y=0 //x2=89.54 //y2=0
r1499 (  149 498 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=87.32 //y=0 //x2=87.32 //y2=0
r1500 (  149 151 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=87.32 //y=0 //x2=88.43 //y2=0
r1501 (  147 492 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=85.84 //y=0 //x2=85.84 //y2=0
r1502 (  147 149 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=85.84 //y=0 //x2=87.32 //y2=0
r1503 (  145 490 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=84.73 //y=0 //x2=84.73 //y2=0
r1504 (  145 147 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=84.73 //y=0 //x2=85.84 //y2=0
r1505 (  143 488 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=83.62 //y=0 //x2=83.62 //y2=0
r1506 (  143 145 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=83.62 //y=0 //x2=84.73 //y2=0
r1507 (  141 480 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.51 //y=0 //x2=82.51 //y2=0
r1508 (  141 143 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=82.51 //y=0 //x2=83.62 //y2=0
r1509 (  139 474 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=81.03 //y=0 //x2=81.03 //y2=0
r1510 (  139 141 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=81.03 //y=0 //x2=82.51 //y2=0
r1511 (  137 472 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=79.92 //y=0 //x2=79.92 //y2=0
r1512 (  137 139 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=79.92 //y=0 //x2=81.03 //y2=0
r1513 (  135 470 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.81 //y=0 //x2=78.81 //y2=0
r1514 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=78.81 //y=0 //x2=79.92 //y2=0
r1515 (  133 462 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=77.7 //y=0 //x2=77.7 //y2=0
r1516 (  133 135 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=77.7 //y=0 //x2=78.81 //y2=0
r1517 (  131 456 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.22 //y=0 //x2=76.22 //y2=0
r1518 (  131 133 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.22 //y=0 //x2=77.7 //y2=0
r1519 (  129 454 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.11 //y=0 //x2=75.11 //y2=0
r1520 (  129 131 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=0 //x2=76.22 //y2=0
r1521 (  127 452 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74 //y=0 //x2=74 //y2=0
r1522 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74 //y=0 //x2=75.11 //y2=0
r1523 (  125 444 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.89 //y=0 //x2=72.89 //y2=0
r1524 (  125 127 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=72.89 //y=0 //x2=74 //y2=0
r1525 (  123 438 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=0 //x2=71.41 //y2=0
r1526 (  123 125 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=0 //x2=72.89 //y2=0
r1527 (  121 436 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=70.3 //y=0 //x2=70.3 //y2=0
r1528 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=70.3 //y=0 //x2=71.41 //y2=0
r1529 (  119 434 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.19 //y=0 //x2=69.19 //y2=0
r1530 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.19 //y=0 //x2=70.3 //y2=0
r1531 (  117 426 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=68.08 //y=0 //x2=68.08 //y2=0
r1532 (  117 119 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=68.08 //y=0 //x2=69.19 //y2=0
r1533 (  115 420 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.6 //y=0 //x2=66.6 //y2=0
r1534 (  115 117 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=66.6 //y=0 //x2=68.08 //y2=0
r1535 (  113 418 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.49 //y=0 //x2=65.49 //y2=0
r1536 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.49 //y=0 //x2=66.6 //y2=0
r1537 (  111 416 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=64.38 //y=0 //x2=64.38 //y2=0
r1538 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=64.38 //y=0 //x2=65.49 //y2=0
r1539 (  109 408 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=63.27 //y=0 //x2=63.27 //y2=0
r1540 (  109 111 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=63.27 //y=0 //x2=64.38 //y2=0
r1541 (  107 402 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.79 //y=0 //x2=61.79 //y2=0
r1542 (  107 109 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.79 //y=0 //x2=63.27 //y2=0
r1543 (  105 400 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=60.68 //y=0 //x2=60.68 //y2=0
r1544 (  105 107 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=60.68 //y=0 //x2=61.79 //y2=0
r1545 (  103 398 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.57 //y=0 //x2=59.57 //y2=0
r1546 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.57 //y=0 //x2=60.68 //y2=0
r1547 (  101 390 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.46 //y=0 //x2=58.46 //y2=0
r1548 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.46 //y=0 //x2=59.57 //y2=0
r1549 (  99 384 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.98 //y=0 //x2=56.98 //y2=0
r1550 (  99 101 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.98 //y=0 //x2=58.46 //y2=0
r1551 (  97 382 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.87 //y=0 //x2=55.87 //y2=0
r1552 (  97 99 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.87 //y=0 //x2=56.98 //y2=0
r1553 (  95 380 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.76 //y=0 //x2=54.76 //y2=0
r1554 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.76 //y=0 //x2=55.87 //y2=0
r1555 (  93 372 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.65 //y=0 //x2=53.65 //y2=0
r1556 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=53.65 //y=0 //x2=54.76 //y2=0
r1557 (  91 366 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=52.17 //y=0 //x2=52.17 //y2=0
r1558 (  91 93 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=52.17 //y=0 //x2=53.65 //y2=0
r1559 (  89 364 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.06 //y=0 //x2=51.06 //y2=0
r1560 (  89 91 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=51.06 //y=0 //x2=52.17 //y2=0
r1561 (  87 362 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.95 //y=0 //x2=49.95 //y2=0
r1562 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.95 //y=0 //x2=51.06 //y2=0
r1563 (  84 354 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.84 //y=0 //x2=48.84 //y2=0
r1564 (  82 348 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=47.36 //y=0 //x2=47.36 //y2=0
r1565 (  82 84 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=47.36 //y=0 //x2=48.84 //y2=0
r1566 (  80 346 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.25 //y=0 //x2=46.25 //y2=0
r1567 (  80 82 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.25 //y=0 //x2=47.36 //y2=0
r1568 (  78 344 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.14 //y=0 //x2=45.14 //y2=0
r1569 (  78 80 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.14 //y=0 //x2=46.25 //y2=0
r1570 (  76 336 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.03 //y=0 //x2=44.03 //y2=0
r1571 (  76 78 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.03 //y=0 //x2=45.14 //y2=0
r1572 (  74 330 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.55 //y=0 //x2=42.55 //y2=0
r1573 (  74 76 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=42.55 //y=0 //x2=44.03 //y2=0
r1574 (  72 328 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.44 //y=0 //x2=41.44 //y2=0
r1575 (  72 74 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.44 //y=0 //x2=42.55 //y2=0
r1576 (  70 326 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=40.33 //y=0 //x2=40.33 //y2=0
r1577 (  70 72 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=40.33 //y=0 //x2=41.44 //y2=0
r1578 (  68 318 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.22 //y=0 //x2=39.22 //y2=0
r1579 (  68 70 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=39.22 //y=0 //x2=40.33 //y2=0
r1580 (  66 312 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37.74 //y=0 //x2=37.74 //y2=0
r1581 (  66 68 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=37.74 //y=0 //x2=39.22 //y2=0
r1582 (  64 310 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=36.63 //y=0 //x2=36.63 //y2=0
r1583 (  64 66 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=36.63 //y=0 //x2=37.74 //y2=0
r1584 (  62 308 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.52 //y=0 //x2=35.52 //y2=0
r1585 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.52 //y=0 //x2=36.63 //y2=0
r1586 (  60 300 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.41 //y=0 //x2=34.41 //y2=0
r1587 (  60 62 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.41 //y=0 //x2=35.52 //y2=0
r1588 (  58 294 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.93 //y=0 //x2=32.93 //y2=0
r1589 (  58 60 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.93 //y=0 //x2=34.41 //y2=0
r1590 (  56 292 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.82 //y=0 //x2=31.82 //y2=0
r1591 (  56 58 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.82 //y=0 //x2=32.93 //y2=0
r1592 (  54 290 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=30.71 //y=0 //x2=30.71 //y2=0
r1593 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=30.71 //y=0 //x2=31.82 //y2=0
r1594 (  52 282 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.6 //y=0 //x2=29.6 //y2=0
r1595 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=29.6 //y=0 //x2=30.71 //y2=0
r1596 (  50 276 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.12 //y=0 //x2=28.12 //y2=0
r1597 (  50 52 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=28.12 //y=0 //x2=29.6 //y2=0
r1598 (  48 274 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.01 //y=0 //x2=27.01 //y2=0
r1599 (  48 50 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.01 //y=0 //x2=28.12 //y2=0
r1600 (  46 272 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.9 //y=0 //x2=25.9 //y2=0
r1601 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.9 //y=0 //x2=27.01 //y2=0
r1602 (  44 264 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=0 //x2=24.79 //y2=0
r1603 (  44 46 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=0 //x2=25.9 //y2=0
r1604 (  42 258 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.31 //y=0 //x2=23.31 //y2=0
r1605 (  42 44 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.31 //y=0 //x2=24.79 //y2=0
r1606 (  40 256 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=0 //x2=22.2 //y2=0
r1607 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=0 //x2=23.31 //y2=0
r1608 (  38 254 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r1609 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=0 //x2=22.2 //y2=0
r1610 (  36 246 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=0 //x2=19.98 //y2=0
r1611 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=0 //x2=21.09 //y2=0
r1612 (  34 240 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=0 //x2=18.5 //y2=0
r1613 (  34 36 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=0 //x2=19.98 //y2=0
r1614 (  32 238 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=0 //x2=17.39 //y2=0
r1615 (  32 34 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=0 //x2=18.5 //y2=0
r1616 (  30 236 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=0 //x2=16.28 //y2=0
r1617 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=0 //x2=17.39 //y2=0
r1618 (  28 228 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r1619 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.28 //y2=0
r1620 (  26 222 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=0 //x2=13.69 //y2=0
r1621 (  26 28 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=0 //x2=15.17 //y2=0
r1622 (  24 220 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r1623 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=0 //x2=13.69 //y2=0
r1624 (  22 218 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r1625 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=0 //x2=12.58 //y2=0
r1626 (  20 210 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r1627 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r1628 (  18 204 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=0 //x2=8.88 //y2=0
r1629 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=0 //x2=10.36 //y2=0
r1630 (  16 202 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r1631 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=8.88 //y2=0
r1632 (  14 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r1633 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r1634 (  12 192 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r1635 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r1636 (  10 186 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r1637 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r1638 (  8 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r1639 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r1640 (  6 182 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r1641 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r1642 (  3 174 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r1643 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r1644 (  1 87 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=49.395 //y=0 //x2=49.95 //y2=0
r1645 (  1 84 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=49.395 //y=0 //x2=48.84 //y2=0
ends PM_TMRDFFSNRNQX1\%GND

subckt PM_TMRDFFSNRNQX1\%VDD ( 1 167 171 174 181 191 199 209 215 225 235 243 \
 253 259 269 279 287 297 303 313 323 331 341 347 357 367 375 385 391 401 411 \
 419 429 435 445 455 463 473 479 489 499 507 517 523 533 543 551 561 567 577 \
 587 595 605 611 621 631 639 649 655 665 675 683 693 699 709 719 727 737 743 \
 753 763 771 781 787 797 807 815 825 831 841 851 859 869 875 885 895 903 913 \
 919 929 939 947 957 963 971 979 989 995 1003 1013 1021 1037 1042 1047 1052 \
 1057 1062 1067 1072 1077 1082 1087 1092 1097 1102 1107 1112 1117 1122 1127 \
 1128 1129 1133 1134 1135 1136 1137 1138 1139 1140 1141 1142 1143 1144 1145 \
 1146 1147 1148 1149 1150 1151 1152 1153 1154 1155 1156 1157 1158 1159 1160 \
 1161 1162 1163 1164 1165 1166 1167 1168 1169 1170 1171 1172 1173 1174 1175 \
 1176 1177 1178 1179 1180 1181 1182 1183 1184 1185 1186 1187 1188 1189 1190 \
 1191 1192 1193 1194 1195 1196 1197 1198 1199 1200 1201 1202 1203 1204 1205 \
 1206 1207 1208 1209 1210 )
c1196 ( 1210 0 ) capacitor c=0.0433929f //x=97.98 //y=5.02
c1197 ( 1209 0 ) capacitor c=0.0420333f //x=97.11 //y=5.02
c1198 ( 1208 0 ) capacitor c=0.0476806f //x=88.985 //y=5.025
c1199 ( 1207 0 ) capacitor c=0.0241714f //x=88.105 //y=5.025
c1200 ( 1206 0 ) capacitor c=0.0467094f //x=87.235 //y=5.025
c1201 ( 1205 0 ) capacitor c=0.0452179f //x=85.355 //y=5.02
c1202 ( 1204 0 ) capacitor c=0.024152f //x=84.475 //y=5.02
c1203 ( 1203 0 ) capacitor c=0.024152f //x=83.595 //y=5.02
c1204 ( 1202 0 ) capacitor c=0.053132f //x=82.725 //y=5.02
c1205 ( 1201 0 ) capacitor c=0.0452179f //x=80.545 //y=5.02
c1206 ( 1200 0 ) capacitor c=0.024152f //x=79.665 //y=5.02
c1207 ( 1199 0 ) capacitor c=0.024152f //x=78.785 //y=5.02
c1208 ( 1198 0 ) capacitor c=0.053132f //x=77.915 //y=5.02
c1209 ( 1197 0 ) capacitor c=0.0452179f //x=75.735 //y=5.02
c1210 ( 1196 0 ) capacitor c=0.0240372f //x=74.855 //y=5.02
c1211 ( 1195 0 ) capacitor c=0.0240372f //x=73.975 //y=5.02
c1212 ( 1194 0 ) capacitor c=0.0530795f //x=73.105 //y=5.02
c1213 ( 1193 0 ) capacitor c=0.0451031f //x=70.925 //y=5.02
c1214 ( 1192 0 ) capacitor c=0.0240372f //x=70.045 //y=5.02
c1215 ( 1191 0 ) capacitor c=0.0240372f //x=69.165 //y=5.02
c1216 ( 1190 0 ) capacitor c=0.0530795f //x=68.295 //y=5.02
c1217 ( 1189 0 ) capacitor c=0.0451031f //x=66.115 //y=5.02
c1218 ( 1188 0 ) capacitor c=0.0240372f //x=65.235 //y=5.02
c1219 ( 1187 0 ) capacitor c=0.0240372f //x=64.355 //y=5.02
c1220 ( 1186 0 ) capacitor c=0.0530795f //x=63.485 //y=5.02
c1221 ( 1185 0 ) capacitor c=0.0451031f //x=61.305 //y=5.02
c1222 ( 1184 0 ) capacitor c=0.0240372f //x=60.425 //y=5.02
c1223 ( 1183 0 ) capacitor c=0.0240372f //x=59.545 //y=5.02
c1224 ( 1182 0 ) capacitor c=0.0530795f //x=58.675 //y=5.02
c1225 ( 1181 0 ) capacitor c=0.0451031f //x=56.495 //y=5.02
c1226 ( 1180 0 ) capacitor c=0.0240372f //x=55.615 //y=5.02
c1227 ( 1179 0 ) capacitor c=0.0240372f //x=54.735 //y=5.02
c1228 ( 1178 0 ) capacitor c=0.0530795f //x=53.865 //y=5.02
c1229 ( 1177 0 ) capacitor c=0.0451031f //x=51.685 //y=5.02
c1230 ( 1176 0 ) capacitor c=0.0240372f //x=50.805 //y=5.02
c1231 ( 1175 0 ) capacitor c=0.0240372f //x=49.925 //y=5.02
c1232 ( 1174 0 ) capacitor c=0.0530795f //x=49.055 //y=5.02
c1233 ( 1173 0 ) capacitor c=0.0451031f //x=46.875 //y=5.02
c1234 ( 1172 0 ) capacitor c=0.0240372f //x=45.995 //y=5.02
c1235 ( 1171 0 ) capacitor c=0.0240372f //x=45.115 //y=5.02
c1236 ( 1170 0 ) capacitor c=0.0530795f //x=44.245 //y=5.02
c1237 ( 1169 0 ) capacitor c=0.0451031f //x=42.065 //y=5.02
c1238 ( 1168 0 ) capacitor c=0.0240372f //x=41.185 //y=5.02
c1239 ( 1167 0 ) capacitor c=0.0240372f //x=40.305 //y=5.02
c1240 ( 1166 0 ) capacitor c=0.0530795f //x=39.435 //y=5.02
c1241 ( 1165 0 ) capacitor c=0.0451031f //x=37.255 //y=5.02
c1242 ( 1164 0 ) capacitor c=0.0240372f //x=36.375 //y=5.02
c1243 ( 1163 0 ) capacitor c=0.0240372f //x=35.495 //y=5.02
c1244 ( 1162 0 ) capacitor c=0.0530795f //x=34.625 //y=5.02
c1245 ( 1161 0 ) capacitor c=0.0451031f //x=32.445 //y=5.02
c1246 ( 1160 0 ) capacitor c=0.0240372f //x=31.565 //y=5.02
c1247 ( 1159 0 ) capacitor c=0.0240372f //x=30.685 //y=5.02
c1248 ( 1158 0 ) capacitor c=0.0530795f //x=29.815 //y=5.02
c1249 ( 1157 0 ) capacitor c=0.0452179f //x=27.635 //y=5.02
c1250 ( 1156 0 ) capacitor c=0.024152f //x=26.755 //y=5.02
c1251 ( 1155 0 ) capacitor c=0.024152f //x=25.875 //y=5.02
c1252 ( 1154 0 ) capacitor c=0.053132f //x=25.005 //y=5.02
c1253 ( 1153 0 ) capacitor c=0.0452179f //x=22.825 //y=5.02
c1254 ( 1152 0 ) capacitor c=0.024152f //x=21.945 //y=5.02
c1255 ( 1151 0 ) capacitor c=0.024152f //x=21.065 //y=5.02
c1256 ( 1150 0 ) capacitor c=0.053132f //x=20.195 //y=5.02
c1257 ( 1149 0 ) capacitor c=0.0452179f //x=18.015 //y=5.02
c1258 ( 1148 0 ) capacitor c=0.024152f //x=17.135 //y=5.02
c1259 ( 1147 0 ) capacitor c=0.024152f //x=16.255 //y=5.02
c1260 ( 1146 0 ) capacitor c=0.053132f //x=15.385 //y=5.02
c1261 ( 1145 0 ) capacitor c=0.0452179f //x=13.205 //y=5.02
c1262 ( 1144 0 ) capacitor c=0.024152f //x=12.325 //y=5.02
c1263 ( 1143 0 ) capacitor c=0.024152f //x=11.445 //y=5.02
c1264 ( 1142 0 ) capacitor c=0.053132f //x=10.575 //y=5.02
c1265 ( 1141 0 ) capacitor c=0.0452179f //x=8.395 //y=5.02
c1266 ( 1140 0 ) capacitor c=0.024152f //x=7.515 //y=5.02
c1267 ( 1139 0 ) capacitor c=0.02424f //x=6.635 //y=5.02
c1268 ( 1138 0 ) capacitor c=0.0531793f //x=5.765 //y=5.02
c1269 ( 1137 0 ) capacitor c=0.0453059f //x=3.585 //y=5.02
c1270 ( 1136 0 ) capacitor c=0.02424f //x=2.705 //y=5.02
c1271 ( 1135 0 ) capacitor c=0.02424f //x=1.825 //y=5.02
c1272 ( 1134 0 ) capacitor c=0.0531407f //x=0.955 //y=5.02
c1273 ( 1133 0 ) capacitor c=0.233995f //x=98.05 //y=7.4
c1274 ( 1131 0 ) capacitor c=0.00591168f //x=97.31 //y=7.4
c1275 ( 1129 0 ) capacitor c=0.107657f //x=96.57 //y=7.4
c1276 ( 1128 0 ) capacitor c=0.113329f //x=93.24 //y=7.4
c1277 ( 1127 0 ) capacitor c=0.121389f //x=89.91 //y=7.4
c1278 ( 1126 0 ) capacitor c=0.00591168f //x=89.13 //y=7.4
c1279 ( 1125 0 ) capacitor c=0.00591168f //x=88.25 //y=7.4
c1280 ( 1124 0 ) capacitor c=0.00591168f //x=87.32 //y=7.4
c1281 ( 1122 0 ) capacitor c=0.132974f //x=86.58 //y=7.4
c1282 ( 1121 0 ) capacitor c=0.00591168f //x=85.5 //y=7.4
c1283 ( 1120 0 ) capacitor c=0.00591168f //x=84.62 //y=7.4
c1284 ( 1119 0 ) capacitor c=0.00591168f //x=83.74 //y=7.4
c1285 ( 1118 0 ) capacitor c=0.00591168f //x=82.86 //y=7.4
c1286 ( 1117 0 ) capacitor c=0.155236f //x=81.77 //y=7.4
c1287 ( 1116 0 ) capacitor c=0.00591168f //x=80.69 //y=7.4
c1288 ( 1115 0 ) capacitor c=0.00591168f //x=79.81 //y=7.4
c1289 ( 1114 0 ) capacitor c=0.00591168f //x=78.93 //y=7.4
c1290 ( 1113 0 ) capacitor c=0.00591168f //x=78.05 //y=7.4
c1291 ( 1112 0 ) capacitor c=0.154686f //x=76.96 //y=7.4
c1292 ( 1111 0 ) capacitor c=0.00591168f //x=75.88 //y=7.4
c1293 ( 1110 0 ) capacitor c=0.00591168f //x=75 //y=7.4
c1294 ( 1109 0 ) capacitor c=0.00591168f //x=74.12 //y=7.4
c1295 ( 1108 0 ) capacitor c=0.00591168f //x=73.24 //y=7.4
c1296 ( 1107 0 ) capacitor c=0.153722f //x=72.15 //y=7.4
c1297 ( 1106 0 ) capacitor c=0.00591168f //x=71.07 //y=7.4
c1298 ( 1105 0 ) capacitor c=0.00591168f //x=70.19 //y=7.4
c1299 ( 1104 0 ) capacitor c=0.00591168f //x=69.31 //y=7.4
c1300 ( 1103 0 ) capacitor c=0.00591168f //x=68.43 //y=7.4
c1301 ( 1102 0 ) capacitor c=0.153803f //x=67.34 //y=7.4
c1302 ( 1101 0 ) capacitor c=0.00591168f //x=66.26 //y=7.4
c1303 ( 1100 0 ) capacitor c=0.00591168f //x=65.38 //y=7.4
c1304 ( 1099 0 ) capacitor c=0.00591168f //x=64.5 //y=7.4
c1305 ( 1098 0 ) capacitor c=0.00591168f //x=63.62 //y=7.4
c1306 ( 1097 0 ) capacitor c=0.158289f //x=62.53 //y=7.4
c1307 ( 1096 0 ) capacitor c=0.00591168f //x=61.45 //y=7.4
c1308 ( 1095 0 ) capacitor c=0.00591168f //x=60.57 //y=7.4
c1309 ( 1094 0 ) capacitor c=0.00591168f //x=59.69 //y=7.4
c1310 ( 1093 0 ) capacitor c=0.00591168f //x=58.81 //y=7.4
c1311 ( 1092 0 ) capacitor c=0.15374f //x=57.72 //y=7.4
c1312 ( 1091 0 ) capacitor c=0.00591168f //x=56.64 //y=7.4
c1313 ( 1090 0 ) capacitor c=0.00591168f //x=55.76 //y=7.4
c1314 ( 1089 0 ) capacitor c=0.00591168f //x=54.88 //y=7.4
c1315 ( 1088 0 ) capacitor c=0.00591168f //x=54 //y=7.4
c1316 ( 1087 0 ) capacitor c=0.15385f //x=52.91 //y=7.4
c1317 ( 1086 0 ) capacitor c=0.00591168f //x=51.83 //y=7.4
c1318 ( 1085 0 ) capacitor c=0.00591168f //x=50.95 //y=7.4
c1319 ( 1084 0 ) capacitor c=0.00591168f //x=50.07 //y=7.4
c1320 ( 1083 0 ) capacitor c=0.00591168f //x=49.19 //y=7.4
c1321 ( 1082 0 ) capacitor c=0.153803f //x=48.1 //y=7.4
c1322 ( 1081 0 ) capacitor c=0.00591168f //x=47.02 //y=7.4
c1323 ( 1080 0 ) capacitor c=0.00591168f //x=46.14 //y=7.4
c1324 ( 1079 0 ) capacitor c=0.00591168f //x=45.26 //y=7.4
c1325 ( 1078 0 ) capacitor c=0.00591168f //x=44.38 //y=7.4
c1326 ( 1077 0 ) capacitor c=0.153779f //x=43.29 //y=7.4
c1327 ( 1076 0 ) capacitor c=0.00591168f //x=42.21 //y=7.4
c1328 ( 1075 0 ) capacitor c=0.00591168f //x=41.33 //y=7.4
c1329 ( 1074 0 ) capacitor c=0.00591168f //x=40.45 //y=7.4
c1330 ( 1073 0 ) capacitor c=0.00591168f //x=39.57 //y=7.4
c1331 ( 1072 0 ) capacitor c=0.153803f //x=38.48 //y=7.4
c1332 ( 1071 0 ) capacitor c=0.00591168f //x=37.4 //y=7.4
c1333 ( 1070 0 ) capacitor c=0.00591168f //x=36.52 //y=7.4
c1334 ( 1069 0 ) capacitor c=0.00591168f //x=35.64 //y=7.4
c1335 ( 1068 0 ) capacitor c=0.00591168f //x=34.76 //y=7.4
c1336 ( 1067 0 ) capacitor c=0.153957f //x=33.67 //y=7.4
c1337 ( 1066 0 ) capacitor c=0.00591168f //x=32.59 //y=7.4
c1338 ( 1065 0 ) capacitor c=0.00591168f //x=31.71 //y=7.4
c1339 ( 1064 0 ) capacitor c=0.00591168f //x=30.83 //y=7.4
c1340 ( 1063 0 ) capacitor c=0.00591168f //x=29.95 //y=7.4
c1341 ( 1062 0 ) capacitor c=0.153836f //x=28.86 //y=7.4
c1342 ( 1061 0 ) capacitor c=0.00591168f //x=27.78 //y=7.4
c1343 ( 1060 0 ) capacitor c=0.00591168f //x=26.9 //y=7.4
c1344 ( 1059 0 ) capacitor c=0.00591168f //x=26.02 //y=7.4
c1345 ( 1058 0 ) capacitor c=0.00591168f //x=25.14 //y=7.4
c1346 ( 1057 0 ) capacitor c=0.155236f //x=24.05 //y=7.4
c1347 ( 1056 0 ) capacitor c=0.00591168f //x=22.97 //y=7.4
c1348 ( 1055 0 ) capacitor c=0.00591168f //x=22.09 //y=7.4
c1349 ( 1054 0 ) capacitor c=0.00591168f //x=21.21 //y=7.4
c1350 ( 1053 0 ) capacitor c=0.00591168f //x=20.33 //y=7.4
c1351 ( 1052 0 ) capacitor c=0.15519f //x=19.24 //y=7.4
c1352 ( 1051 0 ) capacitor c=0.00591168f //x=18.16 //y=7.4
c1353 ( 1050 0 ) capacitor c=0.00591168f //x=17.28 //y=7.4
c1354 ( 1049 0 ) capacitor c=0.00591168f //x=16.4 //y=7.4
c1355 ( 1048 0 ) capacitor c=0.00591168f //x=15.52 //y=7.4
c1356 ( 1047 0 ) capacitor c=0.155166f //x=14.43 //y=7.4
c1357 ( 1046 0 ) capacitor c=0.00591168f //x=13.35 //y=7.4
c1358 ( 1045 0 ) capacitor c=0.00591168f //x=12.47 //y=7.4
c1359 ( 1044 0 ) capacitor c=0.00591168f //x=11.59 //y=7.4
c1360 ( 1043 0 ) capacitor c=0.00591168f //x=10.71 //y=7.4
c1361 ( 1042 0 ) capacitor c=0.15519f //x=9.62 //y=7.4
c1362 ( 1041 0 ) capacitor c=0.00591168f //x=8.54 //y=7.4
c1363 ( 1040 0 ) capacitor c=0.00591168f //x=7.66 //y=7.4
c1364 ( 1039 0 ) capacitor c=0.00591168f //x=6.78 //y=7.4
c1365 ( 1038 0 ) capacitor c=0.00591168f //x=5.9 //y=7.4
c1366 ( 1037 0 ) capacitor c=0.157289f //x=4.81 //y=7.4
c1367 ( 1036 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c1368 ( 1035 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c1369 ( 1034 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c1370 ( 1033 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c1371 ( 1021 0 ) capacitor c=0.028907f //x=98.04 //y=7.4
c1372 ( 1013 0 ) capacitor c=0.0186283f //x=97.16 //y=7.4
c1373 ( 1003 0 ) capacitor c=0.12108f //x=96.4 //y=7.4
c1374 ( 995 0 ) capacitor c=0.120978f //x=93.07 //y=7.4
c1375 ( 989 0 ) capacitor c=0.0236224f //x=89.74 //y=7.4
c1376 ( 979 0 ) capacitor c=0.028539f //x=89.045 //y=7.4
c1377 ( 971 0 ) capacitor c=0.0285075f //x=88.165 //y=7.4
c1378 ( 963 0 ) capacitor c=0.0240981f //x=87.285 //y=7.4
c1379 ( 957 0 ) capacitor c=0.0394667f //x=86.41 //y=7.4
c1380 ( 947 0 ) capacitor c=0.0288488f //x=85.415 //y=7.4
c1381 ( 939 0 ) capacitor c=0.0287514f //x=84.535 //y=7.4
c1382 ( 929 0 ) capacitor c=0.0284966f //x=83.655 //y=7.4
c1383 ( 919 0 ) capacitor c=0.0383672f //x=82.775 //y=7.4
c1384 ( 913 0 ) capacitor c=0.0394667f //x=81.6 //y=7.4
c1385 ( 903 0 ) capacitor c=0.0288488f //x=80.605 //y=7.4
c1386 ( 895 0 ) capacitor c=0.0287514f //x=79.725 //y=7.4
c1387 ( 885 0 ) capacitor c=0.0284966f //x=78.845 //y=7.4
c1388 ( 875 0 ) capacitor c=0.0383672f //x=77.965 //y=7.4
c1389 ( 869 0 ) capacitor c=0.0394667f //x=76.79 //y=7.4
c1390 ( 859 0 ) capacitor c=0.0288466f //x=75.795 //y=7.4
c1391 ( 851 0 ) capacitor c=0.028724f //x=74.915 //y=7.4
c1392 ( 841 0 ) capacitor c=0.0284804f //x=74.035 //y=7.4
c1393 ( 831 0 ) capacitor c=0.0383672f //x=73.155 //y=7.4
c1394 ( 825 0 ) capacitor c=0.0394025f //x=71.98 //y=7.4
c1395 ( 815 0 ) capacitor c=0.0288171f //x=70.985 //y=7.4
c1396 ( 807 0 ) capacitor c=0.028724f //x=70.105 //y=7.4
c1397 ( 797 0 ) capacitor c=0.0284804f //x=69.225 //y=7.4
c1398 ( 787 0 ) capacitor c=0.0383672f //x=68.345 //y=7.4
c1399 ( 781 0 ) capacitor c=0.0394025f //x=67.17 //y=7.4
c1400 ( 771 0 ) capacitor c=0.0288171f //x=66.175 //y=7.4
c1401 ( 763 0 ) capacitor c=0.028724f //x=65.295 //y=7.4
c1402 ( 753 0 ) capacitor c=0.0284804f //x=64.415 //y=7.4
c1403 ( 743 0 ) capacitor c=0.0383672f //x=63.535 //y=7.4
c1404 ( 737 0 ) capacitor c=0.0394025f //x=62.36 //y=7.4
c1405 ( 727 0 ) capacitor c=0.0288171f //x=61.365 //y=7.4
c1406 ( 719 0 ) capacitor c=0.028724f //x=60.485 //y=7.4
c1407 ( 709 0 ) capacitor c=0.0284804f //x=59.605 //y=7.4
c1408 ( 699 0 ) capacitor c=0.0383672f //x=58.725 //y=7.4
c1409 ( 693 0 ) capacitor c=0.0394025f //x=57.55 //y=7.4
c1410 ( 683 0 ) capacitor c=0.0288171f //x=56.555 //y=7.4
c1411 ( 675 0 ) capacitor c=0.028724f //x=55.675 //y=7.4
c1412 ( 665 0 ) capacitor c=0.0284804f //x=54.795 //y=7.4
c1413 ( 655 0 ) capacitor c=0.0383672f //x=53.915 //y=7.4
c1414 ( 649 0 ) capacitor c=0.0394025f //x=52.74 //y=7.4
c1415 ( 639 0 ) capacitor c=0.0288171f //x=51.745 //y=7.4
c1416 ( 631 0 ) capacitor c=0.028724f //x=50.865 //y=7.4
c1417 ( 621 0 ) capacitor c=0.0284804f //x=49.985 //y=7.4
c1418 ( 611 0 ) capacitor c=0.0383672f //x=49.105 //y=7.4
c1419 ( 605 0 ) capacitor c=0.0394025f //x=47.93 //y=7.4
c1420 ( 595 0 ) capacitor c=0.0288171f //x=46.935 //y=7.4
c1421 ( 587 0 ) capacitor c=0.028724f //x=46.055 //y=7.4
c1422 ( 577 0 ) capacitor c=0.0284804f //x=45.175 //y=7.4
c1423 ( 567 0 ) capacitor c=0.0383672f //x=44.295 //y=7.4
c1424 ( 561 0 ) capacitor c=0.0394025f //x=43.12 //y=7.4
c1425 ( 551 0 ) capacitor c=0.0288171f //x=42.125 //y=7.4
c1426 ( 543 0 ) capacitor c=0.028724f //x=41.245 //y=7.4
c1427 ( 533 0 ) capacitor c=0.0284804f //x=40.365 //y=7.4
c1428 ( 523 0 ) capacitor c=0.0383672f //x=39.485 //y=7.4
c1429 ( 517 0 ) capacitor c=0.0394025f //x=38.31 //y=7.4
c1430 ( 507 0 ) capacitor c=0.0288171f //x=37.315 //y=7.4
c1431 ( 499 0 ) capacitor c=0.028724f //x=36.435 //y=7.4
c1432 ( 489 0 ) capacitor c=0.0284804f //x=35.555 //y=7.4
c1433 ( 479 0 ) capacitor c=0.0383672f //x=34.675 //y=7.4
c1434 ( 473 0 ) capacitor c=0.0394025f //x=33.5 //y=7.4
c1435 ( 463 0 ) capacitor c=0.0288171f //x=32.505 //y=7.4
c1436 ( 455 0 ) capacitor c=0.028724f //x=31.625 //y=7.4
c1437 ( 445 0 ) capacitor c=0.0284804f //x=30.745 //y=7.4
c1438 ( 435 0 ) capacitor c=0.0383672f //x=29.865 //y=7.4
c1439 ( 429 0 ) capacitor c=0.0394119f //x=28.69 //y=7.4
c1440 ( 419 0 ) capacitor c=0.0288488f //x=27.695 //y=7.4
c1441 ( 411 0 ) capacitor c=0.0287514f //x=26.815 //y=7.4
c1442 ( 401 0 ) capacitor c=0.0284966f //x=25.935 //y=7.4
c1443 ( 391 0 ) capacitor c=0.0383672f //x=25.055 //y=7.4
c1444 ( 385 0 ) capacitor c=0.0394667f //x=23.88 //y=7.4
c1445 ( 375 0 ) capacitor c=0.0288488f //x=22.885 //y=7.4
c1446 ( 367 0 ) capacitor c=0.0287514f //x=22.005 //y=7.4
c1447 ( 357 0 ) capacitor c=0.0284966f //x=21.125 //y=7.4
c1448 ( 347 0 ) capacitor c=0.0383672f //x=20.245 //y=7.4
c1449 ( 341 0 ) capacitor c=0.0394667f //x=19.07 //y=7.4
c1450 ( 331 0 ) capacitor c=0.0288488f //x=18.075 //y=7.4
c1451 ( 323 0 ) capacitor c=0.0287505f //x=17.195 //y=7.4
c1452 ( 313 0 ) capacitor c=0.0284966f //x=16.315 //y=7.4
c1453 ( 303 0 ) capacitor c=0.0383672f //x=15.435 //y=7.4
c1454 ( 297 0 ) capacitor c=0.0394667f //x=14.26 //y=7.4
c1455 ( 287 0 ) capacitor c=0.0288488f //x=13.265 //y=7.4
c1456 ( 279 0 ) capacitor c=0.0287514f //x=12.385 //y=7.4
c1457 ( 269 0 ) capacitor c=0.0284966f //x=11.505 //y=7.4
c1458 ( 259 0 ) capacitor c=0.0383672f //x=10.625 //y=7.4
c1459 ( 253 0 ) capacitor c=0.0394667f //x=9.45 //y=7.4
c1460 ( 243 0 ) capacitor c=0.0288488f //x=8.455 //y=7.4
c1461 ( 235 0 ) capacitor c=0.0287505f //x=7.575 //y=7.4
c1462 ( 225 0 ) capacitor c=0.028511f //x=6.695 //y=7.4
c1463 ( 215 0 ) capacitor c=0.0383672f //x=5.815 //y=7.4
c1464 ( 209 0 ) capacitor c=0.0395236f //x=4.64 //y=7.4
c1465 ( 199 0 ) capacitor c=0.0288769f //x=3.645 //y=7.4
c1466 ( 191 0 ) capacitor c=0.0287757f //x=2.765 //y=7.4
c1467 ( 181 0 ) capacitor c=0.028511f //x=1.885 //y=7.4
c1468 ( 174 0 ) capacitor c=0.234727f //x=0.74 //y=7.4
c1469 ( 171 0 ) capacitor c=0.0441843f //x=1.005 //y=7.4
c1470 ( 167 0 ) capacitor c=3.25525f //x=98.05 //y=7.4
r1471 (  1023 1133 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=98.125 //y=7.23 //x2=98.125 //y2=7.4
r1472 (  1023 1210 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=98.125 //y=7.23 //x2=98.125 //y2=6.405
r1473 (  1022 1131 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=97.33 //y=7.4 //x2=97.245 //y2=7.4
r1474 (  1021 1133 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=98.04 //y=7.4 //x2=98.125 //y2=7.4
r1475 (  1021 1022 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=98.04 //y=7.4 //x2=97.33 //y2=7.4
r1476 (  1015 1131 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=97.245 //y=7.23 //x2=97.245 //y2=7.4
r1477 (  1015 1209 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=97.245 //y=7.23 //x2=97.245 //y2=6.405
r1478 (  1014 1129 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=96.74 //y=7.4 //x2=96.57 //y2=7.4
r1479 (  1013 1131 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=97.16 //y=7.4 //x2=97.245 //y2=7.4
r1480 (  1013 1014 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=97.16 //y=7.4 //x2=96.74 //y2=7.4
r1481 (  1008 1010 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=94.72 //y=7.4 //x2=95.83 //y2=7.4
r1482 (  1006 1008 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=93.61 //y=7.4 //x2=94.72 //y2=7.4
r1483 (  1004 1128 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=93.41 //y=7.4 //x2=93.24 //y2=7.4
r1484 (  1004 1006 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=93.41 //y=7.4 //x2=93.61 //y2=7.4
r1485 (  1003 1129 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=96.4 //y=7.4 //x2=96.57 //y2=7.4
r1486 (  1003 1010 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=96.4 //y=7.4 //x2=95.83 //y2=7.4
r1487 (  998 1000 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=91.02 //y=7.4 //x2=92.13 //y2=7.4
r1488 (  996 1127 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=90.08 //y=7.4 //x2=89.91 //y2=7.4
r1489 (  996 998 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=90.08 //y=7.4 //x2=91.02 //y2=7.4
r1490 (  995 1128 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=93.07 //y=7.4 //x2=93.24 //y2=7.4
r1491 (  995 1000 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=93.07 //y=7.4 //x2=92.13 //y2=7.4
r1492 (  990 1126 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=89.215 //y=7.4 //x2=89.13 //y2=7.4
r1493 (  990 992 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=89.215 //y=7.4 //x2=89.54 //y2=7.4
r1494 (  989 1127 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=89.74 //y=7.4 //x2=89.91 //y2=7.4
r1495 (  989 992 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=89.74 //y=7.4 //x2=89.54 //y2=7.4
r1496 (  983 1126 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=89.13 //y=7.23 //x2=89.13 //y2=7.4
r1497 (  983 1208 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=89.13 //y=7.23 //x2=89.13 //y2=6.4
r1498 (  980 1125 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=88.335 //y=7.4 //x2=88.25 //y2=7.4
r1499 (  980 982 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=88.335 //y=7.4 //x2=88.43 //y2=7.4
r1500 (  979 1126 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=89.045 //y=7.4 //x2=89.13 //y2=7.4
r1501 (  979 982 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=89.045 //y=7.4 //x2=88.43 //y2=7.4
r1502 (  973 1125 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=88.25 //y=7.23 //x2=88.25 //y2=7.4
r1503 (  973 1207 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=88.25 //y=7.23 //x2=88.25 //y2=6.74
r1504 (  972 1124 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=87.455 //y=7.4 //x2=87.37 //y2=7.4
r1505 (  971 1125 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=88.165 //y=7.4 //x2=88.25 //y2=7.4
r1506 (  971 972 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=88.165 //y=7.4 //x2=87.455 //y2=7.4
r1507 (  965 1124 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=87.37 //y=7.23 //x2=87.37 //y2=7.4
r1508 (  965 1206 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=87.37 //y=7.23 //x2=87.37 //y2=6.4
r1509 (  964 1122 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=86.75 //y=7.4 //x2=86.58 //y2=7.4
r1510 (  963 1124 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=87.285 //y=7.4 //x2=87.37 //y2=7.4
r1511 (  963 964 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=87.285 //y=7.4 //x2=86.75 //y2=7.4
r1512 (  958 1121 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.585 //y=7.4 //x2=85.5 //y2=7.4
r1513 (  958 960 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=85.585 //y=7.4 //x2=85.84 //y2=7.4
r1514 (  957 1122 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=86.41 //y=7.4 //x2=86.58 //y2=7.4
r1515 (  957 960 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=86.41 //y=7.4 //x2=85.84 //y2=7.4
r1516 (  951 1121 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=85.5 //y=7.23 //x2=85.5 //y2=7.4
r1517 (  951 1205 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=85.5 //y=7.23 //x2=85.5 //y2=6.745
r1518 (  948 1120 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.705 //y=7.4 //x2=84.62 //y2=7.4
r1519 (  948 950 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=84.705 //y=7.4 //x2=84.73 //y2=7.4
r1520 (  947 1121 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.415 //y=7.4 //x2=85.5 //y2=7.4
r1521 (  947 950 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=85.415 //y=7.4 //x2=84.73 //y2=7.4
r1522 (  941 1120 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=84.62 //y=7.23 //x2=84.62 //y2=7.4
r1523 (  941 1204 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=84.62 //y=7.23 //x2=84.62 //y2=6.745
r1524 (  940 1119 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.825 //y=7.4 //x2=83.74 //y2=7.4
r1525 (  939 1120 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.535 //y=7.4 //x2=84.62 //y2=7.4
r1526 (  939 940 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=84.535 //y=7.4 //x2=83.825 //y2=7.4
r1527 (  933 1119 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=83.74 //y=7.23 //x2=83.74 //y2=7.4
r1528 (  933 1203 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=83.74 //y=7.23 //x2=83.74 //y2=6.745
r1529 (  930 1118 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.945 //y=7.4 //x2=82.86 //y2=7.4
r1530 (  930 932 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=82.945 //y=7.4 //x2=83.62 //y2=7.4
r1531 (  929 1119 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.655 //y=7.4 //x2=83.74 //y2=7.4
r1532 (  929 932 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=83.655 //y=7.4 //x2=83.62 //y2=7.4
r1533 (  923 1118 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=82.86 //y=7.23 //x2=82.86 //y2=7.4
r1534 (  923 1202 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=82.86 //y=7.23 //x2=82.86 //y2=6.405
r1535 (  920 1117 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.94 //y=7.4 //x2=81.77 //y2=7.4
r1536 (  920 922 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=81.94 //y=7.4 //x2=82.51 //y2=7.4
r1537 (  919 1118 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.775 //y=7.4 //x2=82.86 //y2=7.4
r1538 (  919 922 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=82.775 //y=7.4 //x2=82.51 //y2=7.4
r1539 (  914 1116 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.775 //y=7.4 //x2=80.69 //y2=7.4
r1540 (  914 916 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=80.775 //y=7.4 //x2=81.03 //y2=7.4
r1541 (  913 1117 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.6 //y=7.4 //x2=81.77 //y2=7.4
r1542 (  913 916 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=81.6 //y=7.4 //x2=81.03 //y2=7.4
r1543 (  907 1116 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=80.69 //y=7.23 //x2=80.69 //y2=7.4
r1544 (  907 1201 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=80.69 //y=7.23 //x2=80.69 //y2=6.745
r1545 (  904 1115 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.895 //y=7.4 //x2=79.81 //y2=7.4
r1546 (  904 906 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=79.895 //y=7.4 //x2=79.92 //y2=7.4
r1547 (  903 1116 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.605 //y=7.4 //x2=80.69 //y2=7.4
r1548 (  903 906 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=80.605 //y=7.4 //x2=79.92 //y2=7.4
r1549 (  897 1115 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=79.81 //y=7.23 //x2=79.81 //y2=7.4
r1550 (  897 1200 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=79.81 //y=7.23 //x2=79.81 //y2=6.745
r1551 (  896 1114 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.015 //y=7.4 //x2=78.93 //y2=7.4
r1552 (  895 1115 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.725 //y=7.4 //x2=79.81 //y2=7.4
r1553 (  895 896 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=79.725 //y=7.4 //x2=79.015 //y2=7.4
r1554 (  889 1114 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=78.93 //y=7.23 //x2=78.93 //y2=7.4
r1555 (  889 1199 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=78.93 //y=7.23 //x2=78.93 //y2=6.745
r1556 (  886 1113 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.135 //y=7.4 //x2=78.05 //y2=7.4
r1557 (  886 888 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=78.135 //y=7.4 //x2=78.81 //y2=7.4
r1558 (  885 1114 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.845 //y=7.4 //x2=78.93 //y2=7.4
r1559 (  885 888 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=78.845 //y=7.4 //x2=78.81 //y2=7.4
r1560 (  879 1113 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=78.05 //y=7.23 //x2=78.05 //y2=7.4
r1561 (  879 1198 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=78.05 //y=7.23 //x2=78.05 //y2=6.405
r1562 (  876 1112 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.13 //y=7.4 //x2=76.96 //y2=7.4
r1563 (  876 878 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=77.13 //y=7.4 //x2=77.7 //y2=7.4
r1564 (  875 1113 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.965 //y=7.4 //x2=78.05 //y2=7.4
r1565 (  875 878 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=77.965 //y=7.4 //x2=77.7 //y2=7.4
r1566 (  870 1111 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.965 //y=7.4 //x2=75.88 //y2=7.4
r1567 (  870 872 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=75.965 //y=7.4 //x2=76.22 //y2=7.4
r1568 (  869 1112 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.79 //y=7.4 //x2=76.96 //y2=7.4
r1569 (  869 872 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=76.79 //y=7.4 //x2=76.22 //y2=7.4
r1570 (  863 1111 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=75.88 //y=7.23 //x2=75.88 //y2=7.4
r1571 (  863 1197 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=75.88 //y=7.23 //x2=75.88 //y2=6.745
r1572 (  860 1110 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.085 //y=7.4 //x2=75 //y2=7.4
r1573 (  860 862 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=75.085 //y=7.4 //x2=75.11 //y2=7.4
r1574 (  859 1111 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.795 //y=7.4 //x2=75.88 //y2=7.4
r1575 (  859 862 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=75.795 //y=7.4 //x2=75.11 //y2=7.4
r1576 (  853 1110 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=75 //y=7.23 //x2=75 //y2=7.4
r1577 (  853 1196 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=75 //y=7.23 //x2=75 //y2=6.745
r1578 (  852 1109 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.205 //y=7.4 //x2=74.12 //y2=7.4
r1579 (  851 1110 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.915 //y=7.4 //x2=75 //y2=7.4
r1580 (  851 852 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=74.915 //y=7.4 //x2=74.205 //y2=7.4
r1581 (  845 1109 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.12 //y=7.23 //x2=74.12 //y2=7.4
r1582 (  845 1195 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=74.12 //y=7.23 //x2=74.12 //y2=6.745
r1583 (  842 1108 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.325 //y=7.4 //x2=73.24 //y2=7.4
r1584 (  842 844 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=73.325 //y=7.4 //x2=74 //y2=7.4
r1585 (  841 1109 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.035 //y=7.4 //x2=74.12 //y2=7.4
r1586 (  841 844 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=74.035 //y=7.4 //x2=74 //y2=7.4
r1587 (  835 1108 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.24 //y=7.23 //x2=73.24 //y2=7.4
r1588 (  835 1194 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=73.24 //y=7.23 //x2=73.24 //y2=6.405
r1589 (  832 1107 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=72.32 //y=7.4 //x2=72.15 //y2=7.4
r1590 (  832 834 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=72.32 //y=7.4 //x2=72.89 //y2=7.4
r1591 (  831 1108 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.155 //y=7.4 //x2=73.24 //y2=7.4
r1592 (  831 834 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=73.155 //y=7.4 //x2=72.89 //y2=7.4
r1593 (  826 1106 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.155 //y=7.4 //x2=71.07 //y2=7.4
r1594 (  826 828 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=71.155 //y=7.4 //x2=71.41 //y2=7.4
r1595 (  825 1107 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.98 //y=7.4 //x2=72.15 //y2=7.4
r1596 (  825 828 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=71.98 //y=7.4 //x2=71.41 //y2=7.4
r1597 (  819 1106 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.07 //y=7.23 //x2=71.07 //y2=7.4
r1598 (  819 1193 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=71.07 //y=7.23 //x2=71.07 //y2=6.745
r1599 (  816 1105 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.275 //y=7.4 //x2=70.19 //y2=7.4
r1600 (  816 818 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=70.275 //y=7.4 //x2=70.3 //y2=7.4
r1601 (  815 1106 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.985 //y=7.4 //x2=71.07 //y2=7.4
r1602 (  815 818 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=70.985 //y=7.4 //x2=70.3 //y2=7.4
r1603 (  809 1105 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=70.19 //y=7.23 //x2=70.19 //y2=7.4
r1604 (  809 1192 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=70.19 //y=7.23 //x2=70.19 //y2=6.745
r1605 (  808 1104 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.395 //y=7.4 //x2=69.31 //y2=7.4
r1606 (  807 1105 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.105 //y=7.4 //x2=70.19 //y2=7.4
r1607 (  807 808 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=70.105 //y=7.4 //x2=69.395 //y2=7.4
r1608 (  801 1104 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.31 //y=7.23 //x2=69.31 //y2=7.4
r1609 (  801 1191 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=69.31 //y=7.23 //x2=69.31 //y2=6.745
r1610 (  798 1103 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.515 //y=7.4 //x2=68.43 //y2=7.4
r1611 (  798 800 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=68.515 //y=7.4 //x2=69.19 //y2=7.4
r1612 (  797 1104 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.225 //y=7.4 //x2=69.31 //y2=7.4
r1613 (  797 800 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=69.225 //y=7.4 //x2=69.19 //y2=7.4
r1614 (  791 1103 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.43 //y=7.23 //x2=68.43 //y2=7.4
r1615 (  791 1190 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=68.43 //y=7.23 //x2=68.43 //y2=6.405
r1616 (  788 1102 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.51 //y=7.4 //x2=67.34 //y2=7.4
r1617 (  788 790 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.51 //y=7.4 //x2=68.08 //y2=7.4
r1618 (  787 1103 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.345 //y=7.4 //x2=68.43 //y2=7.4
r1619 (  787 790 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=68.345 //y=7.4 //x2=68.08 //y2=7.4
r1620 (  782 1101 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.345 //y=7.4 //x2=66.26 //y2=7.4
r1621 (  782 784 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=66.345 //y=7.4 //x2=66.6 //y2=7.4
r1622 (  781 1102 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.17 //y=7.4 //x2=67.34 //y2=7.4
r1623 (  781 784 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.17 //y=7.4 //x2=66.6 //y2=7.4
r1624 (  775 1101 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=66.26 //y=7.23 //x2=66.26 //y2=7.4
r1625 (  775 1189 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=66.26 //y=7.23 //x2=66.26 //y2=6.745
r1626 (  772 1100 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.465 //y=7.4 //x2=65.38 //y2=7.4
r1627 (  772 774 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=65.465 //y=7.4 //x2=65.49 //y2=7.4
r1628 (  771 1101 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.175 //y=7.4 //x2=66.26 //y2=7.4
r1629 (  771 774 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=66.175 //y=7.4 //x2=65.49 //y2=7.4
r1630 (  765 1100 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.38 //y=7.23 //x2=65.38 //y2=7.4
r1631 (  765 1188 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=65.38 //y=7.23 //x2=65.38 //y2=6.745
r1632 (  764 1099 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.585 //y=7.4 //x2=64.5 //y2=7.4
r1633 (  763 1100 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.295 //y=7.4 //x2=65.38 //y2=7.4
r1634 (  763 764 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=65.295 //y=7.4 //x2=64.585 //y2=7.4
r1635 (  757 1099 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.5 //y=7.23 //x2=64.5 //y2=7.4
r1636 (  757 1187 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=64.5 //y=7.23 //x2=64.5 //y2=6.745
r1637 (  754 1098 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.705 //y=7.4 //x2=63.62 //y2=7.4
r1638 (  754 756 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=63.705 //y=7.4 //x2=64.38 //y2=7.4
r1639 (  753 1099 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.415 //y=7.4 //x2=64.5 //y2=7.4
r1640 (  753 756 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=64.415 //y=7.4 //x2=64.38 //y2=7.4
r1641 (  747 1098 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=63.62 //y=7.23 //x2=63.62 //y2=7.4
r1642 (  747 1186 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=63.62 //y=7.23 //x2=63.62 //y2=6.405
r1643 (  744 1097 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.7 //y=7.4 //x2=62.53 //y2=7.4
r1644 (  744 746 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=62.7 //y=7.4 //x2=63.27 //y2=7.4
r1645 (  743 1098 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.535 //y=7.4 //x2=63.62 //y2=7.4
r1646 (  743 746 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=63.535 //y=7.4 //x2=63.27 //y2=7.4
r1647 (  738 1096 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.535 //y=7.4 //x2=61.45 //y2=7.4
r1648 (  738 740 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=61.535 //y=7.4 //x2=61.79 //y2=7.4
r1649 (  737 1097 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.36 //y=7.4 //x2=62.53 //y2=7.4
r1650 (  737 740 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=62.36 //y=7.4 //x2=61.79 //y2=7.4
r1651 (  731 1096 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.45 //y=7.23 //x2=61.45 //y2=7.4
r1652 (  731 1185 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=61.45 //y=7.23 //x2=61.45 //y2=6.745
r1653 (  728 1095 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.655 //y=7.4 //x2=60.57 //y2=7.4
r1654 (  728 730 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=60.655 //y=7.4 //x2=60.68 //y2=7.4
r1655 (  727 1096 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.365 //y=7.4 //x2=61.45 //y2=7.4
r1656 (  727 730 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=61.365 //y=7.4 //x2=60.68 //y2=7.4
r1657 (  721 1095 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=60.57 //y=7.23 //x2=60.57 //y2=7.4
r1658 (  721 1184 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.57 //y=7.23 //x2=60.57 //y2=6.745
r1659 (  720 1094 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.775 //y=7.4 //x2=59.69 //y2=7.4
r1660 (  719 1095 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.485 //y=7.4 //x2=60.57 //y2=7.4
r1661 (  719 720 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=60.485 //y=7.4 //x2=59.775 //y2=7.4
r1662 (  713 1094 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=59.69 //y=7.23 //x2=59.69 //y2=7.4
r1663 (  713 1183 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.69 //y=7.23 //x2=59.69 //y2=6.745
r1664 (  710 1093 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.895 //y=7.4 //x2=58.81 //y2=7.4
r1665 (  710 712 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=58.895 //y=7.4 //x2=59.57 //y2=7.4
r1666 (  709 1094 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.605 //y=7.4 //x2=59.69 //y2=7.4
r1667 (  709 712 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=59.605 //y=7.4 //x2=59.57 //y2=7.4
r1668 (  703 1093 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.81 //y=7.23 //x2=58.81 //y2=7.4
r1669 (  703 1182 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=58.81 //y=7.23 //x2=58.81 //y2=6.405
r1670 (  700 1092 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.89 //y=7.4 //x2=57.72 //y2=7.4
r1671 (  700 702 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=57.89 //y=7.4 //x2=58.46 //y2=7.4
r1672 (  699 1093 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.725 //y=7.4 //x2=58.81 //y2=7.4
r1673 (  699 702 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=58.725 //y=7.4 //x2=58.46 //y2=7.4
r1674 (  694 1091 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.725 //y=7.4 //x2=56.64 //y2=7.4
r1675 (  694 696 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=56.725 //y=7.4 //x2=56.98 //y2=7.4
r1676 (  693 1092 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.55 //y=7.4 //x2=57.72 //y2=7.4
r1677 (  693 696 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=57.55 //y=7.4 //x2=56.98 //y2=7.4
r1678 (  687 1091 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.64 //y=7.23 //x2=56.64 //y2=7.4
r1679 (  687 1181 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=56.64 //y=7.23 //x2=56.64 //y2=6.745
r1680 (  684 1090 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.845 //y=7.4 //x2=55.76 //y2=7.4
r1681 (  684 686 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=55.845 //y=7.4 //x2=55.87 //y2=7.4
r1682 (  683 1091 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.555 //y=7.4 //x2=56.64 //y2=7.4
r1683 (  683 686 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=56.555 //y=7.4 //x2=55.87 //y2=7.4
r1684 (  677 1090 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=55.76 //y=7.23 //x2=55.76 //y2=7.4
r1685 (  677 1180 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.76 //y=7.23 //x2=55.76 //y2=6.745
r1686 (  676 1089 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.965 //y=7.4 //x2=54.88 //y2=7.4
r1687 (  675 1090 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.675 //y=7.4 //x2=55.76 //y2=7.4
r1688 (  675 676 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=55.675 //y=7.4 //x2=54.965 //y2=7.4
r1689 (  669 1089 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=54.88 //y=7.23 //x2=54.88 //y2=7.4
r1690 (  669 1179 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.88 //y=7.23 //x2=54.88 //y2=6.745
r1691 (  666 1088 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.085 //y=7.4 //x2=54 //y2=7.4
r1692 (  666 668 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=54.085 //y=7.4 //x2=54.76 //y2=7.4
r1693 (  665 1089 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.795 //y=7.4 //x2=54.88 //y2=7.4
r1694 (  665 668 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=54.795 //y=7.4 //x2=54.76 //y2=7.4
r1695 (  659 1088 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=54 //y=7.23 //x2=54 //y2=7.4
r1696 (  659 1178 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=54 //y=7.23 //x2=54 //y2=6.405
r1697 (  656 1087 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.08 //y=7.4 //x2=52.91 //y2=7.4
r1698 (  656 658 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=53.08 //y=7.4 //x2=53.65 //y2=7.4
r1699 (  655 1088 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.915 //y=7.4 //x2=54 //y2=7.4
r1700 (  655 658 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=53.915 //y=7.4 //x2=53.65 //y2=7.4
r1701 (  650 1086 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.915 //y=7.4 //x2=51.83 //y2=7.4
r1702 (  650 652 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=51.915 //y=7.4 //x2=52.17 //y2=7.4
r1703 (  649 1087 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.74 //y=7.4 //x2=52.91 //y2=7.4
r1704 (  649 652 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=52.74 //y=7.4 //x2=52.17 //y2=7.4
r1705 (  643 1086 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.83 //y=7.23 //x2=51.83 //y2=7.4
r1706 (  643 1177 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=51.83 //y=7.23 //x2=51.83 //y2=6.745
r1707 (  640 1085 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.035 //y=7.4 //x2=50.95 //y2=7.4
r1708 (  640 642 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=51.035 //y=7.4 //x2=51.06 //y2=7.4
r1709 (  639 1086 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.745 //y=7.4 //x2=51.83 //y2=7.4
r1710 (  639 642 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=51.745 //y=7.4 //x2=51.06 //y2=7.4
r1711 (  633 1085 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.95 //y=7.23 //x2=50.95 //y2=7.4
r1712 (  633 1176 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.95 //y=7.23 //x2=50.95 //y2=6.745
r1713 (  632 1084 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.155 //y=7.4 //x2=50.07 //y2=7.4
r1714 (  631 1085 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.865 //y=7.4 //x2=50.95 //y2=7.4
r1715 (  631 632 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.865 //y=7.4 //x2=50.155 //y2=7.4
r1716 (  625 1084 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.07 //y=7.23 //x2=50.07 //y2=7.4
r1717 (  625 1175 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.07 //y=7.23 //x2=50.07 //y2=6.745
r1718 (  622 1083 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.275 //y=7.4 //x2=49.19 //y2=7.4
r1719 (  622 624 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=49.275 //y=7.4 //x2=49.95 //y2=7.4
r1720 (  621 1084 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.985 //y=7.4 //x2=50.07 //y2=7.4
r1721 (  621 624 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=49.985 //y=7.4 //x2=49.95 //y2=7.4
r1722 (  615 1083 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.19 //y=7.23 //x2=49.19 //y2=7.4
r1723 (  615 1174 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=49.19 //y=7.23 //x2=49.19 //y2=6.405
r1724 (  612 1082 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.27 //y=7.4 //x2=48.1 //y2=7.4
r1725 (  612 614 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.27 //y=7.4 //x2=48.84 //y2=7.4
r1726 (  611 1083 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.105 //y=7.4 //x2=49.19 //y2=7.4
r1727 (  611 614 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=49.105 //y=7.4 //x2=48.84 //y2=7.4
r1728 (  606 1081 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.105 //y=7.4 //x2=47.02 //y2=7.4
r1729 (  606 608 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=47.105 //y=7.4 //x2=47.36 //y2=7.4
r1730 (  605 1082 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.93 //y=7.4 //x2=48.1 //y2=7.4
r1731 (  605 608 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=47.93 //y=7.4 //x2=47.36 //y2=7.4
r1732 (  599 1081 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.02 //y=7.23 //x2=47.02 //y2=7.4
r1733 (  599 1173 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=47.02 //y=7.23 //x2=47.02 //y2=6.745
r1734 (  596 1080 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.225 //y=7.4 //x2=46.14 //y2=7.4
r1735 (  596 598 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=46.225 //y=7.4 //x2=46.25 //y2=7.4
r1736 (  595 1081 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.935 //y=7.4 //x2=47.02 //y2=7.4
r1737 (  595 598 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=46.935 //y=7.4 //x2=46.25 //y2=7.4
r1738 (  589 1080 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=46.14 //y=7.23 //x2=46.14 //y2=7.4
r1739 (  589 1172 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.14 //y=7.23 //x2=46.14 //y2=6.745
r1740 (  588 1079 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.345 //y=7.4 //x2=45.26 //y2=7.4
r1741 (  587 1080 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.055 //y=7.4 //x2=46.14 //y2=7.4
r1742 (  587 588 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.055 //y=7.4 //x2=45.345 //y2=7.4
r1743 (  581 1079 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=45.26 //y=7.23 //x2=45.26 //y2=7.4
r1744 (  581 1171 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.26 //y=7.23 //x2=45.26 //y2=6.745
r1745 (  578 1078 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.465 //y=7.4 //x2=44.38 //y2=7.4
r1746 (  578 580 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=44.465 //y=7.4 //x2=45.14 //y2=7.4
r1747 (  577 1079 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.175 //y=7.4 //x2=45.26 //y2=7.4
r1748 (  577 580 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=45.175 //y=7.4 //x2=45.14 //y2=7.4
r1749 (  571 1078 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.38 //y=7.23 //x2=44.38 //y2=7.4
r1750 (  571 1170 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=44.38 //y=7.23 //x2=44.38 //y2=6.405
r1751 (  568 1077 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.46 //y=7.4 //x2=43.29 //y2=7.4
r1752 (  568 570 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.46 //y=7.4 //x2=44.03 //y2=7.4
r1753 (  567 1078 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.295 //y=7.4 //x2=44.38 //y2=7.4
r1754 (  567 570 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=44.295 //y=7.4 //x2=44.03 //y2=7.4
r1755 (  562 1076 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.295 //y=7.4 //x2=42.21 //y2=7.4
r1756 (  562 564 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=42.295 //y=7.4 //x2=42.55 //y2=7.4
r1757 (  561 1077 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.12 //y=7.4 //x2=43.29 //y2=7.4
r1758 (  561 564 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.12 //y=7.4 //x2=42.55 //y2=7.4
r1759 (  555 1076 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=42.21 //y=7.23 //x2=42.21 //y2=7.4
r1760 (  555 1169 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=42.21 //y=7.23 //x2=42.21 //y2=6.745
r1761 (  552 1075 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.415 //y=7.4 //x2=41.33 //y2=7.4
r1762 (  552 554 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=41.415 //y=7.4 //x2=41.44 //y2=7.4
r1763 (  551 1076 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.125 //y=7.4 //x2=42.21 //y2=7.4
r1764 (  551 554 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=42.125 //y=7.4 //x2=41.44 //y2=7.4
r1765 (  545 1075 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=41.33 //y=7.23 //x2=41.33 //y2=7.4
r1766 (  545 1168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=41.33 //y=7.23 //x2=41.33 //y2=6.745
r1767 (  544 1074 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.535 //y=7.4 //x2=40.45 //y2=7.4
r1768 (  543 1075 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.245 //y=7.4 //x2=41.33 //y2=7.4
r1769 (  543 544 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=41.245 //y=7.4 //x2=40.535 //y2=7.4
r1770 (  537 1074 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.45 //y=7.23 //x2=40.45 //y2=7.4
r1771 (  537 1167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=40.45 //y=7.23 //x2=40.45 //y2=6.745
r1772 (  534 1073 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.655 //y=7.4 //x2=39.57 //y2=7.4
r1773 (  534 536 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=39.655 //y=7.4 //x2=40.33 //y2=7.4
r1774 (  533 1074 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.365 //y=7.4 //x2=40.45 //y2=7.4
r1775 (  533 536 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=40.365 //y=7.4 //x2=40.33 //y2=7.4
r1776 (  527 1073 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.57 //y=7.23 //x2=39.57 //y2=7.4
r1777 (  527 1166 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=39.57 //y=7.23 //x2=39.57 //y2=6.405
r1778 (  524 1072 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.65 //y=7.4 //x2=38.48 //y2=7.4
r1779 (  524 526 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.65 //y=7.4 //x2=39.22 //y2=7.4
r1780 (  523 1073 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.485 //y=7.4 //x2=39.57 //y2=7.4
r1781 (  523 526 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=39.485 //y=7.4 //x2=39.22 //y2=7.4
r1782 (  518 1071 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.485 //y=7.4 //x2=37.4 //y2=7.4
r1783 (  518 520 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=37.485 //y=7.4 //x2=37.74 //y2=7.4
r1784 (  517 1072 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.31 //y=7.4 //x2=38.48 //y2=7.4
r1785 (  517 520 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.31 //y=7.4 //x2=37.74 //y2=7.4
r1786 (  511 1071 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.4 //y=7.23 //x2=37.4 //y2=7.4
r1787 (  511 1165 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=37.4 //y=7.23 //x2=37.4 //y2=6.745
r1788 (  508 1070 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.605 //y=7.4 //x2=36.52 //y2=7.4
r1789 (  508 510 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=36.605 //y=7.4 //x2=36.63 //y2=7.4
r1790 (  507 1071 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.315 //y=7.4 //x2=37.4 //y2=7.4
r1791 (  507 510 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=37.315 //y=7.4 //x2=36.63 //y2=7.4
r1792 (  501 1070 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.52 //y=7.23 //x2=36.52 //y2=7.4
r1793 (  501 1164 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=36.52 //y=7.23 //x2=36.52 //y2=6.745
r1794 (  500 1069 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.725 //y=7.4 //x2=35.64 //y2=7.4
r1795 (  499 1070 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.435 //y=7.4 //x2=36.52 //y2=7.4
r1796 (  499 500 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=36.435 //y=7.4 //x2=35.725 //y2=7.4
r1797 (  493 1069 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.64 //y=7.23 //x2=35.64 //y2=7.4
r1798 (  493 1163 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.64 //y=7.23 //x2=35.64 //y2=6.745
r1799 (  490 1068 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.845 //y=7.4 //x2=34.76 //y2=7.4
r1800 (  490 492 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=34.845 //y=7.4 //x2=35.52 //y2=7.4
r1801 (  489 1069 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.555 //y=7.4 //x2=35.64 //y2=7.4
r1802 (  489 492 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=35.555 //y=7.4 //x2=35.52 //y2=7.4
r1803 (  483 1068 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.76 //y=7.23 //x2=34.76 //y2=7.4
r1804 (  483 1162 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=34.76 //y=7.23 //x2=34.76 //y2=6.405
r1805 (  480 1067 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.84 //y=7.4 //x2=33.67 //y2=7.4
r1806 (  480 482 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=33.84 //y=7.4 //x2=34.41 //y2=7.4
r1807 (  479 1068 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.675 //y=7.4 //x2=34.76 //y2=7.4
r1808 (  479 482 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=34.675 //y=7.4 //x2=34.41 //y2=7.4
r1809 (  474 1066 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.675 //y=7.4 //x2=32.59 //y2=7.4
r1810 (  474 476 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=32.675 //y=7.4 //x2=32.93 //y2=7.4
r1811 (  473 1067 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.5 //y=7.4 //x2=33.67 //y2=7.4
r1812 (  473 476 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=33.5 //y=7.4 //x2=32.93 //y2=7.4
r1813 (  467 1066 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.59 //y=7.23 //x2=32.59 //y2=7.4
r1814 (  467 1161 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=32.59 //y=7.23 //x2=32.59 //y2=6.745
r1815 (  464 1065 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.795 //y=7.4 //x2=31.71 //y2=7.4
r1816 (  464 466 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=31.795 //y=7.4 //x2=31.82 //y2=7.4
r1817 (  463 1066 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.505 //y=7.4 //x2=32.59 //y2=7.4
r1818 (  463 466 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=32.505 //y=7.4 //x2=31.82 //y2=7.4
r1819 (  457 1065 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.71 //y=7.23 //x2=31.71 //y2=7.4
r1820 (  457 1160 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.71 //y=7.23 //x2=31.71 //y2=6.745
r1821 (  456 1064 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.915 //y=7.4 //x2=30.83 //y2=7.4
r1822 (  455 1065 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.625 //y=7.4 //x2=31.71 //y2=7.4
r1823 (  455 456 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=31.625 //y=7.4 //x2=30.915 //y2=7.4
r1824 (  449 1064 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.83 //y=7.23 //x2=30.83 //y2=7.4
r1825 (  449 1159 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=30.83 //y=7.23 //x2=30.83 //y2=6.745
r1826 (  446 1063 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.035 //y=7.4 //x2=29.95 //y2=7.4
r1827 (  446 448 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=30.035 //y=7.4 //x2=30.71 //y2=7.4
r1828 (  445 1064 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.745 //y=7.4 //x2=30.83 //y2=7.4
r1829 (  445 448 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=30.745 //y=7.4 //x2=30.71 //y2=7.4
r1830 (  439 1063 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.95 //y=7.23 //x2=29.95 //y2=7.4
r1831 (  439 1158 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=29.95 //y=7.23 //x2=29.95 //y2=6.405
r1832 (  436 1062 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.03 //y=7.4 //x2=28.86 //y2=7.4
r1833 (  436 438 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=29.03 //y=7.4 //x2=29.6 //y2=7.4
r1834 (  435 1063 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.865 //y=7.4 //x2=29.95 //y2=7.4
r1835 (  435 438 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=29.865 //y=7.4 //x2=29.6 //y2=7.4
r1836 (  430 1061 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.865 //y=7.4 //x2=27.78 //y2=7.4
r1837 (  430 432 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=27.865 //y=7.4 //x2=28.12 //y2=7.4
r1838 (  429 1062 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.69 //y=7.4 //x2=28.86 //y2=7.4
r1839 (  429 432 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=28.69 //y=7.4 //x2=28.12 //y2=7.4
r1840 (  423 1061 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.78 //y=7.23 //x2=27.78 //y2=7.4
r1841 (  423 1157 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.78 //y=7.23 //x2=27.78 //y2=6.745
r1842 (  420 1060 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.985 //y=7.4 //x2=26.9 //y2=7.4
r1843 (  420 422 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=26.985 //y=7.4 //x2=27.01 //y2=7.4
r1844 (  419 1061 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.695 //y=7.4 //x2=27.78 //y2=7.4
r1845 (  419 422 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=27.695 //y=7.4 //x2=27.01 //y2=7.4
r1846 (  413 1060 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.9 //y=7.23 //x2=26.9 //y2=7.4
r1847 (  413 1156 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.9 //y=7.23 //x2=26.9 //y2=6.745
r1848 (  412 1059 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.105 //y=7.4 //x2=26.02 //y2=7.4
r1849 (  411 1060 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.815 //y=7.4 //x2=26.9 //y2=7.4
r1850 (  411 412 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.815 //y=7.4 //x2=26.105 //y2=7.4
r1851 (  405 1059 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.02 //y=7.23 //x2=26.02 //y2=7.4
r1852 (  405 1155 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.02 //y=7.23 //x2=26.02 //y2=6.745
r1853 (  402 1058 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.225 //y=7.4 //x2=25.14 //y2=7.4
r1854 (  402 404 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=25.225 //y=7.4 //x2=25.9 //y2=7.4
r1855 (  401 1059 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.935 //y=7.4 //x2=26.02 //y2=7.4
r1856 (  401 404 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=25.935 //y=7.4 //x2=25.9 //y2=7.4
r1857 (  395 1058 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.14 //y=7.23 //x2=25.14 //y2=7.4
r1858 (  395 1154 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=25.14 //y=7.23 //x2=25.14 //y2=6.405
r1859 (  392 1057 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.22 //y=7.4 //x2=24.05 //y2=7.4
r1860 (  392 394 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.22 //y=7.4 //x2=24.79 //y2=7.4
r1861 (  391 1058 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.055 //y=7.4 //x2=25.14 //y2=7.4
r1862 (  391 394 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=25.055 //y=7.4 //x2=24.79 //y2=7.4
r1863 (  386 1056 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.055 //y=7.4 //x2=22.97 //y2=7.4
r1864 (  386 388 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=23.055 //y=7.4 //x2=23.31 //y2=7.4
r1865 (  385 1057 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.88 //y=7.4 //x2=24.05 //y2=7.4
r1866 (  385 388 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.88 //y=7.4 //x2=23.31 //y2=7.4
r1867 (  379 1056 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.97 //y=7.23 //x2=22.97 //y2=7.4
r1868 (  379 1153 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.97 //y=7.23 //x2=22.97 //y2=6.745
r1869 (  376 1055 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.175 //y=7.4 //x2=22.09 //y2=7.4
r1870 (  376 378 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=22.175 //y=7.4 //x2=22.2 //y2=7.4
r1871 (  375 1056 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.885 //y=7.4 //x2=22.97 //y2=7.4
r1872 (  375 378 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=22.885 //y=7.4 //x2=22.2 //y2=7.4
r1873 (  369 1055 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.09 //y=7.23 //x2=22.09 //y2=7.4
r1874 (  369 1152 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.09 //y=7.23 //x2=22.09 //y2=6.745
r1875 (  368 1054 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.295 //y=7.4 //x2=21.21 //y2=7.4
r1876 (  367 1055 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.005 //y=7.4 //x2=22.09 //y2=7.4
r1877 (  367 368 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.005 //y=7.4 //x2=21.295 //y2=7.4
r1878 (  361 1054 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.21 //y=7.23 //x2=21.21 //y2=7.4
r1879 (  361 1151 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.21 //y=7.23 //x2=21.21 //y2=6.745
r1880 (  358 1053 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.415 //y=7.4 //x2=20.33 //y2=7.4
r1881 (  358 360 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=20.415 //y=7.4 //x2=21.09 //y2=7.4
r1882 (  357 1054 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.125 //y=7.4 //x2=21.21 //y2=7.4
r1883 (  357 360 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=21.125 //y=7.4 //x2=21.09 //y2=7.4
r1884 (  351 1053 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.33 //y=7.23 //x2=20.33 //y2=7.4
r1885 (  351 1150 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=20.33 //y=7.23 //x2=20.33 //y2=6.405
r1886 (  348 1052 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.41 //y=7.4 //x2=19.24 //y2=7.4
r1887 (  348 350 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.41 //y=7.4 //x2=19.98 //y2=7.4
r1888 (  347 1053 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.245 //y=7.4 //x2=20.33 //y2=7.4
r1889 (  347 350 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.245 //y=7.4 //x2=19.98 //y2=7.4
r1890 (  342 1051 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.245 //y=7.4 //x2=18.16 //y2=7.4
r1891 (  342 344 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=18.245 //y=7.4 //x2=18.5 //y2=7.4
r1892 (  341 1052 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.07 //y=7.4 //x2=19.24 //y2=7.4
r1893 (  341 344 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.07 //y=7.4 //x2=18.5 //y2=7.4
r1894 (  335 1051 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.16 //y=7.23 //x2=18.16 //y2=7.4
r1895 (  335 1149 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=18.16 //y=7.23 //x2=18.16 //y2=6.745
r1896 (  332 1050 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.365 //y=7.4 //x2=17.28 //y2=7.4
r1897 (  332 334 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=17.365 //y=7.4 //x2=17.39 //y2=7.4
r1898 (  331 1051 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.075 //y=7.4 //x2=18.16 //y2=7.4
r1899 (  331 334 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=18.075 //y=7.4 //x2=17.39 //y2=7.4
r1900 (  325 1050 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.28 //y=7.23 //x2=17.28 //y2=7.4
r1901 (  325 1148 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.28 //y=7.23 //x2=17.28 //y2=6.745
r1902 (  324 1049 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.485 //y=7.4 //x2=16.4 //y2=7.4
r1903 (  323 1050 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.195 //y=7.4 //x2=17.28 //y2=7.4
r1904 (  323 324 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=17.195 //y=7.4 //x2=16.485 //y2=7.4
r1905 (  317 1049 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.4 //y=7.23 //x2=16.4 //y2=7.4
r1906 (  317 1147 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.4 //y=7.23 //x2=16.4 //y2=6.745
r1907 (  314 1048 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.605 //y=7.4 //x2=15.52 //y2=7.4
r1908 (  314 316 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=15.605 //y=7.4 //x2=16.28 //y2=7.4
r1909 (  313 1049 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.315 //y=7.4 //x2=16.4 //y2=7.4
r1910 (  313 316 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=16.315 //y=7.4 //x2=16.28 //y2=7.4
r1911 (  307 1048 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.52 //y=7.23 //x2=15.52 //y2=7.4
r1912 (  307 1146 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=15.52 //y=7.23 //x2=15.52 //y2=6.405
r1913 (  304 1047 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=14.43 //y2=7.4
r1914 (  304 306 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=15.17 //y2=7.4
r1915 (  303 1048 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.435 //y=7.4 //x2=15.52 //y2=7.4
r1916 (  303 306 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.435 //y=7.4 //x2=15.17 //y2=7.4
r1917 (  298 1046 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.435 //y=7.4 //x2=13.35 //y2=7.4
r1918 (  298 300 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=13.435 //y=7.4 //x2=13.69 //y2=7.4
r1919 (  297 1047 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=14.43 //y2=7.4
r1920 (  297 300 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=13.69 //y2=7.4
r1921 (  291 1046 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.35 //y=7.23 //x2=13.35 //y2=7.4
r1922 (  291 1145 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=13.35 //y=7.23 //x2=13.35 //y2=6.745
r1923 (  288 1045 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.555 //y=7.4 //x2=12.47 //y2=7.4
r1924 (  288 290 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=12.555 //y=7.4 //x2=12.58 //y2=7.4
r1925 (  287 1046 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.265 //y=7.4 //x2=13.35 //y2=7.4
r1926 (  287 290 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=13.265 //y=7.4 //x2=12.58 //y2=7.4
r1927 (  281 1045 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.47 //y=7.23 //x2=12.47 //y2=7.4
r1928 (  281 1144 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.47 //y=7.23 //x2=12.47 //y2=6.745
r1929 (  280 1044 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.675 //y=7.4 //x2=11.59 //y2=7.4
r1930 (  279 1045 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.385 //y=7.4 //x2=12.47 //y2=7.4
r1931 (  279 280 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=12.385 //y=7.4 //x2=11.675 //y2=7.4
r1932 (  273 1044 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.59 //y=7.23 //x2=11.59 //y2=7.4
r1933 (  273 1143 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.59 //y=7.23 //x2=11.59 //y2=6.745
r1934 (  270 1043 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.795 //y=7.4 //x2=10.71 //y2=7.4
r1935 (  270 272 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=10.795 //y=7.4 //x2=11.47 //y2=7.4
r1936 (  269 1044 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.505 //y=7.4 //x2=11.59 //y2=7.4
r1937 (  269 272 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=11.505 //y=7.4 //x2=11.47 //y2=7.4
r1938 (  263 1043 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.71 //y=7.23 //x2=10.71 //y2=7.4
r1939 (  263 1142 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.71 //y=7.23 //x2=10.71 //y2=6.405
r1940 (  260 1042 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=9.62 //y2=7.4
r1941 (  260 262 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=10.36 //y2=7.4
r1942 (  259 1043 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.625 //y=7.4 //x2=10.71 //y2=7.4
r1943 (  259 262 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=10.625 //y=7.4 //x2=10.36 //y2=7.4
r1944 (  254 1041 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.54 //y2=7.4
r1945 (  254 256 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.88 //y2=7.4
r1946 (  253 1042 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=9.62 //y2=7.4
r1947 (  253 256 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=8.88 //y2=7.4
r1948 (  247 1041 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=7.4
r1949 (  247 1141 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=6.745
r1950 (  244 1040 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.66 //y2=7.4
r1951 (  244 246 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.77 //y2=7.4
r1952 (  243 1041 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=8.54 //y2=7.4
r1953 (  243 246 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=7.77 //y2=7.4
r1954 (  237 1040 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=7.4
r1955 (  237 1140 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=6.745
r1956 (  236 1039 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=6.78 //y2=7.4
r1957 (  235 1040 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=7.66 //y2=7.4
r1958 (  235 236 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=6.865 //y2=7.4
r1959 (  229 1039 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=7.4
r1960 (  229 1139 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=6.745
r1961 (  226 1038 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=5.9 //y2=7.4
r1962 (  226 228 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=6.66 //y2=7.4
r1963 (  225 1039 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.78 //y2=7.4
r1964 (  225 228 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.66 //y2=7.4
r1965 (  219 1038 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=7.4
r1966 (  219 1138 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=6.405
r1967 (  216 1037 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r1968 (  216 218 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=5.55 //y2=7.4
r1969 (  215 1038 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.9 //y2=7.4
r1970 (  215 218 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.55 //y2=7.4
r1971 (  210 1036 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r1972 (  210 212 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r1973 (  209 1037 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r1974 (  209 212 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r1975 (  203 1036 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r1976 (  203 1137 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r1977 (  200 1035 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r1978 (  200 202 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r1979 (  199 1036 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r1980 (  199 202 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r1981 (  193 1035 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r1982 (  193 1136 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r1983 (  192 1034 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r1984 (  191 1035 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r1985 (  191 192 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r1986 (  185 1034 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r1987 (  185 1135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r1988 (  182 1033 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r1989 (  182 184 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r1990 (  181 1034 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r1991 (  181 184 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r1992 (  175 1033 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r1993 (  175 1134 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r1994 (  171 1033 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r1995 (  171 174 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r1996 (  167 1133 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=98.05 //y=7.4 //x2=98.05 //y2=7.4
r1997 (  165 1131 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=97.31 //y=7.4 //x2=97.31 //y2=7.4
r1998 (  165 167 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=97.31 //y=7.4 //x2=98.05 //y2=7.4
r1999 (  163 1010 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=95.83 //y=7.4 //x2=95.83 //y2=7.4
r2000 (  163 165 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=95.83 //y=7.4 //x2=97.31 //y2=7.4
r2001 (  161 1008 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=94.72 //y=7.4 //x2=94.72 //y2=7.4
r2002 (  161 163 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=94.72 //y=7.4 //x2=95.83 //y2=7.4
r2003 (  159 1006 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=93.61 //y=7.4 //x2=93.61 //y2=7.4
r2004 (  159 161 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=93.61 //y=7.4 //x2=94.72 //y2=7.4
r2005 (  157 1000 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=92.13 //y=7.4 //x2=92.13 //y2=7.4
r2006 (  157 159 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=92.13 //y=7.4 //x2=93.61 //y2=7.4
r2007 (  155 998 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=91.02 //y=7.4 //x2=91.02 //y2=7.4
r2008 (  155 157 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=91.02 //y=7.4 //x2=92.13 //y2=7.4
r2009 (  153 992 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=89.54 //y=7.4 //x2=89.54 //y2=7.4
r2010 (  153 155 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=89.54 //y=7.4 //x2=91.02 //y2=7.4
r2011 (  151 982 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=88.43 //y=7.4 //x2=88.43 //y2=7.4
r2012 (  151 153 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=88.43 //y=7.4 //x2=89.54 //y2=7.4
r2013 (  149 1124 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=87.32 //y=7.4 //x2=87.32 //y2=7.4
r2014 (  149 151 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=87.32 //y=7.4 //x2=88.43 //y2=7.4
r2015 (  147 960 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=85.84 //y=7.4 //x2=85.84 //y2=7.4
r2016 (  147 149 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=85.84 //y=7.4 //x2=87.32 //y2=7.4
r2017 (  145 950 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=84.73 //y=7.4 //x2=84.73 //y2=7.4
r2018 (  145 147 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=84.73 //y=7.4 //x2=85.84 //y2=7.4
r2019 (  143 932 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=83.62 //y=7.4 //x2=83.62 //y2=7.4
r2020 (  143 145 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=83.62 //y=7.4 //x2=84.73 //y2=7.4
r2021 (  141 922 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.51 //y=7.4 //x2=82.51 //y2=7.4
r2022 (  141 143 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=82.51 //y=7.4 //x2=83.62 //y2=7.4
r2023 (  139 916 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=81.03 //y=7.4 //x2=81.03 //y2=7.4
r2024 (  139 141 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=81.03 //y=7.4 //x2=82.51 //y2=7.4
r2025 (  137 906 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=79.92 //y=7.4 //x2=79.92 //y2=7.4
r2026 (  137 139 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=79.92 //y=7.4 //x2=81.03 //y2=7.4
r2027 (  135 888 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.81 //y=7.4 //x2=78.81 //y2=7.4
r2028 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=78.81 //y=7.4 //x2=79.92 //y2=7.4
r2029 (  133 878 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=77.7 //y=7.4 //x2=77.7 //y2=7.4
r2030 (  133 135 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=77.7 //y=7.4 //x2=78.81 //y2=7.4
r2031 (  131 872 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.22 //y=7.4 //x2=76.22 //y2=7.4
r2032 (  131 133 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.22 //y=7.4 //x2=77.7 //y2=7.4
r2033 (  129 862 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.11 //y=7.4 //x2=75.11 //y2=7.4
r2034 (  129 131 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=7.4 //x2=76.22 //y2=7.4
r2035 (  127 844 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74 //y=7.4 //x2=74 //y2=7.4
r2036 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74 //y=7.4 //x2=75.11 //y2=7.4
r2037 (  125 834 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.89 //y=7.4 //x2=72.89 //y2=7.4
r2038 (  125 127 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=72.89 //y=7.4 //x2=74 //y2=7.4
r2039 (  123 828 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=7.4 //x2=71.41 //y2=7.4
r2040 (  123 125 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=7.4 //x2=72.89 //y2=7.4
r2041 (  121 818 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=70.3 //y=7.4 //x2=70.3 //y2=7.4
r2042 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=70.3 //y=7.4 //x2=71.41 //y2=7.4
r2043 (  119 800 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.19 //y=7.4 //x2=69.19 //y2=7.4
r2044 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.19 //y=7.4 //x2=70.3 //y2=7.4
r2045 (  117 790 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=68.08 //y=7.4 //x2=68.08 //y2=7.4
r2046 (  117 119 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=68.08 //y=7.4 //x2=69.19 //y2=7.4
r2047 (  115 784 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.6 //y=7.4 //x2=66.6 //y2=7.4
r2048 (  115 117 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=66.6 //y=7.4 //x2=68.08 //y2=7.4
r2049 (  113 774 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.49 //y=7.4 //x2=65.49 //y2=7.4
r2050 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.49 //y=7.4 //x2=66.6 //y2=7.4
r2051 (  111 756 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=64.38 //y=7.4 //x2=64.38 //y2=7.4
r2052 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=64.38 //y=7.4 //x2=65.49 //y2=7.4
r2053 (  109 746 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=63.27 //y=7.4 //x2=63.27 //y2=7.4
r2054 (  109 111 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=63.27 //y=7.4 //x2=64.38 //y2=7.4
r2055 (  107 740 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.79 //y=7.4 //x2=61.79 //y2=7.4
r2056 (  107 109 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.79 //y=7.4 //x2=63.27 //y2=7.4
r2057 (  105 730 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=60.68 //y=7.4 //x2=60.68 //y2=7.4
r2058 (  105 107 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=60.68 //y=7.4 //x2=61.79 //y2=7.4
r2059 (  103 712 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.57 //y=7.4 //x2=59.57 //y2=7.4
r2060 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.57 //y=7.4 //x2=60.68 //y2=7.4
r2061 (  101 702 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.46 //y=7.4 //x2=58.46 //y2=7.4
r2062 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.46 //y=7.4 //x2=59.57 //y2=7.4
r2063 (  99 696 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.98 //y=7.4 //x2=56.98 //y2=7.4
r2064 (  99 101 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.98 //y=7.4 //x2=58.46 //y2=7.4
r2065 (  97 686 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.87 //y=7.4 //x2=55.87 //y2=7.4
r2066 (  97 99 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.87 //y=7.4 //x2=56.98 //y2=7.4
r2067 (  95 668 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.76 //y=7.4 //x2=54.76 //y2=7.4
r2068 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.76 //y=7.4 //x2=55.87 //y2=7.4
r2069 (  93 658 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.65 //y=7.4 //x2=53.65 //y2=7.4
r2070 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=53.65 //y=7.4 //x2=54.76 //y2=7.4
r2071 (  91 652 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=52.17 //y=7.4 //x2=52.17 //y2=7.4
r2072 (  91 93 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=52.17 //y=7.4 //x2=53.65 //y2=7.4
r2073 (  89 642 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.06 //y=7.4 //x2=51.06 //y2=7.4
r2074 (  89 91 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=51.06 //y=7.4 //x2=52.17 //y2=7.4
r2075 (  87 624 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.95 //y=7.4 //x2=49.95 //y2=7.4
r2076 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.95 //y=7.4 //x2=51.06 //y2=7.4
r2077 (  84 614 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.84 //y=7.4 //x2=48.84 //y2=7.4
r2078 (  82 608 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=47.36 //y=7.4 //x2=47.36 //y2=7.4
r2079 (  82 84 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=47.36 //y=7.4 //x2=48.84 //y2=7.4
r2080 (  80 598 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.25 //y=7.4 //x2=46.25 //y2=7.4
r2081 (  80 82 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.25 //y=7.4 //x2=47.36 //y2=7.4
r2082 (  78 580 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.14 //y=7.4 //x2=45.14 //y2=7.4
r2083 (  78 80 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.14 //y=7.4 //x2=46.25 //y2=7.4
r2084 (  76 570 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.03 //y=7.4 //x2=44.03 //y2=7.4
r2085 (  76 78 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.03 //y=7.4 //x2=45.14 //y2=7.4
r2086 (  74 564 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.55 //y=7.4 //x2=42.55 //y2=7.4
r2087 (  74 76 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=42.55 //y=7.4 //x2=44.03 //y2=7.4
r2088 (  72 554 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.44 //y=7.4 //x2=41.44 //y2=7.4
r2089 (  72 74 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.44 //y=7.4 //x2=42.55 //y2=7.4
r2090 (  70 536 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=40.33 //y=7.4 //x2=40.33 //y2=7.4
r2091 (  70 72 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=40.33 //y=7.4 //x2=41.44 //y2=7.4
r2092 (  68 526 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.22 //y=7.4 //x2=39.22 //y2=7.4
r2093 (  68 70 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=39.22 //y=7.4 //x2=40.33 //y2=7.4
r2094 (  66 520 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37.74 //y=7.4 //x2=37.74 //y2=7.4
r2095 (  66 68 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=37.74 //y=7.4 //x2=39.22 //y2=7.4
r2096 (  64 510 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=36.63 //y=7.4 //x2=36.63 //y2=7.4
r2097 (  64 66 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=36.63 //y=7.4 //x2=37.74 //y2=7.4
r2098 (  62 492 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.52 //y=7.4 //x2=35.52 //y2=7.4
r2099 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.52 //y=7.4 //x2=36.63 //y2=7.4
r2100 (  60 482 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.41 //y=7.4 //x2=34.41 //y2=7.4
r2101 (  60 62 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.41 //y=7.4 //x2=35.52 //y2=7.4
r2102 (  58 476 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.93 //y=7.4 //x2=32.93 //y2=7.4
r2103 (  58 60 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.93 //y=7.4 //x2=34.41 //y2=7.4
r2104 (  56 466 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.82 //y=7.4 //x2=31.82 //y2=7.4
r2105 (  56 58 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.82 //y=7.4 //x2=32.93 //y2=7.4
r2106 (  54 448 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=30.71 //y=7.4 //x2=30.71 //y2=7.4
r2107 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=30.71 //y=7.4 //x2=31.82 //y2=7.4
r2108 (  52 438 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.6 //y=7.4 //x2=29.6 //y2=7.4
r2109 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=29.6 //y=7.4 //x2=30.71 //y2=7.4
r2110 (  50 432 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.12 //y=7.4 //x2=28.12 //y2=7.4
r2111 (  50 52 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=28.12 //y=7.4 //x2=29.6 //y2=7.4
r2112 (  48 422 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.01 //y=7.4 //x2=27.01 //y2=7.4
r2113 (  48 50 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.01 //y=7.4 //x2=28.12 //y2=7.4
r2114 (  46 404 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.9 //y=7.4 //x2=25.9 //y2=7.4
r2115 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.9 //y=7.4 //x2=27.01 //y2=7.4
r2116 (  44 394 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=7.4 //x2=24.79 //y2=7.4
r2117 (  44 46 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=7.4 //x2=25.9 //y2=7.4
r2118 (  42 388 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.31 //y=7.4 //x2=23.31 //y2=7.4
r2119 (  42 44 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.31 //y=7.4 //x2=24.79 //y2=7.4
r2120 (  40 378 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=7.4 //x2=22.2 //y2=7.4
r2121 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=7.4 //x2=23.31 //y2=7.4
r2122 (  38 360 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=7.4 //x2=21.09 //y2=7.4
r2123 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=7.4 //x2=22.2 //y2=7.4
r2124 (  36 350 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=7.4 //x2=19.98 //y2=7.4
r2125 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=7.4 //x2=21.09 //y2=7.4
r2126 (  34 344 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=7.4 //x2=18.5 //y2=7.4
r2127 (  34 36 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=7.4 //x2=19.98 //y2=7.4
r2128 (  32 334 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r2129 (  32 34 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.4 //x2=18.5 //y2=7.4
r2130 (  30 316 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=7.4 //x2=16.28 //y2=7.4
r2131 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=7.4 //x2=17.39 //y2=7.4
r2132 (  28 306 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r2133 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.28 //y2=7.4
r2134 (  26 300 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=7.4 //x2=13.69 //y2=7.4
r2135 (  26 28 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=7.4 //x2=15.17 //y2=7.4
r2136 (  24 290 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r2137 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.4 //x2=13.69 //y2=7.4
r2138 (  22 272 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r2139 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=7.4 //x2=12.58 //y2=7.4
r2140 (  20 262 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r2141 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r2142 (  18 256 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=7.4 //x2=8.88 //y2=7.4
r2143 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=7.4 //x2=10.36 //y2=7.4
r2144 (  16 246 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r2145 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=8.88 //y2=7.4
r2146 (  14 228 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r2147 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r2148 (  12 218 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r2149 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r2150 (  10 212 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r2151 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.4 //x2=5.55 //y2=7.4
r2152 (  8 202 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r2153 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r2154 (  6 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r2155 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r2156 (  3 174 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r2157 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r2158 (  1 87 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=49.395 //y=7.4 //x2=49.95 //y2=7.4
r2159 (  1 84 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=49.395 //y=7.4 //x2=48.84 //y2=7.4
ends PM_TMRDFFSNRNQX1\%VDD

subckt PM_TMRDFFSNRNQX1\%noxref_3 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 \
 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c240 ( 127 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c241 ( 126 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c242 ( 125 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c243 ( 123 0 ) capacitor c=0.00853354f //x=3.395 //y=0.915
c244 ( 103 0 ) capacitor c=0.0556143f //x=11.005 //y=4.79
c245 ( 102 0 ) capacitor c=0.0293157f //x=11.295 //y=4.79
c246 ( 101 0 ) capacitor c=0.0347816f //x=10.96 //y=1.22
c247 ( 100 0 ) capacitor c=0.0187487f //x=10.96 //y=0.875
c248 ( 94 0 ) capacitor c=0.0137055f //x=10.805 //y=1.375
c249 ( 92 0 ) capacitor c=0.0149861f //x=10.805 //y=0.72
c250 ( 91 0 ) capacitor c=0.096037f //x=10.43 //y=1.915
c251 ( 90 0 ) capacitor c=0.0228993f //x=10.43 //y=1.53
c252 ( 89 0 ) capacitor c=0.0234352f //x=10.43 //y=1.22
c253 ( 88 0 ) capacitor c=0.0198724f //x=10.43 //y=0.875
c254 ( 84 0 ) capacitor c=0.055995f //x=6.195 //y=4.79
c255 ( 83 0 ) capacitor c=0.0298189f //x=6.485 //y=4.79
c256 ( 82 0 ) capacitor c=0.0347816f //x=6.15 //y=1.22
c257 ( 81 0 ) capacitor c=0.0187487f //x=6.15 //y=0.875
c258 ( 75 0 ) capacitor c=0.0137055f //x=5.995 //y=1.375
c259 ( 73 0 ) capacitor c=0.0149861f //x=5.995 //y=0.72
c260 ( 72 0 ) capacitor c=0.096037f //x=5.62 //y=1.915
c261 ( 71 0 ) capacitor c=0.0228993f //x=5.62 //y=1.53
c262 ( 70 0 ) capacitor c=0.0234352f //x=5.62 //y=1.22
c263 ( 69 0 ) capacitor c=0.0198724f //x=5.62 //y=0.875
c264 ( 68 0 ) capacitor c=0.110114f //x=11.37 //y=6.02
c265 ( 67 0 ) capacitor c=0.158956f //x=10.93 //y=6.02
c266 ( 66 0 ) capacitor c=0.110114f //x=6.56 //y=6.02
c267 ( 65 0 ) capacitor c=0.158956f //x=6.12 //y=6.02
c268 ( 62 0 ) capacitor c=0.00116729f //x=3.29 //y=5.155
c269 ( 61 0 ) capacitor c=0.00226015f //x=2.41 //y=5.155
c270 ( 54 0 ) capacitor c=0.0970684f //x=10.73 //y=2.08
c271 ( 46 0 ) capacitor c=0.102314f //x=5.92 //y=2.08
c272 ( 44 0 ) capacitor c=0.111586f //x=4.07 //y=2.59
c273 ( 40 0 ) capacitor c=0.00398962f //x=3.67 //y=1.665
c274 ( 39 0 ) capacitor c=0.0137288f //x=3.985 //y=1.665
c275 ( 33 0 ) capacitor c=0.0291119f //x=3.985 //y=5.155
c276 ( 25 0 ) capacitor c=0.0184197f //x=3.205 //y=5.155
c277 ( 18 0 ) capacitor c=0.00351598f //x=1.615 //y=5.155
c278 ( 17 0 ) capacitor c=0.0155255f //x=2.325 //y=5.155
c279 ( 4 0 ) capacitor c=0.00440131f //x=6.035 //y=2.59
c280 ( 3 0 ) capacitor c=0.0870935f //x=10.615 //y=2.59
c281 ( 2 0 ) capacitor c=0.0124623f //x=4.185 //y=2.59
c282 ( 1 0 ) capacitor c=0.0300768f //x=5.805 //y=2.59
r283 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.295 //y=4.79 //x2=11.37 //y2=4.865
r284 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=11.295 //y=4.79 //x2=11.005 //y2=4.79
r285 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.96 //y=1.22 //x2=10.92 //y2=1.375
r286 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.96 //y=0.875 //x2=10.92 //y2=0.72
r287 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.96 //y=0.875 //x2=10.96 //y2=1.22
r288 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.93 //y=4.865 //x2=11.005 //y2=4.79
r289 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=10.93 //y=4.865 //x2=10.73 //y2=4.7
r290 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.585 //y=1.375 //x2=10.47 //y2=1.375
r291 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.805 //y=1.375 //x2=10.92 //y2=1.375
r292 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.585 //y=0.72 //x2=10.47 //y2=0.72
r293 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.805 //y=0.72 //x2=10.92 //y2=0.72
r294 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.805 //y=0.72 //x2=10.585 //y2=0.72
r295 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.915 //x2=10.73 //y2=2.08
r296 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.53 //x2=10.47 //y2=1.375
r297 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.53 //x2=10.43 //y2=1.915
r298 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.22 //x2=10.47 //y2=1.375
r299 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=0.875 //x2=10.47 //y2=0.72
r300 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.43 //y=0.875 //x2=10.43 //y2=1.22
r301 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.56 //y2=4.865
r302 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.195 //y2=4.79
r303 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=1.22 //x2=6.11 //y2=1.375
r304 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.11 //y2=0.72
r305 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.15 //y2=1.22
r306 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=6.195 //y2=4.79
r307 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=5.92 //y2=4.7
r308 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=1.375 //x2=5.66 //y2=1.375
r309 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=1.375 //x2=6.11 //y2=1.375
r310 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=0.72 //x2=5.66 //y2=0.72
r311 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=6.11 //y2=0.72
r312 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=5.775 //y2=0.72
r313 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.915 //x2=5.92 //y2=2.08
r314 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.66 //y2=1.375
r315 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.62 //y2=1.915
r316 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.22 //x2=5.66 //y2=1.375
r317 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.66 //y2=0.72
r318 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.62 //y2=1.22
r319 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.37 //y=6.02 //x2=11.37 //y2=4.865
r320 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.93 //y=6.02 //x2=10.93 //y2=4.865
r321 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.56 //y=6.02 //x2=6.56 //y2=4.865
r322 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.12 //y=6.02 //x2=6.12 //y2=4.865
r323 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.695 //y=1.375 //x2=10.805 //y2=1.375
r324 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.695 //y=1.375 //x2=10.585 //y2=1.375
r325 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.995 //y2=1.375
r326 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.775 //y2=1.375
r327 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=4.7 //x2=10.73 //y2=4.7
r328 (  57 59 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.59 //x2=10.73 //y2=4.7
r329 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=2.08 //x2=10.73 //y2=2.08
r330 (  54 57 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.08 //x2=10.73 //y2=2.59
r331 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.7 //x2=5.92 //y2=4.7
r332 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.59 //x2=5.92 //y2=4.7
r333 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r334 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=2.59
r335 (  42 44 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=2.59
r336 (  41 44 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=2.59
r337 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r338 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r339 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r340 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r341 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r342 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r343 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r344 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r345 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r346 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r347 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r348 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r349 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r350 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r351 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r352 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r353 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r354 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r355 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=2.59 //x2=10.73 //y2=2.59
r356 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=2.59 //x2=5.92 //y2=2.59
r357 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=2.59 //x2=4.07 //y2=2.59
r358 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=2.59 //x2=5.92 //y2=2.59
r359 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.59 //x2=10.73 //y2=2.59
r360 (  3 4 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.59 //x2=6.035 //y2=2.59
r361 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=2.59 //x2=4.07 //y2=2.59
r362 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.805 //y=2.59 //x2=5.92 //y2=2.59
r363 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.805 //y=2.59 //x2=4.185 //y2=2.59
ends PM_TMRDFFSNRNQX1\%noxref_3

subckt PM_TMRDFFSNRNQX1\%noxref_4 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c165 ( 85 0 ) capacitor c=0.023087f //x=12.765 //y=5.02
c166 ( 84 0 ) capacitor c=0.023519f //x=11.885 //y=5.02
c167 ( 83 0 ) capacitor c=0.0224735f //x=11.005 //y=5.02
c168 ( 81 0 ) capacitor c=0.00853354f //x=13.015 //y=0.915
c169 ( 69 0 ) capacitor c=0.0557698f //x=15.815 //y=4.79
c170 ( 68 0 ) capacitor c=0.0293157f //x=16.105 //y=4.79
c171 ( 67 0 ) capacitor c=0.0347816f //x=15.77 //y=1.22
c172 ( 66 0 ) capacitor c=0.0187487f //x=15.77 //y=0.875
c173 ( 60 0 ) capacitor c=0.0137055f //x=15.615 //y=1.375
c174 ( 58 0 ) capacitor c=0.0149861f //x=15.615 //y=0.72
c175 ( 57 0 ) capacitor c=0.096037f //x=15.24 //y=1.915
c176 ( 56 0 ) capacitor c=0.0228993f //x=15.24 //y=1.53
c177 ( 55 0 ) capacitor c=0.0234352f //x=15.24 //y=1.22
c178 ( 54 0 ) capacitor c=0.0198724f //x=15.24 //y=0.875
c179 ( 53 0 ) capacitor c=0.110114f //x=16.18 //y=6.02
c180 ( 52 0 ) capacitor c=0.158956f //x=15.74 //y=6.02
c181 ( 50 0 ) capacitor c=0.00106608f //x=12.91 //y=5.155
c182 ( 49 0 ) capacitor c=0.00207319f //x=12.03 //y=5.155
c183 ( 42 0 ) capacitor c=0.0939064f //x=15.54 //y=2.08
c184 ( 40 0 ) capacitor c=0.10406f //x=13.69 //y=2.59
c185 ( 36 0 ) capacitor c=0.00398962f //x=13.29 //y=1.665
c186 ( 35 0 ) capacitor c=0.0137288f //x=13.605 //y=1.665
c187 ( 29 0 ) capacitor c=0.0283082f //x=13.605 //y=5.155
c188 ( 21 0 ) capacitor c=0.0176454f //x=12.825 //y=5.155
c189 ( 14 0 ) capacitor c=0.00332903f //x=11.235 //y=5.155
c190 ( 13 0 ) capacitor c=0.0148427f //x=11.945 //y=5.155
c191 ( 2 0 ) capacitor c=0.00808366f //x=13.805 //y=2.59
c192 ( 1 0 ) capacitor c=0.0352679f //x=15.425 //y=2.59
r193 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=16.105 //y=4.79 //x2=16.18 //y2=4.865
r194 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=16.105 //y=4.79 //x2=15.815 //y2=4.79
r195 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.77 //y=1.22 //x2=15.73 //y2=1.375
r196 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.77 //y=0.875 //x2=15.73 //y2=0.72
r197 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.77 //y=0.875 //x2=15.77 //y2=1.22
r198 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.74 //y=4.865 //x2=15.815 //y2=4.79
r199 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=15.74 //y=4.865 //x2=15.54 //y2=4.7
r200 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.395 //y=1.375 //x2=15.28 //y2=1.375
r201 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.615 //y=1.375 //x2=15.73 //y2=1.375
r202 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.395 //y=0.72 //x2=15.28 //y2=0.72
r203 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.615 //y=0.72 //x2=15.73 //y2=0.72
r204 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.615 //y=0.72 //x2=15.395 //y2=0.72
r205 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.915 //x2=15.54 //y2=2.08
r206 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.53 //x2=15.28 //y2=1.375
r207 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.53 //x2=15.24 //y2=1.915
r208 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.22 //x2=15.28 //y2=1.375
r209 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=0.875 //x2=15.28 //y2=0.72
r210 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.24 //y=0.875 //x2=15.24 //y2=1.22
r211 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.18 //y=6.02 //x2=16.18 //y2=4.865
r212 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.74 //y=6.02 //x2=15.74 //y2=4.865
r213 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.505 //y=1.375 //x2=15.615 //y2=1.375
r214 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.505 //y=1.375 //x2=15.395 //y2=1.375
r215 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=4.7 //x2=15.54 //y2=4.7
r216 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=15.54 //y=2.59 //x2=15.54 //y2=4.7
r217 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=2.08 //x2=15.54 //y2=2.08
r218 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=15.54 //y=2.08 //x2=15.54 //y2=2.59
r219 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=13.69 //y=5.07 //x2=13.69 //y2=2.59
r220 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=13.69 //y=1.75 //x2=13.69 //y2=2.59
r221 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.665 //x2=13.69 //y2=1.75
r222 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.665 //x2=13.29 //y2=1.665
r223 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.205 //y=1.58 //x2=13.29 //y2=1.665
r224 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=13.205 //y=1.58 //x2=13.205 //y2=1.01
r225 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.995 //y=5.155 //x2=12.91 //y2=5.155
r226 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.155 //x2=13.69 //y2=5.07
r227 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.155 //x2=12.995 //y2=5.155
r228 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.91 //y=5.24 //x2=12.91 //y2=5.155
r229 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.91 //y=5.24 //x2=12.91 //y2=5.725
r230 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.115 //y=5.155 //x2=12.03 //y2=5.155
r231 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.825 //y=5.155 //x2=12.91 //y2=5.155
r232 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=12.825 //y=5.155 //x2=12.115 //y2=5.155
r233 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.03 //y=5.24 //x2=12.03 //y2=5.155
r234 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.03 //y=5.24 //x2=12.03 //y2=5.725
r235 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.945 //y=5.155 //x2=12.03 //y2=5.155
r236 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.945 //y=5.155 //x2=11.235 //y2=5.155
r237 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.15 //y=5.24 //x2=11.235 //y2=5.155
r238 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.15 //y=5.24 //x2=11.15 //y2=5.725
r239 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=2.59 //x2=15.54 //y2=2.59
r240 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=13.69 //y=2.59 //x2=13.69 //y2=2.59
r241 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.805 //y=2.59 //x2=13.69 //y2=2.59
r242 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=2.59 //x2=15.54 //y2=2.59
r243 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=15.425 //y=2.59 //x2=13.805 //y2=2.59
ends PM_TMRDFFSNRNQX1\%noxref_4

subckt PM_TMRDFFSNRNQX1\%noxref_5 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 \
 63 64 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 90 92 98 99 100 101 106 \
 107 112 123 125 126 127 )
c267 ( 127 0 ) capacitor c=0.023087f //x=7.955 //y=5.02
c268 ( 126 0 ) capacitor c=0.023519f //x=7.075 //y=5.02
c269 ( 125 0 ) capacitor c=0.0224735f //x=6.195 //y=5.02
c270 ( 123 0 ) capacitor c=0.00853354f //x=8.205 //y=0.915
c271 ( 112 0 ) capacitor c=0.059212f //x=3.33 //y=4.7
c272 ( 107 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c273 ( 106 0 ) capacitor c=0.045877f //x=3.33 //y=2.08
c274 ( 101 0 ) capacitor c=0.0556143f //x=20.625 //y=4.79
c275 ( 100 0 ) capacitor c=0.0293157f //x=20.915 //y=4.79
c276 ( 99 0 ) capacitor c=0.0347816f //x=20.58 //y=1.22
c277 ( 98 0 ) capacitor c=0.0187487f //x=20.58 //y=0.875
c278 ( 92 0 ) capacitor c=0.0137055f //x=20.425 //y=1.375
c279 ( 90 0 ) capacitor c=0.0149861f //x=20.425 //y=0.72
c280 ( 89 0 ) capacitor c=0.096037f //x=20.05 //y=1.915
c281 ( 88 0 ) capacitor c=0.0228993f //x=20.05 //y=1.53
c282 ( 87 0 ) capacitor c=0.0234352f //x=20.05 //y=1.22
c283 ( 86 0 ) capacitor c=0.0198724f //x=20.05 //y=0.875
c284 ( 85 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c285 ( 84 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c286 ( 81 0 ) capacitor c=0.0148873f //x=3.695 //y=1.415
c287 ( 79 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c288 ( 74 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c289 ( 73 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c290 ( 72 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c291 ( 68 0 ) capacitor c=0.110114f //x=20.99 //y=6.02
c292 ( 67 0 ) capacitor c=0.158956f //x=20.55 //y=6.02
c293 ( 66 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c294 ( 65 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c295 ( 62 0 ) capacitor c=0.00106608f //x=8.1 //y=5.155
c296 ( 61 0 ) capacitor c=0.00207162f //x=7.22 //y=5.155
c297 ( 54 0 ) capacitor c=0.0965808f //x=20.35 //y=2.08
c298 ( 52 0 ) capacitor c=0.10653f //x=8.88 //y=3.33
c299 ( 48 0 ) capacitor c=0.00398962f //x=8.48 //y=1.665
c300 ( 47 0 ) capacitor c=0.0137288f //x=8.795 //y=1.665
c301 ( 41 0 ) capacitor c=0.0283082f //x=8.795 //y=5.155
c302 ( 33 0 ) capacitor c=0.0176454f //x=8.015 //y=5.155
c303 ( 26 0 ) capacitor c=0.00351598f //x=6.425 //y=5.155
c304 ( 25 0 ) capacitor c=0.0154196f //x=7.135 //y=5.155
c305 ( 12 0 ) capacitor c=0.0883624f //x=3.33 //y=2.08
c306 ( 4 0 ) capacitor c=0.00578611f //x=8.995 //y=3.33
c307 ( 3 0 ) capacitor c=0.184375f //x=20.235 //y=3.33
c308 ( 2 0 ) capacitor c=0.0148738f //x=3.445 //y=3.33
c309 ( 1 0 ) capacitor c=0.107193f //x=8.765 //y=3.33
r310 (  106 107 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r311 (  100 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.915 //y=4.79 //x2=20.99 //y2=4.865
r312 (  100 101 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=20.915 //y=4.79 //x2=20.625 //y2=4.79
r313 (  99 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.58 //y=1.22 //x2=20.54 //y2=1.375
r314 (  98 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.58 //y=0.875 //x2=20.54 //y2=0.72
r315 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.58 //y=0.875 //x2=20.58 //y2=1.22
r316 (  95 101 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.55 //y=4.865 //x2=20.625 //y2=4.79
r317 (  95 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=20.55 //y=4.865 //x2=20.35 //y2=4.7
r318 (  93 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.205 //y=1.375 //x2=20.09 //y2=1.375
r319 (  92 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.425 //y=1.375 //x2=20.54 //y2=1.375
r320 (  91 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.205 //y=0.72 //x2=20.09 //y2=0.72
r321 (  90 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.425 //y=0.72 //x2=20.54 //y2=0.72
r322 (  90 91 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.425 //y=0.72 //x2=20.205 //y2=0.72
r323 (  89 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.915 //x2=20.35 //y2=2.08
r324 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.53 //x2=20.09 //y2=1.375
r325 (  88 89 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.53 //x2=20.05 //y2=1.915
r326 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.22 //x2=20.09 //y2=1.375
r327 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=0.875 //x2=20.09 //y2=0.72
r328 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.05 //y=0.875 //x2=20.05 //y2=1.22
r329 (  85 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r330 (  84 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r331 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r332 (  82 110 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r333 (  81 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r334 (  80 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r335 (  79 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r336 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r337 (  76 112 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r338 (  74 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r339 (  74 107 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r340 (  73 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r341 (  72 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r342 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r343 (  69 112 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r344 (  68 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.99 //y=6.02 //x2=20.99 //y2=4.865
r345 (  67 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.55 //y=6.02 //x2=20.55 //y2=4.865
r346 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r347 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r348 (  64 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.315 //y=1.375 //x2=20.425 //y2=1.375
r349 (  64 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.315 //y=1.375 //x2=20.205 //y2=1.375
r350 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r351 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r352 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.35 //y=4.7 //x2=20.35 //y2=4.7
r353 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=20.35 //y=3.33 //x2=20.35 //y2=4.7
r354 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.35 //y=2.08 //x2=20.35 //y2=2.08
r355 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=20.35 //y=2.08 //x2=20.35 //y2=3.33
r356 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=8.88 //y=5.07 //x2=8.88 //y2=3.33
r357 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=8.88 //y=1.75 //x2=8.88 //y2=3.33
r358 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.88 //y2=1.75
r359 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.48 //y2=1.665
r360 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.48 //y2=1.665
r361 (  43 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.395 //y2=1.01
r362 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.185 //y=5.155 //x2=8.1 //y2=5.155
r363 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.88 //y2=5.07
r364 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.185 //y2=5.155
r365 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.155
r366 (  35 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.725
r367 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.305 //y=5.155 //x2=7.22 //y2=5.155
r368 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=8.1 //y2=5.155
r369 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=7.305 //y2=5.155
r370 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.155
r371 (  27 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.725
r372 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=7.22 //y2=5.155
r373 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=6.425 //y2=5.155
r374 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.425 //y2=5.155
r375 (  19 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.34 //y2=5.725
r376 (  17 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r377 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.33 //x2=3.33 //y2=4.7
r378 (  12 106 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r379 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.33
r380 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.35 //y=3.33 //x2=20.35 //y2=3.33
r381 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.88 //y=3.33 //x2=8.88 //y2=3.33
r382 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.33 //x2=3.33 //y2=3.33
r383 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.995 //y=3.33 //x2=8.88 //y2=3.33
r384 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.235 //y=3.33 //x2=20.35 //y2=3.33
r385 (  3 4 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=20.235 //y=3.33 //x2=8.995 //y2=3.33
r386 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.445 //y=3.33 //x2=3.33 //y2=3.33
r387 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=8.88 //y2=3.33
r388 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=3.445 //y2=3.33
ends PM_TMRDFFSNRNQX1\%noxref_5

subckt PM_TMRDFFSNRNQX1\%noxref_6 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c164 ( 85 0 ) capacitor c=0.023087f //x=22.385 //y=5.02
c165 ( 84 0 ) capacitor c=0.023519f //x=21.505 //y=5.02
c166 ( 83 0 ) capacitor c=0.0224735f //x=20.625 //y=5.02
c167 ( 81 0 ) capacitor c=0.00853354f //x=22.635 //y=0.915
c168 ( 69 0 ) capacitor c=0.0556143f //x=25.435 //y=4.79
c169 ( 68 0 ) capacitor c=0.0293157f //x=25.725 //y=4.79
c170 ( 67 0 ) capacitor c=0.0347816f //x=25.39 //y=1.22
c171 ( 66 0 ) capacitor c=0.0187487f //x=25.39 //y=0.875
c172 ( 60 0 ) capacitor c=0.0137055f //x=25.235 //y=1.375
c173 ( 58 0 ) capacitor c=0.0149861f //x=25.235 //y=0.72
c174 ( 57 0 ) capacitor c=0.096037f //x=24.86 //y=1.915
c175 ( 56 0 ) capacitor c=0.0228993f //x=24.86 //y=1.53
c176 ( 55 0 ) capacitor c=0.0234352f //x=24.86 //y=1.22
c177 ( 54 0 ) capacitor c=0.0198724f //x=24.86 //y=0.875
c178 ( 53 0 ) capacitor c=0.110114f //x=25.8 //y=6.02
c179 ( 52 0 ) capacitor c=0.158956f //x=25.36 //y=6.02
c180 ( 50 0 ) capacitor c=0.00106608f //x=22.53 //y=5.155
c181 ( 49 0 ) capacitor c=0.00207319f //x=21.65 //y=5.155
c182 ( 42 0 ) capacitor c=0.0937944f //x=25.16 //y=2.08
c183 ( 40 0 ) capacitor c=0.103719f //x=23.31 //y=2.59
c184 ( 36 0 ) capacitor c=0.00398962f //x=22.91 //y=1.665
c185 ( 35 0 ) capacitor c=0.0137288f //x=23.225 //y=1.665
c186 ( 29 0 ) capacitor c=0.0283082f //x=23.225 //y=5.155
c187 ( 21 0 ) capacitor c=0.0176454f //x=22.445 //y=5.155
c188 ( 14 0 ) capacitor c=0.00332903f //x=20.855 //y=5.155
c189 ( 13 0 ) capacitor c=0.0148427f //x=21.565 //y=5.155
c190 ( 2 0 ) capacitor c=0.0116088f //x=23.425 //y=2.59
c191 ( 1 0 ) capacitor c=0.0352679f //x=25.045 //y=2.59
r192 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=25.725 //y=4.79 //x2=25.8 //y2=4.865
r193 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=25.725 //y=4.79 //x2=25.435 //y2=4.79
r194 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.39 //y=1.22 //x2=25.35 //y2=1.375
r195 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.39 //y=0.875 //x2=25.35 //y2=0.72
r196 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=25.39 //y=0.875 //x2=25.39 //y2=1.22
r197 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=25.36 //y=4.865 //x2=25.435 //y2=4.79
r198 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=25.36 //y=4.865 //x2=25.16 //y2=4.7
r199 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.015 //y=1.375 //x2=24.9 //y2=1.375
r200 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.235 //y=1.375 //x2=25.35 //y2=1.375
r201 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.015 //y=0.72 //x2=24.9 //y2=0.72
r202 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.235 //y=0.72 //x2=25.35 //y2=0.72
r203 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=25.235 //y=0.72 //x2=25.015 //y2=0.72
r204 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.915 //x2=25.16 //y2=2.08
r205 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.53 //x2=24.9 //y2=1.375
r206 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.53 //x2=24.86 //y2=1.915
r207 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.22 //x2=24.9 //y2=1.375
r208 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=0.875 //x2=24.9 //y2=0.72
r209 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.86 //y=0.875 //x2=24.86 //y2=1.22
r210 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.8 //y=6.02 //x2=25.8 //y2=4.865
r211 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.36 //y=6.02 //x2=25.36 //y2=4.865
r212 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.125 //y=1.375 //x2=25.235 //y2=1.375
r213 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.125 //y=1.375 //x2=25.015 //y2=1.375
r214 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.16 //y=4.7 //x2=25.16 //y2=4.7
r215 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.59 //x2=25.16 //y2=4.7
r216 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.16 //y=2.08 //x2=25.16 //y2=2.08
r217 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.08 //x2=25.16 //y2=2.59
r218 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=23.31 //y=5.07 //x2=23.31 //y2=2.59
r219 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=23.31 //y=1.75 //x2=23.31 //y2=2.59
r220 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.225 //y=1.665 //x2=23.31 //y2=1.75
r221 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=23.225 //y=1.665 //x2=22.91 //y2=1.665
r222 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=22.825 //y=1.58 //x2=22.91 //y2=1.665
r223 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=22.825 //y=1.58 //x2=22.825 //y2=1.01
r224 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.615 //y=5.155 //x2=22.53 //y2=5.155
r225 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.225 //y=5.155 //x2=23.31 //y2=5.07
r226 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=23.225 //y=5.155 //x2=22.615 //y2=5.155
r227 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.53 //y=5.24 //x2=22.53 //y2=5.155
r228 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.53 //y=5.24 //x2=22.53 //y2=5.725
r229 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.735 //y=5.155 //x2=21.65 //y2=5.155
r230 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.445 //y=5.155 //x2=22.53 //y2=5.155
r231 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.445 //y=5.155 //x2=21.735 //y2=5.155
r232 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.65 //y=5.24 //x2=21.65 //y2=5.155
r233 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.65 //y=5.24 //x2=21.65 //y2=5.725
r234 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.565 //y=5.155 //x2=21.65 //y2=5.155
r235 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=21.565 //y=5.155 //x2=20.855 //y2=5.155
r236 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.77 //y=5.24 //x2=20.855 //y2=5.155
r237 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.77 //y=5.24 //x2=20.77 //y2=5.725
r238 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.16 //y=2.59 //x2=25.16 //y2=2.59
r239 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.31 //y=2.59 //x2=23.31 //y2=2.59
r240 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.425 //y=2.59 //x2=23.31 //y2=2.59
r241 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.045 //y=2.59 //x2=25.16 //y2=2.59
r242 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=25.045 //y=2.59 //x2=23.425 //y2=2.59
ends PM_TMRDFFSNRNQX1\%noxref_6

subckt PM_TMRDFFSNRNQX1\%noxref_7 ( 1 2 3 4 5 6 16 24 37 38 45 53 59 60 64 66 \
 73 74 75 76 77 78 79 80 81 82 83 87 88 89 94 96 99 100 104 105 106 111 113 \
 116 117 121 122 123 128 130 133 134 136 137 142 146 147 152 156 157 162 165 \
 167 168 169 )
c338 ( 169 0 ) capacitor c=0.023087f //x=17.575 //y=5.02
c339 ( 168 0 ) capacitor c=0.023519f //x=16.695 //y=5.02
c340 ( 167 0 ) capacitor c=0.0224735f //x=15.815 //y=5.02
c341 ( 165 0 ) capacitor c=0.00853354f //x=17.825 //y=0.915
c342 ( 162 0 ) capacitor c=0.0587755f //x=27.38 //y=4.7
c343 ( 157 0 ) capacitor c=0.0273931f //x=27.38 //y=1.915
c344 ( 156 0 ) capacitor c=0.0456313f //x=27.38 //y=2.08
c345 ( 152 0 ) capacitor c=0.0587755f //x=12.95 //y=4.7
c346 ( 147 0 ) capacitor c=0.0273931f //x=12.95 //y=1.915
c347 ( 146 0 ) capacitor c=0.0456313f //x=12.95 //y=2.08
c348 ( 142 0 ) capacitor c=0.058931f //x=8.14 //y=4.7
c349 ( 137 0 ) capacitor c=0.0273931f //x=8.14 //y=1.915
c350 ( 136 0 ) capacitor c=0.0456313f //x=8.14 //y=2.08
c351 ( 134 0 ) capacitor c=0.0432517f //x=27.9 //y=1.26
c352 ( 133 0 ) capacitor c=0.0200379f //x=27.9 //y=0.915
c353 ( 130 0 ) capacitor c=0.0148873f //x=27.745 //y=1.415
c354 ( 128 0 ) capacitor c=0.0157803f //x=27.745 //y=0.76
c355 ( 123 0 ) capacitor c=0.0218028f //x=27.37 //y=1.57
c356 ( 122 0 ) capacitor c=0.0207459f //x=27.37 //y=1.26
c357 ( 121 0 ) capacitor c=0.0194308f //x=27.37 //y=0.915
c358 ( 117 0 ) capacitor c=0.0432517f //x=13.47 //y=1.26
c359 ( 116 0 ) capacitor c=0.0200379f //x=13.47 //y=0.915
c360 ( 113 0 ) capacitor c=0.0148873f //x=13.315 //y=1.415
c361 ( 111 0 ) capacitor c=0.0157803f //x=13.315 //y=0.76
c362 ( 106 0 ) capacitor c=0.0218028f //x=12.94 //y=1.57
c363 ( 105 0 ) capacitor c=0.0207459f //x=12.94 //y=1.26
c364 ( 104 0 ) capacitor c=0.0194308f //x=12.94 //y=0.915
c365 ( 100 0 ) capacitor c=0.0432517f //x=8.66 //y=1.26
c366 ( 99 0 ) capacitor c=0.0200379f //x=8.66 //y=0.915
c367 ( 96 0 ) capacitor c=0.0148873f //x=8.505 //y=1.415
c368 ( 94 0 ) capacitor c=0.0157803f //x=8.505 //y=0.76
c369 ( 89 0 ) capacitor c=0.0218028f //x=8.13 //y=1.57
c370 ( 88 0 ) capacitor c=0.0207459f //x=8.13 //y=1.26
c371 ( 87 0 ) capacitor c=0.0194308f //x=8.13 //y=0.915
c372 ( 83 0 ) capacitor c=0.158794f //x=27.56 //y=6.02
c373 ( 82 0 ) capacitor c=0.110114f //x=27.12 //y=6.02
c374 ( 81 0 ) capacitor c=0.158794f //x=13.13 //y=6.02
c375 ( 80 0 ) capacitor c=0.110114f //x=12.69 //y=6.02
c376 ( 79 0 ) capacitor c=0.158794f //x=8.32 //y=6.02
c377 ( 78 0 ) capacitor c=0.110114f //x=7.88 //y=6.02
c378 ( 74 0 ) capacitor c=0.00106608f //x=17.72 //y=5.155
c379 ( 73 0 ) capacitor c=0.00207162f //x=16.84 //y=5.155
c380 ( 66 0 ) capacitor c=0.0816644f //x=27.38 //y=2.08
c381 ( 64 0 ) capacitor c=0.105458f //x=18.5 //y=3.7
c382 ( 60 0 ) capacitor c=0.00398962f //x=18.1 //y=1.665
c383 ( 59 0 ) capacitor c=0.0137288f //x=18.415 //y=1.665
c384 ( 53 0 ) capacitor c=0.0283082f //x=18.415 //y=5.155
c385 ( 45 0 ) capacitor c=0.0176454f //x=17.635 //y=5.155
c386 ( 38 0 ) capacitor c=0.00332903f //x=16.045 //y=5.155
c387 ( 37 0 ) capacitor c=0.014837f //x=16.755 //y=5.155
c388 ( 24 0 ) capacitor c=0.0810736f //x=12.95 //y=2.08
c389 ( 16 0 ) capacitor c=0.0819749f //x=8.14 //y=2.08
c390 ( 6 0 ) capacitor c=0.0055354f //x=18.615 //y=3.7
c391 ( 5 0 ) capacitor c=0.146292f //x=27.265 //y=3.7
c392 ( 4 0 ) capacitor c=0.00556898f //x=13.065 //y=3.7
c393 ( 3 0 ) capacitor c=0.0758356f //x=18.385 //y=3.7
c394 ( 2 0 ) capacitor c=0.0138772f //x=8.255 //y=3.7
c395 ( 1 0 ) capacitor c=0.067053f //x=12.835 //y=3.7
r396 (  156 157 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=27.38 //y=2.08 //x2=27.38 //y2=1.915
r397 (  146 147 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=12.95 //y=2.08 //x2=12.95 //y2=1.915
r398 (  136 137 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.14 //y=2.08 //x2=8.14 //y2=1.915
r399 (  134 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.9 //y=1.26 //x2=27.86 //y2=1.415
r400 (  133 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.9 //y=0.915 //x2=27.86 //y2=0.76
r401 (  133 134 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.9 //y=0.915 //x2=27.9 //y2=1.26
r402 (  131 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.525 //y=1.415 //x2=27.41 //y2=1.415
r403 (  130 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.745 //y=1.415 //x2=27.86 //y2=1.415
r404 (  129 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.525 //y=0.76 //x2=27.41 //y2=0.76
r405 (  128 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.745 //y=0.76 //x2=27.86 //y2=0.76
r406 (  128 129 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=27.745 //y=0.76 //x2=27.525 //y2=0.76
r407 (  125 162 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=27.56 //y=4.865 //x2=27.38 //y2=4.7
r408 (  123 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.57 //x2=27.41 //y2=1.415
r409 (  123 157 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.57 //x2=27.37 //y2=1.915
r410 (  122 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.26 //x2=27.41 //y2=1.415
r411 (  121 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=0.915 //x2=27.41 //y2=0.76
r412 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.37 //y=0.915 //x2=27.37 //y2=1.26
r413 (  118 162 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=27.12 //y=4.865 //x2=27.38 //y2=4.7
r414 (  117 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.47 //y=1.26 //x2=13.43 //y2=1.415
r415 (  116 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.47 //y=0.915 //x2=13.43 //y2=0.76
r416 (  116 117 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.47 //y=0.915 //x2=13.47 //y2=1.26
r417 (  114 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.095 //y=1.415 //x2=12.98 //y2=1.415
r418 (  113 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.315 //y=1.415 //x2=13.43 //y2=1.415
r419 (  112 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.095 //y=0.76 //x2=12.98 //y2=0.76
r420 (  111 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.315 //y=0.76 //x2=13.43 //y2=0.76
r421 (  111 112 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=13.315 //y=0.76 //x2=13.095 //y2=0.76
r422 (  108 152 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=13.13 //y=4.865 //x2=12.95 //y2=4.7
r423 (  106 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.57 //x2=12.98 //y2=1.415
r424 (  106 147 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.57 //x2=12.94 //y2=1.915
r425 (  105 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.26 //x2=12.98 //y2=1.415
r426 (  104 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=0.915 //x2=12.98 //y2=0.76
r427 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.94 //y=0.915 //x2=12.94 //y2=1.26
r428 (  101 152 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=12.69 //y=4.865 //x2=12.95 //y2=4.7
r429 (  100 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=1.26 //x2=8.62 //y2=1.415
r430 (  99 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.62 //y2=0.76
r431 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.66 //y2=1.26
r432 (  97 140 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=1.415 //x2=8.17 //y2=1.415
r433 (  96 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=1.415 //x2=8.62 //y2=1.415
r434 (  95 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=0.76 //x2=8.17 //y2=0.76
r435 (  94 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.62 //y2=0.76
r436 (  94 95 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.285 //y2=0.76
r437 (  91 142 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=8.32 //y=4.865 //x2=8.14 //y2=4.7
r438 (  89 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.17 //y2=1.415
r439 (  89 137 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.13 //y2=1.915
r440 (  88 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.26 //x2=8.17 //y2=1.415
r441 (  87 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.17 //y2=0.76
r442 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.13 //y2=1.26
r443 (  84 142 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=7.88 //y=4.865 //x2=8.14 //y2=4.7
r444 (  83 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.56 //y=6.02 //x2=27.56 //y2=4.865
r445 (  82 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.12 //y=6.02 //x2=27.12 //y2=4.865
r446 (  81 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.13 //y=6.02 //x2=13.13 //y2=4.865
r447 (  80 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.69 //y=6.02 //x2=12.69 //y2=4.865
r448 (  79 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.32 //y=6.02 //x2=8.32 //y2=4.865
r449 (  78 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.88 //y=6.02 //x2=7.88 //y2=4.865
r450 (  77 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.635 //y=1.415 //x2=27.745 //y2=1.415
r451 (  77 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.635 //y=1.415 //x2=27.525 //y2=1.415
r452 (  76 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.205 //y=1.415 //x2=13.315 //y2=1.415
r453 (  76 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.205 //y=1.415 //x2=13.095 //y2=1.415
r454 (  75 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.505 //y2=1.415
r455 (  75 97 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.285 //y2=1.415
r456 (  71 162 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=4.7 //x2=27.38 //y2=4.7
r457 (  69 71 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=27.38 //y=3.7 //x2=27.38 //y2=4.7
r458 (  66 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=2.08 //x2=27.38 //y2=2.08
r459 (  66 69 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=27.38 //y=2.08 //x2=27.38 //y2=3.7
r460 (  62 64 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=18.5 //y=5.07 //x2=18.5 //y2=3.7
r461 (  61 64 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=18.5 //y=1.75 //x2=18.5 //y2=3.7
r462 (  59 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.415 //y=1.665 //x2=18.5 //y2=1.75
r463 (  59 60 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=18.415 //y=1.665 //x2=18.1 //y2=1.665
r464 (  55 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.015 //y=1.58 //x2=18.1 //y2=1.665
r465 (  55 165 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=18.015 //y=1.58 //x2=18.015 //y2=1.01
r466 (  54 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.805 //y=5.155 //x2=17.72 //y2=5.155
r467 (  53 62 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.415 //y=5.155 //x2=18.5 //y2=5.07
r468 (  53 54 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=18.415 //y=5.155 //x2=17.805 //y2=5.155
r469 (  47 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.72 //y=5.24 //x2=17.72 //y2=5.155
r470 (  47 169 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.72 //y=5.24 //x2=17.72 //y2=5.725
r471 (  46 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.925 //y=5.155 //x2=16.84 //y2=5.155
r472 (  45 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.635 //y=5.155 //x2=17.72 //y2=5.155
r473 (  45 46 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=17.635 //y=5.155 //x2=16.925 //y2=5.155
r474 (  39 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.84 //y=5.24 //x2=16.84 //y2=5.155
r475 (  39 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.84 //y=5.24 //x2=16.84 //y2=5.725
r476 (  37 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.755 //y=5.155 //x2=16.84 //y2=5.155
r477 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.755 //y=5.155 //x2=16.045 //y2=5.155
r478 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.96 //y=5.24 //x2=16.045 //y2=5.155
r479 (  31 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.96 //y=5.24 //x2=15.96 //y2=5.725
r480 (  29 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.95 //y=4.7 //x2=12.95 //y2=4.7
r481 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=12.95 //y=3.7 //x2=12.95 //y2=4.7
r482 (  24 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.95 //y=2.08 //x2=12.95 //y2=2.08
r483 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=12.95 //y=2.08 //x2=12.95 //y2=3.7
r484 (  21 142 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=4.7 //x2=8.14 //y2=4.7
r485 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=8.14 //y=3.7 //x2=8.14 //y2=4.7
r486 (  16 136 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=2.08 //x2=8.14 //y2=2.08
r487 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.08 //x2=8.14 //y2=3.7
r488 (  14 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=27.38 //y=3.7 //x2=27.38 //y2=3.7
r489 (  12 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.5 //y=3.7 //x2=18.5 //y2=3.7
r490 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.95 //y=3.7 //x2=12.95 //y2=3.7
r491 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.14 //y=3.7 //x2=8.14 //y2=3.7
r492 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.615 //y=3.7 //x2=18.5 //y2=3.7
r493 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.265 //y=3.7 //x2=27.38 //y2=3.7
r494 (  5 6 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=27.265 //y=3.7 //x2=18.615 //y2=3.7
r495 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.065 //y=3.7 //x2=12.95 //y2=3.7
r496 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=3.7 //x2=18.5 //y2=3.7
r497 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=3.7 //x2=13.065 //y2=3.7
r498 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.255 //y=3.7 //x2=8.14 //y2=3.7
r499 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.835 //y=3.7 //x2=12.95 //y2=3.7
r500 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=12.835 //y=3.7 //x2=8.255 //y2=3.7
ends PM_TMRDFFSNRNQX1\%noxref_7

subckt PM_TMRDFFSNRNQX1\%noxref_8 ( 1 2 3 4 6 7 8 9 10 22 35 36 43 51 57 58 62 \
 66 74 81 82 83 84 85 86 87 88 89 90 91 95 96 97 102 104 107 108 109 110 111 \
 112 116 118 121 122 123 124 128 129 130 131 135 137 143 144 146 147 152 156 \
 169 172 174 175 176 )
c629 ( 176 0 ) capacitor c=0.023087f //x=27.195 //y=5.02
c630 ( 175 0 ) capacitor c=0.023519f //x=26.315 //y=5.02
c631 ( 174 0 ) capacitor c=0.0224735f //x=25.435 //y=5.02
c632 ( 172 0 ) capacitor c=0.00853354f //x=27.445 //y=0.915
c633 ( 169 0 ) capacitor c=0.0655948f //x=91.02 //y=4.705
c634 ( 156 0 ) capacitor c=0.054113f //x=87.32 //y=2.08
c635 ( 152 0 ) capacitor c=0.0587755f //x=22.57 //y=4.7
c636 ( 147 0 ) capacitor c=0.0273931f //x=22.57 //y=1.915
c637 ( 146 0 ) capacitor c=0.0456313f //x=22.57 //y=2.08
c638 ( 144 0 ) capacitor c=0.0342409f //x=91.355 //y=1.21
c639 ( 143 0 ) capacitor c=0.0187384f //x=91.355 //y=0.865
c640 ( 137 0 ) capacitor c=0.0141797f //x=91.2 //y=1.365
c641 ( 135 0 ) capacitor c=0.0149844f //x=91.2 //y=0.71
c642 ( 131 0 ) capacitor c=0.0954119f //x=90.825 //y=1.915
c643 ( 130 0 ) capacitor c=0.022465f //x=90.825 //y=1.52
c644 ( 129 0 ) capacitor c=0.0234376f //x=90.825 //y=1.21
c645 ( 128 0 ) capacitor c=0.0199343f //x=90.825 //y=0.865
c646 ( 124 0 ) capacitor c=0.0318948f //x=88.025 //y=1.21
c647 ( 123 0 ) capacitor c=0.0187384f //x=88.025 //y=0.865
c648 ( 122 0 ) capacitor c=0.0605713f //x=87.665 //y=4.795
c649 ( 121 0 ) capacitor c=0.0292043f //x=87.955 //y=4.795
c650 ( 118 0 ) capacitor c=0.0157913f //x=87.87 //y=1.365
c651 ( 116 0 ) capacitor c=0.0149844f //x=87.87 //y=0.71
c652 ( 112 0 ) capacitor c=0.0302441f //x=87.495 //y=1.915
c653 ( 111 0 ) capacitor c=0.0237559f //x=87.495 //y=1.52
c654 ( 110 0 ) capacitor c=0.0234352f //x=87.495 //y=1.21
c655 ( 109 0 ) capacitor c=0.0199931f //x=87.495 //y=0.865
c656 ( 108 0 ) capacitor c=0.0432517f //x=23.09 //y=1.26
c657 ( 107 0 ) capacitor c=0.0200379f //x=23.09 //y=0.915
c658 ( 104 0 ) capacitor c=0.0148873f //x=22.935 //y=1.415
c659 ( 102 0 ) capacitor c=0.0157803f //x=22.935 //y=0.76
c660 ( 97 0 ) capacitor c=0.0218028f //x=22.56 //y=1.57
c661 ( 96 0 ) capacitor c=0.0207459f //x=22.56 //y=1.26
c662 ( 95 0 ) capacitor c=0.0194308f //x=22.56 //y=0.915
c663 ( 91 0 ) capacitor c=0.110336f //x=91.35 //y=6.025
c664 ( 90 0 ) capacitor c=0.154049f //x=90.91 //y=6.025
c665 ( 89 0 ) capacitor c=0.110003f //x=88.03 //y=6.025
c666 ( 88 0 ) capacitor c=0.15424f //x=87.59 //y=6.025
c667 ( 87 0 ) capacitor c=0.158794f //x=22.75 //y=6.02
c668 ( 86 0 ) capacitor c=0.110114f //x=22.31 //y=6.02
c669 ( 82 0 ) capacitor c=0.00106608f //x=27.34 //y=5.155
c670 ( 81 0 ) capacitor c=0.00207319f //x=26.46 //y=5.155
c671 ( 74 0 ) capacitor c=0.119551f //x=91.02 //y=2.08
c672 ( 66 0 ) capacitor c=0.0994818f //x=87.32 //y=2.08
c673 ( 62 0 ) capacitor c=0.106944f //x=28.12 //y=3.33
c674 ( 58 0 ) capacitor c=0.00398962f //x=27.72 //y=1.665
c675 ( 57 0 ) capacitor c=0.0137288f //x=28.035 //y=1.665
c676 ( 51 0 ) capacitor c=0.0282124f //x=28.035 //y=5.155
c677 ( 43 0 ) capacitor c=0.0176454f //x=27.255 //y=5.155
c678 ( 36 0 ) capacitor c=0.00332903f //x=25.665 //y=5.155
c679 ( 35 0 ) capacitor c=0.0148427f //x=26.375 //y=5.155
c680 ( 22 0 ) capacitor c=0.0820026f //x=22.57 //y=2.08
c681 ( 10 0 ) capacitor c=0.00638553f //x=87.435 //y=4.44
c682 ( 9 0 ) capacitor c=0.0799095f //x=90.905 //y=4.44
c683 ( 8 0 ) capacitor c=0.00309768f //x=75.195 //y=4.44
c684 ( 7 0 ) capacitor c=0.267484f //x=87.205 //y=4.44
c685 ( 6 0 ) capacitor c=0.00718365f //x=75.11 //y=4.725
c686 ( 4 0 ) capacitor c=0.0158574f //x=28.235 //y=4.81
c687 ( 3 0 ) capacitor c=0.852749f //x=75.025 //y=4.81
c688 ( 2 0 ) capacitor c=0.00906635f //x=22.685 //y=3.33
c689 ( 1 0 ) capacitor c=0.0889942f //x=28.005 //y=3.33
r690 (  167 169 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=90.91 //y=4.705 //x2=91.02 //y2=4.705
r691 (  146 147 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=22.57 //y=2.08 //x2=22.57 //y2=1.915
r692 (  144 171 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=91.355 //y=1.21 //x2=91.315 //y2=1.365
r693 (  143 170 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=91.355 //y=0.865 //x2=91.315 //y2=0.71
r694 (  143 144 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=91.355 //y=0.865 //x2=91.355 //y2=1.21
r695 (  140 169 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=91.35 //y=4.87 //x2=91.02 //y2=4.705
r696 (  138 166 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=90.98 //y=1.365 //x2=90.865 //y2=1.365
r697 (  137 171 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=91.2 //y=1.365 //x2=91.315 //y2=1.365
r698 (  136 165 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=90.98 //y=0.71 //x2=90.865 //y2=0.71
r699 (  135 170 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=91.2 //y=0.71 //x2=91.315 //y2=0.71
r700 (  135 136 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=91.2 //y=0.71 //x2=90.98 //y2=0.71
r701 (  132 167 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=90.91 //y=4.87 //x2=90.91 //y2=4.705
r702 (  131 164 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=90.825 //y=1.915 //x2=91.02 //y2=2.08
r703 (  130 166 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=90.825 //y=1.52 //x2=90.865 //y2=1.365
r704 (  130 131 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=90.825 //y=1.52 //x2=90.825 //y2=1.915
r705 (  129 166 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=90.825 //y=1.21 //x2=90.865 //y2=1.365
r706 (  128 165 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=90.825 //y=0.865 //x2=90.865 //y2=0.71
r707 (  128 129 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=90.825 //y=0.865 //x2=90.825 //y2=1.21
r708 (  124 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.025 //y=1.21 //x2=87.985 //y2=1.365
r709 (  123 161 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.025 //y=0.865 //x2=87.985 //y2=0.71
r710 (  123 124 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=88.025 //y=0.865 //x2=88.025 //y2=1.21
r711 (  121 125 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=87.955 //y=4.795 //x2=88.03 //y2=4.87
r712 (  121 122 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=87.955 //y=4.795 //x2=87.665 //y2=4.795
r713 (  119 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=87.65 //y=1.365 //x2=87.535 //y2=1.365
r714 (  118 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=87.87 //y=1.365 //x2=87.985 //y2=1.365
r715 (  117 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=87.65 //y=0.71 //x2=87.535 //y2=0.71
r716 (  116 161 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=87.87 //y=0.71 //x2=87.985 //y2=0.71
r717 (  116 117 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=87.87 //y=0.71 //x2=87.65 //y2=0.71
r718 (  113 122 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=87.59 //y=4.87 //x2=87.665 //y2=4.795
r719 (  113 158 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=87.59 //y=4.87 //x2=87.32 //y2=4.705
r720 (  112 156 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=87.495 //y=1.915 //x2=87.32 //y2=2.08
r721 (  111 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=87.495 //y=1.52 //x2=87.535 //y2=1.365
r722 (  111 112 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=87.495 //y=1.52 //x2=87.495 //y2=1.915
r723 (  110 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=87.495 //y=1.21 //x2=87.535 //y2=1.365
r724 (  109 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=87.495 //y=0.865 //x2=87.535 //y2=0.71
r725 (  109 110 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=87.495 //y=0.865 //x2=87.495 //y2=1.21
r726 (  108 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.09 //y=1.26 //x2=23.05 //y2=1.415
r727 (  107 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.09 //y=0.915 //x2=23.05 //y2=0.76
r728 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.09 //y=0.915 //x2=23.09 //y2=1.26
r729 (  105 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.715 //y=1.415 //x2=22.6 //y2=1.415
r730 (  104 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.935 //y=1.415 //x2=23.05 //y2=1.415
r731 (  103 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.715 //y=0.76 //x2=22.6 //y2=0.76
r732 (  102 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.935 //y=0.76 //x2=23.05 //y2=0.76
r733 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=22.935 //y=0.76 //x2=22.715 //y2=0.76
r734 (  99 152 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=22.75 //y=4.865 //x2=22.57 //y2=4.7
r735 (  97 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.57 //x2=22.6 //y2=1.415
r736 (  97 147 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.57 //x2=22.56 //y2=1.915
r737 (  96 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.26 //x2=22.6 //y2=1.415
r738 (  95 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=0.915 //x2=22.6 //y2=0.76
r739 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.56 //y=0.915 //x2=22.56 //y2=1.26
r740 (  92 152 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=22.31 //y=4.865 //x2=22.57 //y2=4.7
r741 (  91 140 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=91.35 //y=6.025 //x2=91.35 //y2=4.87
r742 (  90 132 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=90.91 //y=6.025 //x2=90.91 //y2=4.87
r743 (  89 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=88.03 //y=6.025 //x2=88.03 //y2=4.87
r744 (  88 113 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=87.59 //y=6.025 //x2=87.59 //y2=4.87
r745 (  87 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.75 //y=6.02 //x2=22.75 //y2=4.865
r746 (  86 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.31 //y=6.02 //x2=22.31 //y2=4.865
r747 (  85 137 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=91.09 //y=1.365 //x2=91.2 //y2=1.365
r748 (  85 138 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=91.09 //y=1.365 //x2=90.98 //y2=1.365
r749 (  84 118 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=87.76 //y=1.365 //x2=87.87 //y2=1.365
r750 (  84 119 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=87.76 //y=1.365 //x2=87.65 //y2=1.365
r751 (  83 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.825 //y=1.415 //x2=22.935 //y2=1.415
r752 (  83 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.825 //y=1.415 //x2=22.715 //y2=1.415
r753 (  79 169 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=91.02 //y=4.705 //x2=91.02 //y2=4.705
r754 (  77 79 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=91.02 //y=4.44 //x2=91.02 //y2=4.705
r755 (  74 164 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=91.02 //y=2.08 //x2=91.02 //y2=2.08
r756 (  74 77 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=91.02 //y=2.08 //x2=91.02 //y2=4.44
r757 (  71 158 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=87.32 //y=4.705 //x2=87.32 //y2=4.705
r758 (  69 71 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=87.32 //y=4.44 //x2=87.32 //y2=4.705
r759 (  66 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=87.32 //y=2.08 //x2=87.32 //y2=2.08
r760 (  66 69 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=87.32 //y=2.08 //x2=87.32 //y2=4.44
r761 (  62 64 ) resistor r=101.305 //w=0.187 //l=1.48 //layer=li \
 //thickness=0.1 //x=28.12 //y=3.33 //x2=28.12 //y2=4.81
r762 (  60 64 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=28.12 //y=5.07 //x2=28.12 //y2=4.81
r763 (  59 62 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=28.12 //y=1.75 //x2=28.12 //y2=3.33
r764 (  57 59 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.035 //y=1.665 //x2=28.12 //y2=1.75
r765 (  57 58 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=28.035 //y=1.665 //x2=27.72 //y2=1.665
r766 (  53 58 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=27.635 //y=1.58 //x2=27.72 //y2=1.665
r767 (  53 172 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=27.635 //y=1.58 //x2=27.635 //y2=1.01
r768 (  52 82 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.425 //y=5.155 //x2=27.34 //y2=5.155
r769 (  51 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.035 //y=5.155 //x2=28.12 //y2=5.07
r770 (  51 52 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=28.035 //y=5.155 //x2=27.425 //y2=5.155
r771 (  45 82 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.34 //y=5.24 //x2=27.34 //y2=5.155
r772 (  45 176 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.34 //y=5.24 //x2=27.34 //y2=5.725
r773 (  44 81 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.545 //y=5.155 //x2=26.46 //y2=5.155
r774 (  43 82 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.255 //y=5.155 //x2=27.34 //y2=5.155
r775 (  43 44 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=27.255 //y=5.155 //x2=26.545 //y2=5.155
r776 (  37 81 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.46 //y=5.24 //x2=26.46 //y2=5.155
r777 (  37 175 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.46 //y=5.24 //x2=26.46 //y2=5.725
r778 (  35 81 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.375 //y=5.155 //x2=26.46 //y2=5.155
r779 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.375 //y=5.155 //x2=25.665 //y2=5.155
r780 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.58 //y=5.24 //x2=25.665 //y2=5.155
r781 (  29 174 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=25.58 //y=5.24 //x2=25.58 //y2=5.725
r782 (  27 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=4.7 //x2=22.57 //y2=4.7
r783 (  25 27 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=22.57 //y=3.33 //x2=22.57 //y2=4.7
r784 (  22 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=2.08 //x2=22.57 //y2=2.08
r785 (  22 25 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=22.57 //y=2.08 //x2=22.57 //y2=3.33
r786 (  20 77 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=91.02 //y=4.44 //x2=91.02 //y2=4.44
r787 (  18 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=87.32 //y=4.44 //x2=87.32 //y2=4.44
r788 (  16 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.12 //y=3.33 //x2=28.12 //y2=3.33
r789 (  14 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.12 //y=4.81 //x2=28.12 //y2=4.81
r790 (  12 25 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=22.57 //y=3.33 //x2=22.57 //y2=3.33
r791 (  10 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=87.435 //y=4.44 //x2=87.32 //y2=4.44
r792 (  9 20 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=90.905 //y=4.44 //x2=91.02 //y2=4.44
r793 (  9 10 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=90.905 //y=4.44 //x2=87.435 //y2=4.44
r794 (  7 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=87.205 //y=4.44 //x2=87.32 //y2=4.44
r795 (  7 8 ) resistor r=11.4599 //w=0.131 //l=12.01 //layer=m1 \
 //thickness=0.36 //x=87.205 //y=4.44 //x2=75.195 //y2=4.44
r796 (  5 8 ) resistor r=0.0718295 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=4.525 //x2=75.195 //y2=4.44
r797 (  5 6 ) resistor r=0.19084 //w=0.131 //l=0.2 //layer=m1 //thickness=0.36 \
 //x=75.11 //y=4.525 //x2=75.11 //y2=4.725
r798 (  4 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.235 //y=4.81 //x2=28.12 //y2=4.81
r799 (  3 6 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=75.025 //y=4.81 //x2=75.11 //y2=4.725
r800 (  3 4 ) resistor r=44.6469 //w=0.131 //l=46.79 //layer=m1 \
 //thickness=0.36 //x=75.025 //y=4.81 //x2=28.235 //y2=4.81
r801 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=22.685 //y=3.33 //x2=22.57 //y2=3.33
r802 (  1 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=3.33 //x2=28.12 //y2=3.33
r803 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=3.33 //x2=22.685 //y2=3.33
ends PM_TMRDFFSNRNQX1\%noxref_8

subckt PM_TMRDFFSNRNQX1\%noxref_9 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 \
 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c253 ( 127 0 ) capacitor c=0.023087f //x=32.005 //y=5.02
c254 ( 126 0 ) capacitor c=0.023519f //x=31.125 //y=5.02
c255 ( 125 0 ) capacitor c=0.0224735f //x=30.245 //y=5.02
c256 ( 123 0 ) capacitor c=0.00853354f //x=32.255 //y=0.915
c257 ( 103 0 ) capacitor c=0.0547611f //x=39.865 //y=4.79
c258 ( 102 0 ) capacitor c=0.0294456f //x=40.155 //y=4.79
c259 ( 101 0 ) capacitor c=0.0347816f //x=39.82 //y=1.22
c260 ( 100 0 ) capacitor c=0.0187487f //x=39.82 //y=0.875
c261 ( 94 0 ) capacitor c=0.0137055f //x=39.665 //y=1.375
c262 ( 92 0 ) capacitor c=0.0149861f //x=39.665 //y=0.72
c263 ( 91 0 ) capacitor c=0.096037f //x=39.29 //y=1.915
c264 ( 90 0 ) capacitor c=0.0228993f //x=39.29 //y=1.53
c265 ( 89 0 ) capacitor c=0.0234352f //x=39.29 //y=1.22
c266 ( 88 0 ) capacitor c=0.0198724f //x=39.29 //y=0.875
c267 ( 84 0 ) capacitor c=0.0549166f //x=35.055 //y=4.79
c268 ( 83 0 ) capacitor c=0.0294456f //x=35.345 //y=4.79
c269 ( 82 0 ) capacitor c=0.0347816f //x=35.01 //y=1.22
c270 ( 81 0 ) capacitor c=0.0187487f //x=35.01 //y=0.875
c271 ( 75 0 ) capacitor c=0.0137055f //x=34.855 //y=1.375
c272 ( 73 0 ) capacitor c=0.0149861f //x=34.855 //y=0.72
c273 ( 72 0 ) capacitor c=0.096037f //x=34.48 //y=1.915
c274 ( 71 0 ) capacitor c=0.0228993f //x=34.48 //y=1.53
c275 ( 70 0 ) capacitor c=0.0234352f //x=34.48 //y=1.22
c276 ( 69 0 ) capacitor c=0.0198724f //x=34.48 //y=0.875
c277 ( 68 0 ) capacitor c=0.109949f //x=40.23 //y=6.02
c278 ( 67 0 ) capacitor c=0.158483f //x=39.79 //y=6.02
c279 ( 66 0 ) capacitor c=0.109949f //x=35.42 //y=6.02
c280 ( 65 0 ) capacitor c=0.158483f //x=34.98 //y=6.02
c281 ( 62 0 ) capacitor c=9.74268e-19 //x=32.15 //y=5.155
c282 ( 61 0 ) capacitor c=0.00191414f //x=31.27 //y=5.155
c283 ( 54 0 ) capacitor c=0.0914984f //x=39.59 //y=2.08
c284 ( 46 0 ) capacitor c=0.0942434f //x=34.78 //y=2.08
c285 ( 44 0 ) capacitor c=0.106133f //x=32.93 //y=2.59
c286 ( 40 0 ) capacitor c=0.00398962f //x=32.53 //y=1.665
c287 ( 39 0 ) capacitor c=0.0137288f //x=32.845 //y=1.665
c288 ( 33 0 ) capacitor c=0.0276208f //x=32.845 //y=5.155
c289 ( 25 0 ) capacitor c=0.0169868f //x=32.065 //y=5.155
c290 ( 18 0 ) capacitor c=0.00316998f //x=30.475 //y=5.155
c291 ( 17 0 ) capacitor c=0.014258f //x=31.185 //y=5.155
c292 ( 4 0 ) capacitor c=0.00401138f //x=34.895 //y=2.59
c293 ( 3 0 ) capacitor c=0.0706637f //x=39.475 //y=2.59
c294 ( 2 0 ) capacitor c=0.0120752f //x=33.045 //y=2.59
c295 ( 1 0 ) capacitor c=0.0233554f //x=34.665 //y=2.59
r296 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=40.155 //y=4.79 //x2=40.23 //y2=4.865
r297 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=40.155 //y=4.79 //x2=39.865 //y2=4.79
r298 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.82 //y=1.22 //x2=39.78 //y2=1.375
r299 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.82 //y=0.875 //x2=39.78 //y2=0.72
r300 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=39.82 //y=0.875 //x2=39.82 //y2=1.22
r301 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=39.79 //y=4.865 //x2=39.865 //y2=4.79
r302 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=39.79 //y=4.865 //x2=39.59 //y2=4.7
r303 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.445 //y=1.375 //x2=39.33 //y2=1.375
r304 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.665 //y=1.375 //x2=39.78 //y2=1.375
r305 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.445 //y=0.72 //x2=39.33 //y2=0.72
r306 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.665 //y=0.72 //x2=39.78 //y2=0.72
r307 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=39.665 //y=0.72 //x2=39.445 //y2=0.72
r308 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=39.29 //y=1.915 //x2=39.59 //y2=2.08
r309 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.29 //y=1.53 //x2=39.33 //y2=1.375
r310 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=39.29 //y=1.53 //x2=39.29 //y2=1.915
r311 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.29 //y=1.22 //x2=39.33 //y2=1.375
r312 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.29 //y=0.875 //x2=39.33 //y2=0.72
r313 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=39.29 //y=0.875 //x2=39.29 //y2=1.22
r314 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=35.345 //y=4.79 //x2=35.42 //y2=4.865
r315 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=35.345 //y=4.79 //x2=35.055 //y2=4.79
r316 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.01 //y=1.22 //x2=34.97 //y2=1.375
r317 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.01 //y=0.875 //x2=34.97 //y2=0.72
r318 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=35.01 //y=0.875 //x2=35.01 //y2=1.22
r319 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=34.98 //y=4.865 //x2=35.055 //y2=4.79
r320 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=34.98 //y=4.865 //x2=34.78 //y2=4.7
r321 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.635 //y=1.375 //x2=34.52 //y2=1.375
r322 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.855 //y=1.375 //x2=34.97 //y2=1.375
r323 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.635 //y=0.72 //x2=34.52 //y2=0.72
r324 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.855 //y=0.72 //x2=34.97 //y2=0.72
r325 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=34.855 //y=0.72 //x2=34.635 //y2=0.72
r326 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.915 //x2=34.78 //y2=2.08
r327 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.53 //x2=34.52 //y2=1.375
r328 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.53 //x2=34.48 //y2=1.915
r329 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.22 //x2=34.52 //y2=1.375
r330 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.48 //y=0.875 //x2=34.52 //y2=0.72
r331 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=34.48 //y=0.875 //x2=34.48 //y2=1.22
r332 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=40.23 //y=6.02 //x2=40.23 //y2=4.865
r333 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=39.79 //y=6.02 //x2=39.79 //y2=4.865
r334 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.42 //y=6.02 //x2=35.42 //y2=4.865
r335 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.98 //y=6.02 //x2=34.98 //y2=4.865
r336 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.555 //y=1.375 //x2=39.665 //y2=1.375
r337 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.555 //y=1.375 //x2=39.445 //y2=1.375
r338 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.745 //y=1.375 //x2=34.855 //y2=1.375
r339 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.745 //y=1.375 //x2=34.635 //y2=1.375
r340 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.59 //y=4.7 //x2=39.59 //y2=4.7
r341 (  57 59 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=39.59 //y=2.59 //x2=39.59 //y2=4.7
r342 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.59 //y=2.08 //x2=39.59 //y2=2.08
r343 (  54 57 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=39.59 //y=2.08 //x2=39.59 //y2=2.59
r344 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.78 //y=4.7 //x2=34.78 //y2=4.7
r345 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=34.78 //y=2.59 //x2=34.78 //y2=4.7
r346 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.78 //y=2.08 //x2=34.78 //y2=2.08
r347 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=34.78 //y=2.08 //x2=34.78 //y2=2.59
r348 (  42 44 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=32.93 //y=5.07 //x2=32.93 //y2=2.59
r349 (  41 44 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=32.93 //y=1.75 //x2=32.93 //y2=2.59
r350 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.845 //y=1.665 //x2=32.93 //y2=1.75
r351 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=32.845 //y=1.665 //x2=32.53 //y2=1.665
r352 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.445 //y=1.58 //x2=32.53 //y2=1.665
r353 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=32.445 //y=1.58 //x2=32.445 //y2=1.01
r354 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.235 //y=5.155 //x2=32.15 //y2=5.155
r355 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.845 //y=5.155 //x2=32.93 //y2=5.07
r356 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=32.845 //y=5.155 //x2=32.235 //y2=5.155
r357 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.15 //y=5.24 //x2=32.15 //y2=5.155
r358 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=32.15 //y=5.24 //x2=32.15 //y2=5.725
r359 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.355 //y=5.155 //x2=31.27 //y2=5.155
r360 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.065 //y=5.155 //x2=32.15 //y2=5.155
r361 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=32.065 //y=5.155 //x2=31.355 //y2=5.155
r362 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.27 //y=5.24 //x2=31.27 //y2=5.155
r363 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.27 //y=5.24 //x2=31.27 //y2=5.725
r364 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.185 //y=5.155 //x2=31.27 //y2=5.155
r365 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=31.185 //y=5.155 //x2=30.475 //y2=5.155
r366 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=30.39 //y=5.24 //x2=30.475 //y2=5.155
r367 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=30.39 //y=5.24 //x2=30.39 //y2=5.725
r368 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=39.59 //y=2.59 //x2=39.59 //y2=2.59
r369 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=34.78 //y=2.59 //x2=34.78 //y2=2.59
r370 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=32.93 //y=2.59 //x2=32.93 //y2=2.59
r371 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.895 //y=2.59 //x2=34.78 //y2=2.59
r372 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=39.475 //y=2.59 //x2=39.59 //y2=2.59
r373 (  3 4 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=39.475 //y=2.59 //x2=34.895 //y2=2.59
r374 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=33.045 //y=2.59 //x2=32.93 //y2=2.59
r375 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=2.59 //x2=34.78 //y2=2.59
r376 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=34.665 //y=2.59 //x2=33.045 //y2=2.59
ends PM_TMRDFFSNRNQX1\%noxref_9

subckt PM_TMRDFFSNRNQX1\%noxref_10 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 \
 53 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c169 ( 85 0 ) capacitor c=0.023087f //x=41.625 //y=5.02
c170 ( 84 0 ) capacitor c=0.023519f //x=40.745 //y=5.02
c171 ( 83 0 ) capacitor c=0.0224735f //x=39.865 //y=5.02
c172 ( 81 0 ) capacitor c=0.00853354f //x=41.875 //y=0.915
c173 ( 69 0 ) capacitor c=0.0549166f //x=44.675 //y=4.79
c174 ( 68 0 ) capacitor c=0.0294456f //x=44.965 //y=4.79
c175 ( 67 0 ) capacitor c=0.0347816f //x=44.63 //y=1.22
c176 ( 66 0 ) capacitor c=0.0187487f //x=44.63 //y=0.875
c177 ( 60 0 ) capacitor c=0.0137055f //x=44.475 //y=1.375
c178 ( 58 0 ) capacitor c=0.0149861f //x=44.475 //y=0.72
c179 ( 57 0 ) capacitor c=0.096037f //x=44.1 //y=1.915
c180 ( 56 0 ) capacitor c=0.0228993f //x=44.1 //y=1.53
c181 ( 55 0 ) capacitor c=0.0234352f //x=44.1 //y=1.22
c182 ( 54 0 ) capacitor c=0.0198724f //x=44.1 //y=0.875
c183 ( 53 0 ) capacitor c=0.109949f //x=45.04 //y=6.02
c184 ( 52 0 ) capacitor c=0.158483f //x=44.6 //y=6.02
c185 ( 50 0 ) capacitor c=9.74268e-19 //x=41.77 //y=5.155
c186 ( 49 0 ) capacitor c=0.00191414f //x=40.89 //y=5.155
c187 ( 42 0 ) capacitor c=0.0911502f //x=44.4 //y=2.08
c188 ( 40 0 ) capacitor c=0.103494f //x=42.55 //y=2.59
c189 ( 36 0 ) capacitor c=0.00398962f //x=42.15 //y=1.665
c190 ( 35 0 ) capacitor c=0.0137288f //x=42.465 //y=1.665
c191 ( 29 0 ) capacitor c=0.0276208f //x=42.465 //y=5.155
c192 ( 21 0 ) capacitor c=0.0169868f //x=41.685 //y=5.155
c193 ( 14 0 ) capacitor c=0.00316998f //x=40.095 //y=5.155
c194 ( 13 0 ) capacitor c=0.014258f //x=40.805 //y=5.155
c195 ( 2 0 ) capacitor c=0.00808366f //x=42.665 //y=2.59
c196 ( 1 0 ) capacitor c=0.0351856f //x=44.285 //y=2.59
r197 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=44.965 //y=4.79 //x2=45.04 //y2=4.865
r198 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=44.965 //y=4.79 //x2=44.675 //y2=4.79
r199 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.63 //y=1.22 //x2=44.59 //y2=1.375
r200 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.63 //y=0.875 //x2=44.59 //y2=0.72
r201 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=44.63 //y=0.875 //x2=44.63 //y2=1.22
r202 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=44.6 //y=4.865 //x2=44.675 //y2=4.79
r203 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=44.6 //y=4.865 //x2=44.4 //y2=4.7
r204 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.255 //y=1.375 //x2=44.14 //y2=1.375
r205 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.475 //y=1.375 //x2=44.59 //y2=1.375
r206 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.255 //y=0.72 //x2=44.14 //y2=0.72
r207 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.475 //y=0.72 //x2=44.59 //y2=0.72
r208 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=44.475 //y=0.72 //x2=44.255 //y2=0.72
r209 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=44.1 //y=1.915 //x2=44.4 //y2=2.08
r210 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.1 //y=1.53 //x2=44.14 //y2=1.375
r211 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=44.1 //y=1.53 //x2=44.1 //y2=1.915
r212 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.1 //y=1.22 //x2=44.14 //y2=1.375
r213 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.1 //y=0.875 //x2=44.14 //y2=0.72
r214 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=44.1 //y=0.875 //x2=44.1 //y2=1.22
r215 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.04 //y=6.02 //x2=45.04 //y2=4.865
r216 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=44.6 //y=6.02 //x2=44.6 //y2=4.865
r217 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=44.365 //y=1.375 //x2=44.475 //y2=1.375
r218 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=44.365 //y=1.375 //x2=44.255 //y2=1.375
r219 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=44.4 //y=4.7 //x2=44.4 //y2=4.7
r220 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=44.4 //y=2.59 //x2=44.4 //y2=4.7
r221 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=44.4 //y=2.08 //x2=44.4 //y2=2.08
r222 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=44.4 //y=2.08 //x2=44.4 //y2=2.59
r223 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=42.55 //y=5.07 //x2=42.55 //y2=2.59
r224 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=42.55 //y=1.75 //x2=42.55 //y2=2.59
r225 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.465 //y=1.665 //x2=42.55 //y2=1.75
r226 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=42.465 //y=1.665 //x2=42.15 //y2=1.665
r227 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.065 //y=1.58 //x2=42.15 //y2=1.665
r228 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=42.065 //y=1.58 //x2=42.065 //y2=1.01
r229 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.855 //y=5.155 //x2=41.77 //y2=5.155
r230 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.465 //y=5.155 //x2=42.55 //y2=5.07
r231 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=42.465 //y=5.155 //x2=41.855 //y2=5.155
r232 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.77 //y=5.24 //x2=41.77 //y2=5.155
r233 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=41.77 //y=5.24 //x2=41.77 //y2=5.725
r234 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.975 //y=5.155 //x2=40.89 //y2=5.155
r235 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.685 //y=5.155 //x2=41.77 //y2=5.155
r236 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=41.685 //y=5.155 //x2=40.975 //y2=5.155
r237 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.89 //y=5.24 //x2=40.89 //y2=5.155
r238 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=40.89 //y=5.24 //x2=40.89 //y2=5.725
r239 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.805 //y=5.155 //x2=40.89 //y2=5.155
r240 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=40.805 //y=5.155 //x2=40.095 //y2=5.155
r241 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=40.01 //y=5.24 //x2=40.095 //y2=5.155
r242 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=40.01 //y=5.24 //x2=40.01 //y2=5.725
r243 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=44.4 //y=2.59 //x2=44.4 //y2=2.59
r244 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=42.55 //y=2.59 //x2=42.55 //y2=2.59
r245 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=42.665 //y=2.59 //x2=42.55 //y2=2.59
r246 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=44.285 //y=2.59 //x2=44.4 //y2=2.59
r247 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=44.285 //y=2.59 //x2=42.665 //y2=2.59
ends PM_TMRDFFSNRNQX1\%noxref_10

subckt PM_TMRDFFSNRNQX1\%noxref_11 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 \
 63 64 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 90 92 98 99 100 101 106 \
 107 112 123 125 126 127 )
c281 ( 127 0 ) capacitor c=0.023087f //x=36.815 //y=5.02
c282 ( 126 0 ) capacitor c=0.023519f //x=35.935 //y=5.02
c283 ( 125 0 ) capacitor c=0.0224735f //x=35.055 //y=5.02
c284 ( 123 0 ) capacitor c=0.00853354f //x=37.065 //y=0.915
c285 ( 112 0 ) capacitor c=0.0588394f //x=32.19 //y=4.7
c286 ( 107 0 ) capacitor c=0.0273931f //x=32.19 //y=1.915
c287 ( 106 0 ) capacitor c=0.0456313f //x=32.19 //y=2.08
c288 ( 101 0 ) capacitor c=0.0547611f //x=49.485 //y=4.79
c289 ( 100 0 ) capacitor c=0.0294456f //x=49.775 //y=4.79
c290 ( 99 0 ) capacitor c=0.0347816f //x=49.44 //y=1.22
c291 ( 98 0 ) capacitor c=0.0187487f //x=49.44 //y=0.875
c292 ( 92 0 ) capacitor c=0.0137055f //x=49.285 //y=1.375
c293 ( 90 0 ) capacitor c=0.0149861f //x=49.285 //y=0.72
c294 ( 89 0 ) capacitor c=0.096037f //x=48.91 //y=1.915
c295 ( 88 0 ) capacitor c=0.0228993f //x=48.91 //y=1.53
c296 ( 87 0 ) capacitor c=0.0234352f //x=48.91 //y=1.22
c297 ( 86 0 ) capacitor c=0.0198724f //x=48.91 //y=0.875
c298 ( 85 0 ) capacitor c=0.0432517f //x=32.71 //y=1.26
c299 ( 84 0 ) capacitor c=0.0200379f //x=32.71 //y=0.915
c300 ( 81 0 ) capacitor c=0.0148873f //x=32.555 //y=1.415
c301 ( 79 0 ) capacitor c=0.0157803f //x=32.555 //y=0.76
c302 ( 74 0 ) capacitor c=0.0218028f //x=32.18 //y=1.57
c303 ( 73 0 ) capacitor c=0.0207459f //x=32.18 //y=1.26
c304 ( 72 0 ) capacitor c=0.0194308f //x=32.18 //y=0.915
c305 ( 68 0 ) capacitor c=0.109949f //x=49.85 //y=6.02
c306 ( 67 0 ) capacitor c=0.158483f //x=49.41 //y=6.02
c307 ( 66 0 ) capacitor c=0.158754f //x=32.37 //y=6.02
c308 ( 65 0 ) capacitor c=0.109949f //x=31.93 //y=6.02
c309 ( 62 0 ) capacitor c=9.74268e-19 //x=36.96 //y=5.155
c310 ( 61 0 ) capacitor c=0.00191414f //x=36.08 //y=5.155
c311 ( 54 0 ) capacitor c=0.0938247f //x=49.21 //y=2.08
c312 ( 52 0 ) capacitor c=0.103032f //x=37.74 //y=3.33
c313 ( 48 0 ) capacitor c=0.00398962f //x=37.34 //y=1.665
c314 ( 47 0 ) capacitor c=0.0137288f //x=37.655 //y=1.665
c315 ( 41 0 ) capacitor c=0.0276208f //x=37.655 //y=5.155
c316 ( 33 0 ) capacitor c=0.0169868f //x=36.875 //y=5.155
c317 ( 26 0 ) capacitor c=0.00316998f //x=35.285 //y=5.155
c318 ( 25 0 ) capacitor c=0.014258f //x=35.995 //y=5.155
c319 ( 12 0 ) capacitor c=0.0816952f //x=32.19 //y=2.08
c320 ( 4 0 ) capacitor c=0.00551333f //x=37.855 //y=3.33
c321 ( 3 0 ) capacitor c=0.173188f //x=49.095 //y=3.33
c322 ( 2 0 ) capacitor c=0.0108616f //x=32.305 //y=3.33
c323 ( 1 0 ) capacitor c=0.0905825f //x=37.625 //y=3.33
r324 (  106 107 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=32.19 //y=2.08 //x2=32.19 //y2=1.915
r325 (  100 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=49.775 //y=4.79 //x2=49.85 //y2=4.865
r326 (  100 101 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=49.775 //y=4.79 //x2=49.485 //y2=4.79
r327 (  99 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.44 //y=1.22 //x2=49.4 //y2=1.375
r328 (  98 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.44 //y=0.875 //x2=49.4 //y2=0.72
r329 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=49.44 //y=0.875 //x2=49.44 //y2=1.22
r330 (  95 101 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=49.41 //y=4.865 //x2=49.485 //y2=4.79
r331 (  95 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=49.41 //y=4.865 //x2=49.21 //y2=4.7
r332 (  93 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.065 //y=1.375 //x2=48.95 //y2=1.375
r333 (  92 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.285 //y=1.375 //x2=49.4 //y2=1.375
r334 (  91 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.065 //y=0.72 //x2=48.95 //y2=0.72
r335 (  90 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.285 //y=0.72 //x2=49.4 //y2=0.72
r336 (  90 91 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=49.285 //y=0.72 //x2=49.065 //y2=0.72
r337 (  89 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.915 //x2=49.21 //y2=2.08
r338 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.53 //x2=48.95 //y2=1.375
r339 (  88 89 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.53 //x2=48.91 //y2=1.915
r340 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.22 //x2=48.95 //y2=1.375
r341 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=48.91 //y=0.875 //x2=48.95 //y2=0.72
r342 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=48.91 //y=0.875 //x2=48.91 //y2=1.22
r343 (  85 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.71 //y=1.26 //x2=32.67 //y2=1.415
r344 (  84 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.71 //y=0.915 //x2=32.67 //y2=0.76
r345 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=32.71 //y=0.915 //x2=32.71 //y2=1.26
r346 (  82 110 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.335 //y=1.415 //x2=32.22 //y2=1.415
r347 (  81 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.555 //y=1.415 //x2=32.67 //y2=1.415
r348 (  80 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.335 //y=0.76 //x2=32.22 //y2=0.76
r349 (  79 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.555 //y=0.76 //x2=32.67 //y2=0.76
r350 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=32.555 //y=0.76 //x2=32.335 //y2=0.76
r351 (  76 112 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=32.37 //y=4.865 //x2=32.19 //y2=4.7
r352 (  74 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.18 //y=1.57 //x2=32.22 //y2=1.415
r353 (  74 107 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=32.18 //y=1.57 //x2=32.18 //y2=1.915
r354 (  73 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.18 //y=1.26 //x2=32.22 //y2=1.415
r355 (  72 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.18 //y=0.915 //x2=32.22 //y2=0.76
r356 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=32.18 //y=0.915 //x2=32.18 //y2=1.26
r357 (  69 112 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=31.93 //y=4.865 //x2=32.19 //y2=4.7
r358 (  68 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.85 //y=6.02 //x2=49.85 //y2=4.865
r359 (  67 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.41 //y=6.02 //x2=49.41 //y2=4.865
r360 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=32.37 //y=6.02 //x2=32.37 //y2=4.865
r361 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.93 //y=6.02 //x2=31.93 //y2=4.865
r362 (  64 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=49.175 //y=1.375 //x2=49.285 //y2=1.375
r363 (  64 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=49.175 //y=1.375 //x2=49.065 //y2=1.375
r364 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=32.445 //y=1.415 //x2=32.555 //y2=1.415
r365 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=32.445 //y=1.415 //x2=32.335 //y2=1.415
r366 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.21 //y=4.7 //x2=49.21 //y2=4.7
r367 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=49.21 //y=3.33 //x2=49.21 //y2=4.7
r368 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.21 //y=2.08 //x2=49.21 //y2=2.08
r369 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=49.21 //y=2.08 //x2=49.21 //y2=3.33
r370 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=37.74 //y=5.07 //x2=37.74 //y2=3.33
r371 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=37.74 //y=1.75 //x2=37.74 //y2=3.33
r372 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.655 //y=1.665 //x2=37.74 //y2=1.75
r373 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=37.655 //y=1.665 //x2=37.34 //y2=1.665
r374 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.255 //y=1.58 //x2=37.34 //y2=1.665
r375 (  43 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=37.255 //y=1.58 //x2=37.255 //y2=1.01
r376 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.045 //y=5.155 //x2=36.96 //y2=5.155
r377 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.655 //y=5.155 //x2=37.74 //y2=5.07
r378 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=37.655 //y=5.155 //x2=37.045 //y2=5.155
r379 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.96 //y=5.24 //x2=36.96 //y2=5.155
r380 (  35 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=36.96 //y=5.24 //x2=36.96 //y2=5.725
r381 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.165 //y=5.155 //x2=36.08 //y2=5.155
r382 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.875 //y=5.155 //x2=36.96 //y2=5.155
r383 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=36.875 //y=5.155 //x2=36.165 //y2=5.155
r384 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.08 //y=5.24 //x2=36.08 //y2=5.155
r385 (  27 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=36.08 //y=5.24 //x2=36.08 //y2=5.725
r386 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.995 //y=5.155 //x2=36.08 //y2=5.155
r387 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=35.995 //y=5.155 //x2=35.285 //y2=5.155
r388 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=35.2 //y=5.24 //x2=35.285 //y2=5.155
r389 (  19 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.2 //y=5.24 //x2=35.2 //y2=5.725
r390 (  17 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=32.19 //y=4.7 //x2=32.19 //y2=4.7
r391 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=32.19 //y=3.33 //x2=32.19 //y2=4.7
r392 (  12 106 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=32.19 //y=2.08 //x2=32.19 //y2=2.08
r393 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=32.19 //y=2.08 //x2=32.19 //y2=3.33
r394 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=49.21 //y=3.33 //x2=49.21 //y2=3.33
r395 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=37.74 //y=3.33 //x2=37.74 //y2=3.33
r396 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=32.19 //y=3.33 //x2=32.19 //y2=3.33
r397 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.855 //y=3.33 //x2=37.74 //y2=3.33
r398 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=49.095 //y=3.33 //x2=49.21 //y2=3.33
r399 (  3 4 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=49.095 //y=3.33 //x2=37.855 //y2=3.33
r400 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=32.305 //y=3.33 //x2=32.19 //y2=3.33
r401 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.625 //y=3.33 //x2=37.74 //y2=3.33
r402 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=37.625 //y=3.33 //x2=32.305 //y2=3.33
ends PM_TMRDFFSNRNQX1\%noxref_11

subckt PM_TMRDFFSNRNQX1\%noxref_12 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 \
 53 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c168 ( 85 0 ) capacitor c=0.023087f //x=51.245 //y=5.02
c169 ( 84 0 ) capacitor c=0.023519f //x=50.365 //y=5.02
c170 ( 83 0 ) capacitor c=0.0224735f //x=49.485 //y=5.02
c171 ( 81 0 ) capacitor c=0.00853354f //x=51.495 //y=0.915
c172 ( 69 0 ) capacitor c=0.0547611f //x=54.295 //y=4.79
c173 ( 68 0 ) capacitor c=0.0294456f //x=54.585 //y=4.79
c174 ( 67 0 ) capacitor c=0.0347816f //x=54.25 //y=1.22
c175 ( 66 0 ) capacitor c=0.0187487f //x=54.25 //y=0.875
c176 ( 60 0 ) capacitor c=0.0137055f //x=54.095 //y=1.375
c177 ( 58 0 ) capacitor c=0.0149861f //x=54.095 //y=0.72
c178 ( 57 0 ) capacitor c=0.096037f //x=53.72 //y=1.915
c179 ( 56 0 ) capacitor c=0.0228993f //x=53.72 //y=1.53
c180 ( 55 0 ) capacitor c=0.0234352f //x=53.72 //y=1.22
c181 ( 54 0 ) capacitor c=0.0198724f //x=53.72 //y=0.875
c182 ( 53 0 ) capacitor c=0.109949f //x=54.66 //y=6.02
c183 ( 52 0 ) capacitor c=0.158483f //x=54.22 //y=6.02
c184 ( 50 0 ) capacitor c=9.74268e-19 //x=51.39 //y=5.155
c185 ( 49 0 ) capacitor c=0.00191414f //x=50.51 //y=5.155
c186 ( 42 0 ) capacitor c=0.0910382f //x=54.02 //y=2.08
c187 ( 40 0 ) capacitor c=0.103154f //x=52.17 //y=2.59
c188 ( 36 0 ) capacitor c=0.00398962f //x=51.77 //y=1.665
c189 ( 35 0 ) capacitor c=0.0137288f //x=52.085 //y=1.665
c190 ( 29 0 ) capacitor c=0.0276208f //x=52.085 //y=5.155
c191 ( 21 0 ) capacitor c=0.0169868f //x=51.305 //y=5.155
c192 ( 14 0 ) capacitor c=0.00316998f //x=49.715 //y=5.155
c193 ( 13 0 ) capacitor c=0.014258f //x=50.425 //y=5.155
c194 ( 2 0 ) capacitor c=0.0116088f //x=52.285 //y=2.59
c195 ( 1 0 ) capacitor c=0.0351856f //x=53.905 //y=2.59
r196 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=54.585 //y=4.79 //x2=54.66 //y2=4.865
r197 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=54.585 //y=4.79 //x2=54.295 //y2=4.79
r198 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.25 //y=1.22 //x2=54.21 //y2=1.375
r199 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.25 //y=0.875 //x2=54.21 //y2=0.72
r200 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=54.25 //y=0.875 //x2=54.25 //y2=1.22
r201 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=54.22 //y=4.865 //x2=54.295 //y2=4.79
r202 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=54.22 //y=4.865 //x2=54.02 //y2=4.7
r203 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.875 //y=1.375 //x2=53.76 //y2=1.375
r204 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.095 //y=1.375 //x2=54.21 //y2=1.375
r205 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.875 //y=0.72 //x2=53.76 //y2=0.72
r206 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.095 //y=0.72 //x2=54.21 //y2=0.72
r207 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=54.095 //y=0.72 //x2=53.875 //y2=0.72
r208 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=53.72 //y=1.915 //x2=54.02 //y2=2.08
r209 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.72 //y=1.53 //x2=53.76 //y2=1.375
r210 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=53.72 //y=1.53 //x2=53.72 //y2=1.915
r211 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.72 //y=1.22 //x2=53.76 //y2=1.375
r212 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.72 //y=0.875 //x2=53.76 //y2=0.72
r213 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=53.72 //y=0.875 //x2=53.72 //y2=1.22
r214 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.66 //y=6.02 //x2=54.66 //y2=4.865
r215 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.22 //y=6.02 //x2=54.22 //y2=4.865
r216 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.985 //y=1.375 //x2=54.095 //y2=1.375
r217 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.985 //y=1.375 //x2=53.875 //y2=1.375
r218 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.02 //y=4.7 //x2=54.02 //y2=4.7
r219 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=54.02 //y=2.59 //x2=54.02 //y2=4.7
r220 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.02 //y=2.08 //x2=54.02 //y2=2.08
r221 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=54.02 //y=2.08 //x2=54.02 //y2=2.59
r222 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=52.17 //y=5.07 //x2=52.17 //y2=2.59
r223 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=52.17 //y=1.75 //x2=52.17 //y2=2.59
r224 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=52.085 //y=1.665 //x2=52.17 //y2=1.75
r225 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=52.085 //y=1.665 //x2=51.77 //y2=1.665
r226 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=51.685 //y=1.58 //x2=51.77 //y2=1.665
r227 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=51.685 //y=1.58 //x2=51.685 //y2=1.01
r228 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.475 //y=5.155 //x2=51.39 //y2=5.155
r229 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=52.085 //y=5.155 //x2=52.17 //y2=5.07
r230 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=52.085 //y=5.155 //x2=51.475 //y2=5.155
r231 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.39 //y=5.24 //x2=51.39 //y2=5.155
r232 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=51.39 //y=5.24 //x2=51.39 //y2=5.725
r233 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.595 //y=5.155 //x2=50.51 //y2=5.155
r234 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.305 //y=5.155 //x2=51.39 //y2=5.155
r235 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=51.305 //y=5.155 //x2=50.595 //y2=5.155
r236 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.51 //y=5.24 //x2=50.51 //y2=5.155
r237 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.51 //y=5.24 //x2=50.51 //y2=5.725
r238 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.425 //y=5.155 //x2=50.51 //y2=5.155
r239 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.425 //y=5.155 //x2=49.715 //y2=5.155
r240 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=49.63 //y=5.24 //x2=49.715 //y2=5.155
r241 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=49.63 //y=5.24 //x2=49.63 //y2=5.725
r242 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=54.02 //y=2.59 //x2=54.02 //y2=2.59
r243 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=52.17 //y=2.59 //x2=52.17 //y2=2.59
r244 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=52.285 //y=2.59 //x2=52.17 //y2=2.59
r245 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=53.905 //y=2.59 //x2=54.02 //y2=2.59
r246 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=53.905 //y=2.59 //x2=52.285 //y2=2.59
ends PM_TMRDFFSNRNQX1\%noxref_12

subckt PM_TMRDFFSNRNQX1\%noxref_13 ( 1 2 3 4 5 6 16 24 37 38 45 53 59 60 64 66 \
 73 74 75 76 77 78 79 80 81 82 83 87 88 89 94 96 99 100 104 105 106 111 113 \
 116 117 121 122 123 128 130 133 134 136 137 142 146 147 152 156 157 162 165 \
 167 168 169 )
c347 ( 169 0 ) capacitor c=0.023087f //x=46.435 //y=5.02
c348 ( 168 0 ) capacitor c=0.023519f //x=45.555 //y=5.02
c349 ( 167 0 ) capacitor c=0.0224735f //x=44.675 //y=5.02
c350 ( 165 0 ) capacitor c=0.00853354f //x=46.685 //y=0.915
c351 ( 162 0 ) capacitor c=0.0588394f //x=56.24 //y=4.7
c352 ( 157 0 ) capacitor c=0.0273931f //x=56.24 //y=1.915
c353 ( 156 0 ) capacitor c=0.0456313f //x=56.24 //y=2.08
c354 ( 152 0 ) capacitor c=0.0588394f //x=41.81 //y=4.7
c355 ( 147 0 ) capacitor c=0.0273931f //x=41.81 //y=1.915
c356 ( 146 0 ) capacitor c=0.0456313f //x=41.81 //y=2.08
c357 ( 142 0 ) capacitor c=0.0589949f //x=37 //y=4.7
c358 ( 137 0 ) capacitor c=0.0273931f //x=37 //y=1.915
c359 ( 136 0 ) capacitor c=0.0456313f //x=37 //y=2.08
c360 ( 134 0 ) capacitor c=0.0432517f //x=56.76 //y=1.26
c361 ( 133 0 ) capacitor c=0.0200379f //x=56.76 //y=0.915
c362 ( 130 0 ) capacitor c=0.0148873f //x=56.605 //y=1.415
c363 ( 128 0 ) capacitor c=0.0157803f //x=56.605 //y=0.76
c364 ( 123 0 ) capacitor c=0.0218028f //x=56.23 //y=1.57
c365 ( 122 0 ) capacitor c=0.0207459f //x=56.23 //y=1.26
c366 ( 121 0 ) capacitor c=0.0194308f //x=56.23 //y=0.915
c367 ( 117 0 ) capacitor c=0.0432517f //x=42.33 //y=1.26
c368 ( 116 0 ) capacitor c=0.0200379f //x=42.33 //y=0.915
c369 ( 113 0 ) capacitor c=0.0148873f //x=42.175 //y=1.415
c370 ( 111 0 ) capacitor c=0.0157803f //x=42.175 //y=0.76
c371 ( 106 0 ) capacitor c=0.0218028f //x=41.8 //y=1.57
c372 ( 105 0 ) capacitor c=0.0207459f //x=41.8 //y=1.26
c373 ( 104 0 ) capacitor c=0.0194308f //x=41.8 //y=0.915
c374 ( 100 0 ) capacitor c=0.0432517f //x=37.52 //y=1.26
c375 ( 99 0 ) capacitor c=0.0200379f //x=37.52 //y=0.915
c376 ( 96 0 ) capacitor c=0.0148873f //x=37.365 //y=1.415
c377 ( 94 0 ) capacitor c=0.0157803f //x=37.365 //y=0.76
c378 ( 89 0 ) capacitor c=0.0218028f //x=36.99 //y=1.57
c379 ( 88 0 ) capacitor c=0.0207459f //x=36.99 //y=1.26
c380 ( 87 0 ) capacitor c=0.0194308f //x=36.99 //y=0.915
c381 ( 83 0 ) capacitor c=0.158754f //x=56.42 //y=6.02
c382 ( 82 0 ) capacitor c=0.109949f //x=55.98 //y=6.02
c383 ( 81 0 ) capacitor c=0.158754f //x=41.99 //y=6.02
c384 ( 80 0 ) capacitor c=0.109949f //x=41.55 //y=6.02
c385 ( 79 0 ) capacitor c=0.158754f //x=37.18 //y=6.02
c386 ( 78 0 ) capacitor c=0.109949f //x=36.74 //y=6.02
c387 ( 74 0 ) capacitor c=9.74268e-19 //x=46.58 //y=5.155
c388 ( 73 0 ) capacitor c=0.00191414f //x=45.7 //y=5.155
c389 ( 66 0 ) capacitor c=0.0797834f //x=56.24 //y=2.08
c390 ( 64 0 ) capacitor c=0.104892f //x=47.36 //y=3.7
c391 ( 60 0 ) capacitor c=0.00398962f //x=46.96 //y=1.665
c392 ( 59 0 ) capacitor c=0.0137288f //x=47.275 //y=1.665
c393 ( 53 0 ) capacitor c=0.0276208f //x=47.275 //y=5.155
c394 ( 45 0 ) capacitor c=0.0169868f //x=46.495 //y=5.155
c395 ( 38 0 ) capacitor c=0.00316998f //x=44.905 //y=5.155
c396 ( 37 0 ) capacitor c=0.014258f //x=45.615 //y=5.155
c397 ( 24 0 ) capacitor c=0.0790362f //x=41.81 //y=2.08
c398 ( 16 0 ) capacitor c=0.0776243f //x=37 //y=2.08
c399 ( 6 0 ) capacitor c=0.0055354f //x=47.475 //y=3.7
c400 ( 5 0 ) capacitor c=0.137252f //x=56.125 //y=3.7
c401 ( 4 0 ) capacitor c=0.00533183f //x=41.925 //y=3.7
c402 ( 3 0 ) capacitor c=0.0751185f //x=47.245 //y=3.7
c403 ( 2 0 ) capacitor c=0.01364f //x=37.115 //y=3.7
c404 ( 1 0 ) capacitor c=0.0665749f //x=41.695 //y=3.7
r405 (  156 157 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=56.24 //y=2.08 //x2=56.24 //y2=1.915
r406 (  146 147 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=41.81 //y=2.08 //x2=41.81 //y2=1.915
r407 (  136 137 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=37 //y=2.08 //x2=37 //y2=1.915
r408 (  134 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.76 //y=1.26 //x2=56.72 //y2=1.415
r409 (  133 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.76 //y=0.915 //x2=56.72 //y2=0.76
r410 (  133 134 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.76 //y=0.915 //x2=56.76 //y2=1.26
r411 (  131 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.385 //y=1.415 //x2=56.27 //y2=1.415
r412 (  130 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.605 //y=1.415 //x2=56.72 //y2=1.415
r413 (  129 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.385 //y=0.76 //x2=56.27 //y2=0.76
r414 (  128 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.605 //y=0.76 //x2=56.72 //y2=0.76
r415 (  128 129 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=56.605 //y=0.76 //x2=56.385 //y2=0.76
r416 (  125 162 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=56.42 //y=4.865 //x2=56.24 //y2=4.7
r417 (  123 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.23 //y=1.57 //x2=56.27 //y2=1.415
r418 (  123 157 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.23 //y=1.57 //x2=56.23 //y2=1.915
r419 (  122 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.23 //y=1.26 //x2=56.27 //y2=1.415
r420 (  121 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.23 //y=0.915 //x2=56.27 //y2=0.76
r421 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.23 //y=0.915 //x2=56.23 //y2=1.26
r422 (  118 162 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=55.98 //y=4.865 //x2=56.24 //y2=4.7
r423 (  117 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.33 //y=1.26 //x2=42.29 //y2=1.415
r424 (  116 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.33 //y=0.915 //x2=42.29 //y2=0.76
r425 (  116 117 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.33 //y=0.915 //x2=42.33 //y2=1.26
r426 (  114 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.955 //y=1.415 //x2=41.84 //y2=1.415
r427 (  113 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.175 //y=1.415 //x2=42.29 //y2=1.415
r428 (  112 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.955 //y=0.76 //x2=41.84 //y2=0.76
r429 (  111 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.175 //y=0.76 //x2=42.29 //y2=0.76
r430 (  111 112 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=42.175 //y=0.76 //x2=41.955 //y2=0.76
r431 (  108 152 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=41.99 //y=4.865 //x2=41.81 //y2=4.7
r432 (  106 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.8 //y=1.57 //x2=41.84 //y2=1.415
r433 (  106 147 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=41.8 //y=1.57 //x2=41.8 //y2=1.915
r434 (  105 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.8 //y=1.26 //x2=41.84 //y2=1.415
r435 (  104 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.8 //y=0.915 //x2=41.84 //y2=0.76
r436 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=41.8 //y=0.915 //x2=41.8 //y2=1.26
r437 (  101 152 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=41.55 //y=4.865 //x2=41.81 //y2=4.7
r438 (  100 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.52 //y=1.26 //x2=37.48 //y2=1.415
r439 (  99 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.52 //y=0.915 //x2=37.48 //y2=0.76
r440 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=37.52 //y=0.915 //x2=37.52 //y2=1.26
r441 (  97 140 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.145 //y=1.415 //x2=37.03 //y2=1.415
r442 (  96 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.365 //y=1.415 //x2=37.48 //y2=1.415
r443 (  95 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.145 //y=0.76 //x2=37.03 //y2=0.76
r444 (  94 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.365 //y=0.76 //x2=37.48 //y2=0.76
r445 (  94 95 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=37.365 //y=0.76 //x2=37.145 //y2=0.76
r446 (  91 142 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=37.18 //y=4.865 //x2=37 //y2=4.7
r447 (  89 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.99 //y=1.57 //x2=37.03 //y2=1.415
r448 (  89 137 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=36.99 //y=1.57 //x2=36.99 //y2=1.915
r449 (  88 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.99 //y=1.26 //x2=37.03 //y2=1.415
r450 (  87 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.99 //y=0.915 //x2=37.03 //y2=0.76
r451 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=36.99 //y=0.915 //x2=36.99 //y2=1.26
r452 (  84 142 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=36.74 //y=4.865 //x2=37 //y2=4.7
r453 (  83 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=56.42 //y=6.02 //x2=56.42 //y2=4.865
r454 (  82 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.98 //y=6.02 //x2=55.98 //y2=4.865
r455 (  81 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.99 //y=6.02 //x2=41.99 //y2=4.865
r456 (  80 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.55 //y=6.02 //x2=41.55 //y2=4.865
r457 (  79 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=37.18 //y=6.02 //x2=37.18 //y2=4.865
r458 (  78 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=36.74 //y=6.02 //x2=36.74 //y2=4.865
r459 (  77 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=56.495 //y=1.415 //x2=56.605 //y2=1.415
r460 (  77 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=56.495 //y=1.415 //x2=56.385 //y2=1.415
r461 (  76 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.065 //y=1.415 //x2=42.175 //y2=1.415
r462 (  76 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.065 //y=1.415 //x2=41.955 //y2=1.415
r463 (  75 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.255 //y=1.415 //x2=37.365 //y2=1.415
r464 (  75 97 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.255 //y=1.415 //x2=37.145 //y2=1.415
r465 (  71 162 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=56.24 //y=4.7 //x2=56.24 //y2=4.7
r466 (  69 71 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=56.24 //y=3.7 //x2=56.24 //y2=4.7
r467 (  66 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=56.24 //y=2.08 //x2=56.24 //y2=2.08
r468 (  66 69 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=56.24 //y=2.08 //x2=56.24 //y2=3.7
r469 (  62 64 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=47.36 //y=5.07 //x2=47.36 //y2=3.7
r470 (  61 64 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=47.36 //y=1.75 //x2=47.36 //y2=3.7
r471 (  59 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=47.275 //y=1.665 //x2=47.36 //y2=1.75
r472 (  59 60 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=47.275 //y=1.665 //x2=46.96 //y2=1.665
r473 (  55 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=46.875 //y=1.58 //x2=46.96 //y2=1.665
r474 (  55 165 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=46.875 //y=1.58 //x2=46.875 //y2=1.01
r475 (  54 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.665 //y=5.155 //x2=46.58 //y2=5.155
r476 (  53 62 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=47.275 //y=5.155 //x2=47.36 //y2=5.07
r477 (  53 54 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=47.275 //y=5.155 //x2=46.665 //y2=5.155
r478 (  47 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.58 //y=5.24 //x2=46.58 //y2=5.155
r479 (  47 169 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.58 //y=5.24 //x2=46.58 //y2=5.725
r480 (  46 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.785 //y=5.155 //x2=45.7 //y2=5.155
r481 (  45 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.495 //y=5.155 //x2=46.58 //y2=5.155
r482 (  45 46 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.495 //y=5.155 //x2=45.785 //y2=5.155
r483 (  39 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.7 //y=5.24 //x2=45.7 //y2=5.155
r484 (  39 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.7 //y=5.24 //x2=45.7 //y2=5.725
r485 (  37 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.615 //y=5.155 //x2=45.7 //y2=5.155
r486 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=45.615 //y=5.155 //x2=44.905 //y2=5.155
r487 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=44.82 //y=5.24 //x2=44.905 //y2=5.155
r488 (  31 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=44.82 //y=5.24 //x2=44.82 //y2=5.725
r489 (  29 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.81 //y=4.7 //x2=41.81 //y2=4.7
r490 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=41.81 //y=3.7 //x2=41.81 //y2=4.7
r491 (  24 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.81 //y=2.08 //x2=41.81 //y2=2.08
r492 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=41.81 //y=2.08 //x2=41.81 //y2=3.7
r493 (  21 142 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37 //y=4.7 //x2=37 //y2=4.7
r494 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=37 //y=3.7 //x2=37 //y2=4.7
r495 (  16 136 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37 //y=2.08 //x2=37 //y2=2.08
r496 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=37 //y=2.08 //x2=37 //y2=3.7
r497 (  14 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=56.24 //y=3.7 //x2=56.24 //y2=3.7
r498 (  12 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=47.36 //y=3.7 //x2=47.36 //y2=3.7
r499 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=41.81 //y=3.7 //x2=41.81 //y2=3.7
r500 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=37 \
 //y=3.7 //x2=37 //y2=3.7
r501 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.475 //y=3.7 //x2=47.36 //y2=3.7
r502 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.125 //y=3.7 //x2=56.24 //y2=3.7
r503 (  5 6 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=56.125 //y=3.7 //x2=47.475 //y2=3.7
r504 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=41.925 //y=3.7 //x2=41.81 //y2=3.7
r505 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.245 //y=3.7 //x2=47.36 //y2=3.7
r506 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=47.245 //y=3.7 //x2=41.925 //y2=3.7
r507 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.115 //y=3.7 //x2=37 //y2=3.7
r508 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=41.695 //y=3.7 //x2=41.81 //y2=3.7
r509 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=41.695 //y=3.7 //x2=37.115 //y2=3.7
ends PM_TMRDFFSNRNQX1\%noxref_13

subckt PM_TMRDFFSNRNQX1\%noxref_14 ( 1 2 3 4 6 7 8 9 10 22 35 36 43 51 57 58 \
 62 65 67 73 77 78 82 85 86 87 88 89 90 91 92 93 97 98 99 104 106 109 110 111 \
 112 113 118 120 122 128 129 130 131 132 137 139 141 147 148 150 151 156 160 \
 161 164 172 173 176 184 186 187 188 )
c450 ( 188 0 ) capacitor c=0.023087f //x=56.055 //y=5.02
c451 ( 187 0 ) capacitor c=0.023519f //x=55.175 //y=5.02
c452 ( 186 0 ) capacitor c=0.0224735f //x=54.295 //y=5.02
c453 ( 184 0 ) capacitor c=0.00853354f //x=56.305 //y=0.915
c454 ( 176 0 ) capacitor c=0.0352016f //x=95.11 //y=4.705
c455 ( 173 0 ) capacitor c=0.0279733f //x=95.09 //y=1.915
c456 ( 172 0 ) capacitor c=0.0467621f //x=95.09 //y=2.08
c457 ( 164 0 ) capacitor c=0.03845f //x=88.47 //y=4.705
c458 ( 161 0 ) capacitor c=0.0300885f //x=88.43 //y=1.915
c459 ( 160 0 ) capacitor c=0.0504818f //x=88.43 //y=2.08
c460 ( 156 0 ) capacitor c=0.0588394f //x=51.43 //y=4.7
c461 ( 151 0 ) capacitor c=0.0273931f //x=51.43 //y=1.915
c462 ( 150 0 ) capacitor c=0.0456313f //x=51.43 //y=2.08
c463 ( 148 0 ) capacitor c=0.0237734f //x=95.655 //y=1.255
c464 ( 147 0 ) capacitor c=0.0191782f //x=95.655 //y=0.905
c465 ( 141 0 ) capacitor c=0.0351663f //x=95.5 //y=1.405
c466 ( 139 0 ) capacitor c=0.0157803f //x=95.5 //y=0.75
c467 ( 137 0 ) capacitor c=0.0374703f //x=95.495 //y=4.795
c468 ( 132 0 ) capacitor c=0.0200628f //x=95.125 //y=1.56
c469 ( 131 0 ) capacitor c=0.0168575f //x=95.125 //y=1.255
c470 ( 130 0 ) capacitor c=0.0174993f //x=95.125 //y=0.905
c471 ( 129 0 ) capacitor c=0.0435065f //x=88.995 //y=1.25
c472 ( 128 0 ) capacitor c=0.019286f //x=88.995 //y=0.905
c473 ( 122 0 ) capacitor c=0.0164316f //x=88.84 //y=1.405
c474 ( 120 0 ) capacitor c=0.0157795f //x=88.84 //y=0.75
c475 ( 118 0 ) capacitor c=0.029531f //x=88.835 //y=4.795
c476 ( 113 0 ) capacitor c=0.0206178f //x=88.465 //y=1.56
c477 ( 112 0 ) capacitor c=0.016848f //x=88.465 //y=1.25
c478 ( 111 0 ) capacitor c=0.0174777f //x=88.465 //y=0.905
c479 ( 110 0 ) capacitor c=0.0432517f //x=51.95 //y=1.26
c480 ( 109 0 ) capacitor c=0.0200379f //x=51.95 //y=0.915
c481 ( 106 0 ) capacitor c=0.0148873f //x=51.795 //y=1.415
c482 ( 104 0 ) capacitor c=0.0157803f //x=51.795 //y=0.76
c483 ( 99 0 ) capacitor c=0.0218028f //x=51.42 //y=1.57
c484 ( 98 0 ) capacitor c=0.0207459f //x=51.42 //y=1.26
c485 ( 97 0 ) capacitor c=0.0194308f //x=51.42 //y=0.915
c486 ( 93 0 ) capacitor c=0.15325f //x=95.57 //y=6.025
c487 ( 92 0 ) capacitor c=0.110411f //x=95.13 //y=6.025
c488 ( 91 0 ) capacitor c=0.154236f //x=88.91 //y=6.025
c489 ( 90 0 ) capacitor c=0.110294f //x=88.47 //y=6.025
c490 ( 89 0 ) capacitor c=0.158754f //x=51.61 //y=6.02
c491 ( 88 0 ) capacitor c=0.109949f //x=51.17 //y=6.02
c492 ( 82 0 ) capacitor c=0.00501304f //x=95.11 //y=4.705
c493 ( 78 0 ) capacitor c=9.74268e-19 //x=56.2 //y=5.155
c494 ( 77 0 ) capacitor c=0.00191414f //x=55.32 //y=5.155
c495 ( 73 0 ) capacitor c=0.0903046f //x=95.09 //y=2.08
c496 ( 67 0 ) capacitor c=0.110253f //x=88.43 //y=2.08
c497 ( 65 0 ) capacitor c=0.00669947f //x=88.43 //y=4.54
c498 ( 62 0 ) capacitor c=0.104652f //x=56.98 //y=3.33
c499 ( 58 0 ) capacitor c=0.00398962f //x=56.58 //y=1.665
c500 ( 57 0 ) capacitor c=0.0137288f //x=56.895 //y=1.665
c501 ( 51 0 ) capacitor c=0.0276208f //x=56.895 //y=5.155
c502 ( 43 0 ) capacitor c=0.0169868f //x=56.115 //y=5.155
c503 ( 36 0 ) capacitor c=0.00316998f //x=54.525 //y=5.155
c504 ( 35 0 ) capacitor c=0.014258f //x=55.235 //y=5.155
c505 ( 22 0 ) capacitor c=0.0799652f //x=51.43 //y=2.08
c506 ( 10 0 ) capacitor c=0.00672327f //x=88.545 //y=4.07
c507 ( 9 0 ) capacitor c=0.213063f //x=94.975 //y=4.07
c508 ( 8 0 ) capacitor c=0.004561f //x=65.205 //y=4.07
c509 ( 7 0 ) capacitor c=0.347024f //x=88.315 //y=4.07
c510 ( 6 0 ) capacitor c=0.00784097f //x=65.12 //y=3.985
c511 ( 4 0 ) capacitor c=0.00594726f //x=57.095 //y=3.7
c512 ( 3 0 ) capacitor c=0.14546f //x=65.035 //y=3.7
c513 ( 2 0 ) capacitor c=0.00889972f //x=51.545 //y=3.33
c514 ( 1 0 ) capacitor c=0.0876378f //x=56.865 //y=3.33
r515 (  178 179 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=95.11 //y=4.795 //x2=95.11 //y2=4.87
r516 (  176 178 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=95.11 //y=4.705 //x2=95.11 //y2=4.795
r517 (  172 173 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=95.09 //y=2.08 //x2=95.09 //y2=1.915
r518 (  164 166 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=88.47 //y=4.705 //x2=88.47 //y2=4.795
r519 (  160 161 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=88.43 //y=2.08 //x2=88.43 //y2=1.915
r520 (  150 151 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=51.43 //y=2.08 //x2=51.43 //y2=1.915
r521 (  148 183 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=95.655 //y=1.255 //x2=95.655 //y2=1.367
r522 (  147 182 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=95.655 //y=0.905 //x2=95.615 //y2=0.75
r523 (  147 148 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=95.655 //y=0.905 //x2=95.655 //y2=1.255
r524 (  142 181 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=95.28 //y=1.405 //x2=95.165 //y2=1.405
r525 (  141 183 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=95.5 //y=1.405 //x2=95.655 //y2=1.367
r526 (  140 180 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=95.28 //y=0.75 //x2=95.165 //y2=0.75
r527 (  139 182 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=95.5 //y=0.75 //x2=95.615 //y2=0.75
r528 (  139 140 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=95.5 //y=0.75 //x2=95.28 //y2=0.75
r529 (  138 178 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=95.245 //y=4.795 //x2=95.11 //y2=4.795
r530 (  137 144 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=95.495 //y=4.795 //x2=95.57 //y2=4.87
r531 (  137 138 ) resistor r=128.191 //w=0.094 //l=0.25 //layer=ply \
 //thickness=0.18 //x=95.495 //y=4.795 //x2=95.245 //y2=4.795
r532 (  132 181 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=95.125 //y=1.56 //x2=95.165 //y2=1.405
r533 (  132 173 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=95.125 //y=1.56 //x2=95.125 //y2=1.915
r534 (  131 181 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=95.125 //y=1.255 //x2=95.165 //y2=1.405
r535 (  130 180 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=95.125 //y=0.905 //x2=95.165 //y2=0.75
r536 (  130 131 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=95.125 //y=0.905 //x2=95.125 //y2=1.255
r537 (  129 170 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.995 //y=1.25 //x2=88.955 //y2=1.405
r538 (  128 169 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.995 //y=0.905 //x2=88.955 //y2=0.75
r539 (  128 129 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=88.995 //y=0.905 //x2=88.995 //y2=1.25
r540 (  123 168 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=88.62 //y=1.405 //x2=88.505 //y2=1.405
r541 (  122 170 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=88.84 //y=1.405 //x2=88.955 //y2=1.405
r542 (  121 167 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=88.62 //y=0.75 //x2=88.505 //y2=0.75
r543 (  120 169 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=88.84 //y=0.75 //x2=88.955 //y2=0.75
r544 (  120 121 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=88.84 //y=0.75 //x2=88.62 //y2=0.75
r545 (  119 166 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=88.605 //y=4.795 //x2=88.47 //y2=4.795
r546 (  118 125 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=88.835 //y=4.795 //x2=88.91 //y2=4.87
r547 (  118 119 ) resistor r=117.936 //w=0.094 //l=0.23 //layer=ply \
 //thickness=0.18 //x=88.835 //y=4.795 //x2=88.605 //y2=4.795
r548 (  115 166 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=88.47 //y=4.87 //x2=88.47 //y2=4.795
r549 (  113 168 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.465 //y=1.56 //x2=88.505 //y2=1.405
r550 (  113 161 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=88.465 //y=1.56 //x2=88.465 //y2=1.915
r551 (  112 168 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.465 //y=1.25 //x2=88.505 //y2=1.405
r552 (  111 167 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=88.465 //y=0.905 //x2=88.505 //y2=0.75
r553 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=88.465 //y=0.905 //x2=88.465 //y2=1.25
r554 (  110 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.95 //y=1.26 //x2=51.91 //y2=1.415
r555 (  109 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.95 //y=0.915 //x2=51.91 //y2=0.76
r556 (  109 110 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=51.95 //y=0.915 //x2=51.95 //y2=1.26
r557 (  107 154 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.575 //y=1.415 //x2=51.46 //y2=1.415
r558 (  106 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.795 //y=1.415 //x2=51.91 //y2=1.415
r559 (  105 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.575 //y=0.76 //x2=51.46 //y2=0.76
r560 (  104 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.795 //y=0.76 //x2=51.91 //y2=0.76
r561 (  104 105 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=51.795 //y=0.76 //x2=51.575 //y2=0.76
r562 (  101 156 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=51.61 //y=4.865 //x2=51.43 //y2=4.7
r563 (  99 154 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.42 //y=1.57 //x2=51.46 //y2=1.415
r564 (  99 151 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=51.42 //y=1.57 //x2=51.42 //y2=1.915
r565 (  98 154 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.42 //y=1.26 //x2=51.46 //y2=1.415
r566 (  97 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.42 //y=0.915 //x2=51.46 //y2=0.76
r567 (  97 98 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=51.42 //y=0.915 //x2=51.42 //y2=1.26
r568 (  94 156 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=51.17 //y=4.865 //x2=51.43 //y2=4.7
r569 (  93 144 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=95.57 //y=6.025 //x2=95.57 //y2=4.87
r570 (  92 179 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=95.13 //y=6.025 //x2=95.13 //y2=4.87
r571 (  91 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=88.91 //y=6.025 //x2=88.91 //y2=4.87
r572 (  90 115 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=88.47 //y=6.025 //x2=88.47 //y2=4.87
r573 (  89 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=51.61 //y=6.02 //x2=51.61 //y2=4.865
r574 (  88 94 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=51.17 //y=6.02 //x2=51.17 //y2=4.865
r575 (  87 141 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=95.39 //y=1.405 //x2=95.5 //y2=1.405
r576 (  87 142 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=95.39 //y=1.405 //x2=95.28 //y2=1.405
r577 (  86 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=88.73 //y=1.405 //x2=88.84 //y2=1.405
r578 (  86 123 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=88.73 //y=1.405 //x2=88.62 //y2=1.405
r579 (  85 106 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=51.685 //y=1.415 //x2=51.795 //y2=1.415
r580 (  85 107 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=51.685 //y=1.415 //x2=51.575 //y2=1.415
r581 (  82 176 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=95.11 //y=4.705 //x2=95.11 //y2=4.705
r582 (  82 83 ) resistor r=10.3507 //w=0.207 //l=0.165 //layer=li \
 //thickness=0.1 //x=95.1 //y=4.705 //x2=95.1 //y2=4.54
r583 (  80 164 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=88.47 //y=4.705 //x2=88.47 //y2=4.705
r584 (  76 83 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=95.09 //y=4.07 //x2=95.09 //y2=4.54
r585 (  73 172 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=95.09 //y=2.08 //x2=95.09 //y2=2.08
r586 (  73 76 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=95.09 //y=2.08 //x2=95.09 //y2=4.07
r587 (  67 160 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=88.43 //y=2.08 //x2=88.43 //y2=2.08
r588 (  67 70 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=88.43 //y=2.08 //x2=88.43 //y2=4.07
r589 (  65 80 ) resistor r=11.2426 //w=0.191 //l=0.174714 //layer=li \
 //thickness=0.1 //x=88.43 //y=4.54 //x2=88.45 //y2=4.705
r590 (  65 70 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=88.43 //y=4.54 //x2=88.43 //y2=4.07
r591 (  62 64 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=56.98 //y=3.33 //x2=56.98 //y2=3.7
r592 (  60 64 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=56.98 //y=5.07 //x2=56.98 //y2=3.7
r593 (  59 62 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=56.98 //y=1.75 //x2=56.98 //y2=3.33
r594 (  57 59 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.895 //y=1.665 //x2=56.98 //y2=1.75
r595 (  57 58 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=56.895 //y=1.665 //x2=56.58 //y2=1.665
r596 (  53 58 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.495 //y=1.58 //x2=56.58 //y2=1.665
r597 (  53 184 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=56.495 //y=1.58 //x2=56.495 //y2=1.01
r598 (  52 78 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.285 //y=5.155 //x2=56.2 //y2=5.155
r599 (  51 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.895 //y=5.155 //x2=56.98 //y2=5.07
r600 (  51 52 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=56.895 //y=5.155 //x2=56.285 //y2=5.155
r601 (  45 78 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.2 //y=5.24 //x2=56.2 //y2=5.155
r602 (  45 188 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=56.2 //y=5.24 //x2=56.2 //y2=5.725
r603 (  44 77 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.405 //y=5.155 //x2=55.32 //y2=5.155
r604 (  43 78 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.115 //y=5.155 //x2=56.2 //y2=5.155
r605 (  43 44 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=56.115 //y=5.155 //x2=55.405 //y2=5.155
r606 (  37 77 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.32 //y=5.24 //x2=55.32 //y2=5.155
r607 (  37 187 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.32 //y=5.24 //x2=55.32 //y2=5.725
r608 (  35 77 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.235 //y=5.155 //x2=55.32 //y2=5.155
r609 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=55.235 //y=5.155 //x2=54.525 //y2=5.155
r610 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=54.44 //y=5.24 //x2=54.525 //y2=5.155
r611 (  29 186 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.44 //y=5.24 //x2=54.44 //y2=5.725
r612 (  27 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=51.43 //y=4.7 //x2=51.43 //y2=4.7
r613 (  25 27 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=51.43 //y=3.33 //x2=51.43 //y2=4.7
r614 (  22 150 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=51.43 //y=2.08 //x2=51.43 //y2=2.08
r615 (  22 25 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=51.43 //y=2.08 //x2=51.43 //y2=3.33
r616 (  20 76 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=95.09 //y=4.07 //x2=95.09 //y2=4.07
r617 (  18 70 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=88.43 //y=4.07 //x2=88.43 //y2=4.07
r618 (  16 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=56.98 //y=3.33 //x2=56.98 //y2=3.33
r619 (  14 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=56.98 //y=3.7 //x2=56.98 //y2=3.7
r620 (  12 25 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=51.43 //y=3.33 //x2=51.43 //y2=3.33
r621 (  10 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=88.545 //y=4.07 //x2=88.43 //y2=4.07
r622 (  9 20 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=94.975 //y=4.07 //x2=95.09 //y2=4.07
r623 (  9 10 ) resistor r=6.1355 //w=0.131 //l=6.43 //layer=m1 \
 //thickness=0.36 //x=94.975 //y=4.07 //x2=88.545 //y2=4.07
r624 (  7 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=88.315 //y=4.07 //x2=88.43 //y2=4.07
r625 (  7 8 ) resistor r=22.0515 //w=0.131 //l=23.11 //layer=m1 \
 //thickness=0.36 //x=88.315 //y=4.07 //x2=65.205 //y2=4.07
r626 (  6 8 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=65.12 //y=3.985 //x2=65.205 //y2=4.07
r627 (  5 6 ) resistor r=0.19084 //w=0.131 //l=0.2 //layer=m1 //thickness=0.36 \
 //x=65.12 //y=3.785 //x2=65.12 //y2=3.985
r628 (  4 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=57.095 //y=3.7 //x2=56.98 //y2=3.7
r629 (  3 5 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=65.035 //y=3.7 //x2=65.12 //y2=3.785
r630 (  3 4 ) resistor r=7.57634 //w=0.131 //l=7.94 //layer=m1 \
 //thickness=0.36 //x=65.035 //y=3.7 //x2=57.095 //y2=3.7
r631 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=51.545 //y=3.33 //x2=51.43 //y2=3.33
r632 (  1 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.865 //y=3.33 //x2=56.98 //y2=3.33
r633 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=56.865 //y=3.33 //x2=51.545 //y2=3.33
ends PM_TMRDFFSNRNQX1\%noxref_14

subckt PM_TMRDFFSNRNQX1\%D ( 1 2 3 4 11 12 13 14 15 16 17 18 19 20 21 22 23 24 \
 26 40 51 60 61 62 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 \
 92 94 100 101 102 103 107 108 109 110 111 113 119 120 121 122 )
c341 ( 122 0 ) capacitor c=0.0547611f //x=59.105 //y=4.79
c342 ( 121 0 ) capacitor c=0.0294456f //x=59.395 //y=4.79
c343 ( 120 0 ) capacitor c=0.0347816f //x=59.06 //y=1.22
c344 ( 119 0 ) capacitor c=0.0187487f //x=59.06 //y=0.875
c345 ( 113 0 ) capacitor c=0.0137055f //x=58.905 //y=1.375
c346 ( 111 0 ) capacitor c=0.0149861f //x=58.905 //y=0.72
c347 ( 110 0 ) capacitor c=0.096037f //x=58.53 //y=1.915
c348 ( 109 0 ) capacitor c=0.0228993f //x=58.53 //y=1.53
c349 ( 108 0 ) capacitor c=0.0234352f //x=58.53 //y=1.22
c350 ( 107 0 ) capacitor c=0.0198724f //x=58.53 //y=0.875
c351 ( 103 0 ) capacitor c=0.0547611f //x=30.245 //y=4.79
c352 ( 102 0 ) capacitor c=0.0294456f //x=30.535 //y=4.79
c353 ( 101 0 ) capacitor c=0.0347816f //x=30.2 //y=1.22
c354 ( 100 0 ) capacitor c=0.0187487f //x=30.2 //y=0.875
c355 ( 94 0 ) capacitor c=0.0137055f //x=30.045 //y=1.375
c356 ( 92 0 ) capacitor c=0.0149861f //x=30.045 //y=0.72
c357 ( 91 0 ) capacitor c=0.096037f //x=29.67 //y=1.915
c358 ( 90 0 ) capacitor c=0.0228993f //x=29.67 //y=1.53
c359 ( 89 0 ) capacitor c=0.0234352f //x=29.67 //y=1.22
c360 ( 88 0 ) capacitor c=0.0198724f //x=29.67 //y=0.875
c361 ( 84 0 ) capacitor c=0.0558341f //x=1.385 //y=4.79
c362 ( 83 0 ) capacitor c=0.0298189f //x=1.675 //y=4.79
c363 ( 82 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c364 ( 81 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c365 ( 75 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c366 ( 73 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c367 ( 72 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c368 ( 71 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c369 ( 70 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c370 ( 69 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c371 ( 68 0 ) capacitor c=0.109949f //x=59.47 //y=6.02
c372 ( 67 0 ) capacitor c=0.158483f //x=59.03 //y=6.02
c373 ( 66 0 ) capacitor c=0.109949f //x=30.61 //y=6.02
c374 ( 65 0 ) capacitor c=0.158483f //x=30.17 //y=6.02
c375 ( 64 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c376 ( 63 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c377 ( 51 0 ) capacitor c=0.0959046f //x=58.83 //y=2.08
c378 ( 40 0 ) capacitor c=0.0991769f //x=29.97 //y=2.08
c379 ( 26 0 ) capacitor c=0.124371f //x=1.11 //y=2.08
c380 ( 4 0 ) capacitor c=0.00590384f //x=30.085 //y=4.07
c381 ( 3 0 ) capacitor c=0.426259f //x=58.715 //y=4.07
c382 ( 2 0 ) capacitor c=0.0231516f //x=1.225 //y=4.07
c383 ( 1 0 ) capacitor c=0.512603f //x=29.855 //y=4.07
r384 (  121 123 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=59.395 //y=4.79 //x2=59.47 //y2=4.865
r385 (  121 122 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=59.395 //y=4.79 //x2=59.105 //y2=4.79
r386 (  120 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.06 //y=1.22 //x2=59.02 //y2=1.375
r387 (  119 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.06 //y=0.875 //x2=59.02 //y2=0.72
r388 (  119 120 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=59.06 //y=0.875 //x2=59.06 //y2=1.22
r389 (  116 122 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=59.03 //y=4.865 //x2=59.105 //y2=4.79
r390 (  116 147 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=59.03 //y=4.865 //x2=58.83 //y2=4.7
r391 (  114 143 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.685 //y=1.375 //x2=58.57 //y2=1.375
r392 (  113 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.905 //y=1.375 //x2=59.02 //y2=1.375
r393 (  112 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.685 //y=0.72 //x2=58.57 //y2=0.72
r394 (  111 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.905 //y=0.72 //x2=59.02 //y2=0.72
r395 (  111 112 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=58.905 //y=0.72 //x2=58.685 //y2=0.72
r396 (  110 145 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=58.53 //y=1.915 //x2=58.83 //y2=2.08
r397 (  109 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.53 //y=1.53 //x2=58.57 //y2=1.375
r398 (  109 110 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=58.53 //y=1.53 //x2=58.53 //y2=1.915
r399 (  108 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.53 //y=1.22 //x2=58.57 //y2=1.375
r400 (  107 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.53 //y=0.875 //x2=58.57 //y2=0.72
r401 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=58.53 //y=0.875 //x2=58.53 //y2=1.22
r402 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=30.535 //y=4.79 //x2=30.61 //y2=4.865
r403 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=30.535 //y=4.79 //x2=30.245 //y2=4.79
r404 (  101 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.2 //y=1.22 //x2=30.16 //y2=1.375
r405 (  100 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.2 //y=0.875 //x2=30.16 //y2=0.72
r406 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=30.2 //y=0.875 //x2=30.2 //y2=1.22
r407 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=30.17 //y=4.865 //x2=30.245 //y2=4.79
r408 (  97 139 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=30.17 //y=4.865 //x2=29.97 //y2=4.7
r409 (  95 135 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.825 //y=1.375 //x2=29.71 //y2=1.375
r410 (  94 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.045 //y=1.375 //x2=30.16 //y2=1.375
r411 (  93 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.825 //y=0.72 //x2=29.71 //y2=0.72
r412 (  92 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.045 //y=0.72 //x2=30.16 //y2=0.72
r413 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=30.045 //y=0.72 //x2=29.825 //y2=0.72
r414 (  91 137 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=29.67 //y=1.915 //x2=29.97 //y2=2.08
r415 (  90 135 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.67 //y=1.53 //x2=29.71 //y2=1.375
r416 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=29.67 //y=1.53 //x2=29.67 //y2=1.915
r417 (  89 135 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.67 //y=1.22 //x2=29.71 //y2=1.375
r418 (  88 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.67 //y=0.875 //x2=29.71 //y2=0.72
r419 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=29.67 //y=0.875 //x2=29.67 //y2=1.22
r420 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r421 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r422 (  82 133 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r423 (  81 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r424 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r425 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r426 (  78 131 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r427 (  76 127 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r428 (  75 133 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r429 (  74 126 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r430 (  73 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r431 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r432 (  72 129 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r433 (  71 127 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r434 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r435 (  70 127 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r436 (  69 126 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r437 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r438 (  68 123 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.47 //y=6.02 //x2=59.47 //y2=4.865
r439 (  67 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.03 //y=6.02 //x2=59.03 //y2=4.865
r440 (  66 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.61 //y=6.02 //x2=30.61 //y2=4.865
r441 (  65 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.17 //y=6.02 //x2=30.17 //y2=4.865
r442 (  64 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r443 (  63 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r444 (  62 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.795 //y=1.375 //x2=58.905 //y2=1.375
r445 (  62 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.795 //y=1.375 //x2=58.685 //y2=1.375
r446 (  61 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=29.935 //y=1.375 //x2=30.045 //y2=1.375
r447 (  61 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=29.935 //y=1.375 //x2=29.825 //y2=1.375
r448 (  60 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r449 (  60 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r450 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.83 //y=4.7 //x2=58.83 //y2=4.7
r451 (  51 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.83 //y=2.08 //x2=58.83 //y2=2.08
r452 (  48 139 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.97 //y=4.7 //x2=29.97 //y2=4.7
r453 (  40 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.97 //y=2.08 //x2=29.97 //y2=2.08
r454 (  37 131 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r455 (  26 129 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r456 (  24 58 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=58.83 //y=4.07 //x2=58.83 //y2=4.7
r457 (  23 24 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=58.83 //y=3.33 //x2=58.83 //y2=4.07
r458 (  22 23 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=58.83 //y=2.59 //x2=58.83 //y2=3.33
r459 (  22 51 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=58.83 //y=2.59 //x2=58.83 //y2=2.08
r460 (  21 48 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=29.97 //y=4.07 //x2=29.97 //y2=4.7
r461 (  20 21 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=29.97 //y=3.7 //x2=29.97 //y2=4.07
r462 (  19 20 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=29.97 //y=3.33 //x2=29.97 //y2=3.7
r463 (  18 19 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=29.97 //y=2.59 //x2=29.97 //y2=3.33
r464 (  18 40 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=29.97 //y=2.59 //x2=29.97 //y2=2.08
r465 (  17 37 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.44 //x2=1.11 //y2=4.7
r466 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r467 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r468 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r469 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r470 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r471 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.22 //x2=1.11 //y2=2.59
r472 (  11 26 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.22 //x2=1.11 //y2=2.08
r473 (  10 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=58.83 //y=4.07 //x2=58.83 //y2=4.07
r474 (  8 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=29.97 //y=4.07 //x2=29.97 //y2=4.07
r475 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.07
r476 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=30.085 //y=4.07 //x2=29.97 //y2=4.07
r477 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=58.715 //y=4.07 //x2=58.83 //y2=4.07
r478 (  3 4 ) resistor r=27.3187 //w=0.131 //l=28.63 //layer=m1 \
 //thickness=0.36 //x=58.715 //y=4.07 //x2=30.085 //y2=4.07
r479 (  2 6 ) resistor r=0.0738079 //w=0.207 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=4.07 //x2=1.11 //y2=4.07
r480 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=29.855 //y=4.07 //x2=29.97 //y2=4.07
r481 (  1 2 ) resistor r=27.3187 //w=0.131 //l=28.63 //layer=m1 \
 //thickness=0.36 //x=29.855 //y=4.07 //x2=1.225 //y2=4.07
ends PM_TMRDFFSNRNQX1\%D

subckt PM_TMRDFFSNRNQX1\%noxref_16 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 \
 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c253 ( 127 0 ) capacitor c=0.023087f //x=60.865 //y=5.02
c254 ( 126 0 ) capacitor c=0.023519f //x=59.985 //y=5.02
c255 ( 125 0 ) capacitor c=0.0224735f //x=59.105 //y=5.02
c256 ( 123 0 ) capacitor c=0.00853354f //x=61.115 //y=0.915
c257 ( 103 0 ) capacitor c=0.0547611f //x=68.725 //y=4.79
c258 ( 102 0 ) capacitor c=0.0294456f //x=69.015 //y=4.79
c259 ( 101 0 ) capacitor c=0.0347816f //x=68.68 //y=1.22
c260 ( 100 0 ) capacitor c=0.0187487f //x=68.68 //y=0.875
c261 ( 94 0 ) capacitor c=0.0137055f //x=68.525 //y=1.375
c262 ( 92 0 ) capacitor c=0.0149861f //x=68.525 //y=0.72
c263 ( 91 0 ) capacitor c=0.096037f //x=68.15 //y=1.915
c264 ( 90 0 ) capacitor c=0.0228993f //x=68.15 //y=1.53
c265 ( 89 0 ) capacitor c=0.0234352f //x=68.15 //y=1.22
c266 ( 88 0 ) capacitor c=0.0198724f //x=68.15 //y=0.875
c267 ( 84 0 ) capacitor c=0.0549166f //x=63.915 //y=4.79
c268 ( 83 0 ) capacitor c=0.0294456f //x=64.205 //y=4.79
c269 ( 82 0 ) capacitor c=0.0347816f //x=63.87 //y=1.22
c270 ( 81 0 ) capacitor c=0.0187487f //x=63.87 //y=0.875
c271 ( 75 0 ) capacitor c=0.0137055f //x=63.715 //y=1.375
c272 ( 73 0 ) capacitor c=0.0149861f //x=63.715 //y=0.72
c273 ( 72 0 ) capacitor c=0.096037f //x=63.34 //y=1.915
c274 ( 71 0 ) capacitor c=0.0228993f //x=63.34 //y=1.53
c275 ( 70 0 ) capacitor c=0.0234352f //x=63.34 //y=1.22
c276 ( 69 0 ) capacitor c=0.0198724f //x=63.34 //y=0.875
c277 ( 68 0 ) capacitor c=0.109949f //x=69.09 //y=6.02
c278 ( 67 0 ) capacitor c=0.158483f //x=68.65 //y=6.02
c279 ( 66 0 ) capacitor c=0.109949f //x=64.28 //y=6.02
c280 ( 65 0 ) capacitor c=0.158483f //x=63.84 //y=6.02
c281 ( 62 0 ) capacitor c=9.74268e-19 //x=61.01 //y=5.155
c282 ( 61 0 ) capacitor c=0.00191414f //x=60.13 //y=5.155
c283 ( 54 0 ) capacitor c=0.0913827f //x=68.45 //y=2.08
c284 ( 46 0 ) capacitor c=0.093372f //x=63.64 //y=2.08
c285 ( 44 0 ) capacitor c=0.105725f //x=61.79 //y=2.59
c286 ( 40 0 ) capacitor c=0.00398962f //x=61.39 //y=1.665
c287 ( 39 0 ) capacitor c=0.0137288f //x=61.705 //y=1.665
c288 ( 33 0 ) capacitor c=0.0276208f //x=61.705 //y=5.155
c289 ( 25 0 ) capacitor c=0.0169868f //x=60.925 //y=5.155
c290 ( 18 0 ) capacitor c=0.00316998f //x=59.335 //y=5.155
c291 ( 17 0 ) capacitor c=0.014258f //x=60.045 //y=5.155
c292 ( 4 0 ) capacitor c=0.00401138f //x=63.755 //y=2.59
c293 ( 3 0 ) capacitor c=0.0706637f //x=68.335 //y=2.59
c294 ( 2 0 ) capacitor c=0.0120752f //x=61.905 //y=2.59
c295 ( 1 0 ) capacitor c=0.0233554f //x=63.525 //y=2.59
r296 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=69.015 //y=4.79 //x2=69.09 //y2=4.865
r297 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=69.015 //y=4.79 //x2=68.725 //y2=4.79
r298 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.68 //y=1.22 //x2=68.64 //y2=1.375
r299 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.68 //y=0.875 //x2=68.64 //y2=0.72
r300 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=68.68 //y=0.875 //x2=68.68 //y2=1.22
r301 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=68.65 //y=4.865 //x2=68.725 //y2=4.79
r302 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=68.65 //y=4.865 //x2=68.45 //y2=4.7
r303 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.305 //y=1.375 //x2=68.19 //y2=1.375
r304 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.525 //y=1.375 //x2=68.64 //y2=1.375
r305 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.305 //y=0.72 //x2=68.19 //y2=0.72
r306 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.525 //y=0.72 //x2=68.64 //y2=0.72
r307 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=68.525 //y=0.72 //x2=68.305 //y2=0.72
r308 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=68.15 //y=1.915 //x2=68.45 //y2=2.08
r309 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.15 //y=1.53 //x2=68.19 //y2=1.375
r310 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=68.15 //y=1.53 //x2=68.15 //y2=1.915
r311 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.15 //y=1.22 //x2=68.19 //y2=1.375
r312 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.15 //y=0.875 //x2=68.19 //y2=0.72
r313 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=68.15 //y=0.875 //x2=68.15 //y2=1.22
r314 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=64.205 //y=4.79 //x2=64.28 //y2=4.865
r315 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=64.205 //y=4.79 //x2=63.915 //y2=4.79
r316 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.87 //y=1.22 //x2=63.83 //y2=1.375
r317 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.87 //y=0.875 //x2=63.83 //y2=0.72
r318 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.87 //y=0.875 //x2=63.87 //y2=1.22
r319 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=63.84 //y=4.865 //x2=63.915 //y2=4.79
r320 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=63.84 //y=4.865 //x2=63.64 //y2=4.7
r321 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.495 //y=1.375 //x2=63.38 //y2=1.375
r322 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.715 //y=1.375 //x2=63.83 //y2=1.375
r323 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.495 //y=0.72 //x2=63.38 //y2=0.72
r324 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.715 //y=0.72 //x2=63.83 //y2=0.72
r325 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=63.715 //y=0.72 //x2=63.495 //y2=0.72
r326 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=63.34 //y=1.915 //x2=63.64 //y2=2.08
r327 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.34 //y=1.53 //x2=63.38 //y2=1.375
r328 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=63.34 //y=1.53 //x2=63.34 //y2=1.915
r329 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.34 //y=1.22 //x2=63.38 //y2=1.375
r330 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.34 //y=0.875 //x2=63.38 //y2=0.72
r331 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.34 //y=0.875 //x2=63.34 //y2=1.22
r332 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.09 //y=6.02 //x2=69.09 //y2=4.865
r333 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=68.65 //y=6.02 //x2=68.65 //y2=4.865
r334 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=64.28 //y=6.02 //x2=64.28 //y2=4.865
r335 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=63.84 //y=6.02 //x2=63.84 //y2=4.865
r336 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=68.415 //y=1.375 //x2=68.525 //y2=1.375
r337 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=68.415 //y=1.375 //x2=68.305 //y2=1.375
r338 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.605 //y=1.375 //x2=63.715 //y2=1.375
r339 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.605 //y=1.375 //x2=63.495 //y2=1.375
r340 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=68.45 //y=4.7 //x2=68.45 //y2=4.7
r341 (  57 59 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=68.45 //y=2.59 //x2=68.45 //y2=4.7
r342 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=68.45 //y=2.08 //x2=68.45 //y2=2.08
r343 (  54 57 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=68.45 //y=2.08 //x2=68.45 //y2=2.59
r344 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.64 //y=4.7 //x2=63.64 //y2=4.7
r345 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=63.64 //y=2.59 //x2=63.64 //y2=4.7
r346 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.64 //y=2.08 //x2=63.64 //y2=2.08
r347 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=63.64 //y=2.08 //x2=63.64 //y2=2.59
r348 (  42 44 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=61.79 //y=5.07 //x2=61.79 //y2=2.59
r349 (  41 44 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=61.79 //y=1.75 //x2=61.79 //y2=2.59
r350 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=61.705 //y=1.665 //x2=61.79 //y2=1.75
r351 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=61.705 //y=1.665 //x2=61.39 //y2=1.665
r352 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=61.305 //y=1.58 //x2=61.39 //y2=1.665
r353 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=61.305 //y=1.58 //x2=61.305 //y2=1.01
r354 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.095 //y=5.155 //x2=61.01 //y2=5.155
r355 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=61.705 //y=5.155 //x2=61.79 //y2=5.07
r356 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=61.705 //y=5.155 //x2=61.095 //y2=5.155
r357 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.01 //y=5.24 //x2=61.01 //y2=5.155
r358 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=61.01 //y=5.24 //x2=61.01 //y2=5.725
r359 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.215 //y=5.155 //x2=60.13 //y2=5.155
r360 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.925 //y=5.155 //x2=61.01 //y2=5.155
r361 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=60.925 //y=5.155 //x2=60.215 //y2=5.155
r362 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.13 //y=5.24 //x2=60.13 //y2=5.155
r363 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.13 //y=5.24 //x2=60.13 //y2=5.725
r364 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.045 //y=5.155 //x2=60.13 //y2=5.155
r365 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=60.045 //y=5.155 //x2=59.335 //y2=5.155
r366 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=59.25 //y=5.24 //x2=59.335 //y2=5.155
r367 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.25 //y=5.24 //x2=59.25 //y2=5.725
r368 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=68.45 //y=2.59 //x2=68.45 //y2=2.59
r369 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=63.64 //y=2.59 //x2=63.64 //y2=2.59
r370 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=61.79 //y=2.59 //x2=61.79 //y2=2.59
r371 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.755 //y=2.59 //x2=63.64 //y2=2.59
r372 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=68.335 //y=2.59 //x2=68.45 //y2=2.59
r373 (  3 4 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=68.335 //y=2.59 //x2=63.755 //y2=2.59
r374 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=61.905 //y=2.59 //x2=61.79 //y2=2.59
r375 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.525 //y=2.59 //x2=63.64 //y2=2.59
r376 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=63.525 //y=2.59 //x2=61.905 //y2=2.59
ends PM_TMRDFFSNRNQX1\%noxref_16

subckt PM_TMRDFFSNRNQX1\%noxref_17 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 \
 53 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c168 ( 85 0 ) capacitor c=0.023087f //x=70.485 //y=5.02
c169 ( 84 0 ) capacitor c=0.023519f //x=69.605 //y=5.02
c170 ( 83 0 ) capacitor c=0.0224735f //x=68.725 //y=5.02
c171 ( 81 0 ) capacitor c=0.00853354f //x=70.735 //y=0.915
c172 ( 69 0 ) capacitor c=0.0547611f //x=73.535 //y=4.79
c173 ( 68 0 ) capacitor c=0.0294456f //x=73.825 //y=4.79
c174 ( 67 0 ) capacitor c=0.0347816f //x=73.49 //y=1.22
c175 ( 66 0 ) capacitor c=0.0187487f //x=73.49 //y=0.875
c176 ( 60 0 ) capacitor c=0.0137055f //x=73.335 //y=1.375
c177 ( 58 0 ) capacitor c=0.0149861f //x=73.335 //y=0.72
c178 ( 57 0 ) capacitor c=0.096037f //x=72.96 //y=1.915
c179 ( 56 0 ) capacitor c=0.0228993f //x=72.96 //y=1.53
c180 ( 55 0 ) capacitor c=0.0234352f //x=72.96 //y=1.22
c181 ( 54 0 ) capacitor c=0.0198724f //x=72.96 //y=0.875
c182 ( 53 0 ) capacitor c=0.109949f //x=73.9 //y=6.02
c183 ( 52 0 ) capacitor c=0.158483f //x=73.46 //y=6.02
c184 ( 50 0 ) capacitor c=9.74268e-19 //x=70.63 //y=5.155
c185 ( 49 0 ) capacitor c=0.00191414f //x=69.75 //y=5.155
c186 ( 42 0 ) capacitor c=0.0911502f //x=73.26 //y=2.08
c187 ( 40 0 ) capacitor c=0.103494f //x=71.41 //y=2.59
c188 ( 36 0 ) capacitor c=0.00398962f //x=71.01 //y=1.665
c189 ( 35 0 ) capacitor c=0.0137288f //x=71.325 //y=1.665
c190 ( 29 0 ) capacitor c=0.0276208f //x=71.325 //y=5.155
c191 ( 21 0 ) capacitor c=0.0169868f //x=70.545 //y=5.155
c192 ( 14 0 ) capacitor c=0.00316998f //x=68.955 //y=5.155
c193 ( 13 0 ) capacitor c=0.014258f //x=69.665 //y=5.155
c194 ( 2 0 ) capacitor c=0.00808366f //x=71.525 //y=2.59
c195 ( 1 0 ) capacitor c=0.0351856f //x=73.145 //y=2.59
r196 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=73.825 //y=4.79 //x2=73.9 //y2=4.865
r197 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=73.825 //y=4.79 //x2=73.535 //y2=4.79
r198 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.49 //y=1.22 //x2=73.45 //y2=1.375
r199 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.49 //y=0.875 //x2=73.45 //y2=0.72
r200 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=73.49 //y=0.875 //x2=73.49 //y2=1.22
r201 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=73.46 //y=4.865 //x2=73.535 //y2=4.79
r202 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=73.46 //y=4.865 //x2=73.26 //y2=4.7
r203 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.115 //y=1.375 //x2=73 //y2=1.375
r204 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.335 //y=1.375 //x2=73.45 //y2=1.375
r205 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.115 //y=0.72 //x2=73 //y2=0.72
r206 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.335 //y=0.72 //x2=73.45 //y2=0.72
r207 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=73.335 //y=0.72 //x2=73.115 //y2=0.72
r208 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=72.96 //y=1.915 //x2=73.26 //y2=2.08
r209 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.96 //y=1.53 //x2=73 //y2=1.375
r210 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=72.96 //y=1.53 //x2=72.96 //y2=1.915
r211 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.96 //y=1.22 //x2=73 //y2=1.375
r212 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.96 //y=0.875 //x2=73 //y2=0.72
r213 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=72.96 //y=0.875 //x2=72.96 //y2=1.22
r214 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=73.9 //y=6.02 //x2=73.9 //y2=4.865
r215 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=73.46 //y=6.02 //x2=73.46 //y2=4.865
r216 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=73.225 //y=1.375 //x2=73.335 //y2=1.375
r217 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=73.225 //y=1.375 //x2=73.115 //y2=1.375
r218 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=73.26 //y=4.7 //x2=73.26 //y2=4.7
r219 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=73.26 //y=2.59 //x2=73.26 //y2=4.7
r220 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=73.26 //y=2.08 //x2=73.26 //y2=2.08
r221 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=73.26 //y=2.08 //x2=73.26 //y2=2.59
r222 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=71.41 //y=5.07 //x2=71.41 //y2=2.59
r223 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=71.41 //y=1.75 //x2=71.41 //y2=2.59
r224 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=71.325 //y=1.665 //x2=71.41 //y2=1.75
r225 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=71.325 //y=1.665 //x2=71.01 //y2=1.665
r226 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=70.925 //y=1.58 //x2=71.01 //y2=1.665
r227 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=70.925 //y=1.58 //x2=70.925 //y2=1.01
r228 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.715 //y=5.155 //x2=70.63 //y2=5.155
r229 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=71.325 //y=5.155 //x2=71.41 //y2=5.07
r230 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=71.325 //y=5.155 //x2=70.715 //y2=5.155
r231 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.63 //y=5.24 //x2=70.63 //y2=5.155
r232 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=70.63 //y=5.24 //x2=70.63 //y2=5.725
r233 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.835 //y=5.155 //x2=69.75 //y2=5.155
r234 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.545 //y=5.155 //x2=70.63 //y2=5.155
r235 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=70.545 //y=5.155 //x2=69.835 //y2=5.155
r236 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.75 //y=5.24 //x2=69.75 //y2=5.155
r237 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=69.75 //y=5.24 //x2=69.75 //y2=5.725
r238 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.665 //y=5.155 //x2=69.75 //y2=5.155
r239 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=69.665 //y=5.155 //x2=68.955 //y2=5.155
r240 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=68.87 //y=5.24 //x2=68.955 //y2=5.155
r241 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=68.87 //y=5.24 //x2=68.87 //y2=5.725
r242 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=73.26 //y=2.59 //x2=73.26 //y2=2.59
r243 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=71.41 //y=2.59 //x2=71.41 //y2=2.59
r244 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=71.525 //y=2.59 //x2=71.41 //y2=2.59
r245 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=73.145 //y=2.59 //x2=73.26 //y2=2.59
r246 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=73.145 //y=2.59 //x2=71.525 //y2=2.59
ends PM_TMRDFFSNRNQX1\%noxref_17

subckt PM_TMRDFFSNRNQX1\%CLK ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 31 \
 32 33 34 36 46 55 64 73 81 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 \
 104 105 106 107 108 109 111 117 118 119 120 121 126 127 128 130 136 137 138 \
 139 140 145 146 147 149 155 156 157 158 159 164 165 166 168 174 175 176 177 \
 178 183 184 185 187 193 194 195 196 197 202 203 204 206 212 213 214 215 216 \
 224 235 246 257 268 279 )
c715 ( 279 0 ) capacitor c=0.0333177f //x=74.37 //y=4.7
c716 ( 268 0 ) capacitor c=0.0333177f //x=64.75 //y=4.7
c717 ( 257 0 ) capacitor c=0.0333177f //x=45.51 //y=4.7
c718 ( 246 0 ) capacitor c=0.0333177f //x=35.89 //y=4.7
c719 ( 235 0 ) capacitor c=0.0334842f //x=16.65 //y=4.7
c720 ( 224 0 ) capacitor c=0.0334842f //x=7.03 //y=4.7
c721 ( 216 0 ) capacitor c=0.0252241f //x=74.705 //y=4.79
c722 ( 215 0 ) capacitor c=0.0825763f //x=74.46 //y=1.915
c723 ( 214 0 ) capacitor c=0.0170266f //x=74.46 //y=1.45
c724 ( 213 0 ) capacitor c=0.018609f //x=74.46 //y=1.22
c725 ( 212 0 ) capacitor c=0.0187309f //x=74.46 //y=0.91
c726 ( 206 0 ) capacitor c=0.014725f //x=74.305 //y=1.375
c727 ( 204 0 ) capacitor c=0.0146567f //x=74.305 //y=0.755
c728 ( 203 0 ) capacitor c=0.0335408f //x=73.935 //y=1.22
c729 ( 202 0 ) capacitor c=0.0173761f //x=73.935 //y=0.91
c730 ( 197 0 ) capacitor c=0.0246783f //x=65.085 //y=4.79
c731 ( 196 0 ) capacitor c=0.0825763f //x=64.84 //y=1.915
c732 ( 195 0 ) capacitor c=0.0170266f //x=64.84 //y=1.45
c733 ( 194 0 ) capacitor c=0.018609f //x=64.84 //y=1.22
c734 ( 193 0 ) capacitor c=0.0187309f //x=64.84 //y=0.91
c735 ( 187 0 ) capacitor c=0.014725f //x=64.685 //y=1.375
c736 ( 185 0 ) capacitor c=0.0146567f //x=64.685 //y=0.755
c737 ( 184 0 ) capacitor c=0.0335408f //x=64.315 //y=1.22
c738 ( 183 0 ) capacitor c=0.0173761f //x=64.315 //y=0.91
c739 ( 178 0 ) capacitor c=0.0246783f //x=45.845 //y=4.79
c740 ( 177 0 ) capacitor c=0.0825763f //x=45.6 //y=1.915
c741 ( 176 0 ) capacitor c=0.0170266f //x=45.6 //y=1.45
c742 ( 175 0 ) capacitor c=0.018609f //x=45.6 //y=1.22
c743 ( 174 0 ) capacitor c=0.0187309f //x=45.6 //y=0.91
c744 ( 168 0 ) capacitor c=0.014725f //x=45.445 //y=1.375
c745 ( 166 0 ) capacitor c=0.0146567f //x=45.445 //y=0.755
c746 ( 165 0 ) capacitor c=0.0335408f //x=45.075 //y=1.22
c747 ( 164 0 ) capacitor c=0.0173761f //x=45.075 //y=0.91
c748 ( 159 0 ) capacitor c=0.0246783f //x=36.225 //y=4.79
c749 ( 158 0 ) capacitor c=0.0825763f //x=35.98 //y=1.915
c750 ( 157 0 ) capacitor c=0.0170266f //x=35.98 //y=1.45
c751 ( 156 0 ) capacitor c=0.018609f //x=35.98 //y=1.22
c752 ( 155 0 ) capacitor c=0.0187309f //x=35.98 //y=0.91
c753 ( 149 0 ) capacitor c=0.014725f //x=35.825 //y=1.375
c754 ( 147 0 ) capacitor c=0.0146567f //x=35.825 //y=0.755
c755 ( 146 0 ) capacitor c=0.0335408f //x=35.455 //y=1.22
c756 ( 145 0 ) capacitor c=0.0173761f //x=35.455 //y=0.91
c757 ( 140 0 ) capacitor c=0.0245352f //x=16.985 //y=4.79
c758 ( 139 0 ) capacitor c=0.0825763f //x=16.74 //y=1.915
c759 ( 138 0 ) capacitor c=0.0170266f //x=16.74 //y=1.45
c760 ( 137 0 ) capacitor c=0.018609f //x=16.74 //y=1.22
c761 ( 136 0 ) capacitor c=0.0187309f //x=16.74 //y=0.91
c762 ( 130 0 ) capacitor c=0.014725f //x=16.585 //y=1.375
c763 ( 128 0 ) capacitor c=0.0146567f //x=16.585 //y=0.755
c764 ( 127 0 ) capacitor c=0.0335408f //x=16.215 //y=1.22
c765 ( 126 0 ) capacitor c=0.0173761f //x=16.215 //y=0.91
c766 ( 121 0 ) capacitor c=0.0245352f //x=7.365 //y=4.79
c767 ( 120 0 ) capacitor c=0.0825763f //x=7.12 //y=1.915
c768 ( 119 0 ) capacitor c=0.0170266f //x=7.12 //y=1.45
c769 ( 118 0 ) capacitor c=0.018609f //x=7.12 //y=1.22
c770 ( 117 0 ) capacitor c=0.0187309f //x=7.12 //y=0.91
c771 ( 111 0 ) capacitor c=0.014725f //x=6.965 //y=1.375
c772 ( 109 0 ) capacitor c=0.0146567f //x=6.965 //y=0.755
c773 ( 108 0 ) capacitor c=0.0335408f //x=6.595 //y=1.22
c774 ( 107 0 ) capacitor c=0.0173761f //x=6.595 //y=0.91
c775 ( 106 0 ) capacitor c=0.109949f //x=74.78 //y=6.02
c776 ( 105 0 ) capacitor c=0.109956f //x=74.34 //y=6.02
c777 ( 104 0 ) capacitor c=0.109949f //x=65.16 //y=6.02
c778 ( 103 0 ) capacitor c=0.109956f //x=64.72 //y=6.02
c779 ( 102 0 ) capacitor c=0.109949f //x=45.92 //y=6.02
c780 ( 101 0 ) capacitor c=0.109956f //x=45.48 //y=6.02
c781 ( 100 0 ) capacitor c=0.109949f //x=36.3 //y=6.02
c782 ( 99 0 ) capacitor c=0.109956f //x=35.86 //y=6.02
c783 ( 98 0 ) capacitor c=0.110114f //x=17.06 //y=6.02
c784 ( 97 0 ) capacitor c=0.11012f //x=16.62 //y=6.02
c785 ( 96 0 ) capacitor c=0.110114f //x=7.44 //y=6.02
c786 ( 95 0 ) capacitor c=0.11012f //x=7 //y=6.02
c787 ( 81 0 ) capacitor c=0.0880092f //x=74.37 //y=2.08
c788 ( 73 0 ) capacitor c=0.0867127f //x=64.75 //y=2.08
c789 ( 64 0 ) capacitor c=0.0882702f //x=45.51 //y=2.08
c790 ( 55 0 ) capacitor c=0.088164f //x=35.89 //y=2.08
c791 ( 46 0 ) capacitor c=0.0899873f //x=16.65 //y=2.08
c792 ( 36 0 ) capacitor c=0.0925246f //x=7.03 //y=2.08
c793 ( 10 0 ) capacitor c=0.0052048f //x=64.865 //y=4.44
c794 ( 9 0 ) capacitor c=0.124137f //x=74.255 //y=4.44
c795 ( 8 0 ) capacitor c=0.00494979f //x=45.625 //y=4.44
c796 ( 7 0 ) capacitor c=0.255004f //x=64.635 //y=4.44
c797 ( 6 0 ) capacitor c=0.00494979f //x=36.005 //y=4.44
c798 ( 5 0 ) capacitor c=0.117333f //x=45.395 //y=4.44
c799 ( 4 0 ) capacitor c=0.00697397f //x=16.765 //y=4.44
c800 ( 3 0 ) capacitor c=0.345925f //x=35.775 //y=4.44
c801 ( 2 0 ) capacitor c=0.0154455f //x=7.145 //y=4.44
c802 ( 1 0 ) capacitor c=0.212324f //x=16.535 //y=4.44
r803 (  281 282 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=74.37 //y=4.79 //x2=74.37 //y2=4.865
r804 (  279 281 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=74.37 //y=4.7 //x2=74.37 //y2=4.79
r805 (  270 271 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=64.75 //y=4.79 //x2=64.75 //y2=4.865
r806 (  268 270 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=64.75 //y=4.7 //x2=64.75 //y2=4.79
r807 (  259 260 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=45.51 //y=4.79 //x2=45.51 //y2=4.865
r808 (  257 259 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=45.51 //y=4.7 //x2=45.51 //y2=4.79
r809 (  248 249 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=35.89 //y=4.79 //x2=35.89 //y2=4.865
r810 (  246 248 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=35.89 //y=4.7 //x2=35.89 //y2=4.79
r811 (  237 238 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=16.65 //y=4.79 //x2=16.65 //y2=4.865
r812 (  235 237 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=16.65 //y=4.7 //x2=16.65 //y2=4.79
r813 (  226 227 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.79 //x2=7.03 //y2=4.865
r814 (  224 226 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.7 //x2=7.03 //y2=4.79
r815 (  217 281 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=74.505 //y=4.79 //x2=74.37 //y2=4.79
r816 (  216 218 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=74.705 //y=4.79 //x2=74.78 //y2=4.865
r817 (  216 217 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=74.705 //y=4.79 //x2=74.505 //y2=4.79
r818 (  215 286 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=74.46 //y=1.915 //x2=74.385 //y2=2.08
r819 (  214 284 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=74.46 //y=1.45 //x2=74.42 //y2=1.375
r820 (  214 215 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=74.46 //y=1.45 //x2=74.46 //y2=1.915
r821 (  213 284 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.46 //y=1.22 //x2=74.42 //y2=1.375
r822 (  212 283 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.46 //y=0.91 //x2=74.42 //y2=0.755
r823 (  212 213 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=74.46 //y=0.91 //x2=74.46 //y2=1.22
r824 (  207 277 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.09 //y=1.375 //x2=73.975 //y2=1.375
r825 (  206 284 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.305 //y=1.375 //x2=74.42 //y2=1.375
r826 (  205 276 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.09 //y=0.755 //x2=73.975 //y2=0.755
r827 (  204 283 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.305 //y=0.755 //x2=74.42 //y2=0.755
r828 (  204 205 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=74.305 //y=0.755 //x2=74.09 //y2=0.755
r829 (  203 277 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.935 //y=1.22 //x2=73.975 //y2=1.375
r830 (  202 276 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.935 //y=0.91 //x2=73.975 //y2=0.755
r831 (  202 203 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=73.935 //y=0.91 //x2=73.935 //y2=1.22
r832 (  198 270 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=64.885 //y=4.79 //x2=64.75 //y2=4.79
r833 (  197 199 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=65.085 //y=4.79 //x2=65.16 //y2=4.865
r834 (  197 198 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=65.085 //y=4.79 //x2=64.885 //y2=4.79
r835 (  196 275 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=64.84 //y=1.915 //x2=64.765 //y2=2.08
r836 (  195 273 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=64.84 //y=1.45 //x2=64.8 //y2=1.375
r837 (  195 196 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=64.84 //y=1.45 //x2=64.84 //y2=1.915
r838 (  194 273 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.84 //y=1.22 //x2=64.8 //y2=1.375
r839 (  193 272 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.84 //y=0.91 //x2=64.8 //y2=0.755
r840 (  193 194 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=64.84 //y=0.91 //x2=64.84 //y2=1.22
r841 (  188 266 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.47 //y=1.375 //x2=64.355 //y2=1.375
r842 (  187 273 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.685 //y=1.375 //x2=64.8 //y2=1.375
r843 (  186 265 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.47 //y=0.755 //x2=64.355 //y2=0.755
r844 (  185 272 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.685 //y=0.755 //x2=64.8 //y2=0.755
r845 (  185 186 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=64.685 //y=0.755 //x2=64.47 //y2=0.755
r846 (  184 266 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.315 //y=1.22 //x2=64.355 //y2=1.375
r847 (  183 265 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.315 //y=0.91 //x2=64.355 //y2=0.755
r848 (  183 184 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=64.315 //y=0.91 //x2=64.315 //y2=1.22
r849 (  179 259 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=45.645 //y=4.79 //x2=45.51 //y2=4.79
r850 (  178 180 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=45.845 //y=4.79 //x2=45.92 //y2=4.865
r851 (  178 179 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=45.845 //y=4.79 //x2=45.645 //y2=4.79
r852 (  177 264 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=45.6 //y=1.915 //x2=45.525 //y2=2.08
r853 (  176 262 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=45.6 //y=1.45 //x2=45.56 //y2=1.375
r854 (  176 177 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=45.6 //y=1.45 //x2=45.6 //y2=1.915
r855 (  175 262 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.6 //y=1.22 //x2=45.56 //y2=1.375
r856 (  174 261 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.6 //y=0.91 //x2=45.56 //y2=0.755
r857 (  174 175 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=45.6 //y=0.91 //x2=45.6 //y2=1.22
r858 (  169 255 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.23 //y=1.375 //x2=45.115 //y2=1.375
r859 (  168 262 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.445 //y=1.375 //x2=45.56 //y2=1.375
r860 (  167 254 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.23 //y=0.755 //x2=45.115 //y2=0.755
r861 (  166 261 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.445 //y=0.755 //x2=45.56 //y2=0.755
r862 (  166 167 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=45.445 //y=0.755 //x2=45.23 //y2=0.755
r863 (  165 255 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.075 //y=1.22 //x2=45.115 //y2=1.375
r864 (  164 254 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.075 //y=0.91 //x2=45.115 //y2=0.755
r865 (  164 165 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=45.075 //y=0.91 //x2=45.075 //y2=1.22
r866 (  160 248 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=36.025 //y=4.79 //x2=35.89 //y2=4.79
r867 (  159 161 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=36.225 //y=4.79 //x2=36.3 //y2=4.865
r868 (  159 160 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=36.225 //y=4.79 //x2=36.025 //y2=4.79
r869 (  158 253 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=35.98 //y=1.915 //x2=35.905 //y2=2.08
r870 (  157 251 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=35.98 //y=1.45 //x2=35.94 //y2=1.375
r871 (  157 158 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=35.98 //y=1.45 //x2=35.98 //y2=1.915
r872 (  156 251 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.98 //y=1.22 //x2=35.94 //y2=1.375
r873 (  155 250 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.98 //y=0.91 //x2=35.94 //y2=0.755
r874 (  155 156 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=35.98 //y=0.91 //x2=35.98 //y2=1.22
r875 (  150 244 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.61 //y=1.375 //x2=35.495 //y2=1.375
r876 (  149 251 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.825 //y=1.375 //x2=35.94 //y2=1.375
r877 (  148 243 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.61 //y=0.755 //x2=35.495 //y2=0.755
r878 (  147 250 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.825 //y=0.755 //x2=35.94 //y2=0.755
r879 (  147 148 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=35.825 //y=0.755 //x2=35.61 //y2=0.755
r880 (  146 244 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.455 //y=1.22 //x2=35.495 //y2=1.375
r881 (  145 243 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.455 //y=0.91 //x2=35.495 //y2=0.755
r882 (  145 146 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=35.455 //y=0.91 //x2=35.455 //y2=1.22
r883 (  141 237 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=16.785 //y=4.79 //x2=16.65 //y2=4.79
r884 (  140 142 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=16.985 //y=4.79 //x2=17.06 //y2=4.865
r885 (  140 141 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=16.985 //y=4.79 //x2=16.785 //y2=4.79
r886 (  139 242 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.915 //x2=16.665 //y2=2.08
r887 (  138 240 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.45 //x2=16.7 //y2=1.375
r888 (  138 139 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.45 //x2=16.74 //y2=1.915
r889 (  137 240 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.22 //x2=16.7 //y2=1.375
r890 (  136 239 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.74 //y=0.91 //x2=16.7 //y2=0.755
r891 (  136 137 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=16.74 //y=0.91 //x2=16.74 //y2=1.22
r892 (  131 233 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.37 //y=1.375 //x2=16.255 //y2=1.375
r893 (  130 240 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.585 //y=1.375 //x2=16.7 //y2=1.375
r894 (  129 232 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.37 //y=0.755 //x2=16.255 //y2=0.755
r895 (  128 239 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.585 //y=0.755 //x2=16.7 //y2=0.755
r896 (  128 129 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=16.585 //y=0.755 //x2=16.37 //y2=0.755
r897 (  127 233 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.215 //y=1.22 //x2=16.255 //y2=1.375
r898 (  126 232 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.215 //y=0.91 //x2=16.255 //y2=0.755
r899 (  126 127 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=16.215 //y=0.91 //x2=16.215 //y2=1.22
r900 (  122 226 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=7.165 //y=4.79 //x2=7.03 //y2=4.79
r901 (  121 123 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.44 //y2=4.865
r902 (  121 122 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.165 //y2=4.79
r903 (  120 231 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.915 //x2=7.045 //y2=2.08
r904 (  119 229 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.08 //y2=1.375
r905 (  119 120 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.12 //y2=1.915
r906 (  118 229 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.22 //x2=7.08 //y2=1.375
r907 (  117 228 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.08 //y2=0.755
r908 (  117 118 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.12 //y2=1.22
r909 (  112 222 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=1.375 //x2=6.635 //y2=1.375
r910 (  111 229 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=1.375 //x2=7.08 //y2=1.375
r911 (  110 221 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=0.755 //x2=6.635 //y2=0.755
r912 (  109 228 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=7.08 //y2=0.755
r913 (  109 110 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=6.75 //y2=0.755
r914 (  108 222 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=1.22 //x2=6.635 //y2=1.375
r915 (  107 221 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.635 //y2=0.755
r916 (  107 108 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.595 //y2=1.22
r917 (  106 218 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=74.78 //y=6.02 //x2=74.78 //y2=4.865
r918 (  105 282 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=74.34 //y=6.02 //x2=74.34 //y2=4.865
r919 (  104 199 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=65.16 //y=6.02 //x2=65.16 //y2=4.865
r920 (  103 271 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=64.72 //y=6.02 //x2=64.72 //y2=4.865
r921 (  102 180 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.92 //y=6.02 //x2=45.92 //y2=4.865
r922 (  101 260 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.48 //y=6.02 //x2=45.48 //y2=4.865
r923 (  100 161 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=36.3 //y=6.02 //x2=36.3 //y2=4.865
r924 (  99 249 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.86 //y=6.02 //x2=35.86 //y2=4.865
r925 (  98 142 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.06 //y=6.02 //x2=17.06 //y2=4.865
r926 (  97 238 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.62 //y=6.02 //x2=16.62 //y2=4.865
r927 (  96 123 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.44 //y=6.02 //x2=7.44 //y2=4.865
r928 (  95 227 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7 //y=6.02 //x2=7 //y2=4.865
r929 (  94 206 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=74.197 //y=1.375 //x2=74.305 //y2=1.375
r930 (  94 207 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=74.197 //y=1.375 //x2=74.09 //y2=1.375
r931 (  93 187 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=64.577 //y=1.375 //x2=64.685 //y2=1.375
r932 (  93 188 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=64.577 //y=1.375 //x2=64.47 //y2=1.375
r933 (  92 168 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=45.337 //y=1.375 //x2=45.445 //y2=1.375
r934 (  92 169 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=45.337 //y=1.375 //x2=45.23 //y2=1.375
r935 (  91 149 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=35.717 //y=1.375 //x2=35.825 //y2=1.375
r936 (  91 150 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=35.717 //y=1.375 //x2=35.61 //y2=1.375
r937 (  90 130 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=16.477 //y=1.375 //x2=16.585 //y2=1.375
r938 (  90 131 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=16.477 //y=1.375 //x2=16.37 //y2=1.375
r939 (  89 111 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.965 //y2=1.375
r940 (  89 112 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.75 //y2=1.375
r941 (  87 279 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=74.37 //y=4.7 //x2=74.37 //y2=4.7
r942 (  81 286 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=74.37 //y=2.08 //x2=74.37 //y2=2.08
r943 (  78 268 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=64.75 //y=4.7 //x2=64.75 //y2=4.7
r944 (  73 275 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=64.75 //y=2.08 //x2=64.75 //y2=2.08
r945 (  70 257 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.51 //y=4.7 //x2=45.51 //y2=4.7
r946 (  64 264 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.51 //y=2.08 //x2=45.51 //y2=2.08
r947 (  61 246 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.89 //y=4.7 //x2=35.89 //y2=4.7
r948 (  55 253 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.89 //y=2.08 //x2=35.89 //y2=2.08
r949 (  52 235 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=4.7 //x2=16.65 //y2=4.7
r950 (  46 242 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=2.08 //x2=16.65 //y2=2.08
r951 (  43 224 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=4.7 //x2=7.03 //y2=4.7
r952 (  36 231 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=2.08 //x2=7.03 //y2=2.08
r953 (  34 87 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=74.37 //y=4.44 //x2=74.37 //y2=4.7
r954 (  33 34 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=74.37 //y=2.59 //x2=74.37 //y2=4.44
r955 (  33 81 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=74.37 //y=2.59 //x2=74.37 //y2=2.08
r956 (  32 78 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=64.75 //y=4.44 //x2=64.75 //y2=4.7
r957 (  32 73 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=64.75 //y=4.44 //x2=64.75 //y2=2.08
r958 (  31 70 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=45.51 //y=4.44 //x2=45.51 //y2=4.7
r959 (  30 31 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=45.51 //y=2.59 //x2=45.51 //y2=4.44
r960 (  30 64 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=45.51 //y=2.59 //x2=45.51 //y2=2.08
r961 (  29 61 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=35.89 //y=4.44 //x2=35.89 //y2=4.7
r962 (  28 29 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=35.89 //y=3.7 //x2=35.89 //y2=4.44
r963 (  28 55 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=35.89 //y=3.7 //x2=35.89 //y2=2.08
r964 (  27 52 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.44 //x2=16.65 //y2=4.7
r965 (  26 27 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.59 //x2=16.65 //y2=4.44
r966 (  26 46 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.59 //x2=16.65 //y2=2.08
r967 (  25 43 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=7.03 //y=4.44 //x2=7.03 //y2=4.7
r968 (  24 25 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=7.03 //y=3.7 //x2=7.03 //y2=4.44
r969 (  23 24 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.96 //x2=7.03 //y2=3.7
r970 (  23 36 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.96 //x2=7.03 //y2=2.08
r971 (  22 34 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=74.37 //y=4.44 //x2=74.37 //y2=4.44
r972 (  20 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=64.75 //y=4.44 //x2=64.75 //y2=4.44
r973 (  18 31 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=45.51 //y=4.44 //x2=45.51 //y2=4.44
r974 (  16 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=35.89 //y=4.44 //x2=35.89 //y2=4.44
r975 (  14 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=16.65 //y=4.44 //x2=16.65 //y2=4.44
r976 (  12 25 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.03 //y=4.44 //x2=7.03 //y2=4.44
r977 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=64.865 //y=4.44 //x2=64.75 //y2=4.44
r978 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=74.255 //y=4.44 //x2=74.37 //y2=4.44
r979 (  9 10 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=74.255 //y=4.44 //x2=64.865 //y2=4.44
r980 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.625 //y=4.44 //x2=45.51 //y2=4.44
r981 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=64.635 //y=4.44 //x2=64.75 //y2=4.44
r982 (  7 8 ) resistor r=18.1393 //w=0.131 //l=19.01 //layer=m1 \
 //thickness=0.36 //x=64.635 //y=4.44 //x2=45.625 //y2=4.44
r983 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=36.005 //y=4.44 //x2=35.89 //y2=4.44
r984 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.395 //y=4.44 //x2=45.51 //y2=4.44
r985 (  5 6 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=45.395 //y=4.44 //x2=36.005 //y2=4.44
r986 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.765 //y=4.44 //x2=16.65 //y2=4.44
r987 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=35.775 //y=4.44 //x2=35.89 //y2=4.44
r988 (  3 4 ) resistor r=18.1393 //w=0.131 //l=19.01 //layer=m1 \
 //thickness=0.36 //x=35.775 //y=4.44 //x2=16.765 //y2=4.44
r989 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.145 //y=4.44 //x2=7.03 //y2=4.44
r990 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.535 //y=4.44 //x2=16.65 //y2=4.44
r991 (  1 2 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=16.535 //y=4.44 //x2=7.145 //y2=4.44
ends PM_TMRDFFSNRNQX1\%CLK

subckt PM_TMRDFFSNRNQX1\%noxref_19 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 \
 63 64 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 90 92 98 99 100 101 106 \
 107 112 123 125 126 127 )
c274 ( 127 0 ) capacitor c=0.023087f //x=65.675 //y=5.02
c275 ( 126 0 ) capacitor c=0.023519f //x=64.795 //y=5.02
c276 ( 125 0 ) capacitor c=0.0224735f //x=63.915 //y=5.02
c277 ( 123 0 ) capacitor c=0.00853354f //x=65.925 //y=0.915
c278 ( 112 0 ) capacitor c=0.0588394f //x=61.05 //y=4.7
c279 ( 107 0 ) capacitor c=0.0273931f //x=61.05 //y=1.915
c280 ( 106 0 ) capacitor c=0.0456313f //x=61.05 //y=2.08
c281 ( 101 0 ) capacitor c=0.0556143f //x=78.345 //y=4.79
c282 ( 100 0 ) capacitor c=0.0293157f //x=78.635 //y=4.79
c283 ( 99 0 ) capacitor c=0.0347816f //x=78.3 //y=1.22
c284 ( 98 0 ) capacitor c=0.0187487f //x=78.3 //y=0.875
c285 ( 92 0 ) capacitor c=0.0137055f //x=78.145 //y=1.375
c286 ( 90 0 ) capacitor c=0.0149861f //x=78.145 //y=0.72
c287 ( 89 0 ) capacitor c=0.096037f //x=77.77 //y=1.915
c288 ( 88 0 ) capacitor c=0.0228993f //x=77.77 //y=1.53
c289 ( 87 0 ) capacitor c=0.0234352f //x=77.77 //y=1.22
c290 ( 86 0 ) capacitor c=0.0198724f //x=77.77 //y=0.875
c291 ( 85 0 ) capacitor c=0.0432517f //x=61.57 //y=1.26
c292 ( 84 0 ) capacitor c=0.0200379f //x=61.57 //y=0.915
c293 ( 81 0 ) capacitor c=0.0148873f //x=61.415 //y=1.415
c294 ( 79 0 ) capacitor c=0.0157803f //x=61.415 //y=0.76
c295 ( 74 0 ) capacitor c=0.0218028f //x=61.04 //y=1.57
c296 ( 73 0 ) capacitor c=0.0207459f //x=61.04 //y=1.26
c297 ( 72 0 ) capacitor c=0.0194308f //x=61.04 //y=0.915
c298 ( 68 0 ) capacitor c=0.110114f //x=78.71 //y=6.02
c299 ( 67 0 ) capacitor c=0.158956f //x=78.27 //y=6.02
c300 ( 66 0 ) capacitor c=0.158754f //x=61.23 //y=6.02
c301 ( 65 0 ) capacitor c=0.109949f //x=60.79 //y=6.02
c302 ( 62 0 ) capacitor c=9.74268e-19 //x=65.82 //y=5.155
c303 ( 61 0 ) capacitor c=0.00191414f //x=64.94 //y=5.155
c304 ( 54 0 ) capacitor c=0.0959558f //x=78.07 //y=2.08
c305 ( 52 0 ) capacitor c=0.1027f //x=66.6 //y=3.33
c306 ( 48 0 ) capacitor c=0.00398962f //x=66.2 //y=1.665
c307 ( 47 0 ) capacitor c=0.0137288f //x=66.515 //y=1.665
c308 ( 41 0 ) capacitor c=0.0276208f //x=66.515 //y=5.155
c309 ( 33 0 ) capacitor c=0.0169868f //x=65.735 //y=5.155
c310 ( 26 0 ) capacitor c=0.00316998f //x=64.145 //y=5.155
c311 ( 25 0 ) capacitor c=0.014258f //x=64.855 //y=5.155
c312 ( 12 0 ) capacitor c=0.0814556f //x=61.05 //y=2.08
c313 ( 4 0 ) capacitor c=0.00551333f //x=66.715 //y=3.33
c314 ( 3 0 ) capacitor c=0.17826f //x=77.955 //y=3.33
c315 ( 2 0 ) capacitor c=0.0105808f //x=61.165 //y=3.33
c316 ( 1 0 ) capacitor c=0.077341f //x=66.485 //y=3.33
r317 (  106 107 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=61.05 //y=2.08 //x2=61.05 //y2=1.915
r318 (  100 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=78.635 //y=4.79 //x2=78.71 //y2=4.865
r319 (  100 101 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=78.635 //y=4.79 //x2=78.345 //y2=4.79
r320 (  99 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.3 //y=1.22 //x2=78.26 //y2=1.375
r321 (  98 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.3 //y=0.875 //x2=78.26 //y2=0.72
r322 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=78.3 //y=0.875 //x2=78.3 //y2=1.22
r323 (  95 101 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=78.27 //y=4.865 //x2=78.345 //y2=4.79
r324 (  95 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=78.27 //y=4.865 //x2=78.07 //y2=4.7
r325 (  93 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.925 //y=1.375 //x2=77.81 //y2=1.375
r326 (  92 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.145 //y=1.375 //x2=78.26 //y2=1.375
r327 (  91 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.925 //y=0.72 //x2=77.81 //y2=0.72
r328 (  90 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.145 //y=0.72 //x2=78.26 //y2=0.72
r329 (  90 91 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=78.145 //y=0.72 //x2=77.925 //y2=0.72
r330 (  89 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.915 //x2=78.07 //y2=2.08
r331 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.53 //x2=77.81 //y2=1.375
r332 (  88 89 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.53 //x2=77.77 //y2=1.915
r333 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.22 //x2=77.81 //y2=1.375
r334 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.77 //y=0.875 //x2=77.81 //y2=0.72
r335 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=77.77 //y=0.875 //x2=77.77 //y2=1.22
r336 (  85 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.57 //y=1.26 //x2=61.53 //y2=1.415
r337 (  84 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.57 //y=0.915 //x2=61.53 //y2=0.76
r338 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=61.57 //y=0.915 //x2=61.57 //y2=1.26
r339 (  82 110 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=61.195 //y=1.415 //x2=61.08 //y2=1.415
r340 (  81 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=61.415 //y=1.415 //x2=61.53 //y2=1.415
r341 (  80 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=61.195 //y=0.76 //x2=61.08 //y2=0.76
r342 (  79 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=61.415 //y=0.76 //x2=61.53 //y2=0.76
r343 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=61.415 //y=0.76 //x2=61.195 //y2=0.76
r344 (  76 112 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=61.23 //y=4.865 //x2=61.05 //y2=4.7
r345 (  74 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.04 //y=1.57 //x2=61.08 //y2=1.415
r346 (  74 107 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=61.04 //y=1.57 //x2=61.04 //y2=1.915
r347 (  73 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.04 //y=1.26 //x2=61.08 //y2=1.415
r348 (  72 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.04 //y=0.915 //x2=61.08 //y2=0.76
r349 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=61.04 //y=0.915 //x2=61.04 //y2=1.26
r350 (  69 112 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=60.79 //y=4.865 //x2=61.05 //y2=4.7
r351 (  68 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.71 //y=6.02 //x2=78.71 //y2=4.865
r352 (  67 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.27 //y=6.02 //x2=78.27 //y2=4.865
r353 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=61.23 //y=6.02 //x2=61.23 //y2=4.865
r354 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.79 //y=6.02 //x2=60.79 //y2=4.865
r355 (  64 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.035 //y=1.375 //x2=78.145 //y2=1.375
r356 (  64 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.035 //y=1.375 //x2=77.925 //y2=1.375
r357 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=61.305 //y=1.415 //x2=61.415 //y2=1.415
r358 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=61.305 //y=1.415 //x2=61.195 //y2=1.415
r359 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=78.07 //y=4.7 //x2=78.07 //y2=4.7
r360 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=78.07 //y=3.33 //x2=78.07 //y2=4.7
r361 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=78.07 //y=2.08 //x2=78.07 //y2=2.08
r362 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=78.07 //y=2.08 //x2=78.07 //y2=3.33
r363 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=66.6 //y=5.07 //x2=66.6 //y2=3.33
r364 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=66.6 //y=1.75 //x2=66.6 //y2=3.33
r365 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=66.515 //y=1.665 //x2=66.6 //y2=1.75
r366 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=66.515 //y=1.665 //x2=66.2 //y2=1.665
r367 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=66.115 //y=1.58 //x2=66.2 //y2=1.665
r368 (  43 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=66.115 //y=1.58 //x2=66.115 //y2=1.01
r369 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.905 //y=5.155 //x2=65.82 //y2=5.155
r370 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=66.515 //y=5.155 //x2=66.6 //y2=5.07
r371 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=66.515 //y=5.155 //x2=65.905 //y2=5.155
r372 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.82 //y=5.24 //x2=65.82 //y2=5.155
r373 (  35 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=65.82 //y=5.24 //x2=65.82 //y2=5.725
r374 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.025 //y=5.155 //x2=64.94 //y2=5.155
r375 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.735 //y=5.155 //x2=65.82 //y2=5.155
r376 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=65.735 //y=5.155 //x2=65.025 //y2=5.155
r377 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.94 //y=5.24 //x2=64.94 //y2=5.155
r378 (  27 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=64.94 //y=5.24 //x2=64.94 //y2=5.725
r379 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.855 //y=5.155 //x2=64.94 //y2=5.155
r380 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=64.855 //y=5.155 //x2=64.145 //y2=5.155
r381 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=64.06 //y=5.24 //x2=64.145 //y2=5.155
r382 (  19 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=64.06 //y=5.24 //x2=64.06 //y2=5.725
r383 (  17 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=61.05 //y=4.7 //x2=61.05 //y2=4.7
r384 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=61.05 //y=3.33 //x2=61.05 //y2=4.7
r385 (  12 106 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=61.05 //y=2.08 //x2=61.05 //y2=2.08
r386 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=61.05 //y=2.08 //x2=61.05 //y2=3.33
r387 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=78.07 //y=3.33 //x2=78.07 //y2=3.33
r388 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.6 //y=3.33 //x2=66.6 //y2=3.33
r389 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=61.05 //y=3.33 //x2=61.05 //y2=3.33
r390 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.715 //y=3.33 //x2=66.6 //y2=3.33
r391 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=77.955 //y=3.33 //x2=78.07 //y2=3.33
r392 (  3 4 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=77.955 //y=3.33 //x2=66.715 //y2=3.33
r393 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=61.165 //y=3.33 //x2=61.05 //y2=3.33
r394 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.485 //y=3.33 //x2=66.6 //y2=3.33
r395 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=66.485 //y=3.33 //x2=61.165 //y2=3.33
ends PM_TMRDFFSNRNQX1\%noxref_19

subckt PM_TMRDFFSNRNQX1\%RN ( 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 35 36 37 \
 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 \
 65 78 87 97 108 117 127 138 147 156 157 158 159 160 161 162 163 164 165 166 \
 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 \
 187 193 194 195 196 197 205 206 207 212 214 217 218 219 220 221 223 229 230 \
 231 232 233 238 239 240 242 248 249 250 251 252 260 261 262 267 269 272 273 \
 274 275 276 278 284 285 286 287 288 293 294 295 297 303 304 305 306 307 315 \
 316 317 322 324 327 328 329 330 331 333 339 340 341 342 343 351 360 361 366 \
 372 383 392 393 398 404 415 424 425 430 436 )
c1111 ( 436 0 ) capacitor c=0.0335551f //x=79.18 //y=4.7
c1112 ( 430 0 ) capacitor c=0.0584472f //x=75.48 //y=4.7
c1113 ( 425 0 ) capacitor c=0.0273931f //x=75.48 //y=1.915
c1114 ( 424 0 ) capacitor c=0.0455604f //x=75.48 //y=2.08
c1115 ( 415 0 ) capacitor c=0.0333886f //x=59.94 //y=4.7
c1116 ( 404 0 ) capacitor c=0.0333886f //x=50.32 //y=4.7
c1117 ( 398 0 ) capacitor c=0.0589949f //x=46.62 //y=4.7
c1118 ( 393 0 ) capacitor c=0.0273931f //x=46.62 //y=1.915
c1119 ( 392 0 ) capacitor c=0.0455604f //x=46.62 //y=2.08
c1120 ( 383 0 ) capacitor c=0.0333886f //x=31.08 //y=4.7
c1121 ( 372 0 ) capacitor c=0.0335551f //x=21.46 //y=4.7
c1122 ( 366 0 ) capacitor c=0.058931f //x=17.76 //y=4.7
c1123 ( 361 0 ) capacitor c=0.0273931f //x=17.76 //y=1.915
c1124 ( 360 0 ) capacitor c=0.0455604f //x=17.76 //y=2.08
c1125 ( 351 0 ) capacitor c=0.0336203f //x=2.22 //y=4.7
c1126 ( 343 0 ) capacitor c=0.0245352f //x=79.515 //y=4.79
c1127 ( 342 0 ) capacitor c=0.0827272f //x=79.27 //y=1.915
c1128 ( 341 0 ) capacitor c=0.0170266f //x=79.27 //y=1.45
c1129 ( 340 0 ) capacitor c=0.018609f //x=79.27 //y=1.22
c1130 ( 339 0 ) capacitor c=0.0187309f //x=79.27 //y=0.91
c1131 ( 333 0 ) capacitor c=0.014725f //x=79.115 //y=1.375
c1132 ( 331 0 ) capacitor c=0.0146567f //x=79.115 //y=0.755
c1133 ( 330 0 ) capacitor c=0.0335408f //x=78.745 //y=1.22
c1134 ( 329 0 ) capacitor c=0.0173761f //x=78.745 //y=0.91
c1135 ( 328 0 ) capacitor c=0.0432517f //x=76 //y=1.26
c1136 ( 327 0 ) capacitor c=0.0200379f //x=76 //y=0.915
c1137 ( 324 0 ) capacitor c=0.0148873f //x=75.845 //y=1.415
c1138 ( 322 0 ) capacitor c=0.0157803f //x=75.845 //y=0.76
c1139 ( 317 0 ) capacitor c=0.0218028f //x=75.47 //y=1.57
c1140 ( 316 0 ) capacitor c=0.0207459f //x=75.47 //y=1.26
c1141 ( 315 0 ) capacitor c=0.0194308f //x=75.47 //y=0.915
c1142 ( 307 0 ) capacitor c=0.0246783f //x=60.275 //y=4.79
c1143 ( 306 0 ) capacitor c=0.0825033f //x=60.03 //y=1.915
c1144 ( 305 0 ) capacitor c=0.0170266f //x=60.03 //y=1.45
c1145 ( 304 0 ) capacitor c=0.018609f //x=60.03 //y=1.22
c1146 ( 303 0 ) capacitor c=0.0187309f //x=60.03 //y=0.91
c1147 ( 297 0 ) capacitor c=0.014725f //x=59.875 //y=1.375
c1148 ( 295 0 ) capacitor c=0.0146567f //x=59.875 //y=0.755
c1149 ( 294 0 ) capacitor c=0.0335408f //x=59.505 //y=1.22
c1150 ( 293 0 ) capacitor c=0.0173761f //x=59.505 //y=0.91
c1151 ( 288 0 ) capacitor c=0.0246783f //x=50.655 //y=4.79
c1152 ( 287 0 ) capacitor c=0.0825033f //x=50.41 //y=1.915
c1153 ( 286 0 ) capacitor c=0.0170266f //x=50.41 //y=1.45
c1154 ( 285 0 ) capacitor c=0.018609f //x=50.41 //y=1.22
c1155 ( 284 0 ) capacitor c=0.0187309f //x=50.41 //y=0.91
c1156 ( 278 0 ) capacitor c=0.014725f //x=50.255 //y=1.375
c1157 ( 276 0 ) capacitor c=0.0146567f //x=50.255 //y=0.755
c1158 ( 275 0 ) capacitor c=0.0335408f //x=49.885 //y=1.22
c1159 ( 274 0 ) capacitor c=0.0173761f //x=49.885 //y=0.91
c1160 ( 273 0 ) capacitor c=0.0432517f //x=47.14 //y=1.26
c1161 ( 272 0 ) capacitor c=0.0200379f //x=47.14 //y=0.915
c1162 ( 269 0 ) capacitor c=0.0148873f //x=46.985 //y=1.415
c1163 ( 267 0 ) capacitor c=0.0157803f //x=46.985 //y=0.76
c1164 ( 262 0 ) capacitor c=0.0218028f //x=46.61 //y=1.57
c1165 ( 261 0 ) capacitor c=0.0207459f //x=46.61 //y=1.26
c1166 ( 260 0 ) capacitor c=0.0194308f //x=46.61 //y=0.915
c1167 ( 252 0 ) capacitor c=0.0246783f //x=31.415 //y=4.79
c1168 ( 251 0 ) capacitor c=0.0825033f //x=31.17 //y=1.915
c1169 ( 250 0 ) capacitor c=0.0170266f //x=31.17 //y=1.45
c1170 ( 249 0 ) capacitor c=0.018609f //x=31.17 //y=1.22
c1171 ( 248 0 ) capacitor c=0.0187309f //x=31.17 //y=0.91
c1172 ( 242 0 ) capacitor c=0.014725f //x=31.015 //y=1.375
c1173 ( 240 0 ) capacitor c=0.0146567f //x=31.015 //y=0.755
c1174 ( 239 0 ) capacitor c=0.0335408f //x=30.645 //y=1.22
c1175 ( 238 0 ) capacitor c=0.0173761f //x=30.645 //y=0.91
c1176 ( 233 0 ) capacitor c=0.0245352f //x=21.795 //y=4.79
c1177 ( 232 0 ) capacitor c=0.0825033f //x=21.55 //y=1.915
c1178 ( 231 0 ) capacitor c=0.0170266f //x=21.55 //y=1.45
c1179 ( 230 0 ) capacitor c=0.018609f //x=21.55 //y=1.22
c1180 ( 229 0 ) capacitor c=0.0187309f //x=21.55 //y=0.91
c1181 ( 223 0 ) capacitor c=0.014725f //x=21.395 //y=1.375
c1182 ( 221 0 ) capacitor c=0.0146567f //x=21.395 //y=0.755
c1183 ( 220 0 ) capacitor c=0.0335408f //x=21.025 //y=1.22
c1184 ( 219 0 ) capacitor c=0.0173761f //x=21.025 //y=0.91
c1185 ( 218 0 ) capacitor c=0.0432517f //x=18.28 //y=1.26
c1186 ( 217 0 ) capacitor c=0.0200379f //x=18.28 //y=0.915
c1187 ( 214 0 ) capacitor c=0.0148873f //x=18.125 //y=1.415
c1188 ( 212 0 ) capacitor c=0.0157803f //x=18.125 //y=0.76
c1189 ( 207 0 ) capacitor c=0.0218028f //x=17.75 //y=1.57
c1190 ( 206 0 ) capacitor c=0.0207459f //x=17.75 //y=1.26
c1191 ( 205 0 ) capacitor c=0.0194308f //x=17.75 //y=0.915
c1192 ( 197 0 ) capacitor c=0.024933f //x=2.555 //y=4.79
c1193 ( 196 0 ) capacitor c=0.0826756f //x=2.31 //y=1.915
c1194 ( 195 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c1195 ( 194 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c1196 ( 193 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c1197 ( 187 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c1198 ( 185 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c1199 ( 184 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c1200 ( 183 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c1201 ( 182 0 ) capacitor c=0.110114f //x=79.59 //y=6.02
c1202 ( 181 0 ) capacitor c=0.11012f //x=79.15 //y=6.02
c1203 ( 180 0 ) capacitor c=0.158794f //x=75.66 //y=6.02
c1204 ( 179 0 ) capacitor c=0.11002f //x=75.22 //y=6.02
c1205 ( 178 0 ) capacitor c=0.109949f //x=60.35 //y=6.02
c1206 ( 177 0 ) capacitor c=0.109956f //x=59.91 //y=6.02
c1207 ( 176 0 ) capacitor c=0.109949f //x=50.73 //y=6.02
c1208 ( 175 0 ) capacitor c=0.109956f //x=50.29 //y=6.02
c1209 ( 174 0 ) capacitor c=0.158754f //x=46.8 //y=6.02
c1210 ( 173 0 ) capacitor c=0.109949f //x=46.36 //y=6.02
c1211 ( 172 0 ) capacitor c=0.109949f //x=31.49 //y=6.02
c1212 ( 171 0 ) capacitor c=0.109956f //x=31.05 //y=6.02
c1213 ( 170 0 ) capacitor c=0.110114f //x=21.87 //y=6.02
c1214 ( 169 0 ) capacitor c=0.11012f //x=21.43 //y=6.02
c1215 ( 168 0 ) capacitor c=0.158794f //x=17.94 //y=6.02
c1216 ( 167 0 ) capacitor c=0.110114f //x=17.5 //y=6.02
c1217 ( 166 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c1218 ( 165 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c1219 ( 147 0 ) capacitor c=0.0925003f //x=79.18 //y=2.08
c1220 ( 138 0 ) capacitor c=0.0818106f //x=75.48 //y=2.08
c1221 ( 127 0 ) capacitor c=0.092289f //x=59.94 //y=2.08
c1222 ( 117 0 ) capacitor c=0.0898148f //x=50.32 //y=2.08
c1223 ( 108 0 ) capacitor c=0.0797966f //x=46.62 //y=2.08
c1224 ( 97 0 ) capacitor c=0.092949f //x=31.08 //y=2.08
c1225 ( 87 0 ) capacitor c=0.0915318f //x=21.46 //y=2.08
c1226 ( 78 0 ) capacitor c=0.081834f //x=17.76 //y=2.08
c1227 ( 65 0 ) capacitor c=0.100124f //x=2.22 //y=2.08
c1228 ( 16 0 ) capacitor c=0.00626813f //x=75.595 //y=2.22
c1229 ( 15 0 ) capacitor c=0.0882914f //x=79.065 //y=2.22
c1230 ( 14 0 ) capacitor c=0.00683472f //x=60.055 //y=2.22
c1231 ( 13 0 ) capacitor c=0.318477f //x=75.365 //y=2.22
c1232 ( 12 0 ) capacitor c=0.0059254f //x=50.435 //y=2.22
c1233 ( 11 0 ) capacitor c=0.207602f //x=59.825 //y=2.22
c1234 ( 10 0 ) capacitor c=0.00618148f //x=46.735 //y=2.22
c1235 ( 9 0 ) capacitor c=0.0804516f //x=50.205 //y=2.22
c1236 ( 8 0 ) capacitor c=0.00683472f //x=31.195 //y=2.22
c1237 ( 7 0 ) capacitor c=0.318477f //x=46.505 //y=2.22
c1238 ( 6 0 ) capacitor c=0.00601205f //x=21.575 //y=2.22
c1239 ( 5 0 ) capacitor c=0.208107f //x=30.965 //y=2.22
c1240 ( 4 0 ) capacitor c=0.00626813f //x=17.875 //y=2.22
c1241 ( 3 0 ) capacitor c=0.0805381f //x=21.345 //y=2.22
c1242 ( 2 0 ) capacitor c=0.0163048f //x=2.335 //y=2.22
c1243 ( 1 0 ) capacitor c=0.330466f //x=17.645 //y=2.22
r1244 (  438 439 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=79.18 //y=4.79 //x2=79.18 //y2=4.865
r1245 (  436 438 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=79.18 //y=4.7 //x2=79.18 //y2=4.79
r1246 (  424 425 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=75.48 //y=2.08 //x2=75.48 //y2=1.915
r1247 (  417 418 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=59.94 //y=4.79 //x2=59.94 //y2=4.865
r1248 (  415 417 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=59.94 //y=4.7 //x2=59.94 //y2=4.79
r1249 (  406 407 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=50.32 //y=4.79 //x2=50.32 //y2=4.865
r1250 (  404 406 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=50.32 //y=4.7 //x2=50.32 //y2=4.79
r1251 (  392 393 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=46.62 //y=2.08 //x2=46.62 //y2=1.915
r1252 (  385 386 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=31.08 //y=4.79 //x2=31.08 //y2=4.865
r1253 (  383 385 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=31.08 //y=4.7 //x2=31.08 //y2=4.79
r1254 (  374 375 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=21.46 //y=4.79 //x2=21.46 //y2=4.865
r1255 (  372 374 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=21.46 //y=4.7 //x2=21.46 //y2=4.79
r1256 (  360 361 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.76 //y=2.08 //x2=17.76 //y2=1.915
r1257 (  353 354 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r1258 (  351 353 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r1259 (  344 438 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=79.315 //y=4.79 //x2=79.18 //y2=4.79
r1260 (  343 345 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=79.515 //y=4.79 //x2=79.59 //y2=4.865
r1261 (  343 344 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=79.515 //y=4.79 //x2=79.315 //y2=4.79
r1262 (  342 443 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=79.27 //y=1.915 //x2=79.195 //y2=2.08
r1263 (  341 441 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=79.27 //y=1.45 //x2=79.23 //y2=1.375
r1264 (  341 342 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=79.27 //y=1.45 //x2=79.27 //y2=1.915
r1265 (  340 441 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.27 //y=1.22 //x2=79.23 //y2=1.375
r1266 (  339 440 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.27 //y=0.91 //x2=79.23 //y2=0.755
r1267 (  339 340 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=79.27 //y=0.91 //x2=79.27 //y2=1.22
r1268 (  334 434 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.9 //y=1.375 //x2=78.785 //y2=1.375
r1269 (  333 441 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=79.115 //y=1.375 //x2=79.23 //y2=1.375
r1270 (  332 433 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.9 //y=0.755 //x2=78.785 //y2=0.755
r1271 (  331 440 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=79.115 //y=0.755 //x2=79.23 //y2=0.755
r1272 (  331 332 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=79.115 //y=0.755 //x2=78.9 //y2=0.755
r1273 (  330 434 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.745 //y=1.22 //x2=78.785 //y2=1.375
r1274 (  329 433 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.745 //y=0.91 //x2=78.785 //y2=0.755
r1275 (  329 330 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=78.745 //y=0.91 //x2=78.745 //y2=1.22
r1276 (  328 432 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=76 //y=1.26 //x2=75.96 //y2=1.415
r1277 (  327 431 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=76 //y=0.915 //x2=75.96 //y2=0.76
r1278 (  327 328 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=76 //y=0.915 //x2=76 //y2=1.26
r1279 (  325 428 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.625 //y=1.415 //x2=75.51 //y2=1.415
r1280 (  324 432 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.845 //y=1.415 //x2=75.96 //y2=1.415
r1281 (  323 427 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.625 //y=0.76 //x2=75.51 //y2=0.76
r1282 (  322 431 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.845 //y=0.76 //x2=75.96 //y2=0.76
r1283 (  322 323 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=75.845 //y=0.76 //x2=75.625 //y2=0.76
r1284 (  319 430 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=75.66 //y=4.865 //x2=75.48 //y2=4.7
r1285 (  317 428 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.47 //y=1.57 //x2=75.51 //y2=1.415
r1286 (  317 425 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.47 //y=1.57 //x2=75.47 //y2=1.915
r1287 (  316 428 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.47 //y=1.26 //x2=75.51 //y2=1.415
r1288 (  315 427 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.47 //y=0.915 //x2=75.51 //y2=0.76
r1289 (  315 316 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.47 //y=0.915 //x2=75.47 //y2=1.26
r1290 (  312 430 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=75.22 //y=4.865 //x2=75.48 //y2=4.7
r1291 (  308 417 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=60.075 //y=4.79 //x2=59.94 //y2=4.79
r1292 (  307 309 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=60.275 //y=4.79 //x2=60.35 //y2=4.865
r1293 (  307 308 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=60.275 //y=4.79 //x2=60.075 //y2=4.79
r1294 (  306 422 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=60.03 //y=1.915 //x2=59.955 //y2=2.08
r1295 (  305 420 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=60.03 //y=1.45 //x2=59.99 //y2=1.375
r1296 (  305 306 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=60.03 //y=1.45 //x2=60.03 //y2=1.915
r1297 (  304 420 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.03 //y=1.22 //x2=59.99 //y2=1.375
r1298 (  303 419 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.03 //y=0.91 //x2=59.99 //y2=0.755
r1299 (  303 304 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=60.03 //y=0.91 //x2=60.03 //y2=1.22
r1300 (  298 413 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.66 //y=1.375 //x2=59.545 //y2=1.375
r1301 (  297 420 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.875 //y=1.375 //x2=59.99 //y2=1.375
r1302 (  296 412 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.66 //y=0.755 //x2=59.545 //y2=0.755
r1303 (  295 419 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.875 //y=0.755 //x2=59.99 //y2=0.755
r1304 (  295 296 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=59.875 //y=0.755 //x2=59.66 //y2=0.755
r1305 (  294 413 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.505 //y=1.22 //x2=59.545 //y2=1.375
r1306 (  293 412 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.505 //y=0.91 //x2=59.545 //y2=0.755
r1307 (  293 294 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=59.505 //y=0.91 //x2=59.505 //y2=1.22
r1308 (  289 406 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=50.455 //y=4.79 //x2=50.32 //y2=4.79
r1309 (  288 290 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=50.655 //y=4.79 //x2=50.73 //y2=4.865
r1310 (  288 289 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=50.655 //y=4.79 //x2=50.455 //y2=4.79
r1311 (  287 411 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=50.41 //y=1.915 //x2=50.335 //y2=2.08
r1312 (  286 409 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=50.41 //y=1.45 //x2=50.37 //y2=1.375
r1313 (  286 287 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=50.41 //y=1.45 //x2=50.41 //y2=1.915
r1314 (  285 409 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.41 //y=1.22 //x2=50.37 //y2=1.375
r1315 (  284 408 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.41 //y=0.91 //x2=50.37 //y2=0.755
r1316 (  284 285 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=50.41 //y=0.91 //x2=50.41 //y2=1.22
r1317 (  279 402 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.04 //y=1.375 //x2=49.925 //y2=1.375
r1318 (  278 409 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.255 //y=1.375 //x2=50.37 //y2=1.375
r1319 (  277 401 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.04 //y=0.755 //x2=49.925 //y2=0.755
r1320 (  276 408 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.255 //y=0.755 //x2=50.37 //y2=0.755
r1321 (  276 277 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=50.255 //y=0.755 //x2=50.04 //y2=0.755
r1322 (  275 402 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.885 //y=1.22 //x2=49.925 //y2=1.375
r1323 (  274 401 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.885 //y=0.91 //x2=49.925 //y2=0.755
r1324 (  274 275 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=49.885 //y=0.91 //x2=49.885 //y2=1.22
r1325 (  273 400 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.14 //y=1.26 //x2=47.1 //y2=1.415
r1326 (  272 399 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.14 //y=0.915 //x2=47.1 //y2=0.76
r1327 (  272 273 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=47.14 //y=0.915 //x2=47.14 //y2=1.26
r1328 (  270 396 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.765 //y=1.415 //x2=46.65 //y2=1.415
r1329 (  269 400 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.985 //y=1.415 //x2=47.1 //y2=1.415
r1330 (  268 395 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.765 //y=0.76 //x2=46.65 //y2=0.76
r1331 (  267 399 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.985 //y=0.76 //x2=47.1 //y2=0.76
r1332 (  267 268 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=46.985 //y=0.76 //x2=46.765 //y2=0.76
r1333 (  264 398 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=46.8 //y=4.865 //x2=46.62 //y2=4.7
r1334 (  262 396 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.61 //y=1.57 //x2=46.65 //y2=1.415
r1335 (  262 393 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=46.61 //y=1.57 //x2=46.61 //y2=1.915
r1336 (  261 396 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.61 //y=1.26 //x2=46.65 //y2=1.415
r1337 (  260 395 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.61 //y=0.915 //x2=46.65 //y2=0.76
r1338 (  260 261 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=46.61 //y=0.915 //x2=46.61 //y2=1.26
r1339 (  257 398 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=46.36 //y=4.865 //x2=46.62 //y2=4.7
r1340 (  253 385 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=31.215 //y=4.79 //x2=31.08 //y2=4.79
r1341 (  252 254 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=31.415 //y=4.79 //x2=31.49 //y2=4.865
r1342 (  252 253 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=31.415 //y=4.79 //x2=31.215 //y2=4.79
r1343 (  251 390 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=31.17 //y=1.915 //x2=31.095 //y2=2.08
r1344 (  250 388 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=31.17 //y=1.45 //x2=31.13 //y2=1.375
r1345 (  250 251 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=31.17 //y=1.45 //x2=31.17 //y2=1.915
r1346 (  249 388 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.17 //y=1.22 //x2=31.13 //y2=1.375
r1347 (  248 387 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.17 //y=0.91 //x2=31.13 //y2=0.755
r1348 (  248 249 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=31.17 //y=0.91 //x2=31.17 //y2=1.22
r1349 (  243 381 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.8 //y=1.375 //x2=30.685 //y2=1.375
r1350 (  242 388 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.015 //y=1.375 //x2=31.13 //y2=1.375
r1351 (  241 380 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.8 //y=0.755 //x2=30.685 //y2=0.755
r1352 (  240 387 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.015 //y=0.755 //x2=31.13 //y2=0.755
r1353 (  240 241 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=31.015 //y=0.755 //x2=30.8 //y2=0.755
r1354 (  239 381 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.645 //y=1.22 //x2=30.685 //y2=1.375
r1355 (  238 380 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.645 //y=0.91 //x2=30.685 //y2=0.755
r1356 (  238 239 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=30.645 //y=0.91 //x2=30.645 //y2=1.22
r1357 (  234 374 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=21.595 //y=4.79 //x2=21.46 //y2=4.79
r1358 (  233 235 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.795 //y=4.79 //x2=21.87 //y2=4.865
r1359 (  233 234 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=21.795 //y=4.79 //x2=21.595 //y2=4.79
r1360 (  232 379 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.915 //x2=21.475 //y2=2.08
r1361 (  231 377 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.45 //x2=21.51 //y2=1.375
r1362 (  231 232 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.45 //x2=21.55 //y2=1.915
r1363 (  230 377 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.22 //x2=21.51 //y2=1.375
r1364 (  229 376 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.91 //x2=21.51 //y2=0.755
r1365 (  229 230 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.91 //x2=21.55 //y2=1.22
r1366 (  224 370 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.18 //y=1.375 //x2=21.065 //y2=1.375
r1367 (  223 377 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.395 //y=1.375 //x2=21.51 //y2=1.375
r1368 (  222 369 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.18 //y=0.755 //x2=21.065 //y2=0.755
r1369 (  221 376 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.755 //x2=21.51 //y2=0.755
r1370 (  221 222 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.755 //x2=21.18 //y2=0.755
r1371 (  220 370 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.025 //y=1.22 //x2=21.065 //y2=1.375
r1372 (  219 369 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.025 //y=0.91 //x2=21.065 //y2=0.755
r1373 (  219 220 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.025 //y=0.91 //x2=21.025 //y2=1.22
r1374 (  218 368 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.28 //y=1.26 //x2=18.24 //y2=1.415
r1375 (  217 367 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.28 //y=0.915 //x2=18.24 //y2=0.76
r1376 (  217 218 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.28 //y=0.915 //x2=18.28 //y2=1.26
r1377 (  215 364 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.905 //y=1.415 //x2=17.79 //y2=1.415
r1378 (  214 368 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.125 //y=1.415 //x2=18.24 //y2=1.415
r1379 (  213 363 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.905 //y=0.76 //x2=17.79 //y2=0.76
r1380 (  212 367 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.125 //y=0.76 //x2=18.24 //y2=0.76
r1381 (  212 213 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.125 //y=0.76 //x2=17.905 //y2=0.76
r1382 (  209 366 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=17.94 //y=4.865 //x2=17.76 //y2=4.7
r1383 (  207 364 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.57 //x2=17.79 //y2=1.415
r1384 (  207 361 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.57 //x2=17.75 //y2=1.915
r1385 (  206 364 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.26 //x2=17.79 //y2=1.415
r1386 (  205 363 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=0.915 //x2=17.79 //y2=0.76
r1387 (  205 206 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.75 //y=0.915 //x2=17.75 //y2=1.26
r1388 (  202 366 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=17.5 //y=4.865 //x2=17.76 //y2=4.7
r1389 (  198 353 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r1390 (  197 199 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r1391 (  197 198 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r1392 (  196 358 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r1393 (  195 356 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r1394 (  195 196 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r1395 (  194 356 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r1396 (  193 355 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r1397 (  193 194 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r1398 (  188 349 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r1399 (  187 356 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r1400 (  186 348 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r1401 (  185 355 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r1402 (  185 186 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r1403 (  184 349 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r1404 (  183 348 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r1405 (  183 184 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r1406 (  182 345 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=79.59 //y=6.02 //x2=79.59 //y2=4.865
r1407 (  181 439 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=79.15 //y=6.02 //x2=79.15 //y2=4.865
r1408 (  180 319 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.66 //y=6.02 //x2=75.66 //y2=4.865
r1409 (  179 312 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.22 //y=6.02 //x2=75.22 //y2=4.865
r1410 (  178 309 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.35 //y=6.02 //x2=60.35 //y2=4.865
r1411 (  177 418 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.91 //y=6.02 //x2=59.91 //y2=4.865
r1412 (  176 290 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.73 //y=6.02 //x2=50.73 //y2=4.865
r1413 (  175 407 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.29 //y=6.02 //x2=50.29 //y2=4.865
r1414 (  174 264 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.8 //y=6.02 //x2=46.8 //y2=4.865
r1415 (  173 257 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.36 //y=6.02 //x2=46.36 //y2=4.865
r1416 (  172 254 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.49 //y=6.02 //x2=31.49 //y2=4.865
r1417 (  171 386 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.05 //y=6.02 //x2=31.05 //y2=4.865
r1418 (  170 235 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.87 //y=6.02 //x2=21.87 //y2=4.865
r1419 (  169 375 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.43 //y=6.02 //x2=21.43 //y2=4.865
r1420 (  168 209 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.94 //y=6.02 //x2=17.94 //y2=4.865
r1421 (  167 202 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.5 //y=6.02 //x2=17.5 //y2=4.865
r1422 (  166 199 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r1423 (  165 354 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r1424 (  164 333 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=79.007 //y=1.375 //x2=79.115 //y2=1.375
r1425 (  164 334 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=79.007 //y=1.375 //x2=78.9 //y2=1.375
r1426 (  163 324 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.735 //y=1.415 //x2=75.845 //y2=1.415
r1427 (  163 325 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.735 //y=1.415 //x2=75.625 //y2=1.415
r1428 (  162 297 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=59.767 //y=1.375 //x2=59.875 //y2=1.375
r1429 (  162 298 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=59.767 //y=1.375 //x2=59.66 //y2=1.375
r1430 (  161 278 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=50.147 //y=1.375 //x2=50.255 //y2=1.375
r1431 (  161 279 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=50.147 //y=1.375 //x2=50.04 //y2=1.375
r1432 (  160 269 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=46.875 //y=1.415 //x2=46.985 //y2=1.415
r1433 (  160 270 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=46.875 //y=1.415 //x2=46.765 //y2=1.415
r1434 (  159 242 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=30.907 //y=1.375 //x2=31.015 //y2=1.375
r1435 (  159 243 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=30.907 //y=1.375 //x2=30.8 //y2=1.375
r1436 (  158 223 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=21.287 //y=1.375 //x2=21.395 //y2=1.375
r1437 (  158 224 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=21.287 //y=1.375 //x2=21.18 //y2=1.375
r1438 (  157 214 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.015 //y=1.415 //x2=18.125 //y2=1.415
r1439 (  157 215 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.015 //y=1.415 //x2=17.905 //y2=1.415
r1440 (  156 187 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r1441 (  156 188 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r1442 (  154 436 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.18 //y=4.7 //x2=79.18 //y2=4.7
r1443 (  147 443 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.18 //y=2.08 //x2=79.18 //y2=2.08
r1444 (  144 430 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.48 //y=4.7 //x2=75.48 //y2=4.7
r1445 (  138 424 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.48 //y=2.08 //x2=75.48 //y2=2.08
r1446 (  135 415 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.94 //y=4.7 //x2=59.94 //y2=4.7
r1447 (  127 422 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.94 //y=2.08 //x2=59.94 //y2=2.08
r1448 (  124 404 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.32 //y=4.7 //x2=50.32 //y2=4.7
r1449 (  117 411 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.32 //y=2.08 //x2=50.32 //y2=2.08
r1450 (  114 398 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.62 //y=4.7 //x2=46.62 //y2=4.7
r1451 (  108 392 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.62 //y=2.08 //x2=46.62 //y2=2.08
r1452 (  105 383 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.08 //y=4.7 //x2=31.08 //y2=4.7
r1453 (  97 390 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.08 //y=2.08 //x2=31.08 //y2=2.08
r1454 (  94 372 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=4.7 //x2=21.46 //y2=4.7
r1455 (  87 379 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=2.08 //x2=21.46 //y2=2.08
r1456 (  84 366 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=4.7 //x2=17.76 //y2=4.7
r1457 (  78 360 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=2.08 //x2=17.76 //y2=2.08
r1458 (  75 351 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r1459 (  65 358 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r1460 (  63 154 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=79.18 //y=3.33 //x2=79.18 //y2=4.7
r1461 (  62 63 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=79.18 //y=2.59 //x2=79.18 //y2=3.33
r1462 (  61 62 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=79.18 //y=2.22 //x2=79.18 //y2=2.59
r1463 (  61 147 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=79.18 //y=2.22 //x2=79.18 //y2=2.08
r1464 (  60 144 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=75.48 //y=2.59 //x2=75.48 //y2=4.7
r1465 (  59 60 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=75.48 //y=2.22 //x2=75.48 //y2=2.59
r1466 (  59 138 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=75.48 //y=2.22 //x2=75.48 //y2=2.08
r1467 (  58 135 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=59.94 //y=4.07 //x2=59.94 //y2=4.7
r1468 (  57 58 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=59.94 //y=3.33 //x2=59.94 //y2=4.07
r1469 (  56 57 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=59.94 //y=2.59 //x2=59.94 //y2=3.33
r1470 (  55 56 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=59.94 //y=2.22 //x2=59.94 //y2=2.59
r1471 (  55 127 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=59.94 //y=2.22 //x2=59.94 //y2=2.08
r1472 (  54 124 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=50.32 //y=3.33 //x2=50.32 //y2=4.7
r1473 (  53 54 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=50.32 //y=2.59 //x2=50.32 //y2=3.33
r1474 (  52 53 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=50.32 //y=2.22 //x2=50.32 //y2=2.59
r1475 (  52 117 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=50.32 //y=2.22 //x2=50.32 //y2=2.08
r1476 (  51 114 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=46.62 //y=2.59 //x2=46.62 //y2=4.7
r1477 (  50 51 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=46.62 //y=2.22 //x2=46.62 //y2=2.59
r1478 (  50 108 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=46.62 //y=2.22 //x2=46.62 //y2=2.08
r1479 (  49 105 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li \
 //thickness=0.1 //x=31.08 //y=3.7 //x2=31.08 //y2=4.7
r1480 (  48 49 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=31.08 //y=3.33 //x2=31.08 //y2=3.7
r1481 (  47 48 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=31.08 //y=2.59 //x2=31.08 //y2=3.33
r1482 (  46 47 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=31.08 //y=2.22 //x2=31.08 //y2=2.59
r1483 (  46 97 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=31.08 //y=2.22 //x2=31.08 //y2=2.08
r1484 (  45 94 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=3.33 //x2=21.46 //y2=4.7
r1485 (  44 45 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.59 //x2=21.46 //y2=3.33
r1486 (  43 44 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.22 //x2=21.46 //y2=2.59
r1487 (  43 87 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.22 //x2=21.46 //y2=2.08
r1488 (  42 84 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.59 //x2=17.76 //y2=4.7
r1489 (  41 42 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.22 //x2=17.76 //y2=2.59
r1490 (  41 78 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.22 //x2=17.76 //y2=2.08
r1491 (  40 75 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=2.22 //y=4.44 //x2=2.22 //y2=4.7
r1492 (  39 40 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.7 //x2=2.22 //y2=4.44
r1493 (  38 39 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.33 //x2=2.22 //y2=3.7
r1494 (  37 38 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.96 //x2=2.22 //y2=3.33
r1495 (  36 37 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.59 //x2=2.22 //y2=2.96
r1496 (  35 36 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.22 //x2=2.22 //y2=2.59
r1497 (  35 65 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.22 //x2=2.22 //y2=2.08
r1498 (  34 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.18 //y=2.22 //x2=79.18 //y2=2.22
r1499 (  32 59 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.48 //y=2.22 //x2=75.48 //y2=2.22
r1500 (  30 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=59.94 //y=2.22 //x2=59.94 //y2=2.22
r1501 (  28 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=50.32 //y=2.22 //x2=50.32 //y2=2.22
r1502 (  26 50 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=46.62 //y=2.22 //x2=46.62 //y2=2.22
r1503 (  24 46 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=31.08 //y=2.22 //x2=31.08 //y2=2.22
r1504 (  22 43 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.46 //y=2.22 //x2=21.46 //y2=2.22
r1505 (  20 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.76 //y=2.22 //x2=17.76 //y2=2.22
r1506 (  18 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.22 //y=2.22 //x2=2.22 //y2=2.22
r1507 (  16 32 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.595 //y=2.22 //x2=75.48 //y2=2.22
r1508 (  15 34 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.065 //y=2.22 //x2=79.18 //y2=2.22
r1509 (  15 16 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=79.065 //y=2.22 //x2=75.595 //y2=2.22
r1510 (  14 30 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.055 //y=2.22 //x2=59.94 //y2=2.22
r1511 (  13 32 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.365 //y=2.22 //x2=75.48 //y2=2.22
r1512 (  13 14 ) resistor r=14.6088 //w=0.131 //l=15.31 //layer=m1 \
 //thickness=0.36 //x=75.365 //y=2.22 //x2=60.055 //y2=2.22
r1513 (  12 28 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.435 //y=2.22 //x2=50.32 //y2=2.22
r1514 (  11 30 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=59.825 //y=2.22 //x2=59.94 //y2=2.22
r1515 (  11 12 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=59.825 //y=2.22 //x2=50.435 //y2=2.22
r1516 (  10 26 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=46.735 //y=2.22 //x2=46.62 //y2=2.22
r1517 (  9 28 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.205 //y=2.22 //x2=50.32 //y2=2.22
r1518 (  9 10 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=50.205 //y=2.22 //x2=46.735 //y2=2.22
r1519 (  8 24 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.195 //y=2.22 //x2=31.08 //y2=2.22
r1520 (  7 26 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=46.505 //y=2.22 //x2=46.62 //y2=2.22
r1521 (  7 8 ) resistor r=14.6088 //w=0.131 //l=15.31 //layer=m1 \
 //thickness=0.36 //x=46.505 //y=2.22 //x2=31.195 //y2=2.22
r1522 (  6 22 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.575 //y=2.22 //x2=21.46 //y2=2.22
r1523 (  5 24 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=30.965 //y=2.22 //x2=31.08 //y2=2.22
r1524 (  5 6 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=30.965 //y=2.22 //x2=21.575 //y2=2.22
r1525 (  4 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.875 //y=2.22 //x2=17.76 //y2=2.22
r1526 (  3 22 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=2.22 //x2=21.46 //y2=2.22
r1527 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=2.22 //x2=17.875 //y2=2.22
r1528 (  2 18 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.335 //y=2.22 //x2=2.22 //y2=2.22
r1529 (  1 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.645 //y=2.22 //x2=17.76 //y2=2.22
r1530 (  1 2 ) resistor r=14.6088 //w=0.131 //l=15.31 //layer=m1 \
 //thickness=0.36 //x=17.645 //y=2.22 //x2=2.335 //y2=2.22
ends PM_TMRDFFSNRNQX1\%RN

subckt PM_TMRDFFSNRNQX1\%noxref_21 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 \
 53 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c161 ( 85 0 ) capacitor c=0.023087f //x=80.105 //y=5.02
c162 ( 84 0 ) capacitor c=0.023519f //x=79.225 //y=5.02
c163 ( 83 0 ) capacitor c=0.0224735f //x=78.345 //y=5.02
c164 ( 81 0 ) capacitor c=0.00853354f //x=80.355 //y=0.915
c165 ( 69 0 ) capacitor c=0.0556143f //x=83.155 //y=4.79
c166 ( 68 0 ) capacitor c=0.0293157f //x=83.445 //y=4.79
c167 ( 67 0 ) capacitor c=0.0347816f //x=83.11 //y=1.22
c168 ( 66 0 ) capacitor c=0.0187487f //x=83.11 //y=0.875
c169 ( 60 0 ) capacitor c=0.0137055f //x=82.955 //y=1.375
c170 ( 58 0 ) capacitor c=0.0149861f //x=82.955 //y=0.72
c171 ( 57 0 ) capacitor c=0.096037f //x=82.58 //y=1.915
c172 ( 56 0 ) capacitor c=0.0228993f //x=82.58 //y=1.53
c173 ( 55 0 ) capacitor c=0.0234352f //x=82.58 //y=1.22
c174 ( 54 0 ) capacitor c=0.0198724f //x=82.58 //y=0.875
c175 ( 53 0 ) capacitor c=0.110114f //x=83.52 //y=6.02
c176 ( 52 0 ) capacitor c=0.158956f //x=83.08 //y=6.02
c177 ( 50 0 ) capacitor c=0.00106608f //x=80.25 //y=5.155
c178 ( 49 0 ) capacitor c=0.00207319f //x=79.37 //y=5.155
c179 ( 42 0 ) capacitor c=0.0971623f //x=82.88 //y=2.08
c180 ( 40 0 ) capacitor c=0.106761f //x=81.03 //y=2.59
c181 ( 36 0 ) capacitor c=0.00398962f //x=80.63 //y=1.665
c182 ( 35 0 ) capacitor c=0.0137288f //x=80.945 //y=1.665
c183 ( 29 0 ) capacitor c=0.0283082f //x=80.945 //y=5.155
c184 ( 21 0 ) capacitor c=0.0176454f //x=80.165 //y=5.155
c185 ( 14 0 ) capacitor c=0.00332903f //x=78.575 //y=5.155
c186 ( 13 0 ) capacitor c=0.0148427f //x=79.285 //y=5.155
c187 ( 2 0 ) capacitor c=0.0116088f //x=81.145 //y=2.59
c188 ( 1 0 ) capacitor c=0.0352679f //x=82.765 //y=2.59
r189 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=83.445 //y=4.79 //x2=83.52 //y2=4.865
r190 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=83.445 //y=4.79 //x2=83.155 //y2=4.79
r191 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.11 //y=1.22 //x2=83.07 //y2=1.375
r192 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.11 //y=0.875 //x2=83.07 //y2=0.72
r193 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=83.11 //y=0.875 //x2=83.11 //y2=1.22
r194 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=83.08 //y=4.865 //x2=83.155 //y2=4.79
r195 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=83.08 //y=4.865 //x2=82.88 //y2=4.7
r196 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.735 //y=1.375 //x2=82.62 //y2=1.375
r197 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.955 //y=1.375 //x2=83.07 //y2=1.375
r198 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.735 //y=0.72 //x2=82.62 //y2=0.72
r199 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.955 //y=0.72 //x2=83.07 //y2=0.72
r200 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=82.955 //y=0.72 //x2=82.735 //y2=0.72
r201 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=82.58 //y=1.915 //x2=82.88 //y2=2.08
r202 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.58 //y=1.53 //x2=82.62 //y2=1.375
r203 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=82.58 //y=1.53 //x2=82.58 //y2=1.915
r204 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.58 //y=1.22 //x2=82.62 //y2=1.375
r205 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.58 //y=0.875 //x2=82.62 //y2=0.72
r206 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=82.58 //y=0.875 //x2=82.58 //y2=1.22
r207 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=83.52 //y=6.02 //x2=83.52 //y2=4.865
r208 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=83.08 //y=6.02 //x2=83.08 //y2=4.865
r209 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.845 //y=1.375 //x2=82.955 //y2=1.375
r210 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.845 //y=1.375 //x2=82.735 //y2=1.375
r211 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=82.88 //y=4.7 //x2=82.88 //y2=4.7
r212 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=82.88 //y=2.59 //x2=82.88 //y2=4.7
r213 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=82.88 //y=2.08 //x2=82.88 //y2=2.08
r214 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=82.88 //y=2.08 //x2=82.88 //y2=2.59
r215 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=81.03 //y=5.07 //x2=81.03 //y2=2.59
r216 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=81.03 //y=1.75 //x2=81.03 //y2=2.59
r217 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=80.945 //y=1.665 //x2=81.03 //y2=1.75
r218 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=80.945 //y=1.665 //x2=80.63 //y2=1.665
r219 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=80.545 //y=1.58 //x2=80.63 //y2=1.665
r220 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=80.545 //y=1.58 //x2=80.545 //y2=1.01
r221 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.335 //y=5.155 //x2=80.25 //y2=5.155
r222 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=80.945 //y=5.155 //x2=81.03 //y2=5.07
r223 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=80.945 //y=5.155 //x2=80.335 //y2=5.155
r224 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.25 //y=5.24 //x2=80.25 //y2=5.155
r225 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=80.25 //y=5.24 //x2=80.25 //y2=5.725
r226 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.455 //y=5.155 //x2=79.37 //y2=5.155
r227 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.165 //y=5.155 //x2=80.25 //y2=5.155
r228 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=80.165 //y=5.155 //x2=79.455 //y2=5.155
r229 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.37 //y=5.24 //x2=79.37 //y2=5.155
r230 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=79.37 //y=5.24 //x2=79.37 //y2=5.725
r231 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.285 //y=5.155 //x2=79.37 //y2=5.155
r232 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=79.285 //y=5.155 //x2=78.575 //y2=5.155
r233 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=78.49 //y=5.24 //x2=78.575 //y2=5.155
r234 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=78.49 //y=5.24 //x2=78.49 //y2=5.725
r235 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=82.88 //y=2.59 //x2=82.88 //y2=2.59
r236 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=81.03 //y=2.59 //x2=81.03 //y2=2.59
r237 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=81.145 //y=2.59 //x2=81.03 //y2=2.59
r238 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=82.765 //y=2.59 //x2=82.88 //y2=2.59
r239 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=82.765 //y=2.59 //x2=81.145 //y2=2.59
ends PM_TMRDFFSNRNQX1\%noxref_21

subckt PM_TMRDFFSNRNQX1\%SN ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 31 \
 32 34 43 52 61 70 79 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 \
 103 104 105 106 108 114 115 116 117 118 123 124 125 127 133 134 135 136 137 \
 142 143 144 146 152 153 154 155 156 161 162 163 165 171 172 173 174 175 180 \
 181 182 184 190 191 192 193 194 199 200 201 203 209 210 211 212 213 221 232 \
 243 254 265 276 )
c687 ( 276 0 ) capacitor c=0.0335551f //x=83.99 //y=4.7
c688 ( 265 0 ) capacitor c=0.0333886f //x=69.56 //y=4.7
c689 ( 254 0 ) capacitor c=0.0333886f //x=55.13 //y=4.7
c690 ( 243 0 ) capacitor c=0.0333886f //x=40.7 //y=4.7
c691 ( 232 0 ) capacitor c=0.0335551f //x=26.27 //y=4.7
c692 ( 221 0 ) capacitor c=0.0335551f //x=11.84 //y=4.7
c693 ( 213 0 ) capacitor c=0.0245352f //x=84.325 //y=4.79
c694 ( 212 0 ) capacitor c=0.0825763f //x=84.08 //y=1.915
c695 ( 211 0 ) capacitor c=0.0170266f //x=84.08 //y=1.45
c696 ( 210 0 ) capacitor c=0.018609f //x=84.08 //y=1.22
c697 ( 209 0 ) capacitor c=0.0187309f //x=84.08 //y=0.91
c698 ( 203 0 ) capacitor c=0.014725f //x=83.925 //y=1.375
c699 ( 201 0 ) capacitor c=0.0146567f //x=83.925 //y=0.755
c700 ( 200 0 ) capacitor c=0.0335408f //x=83.555 //y=1.22
c701 ( 199 0 ) capacitor c=0.0173761f //x=83.555 //y=0.91
c702 ( 194 0 ) capacitor c=0.0246783f //x=69.895 //y=4.79
c703 ( 193 0 ) capacitor c=0.0825763f //x=69.65 //y=1.915
c704 ( 192 0 ) capacitor c=0.0170266f //x=69.65 //y=1.45
c705 ( 191 0 ) capacitor c=0.018609f //x=69.65 //y=1.22
c706 ( 190 0 ) capacitor c=0.0187309f //x=69.65 //y=0.91
c707 ( 184 0 ) capacitor c=0.014725f //x=69.495 //y=1.375
c708 ( 182 0 ) capacitor c=0.0146567f //x=69.495 //y=0.755
c709 ( 181 0 ) capacitor c=0.0335408f //x=69.125 //y=1.22
c710 ( 180 0 ) capacitor c=0.0173761f //x=69.125 //y=0.91
c711 ( 175 0 ) capacitor c=0.0246783f //x=55.465 //y=4.79
c712 ( 174 0 ) capacitor c=0.0825763f //x=55.22 //y=1.915
c713 ( 173 0 ) capacitor c=0.0170266f //x=55.22 //y=1.45
c714 ( 172 0 ) capacitor c=0.018609f //x=55.22 //y=1.22
c715 ( 171 0 ) capacitor c=0.0187309f //x=55.22 //y=0.91
c716 ( 165 0 ) capacitor c=0.014725f //x=55.065 //y=1.375
c717 ( 163 0 ) capacitor c=0.0146567f //x=55.065 //y=0.755
c718 ( 162 0 ) capacitor c=0.0335408f //x=54.695 //y=1.22
c719 ( 161 0 ) capacitor c=0.0173761f //x=54.695 //y=0.91
c720 ( 156 0 ) capacitor c=0.0246783f //x=41.035 //y=4.79
c721 ( 155 0 ) capacitor c=0.0825763f //x=40.79 //y=1.915
c722 ( 154 0 ) capacitor c=0.0170266f //x=40.79 //y=1.45
c723 ( 153 0 ) capacitor c=0.018609f //x=40.79 //y=1.22
c724 ( 152 0 ) capacitor c=0.0187309f //x=40.79 //y=0.91
c725 ( 146 0 ) capacitor c=0.014725f //x=40.635 //y=1.375
c726 ( 144 0 ) capacitor c=0.0146567f //x=40.635 //y=0.755
c727 ( 143 0 ) capacitor c=0.0335408f //x=40.265 //y=1.22
c728 ( 142 0 ) capacitor c=0.0173761f //x=40.265 //y=0.91
c729 ( 137 0 ) capacitor c=0.0245352f //x=26.605 //y=4.79
c730 ( 136 0 ) capacitor c=0.0825763f //x=26.36 //y=1.915
c731 ( 135 0 ) capacitor c=0.0170266f //x=26.36 //y=1.45
c732 ( 134 0 ) capacitor c=0.018609f //x=26.36 //y=1.22
c733 ( 133 0 ) capacitor c=0.0187309f //x=26.36 //y=0.91
c734 ( 127 0 ) capacitor c=0.014725f //x=26.205 //y=1.375
c735 ( 125 0 ) capacitor c=0.0146567f //x=26.205 //y=0.755
c736 ( 124 0 ) capacitor c=0.0335408f //x=25.835 //y=1.22
c737 ( 123 0 ) capacitor c=0.0173761f //x=25.835 //y=0.91
c738 ( 118 0 ) capacitor c=0.0245352f //x=12.175 //y=4.79
c739 ( 117 0 ) capacitor c=0.0825763f //x=11.93 //y=1.915
c740 ( 116 0 ) capacitor c=0.0170266f //x=11.93 //y=1.45
c741 ( 115 0 ) capacitor c=0.018609f //x=11.93 //y=1.22
c742 ( 114 0 ) capacitor c=0.0187309f //x=11.93 //y=0.91
c743 ( 108 0 ) capacitor c=0.014725f //x=11.775 //y=1.375
c744 ( 106 0 ) capacitor c=0.0146567f //x=11.775 //y=0.755
c745 ( 105 0 ) capacitor c=0.0335408f //x=11.405 //y=1.22
c746 ( 104 0 ) capacitor c=0.0173761f //x=11.405 //y=0.91
c747 ( 103 0 ) capacitor c=0.110114f //x=84.4 //y=6.02
c748 ( 102 0 ) capacitor c=0.11012f //x=83.96 //y=6.02
c749 ( 101 0 ) capacitor c=0.109949f //x=69.97 //y=6.02
c750 ( 100 0 ) capacitor c=0.109956f //x=69.53 //y=6.02
c751 ( 99 0 ) capacitor c=0.109949f //x=55.54 //y=6.02
c752 ( 98 0 ) capacitor c=0.109956f //x=55.1 //y=6.02
c753 ( 97 0 ) capacitor c=0.109949f //x=41.11 //y=6.02
c754 ( 96 0 ) capacitor c=0.109956f //x=40.67 //y=6.02
c755 ( 95 0 ) capacitor c=0.110114f //x=26.68 //y=6.02
c756 ( 94 0 ) capacitor c=0.11012f //x=26.24 //y=6.02
c757 ( 93 0 ) capacitor c=0.110114f //x=12.25 //y=6.02
c758 ( 92 0 ) capacitor c=0.11012f //x=11.81 //y=6.02
c759 ( 79 0 ) capacitor c=0.0925663f //x=83.99 //y=2.08
c760 ( 70 0 ) capacitor c=0.0877968f //x=69.56 //y=2.08
c761 ( 61 0 ) capacitor c=0.0881699f //x=55.13 //y=2.08
c762 ( 52 0 ) capacitor c=0.0877968f //x=40.7 //y=2.08
c763 ( 43 0 ) capacitor c=0.089887f //x=26.27 //y=2.08
c764 ( 34 0 ) capacitor c=0.0895139f //x=11.84 //y=2.08
c765 ( 10 0 ) capacitor c=0.00568147f //x=69.675 //y=2.96
c766 ( 9 0 ) capacitor c=0.267214f //x=83.875 //y=2.96
c767 ( 8 0 ) capacitor c=0.00568147f //x=55.245 //y=2.96
c768 ( 7 0 ) capacitor c=0.231482f //x=69.445 //y=2.96
c769 ( 6 0 ) capacitor c=0.00568147f //x=40.815 //y=2.96
c770 ( 5 0 ) capacitor c=0.230801f //x=55.015 //y=2.96
c771 ( 4 0 ) capacitor c=0.00579855f //x=26.385 //y=2.96
c772 ( 3 0 ) capacitor c=0.242173f //x=40.585 //y=2.96
c773 ( 2 0 ) capacitor c=0.0141295f //x=11.955 //y=2.96
c774 ( 1 0 ) capacitor c=0.231794f //x=26.155 //y=2.96
r775 (  278 279 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=83.99 //y=4.79 //x2=83.99 //y2=4.865
r776 (  276 278 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=83.99 //y=4.7 //x2=83.99 //y2=4.79
r777 (  267 268 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=69.56 //y=4.79 //x2=69.56 //y2=4.865
r778 (  265 267 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=69.56 //y=4.7 //x2=69.56 //y2=4.79
r779 (  256 257 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=55.13 //y=4.79 //x2=55.13 //y2=4.865
r780 (  254 256 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=55.13 //y=4.7 //x2=55.13 //y2=4.79
r781 (  245 246 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=40.7 //y=4.79 //x2=40.7 //y2=4.865
r782 (  243 245 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=40.7 //y=4.7 //x2=40.7 //y2=4.79
r783 (  234 235 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=26.27 //y=4.79 //x2=26.27 //y2=4.865
r784 (  232 234 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=26.27 //y=4.7 //x2=26.27 //y2=4.79
r785 (  223 224 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=11.84 //y=4.79 //x2=11.84 //y2=4.865
r786 (  221 223 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=11.84 //y=4.7 //x2=11.84 //y2=4.79
r787 (  214 278 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=84.125 //y=4.79 //x2=83.99 //y2=4.79
r788 (  213 215 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=84.325 //y=4.79 //x2=84.4 //y2=4.865
r789 (  213 214 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=84.325 //y=4.79 //x2=84.125 //y2=4.79
r790 (  212 283 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=84.08 //y=1.915 //x2=84.005 //y2=2.08
r791 (  211 281 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=84.08 //y=1.45 //x2=84.04 //y2=1.375
r792 (  211 212 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=84.08 //y=1.45 //x2=84.08 //y2=1.915
r793 (  210 281 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=84.08 //y=1.22 //x2=84.04 //y2=1.375
r794 (  209 280 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=84.08 //y=0.91 //x2=84.04 //y2=0.755
r795 (  209 210 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=84.08 //y=0.91 //x2=84.08 //y2=1.22
r796 (  204 274 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.71 //y=1.375 //x2=83.595 //y2=1.375
r797 (  203 281 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.925 //y=1.375 //x2=84.04 //y2=1.375
r798 (  202 273 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.71 //y=0.755 //x2=83.595 //y2=0.755
r799 (  201 280 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.925 //y=0.755 //x2=84.04 //y2=0.755
r800 (  201 202 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=83.925 //y=0.755 //x2=83.71 //y2=0.755
r801 (  200 274 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.555 //y=1.22 //x2=83.595 //y2=1.375
r802 (  199 273 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.555 //y=0.91 //x2=83.595 //y2=0.755
r803 (  199 200 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=83.555 //y=0.91 //x2=83.555 //y2=1.22
r804 (  195 267 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=69.695 //y=4.79 //x2=69.56 //y2=4.79
r805 (  194 196 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=69.895 //y=4.79 //x2=69.97 //y2=4.865
r806 (  194 195 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=69.895 //y=4.79 //x2=69.695 //y2=4.79
r807 (  193 272 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=69.65 //y=1.915 //x2=69.575 //y2=2.08
r808 (  192 270 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=69.65 //y=1.45 //x2=69.61 //y2=1.375
r809 (  192 193 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=69.65 //y=1.45 //x2=69.65 //y2=1.915
r810 (  191 270 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.65 //y=1.22 //x2=69.61 //y2=1.375
r811 (  190 269 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.65 //y=0.91 //x2=69.61 //y2=0.755
r812 (  190 191 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=69.65 //y=0.91 //x2=69.65 //y2=1.22
r813 (  185 263 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.28 //y=1.375 //x2=69.165 //y2=1.375
r814 (  184 270 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.495 //y=1.375 //x2=69.61 //y2=1.375
r815 (  183 262 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.28 //y=0.755 //x2=69.165 //y2=0.755
r816 (  182 269 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.495 //y=0.755 //x2=69.61 //y2=0.755
r817 (  182 183 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=69.495 //y=0.755 //x2=69.28 //y2=0.755
r818 (  181 263 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.125 //y=1.22 //x2=69.165 //y2=1.375
r819 (  180 262 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.125 //y=0.91 //x2=69.165 //y2=0.755
r820 (  180 181 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=69.125 //y=0.91 //x2=69.125 //y2=1.22
r821 (  176 256 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=55.265 //y=4.79 //x2=55.13 //y2=4.79
r822 (  175 177 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=55.465 //y=4.79 //x2=55.54 //y2=4.865
r823 (  175 176 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=55.465 //y=4.79 //x2=55.265 //y2=4.79
r824 (  174 261 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=55.22 //y=1.915 //x2=55.145 //y2=2.08
r825 (  173 259 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=55.22 //y=1.45 //x2=55.18 //y2=1.375
r826 (  173 174 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=55.22 //y=1.45 //x2=55.22 //y2=1.915
r827 (  172 259 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.22 //y=1.22 //x2=55.18 //y2=1.375
r828 (  171 258 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.22 //y=0.91 //x2=55.18 //y2=0.755
r829 (  171 172 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=55.22 //y=0.91 //x2=55.22 //y2=1.22
r830 (  166 252 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.85 //y=1.375 //x2=54.735 //y2=1.375
r831 (  165 259 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.065 //y=1.375 //x2=55.18 //y2=1.375
r832 (  164 251 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.85 //y=0.755 //x2=54.735 //y2=0.755
r833 (  163 258 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.065 //y=0.755 //x2=55.18 //y2=0.755
r834 (  163 164 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=55.065 //y=0.755 //x2=54.85 //y2=0.755
r835 (  162 252 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.695 //y=1.22 //x2=54.735 //y2=1.375
r836 (  161 251 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.695 //y=0.91 //x2=54.735 //y2=0.755
r837 (  161 162 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=54.695 //y=0.91 //x2=54.695 //y2=1.22
r838 (  157 245 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=40.835 //y=4.79 //x2=40.7 //y2=4.79
r839 (  156 158 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=41.035 //y=4.79 //x2=41.11 //y2=4.865
r840 (  156 157 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=41.035 //y=4.79 //x2=40.835 //y2=4.79
r841 (  155 250 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=40.79 //y=1.915 //x2=40.715 //y2=2.08
r842 (  154 248 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=40.79 //y=1.45 //x2=40.75 //y2=1.375
r843 (  154 155 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=40.79 //y=1.45 //x2=40.79 //y2=1.915
r844 (  153 248 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.79 //y=1.22 //x2=40.75 //y2=1.375
r845 (  152 247 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.79 //y=0.91 //x2=40.75 //y2=0.755
r846 (  152 153 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=40.79 //y=0.91 //x2=40.79 //y2=1.22
r847 (  147 241 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.42 //y=1.375 //x2=40.305 //y2=1.375
r848 (  146 248 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.635 //y=1.375 //x2=40.75 //y2=1.375
r849 (  145 240 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.42 //y=0.755 //x2=40.305 //y2=0.755
r850 (  144 247 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.635 //y=0.755 //x2=40.75 //y2=0.755
r851 (  144 145 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=40.635 //y=0.755 //x2=40.42 //y2=0.755
r852 (  143 241 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.265 //y=1.22 //x2=40.305 //y2=1.375
r853 (  142 240 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.265 //y=0.91 //x2=40.305 //y2=0.755
r854 (  142 143 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=40.265 //y=0.91 //x2=40.265 //y2=1.22
r855 (  138 234 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=26.405 //y=4.79 //x2=26.27 //y2=4.79
r856 (  137 139 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=26.605 //y=4.79 //x2=26.68 //y2=4.865
r857 (  137 138 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=26.605 //y=4.79 //x2=26.405 //y2=4.79
r858 (  136 239 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.915 //x2=26.285 //y2=2.08
r859 (  135 237 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.45 //x2=26.32 //y2=1.375
r860 (  135 136 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.45 //x2=26.36 //y2=1.915
r861 (  134 237 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.22 //x2=26.32 //y2=1.375
r862 (  133 236 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.36 //y=0.91 //x2=26.32 //y2=0.755
r863 (  133 134 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=26.36 //y=0.91 //x2=26.36 //y2=1.22
r864 (  128 230 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.99 //y=1.375 //x2=25.875 //y2=1.375
r865 (  127 237 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.205 //y=1.375 //x2=26.32 //y2=1.375
r866 (  126 229 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.99 //y=0.755 //x2=25.875 //y2=0.755
r867 (  125 236 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.205 //y=0.755 //x2=26.32 //y2=0.755
r868 (  125 126 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=26.205 //y=0.755 //x2=25.99 //y2=0.755
r869 (  124 230 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.835 //y=1.22 //x2=25.875 //y2=1.375
r870 (  123 229 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.835 //y=0.91 //x2=25.875 //y2=0.755
r871 (  123 124 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=25.835 //y=0.91 //x2=25.835 //y2=1.22
r872 (  119 223 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=11.975 //y=4.79 //x2=11.84 //y2=4.79
r873 (  118 120 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=12.175 //y=4.79 //x2=12.25 //y2=4.865
r874 (  118 119 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=12.175 //y=4.79 //x2=11.975 //y2=4.79
r875 (  117 228 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.915 //x2=11.855 //y2=2.08
r876 (  116 226 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.45 //x2=11.89 //y2=1.375
r877 (  116 117 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.45 //x2=11.93 //y2=1.915
r878 (  115 226 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.22 //x2=11.89 //y2=1.375
r879 (  114 225 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.93 //y=0.91 //x2=11.89 //y2=0.755
r880 (  114 115 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=11.93 //y=0.91 //x2=11.93 //y2=1.22
r881 (  109 219 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.56 //y=1.375 //x2=11.445 //y2=1.375
r882 (  108 226 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.775 //y=1.375 //x2=11.89 //y2=1.375
r883 (  107 218 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.56 //y=0.755 //x2=11.445 //y2=0.755
r884 (  106 225 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.775 //y=0.755 //x2=11.89 //y2=0.755
r885 (  106 107 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=11.775 //y=0.755 //x2=11.56 //y2=0.755
r886 (  105 219 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.405 //y=1.22 //x2=11.445 //y2=1.375
r887 (  104 218 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.405 //y=0.91 //x2=11.445 //y2=0.755
r888 (  104 105 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=11.405 //y=0.91 //x2=11.405 //y2=1.22
r889 (  103 215 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=84.4 //y=6.02 //x2=84.4 //y2=4.865
r890 (  102 279 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=83.96 //y=6.02 //x2=83.96 //y2=4.865
r891 (  101 196 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.97 //y=6.02 //x2=69.97 //y2=4.865
r892 (  100 268 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.53 //y=6.02 //x2=69.53 //y2=4.865
r893 (  99 177 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.54 //y=6.02 //x2=55.54 //y2=4.865
r894 (  98 257 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.1 //y=6.02 //x2=55.1 //y2=4.865
r895 (  97 158 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.11 //y=6.02 //x2=41.11 //y2=4.865
r896 (  96 246 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=40.67 //y=6.02 //x2=40.67 //y2=4.865
r897 (  95 139 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.68 //y=6.02 //x2=26.68 //y2=4.865
r898 (  94 235 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.24 //y=6.02 //x2=26.24 //y2=4.865
r899 (  93 120 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.25 //y=6.02 //x2=12.25 //y2=4.865
r900 (  92 224 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.81 //y=6.02 //x2=11.81 //y2=4.865
r901 (  91 203 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=83.817 //y=1.375 //x2=83.925 //y2=1.375
r902 (  91 204 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=83.817 //y=1.375 //x2=83.71 //y2=1.375
r903 (  90 184 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=69.387 //y=1.375 //x2=69.495 //y2=1.375
r904 (  90 185 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=69.387 //y=1.375 //x2=69.28 //y2=1.375
r905 (  89 165 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=54.957 //y=1.375 //x2=55.065 //y2=1.375
r906 (  89 166 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=54.957 //y=1.375 //x2=54.85 //y2=1.375
r907 (  88 146 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=40.527 //y=1.375 //x2=40.635 //y2=1.375
r908 (  88 147 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=40.527 //y=1.375 //x2=40.42 //y2=1.375
r909 (  87 127 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=26.097 //y=1.375 //x2=26.205 //y2=1.375
r910 (  87 128 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=26.097 //y=1.375 //x2=25.99 //y2=1.375
r911 (  86 108 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=11.667 //y=1.375 //x2=11.775 //y2=1.375
r912 (  86 109 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=11.667 //y=1.375 //x2=11.56 //y2=1.375
r913 (  84 276 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=83.99 //y=4.7 //x2=83.99 //y2=4.7
r914 (  82 84 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=83.99 //y=2.96 //x2=83.99 //y2=4.7
r915 (  79 283 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=83.99 //y=2.08 //x2=83.99 //y2=2.08
r916 (  79 82 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=83.99 //y=2.08 //x2=83.99 //y2=2.96
r917 (  76 265 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=69.56 //y=4.7 //x2=69.56 //y2=4.7
r918 (  70 272 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=69.56 //y=2.08 //x2=69.56 //y2=2.08
r919 (  67 254 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.13 //y=4.7 //x2=55.13 //y2=4.7
r920 (  61 261 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.13 //y=2.08 //x2=55.13 //y2=2.08
r921 (  58 243 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=40.7 //y=4.7 //x2=40.7 //y2=4.7
r922 (  52 250 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=40.7 //y=2.08 //x2=40.7 //y2=2.08
r923 (  49 232 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=4.7 //x2=26.27 //y2=4.7
r924 (  43 239 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=2.08 //x2=26.27 //y2=2.08
r925 (  40 221 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=4.7 //x2=11.84 //y2=4.7
r926 (  34 228 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=2.08 //x2=11.84 //y2=2.08
r927 (  32 76 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=69.56 //y=2.96 //x2=69.56 //y2=4.7
r928 (  31 32 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=69.56 //y=2.59 //x2=69.56 //y2=2.96
r929 (  31 70 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=69.56 //y=2.59 //x2=69.56 //y2=2.08
r930 (  30 67 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=55.13 //y=2.96 //x2=55.13 //y2=4.7
r931 (  29 30 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=55.13 //y=2.59 //x2=55.13 //y2=2.96
r932 (  29 61 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=55.13 //y=2.59 //x2=55.13 //y2=2.08
r933 (  28 58 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=40.7 //y=2.96 //x2=40.7 //y2=4.7
r934 (  27 28 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=40.7 //y=2.59 //x2=40.7 //y2=2.96
r935 (  27 52 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=40.7 //y=2.59 //x2=40.7 //y2=2.08
r936 (  26 49 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.96 //x2=26.27 //y2=4.7
r937 (  25 26 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.59 //x2=26.27 //y2=2.96
r938 (  25 43 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.59 //x2=26.27 //y2=2.08
r939 (  24 40 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.96 //x2=11.84 //y2=4.7
r940 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.59 //x2=11.84 //y2=2.96
r941 (  23 34 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.59 //x2=11.84 //y2=2.08
r942 (  22 82 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=83.99 //y=2.96 //x2=83.99 //y2=2.96
r943 (  20 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=69.56 //y=2.96 //x2=69.56 //y2=2.96
r944 (  18 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=55.13 //y=2.96 //x2=55.13 //y2=2.96
r945 (  16 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=40.7 //y=2.96 //x2=40.7 //y2=2.96
r946 (  14 26 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=26.27 //y=2.96 //x2=26.27 //y2=2.96
r947 (  12 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.84 //y=2.96 //x2=11.84 //y2=2.96
r948 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.675 //y=2.96 //x2=69.56 //y2=2.96
r949 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=83.875 //y=2.96 //x2=83.99 //y2=2.96
r950 (  9 10 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=83.875 //y=2.96 //x2=69.675 //y2=2.96
r951 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.245 //y=2.96 //x2=55.13 //y2=2.96
r952 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.445 //y=2.96 //x2=69.56 //y2=2.96
r953 (  7 8 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=69.445 //y=2.96 //x2=55.245 //y2=2.96
r954 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=40.815 //y=2.96 //x2=40.7 //y2=2.96
r955 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.015 //y=2.96 //x2=55.13 //y2=2.96
r956 (  5 6 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=55.015 //y=2.96 //x2=40.815 //y2=2.96
r957 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=26.385 //y=2.96 //x2=26.27 //y2=2.96
r958 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=40.585 //y=2.96 //x2=40.7 //y2=2.96
r959 (  3 4 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=40.585 //y=2.96 //x2=26.385 //y2=2.96
r960 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.955 //y=2.96 //x2=11.84 //y2=2.96
r961 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=2.96 //x2=26.27 //y2=2.96
r962 (  1 2 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=2.96 //x2=11.955 //y2=2.96
ends PM_TMRDFFSNRNQX1\%SN

subckt PM_TMRDFFSNRNQX1\%noxref_23 ( 1 2 3 4 5 6 16 24 37 38 45 53 59 60 64 66 \
 73 74 75 76 77 78 79 80 81 82 83 87 88 89 94 96 99 100 104 105 106 111 113 \
 116 117 121 122 123 128 130 133 134 136 137 142 146 147 152 156 157 162 165 \
 167 168 169 )
c345 ( 169 0 ) capacitor c=0.023087f //x=75.295 //y=5.02
c346 ( 168 0 ) capacitor c=0.023519f //x=74.415 //y=5.02
c347 ( 167 0 ) capacitor c=0.0224735f //x=73.535 //y=5.02
c348 ( 165 0 ) capacitor c=0.00853354f //x=75.545 //y=0.915
c349 ( 162 0 ) capacitor c=0.0587755f //x=85.1 //y=4.7
c350 ( 157 0 ) capacitor c=0.0273931f //x=85.1 //y=1.915
c351 ( 156 0 ) capacitor c=0.0462455f //x=85.1 //y=2.08
c352 ( 152 0 ) capacitor c=0.0588394f //x=70.67 //y=4.7
c353 ( 147 0 ) capacitor c=0.0273931f //x=70.67 //y=1.915
c354 ( 146 0 ) capacitor c=0.0456313f //x=70.67 //y=2.08
c355 ( 142 0 ) capacitor c=0.0589949f //x=65.86 //y=4.7
c356 ( 137 0 ) capacitor c=0.0273931f //x=65.86 //y=1.915
c357 ( 136 0 ) capacitor c=0.0456313f //x=65.86 //y=2.08
c358 ( 134 0 ) capacitor c=0.0432517f //x=85.62 //y=1.26
c359 ( 133 0 ) capacitor c=0.0200379f //x=85.62 //y=0.915
c360 ( 130 0 ) capacitor c=0.0148873f //x=85.465 //y=1.415
c361 ( 128 0 ) capacitor c=0.0157803f //x=85.465 //y=0.76
c362 ( 123 0 ) capacitor c=0.0218028f //x=85.09 //y=1.57
c363 ( 122 0 ) capacitor c=0.0207459f //x=85.09 //y=1.26
c364 ( 121 0 ) capacitor c=0.0194308f //x=85.09 //y=0.915
c365 ( 117 0 ) capacitor c=0.0432517f //x=71.19 //y=1.26
c366 ( 116 0 ) capacitor c=0.0200379f //x=71.19 //y=0.915
c367 ( 113 0 ) capacitor c=0.0148873f //x=71.035 //y=1.415
c368 ( 111 0 ) capacitor c=0.0157803f //x=71.035 //y=0.76
c369 ( 106 0 ) capacitor c=0.0218028f //x=70.66 //y=1.57
c370 ( 105 0 ) capacitor c=0.0207459f //x=70.66 //y=1.26
c371 ( 104 0 ) capacitor c=0.0194308f //x=70.66 //y=0.915
c372 ( 100 0 ) capacitor c=0.0432517f //x=66.38 //y=1.26
c373 ( 99 0 ) capacitor c=0.0200379f //x=66.38 //y=0.915
c374 ( 96 0 ) capacitor c=0.0148873f //x=66.225 //y=1.415
c375 ( 94 0 ) capacitor c=0.0157803f //x=66.225 //y=0.76
c376 ( 89 0 ) capacitor c=0.0218028f //x=65.85 //y=1.57
c377 ( 88 0 ) capacitor c=0.0207459f //x=65.85 //y=1.26
c378 ( 87 0 ) capacitor c=0.0194308f //x=65.85 //y=0.915
c379 ( 83 0 ) capacitor c=0.158794f //x=85.28 //y=6.02
c380 ( 82 0 ) capacitor c=0.110114f //x=84.84 //y=6.02
c381 ( 81 0 ) capacitor c=0.158754f //x=70.85 //y=6.02
c382 ( 80 0 ) capacitor c=0.109949f //x=70.41 //y=6.02
c383 ( 79 0 ) capacitor c=0.158754f //x=66.04 //y=6.02
c384 ( 78 0 ) capacitor c=0.109949f //x=65.6 //y=6.02
c385 ( 74 0 ) capacitor c=0.00106608f //x=75.44 //y=5.155
c386 ( 73 0 ) capacitor c=0.00191414f //x=74.56 //y=5.155
c387 ( 66 0 ) capacitor c=0.0857665f //x=85.1 //y=2.08
c388 ( 64 0 ) capacitor c=0.10494f //x=76.22 //y=3.7
c389 ( 60 0 ) capacitor c=0.00398962f //x=75.82 //y=1.665
c390 ( 59 0 ) capacitor c=0.0137288f //x=76.135 //y=1.665
c391 ( 53 0 ) capacitor c=0.0283082f //x=76.135 //y=5.155
c392 ( 45 0 ) capacitor c=0.0170864f //x=75.355 //y=5.155
c393 ( 38 0 ) capacitor c=0.00316998f //x=73.765 //y=5.155
c394 ( 37 0 ) capacitor c=0.014258f //x=74.475 //y=5.155
c395 ( 24 0 ) capacitor c=0.0790362f //x=70.67 //y=2.08
c396 ( 16 0 ) capacitor c=0.076565f //x=65.86 //y=2.08
c397 ( 6 0 ) capacitor c=0.0055354f //x=76.335 //y=3.7
c398 ( 5 0 ) capacitor c=0.167028f //x=84.985 //y=3.7
c399 ( 4 0 ) capacitor c=0.00533183f //x=70.785 //y=3.7
c400 ( 3 0 ) capacitor c=0.0753575f //x=76.105 //y=3.7
c401 ( 2 0 ) capacitor c=0.00692093f //x=65.975 //y=3.7
c402 ( 1 0 ) capacitor c=0.0665749f //x=70.555 //y=3.7
r403 (  156 157 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=85.1 //y=2.08 //x2=85.1 //y2=1.915
r404 (  146 147 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=70.67 //y=2.08 //x2=70.67 //y2=1.915
r405 (  136 137 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=65.86 //y=2.08 //x2=65.86 //y2=1.915
r406 (  134 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.62 //y=1.26 //x2=85.58 //y2=1.415
r407 (  133 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.62 //y=0.915 //x2=85.58 //y2=0.76
r408 (  133 134 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=85.62 //y=0.915 //x2=85.62 //y2=1.26
r409 (  131 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.245 //y=1.415 //x2=85.13 //y2=1.415
r410 (  130 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.465 //y=1.415 //x2=85.58 //y2=1.415
r411 (  129 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.245 //y=0.76 //x2=85.13 //y2=0.76
r412 (  128 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.465 //y=0.76 //x2=85.58 //y2=0.76
r413 (  128 129 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=85.465 //y=0.76 //x2=85.245 //y2=0.76
r414 (  125 162 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=85.28 //y=4.865 //x2=85.1 //y2=4.7
r415 (  123 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.09 //y=1.57 //x2=85.13 //y2=1.415
r416 (  123 157 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=85.09 //y=1.57 //x2=85.09 //y2=1.915
r417 (  122 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.09 //y=1.26 //x2=85.13 //y2=1.415
r418 (  121 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.09 //y=0.915 //x2=85.13 //y2=0.76
r419 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=85.09 //y=0.915 //x2=85.09 //y2=1.26
r420 (  118 162 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=84.84 //y=4.865 //x2=85.1 //y2=4.7
r421 (  117 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.19 //y=1.26 //x2=71.15 //y2=1.415
r422 (  116 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.19 //y=0.915 //x2=71.15 //y2=0.76
r423 (  116 117 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=71.19 //y=0.915 //x2=71.19 //y2=1.26
r424 (  114 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.815 //y=1.415 //x2=70.7 //y2=1.415
r425 (  113 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.035 //y=1.415 //x2=71.15 //y2=1.415
r426 (  112 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.815 //y=0.76 //x2=70.7 //y2=0.76
r427 (  111 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.035 //y=0.76 //x2=71.15 //y2=0.76
r428 (  111 112 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=71.035 //y=0.76 //x2=70.815 //y2=0.76
r429 (  108 152 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=70.85 //y=4.865 //x2=70.67 //y2=4.7
r430 (  106 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.66 //y=1.57 //x2=70.7 //y2=1.415
r431 (  106 147 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=70.66 //y=1.57 //x2=70.66 //y2=1.915
r432 (  105 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.66 //y=1.26 //x2=70.7 //y2=1.415
r433 (  104 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.66 //y=0.915 //x2=70.7 //y2=0.76
r434 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=70.66 //y=0.915 //x2=70.66 //y2=1.26
r435 (  101 152 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=70.41 //y=4.865 //x2=70.67 //y2=4.7
r436 (  100 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.38 //y=1.26 //x2=66.34 //y2=1.415
r437 (  99 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.38 //y=0.915 //x2=66.34 //y2=0.76
r438 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=66.38 //y=0.915 //x2=66.38 //y2=1.26
r439 (  97 140 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.005 //y=1.415 //x2=65.89 //y2=1.415
r440 (  96 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.225 //y=1.415 //x2=66.34 //y2=1.415
r441 (  95 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.005 //y=0.76 //x2=65.89 //y2=0.76
r442 (  94 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.225 //y=0.76 //x2=66.34 //y2=0.76
r443 (  94 95 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=66.225 //y=0.76 //x2=66.005 //y2=0.76
r444 (  91 142 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=66.04 //y=4.865 //x2=65.86 //y2=4.7
r445 (  89 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.85 //y=1.57 //x2=65.89 //y2=1.415
r446 (  89 137 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=65.85 //y=1.57 //x2=65.85 //y2=1.915
r447 (  88 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.85 //y=1.26 //x2=65.89 //y2=1.415
r448 (  87 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.85 //y=0.915 //x2=65.89 //y2=0.76
r449 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=65.85 //y=0.915 //x2=65.85 //y2=1.26
r450 (  84 142 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=65.6 //y=4.865 //x2=65.86 //y2=4.7
r451 (  83 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=85.28 //y=6.02 //x2=85.28 //y2=4.865
r452 (  82 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=84.84 //y=6.02 //x2=84.84 //y2=4.865
r453 (  81 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.85 //y=6.02 //x2=70.85 //y2=4.865
r454 (  80 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.41 //y=6.02 //x2=70.41 //y2=4.865
r455 (  79 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.04 //y=6.02 //x2=66.04 //y2=4.865
r456 (  78 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=65.6 //y=6.02 //x2=65.6 //y2=4.865
r457 (  77 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=85.355 //y=1.415 //x2=85.465 //y2=1.415
r458 (  77 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=85.355 //y=1.415 //x2=85.245 //y2=1.415
r459 (  76 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=70.925 //y=1.415 //x2=71.035 //y2=1.415
r460 (  76 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=70.925 //y=1.415 //x2=70.815 //y2=1.415
r461 (  75 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.115 //y=1.415 //x2=66.225 //y2=1.415
r462 (  75 97 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.115 //y=1.415 //x2=66.005 //y2=1.415
r463 (  71 162 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=85.1 //y=4.7 //x2=85.1 //y2=4.7
r464 (  69 71 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=85.1 //y=3.7 //x2=85.1 //y2=4.7
r465 (  66 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=85.1 //y=2.08 //x2=85.1 //y2=2.08
r466 (  66 69 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=85.1 //y=2.08 //x2=85.1 //y2=3.7
r467 (  62 64 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=76.22 //y=5.07 //x2=76.22 //y2=3.7
r468 (  61 64 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=76.22 //y=1.75 //x2=76.22 //y2=3.7
r469 (  59 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=76.135 //y=1.665 //x2=76.22 //y2=1.75
r470 (  59 60 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=76.135 //y=1.665 //x2=75.82 //y2=1.665
r471 (  55 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=75.735 //y=1.58 //x2=75.82 //y2=1.665
r472 (  55 165 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=75.735 //y=1.58 //x2=75.735 //y2=1.01
r473 (  54 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.525 //y=5.155 //x2=75.44 //y2=5.155
r474 (  53 62 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=76.135 //y=5.155 //x2=76.22 //y2=5.07
r475 (  53 54 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=76.135 //y=5.155 //x2=75.525 //y2=5.155
r476 (  47 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.44 //y=5.24 //x2=75.44 //y2=5.155
r477 (  47 169 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=75.44 //y=5.24 //x2=75.44 //y2=5.725
r478 (  46 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.645 //y=5.155 //x2=74.56 //y2=5.155
r479 (  45 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.355 //y=5.155 //x2=75.44 //y2=5.155
r480 (  45 46 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=75.355 //y=5.155 //x2=74.645 //y2=5.155
r481 (  39 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.56 //y=5.24 //x2=74.56 //y2=5.155
r482 (  39 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=74.56 //y=5.24 //x2=74.56 //y2=5.725
r483 (  37 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.475 //y=5.155 //x2=74.56 //y2=5.155
r484 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=74.475 //y=5.155 //x2=73.765 //y2=5.155
r485 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=73.68 //y=5.24 //x2=73.765 //y2=5.155
r486 (  31 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=73.68 //y=5.24 //x2=73.68 //y2=5.725
r487 (  29 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=4.7 //x2=70.67 //y2=4.7
r488 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=70.67 //y=3.7 //x2=70.67 //y2=4.7
r489 (  24 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=2.08 //x2=70.67 //y2=2.08
r490 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=70.67 //y=2.08 //x2=70.67 //y2=3.7
r491 (  21 142 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=65.86 //y=4.7 //x2=65.86 //y2=4.7
r492 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=65.86 //y=3.7 //x2=65.86 //y2=4.7
r493 (  16 136 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=65.86 //y=2.08 //x2=65.86 //y2=2.08
r494 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=65.86 //y=2.08 //x2=65.86 //y2=3.7
r495 (  14 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=85.1 //y=3.7 //x2=85.1 //y2=3.7
r496 (  12 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=76.22 //y=3.7 //x2=76.22 //y2=3.7
r497 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=70.67 //y=3.7 //x2=70.67 //y2=3.7
r498 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=65.86 //y=3.7 //x2=65.86 //y2=3.7
r499 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=76.335 //y=3.7 //x2=76.22 //y2=3.7
r500 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=84.985 //y=3.7 //x2=85.1 //y2=3.7
r501 (  5 6 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=84.985 //y=3.7 //x2=76.335 //y2=3.7
r502 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=70.785 //y=3.7 //x2=70.67 //y2=3.7
r503 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=76.105 //y=3.7 //x2=76.22 //y2=3.7
r504 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=76.105 //y=3.7 //x2=70.785 //y2=3.7
r505 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=65.975 //y=3.7 //x2=65.86 //y2=3.7
r506 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=3.7 //x2=70.67 //y2=3.7
r507 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=3.7 //x2=65.975 //y2=3.7
ends PM_TMRDFFSNRNQX1\%noxref_23

subckt PM_TMRDFFSNRNQX1\%noxref_24 ( 1 2 13 14 15 23 29 30 37 50 51 52 53 54 )
c91 ( 54 0 ) capacitor c=0.034295f //x=92.305 //y=5.025
c92 ( 53 0 ) capacitor c=0.0174957f //x=91.425 //y=5.025
c93 ( 51 0 ) capacitor c=0.0214849f //x=88.545 //y=5.025
c94 ( 50 0 ) capacitor c=0.0217161f //x=87.665 //y=5.025
c95 ( 49 0 ) capacitor c=0.00115294f //x=91.57 //y=6.91
c96 ( 37 0 ) capacitor c=0.0131238f //x=92.365 //y=6.91
c97 ( 30 0 ) capacitor c=0.00386507f //x=90.775 //y=6.91
c98 ( 29 0 ) capacitor c=0.00951687f //x=91.485 //y=6.91
c99 ( 23 0 ) capacitor c=0.0455351f //x=90.69 //y=5.21
c100 ( 15 0 ) capacitor c=0.00871244f //x=88.69 //y=5.295
c101 ( 14 0 ) capacitor c=0.00290434f //x=87.895 //y=5.21
c102 ( 13 0 ) capacitor c=0.0139202f //x=88.605 //y=5.21
c103 ( 2 0 ) capacitor c=0.0091252f //x=88.805 //y=5.21
c104 ( 1 0 ) capacitor c=0.0484159f //x=90.575 //y=5.21
r105 (  39 54 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=92.45 //y=6.825 //x2=92.45 //y2=6.74
r106 (  38 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.655 //y=6.91 //x2=91.57 //y2=6.91
r107 (  37 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=92.365 //y=6.91 //x2=92.45 //y2=6.825
r108 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=92.365 //y=6.91 //x2=91.655 //y2=6.91
r109 (  31 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.57 //y=6.825 //x2=91.57 //y2=6.91
r110 (  31 53 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.57 //y=6.825 //x2=91.57 //y2=6.74
r111 (  29 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=91.485 //y=6.91 //x2=91.57 //y2=6.91
r112 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=91.485 //y=6.91 //x2=90.775 //y2=6.91
r113 (  23 52 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=90.69 //y=5.21 //x2=90.69 //y2=6.06
r114 (  21 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=90.69 //y=6.825 //x2=90.775 //y2=6.91
r115 (  21 52 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=90.69 //y=6.825 //x2=90.69 //y2=6.74
r116 (  15 48 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=88.69 //y=5.295 //x2=88.69 //y2=5.17
r117 (  15 51 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=88.69 //y=5.295 //x2=88.69 //y2=6.06
r118 (  13 48 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=88.605 //y=5.21 //x2=88.69 //y2=5.17
r119 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=88.605 //y=5.21 //x2=87.895 //y2=5.21
r120 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=87.81 //y=5.295 //x2=87.895 //y2=5.21
r121 (  7 50 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=87.81 //y=5.295 //x2=87.81 //y2=5.72
r122 (  6 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=90.69 //y=5.21 //x2=90.69 //y2=5.21
r123 (  4 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=88.69 //y=5.21 //x2=88.69 //y2=5.21
r124 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=88.805 //y=5.21 //x2=88.69 //y2=5.21
r125 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=90.575 //y=5.21 //x2=90.69 //y2=5.21
r126 (  1 2 ) resistor r=1.68893 //w=0.131 //l=1.77 //layer=m1 \
 //thickness=0.36 //x=90.575 //y=5.21 //x2=88.805 //y2=5.21
ends PM_TMRDFFSNRNQX1\%noxref_24

subckt PM_TMRDFFSNRNQX1\%noxref_25 ( 1 2 3 4 5 12 17 30 31 38 46 52 53 57 59 \
 66 72 73 74 75 76 77 78 79 80 81 82 86 87 88 93 95 98 99 103 104 105 106 107 \
 109 112 115 116 117 118 119 120 121 122 126 128 131 132 133 134 139 140 145 \
 157 164 166 167 168 )
c390 ( 168 0 ) capacitor c=0.023087f //x=84.915 //y=5.02
c391 ( 167 0 ) capacitor c=0.023519f //x=84.035 //y=5.02
c392 ( 166 0 ) capacitor c=0.0224735f //x=83.155 //y=5.02
c393 ( 164 0 ) capacitor c=0.0087111f //x=85.165 //y=0.915
c394 ( 157 0 ) capacitor c=0.0583848f //x=93.98 //y=2.08
c395 ( 145 0 ) capacitor c=0.0587755f //x=80.29 //y=4.7
c396 ( 140 0 ) capacitor c=0.0273931f //x=80.29 //y=1.915
c397 ( 139 0 ) capacitor c=0.0457326f //x=80.29 //y=2.08
c398 ( 134 0 ) capacitor c=0.0316774f //x=94.685 //y=1.21
c399 ( 133 0 ) capacitor c=0.0187384f //x=94.685 //y=0.865
c400 ( 132 0 ) capacitor c=0.0590362f //x=94.325 //y=4.795
c401 ( 131 0 ) capacitor c=0.0296075f //x=94.615 //y=4.795
c402 ( 128 0 ) capacitor c=0.0157912f //x=94.53 //y=1.365
c403 ( 126 0 ) capacitor c=0.0149844f //x=94.53 //y=0.71
c404 ( 122 0 ) capacitor c=0.0302441f //x=94.155 //y=1.915
c405 ( 121 0 ) capacitor c=0.0234157f //x=94.155 //y=1.52
c406 ( 120 0 ) capacitor c=0.0234376f //x=94.155 //y=1.21
c407 ( 119 0 ) capacitor c=0.0199931f //x=94.155 //y=0.865
c408 ( 118 0 ) capacitor c=0.092271f //x=92.325 //y=1.915
c409 ( 117 0 ) capacitor c=0.0249466f //x=92.325 //y=1.56
c410 ( 116 0 ) capacitor c=0.0234397f //x=92.325 //y=1.25
c411 ( 115 0 ) capacitor c=0.0193195f //x=92.325 //y=0.905
c412 ( 112 0 ) capacitor c=0.0631944f //x=92.23 //y=4.87
c413 ( 109 0 ) capacitor c=0.0164325f //x=92.17 //y=1.405
c414 ( 107 0 ) capacitor c=0.0157803f //x=92.17 //y=0.75
c415 ( 106 0 ) capacitor c=0.010629f //x=91.865 //y=4.795
c416 ( 105 0 ) capacitor c=0.0194269f //x=92.155 //y=4.795
c417 ( 104 0 ) capacitor c=0.0353695f //x=91.795 //y=1.25
c418 ( 103 0 ) capacitor c=0.0175988f //x=91.795 //y=0.905
c419 ( 99 0 ) capacitor c=0.0432517f //x=80.81 //y=1.26
c420 ( 98 0 ) capacitor c=0.0200379f //x=80.81 //y=0.915
c421 ( 95 0 ) capacitor c=0.0148873f //x=80.655 //y=1.415
c422 ( 93 0 ) capacitor c=0.0157803f //x=80.655 //y=0.76
c423 ( 88 0 ) capacitor c=0.0218028f //x=80.28 //y=1.57
c424 ( 87 0 ) capacitor c=0.0207459f //x=80.28 //y=1.26
c425 ( 86 0 ) capacitor c=0.0194308f //x=80.28 //y=0.915
c426 ( 82 0 ) capacitor c=0.110622f //x=94.69 //y=6.025
c427 ( 81 0 ) capacitor c=0.154068f //x=94.25 //y=6.025
c428 ( 80 0 ) capacitor c=0.154291f //x=92.23 //y=6.025
c429 ( 79 0 ) capacitor c=0.110404f //x=91.79 //y=6.025
c430 ( 78 0 ) capacitor c=0.158794f //x=80.47 //y=6.02
c431 ( 77 0 ) capacitor c=0.110114f //x=80.03 //y=6.02
c432 ( 73 0 ) capacitor c=0.00106608f //x=85.06 //y=5.155
c433 ( 72 0 ) capacitor c=0.00207319f //x=84.18 //y=5.155
c434 ( 66 0 ) capacitor c=0.100793f //x=93.98 //y=2.08
c435 ( 59 0 ) capacitor c=0.107544f //x=92.5 //y=2.08
c436 ( 57 0 ) capacitor c=0.110556f //x=85.84 //y=2.22
c437 ( 53 0 ) capacitor c=0.00398962f //x=85.44 //y=1.665
c438 ( 52 0 ) capacitor c=0.0137249f //x=85.755 //y=1.665
c439 ( 46 0 ) capacitor c=0.0281866f //x=85.755 //y=5.155
c440 ( 38 0 ) capacitor c=0.0176454f //x=84.975 //y=5.155
c441 ( 31 0 ) capacitor c=0.00332903f //x=83.385 //y=5.155
c442 ( 30 0 ) capacitor c=0.0148427f //x=84.095 //y=5.155
c443 ( 17 0 ) capacitor c=0.0838223f //x=80.29 //y=2.08
c444 ( 12 0 ) capacitor c=0.0148272f //x=92.5 //y=2.08
c445 ( 5 0 ) capacitor c=0.0465668f //x=93.865 //y=2.08
c446 ( 4 0 ) capacitor c=0.0078573f //x=85.955 //y=2.22
c447 ( 3 0 ) capacitor c=0.190117f //x=92.355 //y=2.22
c448 ( 2 0 ) capacitor c=0.00906111f //x=80.405 //y=2.22
c449 ( 1 0 ) capacitor c=0.122867f //x=85.725 //y=2.22
r450 (  139 140 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=80.29 //y=2.08 //x2=80.29 //y2=1.915
r451 (  134 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.685 //y=1.21 //x2=94.645 //y2=1.365
r452 (  133 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.685 //y=0.865 //x2=94.645 //y2=0.71
r453 (  133 134 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=94.685 //y=0.865 //x2=94.685 //y2=1.21
r454 (  131 135 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=94.615 //y=4.795 //x2=94.69 //y2=4.87
r455 (  131 132 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=94.615 //y=4.795 //x2=94.325 //y2=4.795
r456 (  129 161 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=94.31 //y=1.365 //x2=94.195 //y2=1.365
r457 (  128 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=94.53 //y=1.365 //x2=94.645 //y2=1.365
r458 (  127 160 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=94.31 //y=0.71 //x2=94.195 //y2=0.71
r459 (  126 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=94.53 //y=0.71 //x2=94.645 //y2=0.71
r460 (  126 127 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=94.53 //y=0.71 //x2=94.31 //y2=0.71
r461 (  123 132 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=94.25 //y=4.87 //x2=94.325 //y2=4.795
r462 (  123 159 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=94.25 //y=4.87 //x2=93.98 //y2=4.705
r463 (  122 157 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=94.155 //y=1.915 //x2=93.98 //y2=2.08
r464 (  121 161 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.155 //y=1.52 //x2=94.195 //y2=1.365
r465 (  121 122 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=94.155 //y=1.52 //x2=94.155 //y2=1.915
r466 (  120 161 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.155 //y=1.21 //x2=94.195 //y2=1.365
r467 (  119 160 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=94.155 //y=0.865 //x2=94.195 //y2=0.71
r468 (  119 120 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=94.155 //y=0.865 //x2=94.155 //y2=1.21
r469 (  118 153 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=92.325 //y=1.915 //x2=92.5 //y2=2.08
r470 (  117 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=92.325 //y=1.56 //x2=92.285 //y2=1.405
r471 (  117 118 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=92.325 //y=1.56 //x2=92.325 //y2=1.915
r472 (  116 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=92.325 //y=1.25 //x2=92.285 //y2=1.405
r473 (  115 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=92.325 //y=0.905 //x2=92.285 //y2=0.75
r474 (  115 116 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=92.325 //y=0.905 //x2=92.325 //y2=1.25
r475 (  112 155 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=92.23 //y=4.87 //x2=92.5 //y2=4.705
r476 (  110 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=91.95 //y=1.405 //x2=91.835 //y2=1.405
r477 (  109 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=92.17 //y=1.405 //x2=92.285 //y2=1.405
r478 (  108 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=91.95 //y=0.75 //x2=91.835 //y2=0.75
r479 (  107 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=92.17 //y=0.75 //x2=92.285 //y2=0.75
r480 (  107 108 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=92.17 //y=0.75 //x2=91.95 //y2=0.75
r481 (  105 112 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=92.155 //y=4.795 //x2=92.23 //y2=4.87
r482 (  105 106 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=92.155 //y=4.795 //x2=91.865 //y2=4.795
r483 (  104 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=91.795 //y=1.25 //x2=91.835 //y2=1.405
r484 (  103 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=91.795 //y=0.905 //x2=91.835 //y2=0.75
r485 (  103 104 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=91.795 //y=0.905 //x2=91.795 //y2=1.25
r486 (  100 106 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=91.79 //y=4.87 //x2=91.865 //y2=4.795
r487 (  99 147 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.81 //y=1.26 //x2=80.77 //y2=1.415
r488 (  98 146 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.81 //y=0.915 //x2=80.77 //y2=0.76
r489 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=80.81 //y=0.915 //x2=80.81 //y2=1.26
r490 (  96 143 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.435 //y=1.415 //x2=80.32 //y2=1.415
r491 (  95 147 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.655 //y=1.415 //x2=80.77 //y2=1.415
r492 (  94 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.435 //y=0.76 //x2=80.32 //y2=0.76
r493 (  93 146 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.655 //y=0.76 //x2=80.77 //y2=0.76
r494 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=80.655 //y=0.76 //x2=80.435 //y2=0.76
r495 (  90 145 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=80.47 //y=4.865 //x2=80.29 //y2=4.7
r496 (  88 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.28 //y=1.57 //x2=80.32 //y2=1.415
r497 (  88 140 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=80.28 //y=1.57 //x2=80.28 //y2=1.915
r498 (  87 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.28 //y=1.26 //x2=80.32 //y2=1.415
r499 (  86 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.28 //y=0.915 //x2=80.32 //y2=0.76
r500 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=80.28 //y=0.915 //x2=80.28 //y2=1.26
r501 (  83 145 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=80.03 //y=4.865 //x2=80.29 //y2=4.7
r502 (  82 135 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=94.69 //y=6.025 //x2=94.69 //y2=4.87
r503 (  81 123 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=94.25 //y=6.025 //x2=94.25 //y2=4.87
r504 (  80 112 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=92.23 //y=6.025 //x2=92.23 //y2=4.87
r505 (  79 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=91.79 //y=6.025 //x2=91.79 //y2=4.87
r506 (  78 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=80.47 //y=6.02 //x2=80.47 //y2=4.865
r507 (  77 83 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=80.03 //y=6.02 //x2=80.03 //y2=4.865
r508 (  76 128 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=94.42 //y=1.365 //x2=94.53 //y2=1.365
r509 (  76 129 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=94.42 //y=1.365 //x2=94.31 //y2=1.365
r510 (  75 109 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=92.06 //y=1.405 //x2=92.17 //y2=1.405
r511 (  75 110 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=92.06 //y=1.405 //x2=91.95 //y2=1.405
r512 (  74 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=80.545 //y=1.415 //x2=80.655 //y2=1.415
r513 (  74 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=80.545 //y=1.415 //x2=80.435 //y2=1.415
r514 (  70 159 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=93.98 //y=4.705 //x2=93.98 //y2=4.705
r515 (  66 157 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=93.98 //y=2.08 //x2=93.98 //y2=2.08
r516 (  66 70 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=93.98 //y=2.08 //x2=93.98 //y2=4.705
r517 (  63 155 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=92.5 //y=4.705 //x2=92.5 //y2=4.705
r518 (  59 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=92.5 //y=2.08 //x2=92.5 //y2=2.08
r519 (  59 63 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=92.5 //y=2.08 //x2=92.5 //y2=4.705
r520 (  55 57 ) resistor r=195.08 //w=0.187 //l=2.85 //layer=li \
 //thickness=0.1 //x=85.84 //y=5.07 //x2=85.84 //y2=2.22
r521 (  54 57 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=85.84 //y=1.75 //x2=85.84 //y2=2.22
r522 (  52 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=85.755 //y=1.665 //x2=85.84 //y2=1.75
r523 (  52 53 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=85.755 //y=1.665 //x2=85.44 //y2=1.665
r524 (  48 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=85.355 //y=1.58 //x2=85.44 //y2=1.665
r525 (  48 164 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=85.355 //y=1.58 //x2=85.355 //y2=1.01
r526 (  47 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.145 //y=5.155 //x2=85.06 //y2=5.155
r527 (  46 55 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=85.755 //y=5.155 //x2=85.84 //y2=5.07
r528 (  46 47 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=85.755 //y=5.155 //x2=85.145 //y2=5.155
r529 (  40 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.06 //y=5.24 //x2=85.06 //y2=5.155
r530 (  40 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=85.06 //y=5.24 //x2=85.06 //y2=5.725
r531 (  39 72 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.265 //y=5.155 //x2=84.18 //y2=5.155
r532 (  38 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.975 //y=5.155 //x2=85.06 //y2=5.155
r533 (  38 39 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=84.975 //y=5.155 //x2=84.265 //y2=5.155
r534 (  32 72 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.18 //y=5.24 //x2=84.18 //y2=5.155
r535 (  32 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=84.18 //y=5.24 //x2=84.18 //y2=5.725
r536 (  30 72 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.095 //y=5.155 //x2=84.18 //y2=5.155
r537 (  30 31 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=84.095 //y=5.155 //x2=83.385 //y2=5.155
r538 (  24 31 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=83.3 //y=5.24 //x2=83.385 //y2=5.155
r539 (  24 166 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=83.3 //y=5.24 //x2=83.3 //y2=5.725
r540 (  22 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=80.29 //y=4.7 //x2=80.29 //y2=4.7
r541 (  20 22 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=80.29 //y=2.22 //x2=80.29 //y2=4.7
r542 (  17 139 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=80.29 //y=2.08 //x2=80.29 //y2=2.08
r543 (  17 20 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=80.29 //y=2.08 //x2=80.29 //y2=2.22
r544 (  15 66 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=93.98 //y=2.08 //x2=93.98 //y2=2.08
r545 (  12 59 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=92.5 //y=2.08 //x2=92.5 //y2=2.08
r546 (  12 13 ) resistor r=0.0678295 //w=0.258 //l=0.14 //layer=m1 \
 //thickness=0.36 //x=92.485 //y=2.08 //x2=92.485 //y2=2.22
r547 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=85.84 //y=2.22 //x2=85.84 //y2=2.22
r548 (  8 20 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=80.29 //y=2.22 //x2=80.29 //y2=2.22
r549 (  6 12 ) resistor r=0.032569 //w=0.258 //l=0.13 //layer=m1 \
 //thickness=0.36 //x=92.615 //y=2.08 //x2=92.485 //y2=2.08
r550 (  5 15 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=93.865 //y=2.08 //x2=93.98 //y2=2.08
r551 (  5 6 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=93.865 //y=2.08 //x2=92.615 //y2=2.08
r552 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=85.955 //y=2.22 //x2=85.84 //y2=2.22
r553 (  3 13 ) resistor r=0.032569 //w=0.258 //l=0.13 //layer=m1 \
 //thickness=0.36 //x=92.355 //y=2.22 //x2=92.485 //y2=2.22
r554 (  3 4 ) resistor r=6.10687 //w=0.131 //l=6.4 //layer=m1 //thickness=0.36 \
 //x=92.355 //y=2.22 //x2=85.955 //y2=2.22
r555 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=80.405 //y=2.22 //x2=80.29 //y2=2.22
r556 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=85.725 //y=2.22 //x2=85.84 //y2=2.22
r557 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=85.725 //y=2.22 //x2=80.405 //y2=2.22
ends PM_TMRDFFSNRNQX1\%noxref_25

subckt PM_TMRDFFSNRNQX1\%noxref_26 ( 1 2 13 14 15 21 27 28 35 46 47 48 49 50 )
c90 ( 50 0 ) capacitor c=0.0306574f //x=95.645 //y=5.025
c91 ( 49 0 ) capacitor c=0.0173945f //x=94.765 //y=5.025
c92 ( 47 0 ) capacitor c=0.0169278f //x=91.865 //y=5.025
c93 ( 46 0 ) capacitor c=0.0166762f //x=90.985 //y=5.025
c94 ( 45 0 ) capacitor c=0.00115294f //x=94.91 //y=6.91
c95 ( 35 0 ) capacitor c=0.0132983f //x=95.705 //y=6.91
c96 ( 28 0 ) capacitor c=0.00388794f //x=94.115 //y=6.91
c97 ( 27 0 ) capacitor c=0.00985708f //x=94.825 //y=6.91
c98 ( 21 0 ) capacitor c=0.0442221f //x=94.03 //y=5.21
c99 ( 15 0 ) capacitor c=0.0105083f //x=92.01 //y=5.295
c100 ( 14 0 ) capacitor c=0.00227812f //x=91.215 //y=5.21
c101 ( 13 0 ) capacitor c=0.0174384f //x=91.925 //y=5.21
c102 ( 2 0 ) capacitor c=0.00682032f //x=92.125 //y=5.21
c103 ( 1 0 ) capacitor c=0.0573196f //x=93.915 //y=5.21
r104 (  37 50 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=95.79 //y=6.825 //x2=95.79 //y2=6.74
r105 (  36 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.995 //y=6.91 //x2=94.91 //y2=6.91
r106 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=95.705 //y=6.91 //x2=95.79 //y2=6.825
r107 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=95.705 //y=6.91 //x2=94.995 //y2=6.91
r108 (  29 45 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.91 //y=6.825 //x2=94.91 //y2=6.91
r109 (  29 49 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.91 //y=6.825 //x2=94.91 //y2=6.74
r110 (  27 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.825 //y=6.91 //x2=94.91 //y2=6.91
r111 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=94.825 //y=6.91 //x2=94.115 //y2=6.91
r112 (  21 48 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=94.03 //y=5.21 //x2=94.03 //y2=6.06
r113 (  19 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=94.03 //y=6.825 //x2=94.115 //y2=6.91
r114 (  19 48 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=94.03 //y=6.825 //x2=94.03 //y2=6.74
r115 (  15 44 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=92.01 //y=5.295 //x2=92.01 //y2=5.17
r116 (  15 47 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=92.01 //y=5.295 //x2=92.01 //y2=6.06
r117 (  13 44 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=91.925 //y=5.21 //x2=92.01 //y2=5.17
r118 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=91.925 //y=5.21 //x2=91.215 //y2=5.21
r119 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=91.13 //y=5.295 //x2=91.215 //y2=5.21
r120 (  7 46 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=91.13 //y=5.295 //x2=91.13 //y2=5.72
r121 (  6 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=94.03 //y=5.21 //x2=94.03 //y2=5.21
r122 (  4 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=92.01 //y=5.21 //x2=92.01 //y2=5.21
r123 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=92.125 //y=5.21 //x2=92.01 //y2=5.21
r124 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=93.915 //y=5.21 //x2=94.03 //y2=5.21
r125 (  1 2 ) resistor r=1.70802 //w=0.131 //l=1.79 //layer=m1 \
 //thickness=0.36 //x=93.915 //y=5.21 //x2=92.125 //y2=5.21
ends PM_TMRDFFSNRNQX1\%noxref_26

subckt PM_TMRDFFSNRNQX1\%noxref_27 ( 1 2 3 4 5 6 29 30 43 45 46 50 52 63 64 65 \
 66 67 68 69 70 74 75 76 78 84 85 87 95 96 97 101 102 )
c242 ( 102 0 ) capacitor c=0.0167617f //x=95.205 //y=5.025
c243 ( 101 0 ) capacitor c=0.0164812f //x=94.325 //y=5.025
c244 ( 97 0 ) capacitor c=0.0110092f //x=95.2 //y=0.905
c245 ( 96 0 ) capacitor c=0.0131637f //x=91.87 //y=0.905
c246 ( 95 0 ) capacitor c=0.0131367f //x=88.54 //y=0.905
c247 ( 87 0 ) capacitor c=0.0537799f //x=97.31 //y=2.085
c248 ( 85 0 ) capacitor c=0.0435629f //x=97.95 //y=1.255
c249 ( 84 0 ) capacitor c=0.0200386f //x=97.95 //y=0.91
c250 ( 78 0 ) capacitor c=0.0152946f //x=97.795 //y=1.41
c251 ( 76 0 ) capacitor c=0.0157804f //x=97.795 //y=0.755
c252 ( 75 0 ) capacitor c=0.05065f //x=97.54 //y=4.79
c253 ( 74 0 ) capacitor c=0.0322983f //x=97.83 //y=4.79
c254 ( 70 0 ) capacitor c=0.0290017f //x=97.42 //y=1.92
c255 ( 69 0 ) capacitor c=0.0250027f //x=97.42 //y=1.565
c256 ( 68 0 ) capacitor c=0.0234316f //x=97.42 //y=1.255
c257 ( 67 0 ) capacitor c=0.0200596f //x=97.42 //y=0.91
c258 ( 66 0 ) capacitor c=0.154218f //x=97.905 //y=6.02
c259 ( 65 0 ) capacitor c=0.154243f //x=97.465 //y=6.02
c260 ( 63 0 ) capacitor c=0.00421476f //x=95.35 //y=5.21
c261 ( 52 0 ) capacitor c=0.09442f //x=97.31 //y=2.085
c262 ( 50 0 ) capacitor c=0.113028f //x=95.83 //y=4.07
c263 ( 46 0 ) capacitor c=0.00775877f //x=95.475 //y=1.645
c264 ( 45 0 ) capacitor c=0.0161066f //x=95.745 //y=1.645
c265 ( 43 0 ) capacitor c=0.0151634f //x=95.745 //y=5.21
c266 ( 30 0 ) capacitor c=0.0029383f //x=94.555 //y=5.21
c267 ( 29 0 ) capacitor c=0.0155464f //x=95.265 //y=5.21
c268 ( 6 0 ) capacitor c=0.00875763f //x=95.945 //y=4.07
c269 ( 5 0 ) capacitor c=0.0716061f //x=97.195 //y=4.07
c270 ( 4 0 ) capacitor c=0.00436966f //x=92.175 //y=1.18
c271 ( 3 0 ) capacitor c=0.069473f //x=95.275 //y=1.18
c272 ( 2 0 ) capacitor c=0.0141674f //x=88.845 //y=1.18
c273 ( 1 0 ) capacitor c=0.0494873f //x=91.945 //y=1.18
r274 (  87 88 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=97.31 //y=2.085 //x2=97.42 //y2=2.085
r275 (  85 94 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=97.95 //y=1.255 //x2=97.91 //y2=1.41
r276 (  84 93 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=97.95 //y=0.91 //x2=97.91 //y2=0.755
r277 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=97.95 //y=0.91 //x2=97.95 //y2=1.255
r278 (  79 92 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=97.575 //y=1.41 //x2=97.46 //y2=1.41
r279 (  78 94 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=97.795 //y=1.41 //x2=97.91 //y2=1.41
r280 (  77 91 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=97.575 //y=0.755 //x2=97.46 //y2=0.755
r281 (  76 93 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=97.795 //y=0.755 //x2=97.91 //y2=0.755
r282 (  76 77 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=97.795 //y=0.755 //x2=97.575 //y2=0.755
r283 (  74 81 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=97.83 //y=4.79 //x2=97.905 //y2=4.865
r284 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=97.83 //y=4.79 //x2=97.54 //y2=4.79
r285 (  71 75 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=97.465 //y=4.865 //x2=97.54 //y2=4.79
r286 (  71 90 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=97.465 //y=4.865 //x2=97.31 //y2=4.7
r287 (  70 88 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=97.42 //y=1.92 //x2=97.42 //y2=2.085
r288 (  69 92 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=97.42 //y=1.565 //x2=97.46 //y2=1.41
r289 (  69 70 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=97.42 //y=1.565 //x2=97.42 //y2=1.92
r290 (  68 92 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=97.42 //y=1.255 //x2=97.46 //y2=1.41
r291 (  67 91 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=97.42 //y=0.91 //x2=97.46 //y2=0.755
r292 (  67 68 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=97.42 //y=0.91 //x2=97.42 //y2=1.255
r293 (  66 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=97.905 //y=6.02 //x2=97.905 //y2=4.865
r294 (  65 71 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=97.465 //y=6.02 //x2=97.465 //y2=4.865
r295 (  64 78 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=97.685 //y=1.41 //x2=97.795 //y2=1.41
r296 (  64 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=97.685 //y=1.41 //x2=97.575 //y2=1.41
r297 (  62 95 ) resistor r=13.3953 //w=0.172 //l=0.18 //layer=li \
 //thickness=0.1 //x=88.727 //y=1.18 //x2=88.727 //y2=1
r298 (  57 90 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=97.31 //y=4.7 //x2=97.31 //y2=4.7
r299 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=97.31 //y=4.07 //x2=97.31 //y2=4.7
r300 (  52 87 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=97.31 //y=2.085 //x2=97.31 //y2=2.085
r301 (  52 55 ) resistor r=135.872 //w=0.187 //l=1.985 //layer=li \
 //thickness=0.1 //x=97.31 //y=2.085 //x2=97.31 //y2=4.07
r302 (  48 50 ) resistor r=72.2139 //w=0.187 //l=1.055 //layer=li \
 //thickness=0.1 //x=95.83 //y=5.125 //x2=95.83 //y2=4.07
r303 (  47 50 ) resistor r=160.171 //w=0.187 //l=2.34 //layer=li \
 //thickness=0.1 //x=95.83 //y=1.73 //x2=95.83 //y2=4.07
r304 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=95.745 //y=1.645 //x2=95.83 //y2=1.73
r305 (  45 46 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=95.745 //y=1.645 //x2=95.475 //y2=1.645
r306 (  44 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=95.435 //y=5.21 //x2=95.35 //y2=5.21
r307 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=95.745 //y=5.21 //x2=95.83 //y2=5.125
r308 (  43 44 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=95.745 //y=5.21 //x2=95.435 //y2=5.21
r309 (  42 97 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=95.39 //y=1.18 //x2=95.39 //y2=1
r310 (  37 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=95.39 //y=1.56 //x2=95.475 //y2=1.645
r311 (  37 42 ) resistor r=26.0107 //w=0.187 //l=0.38 //layer=li \
 //thickness=0.1 //x=95.39 //y=1.56 //x2=95.39 //y2=1.18
r312 (  31 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=95.35 //y=5.295 //x2=95.35 //y2=5.21
r313 (  31 102 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=95.35 //y=5.295 //x2=95.35 //y2=5.72
r314 (  29 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=95.265 //y=5.21 //x2=95.35 //y2=5.21
r315 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=95.265 //y=5.21 //x2=94.555 //y2=5.21
r316 (  23 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=94.47 //y=5.295 //x2=94.555 //y2=5.21
r317 (  23 101 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=94.47 //y=5.295 //x2=94.47 //y2=5.72
r318 (  21 96 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=92.06 //y=1.18 //x2=92.06 //y2=1
r319 (  16 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=97.31 //y=4.07 //x2=97.31 //y2=4.07
r320 (  14 50 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=95.83 //y=4.07 //x2=95.83 //y2=4.07
r321 (  12 42 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=95.39 //y=1.18 //x2=95.39 //y2=1.18
r322 (  10 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=92.06 //y=1.18 //x2=92.06 //y2=1.18
r323 (  8 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=88.73 //y=1.18 //x2=88.73 //y2=1.18
r324 (  6 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=95.945 //y=4.07 //x2=95.83 //y2=4.07
r325 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=97.195 //y=4.07 //x2=97.31 //y2=4.07
r326 (  5 6 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=97.195 //y=4.07 //x2=95.945 //y2=4.07
r327 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=92.175 //y=1.18 //x2=92.06 //y2=1.18
r328 (  3 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=95.275 //y=1.18 //x2=95.39 //y2=1.18
r329 (  3 4 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=95.275 //y=1.18 //x2=92.175 //y2=1.18
r330 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=88.845 //y=1.18 //x2=88.73 //y2=1.18
r331 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=91.945 //y=1.18 //x2=92.06 //y2=1.18
r332 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=91.945 //y=1.18 //x2=88.845 //y2=1.18
ends PM_TMRDFFSNRNQX1\%noxref_27

subckt PM_TMRDFFSNRNQX1\%Q ( 1 14 15 16 17 21 22 24 )
c52 ( 24 0 ) capacitor c=0.028734f //x=97.54 //y=5.02
c53 ( 22 0 ) capacitor c=0.0172744f //x=97.495 //y=0.91
c54 ( 21 0 ) capacitor c=0.102881f //x=98.05 //y=4.07
c55 ( 17 0 ) capacitor c=0.00575887f //x=97.77 //y=4.58
c56 ( 16 0 ) capacitor c=0.0131256f //x=97.965 //y=4.58
c57 ( 15 0 ) capacitor c=0.00636159f //x=97.765 //y=2.08
c58 ( 14 0 ) capacitor c=0.0140466f //x=97.965 //y=2.08
c59 ( 1 0 ) capacitor c=0.0237773f //x=98.05 //y=4.07
r60 (  19 21 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=98.05 //y=4.495 //x2=98.05 //y2=4.07
r61 (  18 21 ) resistor r=130.396 //w=0.187 //l=1.905 //layer=li \
 //thickness=0.1 //x=98.05 //y=2.165 //x2=98.05 //y2=4.07
r62 (  16 19 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=97.965 //y=4.58 //x2=98.05 //y2=4.495
r63 (  16 17 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=97.965 //y=4.58 //x2=97.77 //y2=4.58
r64 (  14 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=97.965 //y=2.08 //x2=98.05 //y2=2.165
r65 (  14 15 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=97.965 //y=2.08 //x2=97.765 //y2=2.08
r66 (  8 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=97.685 //y=4.665 //x2=97.77 //y2=4.58
r67 (  8 24 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li //thickness=0.1 \
 //x=97.685 //y=4.665 //x2=97.685 //y2=5.725
r68 (  4 15 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=97.68 //y=1.995 //x2=97.765 //y2=2.08
r69 (  4 22 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=97.68 //y=1.995 //x2=97.68 //y2=1.005
r70 (  1 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=98.05 //y=4.07 //x2=98.05 //y2=4.07
ends PM_TMRDFFSNRNQX1\%Q

subckt PM_TMRDFFSNRNQX1\%noxref_29 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0687824f //x=0.455 //y=0.375
c50 ( 17 0 ) capacitor c=0.0213512f //x=2.445 //y=1.59
c51 ( 13 0 ) capacitor c=0.015523f //x=2.445 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c53 ( 5 0 ) capacitor c=0.0204181f //x=1.475 //y=1.59
c54 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_29

subckt PM_TMRDFFSNRNQX1\%noxref_30 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=2.965 //y=0.375
c53 ( 28 0 ) capacitor c=0.00462395f //x=1.86 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=3.985 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=3.015 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_30

subckt PM_TMRDFFSNRNQX1\%noxref_31 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=5.265 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=7.255 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=7.255 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=6.37 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=6.285 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=5.4 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=1.59 //x2=6.37 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=1.59 //x2=6.855 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=1.59 //x2=7.34 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=1.59 //x2=6.855 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=0.54 //x2=6.37 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=0.54 //x2=6.855 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=0.54 //x2=7.34 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=0.54 //x2=6.855 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.485 //y=1.59 //x2=5.4 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.485 //y=1.59 //x2=5.885 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.285 //y=1.59 //x2=6.37 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.285 //y=1.59 //x2=5.885 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.4 //y=1.505 //x2=5.4 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.4 //y=1.505 //x2=5.4 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_31

subckt PM_TMRDFFSNRNQX1\%noxref_32 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=7.775 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=6.67 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=7.91 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=8.88 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=8.795 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=7.91 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=7.825 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.995 //y=0.54 //x2=7.91 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.995 //y=0.54 //x2=8.395 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.795 //y=0.54 //x2=8.88 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.795 //y=0.54 //x2=8.395 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.945 //y=0.995 //x2=6.86 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=7.91 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=6.945 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_32

subckt PM_TMRDFFSNRNQX1\%noxref_33 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=10.075 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=12.065 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=12.065 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=11.18 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=11.095 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=10.21 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.265 //y=1.59 //x2=11.18 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.265 //y=1.59 //x2=11.665 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.065 //y=1.59 //x2=12.15 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.065 //y=1.59 //x2=11.665 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.265 //y=0.54 //x2=11.18 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.265 //y=0.54 //x2=11.665 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.065 //y=0.54 //x2=12.15 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.065 //y=0.54 //x2=11.665 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=11.18 //y=1.505 //x2=11.18 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=11.18 //y=1.505 //x2=11.18 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.18 //y=0.625 //x2=11.18 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.18 //y=0.625 //x2=11.18 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.295 //y=1.59 //x2=10.21 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.295 //y=1.59 //x2=10.695 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.095 //y=1.59 //x2=11.18 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.095 //y=1.59 //x2=10.695 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=10.21 //y=1.505 //x2=10.21 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.21 //y=1.505 //x2=10.21 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_33

subckt PM_TMRDFFSNRNQX1\%noxref_34 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=12.585 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=11.48 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=12.72 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=13.69 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=13.605 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=12.72 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=12.635 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=13.69 //y=0.625 //x2=13.69 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=13.69 //y=0.625 //x2=13.69 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.805 //y=0.54 //x2=12.72 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.805 //y=0.54 //x2=13.205 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.605 //y=0.54 //x2=13.69 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.605 //y=0.54 //x2=13.205 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.72 //y=1.08 //x2=12.72 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=12.72 //y=1.08 //x2=12.72 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.91 //x2=12.72 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.91 //x2=12.72 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.625 //x2=12.72 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.625 //x2=12.72 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.755 //y=0.995 //x2=11.67 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.635 //y=0.995 //x2=12.72 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=12.635 //y=0.995 //x2=11.755 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_34

subckt PM_TMRDFFSNRNQX1\%noxref_35 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=14.885 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=16.875 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=16.875 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=15.99 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=15.905 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=15.02 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.075 //y=1.59 //x2=15.99 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.075 //y=1.59 //x2=16.475 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.875 //y=1.59 //x2=16.96 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.875 //y=1.59 //x2=16.475 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.075 //y=0.54 //x2=15.99 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.075 //y=0.54 //x2=16.475 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.875 //y=0.54 //x2=16.96 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.875 //y=0.54 //x2=16.475 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=15.99 //y=1.505 //x2=15.99 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.99 //y=1.505 //x2=15.99 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.99 //y=0.625 //x2=15.99 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=15.99 //y=0.625 //x2=15.99 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.105 //y=1.59 //x2=15.02 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.105 //y=1.59 //x2=15.505 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.905 //y=1.59 //x2=15.99 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.905 //y=1.59 //x2=15.505 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.02 //y=1.505 //x2=15.02 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.02 //y=1.505 //x2=15.02 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_35

subckt PM_TMRDFFSNRNQX1\%noxref_36 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=17.395 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=16.29 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=17.53 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=18.5 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=18.415 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=17.53 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=17.445 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=18.5 //y=0.625 //x2=18.5 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.5 //y=0.625 //x2=18.5 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.615 //y=0.54 //x2=17.53 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.615 //y=0.54 //x2=18.015 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.415 //y=0.54 //x2=18.5 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.415 //y=0.54 //x2=18.015 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.53 //y=1.08 //x2=17.53 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=17.53 //y=1.08 //x2=17.53 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.91 //x2=17.53 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.91 //x2=17.53 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.625 //x2=17.53 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.625 //x2=17.53 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.565 //y=0.995 //x2=16.48 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.445 //y=0.995 //x2=17.53 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=17.445 //y=0.995 //x2=16.565 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_36

subckt PM_TMRDFFSNRNQX1\%noxref_37 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=19.695 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=21.685 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=21.685 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=20.8 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=20.715 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=19.83 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.885 //y=1.59 //x2=20.8 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.885 //y=1.59 //x2=21.285 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.685 //y=1.59 //x2=21.77 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.685 //y=1.59 //x2=21.285 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.885 //y=0.54 //x2=20.8 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.885 //y=0.54 //x2=21.285 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.685 //y=0.54 //x2=21.77 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.685 //y=0.54 //x2=21.285 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=20.8 //y=1.505 //x2=20.8 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=20.8 //y=1.505 //x2=20.8 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.8 //y=0.625 //x2=20.8 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=20.8 //y=0.625 //x2=20.8 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.915 //y=1.59 //x2=19.83 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.915 //y=1.59 //x2=20.315 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.715 //y=1.59 //x2=20.8 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.715 //y=1.59 //x2=20.315 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=19.83 //y=1.505 //x2=19.83 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=19.83 //y=1.505 //x2=19.83 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_37

subckt PM_TMRDFFSNRNQX1\%noxref_38 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=22.205 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=21.1 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=22.34 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=23.31 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=23.225 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=22.34 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=22.255 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.31 //y=0.625 //x2=23.31 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=23.31 //y=0.625 //x2=23.31 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.425 //y=0.54 //x2=22.34 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.425 //y=0.54 //x2=22.825 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.225 //y=0.54 //x2=23.31 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.225 //y=0.54 //x2=22.825 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.34 //y=1.08 //x2=22.34 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=22.34 //y=1.08 //x2=22.34 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.91 //x2=22.34 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.91 //x2=22.34 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.625 //x2=22.34 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.625 //x2=22.34 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.375 //y=0.995 //x2=21.29 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.255 //y=0.995 //x2=22.34 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=22.255 //y=0.995 //x2=21.375 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_38

subckt PM_TMRDFFSNRNQX1\%noxref_39 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=24.505 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=26.495 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=26.495 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=25.61 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=25.525 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=24.64 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.695 //y=1.59 //x2=25.61 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.695 //y=1.59 //x2=26.095 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.495 //y=1.59 //x2=26.58 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.495 //y=1.59 //x2=26.095 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.695 //y=0.54 //x2=25.61 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.695 //y=0.54 //x2=26.095 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.495 //y=0.54 //x2=26.58 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.495 //y=0.54 //x2=26.095 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=25.61 //y=1.505 //x2=25.61 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=25.61 //y=1.505 //x2=25.61 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=25.61 //y=0.625 //x2=25.61 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=25.61 //y=0.625 //x2=25.61 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.725 //y=1.59 //x2=24.64 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.725 //y=1.59 //x2=25.125 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.525 //y=1.59 //x2=25.61 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.525 //y=1.59 //x2=25.125 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=24.64 //y=1.505 //x2=24.64 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=24.64 //y=1.505 //x2=24.64 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_39

subckt PM_TMRDFFSNRNQX1\%noxref_40 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=27.015 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=25.91 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=27.15 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=28.12 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=28.035 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=27.15 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=27.065 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=28.12 //y=0.625 //x2=28.12 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=28.12 //y=0.625 //x2=28.12 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=27.235 //y=0.54 //x2=27.15 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=27.235 //y=0.54 //x2=27.635 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=28.035 //y=0.54 //x2=28.12 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.035 //y=0.54 //x2=27.635 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.15 //y=1.08 //x2=27.15 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=27.15 //y=1.08 //x2=27.15 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.91 //x2=27.15 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.91 //x2=27.15 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.625 //x2=27.15 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.625 //x2=27.15 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.185 //y=0.995 //x2=26.1 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.065 //y=0.995 //x2=27.15 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=27.065 //y=0.995 //x2=26.185 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_40

subckt PM_TMRDFFSNRNQX1\%noxref_41 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=29.315 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=31.305 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=31.305 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=30.42 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=30.335 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=29.45 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.505 //y=1.59 //x2=30.42 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.505 //y=1.59 //x2=30.905 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.305 //y=1.59 //x2=31.39 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=31.305 //y=1.59 //x2=30.905 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.505 //y=0.54 //x2=30.42 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.505 //y=0.54 //x2=30.905 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.305 //y=0.54 //x2=31.39 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=31.305 //y=0.54 //x2=30.905 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=30.42 //y=1.505 //x2=30.42 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=30.42 //y=1.505 //x2=30.42 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=30.42 //y=0.625 //x2=30.42 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=30.42 //y=0.625 //x2=30.42 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.535 //y=1.59 //x2=29.45 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.535 //y=1.59 //x2=29.935 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.335 //y=1.59 //x2=30.42 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.335 //y=1.59 //x2=29.935 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=29.45 //y=1.505 //x2=29.45 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=29.45 //y=1.505 //x2=29.45 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_41

subckt PM_TMRDFFSNRNQX1\%noxref_42 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=31.825 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=30.72 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=31.96 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=32.93 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=32.845 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=31.96 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=31.875 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=32.93 //y=0.625 //x2=32.93 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=32.93 //y=0.625 //x2=32.93 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=32.045 //y=0.54 //x2=31.96 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=32.045 //y=0.54 //x2=32.445 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=32.845 //y=0.54 //x2=32.93 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=32.845 //y=0.54 //x2=32.445 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=31.96 //y=1.08 //x2=31.96 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=31.96 //y=1.08 //x2=31.96 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=31.96 //y=0.91 //x2=31.96 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=31.96 //y=0.91 //x2=31.96 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=31.96 //y=0.625 //x2=31.96 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=31.96 //y=0.625 //x2=31.96 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.995 //y=0.995 //x2=30.91 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=31.875 //y=0.995 //x2=31.96 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=31.875 //y=0.995 //x2=30.995 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_42

subckt PM_TMRDFFSNRNQX1\%noxref_43 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=34.125 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=36.115 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=36.115 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=35.23 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=35.145 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=34.26 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=35.315 //y=1.59 //x2=35.23 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.315 //y=1.59 //x2=35.715 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.115 //y=1.59 //x2=36.2 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=36.115 //y=1.59 //x2=35.715 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=35.315 //y=0.54 //x2=35.23 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.315 //y=0.54 //x2=35.715 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.115 //y=0.54 //x2=36.2 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=36.115 //y=0.54 //x2=35.715 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=35.23 //y=1.505 //x2=35.23 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=35.23 //y=1.505 //x2=35.23 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=35.23 //y=0.625 //x2=35.23 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=35.23 //y=0.625 //x2=35.23 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.345 //y=1.59 //x2=34.26 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.345 //y=1.59 //x2=34.745 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=35.145 //y=1.59 //x2=35.23 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.145 //y=1.59 //x2=34.745 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=34.26 //y=1.505 //x2=34.26 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=34.26 //y=1.505 //x2=34.26 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_43

subckt PM_TMRDFFSNRNQX1\%noxref_44 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=36.635 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=35.53 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=36.77 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=37.74 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=37.655 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=36.77 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=36.685 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=37.74 //y=0.625 //x2=37.74 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=37.74 //y=0.625 //x2=37.74 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=36.855 //y=0.54 //x2=36.77 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=36.855 //y=0.54 //x2=37.255 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=37.655 //y=0.54 //x2=37.74 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=37.655 //y=0.54 //x2=37.255 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=36.77 //y=1.08 //x2=36.77 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=36.77 //y=1.08 //x2=36.77 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=36.77 //y=0.91 //x2=36.77 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=36.77 //y=0.91 //x2=36.77 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=36.77 //y=0.625 //x2=36.77 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=36.77 //y=0.625 //x2=36.77 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.805 //y=0.995 //x2=35.72 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=36.685 //y=0.995 //x2=36.77 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=36.685 //y=0.995 //x2=35.805 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_44

subckt PM_TMRDFFSNRNQX1\%noxref_45 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=38.935 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=40.925 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=40.925 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=40.04 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=39.955 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=39.07 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=40.125 //y=1.59 //x2=40.04 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.125 //y=1.59 //x2=40.525 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.925 //y=1.59 //x2=41.01 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.925 //y=1.59 //x2=40.525 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=40.125 //y=0.54 //x2=40.04 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.125 //y=0.54 //x2=40.525 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.925 //y=0.54 //x2=41.01 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.925 //y=0.54 //x2=40.525 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=40.04 //y=1.505 //x2=40.04 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=40.04 //y=1.505 //x2=40.04 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=40.04 //y=0.625 //x2=40.04 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=40.04 //y=0.625 //x2=40.04 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=39.155 //y=1.59 //x2=39.07 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=39.155 //y=1.59 //x2=39.555 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=39.955 //y=1.59 //x2=40.04 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=39.955 //y=1.59 //x2=39.555 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=39.07 //y=1.505 //x2=39.07 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=39.07 //y=1.505 //x2=39.07 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_45

subckt PM_TMRDFFSNRNQX1\%noxref_46 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=41.445 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=40.34 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=41.58 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=42.55 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=42.465 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=41.58 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=41.495 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=42.55 //y=0.625 //x2=42.55 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=42.55 //y=0.625 //x2=42.55 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=41.665 //y=0.54 //x2=41.58 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=41.665 //y=0.54 //x2=42.065 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=42.465 //y=0.54 //x2=42.55 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=42.465 //y=0.54 //x2=42.065 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=41.58 //y=1.08 //x2=41.58 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=41.58 //y=1.08 //x2=41.58 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=41.58 //y=0.91 //x2=41.58 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=41.58 //y=0.91 //x2=41.58 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=41.58 //y=0.625 //x2=41.58 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=41.58 //y=0.625 //x2=41.58 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.615 //y=0.995 //x2=40.53 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=41.495 //y=0.995 //x2=41.58 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=41.495 //y=0.995 //x2=40.615 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_46

subckt PM_TMRDFFSNRNQX1\%noxref_47 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=43.745 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=45.735 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=45.735 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=44.85 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=44.765 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=43.88 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.935 //y=1.59 //x2=44.85 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.935 //y=1.59 //x2=45.335 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.735 //y=1.59 //x2=45.82 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.735 //y=1.59 //x2=45.335 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.935 //y=0.54 //x2=44.85 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.935 //y=0.54 //x2=45.335 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.735 //y=0.54 //x2=45.82 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.735 //y=0.54 //x2=45.335 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=44.85 //y=1.505 //x2=44.85 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=44.85 //y=1.505 //x2=44.85 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=44.85 //y=0.625 //x2=44.85 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=44.85 //y=0.625 //x2=44.85 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=43.965 //y=1.59 //x2=43.88 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=43.965 //y=1.59 //x2=44.365 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.765 //y=1.59 //x2=44.85 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.765 //y=1.59 //x2=44.365 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=43.88 //y=1.505 //x2=43.88 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=43.88 //y=1.505 //x2=43.88 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_47

subckt PM_TMRDFFSNRNQX1\%noxref_48 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=46.255 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=45.15 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=46.39 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=47.36 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=47.275 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=46.39 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=46.305 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=47.36 //y=0.625 //x2=47.36 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=47.36 //y=0.625 //x2=47.36 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=46.475 //y=0.54 //x2=46.39 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.475 //y=0.54 //x2=46.875 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=47.275 //y=0.54 //x2=47.36 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=47.275 //y=0.54 //x2=46.875 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.39 //y=1.08 //x2=46.39 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=46.39 //y=1.08 //x2=46.39 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.39 //y=0.91 //x2=46.39 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=46.39 //y=0.91 //x2=46.39 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=46.39 //y=0.625 //x2=46.39 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=46.39 //y=0.625 //x2=46.39 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.425 //y=0.995 //x2=45.34 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.305 //y=0.995 //x2=46.39 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=46.305 //y=0.995 //x2=45.425 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_48

subckt PM_TMRDFFSNRNQX1\%noxref_49 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=48.555 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=50.545 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=50.545 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=49.66 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=49.575 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=48.69 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.745 //y=1.59 //x2=49.66 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.745 //y=1.59 //x2=50.145 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.545 //y=1.59 //x2=50.63 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.545 //y=1.59 //x2=50.145 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.745 //y=0.54 //x2=49.66 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.745 //y=0.54 //x2=50.145 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.545 //y=0.54 //x2=50.63 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.545 //y=0.54 //x2=50.145 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=49.66 //y=1.505 //x2=49.66 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=49.66 //y=1.505 //x2=49.66 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=49.66 //y=0.625 //x2=49.66 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=49.66 //y=0.625 //x2=49.66 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=48.775 //y=1.59 //x2=48.69 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=48.775 //y=1.59 //x2=49.175 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.575 //y=1.59 //x2=49.66 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.575 //y=1.59 //x2=49.175 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=48.69 //y=1.505 //x2=48.69 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=48.69 //y=1.505 //x2=48.69 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_49

subckt PM_TMRDFFSNRNQX1\%noxref_50 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=51.065 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=49.96 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=51.2 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=52.17 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=52.085 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=51.2 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=51.115 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=52.17 //y=0.625 //x2=52.17 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=52.17 //y=0.625 //x2=52.17 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=51.285 //y=0.54 //x2=51.2 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=51.285 //y=0.54 //x2=51.685 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=52.085 //y=0.54 //x2=52.17 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=52.085 //y=0.54 //x2=51.685 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=51.2 //y=1.08 //x2=51.2 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=51.2 //y=1.08 //x2=51.2 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=51.2 //y=0.91 //x2=51.2 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=51.2 //y=0.91 //x2=51.2 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=51.2 //y=0.625 //x2=51.2 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=51.2 //y=0.625 //x2=51.2 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.235 //y=0.995 //x2=50.15 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=51.115 //y=0.995 //x2=51.2 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=51.115 //y=0.995 //x2=50.235 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_50

subckt PM_TMRDFFSNRNQX1\%noxref_51 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=53.365 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=55.355 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=55.355 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=54.47 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=54.385 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=53.5 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=54.555 //y=1.59 //x2=54.47 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.555 //y=1.59 //x2=54.955 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.355 //y=1.59 //x2=55.44 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=55.355 //y=1.59 //x2=54.955 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=54.555 //y=0.54 //x2=54.47 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.555 //y=0.54 //x2=54.955 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.355 //y=0.54 //x2=55.44 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=55.355 //y=0.54 //x2=54.955 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=54.47 //y=1.505 //x2=54.47 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=54.47 //y=1.505 //x2=54.47 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=54.47 //y=0.625 //x2=54.47 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=54.47 //y=0.625 //x2=54.47 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.585 //y=1.59 //x2=53.5 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.585 //y=1.59 //x2=53.985 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=54.385 //y=1.59 //x2=54.47 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.385 //y=1.59 //x2=53.985 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=53.5 //y=1.505 //x2=53.5 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=53.5 //y=1.505 //x2=53.5 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_51

subckt PM_TMRDFFSNRNQX1\%noxref_52 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=55.875 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=54.77 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=56.01 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=56.98 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=56.895 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=56.01 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=55.925 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=56.98 //y=0.625 //x2=56.98 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=56.98 //y=0.625 //x2=56.98 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=56.095 //y=0.54 //x2=56.01 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=56.095 //y=0.54 //x2=56.495 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=56.895 //y=0.54 //x2=56.98 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=56.895 //y=0.54 //x2=56.495 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=56.01 //y=1.08 //x2=56.01 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=56.01 //y=1.08 //x2=56.01 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=56.01 //y=0.91 //x2=56.01 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=56.01 //y=0.91 //x2=56.01 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=56.01 //y=0.625 //x2=56.01 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=56.01 //y=0.625 //x2=56.01 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.045 //y=0.995 //x2=54.96 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=55.925 //y=0.995 //x2=56.01 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=55.925 //y=0.995 //x2=55.045 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_52

subckt PM_TMRDFFSNRNQX1\%noxref_53 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=58.175 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=60.165 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=60.165 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=59.28 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=59.195 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=58.31 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=59.365 //y=1.59 //x2=59.28 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.365 //y=1.59 //x2=59.765 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.165 //y=1.59 //x2=60.25 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.165 //y=1.59 //x2=59.765 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=59.365 //y=0.54 //x2=59.28 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.365 //y=0.54 //x2=59.765 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.165 //y=0.54 //x2=60.25 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.165 //y=0.54 //x2=59.765 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=59.28 //y=1.505 //x2=59.28 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=59.28 //y=1.505 //x2=59.28 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=59.28 //y=0.625 //x2=59.28 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=59.28 //y=0.625 //x2=59.28 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.395 //y=1.59 //x2=58.31 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.395 //y=1.59 //x2=58.795 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=59.195 //y=1.59 //x2=59.28 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.195 //y=1.59 //x2=58.795 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=58.31 //y=1.505 //x2=58.31 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=58.31 //y=1.505 //x2=58.31 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_53

subckt PM_TMRDFFSNRNQX1\%noxref_54 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=60.685 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=59.58 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=60.82 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=61.79 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=61.705 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=60.82 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=60.735 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=61.79 //y=0.625 //x2=61.79 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=61.79 //y=0.625 //x2=61.79 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=60.905 //y=0.54 //x2=60.82 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.905 //y=0.54 //x2=61.305 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=61.705 //y=0.54 //x2=61.79 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=61.705 //y=0.54 //x2=61.305 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.82 //y=1.08 //x2=60.82 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=60.82 //y=1.08 //x2=60.82 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.82 //y=0.91 //x2=60.82 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=60.82 //y=0.91 //x2=60.82 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=60.82 //y=0.625 //x2=60.82 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=60.82 //y=0.625 //x2=60.82 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.855 //y=0.995 //x2=59.77 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.735 //y=0.995 //x2=60.82 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=60.735 //y=0.995 //x2=59.855 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_54

subckt PM_TMRDFFSNRNQX1\%noxref_55 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=62.985 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=64.975 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=64.975 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=64.09 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=64.005 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=63.12 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=64.175 //y=1.59 //x2=64.09 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.175 //y=1.59 //x2=64.575 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.975 //y=1.59 //x2=65.06 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.975 //y=1.59 //x2=64.575 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=64.175 //y=0.54 //x2=64.09 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.175 //y=0.54 //x2=64.575 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.975 //y=0.54 //x2=65.06 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.975 //y=0.54 //x2=64.575 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=64.09 //y=1.505 //x2=64.09 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=64.09 //y=1.505 //x2=64.09 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=64.09 //y=0.625 //x2=64.09 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=64.09 //y=0.625 //x2=64.09 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63.205 //y=1.59 //x2=63.12 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63.205 //y=1.59 //x2=63.605 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=64.005 //y=1.59 //x2=64.09 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.005 //y=1.59 //x2=63.605 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=63.12 //y=1.505 //x2=63.12 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=63.12 //y=1.505 //x2=63.12 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_55

subckt PM_TMRDFFSNRNQX1\%noxref_56 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=65.495 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=64.39 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=65.63 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=66.6 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=66.515 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=65.63 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=65.545 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=66.6 //y=0.625 //x2=66.6 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=66.6 //y=0.625 //x2=66.6 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=65.715 //y=0.54 //x2=65.63 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=65.715 //y=0.54 //x2=66.115 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.515 //y=0.54 //x2=66.6 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=66.515 //y=0.54 //x2=66.115 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=65.63 //y=1.08 //x2=65.63 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=65.63 //y=1.08 //x2=65.63 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=65.63 //y=0.91 //x2=65.63 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=65.63 //y=0.91 //x2=65.63 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=65.63 //y=0.625 //x2=65.63 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=65.63 //y=0.625 //x2=65.63 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.665 //y=0.995 //x2=64.58 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=65.545 //y=0.995 //x2=65.63 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=65.545 //y=0.995 //x2=64.665 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_56

subckt PM_TMRDFFSNRNQX1\%noxref_57 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=67.795 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=69.785 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=69.785 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=68.9 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=68.815 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=67.93 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.985 //y=1.59 //x2=68.9 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.985 //y=1.59 //x2=69.385 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.785 //y=1.59 //x2=69.87 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.785 //y=1.59 //x2=69.385 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.985 //y=0.54 //x2=68.9 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.985 //y=0.54 //x2=69.385 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.785 //y=0.54 //x2=69.87 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.785 //y=0.54 //x2=69.385 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=68.9 //y=1.505 //x2=68.9 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=68.9 //y=1.505 //x2=68.9 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=68.9 //y=0.625 //x2=68.9 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=68.9 //y=0.625 //x2=68.9 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.015 //y=1.59 //x2=67.93 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.015 //y=1.59 //x2=68.415 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.815 //y=1.59 //x2=68.9 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.815 //y=1.59 //x2=68.415 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=67.93 //y=1.505 //x2=67.93 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=67.93 //y=1.505 //x2=67.93 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_57

subckt PM_TMRDFFSNRNQX1\%noxref_58 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=70.305 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=69.2 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=70.44 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=71.41 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=71.325 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=70.44 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=70.355 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=71.41 //y=0.625 //x2=71.41 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=71.41 //y=0.625 //x2=71.41 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=70.525 //y=0.54 //x2=70.44 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.525 //y=0.54 //x2=70.925 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=71.325 //y=0.54 //x2=71.41 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=71.325 //y=0.54 //x2=70.925 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=70.44 //y=1.08 //x2=70.44 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=70.44 //y=1.08 //x2=70.44 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=70.44 //y=0.91 //x2=70.44 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=70.44 //y=0.91 //x2=70.44 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=70.44 //y=0.625 //x2=70.44 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=70.44 //y=0.625 //x2=70.44 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.475 //y=0.995 //x2=69.39 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=70.355 //y=0.995 //x2=70.44 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=70.355 //y=0.995 //x2=69.475 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_58

subckt PM_TMRDFFSNRNQX1\%noxref_59 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=72.605 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=74.595 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=74.595 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=73.71 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=73.625 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=72.74 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=73.795 //y=1.59 //x2=73.71 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=73.795 //y=1.59 //x2=74.195 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.595 //y=1.59 //x2=74.68 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=74.595 //y=1.59 //x2=74.195 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=73.795 //y=0.54 //x2=73.71 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=73.795 //y=0.54 //x2=74.195 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.595 //y=0.54 //x2=74.68 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=74.595 //y=0.54 //x2=74.195 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=73.71 //y=1.505 //x2=73.71 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=73.71 //y=1.505 //x2=73.71 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=73.71 //y=0.625 //x2=73.71 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=73.71 //y=0.625 //x2=73.71 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=72.825 //y=1.59 //x2=72.74 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=72.825 //y=1.59 //x2=73.225 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=73.625 //y=1.59 //x2=73.71 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=73.625 //y=1.59 //x2=73.225 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=72.74 //y=1.505 //x2=72.74 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=72.74 //y=1.505 //x2=72.74 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_59

subckt PM_TMRDFFSNRNQX1\%noxref_60 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=75.115 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=74.01 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=75.25 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=76.22 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=76.135 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=75.25 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=75.165 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=76.22 //y=0.625 //x2=76.22 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=76.22 //y=0.625 //x2=76.22 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.335 //y=0.54 //x2=75.25 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=75.335 //y=0.54 //x2=75.735 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=76.135 //y=0.54 //x2=76.22 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=76.135 //y=0.54 //x2=75.735 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=75.25 //y=1.08 //x2=75.25 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=75.25 //y=1.08 //x2=75.25 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=75.25 //y=0.91 //x2=75.25 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=75.25 //y=0.91 //x2=75.25 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=75.25 //y=0.625 //x2=75.25 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=75.25 //y=0.625 //x2=75.25 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.285 //y=0.995 //x2=74.2 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=75.165 //y=0.995 //x2=75.25 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=75.165 //y=0.995 //x2=74.285 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_60

subckt PM_TMRDFFSNRNQX1\%noxref_61 ( 1 5 9 13 17 35 )
c51 ( 35 0 ) capacitor c=0.0680259f //x=77.415 //y=0.375
c52 ( 17 0 ) capacitor c=0.0180446f //x=79.405 //y=1.59
c53 ( 13 0 ) capacitor c=0.0155283f //x=79.405 //y=0.54
c54 ( 9 0 ) capacitor c=0.00678203f //x=78.52 //y=0.625
c55 ( 5 0 ) capacitor c=0.0164013f //x=78.435 //y=1.59
c56 ( 1 0 ) capacitor c=0.00696517f //x=77.55 //y=1.505
r57 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.605 //y=1.59 //x2=78.52 //y2=1.63
r58 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.605 //y=1.59 //x2=79.005 //y2=1.59
r59 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.405 //y=1.59 //x2=79.49 //y2=1.59
r60 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=79.405 //y=1.59 //x2=79.005 //y2=1.59
r61 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.605 //y=0.54 //x2=78.52 //y2=0.5
r62 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.605 //y=0.54 //x2=79.005 //y2=0.54
r63 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.405 //y=0.54 //x2=79.49 //y2=0.54
r64 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=79.405 //y=0.54 //x2=79.005 //y2=0.54
r65 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=78.52 //y=1.505 //x2=78.52 //y2=1.63
r66 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=78.52 //y=1.505 //x2=78.52 //y2=0.89
r67 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=78.52 //y=0.625 //x2=78.52 //y2=0.5
r68 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=78.52 //y=0.625 //x2=78.52 //y2=0.89
r69 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=77.635 //y=1.59 //x2=77.55 //y2=1.63
r70 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=77.635 //y=1.59 //x2=78.035 //y2=1.59
r71 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.435 //y=1.59 //x2=78.52 //y2=1.63
r72 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.435 //y=1.59 //x2=78.035 //y2=1.59
r73 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=77.55 //y=1.505 //x2=77.55 //y2=1.63
r74 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=77.55 //y=1.505 //x2=77.55 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_61

subckt PM_TMRDFFSNRNQX1\%noxref_62 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0421259f //x=79.925 //y=0.375
c54 ( 28 0 ) capacitor c=0.00457437f //x=78.82 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=80.06 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=81.03 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=80.945 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=80.06 //y=0.625
c59 ( 1 0 ) capacitor c=0.0234159f //x=79.975 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=81.03 //y=0.625 //x2=81.03 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=81.03 //y=0.625 //x2=81.03 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=80.145 //y=0.54 //x2=80.06 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=80.145 //y=0.54 //x2=80.545 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=80.945 //y=0.54 //x2=81.03 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=80.945 //y=0.54 //x2=80.545 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=80.06 //y=1.08 //x2=80.06 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=80.06 //y=1.08 //x2=80.06 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=80.06 //y=0.91 //x2=80.06 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=80.06 //y=0.91 //x2=80.06 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=80.06 //y=0.625 //x2=80.06 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=80.06 //y=0.625 //x2=80.06 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.095 //y=0.995 //x2=79.01 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=79.975 //y=0.995 //x2=80.06 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=79.975 //y=0.995 //x2=79.095 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_62

subckt PM_TMRDFFSNRNQX1\%noxref_63 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=82.225 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=84.215 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=84.215 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=83.33 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=83.245 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=82.36 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=83.415 //y=1.59 //x2=83.33 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=83.415 //y=1.59 //x2=83.815 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.215 //y=1.59 //x2=84.3 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=84.215 //y=1.59 //x2=83.815 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=83.415 //y=0.54 //x2=83.33 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=83.415 //y=0.54 //x2=83.815 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.215 //y=0.54 //x2=84.3 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=84.215 //y=0.54 //x2=83.815 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=83.33 //y=1.505 //x2=83.33 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=83.33 //y=1.505 //x2=83.33 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=83.33 //y=0.625 //x2=83.33 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=83.33 //y=0.625 //x2=83.33 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=82.445 //y=1.59 //x2=82.36 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=82.445 //y=1.59 //x2=82.845 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=83.245 //y=1.59 //x2=83.33 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=83.245 //y=1.59 //x2=82.845 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=82.36 //y=1.505 //x2=82.36 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=82.36 //y=1.505 //x2=82.36 //y2=0.89
ends PM_TMRDFFSNRNQX1\%noxref_63

subckt PM_TMRDFFSNRNQX1\%noxref_64 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0412521f //x=84.735 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=83.63 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=84.87 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=85.84 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144274f //x=85.755 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=84.87 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=84.785 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=85.84 //y=0.625 //x2=85.84 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=85.84 //y=0.625 //x2=85.84 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=84.955 //y=0.54 //x2=84.87 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=84.955 //y=0.54 //x2=85.355 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=85.755 //y=0.54 //x2=85.84 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=85.755 //y=0.54 //x2=85.355 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=84.87 //y=1.08 //x2=84.87 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=84.87 //y=1.08 //x2=84.87 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=84.87 //y=0.91 //x2=84.87 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=84.87 //y=0.91 //x2=84.87 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=84.87 //y=0.625 //x2=84.87 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=84.87 //y=0.625 //x2=84.87 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.905 //y=0.995 //x2=83.82 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=84.785 //y=0.995 //x2=84.87 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=84.785 //y=0.995 //x2=83.905 //y2=0.995
ends PM_TMRDFFSNRNQX1\%noxref_64

subckt PM_TMRDFFSNRNQX1\%noxref_65 ( 1 5 9 10 13 17 29 )
c57 ( 29 0 ) capacitor c=0.0751624f //x=87.14 //y=0.365
c58 ( 17 0 ) capacitor c=0.0072249f //x=89.215 //y=0.615
c59 ( 13 0 ) capacitor c=0.0152499f //x=89.13 //y=0.53
c60 ( 10 0 ) capacitor c=0.00698291f //x=88.245 //y=1.495
c61 ( 9 0 ) capacitor c=0.006761f //x=88.245 //y=0.615
c62 ( 5 0 ) capacitor c=0.0191191f //x=88.16 //y=1.58
c63 ( 1 0 ) capacitor c=0.00483164f //x=87.275 //y=1.495
r64 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=89.215 //y=0.615 //x2=89.215 //y2=0.49
r65 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=89.215 //y=0.615 //x2=89.215 //y2=1.22
r66 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=88.33 //y=0.53 //x2=88.245 //y2=0.49
r67 (  14 29 ) resistor r=27.0374 //w=0.187 //l=0.395 //layer=li \
 //thickness=0.1 //x=88.33 //y=0.53 //x2=88.725 //y2=0.53
r68 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=89.13 //y=0.53 //x2=89.215 //y2=0.49
r69 (  13 29 ) resistor r=27.7219 //w=0.187 //l=0.405 //layer=li \
 //thickness=0.1 //x=89.13 //y=0.53 //x2=88.725 //y2=0.53
r70 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=88.245 //y=1.495 //x2=88.245 //y2=1.62
r71 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=88.245 //y=1.495 //x2=88.245 //y2=0.88
r72 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=88.245 //y=0.615 //x2=88.245 //y2=0.49
r73 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=88.245 //y=0.615 //x2=88.245 //y2=0.88
r74 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=87.36 //y=1.58 //x2=87.275 //y2=1.62
r75 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=87.36 //y=1.58 //x2=87.76 //y2=1.58
r76 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=88.16 //y=1.58 //x2=88.245 //y2=1.62
r77 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=88.16 //y=1.58 //x2=87.76 //y2=1.58
r78 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=87.275 //y=1.495 //x2=87.275 //y2=1.62
r79 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=87.275 //y=1.495 //x2=87.275 //y2=0.88
ends PM_TMRDFFSNRNQX1\%noxref_65

subckt PM_TMRDFFSNRNQX1\%noxref_66 ( 1 5 9 10 13 17 29 )
c55 ( 29 0 ) capacitor c=0.0723103f //x=90.47 //y=0.365
c56 ( 17 0 ) capacitor c=0.0072249f //x=92.545 //y=0.615
c57 ( 13 0 ) capacitor c=0.0155051f //x=92.46 //y=0.53
c58 ( 10 0 ) capacitor c=0.00811719f //x=91.575 //y=1.495
c59 ( 9 0 ) capacitor c=0.006761f //x=91.575 //y=0.615
c60 ( 5 0 ) capacitor c=0.0166789f //x=91.49 //y=1.58
c61 ( 1 0 ) capacitor c=0.00788388f //x=90.605 //y=1.495
r62 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=92.545 //y=0.615 //x2=92.545 //y2=0.49
r63 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=92.545 //y=0.615 //x2=92.545 //y2=1.22
r64 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=91.66 //y=0.53 //x2=91.575 //y2=0.49
r65 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=91.66 //y=0.53 //x2=92.06 //y2=0.53
r66 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=92.46 //y=0.53 //x2=92.545 //y2=0.49
r67 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=92.46 //y=0.53 //x2=92.06 //y2=0.53
r68 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=91.575 //y=1.495 //x2=91.575 //y2=1.62
r69 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=91.575 //y=1.495 //x2=91.575 //y2=0.88
r70 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=91.575 //y=0.615 //x2=91.575 //y2=0.49
r71 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=91.575 //y=0.615 //x2=91.575 //y2=0.88
r72 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=90.69 //y=1.58 //x2=90.605 //y2=1.62
r73 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=90.69 //y=1.58 //x2=91.09 //y2=1.58
r74 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=91.49 //y=1.58 //x2=91.575 //y2=1.62
r75 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=91.49 //y=1.58 //x2=91.09 //y2=1.58
r76 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=90.605 //y=1.495 //x2=90.605 //y2=1.62
r77 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=90.605 //y=1.495 //x2=90.605 //y2=0.88
ends PM_TMRDFFSNRNQX1\%noxref_66

subckt PM_TMRDFFSNRNQX1\%noxref_67 ( 1 5 9 10 13 17 29 )
c56 ( 29 0 ) capacitor c=0.0637832f //x=93.8 //y=0.365
c57 ( 17 0 ) capacitor c=0.00722228f //x=95.875 //y=0.615
c58 ( 13 0 ) capacitor c=0.0141607f //x=95.79 //y=0.53
c59 ( 10 0 ) capacitor c=0.00712138f //x=94.905 //y=1.495
c60 ( 9 0 ) capacitor c=0.006761f //x=94.905 //y=0.615
c61 ( 5 0 ) capacitor c=0.0233454f //x=94.82 //y=1.58
c62 ( 1 0 ) capacitor c=0.00481264f //x=93.935 //y=1.495
r63 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=95.875 //y=0.615 //x2=95.875 //y2=0.49
r64 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=95.875 //y=0.615 //x2=95.875 //y2=0.88
r65 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=94.99 //y=0.53 //x2=94.905 //y2=0.49
r66 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=94.99 //y=0.53 //x2=95.39 //y2=0.53
r67 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=95.79 //y=0.53 //x2=95.875 //y2=0.49
r68 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=95.79 //y=0.53 //x2=95.39 //y2=0.53
r69 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=94.905 //y=1.495 //x2=94.905 //y2=1.62
r70 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=94.905 //y=1.495 //x2=94.905 //y2=0.88
r71 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=94.905 //y=0.615 //x2=94.905 //y2=0.49
r72 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=94.905 //y=0.615 //x2=94.905 //y2=0.88
r73 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=94.02 //y=1.58 //x2=93.935 //y2=1.62
r74 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=94.02 //y=1.58 //x2=94.42 //y2=1.58
r75 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=94.82 //y=1.58 //x2=94.905 //y2=1.62
r76 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=94.82 //y=1.58 //x2=94.42 //y2=1.58
r77 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=93.935 //y=1.495 //x2=93.935 //y2=1.62
r78 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=93.935 //y=1.495 //x2=93.935 //y2=0.88
ends PM_TMRDFFSNRNQX1\%noxref_67

