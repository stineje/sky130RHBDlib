// File: nand3x1_pcell.spi.NAND3X1_PCELL.pxi
// Created: Tue Oct 15 15:57:52 2024
// 
simulator lang=spectre
x_PM_NAND3X1_PCELL\%noxref_2 ( N_noxref_2_c_59_p N_noxref_2_c_27_n \
 N_noxref_2_c_31_p N_noxref_2_c_38_p N_noxref_2_c_43_p N_noxref_2_c_28_n \
 N_noxref_2_M3_noxref_s N_noxref_2_M4_noxref_d N_noxref_2_M6_noxref_d \
 N_noxref_2_M8_noxref_d )  PM_NAND3X1_PCELL\%noxref_2
x_PM_NAND3X1_PCELL\%noxref_3 ( N_noxref_3_c_74_n N_noxref_3_M0_noxref_g \
 N_noxref_3_M3_noxref_g N_noxref_3_M4_noxref_g N_noxref_3_c_75_n \
 N_noxref_3_c_76_n N_noxref_3_c_77_n N_noxref_3_c_78_n N_noxref_3_c_79_n \
 N_noxref_3_c_80_n N_noxref_3_c_81_n N_noxref_3_c_82_n N_noxref_3_c_93_p \
 N_noxref_3_c_89_n )  PM_NAND3X1_PCELL\%noxref_3
x_PM_NAND3X1_PCELL\%noxref_4 ( N_noxref_4_c_126_n N_noxref_4_M1_noxref_g \
 N_noxref_4_M5_noxref_g N_noxref_4_M6_noxref_g N_noxref_4_c_139_n \
 N_noxref_4_c_142_n N_noxref_4_c_183_p N_noxref_4_c_190_p N_noxref_4_c_144_n \
 N_noxref_4_c_145_n N_noxref_4_c_146_n N_noxref_4_c_147_n N_noxref_4_c_173_p \
 N_noxref_4_c_149_n )  PM_NAND3X1_PCELL\%noxref_4
x_PM_NAND3X1_PCELL\%noxref_5 ( N_noxref_5_c_199_n N_noxref_5_c_195_n \
 N_noxref_5_c_196_n N_noxref_5_c_197_n N_noxref_5_c_211_n \
 N_noxref_5_M0_noxref_s )  PM_NAND3X1_PCELL\%noxref_5
x_PM_NAND3X1_PCELL\%noxref_6 ( N_noxref_6_c_226_n N_noxref_6_M2_noxref_g \
 N_noxref_6_M7_noxref_g N_noxref_6_M8_noxref_g N_noxref_6_c_239_n \
 N_noxref_6_c_240_n N_noxref_6_c_241_n N_noxref_6_c_262_p N_noxref_6_c_251_p \
 N_noxref_6_c_264_p N_noxref_6_c_252_p N_noxref_6_c_242_n N_noxref_6_c_244_n \
 N_noxref_6_c_245_n )  PM_NAND3X1_PCELL\%noxref_6
x_PM_NAND3X1_PCELL\%noxref_7 ( N_noxref_7_c_280_n N_noxref_7_c_283_n \
 N_noxref_7_c_285_n N_noxref_7_c_288_n N_noxref_7_c_278_n N_noxref_7_c_343_p \
 N_noxref_7_c_291_n N_noxref_7_c_316_n N_noxref_7_c_329_n \
 N_noxref_7_M2_noxref_d N_noxref_7_M3_noxref_d N_noxref_7_M5_noxref_d \
 N_noxref_7_M7_noxref_d )  PM_NAND3X1_PCELL\%noxref_7
x_PM_NAND3X1_PCELL\%noxref_8 ( N_noxref_8_c_347_n N_noxref_8_c_348_n \
 N_noxref_8_c_349_n N_noxref_8_c_350_n N_noxref_8_c_377_n \
 N_noxref_8_M1_noxref_d N_noxref_8_M2_noxref_s )  PM_NAND3X1_PCELL\%noxref_8
cc_1 ( noxref_1 N_noxref_2_c_27_n ) capacitor c=0.00989031f //x=0.885 \
 //y=0.875 //x2=0.74 //y2=7.4
cc_2 ( noxref_1 N_noxref_2_c_28_n ) capacitor c=0.00989031f //x=0.885 \
 //y=0.875 //x2=4.07 //y2=7.4
cc_3 ( noxref_1 N_noxref_3_c_74_n ) capacitor c=0.0180363f //x=0.885 //y=0.875 \
 //x2=1.11 //y2=2.08
cc_4 ( noxref_1 N_noxref_3_c_75_n ) capacitor c=0.00344751f //x=0.885 \
 //y=0.875 //x2=0.81 //y2=0.875
cc_5 ( noxref_1 N_noxref_3_c_76_n ) capacitor c=0.00255985f //x=0.885 \
 //y=0.875 //x2=0.81 //y2=1.22
cc_6 ( noxref_1 N_noxref_3_c_77_n ) capacitor c=0.00295461f //x=0.885 \
 //y=0.875 //x2=0.81 //y2=1.53
cc_7 ( noxref_1 N_noxref_3_c_78_n ) capacitor c=0.0134214f //x=0.885 //y=0.875 \
 //x2=0.81 //y2=1.915
cc_8 ( noxref_1 N_noxref_3_c_79_n ) capacitor c=0.0131341f //x=0.885 //y=0.875 \
 //x2=1.185 //y2=0.72
cc_9 ( noxref_1 N_noxref_3_c_80_n ) capacitor c=0.00193146f //x=0.885 \
 //y=0.875 //x2=1.185 //y2=1.375
cc_10 ( noxref_1 N_noxref_3_c_81_n ) capacitor c=0.00386866f //x=0.885 \
 //y=0.875 //x2=1.34 //y2=0.875
cc_11 ( noxref_1 N_noxref_3_c_82_n ) capacitor c=0.00255985f //x=0.885 \
 //y=0.875 //x2=1.34 //y2=1.22
cc_12 ( noxref_1 N_noxref_4_c_126_n ) capacitor c=7.64246e-19 //x=0.885 \
 //y=0.875 //x2=2.22 //y2=2.08
cc_13 ( noxref_1 N_noxref_5_c_195_n ) capacitor c=0.0189984f //x=0.885 \
 //y=0.875 //x2=1.475 //y2=1.59
cc_14 ( noxref_1 N_noxref_5_c_196_n ) capacitor c=0.0564515f //x=0.885 \
 //y=0.875 //x2=1.56 //y2=0.625
cc_15 ( noxref_1 N_noxref_5_c_197_n ) capacitor c=0.0574584f //x=0.885 \
 //y=0.875 //x2=2.445 //y2=0.54
cc_16 ( noxref_1 N_noxref_5_M0_noxref_s ) capacitor c=0.14912f //x=0.885 \
 //y=0.875 //x2=0.455 //y2=0.375
cc_17 ( noxref_1 N_noxref_6_c_226_n ) capacitor c=9.53263e-19 //x=0.885 \
 //y=0.875 //x2=3.33 //y2=2.08
cc_18 ( noxref_1 N_noxref_7_c_278_n ) capacitor c=0.0465819f //x=0.885 \
 //y=0.875 //x2=3.985 //y2=1.665
cc_19 ( noxref_1 N_noxref_7_M2_noxref_d ) capacitor c=0.00593061f //x=0.885 \
 //y=0.875 //x2=3.395 //y2=0.915
cc_20 ( noxref_1 N_noxref_8_c_347_n ) capacitor c=0.0165482f //x=0.885 \
 //y=0.875 //x2=3.015 //y2=0.995
cc_21 ( noxref_1 N_noxref_8_c_348_n ) capacitor c=0.0231189f //x=0.885 \
 //y=0.875 //x2=3.1 //y2=0.625
cc_22 ( noxref_1 N_noxref_8_c_349_n ) capacitor c=0.0584577f //x=0.885 \
 //y=0.875 //x2=3.985 //y2=0.54
cc_23 ( noxref_1 N_noxref_8_c_350_n ) capacitor c=0.0633375f //x=0.885 \
 //y=0.875 //x2=4.07 //y2=0.625
cc_24 ( noxref_1 N_noxref_8_M1_noxref_d ) capacitor c=0.00162435f //x=0.885 \
 //y=0.875 //x2=1.86 //y2=0.91
cc_25 ( noxref_1 N_noxref_8_M2_noxref_s ) capacitor c=0.00265212f //x=0.885 \
 //y=0.875 //x2=2.965 //y2=0.375
cc_26 ( N_noxref_2_c_27_n N_noxref_3_c_74_n ) capacitor c=0.0168497f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_27 ( N_noxref_2_M3_noxref_s N_noxref_3_c_74_n ) capacitor c=0.0128617f \
 //x=0.955 //y=5.02 //x2=1.11 //y2=2.08
cc_28 ( N_noxref_2_c_31_p N_noxref_3_M3_noxref_g ) capacitor c=0.00749687f \
 //x=1.885 //y=7.4 //x2=1.31 //y2=6.02
cc_29 ( N_noxref_2_M3_noxref_s N_noxref_3_M3_noxref_g ) capacitor c=0.0477201f \
 //x=0.955 //y=5.02 //x2=1.31 //y2=6.02
cc_30 ( N_noxref_2_c_31_p N_noxref_3_M4_noxref_g ) capacitor c=0.00675175f \
 //x=1.885 //y=7.4 //x2=1.75 //y2=6.02
cc_31 ( N_noxref_2_M4_noxref_d N_noxref_3_M4_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=1.75 //y2=6.02
cc_32 ( N_noxref_2_c_27_n N_noxref_3_c_89_n ) capacitor c=0.0076931f //x=0.74 \
 //y=7.4 //x2=1.385 //y2=4.79
cc_33 ( N_noxref_2_M3_noxref_s N_noxref_3_c_89_n ) capacitor c=0.00637187f \
 //x=0.955 //y=5.02 //x2=1.385 //y2=4.79
cc_34 ( N_noxref_2_c_27_n N_noxref_4_c_126_n ) capacitor c=7.34553e-19 \
 //x=0.74 //y=7.4 //x2=2.22 //y2=2.08
cc_35 ( N_noxref_2_c_38_p N_noxref_4_M5_noxref_g ) capacitor c=0.00676195f \
 //x=2.765 //y=7.4 //x2=2.19 //y2=6.02
cc_36 ( N_noxref_2_M4_noxref_d N_noxref_4_M5_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=2.19 //y2=6.02
cc_37 ( N_noxref_2_c_38_p N_noxref_4_M6_noxref_g ) capacitor c=0.00675175f \
 //x=2.765 //y=7.4 //x2=2.63 //y2=6.02
cc_38 ( N_noxref_2_M6_noxref_d N_noxref_4_M6_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=2.63 //y2=6.02
cc_39 ( N_noxref_2_c_28_n N_noxref_6_c_226_n ) capacitor c=8.81482e-19 \
 //x=4.07 //y=7.4 //x2=3.33 //y2=2.08
cc_40 ( N_noxref_2_c_43_p N_noxref_6_M7_noxref_g ) capacitor c=0.00675175f \
 //x=3.645 //y=7.4 //x2=3.07 //y2=6.02
cc_41 ( N_noxref_2_M6_noxref_d N_noxref_6_M7_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=3.07 //y2=6.02
cc_42 ( N_noxref_2_c_43_p N_noxref_6_M8_noxref_g ) capacitor c=0.00675379f \
 //x=3.645 //y=7.4 //x2=3.51 //y2=6.02
cc_43 ( N_noxref_2_M8_noxref_d N_noxref_6_M8_noxref_g ) capacitor c=0.0394719f \
 //x=3.585 //y=5.02 //x2=3.51 //y2=6.02
cc_44 ( N_noxref_2_c_31_p N_noxref_7_c_280_n ) capacitor c=5.56103e-19 \
 //x=1.885 //y=7.4 //x2=2.325 //y2=5.155
cc_45 ( N_noxref_2_c_38_p N_noxref_7_c_280_n ) capacitor c=5.56103e-19 \
 //x=2.765 //y=7.4 //x2=2.325 //y2=5.155
cc_46 ( N_noxref_2_M4_noxref_d N_noxref_7_c_280_n ) capacitor c=0.0120385f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_47 ( N_noxref_2_c_27_n N_noxref_7_c_283_n ) capacitor c=0.00880189f \
 //x=0.74 //y=7.4 //x2=1.615 //y2=5.155
cc_48 ( N_noxref_2_M3_noxref_s N_noxref_7_c_283_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_49 ( N_noxref_2_c_38_p N_noxref_7_c_285_n ) capacitor c=5.56103e-19 \
 //x=2.765 //y=7.4 //x2=3.205 //y2=5.155
cc_50 ( N_noxref_2_c_43_p N_noxref_7_c_285_n ) capacitor c=5.56103e-19 \
 //x=3.645 //y=7.4 //x2=3.205 //y2=5.155
cc_51 ( N_noxref_2_M6_noxref_d N_noxref_7_c_285_n ) capacitor c=0.0120385f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_52 ( N_noxref_2_c_43_p N_noxref_7_c_288_n ) capacitor c=8.43508e-19 \
 //x=3.645 //y=7.4 //x2=3.985 //y2=5.155
cc_53 ( N_noxref_2_c_28_n N_noxref_7_c_288_n ) capacitor c=0.00184483f \
 //x=4.07 //y=7.4 //x2=3.985 //y2=5.155
cc_54 ( N_noxref_2_M8_noxref_d N_noxref_7_c_288_n ) capacitor c=0.0120385f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_55 ( N_noxref_2_c_28_n N_noxref_7_c_291_n ) capacitor c=0.046173f //x=4.07 \
 //y=7.4 //x2=4.07 //y2=5.07
cc_56 ( N_noxref_2_c_59_p N_noxref_7_M3_noxref_d ) capacitor c=0.00719816f \
 //x=4.07 //y=7.4 //x2=1.385 //y2=5.02
cc_57 ( N_noxref_2_c_31_p N_noxref_7_M3_noxref_d ) capacitor c=0.0138437f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_58 ( N_noxref_2_c_28_n N_noxref_7_M3_noxref_d ) capacitor c=0.00135292f \
 //x=4.07 //y=7.4 //x2=1.385 //y2=5.02
cc_59 ( N_noxref_2_M4_noxref_d N_noxref_7_M3_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_60 ( N_noxref_2_c_59_p N_noxref_7_M5_noxref_d ) capacitor c=0.00719816f \
 //x=4.07 //y=7.4 //x2=2.265 //y2=5.02
cc_61 ( N_noxref_2_c_38_p N_noxref_7_M5_noxref_d ) capacitor c=0.0138437f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_62 ( N_noxref_2_c_28_n N_noxref_7_M5_noxref_d ) capacitor c=0.00184577f \
 //x=4.07 //y=7.4 //x2=2.265 //y2=5.02
cc_63 ( N_noxref_2_M3_noxref_s N_noxref_7_M5_noxref_d ) capacitor \
 c=0.00130656f //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_64 ( N_noxref_2_M4_noxref_d N_noxref_7_M5_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_65 ( N_noxref_2_M6_noxref_d N_noxref_7_M5_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_66 ( N_noxref_2_c_59_p N_noxref_7_M7_noxref_d ) capacitor c=0.00719816f \
 //x=4.07 //y=7.4 //x2=3.145 //y2=5.02
cc_67 ( N_noxref_2_c_43_p N_noxref_7_M7_noxref_d ) capacitor c=0.0137718f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_68 ( N_noxref_2_c_28_n N_noxref_7_M7_noxref_d ) capacitor c=0.010988f \
 //x=4.07 //y=7.4 //x2=3.145 //y2=5.02
cc_69 ( N_noxref_2_M6_noxref_d N_noxref_7_M7_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_70 ( N_noxref_2_M8_noxref_d N_noxref_7_M7_noxref_d ) capacitor c=0.0664752f \
 //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_71 ( N_noxref_3_c_74_n N_noxref_4_c_126_n ) capacitor c=0.0587479f //x=1.11 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_72 ( N_noxref_3_c_78_n N_noxref_4_c_126_n ) capacitor c=0.00238338f \
 //x=0.81 //y=1.915 //x2=2.22 //y2=2.08
cc_73 ( N_noxref_3_c_93_p N_noxref_4_c_126_n ) capacitor c=0.00147352f \
 //x=1.675 //y=4.79 //x2=2.22 //y2=2.08
cc_74 ( N_noxref_3_c_89_n N_noxref_4_c_126_n ) capacitor c=0.00142741f \
 //x=1.385 //y=4.79 //x2=2.22 //y2=2.08
cc_75 ( N_noxref_3_M3_noxref_g N_noxref_4_M5_noxref_g ) capacitor c=0.0105869f \
 //x=1.31 //y=6.02 //x2=2.19 //y2=6.02
cc_76 ( N_noxref_3_M4_noxref_g N_noxref_4_M5_noxref_g ) capacitor c=0.10632f \
 //x=1.75 //y=6.02 //x2=2.19 //y2=6.02
cc_77 ( N_noxref_3_M4_noxref_g N_noxref_4_M6_noxref_g ) capacitor c=0.0101598f \
 //x=1.75 //y=6.02 //x2=2.63 //y2=6.02
cc_78 ( N_noxref_3_c_75_n N_noxref_4_c_139_n ) capacitor c=5.72482e-19 \
 //x=0.81 //y=0.875 //x2=1.785 //y2=0.91
cc_79 ( N_noxref_3_c_76_n N_noxref_4_c_139_n ) capacitor c=0.00149976f \
 //x=0.81 //y=1.22 //x2=1.785 //y2=0.91
cc_80 ( N_noxref_3_c_81_n N_noxref_4_c_139_n ) capacitor c=0.0160123f //x=1.34 \
 //y=0.875 //x2=1.785 //y2=0.91
cc_81 ( N_noxref_3_c_77_n N_noxref_4_c_142_n ) capacitor c=0.00111227f \
 //x=0.81 //y=1.53 //x2=1.785 //y2=1.22
cc_82 ( N_noxref_3_c_82_n N_noxref_4_c_142_n ) capacitor c=0.0124075f //x=1.34 \
 //y=1.22 //x2=1.785 //y2=1.22
cc_83 ( N_noxref_3_c_81_n N_noxref_4_c_144_n ) capacitor c=0.00103227f \
 //x=1.34 //y=0.875 //x2=2.31 //y2=0.91
cc_84 ( N_noxref_3_c_82_n N_noxref_4_c_145_n ) capacitor c=0.0010154f //x=1.34 \
 //y=1.22 //x2=2.31 //y2=1.22
cc_85 ( N_noxref_3_c_82_n N_noxref_4_c_146_n ) capacitor c=9.23422e-19 \
 //x=1.34 //y=1.22 //x2=2.31 //y2=1.45
cc_86 ( N_noxref_3_c_74_n N_noxref_4_c_147_n ) capacitor c=0.00231304f \
 //x=1.11 //y=2.08 //x2=2.31 //y2=1.915
cc_87 ( N_noxref_3_c_78_n N_noxref_4_c_147_n ) capacitor c=0.00964411f \
 //x=0.81 //y=1.915 //x2=2.31 //y2=1.915
cc_88 ( N_noxref_3_c_74_n N_noxref_4_c_149_n ) capacitor c=0.00183762f \
 //x=1.11 //y=2.08 //x2=2.22 //y2=4.7
cc_89 ( N_noxref_3_c_93_p N_noxref_4_c_149_n ) capacitor c=0.0168581f \
 //x=1.675 //y=4.79 //x2=2.22 //y2=4.7
cc_90 ( N_noxref_3_c_89_n N_noxref_4_c_149_n ) capacitor c=0.00484466f \
 //x=1.385 //y=4.79 //x2=2.22 //y2=4.7
cc_91 ( N_noxref_3_c_78_n N_noxref_5_c_199_n ) capacitor c=0.0034165f //x=0.81 \
 //y=1.915 //x2=0.59 //y2=1.505
cc_92 ( N_noxref_3_c_74_n N_noxref_5_c_195_n ) capacitor c=0.0122915f //x=1.11 \
 //y=2.08 //x2=1.475 //y2=1.59
cc_93 ( N_noxref_3_c_77_n N_noxref_5_c_195_n ) capacitor c=0.00703864f \
 //x=0.81 //y=1.53 //x2=1.475 //y2=1.59
cc_94 ( N_noxref_3_c_78_n N_noxref_5_c_195_n ) capacitor c=0.0259045f //x=0.81 \
 //y=1.915 //x2=1.475 //y2=1.59
cc_95 ( N_noxref_3_c_80_n N_noxref_5_c_195_n ) capacitor c=0.00708583f \
 //x=1.185 //y=1.375 //x2=1.475 //y2=1.59
cc_96 ( N_noxref_3_c_82_n N_noxref_5_c_195_n ) capacitor c=0.00698822f \
 //x=1.34 //y=1.22 //x2=1.475 //y2=1.59
cc_97 ( N_noxref_3_c_75_n N_noxref_5_M0_noxref_s ) capacitor c=0.0327271f \
 //x=0.81 //y=0.875 //x2=0.455 //y2=0.375
cc_98 ( N_noxref_3_c_77_n N_noxref_5_M0_noxref_s ) capacitor c=7.99997e-19 \
 //x=0.81 //y=1.53 //x2=0.455 //y2=0.375
cc_99 ( N_noxref_3_c_78_n N_noxref_5_M0_noxref_s ) capacitor c=0.00122123f \
 //x=0.81 //y=1.915 //x2=0.455 //y2=0.375
cc_100 ( N_noxref_3_c_81_n N_noxref_5_M0_noxref_s ) capacitor c=0.0121427f \
 //x=1.34 //y=0.875 //x2=0.455 //y2=0.375
cc_101 ( N_noxref_3_c_74_n N_noxref_6_c_226_n ) capacitor c=0.00135364f \
 //x=1.11 //y=2.08 //x2=3.33 //y2=2.08
cc_102 ( N_noxref_3_M4_noxref_g N_noxref_7_c_280_n ) capacitor c=0.0204345f \
 //x=1.75 //y=6.02 //x2=2.325 //y2=5.155
cc_103 ( N_noxref_3_M3_noxref_g N_noxref_7_c_283_n ) capacitor c=0.0213876f \
 //x=1.31 //y=6.02 //x2=1.615 //y2=5.155
cc_104 ( N_noxref_3_c_93_p N_noxref_7_c_283_n ) capacitor c=0.0044314f \
 //x=1.675 //y=4.79 //x2=1.615 //y2=5.155
cc_105 ( N_noxref_3_M4_noxref_g N_noxref_7_M3_noxref_d ) capacitor \
 c=0.0180032f //x=1.75 //y=6.02 //x2=1.385 //y2=5.02
cc_106 ( N_noxref_4_c_139_n N_noxref_5_c_197_n ) capacitor c=0.0167228f \
 //x=1.785 //y=0.91 //x2=2.445 //y2=0.54
cc_107 ( N_noxref_4_c_144_n N_noxref_5_c_197_n ) capacitor c=0.00534519f \
 //x=2.31 //y=0.91 //x2=2.445 //y2=0.54
cc_108 ( N_noxref_4_c_126_n N_noxref_5_c_211_n ) capacitor c=0.0124072f \
 //x=2.22 //y=2.08 //x2=2.445 //y2=1.59
cc_109 ( N_noxref_4_c_142_n N_noxref_5_c_211_n ) capacitor c=0.0153476f \
 //x=1.785 //y=1.22 //x2=2.445 //y2=1.59
cc_110 ( N_noxref_4_c_147_n N_noxref_5_c_211_n ) capacitor c=0.023396f \
 //x=2.31 //y=1.915 //x2=2.445 //y2=1.59
cc_111 ( N_noxref_4_c_139_n N_noxref_5_M0_noxref_s ) capacitor c=0.00798959f \
 //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_112 ( N_noxref_4_c_146_n N_noxref_5_M0_noxref_s ) capacitor c=0.00212176f \
 //x=2.31 //y=1.45 //x2=0.455 //y2=0.375
cc_113 ( N_noxref_4_c_147_n N_noxref_5_M0_noxref_s ) capacitor c=0.00298115f \
 //x=2.31 //y=1.915 //x2=0.455 //y2=0.375
cc_114 ( N_noxref_4_c_126_n N_noxref_6_c_226_n ) capacitor c=0.0585754f \
 //x=2.22 //y=2.08 //x2=3.33 //y2=2.08
cc_115 ( N_noxref_4_c_147_n N_noxref_6_c_226_n ) capacitor c=0.0023343f \
 //x=2.31 //y=1.915 //x2=3.33 //y2=2.08
cc_116 ( N_noxref_4_c_149_n N_noxref_6_c_226_n ) capacitor c=0.00142741f \
 //x=2.22 //y=4.7 //x2=3.33 //y2=2.08
cc_117 ( N_noxref_4_M5_noxref_g N_noxref_6_M7_noxref_g ) capacitor \
 c=0.0101598f //x=2.19 //y=6.02 //x2=3.07 //y2=6.02
cc_118 ( N_noxref_4_M6_noxref_g N_noxref_6_M7_noxref_g ) capacitor \
 c=0.0602553f //x=2.63 //y=6.02 //x2=3.07 //y2=6.02
cc_119 ( N_noxref_4_M6_noxref_g N_noxref_6_M8_noxref_g ) capacitor \
 c=0.0101598f //x=2.63 //y=6.02 //x2=3.51 //y2=6.02
cc_120 ( N_noxref_4_c_144_n N_noxref_6_c_239_n ) capacitor c=0.00456962f \
 //x=2.31 //y=0.91 //x2=3.32 //y2=0.915
cc_121 ( N_noxref_4_c_145_n N_noxref_6_c_240_n ) capacitor c=0.00438372f \
 //x=2.31 //y=1.22 //x2=3.32 //y2=1.26
cc_122 ( N_noxref_4_c_146_n N_noxref_6_c_241_n ) capacitor c=0.00438372f \
 //x=2.31 //y=1.45 //x2=3.32 //y2=1.57
cc_123 ( N_noxref_4_c_126_n N_noxref_6_c_242_n ) capacitor c=0.00228632f \
 //x=2.22 //y=2.08 //x2=3.33 //y2=2.08
cc_124 ( N_noxref_4_c_147_n N_noxref_6_c_242_n ) capacitor c=0.00933826f \
 //x=2.31 //y=1.915 //x2=3.33 //y2=2.08
cc_125 ( N_noxref_4_c_147_n N_noxref_6_c_244_n ) capacitor c=0.00438372f \
 //x=2.31 //y=1.915 //x2=3.33 //y2=1.915
cc_126 ( N_noxref_4_c_126_n N_noxref_6_c_245_n ) capacitor c=0.00219458f \
 //x=2.22 //y=2.08 //x2=3.33 //y2=4.7
cc_127 ( N_noxref_4_c_173_p N_noxref_6_c_245_n ) capacitor c=0.0611812f \
 //x=2.555 //y=4.79 //x2=3.33 //y2=4.7
cc_128 ( N_noxref_4_c_149_n N_noxref_6_c_245_n ) capacitor c=0.00487508f \
 //x=2.22 //y=4.7 //x2=3.33 //y2=4.7
cc_129 ( N_noxref_4_c_126_n N_noxref_7_c_280_n ) capacitor c=0.0147127f \
 //x=2.22 //y=2.08 //x2=2.325 //y2=5.155
cc_130 ( N_noxref_4_M5_noxref_g N_noxref_7_c_280_n ) capacitor c=0.0170309f \
 //x=2.19 //y=6.02 //x2=2.325 //y2=5.155
cc_131 ( N_noxref_4_c_149_n N_noxref_7_c_280_n ) capacitor c=0.00325274f \
 //x=2.22 //y=4.7 //x2=2.325 //y2=5.155
cc_132 ( N_noxref_4_M6_noxref_g N_noxref_7_c_285_n ) capacitor c=0.0209597f \
 //x=2.63 //y=6.02 //x2=3.205 //y2=5.155
cc_133 ( N_noxref_4_c_126_n N_noxref_7_c_291_n ) capacitor c=0.003217f \
 //x=2.22 //y=2.08 //x2=4.07 //y2=5.07
cc_134 ( N_noxref_4_c_173_p N_noxref_7_c_316_n ) capacitor c=0.00441288f \
 //x=2.555 //y=4.79 //x2=2.41 //y2=5.155
cc_135 ( N_noxref_4_M5_noxref_g N_noxref_7_M5_noxref_d ) capacitor \
 c=0.0180032f //x=2.19 //y=6.02 //x2=2.265 //y2=5.02
cc_136 ( N_noxref_4_M6_noxref_g N_noxref_7_M5_noxref_d ) capacitor \
 c=0.0180032f //x=2.63 //y=6.02 //x2=2.265 //y2=5.02
cc_137 ( N_noxref_4_c_183_p N_noxref_8_c_347_n ) capacitor c=2.14837e-19 \
 //x=2.155 //y=0.755 //x2=3.015 //y2=0.995
cc_138 ( N_noxref_4_c_144_n N_noxref_8_c_347_n ) capacitor c=0.00123426f \
 //x=2.31 //y=0.91 //x2=3.015 //y2=0.995
cc_139 ( N_noxref_4_c_145_n N_noxref_8_c_347_n ) capacitor c=0.0129288f \
 //x=2.31 //y=1.22 //x2=3.015 //y2=0.995
cc_140 ( N_noxref_4_c_146_n N_noxref_8_c_347_n ) capacitor c=0.00142359f \
 //x=2.31 //y=1.45 //x2=3.015 //y2=0.995
cc_141 ( N_noxref_4_c_139_n N_noxref_8_M1_noxref_d ) capacitor c=0.00223875f \
 //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_142 ( N_noxref_4_c_142_n N_noxref_8_M1_noxref_d ) capacitor c=0.00262485f \
 //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_143 ( N_noxref_4_c_183_p N_noxref_8_M1_noxref_d ) capacitor c=0.00220746f \
 //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_144 ( N_noxref_4_c_190_p N_noxref_8_M1_noxref_d ) capacitor c=0.00194798f \
 //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_145 ( N_noxref_4_c_144_n N_noxref_8_M1_noxref_d ) capacitor c=0.00198465f \
 //x=2.31 //y=0.91 //x2=1.86 //y2=0.91
cc_146 ( N_noxref_4_c_145_n N_noxref_8_M1_noxref_d ) capacitor c=0.00128384f \
 //x=2.31 //y=1.22 //x2=1.86 //y2=0.91
cc_147 ( N_noxref_4_c_144_n N_noxref_8_M2_noxref_s ) capacitor c=7.21316e-19 \
 //x=2.31 //y=0.91 //x2=2.965 //y2=0.375
cc_148 ( N_noxref_4_c_145_n N_noxref_8_M2_noxref_s ) capacitor c=0.00348171f \
 //x=2.31 //y=1.22 //x2=2.965 //y2=0.375
cc_149 ( N_noxref_5_M0_noxref_s N_noxref_7_M2_noxref_d ) capacitor \
 c=0.00309936f //x=0.455 //y=0.375 //x2=3.395 //y2=0.915
cc_150 ( N_noxref_5_c_197_n N_noxref_8_c_347_n ) capacitor c=0.0136048f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_151 ( N_noxref_5_c_211_n N_noxref_8_c_347_n ) capacitor c=0.0102337f \
 //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_152 ( N_noxref_5_M0_noxref_s N_noxref_8_c_347_n ) capacitor c=0.023368f \
 //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_153 ( N_noxref_5_M0_noxref_s N_noxref_8_c_348_n ) capacitor c=0.0180035f \
 //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_154 ( N_noxref_5_c_197_n N_noxref_8_M1_noxref_d ) capacitor c=0.0129526f \
 //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_155 ( N_noxref_5_c_211_n N_noxref_8_M1_noxref_d ) capacitor c=0.0091401f \
 //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_156 ( N_noxref_5_M0_noxref_s N_noxref_8_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_157 ( N_noxref_5_M0_noxref_s N_noxref_8_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_158 ( N_noxref_6_M7_noxref_g N_noxref_7_c_285_n ) capacitor c=0.0209597f \
 //x=3.07 //y=6.02 //x2=3.205 //y2=5.155
cc_159 ( N_noxref_6_M8_noxref_g N_noxref_7_c_288_n ) capacitor c=0.0230978f \
 //x=3.51 //y=6.02 //x2=3.985 //y2=5.155
cc_160 ( N_noxref_6_c_245_n N_noxref_7_c_288_n ) capacitor c=0.00201851f \
 //x=3.33 //y=4.7 //x2=3.985 //y2=5.155
cc_161 ( N_noxref_6_c_251_p N_noxref_7_c_278_n ) capacitor c=0.00359704f \
 //x=3.695 //y=1.415 //x2=3.985 //y2=1.665
cc_162 ( N_noxref_6_c_252_p N_noxref_7_c_278_n ) capacitor c=0.00457401f \
 //x=3.85 //y=1.26 //x2=3.985 //y2=1.665
cc_163 ( N_noxref_6_c_226_n N_noxref_7_c_291_n ) capacitor c=0.0937541f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=5.07
cc_164 ( N_noxref_6_c_242_n N_noxref_7_c_291_n ) capacitor c=0.00877984f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=5.07
cc_165 ( N_noxref_6_c_244_n N_noxref_7_c_291_n ) capacitor c=0.00283672f \
 //x=3.33 //y=1.915 //x2=4.07 //y2=5.07
cc_166 ( N_noxref_6_c_245_n N_noxref_7_c_291_n ) capacitor c=0.013844f \
 //x=3.33 //y=4.7 //x2=4.07 //y2=5.07
cc_167 ( N_noxref_6_c_226_n N_noxref_7_c_329_n ) capacitor c=0.017915f \
 //x=3.33 //y=2.08 //x2=3.29 //y2=5.155
cc_168 ( N_noxref_6_c_245_n N_noxref_7_c_329_n ) capacitor c=0.00625229f \
 //x=3.33 //y=4.7 //x2=3.29 //y2=5.155
cc_169 ( N_noxref_6_c_239_n N_noxref_7_M2_noxref_d ) capacitor c=0.00217566f \
 //x=3.32 //y=0.915 //x2=3.395 //y2=0.915
cc_170 ( N_noxref_6_c_240_n N_noxref_7_M2_noxref_d ) capacitor c=0.0034598f \
 //x=3.32 //y=1.26 //x2=3.395 //y2=0.915
cc_171 ( N_noxref_6_c_241_n N_noxref_7_M2_noxref_d ) capacitor c=0.00544291f \
 //x=3.32 //y=1.57 //x2=3.395 //y2=0.915
cc_172 ( N_noxref_6_c_262_p N_noxref_7_M2_noxref_d ) capacitor c=0.00241102f \
 //x=3.695 //y=0.76 //x2=3.395 //y2=0.915
cc_173 ( N_noxref_6_c_251_p N_noxref_7_M2_noxref_d ) capacitor c=0.0140297f \
 //x=3.695 //y=1.415 //x2=3.395 //y2=0.915
cc_174 ( N_noxref_6_c_264_p N_noxref_7_M2_noxref_d ) capacitor c=0.00219619f \
 //x=3.85 //y=0.915 //x2=3.395 //y2=0.915
cc_175 ( N_noxref_6_c_252_p N_noxref_7_M2_noxref_d ) capacitor c=0.00603828f \
 //x=3.85 //y=1.26 //x2=3.395 //y2=0.915
cc_176 ( N_noxref_6_c_244_n N_noxref_7_M2_noxref_d ) capacitor c=0.00661782f \
 //x=3.33 //y=1.915 //x2=3.395 //y2=0.915
cc_177 ( N_noxref_6_M7_noxref_g N_noxref_7_M7_noxref_d ) capacitor \
 c=0.0180032f //x=3.07 //y=6.02 //x2=3.145 //y2=5.02
cc_178 ( N_noxref_6_M8_noxref_g N_noxref_7_M7_noxref_d ) capacitor \
 c=0.0194246f //x=3.51 //y=6.02 //x2=3.145 //y2=5.02
cc_179 ( N_noxref_6_c_226_n N_noxref_8_c_349_n ) capacitor c=0.00210069f \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_180 ( N_noxref_6_c_239_n N_noxref_8_c_349_n ) capacitor c=0.0192822f \
 //x=3.32 //y=0.915 //x2=3.985 //y2=0.54
cc_181 ( N_noxref_6_c_264_p N_noxref_8_c_349_n ) capacitor c=0.00656458f \
 //x=3.85 //y=0.915 //x2=3.985 //y2=0.54
cc_182 ( N_noxref_6_c_242_n N_noxref_8_c_349_n ) capacitor c=2.20712e-19 \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_183 ( N_noxref_6_c_240_n N_noxref_8_c_377_n ) capacitor c=0.00538829f \
 //x=3.32 //y=1.26 //x2=3.1 //y2=0.995
cc_184 ( N_noxref_6_c_239_n N_noxref_8_M2_noxref_s ) capacitor c=0.00538829f \
 //x=3.32 //y=0.915 //x2=2.965 //y2=0.375
cc_185 ( N_noxref_6_c_241_n N_noxref_8_M2_noxref_s ) capacitor c=0.00538829f \
 //x=3.32 //y=1.57 //x2=2.965 //y2=0.375
cc_186 ( N_noxref_6_c_264_p N_noxref_8_M2_noxref_s ) capacitor c=0.0143002f \
 //x=3.85 //y=0.915 //x2=2.965 //y2=0.375
cc_187 ( N_noxref_6_c_252_p N_noxref_8_M2_noxref_s ) capacitor c=0.00290153f \
 //x=3.85 //y=1.26 //x2=2.965 //y2=0.375
cc_188 ( N_noxref_7_c_278_n N_noxref_8_c_349_n ) capacitor c=0.0046926f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_189 ( N_noxref_7_M2_noxref_d N_noxref_8_c_349_n ) capacitor c=0.0118457f \
 //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_190 ( N_noxref_7_c_343_p N_noxref_8_c_377_n ) capacitor c=0.0200405f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_191 ( N_noxref_7_M2_noxref_d N_noxref_8_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_192 ( N_noxref_7_c_278_n N_noxref_8_M2_noxref_s ) capacitor c=0.0212001f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_193 ( N_noxref_7_M2_noxref_d N_noxref_8_M2_noxref_s ) capacitor \
 c=0.0426368f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
