* SPICE3 file created from DLATCH.ext - technology: sky130A

.subckt DLATCH Q D GATE VDD GND
M1000 a_3461_1051.t1 Q.t4 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VDD.t6 GATE.t0 a_661_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t9 a_1295_209.t3 a_2795_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t4 a_1771_1050.t5 a_2405_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_185_209.t1 D.t1 VDD.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_1295_209.t1 a_661_1050.t5 VDD.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VDD.t10 D.t2 a_1771_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_661_1050.t0 GATE.t1 VDD.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1771_1050.t0 D.t3 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 Q.t1 a_3007_411.t4 a_2795_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_3461_1051.t3 a_2405_209.t3 a_3007_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 GND GATE.t4 a_1666_101.t0 nshort w=-1.605u l=1.765u
+  ad=7.6538p pd=53.32u as=0p ps=0u
M1012 a_661_1050.t4 a_185_209.t4 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1771_1050.t4 GATE.t3 VDD.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_2795_1051.t0 a_1295_209.t4 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD.t3 Q.t6 a_3461_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_2405_209.t0 a_1771_1050.t6 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 Q a_1295_209.t5 GND.t2 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.15u as=0p ps=0u
M1018 Q a_3007_411.t5 GND.t8 nshort w=-1.83u l=2.06u
+  ad=0p pd=0u as=0p ps=0u
M1019 VDD.t5 a_185_209.t5 a_661_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VDD.t15 GATE.t5 a_1771_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t11 D.t4 a_185_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t16 a_661_1050.t7 a_1295_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_3007_411.t1 a_2405_209.t5 a_3461_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 GND a_185_209.t3 a_556_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2795_1051.t3 a_3007_411.t6 Q.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 GATE D 0.58fF
C1 VDD D 0.19fF
C2 GATE VDD 0.15fF
C3 Q VDD 0.33fF
R0 Q.n0 Q.t4 486.819
R1 Q.n0 Q.t6 384.527
R2 Q.n1 Q.t5 250.501
R3 Q.n11 Q.n2 191.889
R4 Q.n11 Q.n10 135.634
R5 Q.n1 Q.n0 133.1
R6 Q.n10 Q.n9 118.016
R7 Q.n5 Q.n3 80.526
R8 Q.n12 Q.n1 77.315
R9 Q.n12 Q.n11 76
R10 Q.n10 Q.n5 48.405
R11 Q.n9 Q.n8 30
R12 Q.n5 Q.n4 30
R13 Q.n7 Q.n6 24.383
R14 Q.n9 Q.n7 23.684
R15 Q.n2 Q.t2 14.282
R16 Q.n2 Q.t1 14.282
R17 Q.n12 Q 0.046
R18 VDD.n242 VDD.n240 144.705
R19 VDD.n304 VDD.n302 144.705
R20 VDD.n184 VDD.n182 144.705
R21 VDD.n371 VDD.n369 144.705
R22 VDD.n138 VDD.n136 144.705
R23 VDD.n80 VDD.n78 144.705
R24 VDD.n143 VDD.n142 77.792
R25 VDD.n152 VDD.n151 77.792
R26 VDD.n340 VDD.n339 77.792
R27 VDD.n330 VDD.n329 77.792
R28 VDD.n232 VDD.n231 77.792
R29 VDD.n221 VDD.n220 77.792
R30 VDD.n40 VDD.n39 76
R31 VDD.n47 VDD.n46 76
R32 VDD.n51 VDD.n50 76
R33 VDD.n55 VDD.n54 76
R34 VDD.n82 VDD.n81 76
R35 VDD.n86 VDD.n85 76
R36 VDD.n90 VDD.n89 76
R37 VDD.n94 VDD.n93 76
R38 VDD.n99 VDD.n98 76
R39 VDD.n106 VDD.n105 76
R40 VDD.n110 VDD.n109 76
R41 VDD.n114 VDD.n113 76
R42 VDD.n140 VDD.n139 76
R43 VDD.n146 VDD.n145 76
R44 VDD.n150 VDD.n149 76
R45 VDD.n156 VDD.n155 76
R46 VDD.n160 VDD.n159 76
R47 VDD.n186 VDD.n185 76
R48 VDD.n191 VDD.n190 76
R49 VDD.n196 VDD.n195 76
R50 VDD.n394 VDD.n393 76
R51 VDD.n388 VDD.n387 76
R52 VDD.n383 VDD.n382 76
R53 VDD.n378 VDD.n377 76
R54 VDD.n373 VDD.n372 76
R55 VDD.n347 VDD.n346 76
R56 VDD.n343 VDD.n342 76
R57 VDD.n337 VDD.n336 76
R58 VDD.n333 VDD.n332 76
R59 VDD.n327 VDD.n326 76
R60 VDD.n301 VDD.n300 76
R61 VDD.n297 VDD.n296 76
R62 VDD.n292 VDD.n291 76
R63 VDD.n287 VDD.n286 76
R64 VDD.n281 VDD.n280 76
R65 VDD.n276 VDD.n275 76
R66 VDD.n271 VDD.n270 76
R67 VDD.n266 VDD.n265 76
R68 VDD.n239 VDD.n238 76
R69 VDD.n235 VDD.n234 76
R70 VDD.n229 VDD.n228 76
R71 VDD.n225 VDD.n224 76
R72 VDD.n219 VDD.n218 76
R73 VDD.n223 VDD.t7 55.106
R74 VDD.n230 VDD.t11 55.106
R75 VDD.n267 VDD.t0 55.106
R76 VDD.n328 VDD.t13 55.106
R77 VDD.n338 VDD.t16 55.106
R78 VDD.n374 VDD.t14 55.106
R79 VDD.n154 VDD.t8 55.106
R80 VDD.n141 VDD.t4 55.106
R81 VDD.n295 VDD.t6 55.106
R82 VDD.n187 VDD.t10 55.106
R83 VDD.n101 VDD.n100 41.183
R84 VDD.n42 VDD.n41 41.183
R85 VDD.n285 VDD.n284 40.824
R86 VDD.n390 VDD.n389 40.824
R87 VDD.n309 VDD.n308 36.774
R88 VDD.n352 VDD.n351 36.774
R89 VDD.n165 VDD.n164 36.774
R90 VDD.n119 VDD.n118 36.774
R91 VDD.n60 VDD.n59 36.774
R92 VDD.n258 VDD.n257 36.774
R93 VDD.n193 VDD.n192 36.608
R94 VDD.n289 VDD.n288 36.608
R95 VDD.n34 VDD.n33 34.942
R96 VDD.n44 VDD.n43 32.032
R97 VDD.n103 VDD.n102 32.032
R98 VDD.n380 VDD.n379 32.032
R99 VDD.n273 VDD.n272 32.032
R100 VDD.n218 VDD.n215 21.841
R101 VDD.n23 VDD.n20 21.841
R102 VDD.n284 VDD.t17 14.282
R103 VDD.n284 VDD.t5 14.282
R104 VDD.n389 VDD.t12 14.282
R105 VDD.n389 VDD.t15 14.282
R106 VDD.n100 VDD.t1 14.282
R107 VDD.n100 VDD.t9 14.282
R108 VDD.n41 VDD.t2 14.282
R109 VDD.n41 VDD.t3 14.282
R110 VDD.n215 VDD.n198 14.167
R111 VDD.n198 VDD.n197 14.167
R112 VDD.n324 VDD.n306 14.167
R113 VDD.n306 VDD.n305 14.167
R114 VDD.n367 VDD.n349 14.167
R115 VDD.n349 VDD.n348 14.167
R116 VDD.n180 VDD.n162 14.167
R117 VDD.n162 VDD.n161 14.167
R118 VDD.n134 VDD.n116 14.167
R119 VDD.n116 VDD.n115 14.167
R120 VDD.n76 VDD.n57 14.167
R121 VDD.n57 VDD.n56 14.167
R122 VDD.n263 VDD.n244 14.167
R123 VDD.n244 VDD.n243 14.167
R124 VDD.n20 VDD.n19 14.167
R125 VDD.n19 VDD.n17 14.167
R126 VDD.n32 VDD.n31 14.167
R127 VDD.n31 VDD.n28 14.167
R128 VDD.n81 VDD.n77 14.167
R129 VDD.n139 VDD.n135 14.167
R130 VDD.n185 VDD.n181 14.167
R131 VDD.n372 VDD.n368 14.167
R132 VDD.n326 VDD.n325 14.167
R133 VDD.n265 VDD.n264 14.167
R134 VDD.n23 VDD.n22 13.653
R135 VDD.n22 VDD.n21 13.653
R136 VDD.n32 VDD.n25 13.653
R137 VDD.n25 VDD.n24 13.653
R138 VDD.n31 VDD.n30 13.653
R139 VDD.n30 VDD.n29 13.653
R140 VDD.n28 VDD.n27 13.653
R141 VDD.n27 VDD.n26 13.653
R142 VDD.n39 VDD.n38 13.653
R143 VDD.n38 VDD.n37 13.653
R144 VDD.n46 VDD.n45 13.653
R145 VDD.n45 VDD.n44 13.653
R146 VDD.n50 VDD.n49 13.653
R147 VDD.n49 VDD.n48 13.653
R148 VDD.n54 VDD.n53 13.653
R149 VDD.n53 VDD.n52 13.653
R150 VDD.n81 VDD.n80 13.653
R151 VDD.n80 VDD.n79 13.653
R152 VDD.n85 VDD.n84 13.653
R153 VDD.n84 VDD.n83 13.653
R154 VDD.n89 VDD.n88 13.653
R155 VDD.n88 VDD.n87 13.653
R156 VDD.n93 VDD.n92 13.653
R157 VDD.n92 VDD.n91 13.653
R158 VDD.n98 VDD.n97 13.653
R159 VDD.n97 VDD.n96 13.653
R160 VDD.n105 VDD.n104 13.653
R161 VDD.n104 VDD.n103 13.653
R162 VDD.n109 VDD.n108 13.653
R163 VDD.n108 VDD.n107 13.653
R164 VDD.n113 VDD.n112 13.653
R165 VDD.n112 VDD.n111 13.653
R166 VDD.n139 VDD.n138 13.653
R167 VDD.n138 VDD.n137 13.653
R168 VDD.n145 VDD.n144 13.653
R169 VDD.n144 VDD.n143 13.653
R170 VDD.n149 VDD.n148 13.653
R171 VDD.n148 VDD.n147 13.653
R172 VDD.n155 VDD.n153 13.653
R173 VDD.n153 VDD.n152 13.653
R174 VDD.n159 VDD.n158 13.653
R175 VDD.n158 VDD.n157 13.653
R176 VDD.n185 VDD.n184 13.653
R177 VDD.n184 VDD.n183 13.653
R178 VDD.n190 VDD.n189 13.653
R179 VDD.n189 VDD.n188 13.653
R180 VDD.n195 VDD.n194 13.653
R181 VDD.n194 VDD.n193 13.653
R182 VDD.n393 VDD.n392 13.653
R183 VDD.n392 VDD.n391 13.653
R184 VDD.n387 VDD.n386 13.653
R185 VDD.n386 VDD.n385 13.653
R186 VDD.n382 VDD.n381 13.653
R187 VDD.n381 VDD.n380 13.653
R188 VDD.n377 VDD.n376 13.653
R189 VDD.n376 VDD.n375 13.653
R190 VDD.n372 VDD.n371 13.653
R191 VDD.n371 VDD.n370 13.653
R192 VDD.n346 VDD.n345 13.653
R193 VDD.n345 VDD.n344 13.653
R194 VDD.n342 VDD.n341 13.653
R195 VDD.n341 VDD.n340 13.653
R196 VDD.n336 VDD.n335 13.653
R197 VDD.n335 VDD.n334 13.653
R198 VDD.n332 VDD.n331 13.653
R199 VDD.n331 VDD.n330 13.653
R200 VDD.n326 VDD.n304 13.653
R201 VDD.n304 VDD.n303 13.653
R202 VDD.n300 VDD.n299 13.653
R203 VDD.n299 VDD.n298 13.653
R204 VDD.n296 VDD.n294 13.653
R205 VDD.n294 VDD.n293 13.653
R206 VDD.n291 VDD.n290 13.653
R207 VDD.n290 VDD.n289 13.653
R208 VDD.n286 VDD.n283 13.653
R209 VDD.n283 VDD.n282 13.653
R210 VDD.n280 VDD.n279 13.653
R211 VDD.n279 VDD.n278 13.653
R212 VDD.n275 VDD.n274 13.653
R213 VDD.n274 VDD.n273 13.653
R214 VDD.n270 VDD.n269 13.653
R215 VDD.n269 VDD.n268 13.653
R216 VDD.n265 VDD.n242 13.653
R217 VDD.n242 VDD.n241 13.653
R218 VDD.n238 VDD.n237 13.653
R219 VDD.n237 VDD.n236 13.653
R220 VDD.n234 VDD.n233 13.653
R221 VDD.n233 VDD.n232 13.653
R222 VDD.n228 VDD.n227 13.653
R223 VDD.n227 VDD.n226 13.653
R224 VDD.n224 VDD.n222 13.653
R225 VDD.n222 VDD.n221 13.653
R226 VDD.n218 VDD.n217 13.653
R227 VDD.n217 VDD.n216 13.653
R228 VDD.n4 VDD.n2 12.915
R229 VDD.n4 VDD.n3 12.66
R230 VDD.n13 VDD.n12 12.343
R231 VDD.n10 VDD.n9 12.343
R232 VDD.n10 VDD.n7 12.343
R233 VDD.n393 VDD.n390 8.658
R234 VDD.n286 VDD.n285 8.658
R235 VDD.n325 VDD.n324 7.674
R236 VDD.n368 VDD.n367 7.674
R237 VDD.n181 VDD.n180 7.674
R238 VDD.n135 VDD.n134 7.674
R239 VDD.n77 VDD.n76 7.674
R240 VDD.n264 VDD.n263 7.674
R241 VDD.n71 VDD.n70 7.5
R242 VDD.n65 VDD.n64 7.5
R243 VDD.n67 VDD.n66 7.5
R244 VDD.n62 VDD.n61 7.5
R245 VDD.n76 VDD.n75 7.5
R246 VDD.n129 VDD.n128 7.5
R247 VDD.n123 VDD.n122 7.5
R248 VDD.n125 VDD.n124 7.5
R249 VDD.n131 VDD.n121 7.5
R250 VDD.n131 VDD.n119 7.5
R251 VDD.n134 VDD.n133 7.5
R252 VDD.n175 VDD.n174 7.5
R253 VDD.n169 VDD.n168 7.5
R254 VDD.n171 VDD.n170 7.5
R255 VDD.n177 VDD.n167 7.5
R256 VDD.n177 VDD.n165 7.5
R257 VDD.n180 VDD.n179 7.5
R258 VDD.n362 VDD.n361 7.5
R259 VDD.n356 VDD.n355 7.5
R260 VDD.n358 VDD.n357 7.5
R261 VDD.n364 VDD.n354 7.5
R262 VDD.n364 VDD.n352 7.5
R263 VDD.n367 VDD.n366 7.5
R264 VDD.n319 VDD.n318 7.5
R265 VDD.n313 VDD.n312 7.5
R266 VDD.n315 VDD.n314 7.5
R267 VDD.n321 VDD.n311 7.5
R268 VDD.n321 VDD.n309 7.5
R269 VDD.n324 VDD.n323 7.5
R270 VDD.n248 VDD.n247 7.5
R271 VDD.n251 VDD.n250 7.5
R272 VDD.n253 VDD.n252 7.5
R273 VDD.n256 VDD.n255 7.5
R274 VDD.n263 VDD.n262 7.5
R275 VDD.n210 VDD.n209 7.5
R276 VDD.n204 VDD.n203 7.5
R277 VDD.n206 VDD.n205 7.5
R278 VDD.n212 VDD.n202 7.5
R279 VDD.n212 VDD.n200 7.5
R280 VDD.n215 VDD.n214 7.5
R281 VDD.n20 VDD.n16 7.5
R282 VDD.n2 VDD.n1 7.5
R283 VDD.n9 VDD.n8 7.5
R284 VDD.n7 VDD.n6 7.5
R285 VDD.n19 VDD.n18 7.5
R286 VDD.n14 VDD.n0 7.5
R287 VDD.n63 VDD.n60 6.772
R288 VDD.n74 VDD.n58 6.772
R289 VDD.n72 VDD.n69 6.772
R290 VDD.n68 VDD.n65 6.772
R291 VDD.n132 VDD.n117 6.772
R292 VDD.n130 VDD.n127 6.772
R293 VDD.n126 VDD.n123 6.772
R294 VDD.n178 VDD.n163 6.772
R295 VDD.n176 VDD.n173 6.772
R296 VDD.n172 VDD.n169 6.772
R297 VDD.n365 VDD.n350 6.772
R298 VDD.n363 VDD.n360 6.772
R299 VDD.n359 VDD.n356 6.772
R300 VDD.n322 VDD.n307 6.772
R301 VDD.n320 VDD.n317 6.772
R302 VDD.n316 VDD.n313 6.772
R303 VDD.n213 VDD.n199 6.772
R304 VDD.n211 VDD.n208 6.772
R305 VDD.n207 VDD.n204 6.772
R306 VDD.n63 VDD.n62 6.772
R307 VDD.n68 VDD.n67 6.772
R308 VDD.n72 VDD.n71 6.772
R309 VDD.n75 VDD.n74 6.772
R310 VDD.n126 VDD.n125 6.772
R311 VDD.n130 VDD.n129 6.772
R312 VDD.n133 VDD.n132 6.772
R313 VDD.n172 VDD.n171 6.772
R314 VDD.n176 VDD.n175 6.772
R315 VDD.n179 VDD.n178 6.772
R316 VDD.n359 VDD.n358 6.772
R317 VDD.n363 VDD.n362 6.772
R318 VDD.n366 VDD.n365 6.772
R319 VDD.n316 VDD.n315 6.772
R320 VDD.n320 VDD.n319 6.772
R321 VDD.n323 VDD.n322 6.772
R322 VDD.n207 VDD.n206 6.772
R323 VDD.n211 VDD.n210 6.772
R324 VDD.n214 VDD.n213 6.772
R325 VDD.n262 VDD.n261 6.772
R326 VDD.n249 VDD.n246 6.772
R327 VDD.n254 VDD.n251 6.772
R328 VDD.n259 VDD.n256 6.772
R329 VDD.n259 VDD.n258 6.772
R330 VDD.n254 VDD.n253 6.772
R331 VDD.n249 VDD.n248 6.772
R332 VDD.n261 VDD.n245 6.772
R333 VDD.n33 VDD.n23 6.487
R334 VDD.n33 VDD.n32 6.475
R335 VDD.n16 VDD.n15 6.458
R336 VDD.n121 VDD.n120 6.202
R337 VDD.n167 VDD.n166 6.202
R338 VDD.n354 VDD.n353 6.202
R339 VDD.n311 VDD.n310 6.202
R340 VDD.n202 VDD.n201 6.202
R341 VDD.n46 VDD.n42 5.903
R342 VDD.n105 VDD.n101 5.903
R343 VDD.n37 VDD.n36 4.576
R344 VDD.n96 VDD.n95 4.576
R345 VDD.n385 VDD.n384 4.576
R346 VDD.n278 VDD.n277 4.576
R347 VDD.n377 VDD.n374 2.754
R348 VDD.n270 VDD.n267 2.754
R349 VDD.n190 VDD.n187 2.361
R350 VDD.n296 VDD.n295 2.361
R351 VDD.n145 VDD.n141 1.967
R352 VDD.n155 VDD.n154 1.967
R353 VDD.n342 VDD.n338 1.967
R354 VDD.n332 VDD.n328 1.967
R355 VDD.n234 VDD.n230 1.967
R356 VDD.n224 VDD.n223 1.967
R357 VDD.n14 VDD.n5 1.329
R358 VDD.n14 VDD.n10 1.329
R359 VDD.n14 VDD.n11 1.329
R360 VDD.n14 VDD.n13 1.329
R361 VDD.n15 VDD.n14 0.696
R362 VDD.n14 VDD.n4 0.696
R363 VDD.n73 VDD.n72 0.365
R364 VDD.n73 VDD.n68 0.365
R365 VDD.n73 VDD.n63 0.365
R366 VDD.n74 VDD.n73 0.365
R367 VDD.n131 VDD.n130 0.365
R368 VDD.n131 VDD.n126 0.365
R369 VDD.n132 VDD.n131 0.365
R370 VDD.n177 VDD.n176 0.365
R371 VDD.n177 VDD.n172 0.365
R372 VDD.n178 VDD.n177 0.365
R373 VDD.n364 VDD.n363 0.365
R374 VDD.n364 VDD.n359 0.365
R375 VDD.n365 VDD.n364 0.365
R376 VDD.n321 VDD.n320 0.365
R377 VDD.n321 VDD.n316 0.365
R378 VDD.n322 VDD.n321 0.365
R379 VDD.n212 VDD.n211 0.365
R380 VDD.n212 VDD.n207 0.365
R381 VDD.n213 VDD.n212 0.365
R382 VDD.n260 VDD.n259 0.365
R383 VDD.n260 VDD.n254 0.365
R384 VDD.n260 VDD.n249 0.365
R385 VDD.n261 VDD.n260 0.365
R386 VDD.n82 VDD.n55 0.29
R387 VDD.n140 VDD.n114 0.29
R388 VDD.n186 VDD.n160 0.29
R389 VDD.n373 VDD.n347 0.29
R390 VDD.n327 VDD.n301 0.29
R391 VDD.n266 VDD.n239 0.29
R392 VDD.n219 VDD 0.207
R393 VDD.n40 VDD.n35 0.181
R394 VDD.n99 VDD.n94 0.181
R395 VDD.n394 VDD.n388 0.181
R396 VDD.n287 VDD.n281 0.181
R397 VDD.n150 VDD.n146 0.157
R398 VDD.n156 VDD.n150 0.157
R399 VDD.n343 VDD.n337 0.157
R400 VDD.n337 VDD.n333 0.157
R401 VDD.n235 VDD.n229 0.157
R402 VDD.n229 VDD.n225 0.157
R403 VDD.n35 VDD.n34 0.145
R404 VDD.n47 VDD.n40 0.145
R405 VDD.n51 VDD.n47 0.145
R406 VDD.n55 VDD.n51 0.145
R407 VDD.n86 VDD.n82 0.145
R408 VDD.n90 VDD.n86 0.145
R409 VDD.n94 VDD.n90 0.145
R410 VDD.n106 VDD.n99 0.145
R411 VDD.n110 VDD.n106 0.145
R412 VDD.n114 VDD.n110 0.145
R413 VDD.n146 VDD.n140 0.145
R414 VDD.n160 VDD.n156 0.145
R415 VDD.n191 VDD.n186 0.145
R416 VDD.n196 VDD.n191 0.145
R417 VDD.n388 VDD.n383 0.145
R418 VDD.n383 VDD.n378 0.145
R419 VDD.n378 VDD.n373 0.145
R420 VDD.n347 VDD.n343 0.145
R421 VDD.n333 VDD.n327 0.145
R422 VDD.n301 VDD.n297 0.145
R423 VDD.n297 VDD.n292 0.145
R424 VDD.n292 VDD.n287 0.145
R425 VDD.n281 VDD.n276 0.145
R426 VDD.n276 VDD.n271 0.145
R427 VDD.n271 VDD.n266 0.145
R428 VDD.n239 VDD.n235 0.145
R429 VDD.n225 VDD.n219 0.145
R430 VDD VDD.n394 0.133
R431 VDD VDD.n196 0.012
R432 a_3461_1051.n0 a_3461_1051.t3 101.66
R433 a_3461_1051.n0 a_3461_1051.t0 101.66
R434 a_3461_1051.n0 a_3461_1051.t2 14.294
R435 a_3461_1051.t1 a_3461_1051.n0 14.282
R436 D.n2 D.t4 512.525
R437 D.n0 D.t2 472.359
R438 D.n0 D.t3 384.527
R439 D.n2 D.t1 371.139
R440 D.n1 D.t5 267.725
R441 D.n3 D.t0 263.54
R442 D.n3 D.n2 120.094
R443 D.n1 D.n0 83.507
R444 D.n4 D.n1 82.484
R445 D.n4 D.n3 76
R446 D.n4 D 0.046
R447 GND.n43 GND.n41 219.745
R448 GND.n165 GND.n164 219.745
R449 GND.n195 GND.n193 219.745
R450 GND.n228 GND.n226 219.745
R451 GND.n120 GND.n118 219.745
R452 GND.n87 GND.n86 219.745
R453 GND.n43 GND.n42 85.529
R454 GND.n165 GND.n163 85.529
R455 GND.n195 GND.n194 85.529
R456 GND.n228 GND.n227 85.529
R457 GND.n120 GND.n119 85.529
R458 GND.n87 GND.n85 85.529
R459 GND.n236 GND.n235 84.842
R460 GND.n173 GND.n172 84.842
R461 GND.n8 GND.n1 76.145
R462 GND.n133 GND.n132 76
R463 GND.n8 GND.n7 76
R464 GND.n14 GND.n13 76
R465 GND.n17 GND.n16 76
R466 GND.n24 GND.n23 76
R467 GND.n30 GND.n29 76
R468 GND.n37 GND.n36 76
R469 GND.n40 GND.n39 76
R470 GND.n47 GND.n46 76
R471 GND.n54 GND.n53 76
R472 GND.n60 GND.n59 76
R473 GND.n63 GND.n62 76
R474 GND.n69 GND.n68 76
R475 GND.n74 GND.n73 76
R476 GND.n81 GND.n80 76
R477 GND.n84 GND.n83 76
R478 GND.n91 GND.n90 76
R479 GND.n99 GND.n98 76
R480 GND.n107 GND.n106 76
R481 GND.n114 GND.n113 76
R482 GND.n117 GND.n116 76
R483 GND.n124 GND.n123 76
R484 GND.n127 GND.n126 76
R485 GND.n130 GND.n129 76
R486 GND.n245 GND.n244 76
R487 GND.n242 GND.n241 76
R488 GND.n239 GND.n238 76
R489 GND.n234 GND.n233 76
R490 GND.n231 GND.n230 76
R491 GND.n224 GND.n223 76
R492 GND.n221 GND.n220 76
R493 GND.n213 GND.n212 76
R494 GND.n205 GND.n204 76
R495 GND.n198 GND.n197 76
R496 GND.n191 GND.n190 76
R497 GND.n188 GND.n187 76
R498 GND.n185 GND.n184 76
R499 GND.n182 GND.n181 76
R500 GND.n179 GND.n178 76
R501 GND.n176 GND.n175 76
R502 GND.n171 GND.n170 76
R503 GND.n168 GND.n167 76
R504 GND.n161 GND.n160 76
R505 GND.n158 GND.n157 76
R506 GND.n150 GND.n149 76
R507 GND.n142 GND.n141 76
R508 GND.n33 GND.t1 39.412
R509 GND.n138 GND.t0 39.412
R510 GND.n95 GND.n94 35.01
R511 GND.n217 GND.n216 35.01
R512 GND.n154 GND.n153 35.01
R513 GND.n93 GND.n92 29.127
R514 GND.n215 GND.n214 29.127
R515 GND.n102 GND.t6 20.794
R516 GND.n208 GND.t3 20.794
R517 GND.n27 GND.n26 19.735
R518 GND.n21 GND.n20 19.735
R519 GND.n12 GND.n11 19.735
R520 GND.n5 GND.n4 19.735
R521 GND.n35 GND.n34 19.735
R522 GND.n71 GND.n70 19.735
R523 GND.n66 GND.n65 19.735
R524 GND.n58 GND.n57 19.735
R525 GND.n51 GND.n50 19.735
R526 GND.n79 GND.n78 19.735
R527 GND.n96 GND.n95 19.735
R528 GND.n104 GND.n103 19.735
R529 GND.n112 GND.n111 19.735
R530 GND.n218 GND.n217 19.735
R531 GND.n210 GND.n209 19.735
R532 GND.n203 GND.n202 19.735
R533 GND.n155 GND.n154 19.735
R534 GND.n147 GND.n146 19.735
R535 GND.n140 GND.n139 19.735
R536 GND.n11 GND.t7 19.724
R537 GND.n57 GND.t8 19.724
R538 GND.n70 GND.t2 19.724
R539 GND.n95 GND.n93 19.017
R540 GND.n217 GND.n215 19.017
R541 GND.n154 GND.n152 19.017
R542 GND.n33 GND.n32 17.185
R543 GND.n138 GND.n137 17.185
R544 GND.n46 GND.n44 14.167
R545 GND.n90 GND.n88 14.167
R546 GND.n123 GND.n121 14.167
R547 GND.n230 GND.n229 14.167
R548 GND.n197 GND.n196 14.167
R549 GND.n167 GND.n166 14.167
R550 GND.n19 GND.n18 13.654
R551 GND.n141 GND.n134 13.653
R552 GND.n149 GND.n148 13.653
R553 GND.n157 GND.n156 13.653
R554 GND.n160 GND.n159 13.653
R555 GND.n167 GND.n162 13.653
R556 GND.n170 GND.n169 13.653
R557 GND.n175 GND.n174 13.653
R558 GND.n178 GND.n177 13.653
R559 GND.n181 GND.n180 13.653
R560 GND.n184 GND.n183 13.653
R561 GND.n187 GND.n186 13.653
R562 GND.n190 GND.n189 13.653
R563 GND.n197 GND.n192 13.653
R564 GND.n204 GND.n199 13.653
R565 GND.n212 GND.n211 13.653
R566 GND.n220 GND.n219 13.653
R567 GND.n223 GND.n222 13.653
R568 GND.n230 GND.n225 13.653
R569 GND.n233 GND.n232 13.653
R570 GND.n238 GND.n237 13.653
R571 GND.n241 GND.n240 13.653
R572 GND.n244 GND.n243 13.653
R573 GND.n129 GND.n128 13.653
R574 GND.n126 GND.n125 13.653
R575 GND.n123 GND.n122 13.653
R576 GND.n116 GND.n115 13.653
R577 GND.n113 GND.n108 13.653
R578 GND.n106 GND.n105 13.653
R579 GND.n98 GND.n97 13.653
R580 GND.n90 GND.n89 13.653
R581 GND.n83 GND.n82 13.653
R582 GND.n80 GND.n75 13.653
R583 GND.n73 GND.n72 13.653
R584 GND.n68 GND.n67 13.653
R585 GND.n62 GND.n61 13.653
R586 GND.n59 GND.n55 13.653
R587 GND.n53 GND.n52 13.653
R588 GND.n46 GND.n45 13.653
R589 GND.n39 GND.n38 13.653
R590 GND.n36 GND.n31 13.653
R591 GND.n29 GND.n28 13.653
R592 GND.n23 GND.n22 13.653
R593 GND.n16 GND.n15 13.653
R594 GND.n13 GND.n9 13.653
R595 GND.n7 GND.n6 13.653
R596 GND.n78 GND.n77 12.837
R597 GND.n111 GND.n110 12.837
R598 GND.n202 GND.n201 12.837
R599 GND.n4 GND.n3 11.605
R600 GND.n50 GND.n49 11.605
R601 GND.n3 GND.n2 9.809
R602 GND.n49 GND.n48 9.809
R603 GND.n23 GND.n21 8.854
R604 GND.n68 GND.n66 8.854
R605 GND.n77 GND.n76 7.566
R606 GND.n110 GND.n109 7.566
R607 GND.n201 GND.n200 7.566
R608 GND.n26 GND.n25 7.5
R609 GND.n152 GND.n151 7.5
R610 GND.n145 GND.n144 7.5
R611 GND.n44 GND.n43 7.312
R612 GND.n166 GND.n165 7.312
R613 GND.n196 GND.n195 7.312
R614 GND.n229 GND.n228 7.312
R615 GND.n121 GND.n120 7.312
R616 GND.n88 GND.n87 7.312
R617 GND.t7 GND.n10 7.04
R618 GND.t8 GND.n56 7.04
R619 GND.n34 GND.n33 6.139
R620 GND.n139 GND.n138 6.139
R621 GND.n20 GND.n19 5.774
R622 GND.n65 GND.n64 5.774
R623 GND.n101 GND.n100 4.551
R624 GND.n207 GND.n206 4.551
R625 GND.n136 GND.n135 4.551
R626 GND.n13 GND.n12 3.935
R627 GND.n29 GND.n27 3.935
R628 GND.n59 GND.n58 3.935
R629 GND.n73 GND.n71 3.935
R630 GND.n98 GND.n96 3.935
R631 GND.n238 GND.n236 3.935
R632 GND.n220 GND.n218 3.935
R633 GND.n175 GND.n173 3.935
R634 GND.n157 GND.n155 3.935
R635 GND.n113 GND.n112 3.541
R636 GND.n204 GND.n203 3.541
R637 GND.n141 GND.n140 3.541
R638 GND.t6 GND.n101 2.238
R639 GND.t3 GND.n207 2.238
R640 GND.t0 GND.n136 2.238
R641 GND.n144 GND.n143 1.935
R642 GND.n7 GND.n5 0.983
R643 GND.n36 GND.n35 0.983
R644 GND.n53 GND.n51 0.983
R645 GND.n80 GND.n79 0.983
R646 GND.n1 GND.n0 0.596
R647 GND.n132 GND.n131 0.596
R648 GND.n103 GND.n102 0.358
R649 GND.n209 GND.n208 0.358
R650 GND.n146 GND.n145 0.358
R651 GND.n47 GND.n40 0.29
R652 GND.n91 GND.n84 0.29
R653 GND.n124 GND.n117 0.29
R654 GND.n231 GND.n224 0.29
R655 GND.n198 GND.n191 0.29
R656 GND.n168 GND.n161 0.29
R657 GND.n133 GND 0.207
R658 GND.n106 GND.n104 0.196
R659 GND.n212 GND.n210 0.196
R660 GND.n149 GND.n147 0.196
R661 GND.n24 GND.n17 0.181
R662 GND.n69 GND.n63 0.181
R663 GND.n245 GND.n242 0.181
R664 GND.n182 GND.n179 0.181
R665 GND.n107 GND.n99 0.157
R666 GND.n114 GND.n107 0.157
R667 GND.n221 GND.n213 0.157
R668 GND.n213 GND.n205 0.157
R669 GND.n158 GND.n150 0.157
R670 GND.n150 GND.n142 0.157
R671 GND.n14 GND.n8 0.145
R672 GND.n17 GND.n14 0.145
R673 GND.n30 GND.n24 0.145
R674 GND.n37 GND.n30 0.145
R675 GND.n40 GND.n37 0.145
R676 GND.n54 GND.n47 0.145
R677 GND.n60 GND.n54 0.145
R678 GND.n63 GND.n60 0.145
R679 GND.n74 GND.n69 0.145
R680 GND.n81 GND.n74 0.145
R681 GND.n84 GND.n81 0.145
R682 GND.n99 GND.n91 0.145
R683 GND.n117 GND.n114 0.145
R684 GND.n127 GND.n124 0.145
R685 GND.n130 GND.n127 0.145
R686 GND.n242 GND.n239 0.145
R687 GND.n239 GND.n234 0.145
R688 GND.n234 GND.n231 0.145
R689 GND.n224 GND.n221 0.145
R690 GND.n205 GND.n198 0.145
R691 GND.n191 GND.n188 0.145
R692 GND.n188 GND.n185 0.145
R693 GND.n185 GND.n182 0.145
R694 GND.n179 GND.n176 0.145
R695 GND.n176 GND.n171 0.145
R696 GND.n171 GND.n168 0.145
R697 GND.n161 GND.n158 0.145
R698 GND.n142 GND.n133 0.145
R699 GND GND.n245 0.133
R700 GND GND.n130 0.012
R701 a_185_209.n0 a_185_209.t5 480.392
R702 a_185_209.n0 a_185_209.t4 403.272
R703 a_185_209.n1 a_185_209.t3 283.48
R704 a_185_209.n3 a_185_209.n2 227.307
R705 a_185_209.n4 a_185_209.n3 157.453
R706 a_185_209.n3 a_185_209.n1 153.315
R707 a_185_209.n1 a_185_209.n0 98.447
R708 a_185_209.n4 a_185_209.t0 14.282
R709 a_185_209.t1 a_185_209.n4 14.282
R710 a_556_101.t0 a_556_101.n1 34.62
R711 a_556_101.t0 a_556_101.n0 8.137
R712 a_556_101.t0 a_556_101.n2 4.69
R713 GATE.n0 GATE.t5 480.392
R714 GATE.n2 GATE.t0 472.359
R715 GATE.n0 GATE.t3 403.272
R716 GATE.n2 GATE.t1 384.527
R717 GATE.n1 GATE.t4 230.374
R718 GATE.n3 GATE.t2 188.066
R719 GATE.n3 GATE.n2 163.166
R720 GATE.n1 GATE.n0 151.553
R721 GATE.n4 GATE.n1 79.491
R722 GATE.n4 GATE.n3 76
R723 GATE.n4 GATE 0.046
R724 a_661_1050.n0 a_661_1050.t7 512.525
R725 a_661_1050.n0 a_661_1050.t5 371.139
R726 a_661_1050.n1 a_661_1050.t6 210.434
R727 a_661_1050.n3 a_661_1050.n2 205.778
R728 a_661_1050.n5 a_661_1050.n3 179.052
R729 a_661_1050.n1 a_661_1050.n0 173.2
R730 a_661_1050.n3 a_661_1050.n1 153.043
R731 a_661_1050.n5 a_661_1050.n4 76.002
R732 a_661_1050.n4 a_661_1050.t3 14.282
R733 a_661_1050.n4 a_661_1050.t4 14.282
R734 a_661_1050.t1 a_661_1050.n6 14.282
R735 a_661_1050.n6 a_661_1050.t0 14.282
R736 a_661_1050.n6 a_661_1050.n5 12.848
R737 a_1295_209.n0 a_1295_209.t4 486.819
R738 a_1295_209.n0 a_1295_209.t3 384.527
R739 a_1295_209.n1 a_1295_209.t5 277.054
R740 a_1295_209.n3 a_1295_209.n2 227.307
R741 a_1295_209.n4 a_1295_209.n3 157.453
R742 a_1295_209.n3 a_1295_209.n1 157.396
R743 a_1295_209.n1 a_1295_209.n0 106.547
R744 a_1295_209.n4 a_1295_209.t0 14.282
R745 a_1295_209.t1 a_1295_209.n4 14.282
R746 a_2795_1051.t1 a_2795_1051.n0 101.66
R747 a_2795_1051.n0 a_2795_1051.t3 101.659
R748 a_2795_1051.n0 a_2795_1051.t2 14.294
R749 a_2795_1051.n0 a_2795_1051.t0 14.282
R750 a_1771_1050.n0 a_1771_1050.t5 512.525
R751 a_1771_1050.n0 a_1771_1050.t6 371.139
R752 a_1771_1050.n1 a_1771_1050.t7 210.434
R753 a_1771_1050.n6 a_1771_1050.n5 184.039
R754 a_1771_1050.n8 a_1771_1050.n6 179.052
R755 a_1771_1050.n1 a_1771_1050.n0 173.2
R756 a_1771_1050.n6 a_1771_1050.n1 153.043
R757 a_1771_1050.n8 a_1771_1050.n7 76.002
R758 a_1771_1050.n5 a_1771_1050.n4 30
R759 a_1771_1050.n3 a_1771_1050.n2 24.383
R760 a_1771_1050.n5 a_1771_1050.n3 23.684
R761 a_1771_1050.n7 a_1771_1050.t3 14.282
R762 a_1771_1050.n7 a_1771_1050.t4 14.282
R763 a_1771_1050.t1 a_1771_1050.n9 14.282
R764 a_1771_1050.n9 a_1771_1050.t0 14.282
R765 a_1771_1050.n9 a_1771_1050.n8 12.848
R766 a_2405_209.n0 a_2405_209.t3 470.752
R767 a_2405_209.n0 a_2405_209.t5 384.527
R768 a_2405_209.n1 a_2405_209.t4 267.725
R769 a_2405_209.n3 a_2405_209.n2 253.86
R770 a_2405_209.n3 a_2405_209.n1 156.307
R771 a_2405_209.n4 a_2405_209.n3 130.9
R772 a_2405_209.n1 a_2405_209.n0 83.62
R773 a_2405_209.t1 a_2405_209.n4 14.282
R774 a_2405_209.n4 a_2405_209.t0 14.282
R775 a_3007_411.n0 a_3007_411.t6 470.752
R776 a_3007_411.n0 a_3007_411.t4 384.527
R777 a_3007_411.n1 a_3007_411.t5 241.172
R778 a_3007_411.n8 a_3007_411.n7 165.335
R779 a_3007_411.n7 a_3007_411.n6 162.187
R780 a_3007_411.n7 a_3007_411.n1 154.947
R781 a_3007_411.n6 a_3007_411.n5 133.539
R782 a_3007_411.n1 a_3007_411.n0 110.173
R783 a_3007_411.n6 a_3007_411.n2 70.262
R784 a_3007_411.n5 a_3007_411.n4 22.578
R785 a_3007_411.t2 a_3007_411.n8 14.282
R786 a_3007_411.n8 a_3007_411.t1 14.282
R787 a_3007_411.n5 a_3007_411.n3 8.58
R788 a_1666_101.t0 a_1666_101.n1 34.62
R789 a_1666_101.t0 a_1666_101.n0 8.137
R790 a_1666_101.t0 a_1666_101.n2 4.69
C4 VDD GND 15.72fF
C5 a_1666_101.n0 GND 0.05fF
C6 a_1666_101.n1 GND 0.12fF
C7 a_1666_101.n2 GND 0.04fF
C8 a_3007_411.n0 GND 0.38fF
C9 a_3007_411.n1 GND 0.84fF
C10 a_3007_411.n2 GND 0.21fF
C11 a_3007_411.n3 GND 0.05fF
C12 a_3007_411.n4 GND 0.06fF
C13 a_3007_411.n5 GND 0.21fF
C14 a_3007_411.n6 GND 0.52fF
C15 a_3007_411.n7 GND 0.84fF
C16 a_3007_411.n8 GND 0.76fF
C17 a_2405_209.n0 GND 0.37fF
C18 a_2405_209.t4 GND 0.67fF
C19 a_2405_209.n1 GND 1.07fF
C20 a_2405_209.n2 GND 0.50fF
C21 a_2405_209.n3 GND 1.18fF
C22 a_2405_209.n4 GND 0.83fF
C23 a_1771_1050.n0 GND 0.33fF
C24 a_1771_1050.t7 GND 0.45fF
C25 a_1771_1050.n1 GND 0.51fF
C26 a_1771_1050.n2 GND 0.04fF
C27 a_1771_1050.n3 GND 0.05fF
C28 a_1771_1050.n4 GND 0.03fF
C29 a_1771_1050.n5 GND 0.24fF
C30 a_1771_1050.n6 GND 0.51fF
C31 a_1771_1050.n7 GND 0.55fF
C32 a_1771_1050.n8 GND 0.30fF
C33 a_1771_1050.n9 GND 0.47fF
C34 a_2795_1051.n0 GND 0.55fF
C35 a_1295_209.n0 GND 0.44fF
C36 a_1295_209.n1 GND 1.26fF
C37 a_1295_209.n2 GND 0.47fF
C38 a_1295_209.n3 GND 1.34fF
C39 a_1295_209.n4 GND 0.88fF
C40 a_661_1050.n0 GND 0.35fF
C41 a_661_1050.t6 GND 0.47fF
C42 a_661_1050.n1 GND 0.53fF
C43 a_661_1050.n2 GND 0.34fF
C44 a_661_1050.n3 GND 0.56fF
C45 a_661_1050.n4 GND 0.58fF
C46 a_661_1050.n5 GND 0.31fF
C47 a_661_1050.n6 GND 0.49fF
C48 a_556_101.n0 GND 0.05fF
C49 a_556_101.n1 GND 0.12fF
C50 a_556_101.n2 GND 0.04fF
C51 a_185_209.n0 GND 0.36fF
C52 a_185_209.n1 GND 0.55fF
C53 a_185_209.n2 GND 0.37fF
C54 a_185_209.n3 GND 0.62fF
C55 a_185_209.n4 GND 0.70fF
C56 a_3461_1051.n0 GND 0.52fF
C57 VDD.n0 GND 0.14fF
C58 VDD.n1 GND 0.02fF
C59 VDD.n2 GND 0.02fF
C60 VDD.n3 GND 0.04fF
C61 VDD.n4 GND 0.01fF
C62 VDD.n6 GND 0.02fF
C63 VDD.n7 GND 0.02fF
C64 VDD.n8 GND 0.02fF
C65 VDD.n9 GND 0.02fF
C66 VDD.n12 GND 0.02fF
C67 VDD.n14 GND 0.43fF
C68 VDD.n16 GND 0.03fF
C69 VDD.n17 GND 0.02fF
C70 VDD.n18 GND 0.02fF
C71 VDD.n19 GND 0.02fF
C72 VDD.n20 GND 0.03fF
C73 VDD.n21 GND 0.26fF
C74 VDD.n22 GND 0.02fF
C75 VDD.n23 GND 0.03fF
C76 VDD.n24 GND 0.26fF
C77 VDD.n25 GND 0.01fF
C78 VDD.n26 GND 0.28fF
C79 VDD.n27 GND 0.01fF
C80 VDD.n28 GND 0.02fF
C81 VDD.n29 GND 0.26fF
C82 VDD.n30 GND 0.01fF
C83 VDD.n31 GND 0.02fF
C84 VDD.n32 GND 0.02fF
C85 VDD.n33 GND 0.00fF
C86 VDD.n34 GND 0.08fF
C87 VDD.n35 GND 0.02fF
C88 VDD.n36 GND 0.16fF
C89 VDD.n37 GND 0.13fF
C90 VDD.n38 GND 0.01fF
C91 VDD.n39 GND 0.02fF
C92 VDD.n40 GND 0.02fF
C93 VDD.n41 GND 0.10fF
C94 VDD.n42 GND 0.02fF
C95 VDD.n43 GND 0.13fF
C96 VDD.n44 GND 0.15fF
C97 VDD.n45 GND 0.01fF
C98 VDD.n46 GND 0.02fF
C99 VDD.n47 GND 0.02fF
C100 VDD.n48 GND 0.23fF
C101 VDD.n49 GND 0.01fF
C102 VDD.n50 GND 0.02fF
C103 VDD.n51 GND 0.02fF
C104 VDD.n52 GND 0.26fF
C105 VDD.n53 GND 0.01fF
C106 VDD.n54 GND 0.02fF
C107 VDD.n55 GND 0.03fF
C108 VDD.n56 GND 0.02fF
C109 VDD.n57 GND 0.02fF
C110 VDD.n58 GND 0.02fF
C111 VDD.n59 GND 0.20fF
C112 VDD.n60 GND 0.04fF
C113 VDD.n61 GND 0.03fF
C114 VDD.n62 GND 0.02fF
C115 VDD.n64 GND 0.02fF
C116 VDD.n65 GND 0.02fF
C117 VDD.n66 GND 0.02fF
C118 VDD.n67 GND 0.02fF
C119 VDD.n69 GND 0.02fF
C120 VDD.n70 GND 0.02fF
C121 VDD.n71 GND 0.02fF
C122 VDD.n73 GND 0.26fF
C123 VDD.n75 GND 0.02fF
C124 VDD.n76 GND 0.02fF
C125 VDD.n77 GND 0.03fF
C126 VDD.n78 GND 0.02fF
C127 VDD.n79 GND 0.26fF
C128 VDD.n80 GND 0.01fF
C129 VDD.n81 GND 0.02fF
C130 VDD.n82 GND 0.03fF
C131 VDD.n83 GND 0.26fF
C132 VDD.n84 GND 0.01fF
C133 VDD.n85 GND 0.02fF
C134 VDD.n86 GND 0.02fF
C135 VDD.n87 GND 0.26fF
C136 VDD.n88 GND 0.01fF
C137 VDD.n89 GND 0.02fF
C138 VDD.n90 GND 0.02fF
C139 VDD.n91 GND 0.28fF
C140 VDD.n92 GND 0.01fF
C141 VDD.n93 GND 0.02fF
C142 VDD.n94 GND 0.02fF
C143 VDD.n95 GND 0.16fF
C144 VDD.n96 GND 0.13fF
C145 VDD.n97 GND 0.01fF
C146 VDD.n98 GND 0.02fF
C147 VDD.n99 GND 0.02fF
C148 VDD.n100 GND 0.10fF
C149 VDD.n101 GND 0.02fF
C150 VDD.n102 GND 0.13fF
C151 VDD.n103 GND 0.15fF
C152 VDD.n104 GND 0.01fF
C153 VDD.n105 GND 0.02fF
C154 VDD.n106 GND 0.02fF
C155 VDD.n107 GND 0.23fF
C156 VDD.n108 GND 0.01fF
C157 VDD.n109 GND 0.02fF
C158 VDD.n110 GND 0.02fF
C159 VDD.n111 GND 0.26fF
C160 VDD.n112 GND 0.01fF
C161 VDD.n113 GND 0.02fF
C162 VDD.n114 GND 0.03fF
C163 VDD.n115 GND 0.02fF
C164 VDD.n116 GND 0.02fF
C165 VDD.n117 GND 0.02fF
C166 VDD.n118 GND 0.17fF
C167 VDD.n119 GND 0.04fF
C168 VDD.n120 GND 0.03fF
C169 VDD.n121 GND 0.02fF
C170 VDD.n122 GND 0.02fF
C171 VDD.n123 GND 0.02fF
C172 VDD.n124 GND 0.02fF
C173 VDD.n125 GND 0.02fF
C174 VDD.n127 GND 0.02fF
C175 VDD.n128 GND 0.02fF
C176 VDD.n129 GND 0.02fF
C177 VDD.n131 GND 0.26fF
C178 VDD.n133 GND 0.02fF
C179 VDD.n134 GND 0.02fF
C180 VDD.n135 GND 0.03fF
C181 VDD.n136 GND 0.02fF
C182 VDD.n137 GND 0.26fF
C183 VDD.n138 GND 0.01fF
C184 VDD.n139 GND 0.02fF
C185 VDD.n140 GND 0.03fF
C186 VDD.n141 GND 0.06fF
C187 VDD.n142 GND 0.14fF
C188 VDD.n143 GND 0.19fF
C189 VDD.n144 GND 0.01fF
C190 VDD.n145 GND 0.01fF
C191 VDD.n146 GND 0.02fF
C192 VDD.n147 GND 0.16fF
C193 VDD.n148 GND 0.01fF
C194 VDD.n149 GND 0.02fF
C195 VDD.n150 GND 0.02fF
C196 VDD.n151 GND 0.14fF
C197 VDD.n152 GND 0.19fF
C198 VDD.n153 GND 0.01fF
C199 VDD.n154 GND 0.06fF
C200 VDD.n155 GND 0.01fF
C201 VDD.n156 GND 0.02fF
C202 VDD.n157 GND 0.26fF
C203 VDD.n158 GND 0.01fF
C204 VDD.n159 GND 0.02fF
C205 VDD.n160 GND 0.03fF
C206 VDD.n161 GND 0.02fF
C207 VDD.n162 GND 0.02fF
C208 VDD.n163 GND 0.02fF
C209 VDD.n164 GND 0.17fF
C210 VDD.n165 GND 0.04fF
C211 VDD.n166 GND 0.03fF
C212 VDD.n167 GND 0.02fF
C213 VDD.n168 GND 0.02fF
C214 VDD.n169 GND 0.02fF
C215 VDD.n170 GND 0.02fF
C216 VDD.n171 GND 0.02fF
C217 VDD.n173 GND 0.02fF
C218 VDD.n174 GND 0.02fF
C219 VDD.n175 GND 0.02fF
C220 VDD.n177 GND 0.26fF
C221 VDD.n179 GND 0.02fF
C222 VDD.n180 GND 0.02fF
C223 VDD.n181 GND 0.03fF
C224 VDD.n182 GND 0.02fF
C225 VDD.n183 GND 0.26fF
C226 VDD.n184 GND 0.01fF
C227 VDD.n185 GND 0.02fF
C228 VDD.n186 GND 0.03fF
C229 VDD.n187 GND 0.05fF
C230 VDD.n188 GND 0.23fF
C231 VDD.n189 GND 0.01fF
C232 VDD.n190 GND 0.01fF
C233 VDD.n191 GND 0.02fF
C234 VDD.n192 GND 0.13fF
C235 VDD.n193 GND 0.16fF
C236 VDD.n194 GND 0.01fF
C237 VDD.n195 GND 0.02fF
C238 VDD.n196 GND 0.01fF
C239 VDD.n197 GND 0.02fF
C240 VDD.n198 GND 0.02fF
C241 VDD.n199 GND 0.02fF
C242 VDD.n200 GND 0.11fF
C243 VDD.n201 GND 0.03fF
C244 VDD.n202 GND 0.02fF
C245 VDD.n203 GND 0.02fF
C246 VDD.n204 GND 0.02fF
C247 VDD.n205 GND 0.02fF
C248 VDD.n206 GND 0.02fF
C249 VDD.n208 GND 0.02fF
C250 VDD.n209 GND 0.02fF
C251 VDD.n210 GND 0.02fF
C252 VDD.n212 GND 0.43fF
C253 VDD.n214 GND 0.03fF
C254 VDD.n215 GND 0.03fF
C255 VDD.n216 GND 0.26fF
C256 VDD.n217 GND 0.02fF
C257 VDD.n218 GND 0.03fF
C258 VDD.n219 GND 0.03fF
C259 VDD.n220 GND 0.14fF
C260 VDD.n221 GND 0.19fF
C261 VDD.n222 GND 0.01fF
C262 VDD.n223 GND 0.06fF
C263 VDD.n224 GND 0.01fF
C264 VDD.n225 GND 0.02fF
C265 VDD.n226 GND 0.16fF
C266 VDD.n227 GND 0.01fF
C267 VDD.n228 GND 0.02fF
C268 VDD.n229 GND 0.02fF
C269 VDD.n230 GND 0.06fF
C270 VDD.n231 GND 0.14fF
C271 VDD.n232 GND 0.19fF
C272 VDD.n233 GND 0.01fF
C273 VDD.n234 GND 0.01fF
C274 VDD.n235 GND 0.02fF
C275 VDD.n236 GND 0.26fF
C276 VDD.n237 GND 0.01fF
C277 VDD.n238 GND 0.02fF
C278 VDD.n239 GND 0.03fF
C279 VDD.n240 GND 0.02fF
C280 VDD.n241 GND 0.26fF
C281 VDD.n242 GND 0.01fF
C282 VDD.n243 GND 0.02fF
C283 VDD.n244 GND 0.02fF
C284 VDD.n245 GND 0.02fF
C285 VDD.n246 GND 0.02fF
C286 VDD.n247 GND 0.02fF
C287 VDD.n248 GND 0.02fF
C288 VDD.n250 GND 0.02fF
C289 VDD.n251 GND 0.02fF
C290 VDD.n252 GND 0.02fF
C291 VDD.n253 GND 0.02fF
C292 VDD.n255 GND 0.03fF
C293 VDD.n256 GND 0.02fF
C294 VDD.n257 GND 0.17fF
C295 VDD.n258 GND 0.04fF
C296 VDD.n260 GND 0.26fF
C297 VDD.n262 GND 0.02fF
C298 VDD.n263 GND 0.02fF
C299 VDD.n264 GND 0.03fF
C300 VDD.n265 GND 0.02fF
C301 VDD.n266 GND 0.03fF
C302 VDD.n267 GND 0.06fF
C303 VDD.n268 GND 0.23fF
C304 VDD.n269 GND 0.01fF
C305 VDD.n270 GND 0.01fF
C306 VDD.n271 GND 0.02fF
C307 VDD.n272 GND 0.13fF
C308 VDD.n273 GND 0.15fF
C309 VDD.n274 GND 0.01fF
C310 VDD.n275 GND 0.02fF
C311 VDD.n276 GND 0.02fF
C312 VDD.n277 GND 0.16fF
C313 VDD.n278 GND 0.13fF
C314 VDD.n279 GND 0.01fF
C315 VDD.n280 GND 0.02fF
C316 VDD.n281 GND 0.02fF
C317 VDD.n282 GND 0.28fF
C318 VDD.n283 GND 0.01fF
C319 VDD.n284 GND 0.10fF
C320 VDD.n285 GND 0.02fF
C321 VDD.n286 GND 0.02fF
C322 VDD.n287 GND 0.02fF
C323 VDD.n288 GND 0.13fF
C324 VDD.n289 GND 0.16fF
C325 VDD.n290 GND 0.01fF
C326 VDD.n291 GND 0.02fF
C327 VDD.n292 GND 0.02fF
C328 VDD.n293 GND 0.23fF
C329 VDD.n294 GND 0.01fF
C330 VDD.n295 GND 0.05fF
C331 VDD.n296 GND 0.01fF
C332 VDD.n297 GND 0.02fF
C333 VDD.n298 GND 0.26fF
C334 VDD.n299 GND 0.01fF
C335 VDD.n300 GND 0.02fF
C336 VDD.n301 GND 0.03fF
C337 VDD.n302 GND 0.02fF
C338 VDD.n303 GND 0.26fF
C339 VDD.n304 GND 0.01fF
C340 VDD.n305 GND 0.02fF
C341 VDD.n306 GND 0.02fF
C342 VDD.n307 GND 0.02fF
C343 VDD.n308 GND 0.17fF
C344 VDD.n309 GND 0.04fF
C345 VDD.n310 GND 0.03fF
C346 VDD.n311 GND 0.02fF
C347 VDD.n312 GND 0.02fF
C348 VDD.n313 GND 0.02fF
C349 VDD.n314 GND 0.02fF
C350 VDD.n315 GND 0.02fF
C351 VDD.n317 GND 0.02fF
C352 VDD.n318 GND 0.02fF
C353 VDD.n319 GND 0.02fF
C354 VDD.n321 GND 0.26fF
C355 VDD.n323 GND 0.02fF
C356 VDD.n324 GND 0.02fF
C357 VDD.n325 GND 0.03fF
C358 VDD.n326 GND 0.02fF
C359 VDD.n327 GND 0.03fF
C360 VDD.n328 GND 0.06fF
C361 VDD.n329 GND 0.14fF
C362 VDD.n330 GND 0.19fF
C363 VDD.n331 GND 0.01fF
C364 VDD.n332 GND 0.01fF
C365 VDD.n333 GND 0.02fF
C366 VDD.n334 GND 0.16fF
C367 VDD.n335 GND 0.01fF
C368 VDD.n336 GND 0.02fF
C369 VDD.n337 GND 0.02fF
C370 VDD.n338 GND 0.06fF
C371 VDD.n339 GND 0.14fF
C372 VDD.n340 GND 0.19fF
C373 VDD.n341 GND 0.01fF
C374 VDD.n342 GND 0.01fF
C375 VDD.n343 GND 0.02fF
C376 VDD.n344 GND 0.26fF
C377 VDD.n345 GND 0.01fF
C378 VDD.n346 GND 0.02fF
C379 VDD.n347 GND 0.03fF
C380 VDD.n348 GND 0.02fF
C381 VDD.n349 GND 0.02fF
C382 VDD.n350 GND 0.02fF
C383 VDD.n351 GND 0.17fF
C384 VDD.n352 GND 0.04fF
C385 VDD.n353 GND 0.03fF
C386 VDD.n354 GND 0.02fF
C387 VDD.n355 GND 0.02fF
C388 VDD.n356 GND 0.02fF
C389 VDD.n357 GND 0.02fF
C390 VDD.n358 GND 0.02fF
C391 VDD.n360 GND 0.02fF
C392 VDD.n361 GND 0.02fF
C393 VDD.n362 GND 0.02fF
C394 VDD.n364 GND 0.26fF
C395 VDD.n366 GND 0.02fF
C396 VDD.n367 GND 0.02fF
C397 VDD.n368 GND 0.03fF
C398 VDD.n369 GND 0.02fF
C399 VDD.n370 GND 0.26fF
C400 VDD.n371 GND 0.01fF
C401 VDD.n372 GND 0.02fF
C402 VDD.n373 GND 0.03fF
C403 VDD.n374 GND 0.06fF
C404 VDD.n375 GND 0.23fF
C405 VDD.n376 GND 0.01fF
C406 VDD.n377 GND 0.01fF
C407 VDD.n378 GND 0.02fF
C408 VDD.n379 GND 0.13fF
C409 VDD.n380 GND 0.15fF
C410 VDD.n381 GND 0.01fF
C411 VDD.n382 GND 0.02fF
C412 VDD.n383 GND 0.02fF
C413 VDD.n384 GND 0.16fF
C414 VDD.n385 GND 0.13fF
C415 VDD.n386 GND 0.01fF
C416 VDD.n387 GND 0.02fF
C417 VDD.n388 GND 0.02fF
C418 VDD.n389 GND 0.10fF
C419 VDD.n390 GND 0.02fF
C420 VDD.n391 GND 0.28fF
C421 VDD.n392 GND 0.01fF
C422 VDD.n393 GND 0.02fF
C423 VDD.n394 GND 0.02fF
C424 Q.n0 GND 0.40fF
C425 Q.t5 GND 0.52fF
C426 Q.n1 GND 0.41fF
C427 Q.n2 GND 0.72fF
C428 Q.n3 GND 0.06fF
C429 Q.n4 GND 0.04fF
C430 Q.n5 GND 0.13fF
C431 Q.n6 GND 0.04fF
C432 Q.n7 GND 0.06fF
C433 Q.n8 GND 0.04fF
C434 Q.n9 GND 0.19fF
C435 Q.n10 GND 0.37fF
C436 Q.n11 GND 0.39fF
C437 Q.n12 GND 0.35fF
.ends
