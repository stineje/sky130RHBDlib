magic
tech sky130A
magscale 1 2
timestamp 1652368010
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 1167 945 1201 979
rect 205 871 239 905
rect 353 871 387 905
rect 1019 871 1053 905
rect 1167 871 1201 905
rect 205 797 239 831
rect 353 797 387 831
rect 1019 797 1053 831
rect 1167 797 1201 831
rect 205 723 239 757
rect 353 723 387 757
rect 1019 723 1053 757
rect 1167 723 1201 757
rect 205 649 239 683
rect 353 649 387 683
rect 1019 649 1053 683
rect 1167 649 1201 683
rect 205 575 239 609
rect 353 575 387 609
rect 1019 575 1053 609
rect 1167 575 1201 609
rect 205 501 239 535
rect 353 501 387 535
rect 1019 501 1053 535
rect 1167 501 1201 535
rect 205 427 239 461
rect 353 427 387 461
rect 1019 427 1053 461
rect 1167 427 1201 461
<< metal1 >>
rect -34 1446 1366 1514
rect -34 -34 1366 34
use aoi3x1_pcell  aoi3x1_pcell_0 pcells
timestamp 1652367586
transform 1 0 0 0 1 0
box -87 -34 1419 1550
<< labels >>
rlabel locali 1167 797 1201 831 1 YN
port 1 nsew signal output
rlabel locali 1167 723 1201 757 1 YN
port 1 nsew signal output
rlabel locali 1167 649 1201 683 1 YN
port 1 nsew signal output
rlabel locali 1167 575 1201 609 1 YN
port 1 nsew signal output
rlabel locali 1167 501 1201 535 1 YN
port 1 nsew signal output
rlabel locali 1167 427 1201 461 1 YN
port 1 nsew signal output
rlabel locali 1167 871 1201 905 1 YN
port 1 nsew signal output
rlabel locali 1167 945 1201 979 1 YN
port 1 nsew signal output
rlabel locali 205 575 239 609 1 A
port 2 nsew signal input
rlabel locali 205 501 239 535 1 A
port 2 nsew signal input
rlabel locali 205 427 239 461 1 A
port 2 nsew signal input
rlabel locali 205 649 239 683 1 A
port 2 nsew signal input
rlabel locali 205 723 239 757 1 A
port 2 nsew signal input
rlabel locali 205 797 239 831 1 A
port 2 nsew signal input
rlabel locali 205 871 239 905 1 A
port 2 nsew signal input
rlabel locali 353 649 387 683 1 B
port 3 nsew signal input
rlabel locali 353 575 387 609 1 B
port 3 nsew signal input
rlabel locali 353 501 387 535 1 B
port 3 nsew signal input
rlabel locali 353 427 387 461 1 B
port 3 nsew signal input
rlabel locali 353 723 387 757 1 B
port 3 nsew signal input
rlabel locali 353 797 387 831 1 B
port 3 nsew signal input
rlabel locali 353 871 387 905 1 B
port 3 nsew signal input
rlabel locali 1019 723 1053 757 1 C
port 4 nsew signal input
rlabel locali 1019 649 1053 683 1 C
port 4 nsew signal input
rlabel locali 1019 575 1053 609 1 C
port 4 nsew signal input
rlabel locali 1019 501 1053 535 1 C
port 4 nsew signal input
rlabel locali 1019 427 1053 461 1 C
port 4 nsew signal input
rlabel locali 1019 797 1053 831 1 C
port 4 nsew signal input
rlabel locali 1019 871 1053 905 1 C
port 4 nsew signal input
rlabel metal1 -34 1446 1366 1514 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 -34 -34 1366 34 1 VGND
port 6 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
port 7 nsew power bidirectional
rlabel pwell 57 -17 91 17 1 VNB
port 8 nsew ground bidirectional
<< properties >>
string LEFsite unithd 
string LEFclass CORE
string FIXED_BBOX 0 0 1332 1480
string LEFsymmetry X Y R90
<< end >>
